module basic_3000_30000_3500_50_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_2203,In_1769);
nand U1 (N_1,In_559,In_1744);
nand U2 (N_2,In_1978,In_1847);
and U3 (N_3,In_733,In_1008);
nor U4 (N_4,In_866,In_18);
xor U5 (N_5,In_1324,In_2063);
xor U6 (N_6,In_2765,In_1401);
nor U7 (N_7,In_1791,In_1384);
nand U8 (N_8,In_423,In_2805);
nand U9 (N_9,In_381,In_269);
or U10 (N_10,In_2755,In_2249);
xnor U11 (N_11,In_651,In_2713);
or U12 (N_12,In_2547,In_263);
nand U13 (N_13,In_1241,In_2836);
and U14 (N_14,In_1131,In_2325);
nor U15 (N_15,In_2436,In_2433);
and U16 (N_16,In_1629,In_1496);
and U17 (N_17,In_1754,In_56);
nor U18 (N_18,In_2988,In_1371);
and U19 (N_19,In_1759,In_189);
and U20 (N_20,In_1670,In_97);
nor U21 (N_21,In_642,In_1739);
or U22 (N_22,In_1969,In_1273);
nor U23 (N_23,In_2862,In_2802);
nor U24 (N_24,In_1330,In_873);
and U25 (N_25,In_336,In_943);
xnor U26 (N_26,In_784,In_1710);
xor U27 (N_27,In_1351,In_57);
or U28 (N_28,In_329,In_1962);
and U29 (N_29,In_1173,In_2303);
xnor U30 (N_30,In_1081,In_2048);
and U31 (N_31,In_2621,In_2894);
nor U32 (N_32,In_1362,In_1167);
xor U33 (N_33,In_1446,In_2425);
or U34 (N_34,In_2013,In_1249);
nor U35 (N_35,In_2105,In_2980);
nor U36 (N_36,In_2218,In_1442);
or U37 (N_37,In_2563,In_193);
nand U38 (N_38,In_272,In_2932);
nand U39 (N_39,In_928,In_506);
and U40 (N_40,In_2523,In_448);
or U41 (N_41,In_1376,In_2597);
xnor U42 (N_42,In_2617,In_2642);
or U43 (N_43,In_509,In_71);
and U44 (N_44,In_4,In_2648);
or U45 (N_45,In_656,In_2993);
nor U46 (N_46,In_229,In_1325);
xor U47 (N_47,In_1368,In_1252);
or U48 (N_48,In_2396,In_195);
and U49 (N_49,In_1530,In_2801);
nand U50 (N_50,In_2797,In_275);
nand U51 (N_51,In_2776,In_863);
and U52 (N_52,In_1660,In_2364);
and U53 (N_53,In_909,In_1303);
and U54 (N_54,In_2450,In_1187);
nor U55 (N_55,In_629,In_1728);
nand U56 (N_56,In_1579,In_2904);
and U57 (N_57,In_1094,In_1863);
and U58 (N_58,In_201,In_1925);
and U59 (N_59,In_988,In_1464);
or U60 (N_60,In_242,In_2674);
and U61 (N_61,In_2457,In_2629);
nor U62 (N_62,In_2769,In_780);
nand U63 (N_63,In_1284,In_2726);
or U64 (N_64,In_2572,In_1866);
and U65 (N_65,In_23,In_1926);
or U66 (N_66,In_1421,In_527);
and U67 (N_67,In_1603,In_1913);
or U68 (N_68,In_2934,In_1043);
and U69 (N_69,In_2069,In_2535);
nand U70 (N_70,In_2373,In_589);
and U71 (N_71,In_816,In_2778);
and U72 (N_72,In_1321,In_2790);
or U73 (N_73,In_1526,In_2973);
xor U74 (N_74,In_1286,In_855);
and U75 (N_75,In_751,In_402);
nand U76 (N_76,In_1860,In_2443);
or U77 (N_77,In_406,In_662);
nand U78 (N_78,In_373,In_1139);
nand U79 (N_79,In_2235,In_2933);
nand U80 (N_80,In_2789,In_566);
or U81 (N_81,In_1200,In_148);
nor U82 (N_82,In_2258,In_2709);
or U83 (N_83,In_1373,In_2500);
and U84 (N_84,In_1428,In_1084);
nor U85 (N_85,In_2925,In_1968);
nand U86 (N_86,In_2283,In_2634);
and U87 (N_87,In_1515,In_1476);
nor U88 (N_88,In_1695,In_1118);
or U89 (N_89,In_2981,In_2109);
xor U90 (N_90,In_1647,In_531);
nor U91 (N_91,In_1210,In_1452);
xor U92 (N_92,In_849,In_996);
and U93 (N_93,In_690,In_142);
or U94 (N_94,In_2407,In_1291);
nand U95 (N_95,In_2897,In_676);
and U96 (N_96,In_515,In_796);
and U97 (N_97,In_1233,In_2290);
and U98 (N_98,In_2170,In_1702);
xor U99 (N_99,In_2078,In_1733);
or U100 (N_100,In_1840,In_2151);
or U101 (N_101,In_1630,In_699);
nor U102 (N_102,In_1290,In_2045);
and U103 (N_103,In_310,In_2846);
and U104 (N_104,In_1775,In_1671);
nand U105 (N_105,In_538,In_1998);
nor U106 (N_106,In_2628,In_2887);
and U107 (N_107,In_313,In_115);
nor U108 (N_108,In_903,In_259);
nor U109 (N_109,In_2056,In_556);
xnor U110 (N_110,In_2935,In_1585);
nor U111 (N_111,In_303,In_1708);
nor U112 (N_112,In_2287,In_2633);
xnor U113 (N_113,In_746,In_2301);
nand U114 (N_114,In_1937,In_1942);
and U115 (N_115,In_1137,In_670);
nor U116 (N_116,In_547,In_404);
and U117 (N_117,In_2233,In_1314);
and U118 (N_118,In_1181,In_990);
and U119 (N_119,In_697,In_1757);
and U120 (N_120,In_2066,In_1356);
nor U121 (N_121,In_1172,In_742);
and U122 (N_122,In_447,In_757);
nand U123 (N_123,In_2391,In_822);
nor U124 (N_124,In_1419,In_2576);
or U125 (N_125,In_1358,In_879);
and U126 (N_126,In_2559,In_1954);
nor U127 (N_127,In_1313,In_2650);
xnor U128 (N_128,In_2867,In_720);
nand U129 (N_129,In_2509,In_2031);
and U130 (N_130,In_1537,In_162);
or U131 (N_131,In_1005,In_557);
and U132 (N_132,In_2546,In_2859);
nand U133 (N_133,In_2575,In_984);
or U134 (N_134,In_734,In_518);
or U135 (N_135,In_1960,In_100);
nand U136 (N_136,In_2868,In_1275);
xor U137 (N_137,In_1653,In_838);
nor U138 (N_138,In_210,In_410);
xnor U139 (N_139,In_1492,In_1527);
and U140 (N_140,In_633,In_440);
nand U141 (N_141,In_1044,In_2794);
and U142 (N_142,In_706,In_2445);
nand U143 (N_143,In_801,In_2505);
nor U144 (N_144,In_2260,In_962);
xnor U145 (N_145,In_109,In_2842);
nor U146 (N_146,In_2912,In_431);
nor U147 (N_147,In_257,In_181);
nor U148 (N_148,In_524,In_326);
nor U149 (N_149,In_1422,In_491);
nor U150 (N_150,In_1773,In_624);
nand U151 (N_151,In_1332,In_1144);
and U152 (N_152,In_1142,In_2543);
xnor U153 (N_153,In_2222,In_1593);
and U154 (N_154,In_537,In_2210);
nand U155 (N_155,In_944,In_282);
or U156 (N_156,In_1209,In_1873);
xnor U157 (N_157,In_2390,In_2308);
and U158 (N_158,In_1770,In_2696);
and U159 (N_159,In_1675,In_2580);
xnor U160 (N_160,In_2122,In_2267);
and U161 (N_161,In_2285,In_2357);
nand U162 (N_162,In_1923,In_1551);
nand U163 (N_163,In_654,In_1498);
or U164 (N_164,In_335,In_1990);
nand U165 (N_165,In_439,In_2092);
nor U166 (N_166,In_896,In_2984);
xor U167 (N_167,In_1891,In_835);
and U168 (N_168,In_1575,In_1615);
and U169 (N_169,In_2051,In_1731);
or U170 (N_170,In_1192,In_2649);
or U171 (N_171,In_991,In_1541);
nor U172 (N_172,In_1590,In_1656);
nor U173 (N_173,In_252,In_542);
or U174 (N_174,In_828,In_2964);
nand U175 (N_175,In_1672,In_1935);
nor U176 (N_176,In_1658,In_316);
or U177 (N_177,In_1936,In_2786);
and U178 (N_178,In_1871,In_1879);
xor U179 (N_179,In_2998,In_2146);
xnor U180 (N_180,In_2018,In_488);
nand U181 (N_181,In_2558,In_1634);
xor U182 (N_182,In_372,In_2888);
or U183 (N_183,In_407,In_1331);
nor U184 (N_184,In_1440,In_2625);
and U185 (N_185,In_1279,In_2100);
xor U186 (N_186,In_2476,In_1943);
nand U187 (N_187,In_1402,In_2914);
or U188 (N_188,In_236,In_17);
nor U189 (N_189,In_867,In_1159);
nor U190 (N_190,In_1269,In_921);
nor U191 (N_191,In_543,In_914);
nor U192 (N_192,In_1763,In_1430);
xor U193 (N_193,In_1302,In_2253);
and U194 (N_194,In_186,In_358);
and U195 (N_195,In_2931,In_2594);
nand U196 (N_196,In_1438,In_2004);
nand U197 (N_197,In_2719,In_2216);
xnor U198 (N_198,In_1189,In_2480);
and U199 (N_199,In_1804,In_2118);
and U200 (N_200,In_191,In_323);
xnor U201 (N_201,In_1857,In_113);
nand U202 (N_202,In_1184,In_179);
nor U203 (N_203,In_992,In_99);
nand U204 (N_204,In_1480,In_738);
xnor U205 (N_205,In_1353,In_964);
xnor U206 (N_206,In_1563,In_1628);
nand U207 (N_207,In_1649,In_360);
or U208 (N_208,In_1031,In_721);
xor U209 (N_209,In_1623,In_2568);
or U210 (N_210,In_2818,In_2102);
nor U211 (N_211,In_615,In_1329);
xor U212 (N_212,In_1732,In_1003);
or U213 (N_213,In_1281,In_998);
nor U214 (N_214,In_2624,In_2660);
nor U215 (N_215,In_603,In_2025);
xnor U216 (N_216,In_2783,In_672);
or U217 (N_217,In_701,In_1668);
xnor U218 (N_218,In_2215,In_52);
nor U219 (N_219,In_1357,In_2471);
and U220 (N_220,In_1705,In_1424);
nand U221 (N_221,In_813,In_1012);
xor U222 (N_222,In_1613,In_541);
xnor U223 (N_223,In_379,In_985);
nand U224 (N_224,In_1479,In_2915);
nor U225 (N_225,In_212,In_1457);
nor U226 (N_226,In_2908,In_2661);
nor U227 (N_227,In_2645,In_2652);
nor U228 (N_228,In_1529,In_2923);
or U229 (N_229,In_1956,In_963);
nor U230 (N_230,In_2737,In_1576);
and U231 (N_231,In_2464,In_333);
and U232 (N_232,In_1963,In_295);
and U233 (N_233,In_2111,In_2144);
or U234 (N_234,In_1341,In_470);
nand U235 (N_235,In_646,In_832);
nand U236 (N_236,In_1343,In_1449);
nand U237 (N_237,In_932,In_1587);
nor U238 (N_238,In_2507,In_1214);
or U239 (N_239,In_869,In_2533);
or U240 (N_240,In_2237,In_735);
nand U241 (N_241,In_254,In_1676);
nor U242 (N_242,In_1699,In_1450);
nand U243 (N_243,In_599,In_2120);
or U244 (N_244,In_1704,In_519);
nand U245 (N_245,In_1104,In_2609);
or U246 (N_246,In_1972,In_839);
nor U247 (N_247,In_123,In_1627);
and U248 (N_248,In_1869,In_2835);
nor U249 (N_249,In_1392,In_1101);
and U250 (N_250,In_724,In_745);
xnor U251 (N_251,In_2740,In_593);
xnor U252 (N_252,In_2968,In_298);
and U253 (N_253,In_1123,In_1100);
nor U254 (N_254,In_2861,In_2462);
nor U255 (N_255,In_552,In_1196);
xnor U256 (N_256,In_2446,In_1298);
nor U257 (N_257,In_2618,In_2343);
xor U258 (N_258,In_2011,In_851);
or U259 (N_259,In_1097,In_1390);
nand U260 (N_260,In_80,In_2340);
and U261 (N_261,In_1211,In_394);
and U262 (N_262,In_1681,In_1523);
xnor U263 (N_263,In_2427,In_1218);
xor U264 (N_264,In_2775,In_1046);
xnor U265 (N_265,In_564,In_2402);
nor U266 (N_266,In_2898,In_235);
xor U267 (N_267,In_571,In_1320);
nor U268 (N_268,In_390,In_622);
xnor U269 (N_269,In_3,In_956);
nand U270 (N_270,In_1415,In_772);
and U271 (N_271,In_1145,In_1793);
nor U272 (N_272,In_1098,In_2161);
nor U273 (N_273,In_340,In_2355);
nor U274 (N_274,In_2224,In_2948);
and U275 (N_275,In_74,In_224);
or U276 (N_276,In_213,In_1489);
xnor U277 (N_277,In_583,In_590);
nand U278 (N_278,In_717,In_2635);
or U279 (N_279,In_199,In_732);
or U280 (N_280,In_1338,In_2536);
or U281 (N_281,In_2125,In_1058);
and U282 (N_282,In_1874,In_411);
nand U283 (N_283,In_675,In_2376);
or U284 (N_284,In_1156,In_1441);
and U285 (N_285,In_2566,In_1451);
xnor U286 (N_286,In_1893,In_467);
nor U287 (N_287,In_819,In_1038);
nand U288 (N_288,In_1293,In_689);
nor U289 (N_289,In_2959,In_1643);
xor U290 (N_290,In_2095,In_1557);
and U291 (N_291,In_1531,In_1999);
and U292 (N_292,In_1133,In_405);
and U293 (N_293,In_2155,In_2971);
or U294 (N_294,In_1635,In_1034);
and U295 (N_295,In_60,In_759);
xor U296 (N_296,In_792,In_2238);
or U297 (N_297,In_1730,In_1856);
nand U298 (N_298,In_793,In_1517);
xor U299 (N_299,In_1177,In_2515);
nand U300 (N_300,In_1746,In_2531);
xnor U301 (N_301,In_1141,In_1818);
and U302 (N_302,In_1932,In_32);
or U303 (N_303,In_1345,In_2681);
xor U304 (N_304,In_51,In_1251);
nand U305 (N_305,In_1577,In_262);
nand U306 (N_306,In_1807,In_249);
nand U307 (N_307,In_73,In_817);
and U308 (N_308,In_2949,In_856);
nor U309 (N_309,In_2437,In_1947);
nor U310 (N_310,In_219,In_1700);
or U311 (N_311,In_637,In_1955);
xor U312 (N_312,In_1662,In_355);
or U313 (N_313,In_584,In_946);
or U314 (N_314,In_2322,In_2207);
xnor U315 (N_315,In_216,In_1598);
nand U316 (N_316,In_172,In_2941);
nor U317 (N_317,In_2495,In_471);
and U318 (N_318,In_2479,In_1912);
xor U319 (N_319,In_1090,In_1347);
and U320 (N_320,In_2008,In_1544);
and U321 (N_321,In_854,In_2229);
nand U322 (N_322,In_299,In_1789);
nand U323 (N_323,In_1154,In_221);
nor U324 (N_324,In_2358,In_465);
nor U325 (N_325,In_605,In_1771);
xnor U326 (N_326,In_2148,In_608);
and U327 (N_327,In_1261,In_444);
nor U328 (N_328,In_1911,In_2254);
nor U329 (N_329,In_2691,In_2418);
nor U330 (N_330,In_2873,In_2721);
or U331 (N_331,In_2664,In_1245);
xnor U332 (N_332,In_886,In_2542);
or U333 (N_333,In_1827,In_1205);
or U334 (N_334,In_2979,In_1334);
nor U335 (N_335,In_1319,In_2697);
nor U336 (N_336,In_1478,In_743);
nand U337 (N_337,In_680,In_1738);
nor U338 (N_338,In_141,In_2110);
nor U339 (N_339,In_818,In_2820);
and U340 (N_340,In_1217,In_1207);
xnor U341 (N_341,In_1375,In_2675);
xnor U342 (N_342,In_321,In_125);
or U343 (N_343,In_460,In_2796);
nor U344 (N_344,In_2647,In_151);
or U345 (N_345,In_1372,In_2885);
nor U346 (N_346,In_1640,In_415);
xor U347 (N_347,In_2298,In_2430);
and U348 (N_348,In_2766,In_2974);
or U349 (N_349,In_43,In_449);
or U350 (N_350,In_1872,In_691);
and U351 (N_351,In_1393,In_859);
xnor U352 (N_352,In_2180,In_764);
or U353 (N_353,In_261,In_107);
or U354 (N_354,In_647,In_2599);
xor U355 (N_355,In_1201,In_2217);
nor U356 (N_356,In_2382,In_558);
and U357 (N_357,In_2982,In_1895);
and U358 (N_358,In_2545,In_2651);
nand U359 (N_359,In_1745,In_2787);
nor U360 (N_360,In_2880,In_1243);
or U361 (N_361,In_2265,In_2379);
xnor U362 (N_362,In_145,In_744);
nand U363 (N_363,In_429,In_2779);
nor U364 (N_364,In_2274,In_2057);
and U365 (N_365,In_1836,In_2150);
xnor U366 (N_366,In_1503,In_1621);
and U367 (N_367,In_1001,In_2960);
or U368 (N_368,In_918,In_1564);
nand U369 (N_369,In_2690,In_89);
and U370 (N_370,In_1089,In_1318);
nand U371 (N_371,In_2774,In_563);
and U372 (N_372,In_1395,In_1583);
and U373 (N_373,In_1722,In_521);
nor U374 (N_374,In_1230,In_174);
nor U375 (N_375,In_2606,In_1425);
nand U376 (N_376,In_1981,In_2183);
and U377 (N_377,In_1801,In_993);
nor U378 (N_378,In_1204,In_1432);
or U379 (N_379,In_177,In_2473);
nand U380 (N_380,In_1514,In_2415);
and U381 (N_381,In_2331,In_2380);
and U382 (N_382,In_975,In_2315);
nand U383 (N_383,In_2307,In_2101);
and U384 (N_384,In_2913,In_951);
nand U385 (N_385,In_905,In_1021);
nand U386 (N_386,In_8,In_1483);
xor U387 (N_387,In_1830,In_1941);
xnor U388 (N_388,In_731,In_2646);
nor U389 (N_389,In_2608,In_858);
nand U390 (N_390,In_476,In_445);
nor U391 (N_391,In_1380,In_752);
and U392 (N_392,In_1032,In_2834);
xor U393 (N_393,In_1158,In_2833);
nand U394 (N_394,In_1661,In_91);
nand U395 (N_395,In_658,In_1108);
xor U396 (N_396,In_2865,In_2196);
nor U397 (N_397,In_2347,In_528);
and U398 (N_398,In_2052,In_237);
or U399 (N_399,In_1533,In_1413);
and U400 (N_400,In_226,In_2041);
nor U401 (N_401,In_1465,In_1988);
or U402 (N_402,In_2097,In_386);
nand U403 (N_403,In_1812,In_1007);
nor U404 (N_404,In_1993,In_2091);
and U405 (N_405,In_1572,In_376);
xnor U406 (N_406,In_2497,In_2541);
xnor U407 (N_407,In_778,In_2942);
nor U408 (N_408,In_718,In_1713);
xnor U409 (N_409,In_370,In_1914);
or U410 (N_410,In_81,In_2389);
nand U411 (N_411,In_325,In_1909);
or U412 (N_412,In_1582,In_2812);
and U413 (N_413,In_630,In_829);
and U414 (N_414,In_119,In_2455);
nand U415 (N_415,In_2975,In_915);
xor U416 (N_416,In_2070,In_1024);
nand U417 (N_417,In_1369,In_2561);
or U418 (N_418,In_1107,In_2593);
xor U419 (N_419,In_2604,In_875);
nand U420 (N_420,In_2967,In_1247);
nand U421 (N_421,In_1254,In_334);
xor U422 (N_422,In_320,In_1294);
nand U423 (N_423,In_904,In_2738);
xnor U424 (N_424,In_1880,In_980);
or U425 (N_425,In_188,In_950);
nand U426 (N_426,In_1176,In_2133);
nand U427 (N_427,In_1469,In_2813);
and U428 (N_428,In_2452,In_805);
nand U429 (N_429,In_1855,In_899);
and U430 (N_430,In_878,In_2901);
or U431 (N_431,In_636,In_957);
xnor U432 (N_432,In_2374,In_2702);
nor U433 (N_433,In_526,In_2037);
and U434 (N_434,In_2996,In_659);
or U435 (N_435,In_1885,In_2192);
or U436 (N_436,In_2295,In_1051);
xnor U437 (N_437,In_285,In_1074);
or U438 (N_438,In_2212,In_2969);
nor U439 (N_439,In_2746,In_2598);
xnor U440 (N_440,In_702,In_2854);
nor U441 (N_441,In_627,In_1690);
xnor U442 (N_442,In_1606,In_610);
and U443 (N_443,In_2548,In_695);
nand U444 (N_444,In_2165,In_536);
or U445 (N_445,In_1121,In_2485);
nor U446 (N_446,In_375,In_1397);
xor U447 (N_447,In_2911,In_1168);
xor U448 (N_448,In_22,In_322);
xor U449 (N_449,In_872,In_1971);
or U450 (N_450,In_1714,In_2451);
nor U451 (N_451,In_1350,In_1930);
xnor U452 (N_452,In_2716,In_218);
and U453 (N_453,In_1813,In_5);
xor U454 (N_454,In_47,In_1578);
nor U455 (N_455,In_368,In_437);
nand U456 (N_456,In_2026,In_880);
nor U457 (N_457,In_1877,In_1803);
and U458 (N_458,In_1625,In_979);
or U459 (N_459,In_1458,In_549);
or U460 (N_460,In_271,In_1228);
nand U461 (N_461,In_388,In_1974);
nand U462 (N_462,In_982,In_2190);
or U463 (N_463,In_1680,In_972);
xor U464 (N_464,In_2491,In_2459);
or U465 (N_465,In_729,In_2760);
xnor U466 (N_466,In_1760,In_1983);
or U467 (N_467,In_1898,In_312);
nor U468 (N_468,In_1786,In_1852);
nand U469 (N_469,In_2429,In_288);
and U470 (N_470,In_952,In_474);
xnor U471 (N_471,In_1427,In_1412);
or U472 (N_472,In_2613,In_280);
nor U473 (N_473,In_508,In_2856);
nand U474 (N_474,In_7,In_2089);
nand U475 (N_475,In_2722,In_902);
nand U476 (N_476,In_1067,In_2135);
xor U477 (N_477,In_1970,In_2119);
and U478 (N_478,In_2785,In_1928);
nor U479 (N_479,In_1042,In_2718);
nor U480 (N_480,In_573,In_1404);
and U481 (N_481,In_1921,In_2706);
and U482 (N_482,In_2910,In_2814);
nand U483 (N_483,In_2084,In_2220);
or U484 (N_484,In_722,In_2784);
and U485 (N_485,In_1654,In_2763);
and U486 (N_486,In_1054,In_1945);
nor U487 (N_487,In_926,In_2397);
xor U488 (N_488,In_1715,In_836);
xnor U489 (N_489,In_419,In_1648);
xor U490 (N_490,In_2073,In_2488);
and U491 (N_491,In_1407,In_2114);
or U492 (N_492,In_2866,In_1366);
nand U493 (N_493,In_1642,In_15);
xnor U494 (N_494,In_2845,In_591);
xnor U495 (N_495,In_2241,In_1619);
nand U496 (N_496,In_959,In_726);
xor U497 (N_497,In_2595,In_1940);
xor U498 (N_498,In_1655,In_233);
nand U499 (N_499,In_2023,In_569);
xnor U500 (N_500,In_1418,In_777);
or U501 (N_501,In_853,In_2244);
nand U502 (N_502,In_727,In_499);
xnor U503 (N_503,In_1231,In_912);
xnor U504 (N_504,In_1934,In_1596);
nand U505 (N_505,In_196,In_2248);
or U506 (N_506,In_2694,In_1272);
or U507 (N_507,In_2416,In_2519);
nor U508 (N_508,In_2257,In_2461);
and U509 (N_509,In_2824,In_791);
nand U510 (N_510,In_1454,In_2058);
xnor U511 (N_511,In_426,In_232);
or U512 (N_512,In_1865,In_924);
or U513 (N_513,In_1363,In_948);
and U514 (N_514,In_1087,In_2759);
and U515 (N_515,In_2731,In_2327);
and U516 (N_516,In_572,In_1161);
nand U517 (N_517,In_580,In_1336);
xnor U518 (N_518,In_1667,In_1811);
and U519 (N_519,In_1109,In_459);
or U520 (N_520,In_2588,In_997);
nand U521 (N_521,In_773,In_1501);
nand U522 (N_522,In_925,In_2349);
and U523 (N_523,In_922,In_652);
nand U524 (N_524,In_606,In_2113);
and U525 (N_525,In_683,In_432);
xnor U526 (N_526,In_2284,In_2992);
and U527 (N_527,In_588,In_2074);
or U528 (N_528,In_2990,In_490);
and U529 (N_529,In_1323,In_2557);
and U530 (N_530,In_941,In_2922);
and U531 (N_531,In_2387,In_723);
and U532 (N_532,In_2838,In_1004);
and U533 (N_533,In_2001,In_2230);
or U534 (N_534,In_1041,In_545);
and U535 (N_535,In_1278,In_2370);
xnor U536 (N_536,In_1982,In_463);
and U537 (N_537,In_2619,In_2749);
nor U538 (N_538,In_2124,In_417);
nor U539 (N_539,In_2456,In_2369);
and U540 (N_540,In_894,In_428);
xnor U541 (N_541,In_2242,In_2453);
nor U542 (N_542,In_1767,In_1795);
nand U543 (N_543,In_1905,In_462);
nor U544 (N_544,In_2064,In_2399);
xor U545 (N_545,In_1453,In_1624);
or U546 (N_546,In_1062,In_2771);
xnor U547 (N_547,In_2361,In_1858);
xor U548 (N_548,In_1057,In_1536);
xor U549 (N_549,In_665,In_1691);
nand U550 (N_550,In_2121,In_1027);
xor U551 (N_551,In_754,In_577);
xor U552 (N_552,In_2999,In_1280);
nand U553 (N_553,In_2022,In_2252);
nand U554 (N_554,In_2677,In_703);
nand U555 (N_555,In_2486,In_1248);
nor U556 (N_556,In_1924,In_671);
nand U557 (N_557,In_2924,In_239);
or U558 (N_558,In_2837,In_2553);
nor U559 (N_559,In_2002,In_639);
nand U560 (N_560,In_2653,In_581);
nor U561 (N_561,In_681,In_2050);
xor U562 (N_562,In_1335,In_1790);
or U563 (N_563,In_30,In_1236);
nand U564 (N_564,In_1602,In_1066);
nor U565 (N_565,In_1721,In_908);
or U566 (N_566,In_436,In_1525);
xor U567 (N_567,In_1386,In_2293);
nand U568 (N_568,In_343,In_2080);
xor U569 (N_569,In_800,In_1882);
xnor U570 (N_570,In_385,In_2130);
or U571 (N_571,In_1305,In_483);
and U572 (N_572,In_2240,In_1841);
xnor U573 (N_573,In_1060,In_1562);
or U574 (N_574,In_2278,In_2075);
xor U575 (N_575,In_1977,In_167);
nor U576 (N_576,In_1806,In_736);
and U577 (N_577,In_967,In_2540);
and U578 (N_578,In_643,In_1796);
or U579 (N_579,In_396,In_2377);
or U580 (N_580,In_2388,In_594);
or U581 (N_581,In_2506,In_1995);
or U582 (N_582,In_291,In_1316);
or U583 (N_583,In_2521,In_2189);
nor U584 (N_584,In_597,In_1663);
and U585 (N_585,In_2909,In_2727);
nor U586 (N_586,In_1194,In_2463);
nand U587 (N_587,In_2123,In_2701);
and U588 (N_588,In_1915,In_1504);
nor U589 (N_589,In_1499,In_850);
and U590 (N_590,In_1216,In_1072);
and U591 (N_591,In_1180,In_821);
or U592 (N_592,In_787,In_931);
nand U593 (N_593,In_2496,In_712);
or U594 (N_594,In_1185,In_2528);
or U595 (N_595,In_1959,In_1006);
or U596 (N_596,In_1741,In_969);
nand U597 (N_597,In_1342,In_2292);
or U598 (N_598,In_1600,In_2966);
or U599 (N_599,In_124,In_2093);
nand U600 (N_600,In_251,N_29);
xnor U601 (N_601,In_238,N_215);
xnor U602 (N_602,N_72,N_447);
nor U603 (N_603,In_166,In_1580);
nor U604 (N_604,N_39,In_1287);
nand U605 (N_605,In_435,In_403);
xnor U606 (N_606,N_155,In_433);
nand U607 (N_607,N_138,In_799);
nand U608 (N_608,In_1025,In_826);
and U609 (N_609,In_1631,In_2302);
nand U610 (N_610,N_135,N_427);
nor U611 (N_611,In_1951,In_2332);
or U612 (N_612,N_53,In_2228);
or U613 (N_613,N_379,In_2406);
xor U614 (N_614,In_438,N_352);
xor U615 (N_615,N_195,N_262);
or U616 (N_616,In_1244,N_394);
nand U617 (N_617,N_228,In_1850);
xor U618 (N_618,N_421,In_1235);
nand U619 (N_619,N_49,In_2279);
or U620 (N_620,In_2305,In_2108);
and U621 (N_621,In_2028,N_524);
and U622 (N_622,N_444,N_187);
nand U623 (N_623,N_400,N_363);
and U624 (N_624,In_1894,In_955);
xor U625 (N_625,In_707,In_1164);
or U626 (N_626,N_376,In_1601);
nor U627 (N_627,N_517,N_176);
nor U628 (N_628,In_2921,In_710);
or U629 (N_629,N_239,In_1125);
nand U630 (N_630,N_289,In_770);
nor U631 (N_631,In_1367,In_768);
nor U632 (N_632,N_383,N_362);
nor U633 (N_633,In_765,N_274);
xnor U634 (N_634,In_2616,In_1414);
nand U635 (N_635,N_461,In_2175);
xnor U636 (N_636,In_1078,In_1919);
and U637 (N_637,In_600,In_2036);
xnor U638 (N_638,In_1651,In_2596);
nand U639 (N_639,In_602,In_458);
xor U640 (N_640,N_514,In_169);
and U641 (N_641,In_2903,N_579);
nor U642 (N_642,In_1720,In_2090);
xor U643 (N_643,In_1238,In_2590);
nand U644 (N_644,N_207,In_2024);
and U645 (N_645,N_593,N_50);
and U646 (N_646,In_2360,In_2665);
xnor U647 (N_647,In_625,N_546);
xnor U648 (N_648,In_2795,In_2158);
nor U649 (N_649,In_669,In_1068);
and U650 (N_650,In_933,In_2348);
nor U651 (N_651,In_2424,N_6);
xnor U652 (N_652,In_2513,In_857);
nor U653 (N_653,In_2534,N_361);
or U654 (N_654,In_827,In_1518);
nand U655 (N_655,In_1276,In_2983);
xor U656 (N_656,N_277,In_1063);
or U657 (N_657,N_17,In_2816);
nand U658 (N_658,In_570,In_789);
nor U659 (N_659,In_1568,In_2640);
nand U660 (N_660,N_157,In_2214);
nor U661 (N_661,In_2261,In_1028);
and U662 (N_662,In_341,In_2823);
xor U663 (N_663,In_283,In_923);
nand U664 (N_664,In_2385,In_684);
xor U665 (N_665,N_345,In_2699);
and U666 (N_666,In_2788,In_2698);
or U667 (N_667,In_1151,N_333);
nor U668 (N_668,In_1588,N_276);
nand U669 (N_669,In_769,In_24);
and U670 (N_670,N_54,In_1864);
and U671 (N_671,In_117,N_2);
nand U672 (N_672,N_93,In_348);
and U673 (N_673,In_1665,N_565);
and U674 (N_674,In_2522,In_250);
or U675 (N_675,In_2466,In_143);
or U676 (N_676,In_974,In_2410);
nor U677 (N_677,In_1815,In_2678);
nand U678 (N_678,N_271,In_661);
nor U679 (N_679,In_1488,N_484);
xnor U680 (N_680,In_1047,In_65);
nand U681 (N_681,In_2483,In_2475);
nor U682 (N_682,In_1826,In_450);
xor U683 (N_683,In_786,In_756);
or U684 (N_684,In_620,In_134);
or U685 (N_685,N_82,In_898);
nand U686 (N_686,N_359,In_1506);
or U687 (N_687,In_657,N_209);
nor U688 (N_688,N_519,In_2319);
xnor U689 (N_689,N_534,N_592);
nor U690 (N_690,In_889,N_453);
nand U691 (N_691,In_1077,In_1213);
or U692 (N_692,In_2346,N_173);
nand U693 (N_693,In_69,In_2945);
nand U694 (N_694,In_159,In_847);
nand U695 (N_695,In_66,In_2670);
or U696 (N_696,In_1299,In_207);
xnor U697 (N_697,In_2872,In_885);
and U698 (N_698,N_386,In_1521);
nand U699 (N_699,In_1764,N_321);
nand U700 (N_700,N_537,In_2712);
or U701 (N_701,In_2147,In_1439);
nor U702 (N_702,In_1119,In_421);
xnor U703 (N_703,In_1470,In_2586);
nor U704 (N_704,In_2003,In_876);
nand U705 (N_705,In_2268,In_240);
nand U706 (N_706,N_268,N_87);
nand U707 (N_707,In_256,In_511);
or U708 (N_708,In_1103,In_126);
or U709 (N_709,N_5,N_42);
xnor U710 (N_710,In_2227,In_705);
xor U711 (N_711,N_512,In_1364);
and U712 (N_712,N_142,In_1174);
nand U713 (N_713,In_1435,In_762);
nor U714 (N_714,In_2939,In_2197);
and U715 (N_715,In_614,In_1365);
xor U716 (N_716,In_130,In_1825);
xnor U717 (N_717,In_1339,In_2209);
xnor U718 (N_718,In_2040,In_164);
nor U719 (N_719,In_493,In_1779);
xnor U720 (N_720,In_108,In_808);
nand U721 (N_721,In_2112,In_362);
nand U722 (N_722,In_2952,In_180);
or U723 (N_723,N_315,In_1875);
or U724 (N_724,In_356,N_481);
or U725 (N_725,In_2520,In_649);
nor U726 (N_726,N_581,N_68);
xor U727 (N_727,In_2438,N_131);
xor U728 (N_728,In_1355,In_1632);
or U729 (N_729,In_1652,N_433);
and U730 (N_730,In_891,In_2870);
xor U731 (N_731,In_2317,In_2306);
or U732 (N_732,N_7,In_2592);
nor U733 (N_733,N_244,In_443);
nor U734 (N_734,In_539,In_2672);
xnor U735 (N_735,In_1333,In_267);
and U736 (N_736,In_478,In_2423);
xnor U737 (N_737,In_364,In_1802);
nor U738 (N_738,In_1405,In_1312);
xor U739 (N_739,In_2527,In_2270);
nand U740 (N_740,In_2490,In_1014);
nand U741 (N_741,In_2489,In_1487);
nand U742 (N_742,In_1765,In_2259);
nand U743 (N_743,In_1429,In_2659);
and U744 (N_744,In_2564,N_1);
xnor U745 (N_745,In_1633,In_2627);
nand U746 (N_746,In_598,In_934);
or U747 (N_747,In_2029,In_2401);
or U748 (N_748,In_2777,In_2806);
nand U749 (N_749,In_482,N_380);
nor U750 (N_750,In_2314,In_2953);
or U751 (N_751,In_55,In_1944);
nor U752 (N_752,N_184,In_1257);
and U753 (N_753,In_2288,In_1697);
nand U754 (N_754,In_781,N_146);
and U755 (N_755,In_2168,In_2087);
nand U756 (N_756,N_77,In_9);
xnor U757 (N_757,In_965,N_285);
or U758 (N_758,In_1182,In_755);
xor U759 (N_759,In_1226,In_865);
and U760 (N_760,N_490,In_2236);
nand U761 (N_761,In_399,In_2683);
or U762 (N_762,N_278,In_2454);
and U763 (N_763,In_122,N_258);
or U764 (N_764,In_1693,N_493);
and U765 (N_765,N_369,In_1933);
nand U766 (N_766,In_2232,In_2098);
nand U767 (N_767,N_62,In_2299);
nand U768 (N_768,In_297,N_74);
and U769 (N_769,In_156,N_381);
nand U770 (N_770,In_1679,In_1571);
nand U771 (N_771,In_2976,N_192);
nor U772 (N_772,N_70,N_165);
and U773 (N_773,N_97,In_354);
nor U774 (N_774,N_250,In_2085);
nor U775 (N_775,In_363,In_361);
nor U776 (N_776,In_1566,N_475);
nand U777 (N_777,In_461,In_2280);
nor U778 (N_778,In_2905,In_366);
and U779 (N_779,In_1052,In_98);
nand U780 (N_780,In_127,In_497);
and U781 (N_781,In_1017,In_2468);
or U782 (N_782,In_296,N_372);
or U783 (N_783,In_2943,N_75);
and U784 (N_784,In_2198,In_479);
and U785 (N_785,In_920,N_27);
nand U786 (N_786,N_334,In_749);
nor U787 (N_787,In_1683,In_2623);
xnor U788 (N_788,In_1637,N_341);
nor U789 (N_789,N_43,In_29);
or U790 (N_790,N_584,In_185);
and U791 (N_791,In_441,N_251);
nor U792 (N_792,N_197,In_2007);
or U793 (N_793,In_2000,In_2498);
and U794 (N_794,In_132,In_2555);
xnor U795 (N_795,In_2071,N_482);
xor U796 (N_796,In_2970,In_1073);
and U797 (N_797,In_1917,In_346);
xnor U798 (N_798,In_2537,In_1524);
nand U799 (N_799,In_1160,In_725);
or U800 (N_800,N_586,N_136);
or U801 (N_801,In_1688,In_1550);
or U802 (N_802,In_2012,In_2067);
nor U803 (N_803,In_901,In_2723);
nor U804 (N_804,In_1573,N_273);
nand U805 (N_805,In_2748,In_2059);
or U806 (N_806,In_814,N_203);
or U807 (N_807,In_1264,In_2264);
or U808 (N_808,In_1758,In_1798);
xnor U809 (N_809,In_1783,In_1788);
xnor U810 (N_810,In_1586,In_1352);
or U811 (N_811,N_476,In_623);
nand U812 (N_812,N_222,In_522);
and U813 (N_813,In_2354,In_2817);
xnor U814 (N_814,N_543,In_357);
xor U815 (N_815,In_2589,In_2469);
xnor U816 (N_816,N_118,N_491);
or U817 (N_817,In_2426,N_230);
nor U818 (N_818,In_49,In_2753);
nor U819 (N_819,In_13,In_1646);
xor U820 (N_820,N_527,In_258);
xor U821 (N_821,In_660,In_2663);
or U822 (N_822,In_844,N_322);
xor U823 (N_823,N_531,In_434);
and U824 (N_824,N_397,In_2356);
nor U825 (N_825,In_840,In_2134);
or U826 (N_826,In_1148,In_995);
and U827 (N_827,In_1886,In_2181);
nor U828 (N_828,In_1761,In_567);
nor U829 (N_829,In_1953,In_25);
nor U830 (N_830,N_237,In_641);
nand U831 (N_831,In_1111,N_407);
nand U832 (N_832,In_1039,In_2096);
nor U833 (N_833,In_1169,N_71);
nand U834 (N_834,N_382,In_674);
and U835 (N_835,In_1884,In_2655);
or U836 (N_836,N_243,In_389);
xor U837 (N_837,In_994,In_621);
xnor U838 (N_838,In_21,In_790);
and U839 (N_839,N_420,N_438);
nor U840 (N_840,N_403,In_140);
nand U841 (N_841,In_862,In_1326);
nand U842 (N_842,In_540,In_1486);
nor U843 (N_843,In_1901,In_1482);
nor U844 (N_844,In_2334,In_2762);
and U845 (N_845,In_345,In_442);
nor U846 (N_846,In_2333,In_328);
or U847 (N_847,In_2160,In_1385);
and U848 (N_848,In_1677,N_159);
or U849 (N_849,In_1106,N_439);
or U850 (N_850,N_233,In_1900);
or U851 (N_851,In_75,In_2883);
xnor U852 (N_852,In_1547,In_1997);
nor U853 (N_853,In_2174,N_545);
or U854 (N_854,In_2398,N_538);
nand U855 (N_855,In_2851,In_42);
nand U856 (N_856,In_2116,N_211);
nand U857 (N_857,In_1502,N_148);
nor U858 (N_858,In_1262,In_2793);
nand U859 (N_859,N_370,N_435);
xnor U860 (N_860,In_1344,In_1558);
or U861 (N_861,In_1946,In_2494);
nand U862 (N_862,N_129,N_123);
or U863 (N_863,In_2128,In_2714);
nand U864 (N_864,In_1186,In_2138);
nor U865 (N_865,N_90,In_895);
xnor U866 (N_866,In_1239,N_511);
and U867 (N_867,In_634,In_40);
or U868 (N_868,In_893,In_2825);
nand U869 (N_869,In_711,In_609);
nand U870 (N_870,In_2899,N_354);
or U871 (N_871,In_2997,N_163);
xnor U872 (N_872,N_521,In_243);
xnor U873 (N_873,In_761,N_120);
xor U874 (N_874,In_175,N_108);
and U875 (N_875,In_1845,In_418);
nor U876 (N_876,In_2853,N_301);
or U877 (N_877,In_1927,In_1069);
xnor U878 (N_878,In_2440,In_2525);
nor U879 (N_879,In_173,N_562);
or U880 (N_880,N_177,In_1082);
nor U881 (N_881,N_254,In_2514);
and U882 (N_882,In_1170,In_2282);
xnor U883 (N_883,In_2467,N_310);
xnor U884 (N_884,In_1595,In_1019);
and U885 (N_885,In_638,In_1706);
and U886 (N_886,In_2350,In_1726);
xnor U887 (N_887,N_181,N_535);
nor U888 (N_888,In_2038,In_954);
or U889 (N_889,In_1639,In_2412);
or U890 (N_890,In_92,In_802);
or U891 (N_891,In_2263,In_2781);
or U892 (N_892,In_2213,In_292);
nor U893 (N_893,In_2583,In_234);
xnor U894 (N_894,In_2200,In_1242);
xnor U895 (N_895,In_278,In_936);
nor U896 (N_896,In_1549,In_812);
nand U897 (N_897,In_1778,N_56);
nor U898 (N_898,N_193,N_448);
xnor U899 (N_899,N_208,In_825);
nand U900 (N_900,N_570,N_540);
nor U901 (N_901,N_216,In_811);
nand U902 (N_902,In_2947,In_1729);
nor U903 (N_903,In_1497,N_249);
xor U904 (N_904,In_494,In_1507);
and U905 (N_905,N_65,In_1820);
and U906 (N_906,In_2246,N_22);
nand U907 (N_907,In_1948,In_2250);
or U908 (N_908,In_307,In_1591);
nand U909 (N_909,In_2009,In_397);
nand U910 (N_910,N_13,In_2858);
nor U911 (N_911,In_2829,N_164);
and U912 (N_912,N_196,In_2449);
nor U913 (N_913,In_1842,In_1215);
nor U914 (N_914,In_2035,In_2710);
or U915 (N_915,In_612,In_2987);
nand U916 (N_916,In_2570,In_2167);
nor U917 (N_917,N_8,In_2149);
or U918 (N_918,In_1618,In_1135);
nand U919 (N_919,N_47,N_314);
nor U920 (N_920,In_1381,N_117);
nand U921 (N_921,N_219,In_1810);
nand U922 (N_922,In_507,In_2730);
nor U923 (N_923,N_557,N_446);
xnor U924 (N_924,N_331,N_293);
or U925 (N_925,In_1644,In_938);
xnor U926 (N_926,In_882,N_469);
or U927 (N_927,In_582,In_874);
or U928 (N_928,N_127,N_202);
and U929 (N_929,N_319,N_459);
or U930 (N_930,N_429,In_2884);
or U931 (N_931,In_276,In_1931);
or U932 (N_932,In_1849,In_2882);
or U933 (N_933,In_1996,In_2231);
nor U934 (N_934,In_2061,In_574);
xor U935 (N_935,In_1361,In_1484);
xnor U936 (N_936,In_2474,In_1297);
and U937 (N_937,In_1834,In_2323);
and U938 (N_938,In_668,In_1692);
and U939 (N_939,In_287,In_1045);
xnor U940 (N_940,In_171,In_1622);
or U941 (N_941,N_480,In_2532);
or U942 (N_942,In_1904,N_455);
xor U943 (N_943,In_152,N_351);
nor U944 (N_944,In_2086,N_201);
or U945 (N_945,In_104,N_101);
nor U946 (N_946,N_158,In_1774);
nor U947 (N_947,In_1015,N_64);
xnor U948 (N_948,In_1270,N_353);
nor U949 (N_949,In_1317,In_2068);
nor U950 (N_950,In_1420,N_297);
or U951 (N_951,In_1611,In_1055);
xnor U952 (N_952,In_503,In_14);
nor U953 (N_953,N_488,In_2739);
nor U954 (N_954,In_253,In_1561);
nand U955 (N_955,In_2892,N_105);
nand U956 (N_956,In_1989,In_2798);
and U957 (N_957,N_89,N_217);
nand U958 (N_958,N_358,In_1225);
xor U959 (N_959,In_617,N_402);
and U960 (N_960,In_2184,In_595);
or U961 (N_961,In_911,In_1829);
nor U962 (N_962,In_2874,In_961);
nand U963 (N_963,In_1939,In_1471);
nor U964 (N_964,In_1950,N_189);
and U965 (N_965,In_1379,In_2658);
xnor U966 (N_966,In_937,In_2033);
or U967 (N_967,In_85,In_12);
xor U968 (N_968,In_2077,N_154);
nand U969 (N_969,In_266,In_737);
xor U970 (N_970,In_1711,In_2309);
nand U971 (N_971,In_2394,N_137);
nand U972 (N_972,N_51,In_2127);
nor U973 (N_973,In_544,In_1036);
and U974 (N_974,In_1129,In_741);
and U975 (N_975,In_2869,N_536);
and U976 (N_976,In_2223,N_539);
or U977 (N_977,In_1166,In_2145);
nor U978 (N_978,In_2417,In_2578);
nand U979 (N_979,In_861,In_2247);
nand U980 (N_980,N_377,In_2179);
or U981 (N_981,N_585,In_2199);
and U982 (N_982,In_2860,In_294);
and U983 (N_983,In_1474,N_458);
or U984 (N_984,N_103,In_2950);
xor U985 (N_985,In_1742,N_445);
xor U986 (N_986,N_3,In_197);
nor U987 (N_987,In_2060,In_820);
nand U988 (N_988,N_205,In_1682);
xor U989 (N_989,In_1134,N_79);
or U990 (N_990,In_205,N_388);
nand U991 (N_991,In_919,N_124);
nor U992 (N_992,In_456,In_2082);
and U993 (N_993,In_716,N_419);
nor U994 (N_994,In_1049,In_1179);
or U995 (N_995,In_2053,In_2808);
nand U996 (N_996,In_178,In_2177);
and U997 (N_997,In_1776,In_28);
or U998 (N_998,In_154,In_2432);
nand U999 (N_999,In_284,In_565);
xor U1000 (N_1000,In_2166,In_870);
and U1001 (N_1001,In_551,N_560);
and U1002 (N_1002,In_2368,N_225);
nor U1003 (N_1003,In_352,In_1736);
and U1004 (N_1004,In_2393,In_217);
xor U1005 (N_1005,N_499,In_2631);
or U1006 (N_1006,In_1782,In_1920);
or U1007 (N_1007,N_503,In_11);
nor U1008 (N_1008,In_2512,In_576);
or U1009 (N_1009,In_1124,In_2729);
or U1010 (N_1010,N_485,N_263);
nor U1011 (N_1011,N_378,In_306);
and U1012 (N_1012,N_151,In_1701);
nand U1013 (N_1013,N_418,In_2117);
and U1014 (N_1014,In_112,In_1887);
xor U1015 (N_1015,In_2544,In_2745);
and U1016 (N_1016,In_837,In_2006);
xor U1017 (N_1017,In_2929,In_2225);
and U1018 (N_1018,In_194,N_357);
and U1019 (N_1019,In_983,In_1455);
nand U1020 (N_1020,In_1426,N_99);
nand U1021 (N_1021,In_1360,N_336);
nand U1022 (N_1022,N_307,In_958);
nand U1023 (N_1023,In_2750,N_513);
or U1024 (N_1024,In_877,N_259);
nor U1025 (N_1025,In_1258,N_568);
or U1026 (N_1026,N_549,In_2920);
or U1027 (N_1027,In_1403,In_1477);
nand U1028 (N_1028,N_141,In_19);
xnor U1029 (N_1029,In_1222,In_136);
nor U1030 (N_1030,In_2927,N_145);
xnor U1031 (N_1031,In_1328,N_431);
or U1032 (N_1032,In_1462,N_212);
nand U1033 (N_1033,N_299,In_498);
and U1034 (N_1034,In_1723,In_782);
xnor U1035 (N_1035,In_1751,In_2239);
and U1036 (N_1036,In_231,In_1659);
or U1037 (N_1037,In_1952,In_845);
xor U1038 (N_1038,In_2384,In_2601);
xnor U1039 (N_1039,In_1510,In_1918);
or U1040 (N_1040,N_257,In_616);
or U1041 (N_1041,In_887,In_1535);
or U1042 (N_1042,N_256,In_2262);
nand U1043 (N_1043,In_1908,In_2501);
or U1044 (N_1044,In_446,In_1641);
and U1045 (N_1045,In_144,In_2800);
or U1046 (N_1046,N_424,In_1117);
xnor U1047 (N_1047,N_21,In_1234);
xnor U1048 (N_1048,In_2956,In_1000);
and U1049 (N_1049,In_1839,In_2700);
nand U1050 (N_1050,N_111,In_1197);
xor U1051 (N_1051,In_1221,In_2219);
and U1052 (N_1052,In_2163,In_677);
xor U1053 (N_1053,In_274,In_1175);
nand U1054 (N_1054,N_45,In_1059);
xnor U1055 (N_1055,In_2470,In_2152);
and U1056 (N_1056,In_1115,In_607);
nor U1057 (N_1057,In_111,In_1540);
nor U1058 (N_1058,In_105,N_561);
xor U1059 (N_1059,N_311,In_1033);
nor U1060 (N_1060,In_110,In_1315);
xor U1061 (N_1061,In_1657,In_939);
nor U1062 (N_1062,In_204,In_2751);
nor U1063 (N_1063,In_1903,In_560);
and U1064 (N_1064,In_314,In_1831);
and U1065 (N_1065,In_2815,N_291);
nand U1066 (N_1066,N_96,In_1468);
and U1067 (N_1067,In_2072,N_86);
nor U1068 (N_1068,In_1190,In_1122);
nand U1069 (N_1069,In_554,In_2164);
or U1070 (N_1070,In_1500,In_2554);
nand U1071 (N_1071,In_888,In_2602);
xor U1072 (N_1072,In_890,N_52);
nor U1073 (N_1073,In_1255,In_2991);
and U1074 (N_1074,In_1817,In_1399);
and U1075 (N_1075,In_1599,N_408);
nor U1076 (N_1076,In_1491,In_1966);
and U1077 (N_1077,In_1843,In_337);
nor U1078 (N_1078,In_1383,In_2320);
nand U1079 (N_1079,In_2918,In_2062);
nor U1080 (N_1080,In_2799,In_1304);
xor U1081 (N_1081,In_2266,In_1346);
and U1082 (N_1082,In_1674,N_309);
or U1083 (N_1083,N_498,In_1916);
and U1084 (N_1084,In_1165,N_204);
xnor U1085 (N_1085,In_2871,In_1556);
and U1086 (N_1086,In_350,In_1436);
or U1087 (N_1087,In_101,In_1560);
nor U1088 (N_1088,N_19,In_1120);
nor U1089 (N_1089,In_486,In_1493);
xnor U1090 (N_1090,N_387,In_1520);
nand U1091 (N_1091,In_36,In_2890);
and U1092 (N_1092,N_150,In_1854);
nand U1093 (N_1093,N_199,In_2782);
and U1094 (N_1094,In_1844,In_2478);
nor U1095 (N_1095,In_492,N_160);
nand U1096 (N_1096,N_279,In_2094);
nand U1097 (N_1097,In_2363,In_1724);
or U1098 (N_1098,N_296,N_34);
nor U1099 (N_1099,In_1553,In_1018);
xor U1100 (N_1100,In_530,N_576);
or U1101 (N_1101,In_1263,In_2695);
and U1102 (N_1102,N_526,N_500);
xor U1103 (N_1103,In_454,In_2573);
and U1104 (N_1104,In_1116,In_155);
and U1105 (N_1105,In_367,N_312);
and U1106 (N_1106,In_1300,In_1819);
nor U1107 (N_1107,In_2375,N_583);
nand U1108 (N_1108,In_2937,N_479);
nor U1109 (N_1109,In_214,N_492);
or U1110 (N_1110,N_390,In_2638);
nand U1111 (N_1111,In_779,N_149);
and U1112 (N_1112,In_2603,In_2877);
nor U1113 (N_1113,N_597,In_54);
or U1114 (N_1114,In_1301,In_2043);
nor U1115 (N_1115,In_1095,In_1559);
nand U1116 (N_1116,N_305,In_1822);
and U1117 (N_1117,In_1957,N_395);
or U1118 (N_1118,In_1752,In_1709);
nor U1119 (N_1119,N_300,N_374);
or U1120 (N_1120,N_32,In_1337);
and U1121 (N_1121,In_1406,In_2685);
xor U1122 (N_1122,In_1899,In_2886);
xor U1123 (N_1123,N_81,In_2431);
or U1124 (N_1124,In_947,In_1718);
and U1125 (N_1125,In_1992,In_687);
and U1126 (N_1126,In_2734,In_1750);
nand U1127 (N_1127,N_59,In_72);
nand U1128 (N_1128,In_1308,N_20);
and U1129 (N_1129,In_1083,In_1022);
nand U1130 (N_1130,In_2442,In_2850);
nor U1131 (N_1131,In_2637,N_183);
nor U1132 (N_1132,In_2193,In_1994);
or U1133 (N_1133,In_2715,N_344);
xor U1134 (N_1134,In_2711,In_70);
or U1135 (N_1135,In_2310,In_114);
or U1136 (N_1136,In_2039,N_404);
nor U1137 (N_1137,In_1567,In_416);
or U1138 (N_1138,N_456,In_585);
nor U1139 (N_1139,In_2958,In_2422);
nand U1140 (N_1140,In_846,In_1892);
or U1141 (N_1141,N_161,In_2275);
nand U1142 (N_1142,In_2995,N_231);
nor U1143 (N_1143,N_450,In_90);
or U1144 (N_1144,In_1382,N_552);
and U1145 (N_1145,In_688,In_1227);
nand U1146 (N_1146,N_116,In_1035);
nand U1147 (N_1147,N_468,In_2054);
xor U1148 (N_1148,In_1717,In_1528);
and U1149 (N_1149,In_1835,In_84);
or U1150 (N_1150,N_206,In_192);
nand U1151 (N_1151,N_422,In_987);
xor U1152 (N_1152,In_940,In_2484);
xnor U1153 (N_1153,In_916,In_1574);
xor U1154 (N_1154,In_2946,In_1552);
nor U1155 (N_1155,N_288,In_2185);
and U1156 (N_1156,In_568,In_2503);
nor U1157 (N_1157,In_2330,N_188);
nor U1158 (N_1158,In_881,In_1698);
nor U1159 (N_1159,N_88,N_320);
and U1160 (N_1160,In_1146,In_2756);
nand U1161 (N_1161,In_1431,In_1434);
and U1162 (N_1162,In_1814,N_194);
and U1163 (N_1163,N_171,In_550);
xnor U1164 (N_1164,In_2221,In_1162);
nand U1165 (N_1165,In_1253,In_2841);
nand U1166 (N_1166,In_1539,In_2027);
or U1167 (N_1167,In_971,In_382);
xnor U1168 (N_1168,In_305,In_1719);
nor U1169 (N_1169,N_236,In_2107);
nand U1170 (N_1170,N_147,In_2188);
and U1171 (N_1171,In_2351,In_6);
xnor U1172 (N_1172,In_2610,N_264);
and U1173 (N_1173,In_2176,In_1126);
nand U1174 (N_1174,N_442,N_281);
nand U1175 (N_1175,N_544,In_76);
or U1176 (N_1176,In_2847,In_1040);
or U1177 (N_1177,N_80,In_44);
nor U1178 (N_1178,N_232,In_1800);
xor U1179 (N_1179,N_572,In_2413);
nor U1180 (N_1180,N_587,In_579);
nand U1181 (N_1181,In_146,In_2081);
nand U1182 (N_1182,In_1370,In_1020);
xnor U1183 (N_1183,In_1570,In_20);
or U1184 (N_1184,In_2764,N_452);
nor U1185 (N_1185,In_46,In_2636);
nand U1186 (N_1186,N_595,N_265);
nor U1187 (N_1187,In_1890,N_487);
or U1188 (N_1188,In_2367,In_2626);
and U1189 (N_1189,In_1448,In_2620);
nor U1190 (N_1190,N_198,In_927);
or U1191 (N_1191,In_1608,In_1678);
or U1192 (N_1192,In_2612,N_384);
or U1193 (N_1193,In_2020,N_467);
or U1194 (N_1194,N_396,In_59);
nand U1195 (N_1195,In_331,In_714);
and U1196 (N_1196,In_809,In_1096);
xor U1197 (N_1197,In_371,In_619);
or U1198 (N_1198,In_533,In_374);
and U1199 (N_1199,N_33,N_113);
xnor U1200 (N_1200,N_708,N_615);
or U1201 (N_1201,N_1096,In_1277);
and U1202 (N_1202,N_182,In_650);
and U1203 (N_1203,In_2611,N_253);
or U1204 (N_1204,In_2341,N_693);
or U1205 (N_1205,N_1118,N_846);
or U1206 (N_1206,In_187,In_484);
xor U1207 (N_1207,N_9,In_1772);
nor U1208 (N_1208,In_2551,N_893);
and U1209 (N_1209,N_744,In_682);
or U1210 (N_1210,In_685,In_694);
xnor U1211 (N_1211,In_2819,In_1433);
nor U1212 (N_1212,In_265,In_1861);
xor U1213 (N_1213,In_2811,In_823);
xor U1214 (N_1214,N_681,N_884);
nor U1215 (N_1215,N_410,In_277);
or U1216 (N_1216,In_1876,N_489);
xnor U1217 (N_1217,In_1749,In_339);
or U1218 (N_1218,N_668,N_152);
xor U1219 (N_1219,N_966,N_731);
nand U1220 (N_1220,N_747,N_272);
nand U1221 (N_1221,In_2300,In_1513);
or U1222 (N_1222,In_830,N_223);
nand U1223 (N_1223,In_945,N_881);
or U1224 (N_1224,In_2395,N_306);
nand U1225 (N_1225,N_355,N_746);
or U1226 (N_1226,N_673,In_2530);
nand U1227 (N_1227,N_1169,N_1135);
nand U1228 (N_1228,In_2895,N_862);
nand U1229 (N_1229,N_718,In_184);
nor U1230 (N_1230,N_776,N_1180);
and U1231 (N_1231,In_1016,N_1076);
xor U1232 (N_1232,In_1208,In_2562);
or U1233 (N_1233,N_601,In_2047);
nand U1234 (N_1234,In_485,In_2518);
xnor U1235 (N_1235,N_892,N_952);
and U1236 (N_1236,N_67,N_782);
or U1237 (N_1237,In_1009,In_1984);
nand U1238 (N_1238,N_698,In_2017);
and U1239 (N_1239,In_806,In_2142);
xnor U1240 (N_1240,N_302,In_977);
xnor U1241 (N_1241,N_1125,In_719);
nor U1242 (N_1242,In_1260,In_424);
nand U1243 (N_1243,N_413,In_1171);
nand U1244 (N_1244,N_94,In_1694);
or U1245 (N_1245,N_722,N_36);
xnor U1246 (N_1246,In_1099,In_2736);
and U1247 (N_1247,N_715,In_2);
and U1248 (N_1248,In_77,In_2392);
nand U1249 (N_1249,N_133,N_1050);
nand U1250 (N_1250,In_1206,In_2345);
nand U1251 (N_1251,N_738,In_2994);
nor U1252 (N_1252,In_2733,N_786);
or U1253 (N_1253,In_94,In_2679);
or U1254 (N_1254,N_1163,N_26);
and U1255 (N_1255,In_1687,N_1168);
nor U1256 (N_1256,N_436,In_1610);
and U1257 (N_1257,In_2574,In_1867);
nor U1258 (N_1258,In_1740,N_855);
nor U1259 (N_1259,In_202,In_942);
or U1260 (N_1260,In_1267,In_1085);
xnor U1261 (N_1261,In_208,In_2630);
nand U1262 (N_1262,In_133,In_1684);
and U1263 (N_1263,In_2552,In_2741);
nor U1264 (N_1264,In_2654,N_778);
nor U1265 (N_1265,In_206,N_261);
or U1266 (N_1266,N_705,N_1032);
and U1267 (N_1267,In_2131,In_2460);
xor U1268 (N_1268,N_750,N_547);
or U1269 (N_1269,N_471,In_160);
and U1270 (N_1270,In_244,N_948);
xnor U1271 (N_1271,In_2409,N_441);
nand U1272 (N_1272,In_2768,In_2157);
or U1273 (N_1273,N_497,N_878);
and U1274 (N_1274,In_523,N_864);
nand U1275 (N_1275,In_1823,In_1605);
nor U1276 (N_1276,In_2584,In_50);
or U1277 (N_1277,N_825,N_247);
xnor U1278 (N_1278,In_1423,In_1645);
xor U1279 (N_1279,N_226,In_2014);
or U1280 (N_1280,In_2316,N_712);
and U1281 (N_1281,In_2208,N_767);
nand U1282 (N_1282,N_774,In_393);
nand U1283 (N_1283,N_507,In_2881);
xor U1284 (N_1284,In_1785,In_2421);
nor U1285 (N_1285,N_1091,N_430);
or U1286 (N_1286,In_241,In_692);
xnor U1287 (N_1287,N_775,In_513);
nor U1288 (N_1288,In_534,N_666);
xor U1289 (N_1289,N_629,In_1673);
nand U1290 (N_1290,In_2747,In_245);
xor U1291 (N_1291,In_2772,N_787);
nor U1292 (N_1292,In_472,N_885);
or U1293 (N_1293,N_662,In_1309);
nand U1294 (N_1294,In_2365,N_719);
xor U1295 (N_1295,In_1445,N_806);
nand U1296 (N_1296,In_842,N_734);
or U1297 (N_1297,In_1387,N_186);
and U1298 (N_1298,In_1809,N_1142);
nand U1299 (N_1299,N_912,N_869);
nor U1300 (N_1300,In_2803,N_868);
nand U1301 (N_1301,In_2477,N_532);
nand U1302 (N_1302,N_753,N_84);
and U1303 (N_1303,N_982,N_1023);
or U1304 (N_1304,N_179,N_889);
nand U1305 (N_1305,N_275,In_45);
nand U1306 (N_1306,N_899,N_770);
xor U1307 (N_1307,In_230,N_1106);
xnor U1308 (N_1308,In_349,N_1019);
nor U1309 (N_1309,N_642,In_2194);
and U1310 (N_1310,N_598,N_1022);
nor U1311 (N_1311,In_632,In_2414);
and U1312 (N_1312,In_1050,N_1016);
or U1313 (N_1313,In_1086,N_663);
nand U1314 (N_1314,In_1064,In_1906);
or U1315 (N_1315,N_682,In_1416);
and U1316 (N_1316,N_1160,In_2129);
nand U1317 (N_1317,N_1147,In_359);
or U1318 (N_1318,N_874,N_802);
nand U1319 (N_1319,N_670,N_832);
and U1320 (N_1320,N_416,N_975);
nand U1321 (N_1321,In_1766,N_858);
xor U1322 (N_1322,N_566,In_477);
nor U1323 (N_1323,N_853,In_2978);
nand U1324 (N_1324,N_974,N_367);
or U1325 (N_1325,In_153,N_1074);
xor U1326 (N_1326,N_529,In_2472);
or U1327 (N_1327,In_408,In_2291);
xnor U1328 (N_1328,N_1020,In_33);
nor U1329 (N_1329,In_897,In_601);
and U1330 (N_1330,N_1053,N_1094);
nand U1331 (N_1331,N_762,N_841);
and U1332 (N_1332,N_654,N_882);
nor U1333 (N_1333,N_440,In_907);
nor U1334 (N_1334,N_934,In_2791);
or U1335 (N_1335,In_500,N_849);
nand U1336 (N_1336,N_988,N_977);
or U1337 (N_1337,In_2591,In_481);
xor U1338 (N_1338,N_1075,N_859);
or U1339 (N_1339,In_2643,N_1171);
and U1340 (N_1340,In_785,N_25);
nor U1341 (N_1341,N_824,In_58);
and U1342 (N_1342,In_38,In_1555);
nand U1343 (N_1343,In_1447,N_340);
nand U1344 (N_1344,In_2447,In_86);
or U1345 (N_1345,In_2587,In_2889);
nand U1346 (N_1346,In_2560,N_1082);
or U1347 (N_1347,N_730,N_1165);
or U1348 (N_1348,In_2344,N_415);
and U1349 (N_1349,N_41,N_895);
nand U1350 (N_1350,In_2720,N_144);
xnor U1351 (N_1351,N_132,In_2849);
nand U1352 (N_1352,N_971,In_1202);
and U1353 (N_1353,N_582,In_968);
nand U1354 (N_1354,N_252,N_925);
xor U1355 (N_1355,N_792,N_867);
or U1356 (N_1356,N_18,In_2226);
and U1357 (N_1357,N_28,In_318);
nor U1358 (N_1358,In_2902,N_830);
nor U1359 (N_1359,In_260,In_2079);
and U1360 (N_1360,N_426,N_63);
or U1361 (N_1361,N_953,N_961);
nand U1362 (N_1362,In_2579,N_796);
or U1363 (N_1363,In_1102,In_384);
xnor U1364 (N_1364,N_496,In_504);
and U1365 (N_1365,In_774,In_2744);
xor U1366 (N_1366,In_999,N_1130);
xnor U1367 (N_1367,In_2632,In_678);
nand U1368 (N_1368,N_240,N_409);
and U1369 (N_1369,N_328,N_104);
xnor U1370 (N_1370,In_1780,N_590);
nor U1371 (N_1371,N_1190,N_1131);
nand U1372 (N_1372,In_1965,N_246);
and U1373 (N_1373,In_1053,N_1126);
or U1374 (N_1374,In_1987,N_1011);
nand U1375 (N_1375,N_643,In_2864);
and U1376 (N_1376,In_1589,In_2313);
xnor U1377 (N_1377,N_1187,In_1030);
nand U1378 (N_1378,In_871,N_835);
xnor U1379 (N_1379,N_789,In_2269);
nor U1380 (N_1380,N_736,N_1060);
and U1381 (N_1381,N_1157,N_900);
nor U1382 (N_1382,In_2272,In_2671);
or U1383 (N_1383,In_116,In_1026);
xor U1384 (N_1384,In_1023,N_365);
or U1385 (N_1385,In_1091,In_1743);
and U1386 (N_1386,In_2962,In_2234);
and U1387 (N_1387,N_818,In_1837);
and U1388 (N_1388,N_857,N_423);
nor U1389 (N_1389,In_149,N_1141);
nor U1390 (N_1390,N_737,In_775);
nand U1391 (N_1391,In_1322,In_2162);
nand U1392 (N_1392,N_1087,In_378);
and U1393 (N_1393,In_2876,In_131);
nor U1394 (N_1394,N_347,In_2271);
or U1395 (N_1395,N_1110,N_1112);
nand U1396 (N_1396,N_614,N_57);
nor U1397 (N_1397,In_978,In_2582);
nand U1398 (N_1398,N_414,In_532);
or U1399 (N_1399,N_627,N_927);
nor U1400 (N_1400,In_496,N_1054);
xnor U1401 (N_1401,In_37,In_1787);
nand U1402 (N_1402,N_577,N_214);
nor U1403 (N_1403,In_1961,N_804);
nand U1404 (N_1404,In_1638,N_360);
or U1405 (N_1405,N_473,In_1797);
and U1406 (N_1406,In_1534,N_640);
nand U1407 (N_1407,In_2855,N_411);
or U1408 (N_1408,N_724,N_495);
xor U1409 (N_1409,In_198,N_78);
or U1410 (N_1410,In_2386,In_1002);
and U1411 (N_1411,N_916,In_2405);
nor U1412 (N_1412,N_375,In_468);
and U1413 (N_1413,N_852,In_39);
nand U1414 (N_1414,In_1183,In_489);
nor U1415 (N_1415,In_225,In_2318);
xnor U1416 (N_1416,N_772,In_1554);
and U1417 (N_1417,N_156,N_323);
and U1418 (N_1418,In_62,N_700);
xnor U1419 (N_1419,N_608,In_1712);
nor U1420 (N_1420,N_564,N_650);
or U1421 (N_1421,In_910,N_958);
nor U1422 (N_1422,In_833,In_1686);
or U1423 (N_1423,In_2878,In_327);
or U1424 (N_1424,In_2614,In_1377);
and U1425 (N_1425,N_1148,In_2556);
nand U1426 (N_1426,N_993,In_2371);
xor U1427 (N_1427,In_1268,In_626);
xor U1428 (N_1428,N_1001,N_260);
nor U1429 (N_1429,In_1237,N_509);
nand U1430 (N_1430,N_733,In_1259);
xnor U1431 (N_1431,N_763,N_876);
nand U1432 (N_1432,In_1157,In_2202);
nor U1433 (N_1433,In_1569,N_992);
or U1434 (N_1434,In_1548,In_1417);
nor U1435 (N_1435,N_1088,N_745);
nand U1436 (N_1436,In_2728,In_1195);
xor U1437 (N_1437,In_2773,N_632);
nor U1438 (N_1438,In_1411,N_1132);
xor U1439 (N_1439,N_1124,In_473);
nand U1440 (N_1440,N_1086,N_520);
nand U1441 (N_1441,N_843,In_308);
nand U1442 (N_1442,In_1594,In_264);
and U1443 (N_1443,In_803,In_1178);
xnor U1444 (N_1444,N_946,In_1964);
nand U1445 (N_1445,N_1017,In_68);
or U1446 (N_1446,In_884,In_332);
or U1447 (N_1447,N_761,In_525);
nand U1448 (N_1448,N_58,In_1929);
and U1449 (N_1449,N_630,In_2891);
nand U1450 (N_1450,N_811,In_2139);
nor U1451 (N_1451,N_817,In_520);
and U1452 (N_1452,In_1029,In_338);
or U1453 (N_1453,In_713,N_1031);
nand U1454 (N_1454,In_2928,In_2688);
nand U1455 (N_1455,N_847,In_106);
and U1456 (N_1456,In_2804,N_871);
or U1457 (N_1457,N_1101,N_1012);
and U1458 (N_1458,In_2502,In_128);
nand U1459 (N_1459,In_2030,N_126);
nand U1460 (N_1460,In_248,N_677);
xnor U1461 (N_1461,N_765,N_60);
or U1462 (N_1462,N_985,N_773);
and U1463 (N_1463,N_917,N_945);
nand U1464 (N_1464,N_965,N_611);
nand U1465 (N_1465,In_2585,In_2822);
nor U1466 (N_1466,N_674,In_286);
or U1467 (N_1467,In_949,N_980);
xnor U1468 (N_1468,In_2930,N_1052);
nor U1469 (N_1469,In_1398,N_687);
nand U1470 (N_1470,In_1768,N_1161);
xor U1471 (N_1471,N_434,In_1716);
or U1472 (N_1472,In_1348,N_938);
and U1473 (N_1473,N_684,In_1132);
or U1474 (N_1474,In_2286,N_1073);
nor U1475 (N_1475,In_2705,In_452);
and U1476 (N_1476,N_449,N_1099);
xor U1477 (N_1477,In_693,In_2140);
or U1478 (N_1478,N_720,N_851);
or U1479 (N_1479,In_673,In_1888);
xor U1480 (N_1480,N_1061,In_1604);
nand U1481 (N_1481,N_652,N_797);
nand U1482 (N_1482,N_588,N_1030);
xnor U1483 (N_1483,In_1409,In_228);
nor U1484 (N_1484,In_270,In_747);
xnor U1485 (N_1485,In_27,In_1516);
and U1486 (N_1486,In_2687,N_555);
nor U1487 (N_1487,In_464,N_15);
xnor U1488 (N_1488,N_556,N_647);
xnor U1489 (N_1489,In_2277,In_666);
nand U1490 (N_1490,In_986,N_143);
xor U1491 (N_1491,In_1076,N_1115);
nor U1492 (N_1492,In_1223,N_1154);
xnor U1493 (N_1493,In_1902,In_1508);
nand U1494 (N_1494,In_380,N_609);
xor U1495 (N_1495,In_1737,N_1102);
and U1496 (N_1496,In_41,In_2042);
nand U1497 (N_1497,N_842,N_888);
and U1498 (N_1498,In_2704,N_292);
and U1499 (N_1499,In_2567,In_2493);
xor U1500 (N_1500,N_840,N_685);
and U1501 (N_1501,N_742,N_553);
or U1502 (N_1502,In_1620,In_767);
xor U1503 (N_1503,N_1174,In_2441);
or U1504 (N_1504,N_478,N_69);
xnor U1505 (N_1505,In_1140,N_589);
nor U1506 (N_1506,In_2156,N_114);
xnor U1507 (N_1507,N_613,In_2321);
nand U1508 (N_1508,N_1029,In_93);
nor U1509 (N_1509,In_1250,N_959);
or U1510 (N_1510,In_61,In_1224);
xor U1511 (N_1511,In_841,N_1105);
nor U1512 (N_1512,In_2676,N_955);
or U1513 (N_1513,N_743,In_2005);
nand U1514 (N_1514,In_2684,In_2757);
nor U1515 (N_1515,In_2428,N_669);
nand U1516 (N_1516,In_2178,N_1145);
nor U1517 (N_1517,In_516,In_67);
nor U1518 (N_1518,In_739,N_472);
nor U1519 (N_1519,N_172,N_502);
nand U1520 (N_1520,N_638,In_2076);
nor U1521 (N_1521,N_741,N_234);
nor U1522 (N_1522,N_594,In_222);
or U1523 (N_1523,In_2792,In_2329);
nand U1524 (N_1524,N_162,In_302);
and U1525 (N_1525,In_176,In_383);
and U1526 (N_1526,In_480,In_868);
or U1527 (N_1527,N_1006,In_1838);
and U1528 (N_1528,N_1136,In_2832);
nor U1529 (N_1529,N_1025,N_998);
nor U1530 (N_1530,In_391,N_617);
nand U1531 (N_1531,In_1461,N_826);
nor U1532 (N_1532,In_414,N_748);
nor U1533 (N_1533,N_428,N_704);
nand U1534 (N_1534,In_2517,N_873);
nand U1535 (N_1535,N_1097,N_861);
xnor U1536 (N_1536,In_512,N_1067);
xor U1537 (N_1537,In_1976,In_824);
nor U1538 (N_1538,In_1851,N_1116);
and U1539 (N_1539,N_1120,In_1282);
nand U1540 (N_1540,N_978,N_740);
and U1541 (N_1541,N_170,N_729);
nor U1542 (N_1542,N_1194,N_870);
xnor U1543 (N_1543,In_1437,N_967);
nor U1544 (N_1544,In_1689,In_2963);
or U1545 (N_1545,In_96,N_1018);
nor U1546 (N_1546,N_723,In_319);
nand U1547 (N_1547,N_373,In_2304);
or U1548 (N_1548,In_2411,N_1043);
or U1549 (N_1549,N_989,N_898);
xnor U1550 (N_1550,In_87,In_2516);
nand U1551 (N_1551,In_1542,In_1543);
or U1552 (N_1552,N_735,N_1137);
or U1553 (N_1553,N_896,In_53);
nand U1554 (N_1554,In_913,In_451);
nor U1555 (N_1555,N_904,In_2046);
xnor U1556 (N_1556,In_1753,In_315);
or U1557 (N_1557,In_1748,N_850);
or U1558 (N_1558,N_432,In_1306);
nor U1559 (N_1559,N_591,In_138);
or U1560 (N_1560,In_2104,N_714);
and U1561 (N_1561,In_215,N_921);
or U1562 (N_1562,In_1199,N_1198);
and U1563 (N_1563,N_935,N_1103);
xor U1564 (N_1564,In_347,In_648);
or U1565 (N_1565,N_255,N_342);
or U1566 (N_1566,In_2848,In_892);
nand U1567 (N_1567,N_909,N_665);
nand U1568 (N_1568,In_2622,N_783);
nand U1569 (N_1569,In_930,N_860);
xor U1570 (N_1570,N_1155,In_2538);
and U1571 (N_1571,In_2335,In_304);
or U1572 (N_1572,In_2936,In_2019);
nand U1573 (N_1573,N_659,N_596);
xnor U1574 (N_1574,N_865,In_2342);
and U1575 (N_1575,N_1085,N_1108);
nand U1576 (N_1576,In_289,N_1038);
nor U1577 (N_1577,In_16,N_604);
xnor U1578 (N_1578,In_409,N_284);
nor U1579 (N_1579,In_900,In_26);
or U1580 (N_1580,N_690,N_914);
nor U1581 (N_1581,N_180,In_2400);
xnor U1582 (N_1582,In_935,In_2673);
xor U1583 (N_1583,N_66,In_2508);
or U1584 (N_1584,N_618,In_776);
xor U1585 (N_1585,N_463,N_1127);
xnor U1586 (N_1586,In_1848,In_1614);
nor U1587 (N_1587,N_1065,In_1075);
nand U1588 (N_1588,N_406,In_2458);
xnor U1589 (N_1589,In_2852,N_1089);
nor U1590 (N_1590,In_2324,In_1538);
nand U1591 (N_1591,N_879,In_387);
and U1592 (N_1592,In_1735,In_2917);
or U1593 (N_1593,N_1037,N_603);
xnor U1594 (N_1594,In_2550,N_339);
xor U1595 (N_1595,N_166,In_529);
nor U1596 (N_1596,In_1650,N_12);
or U1597 (N_1597,In_157,In_1378);
nor U1598 (N_1598,N_11,In_392);
xor U1599 (N_1599,In_2281,In_1792);
nand U1600 (N_1600,In_1289,N_920);
nor U1601 (N_1601,In_852,In_2289);
nand U1602 (N_1602,In_1070,In_457);
and U1603 (N_1603,N_1144,N_1197);
or U1604 (N_1604,In_2010,In_1112);
and U1605 (N_1605,In_555,N_1152);
nor U1606 (N_1606,N_911,N_130);
xnor U1607 (N_1607,In_2957,N_286);
or U1608 (N_1608,N_1119,In_1394);
and U1609 (N_1609,N_522,N_1066);
and U1610 (N_1610,In_2444,N_944);
nand U1611 (N_1611,N_968,N_1179);
or U1612 (N_1612,N_530,N_648);
nand U1613 (N_1613,N_936,In_2944);
and U1614 (N_1614,N_800,N_317);
or U1615 (N_1615,N_294,In_2539);
nor U1616 (N_1616,In_413,N_1150);
nand U1617 (N_1617,N_559,N_812);
and U1618 (N_1618,N_100,N_809);
nor U1619 (N_1619,N_112,N_505);
nor U1620 (N_1620,In_1985,In_2831);
nand U1621 (N_1621,N_661,N_528);
xor U1622 (N_1622,In_2972,In_686);
nand U1623 (N_1623,In_667,In_2276);
nor U1624 (N_1624,N_220,In_1283);
nor U1625 (N_1625,In_1747,N_979);
nor U1626 (N_1626,In_1153,N_46);
nor U1627 (N_1627,N_727,In_2169);
xnor U1628 (N_1628,N_941,In_150);
nor U1629 (N_1629,N_417,N_602);
nand U1630 (N_1630,In_1220,In_2328);
nor U1631 (N_1631,N_1189,N_821);
or U1632 (N_1632,N_248,In_1853);
xnor U1633 (N_1633,In_715,N_766);
and U1634 (N_1634,In_1846,In_2088);
xnor U1635 (N_1635,N_35,N_1033);
and U1636 (N_1636,In_351,N_1095);
nand U1637 (N_1637,N_107,In_220);
nand U1638 (N_1638,N_667,N_894);
and U1639 (N_1639,In_311,N_1191);
and U1640 (N_1640,In_301,In_1288);
or U1641 (N_1641,In_209,N_833);
nor U1642 (N_1642,N_554,In_970);
nor U1643 (N_1643,N_269,N_16);
nor U1644 (N_1644,In_1910,In_430);
or U1645 (N_1645,N_813,N_550);
xor U1646 (N_1646,N_1015,In_1545);
xor U1647 (N_1647,N_115,In_1626);
and U1648 (N_1648,N_574,N_346);
nand U1649 (N_1649,In_728,In_1256);
xnor U1650 (N_1650,In_147,N_392);
and U1651 (N_1651,In_2312,N_739);
and U1652 (N_1652,N_932,In_1246);
nand U1653 (N_1653,In_300,N_756);
nor U1654 (N_1654,N_726,In_2752);
nor U1655 (N_1655,N_751,N_109);
or U1656 (N_1656,N_960,N_819);
nand U1657 (N_1657,In_1065,N_1048);
nor U1658 (N_1658,N_918,In_2434);
nor U1659 (N_1659,In_2439,N_337);
or U1660 (N_1660,N_368,N_1081);
nor U1661 (N_1661,N_1044,N_516);
or U1662 (N_1662,In_1088,N_794);
and U1663 (N_1663,In_420,N_185);
xnor U1664 (N_1664,N_1176,N_1149);
nand U1665 (N_1665,N_725,N_0);
or U1666 (N_1666,In_2465,In_2211);
or U1667 (N_1667,N_121,In_2339);
nand U1668 (N_1668,In_2294,In_797);
and U1669 (N_1669,N_31,In_663);
xor U1670 (N_1670,N_863,In_2378);
and U1671 (N_1671,N_242,In_2182);
nor U1672 (N_1672,N_939,In_561);
xnor U1673 (N_1673,N_644,In_1374);
xnor U1674 (N_1674,In_2754,In_1597);
xnor U1675 (N_1675,N_815,In_1265);
and U1676 (N_1676,In_2605,In_2504);
nor U1677 (N_1677,N_1184,N_525);
nand U1678 (N_1678,In_2907,In_2703);
xor U1679 (N_1679,In_137,N_391);
or U1680 (N_1680,In_843,In_2132);
nor U1681 (N_1681,N_713,In_1859);
and U1682 (N_1682,In_2893,In_88);
nor U1683 (N_1683,In_973,N_641);
or U1684 (N_1684,In_546,N_44);
nor U1685 (N_1685,In_2807,N_599);
xnor U1686 (N_1686,In_1512,In_553);
and U1687 (N_1687,N_836,In_1475);
nor U1688 (N_1688,N_605,N_95);
nor U1689 (N_1689,In_810,In_2154);
nand U1690 (N_1690,In_121,N_425);
and U1691 (N_1691,N_1042,In_10);
nor U1692 (N_1692,N_788,N_1140);
or U1693 (N_1693,In_344,N_92);
xor U1694 (N_1694,N_962,N_645);
xnor U1695 (N_1695,In_2742,In_1110);
or U1696 (N_1696,In_2724,In_1410);
and U1697 (N_1697,N_235,In_1061);
nand U1698 (N_1698,In_103,In_1408);
nand U1699 (N_1699,In_475,N_883);
xnor U1700 (N_1700,N_571,In_1617);
nand U1701 (N_1701,In_1327,N_1004);
nand U1702 (N_1702,In_1607,N_973);
nand U1703 (N_1703,In_1808,N_122);
nor U1704 (N_1704,In_353,N_1070);
nor U1705 (N_1705,In_1219,In_2065);
nand U1706 (N_1706,In_165,In_1193);
and U1707 (N_1707,In_2926,In_548);
xnor U1708 (N_1708,N_1041,N_1098);
xor U1709 (N_1709,In_2032,N_950);
and U1710 (N_1710,N_810,In_753);
nor U1711 (N_1711,N_37,N_1068);
xnor U1712 (N_1712,In_2099,N_689);
and U1713 (N_1713,N_963,In_2565);
nand U1714 (N_1714,N_707,N_908);
nand U1715 (N_1715,In_1828,N_732);
nor U1716 (N_1716,In_1979,N_970);
or U1717 (N_1717,In_2810,N_267);
or U1718 (N_1718,N_634,N_474);
or U1719 (N_1719,In_1609,In_1163);
or U1720 (N_1720,N_1064,In_1490);
or U1721 (N_1721,N_1035,N_1028);
nand U1722 (N_1722,In_281,In_2186);
xor U1723 (N_1723,In_2839,N_1046);
or U1724 (N_1724,N_626,In_1616);
and U1725 (N_1725,In_1781,In_1296);
or U1726 (N_1726,In_1,In_640);
and U1727 (N_1727,In_2044,In_79);
nor U1728 (N_1728,In_1048,N_569);
xor U1729 (N_1729,In_2487,In_1130);
nand U1730 (N_1730,In_120,In_740);
and U1731 (N_1731,N_897,N_951);
nand U1732 (N_1732,In_1878,N_551);
or U1733 (N_1733,N_1063,In_163);
nor U1734 (N_1734,In_655,N_393);
nor U1735 (N_1735,N_167,N_332);
and U1736 (N_1736,N_679,In_1138);
nor U1737 (N_1737,N_175,In_981);
xnor U1738 (N_1738,In_2549,N_91);
xor U1739 (N_1739,In_2195,In_2404);
xor U1740 (N_1740,N_814,N_1196);
or U1741 (N_1741,N_227,In_2510);
nand U1742 (N_1742,In_2607,In_1636);
xor U1743 (N_1743,N_799,In_604);
or U1744 (N_1744,In_246,In_628);
and U1745 (N_1745,In_1832,N_915);
and U1746 (N_1746,In_2243,N_688);
xor U1747 (N_1747,In_2989,N_1107);
nor U1748 (N_1748,N_910,N_805);
or U1749 (N_1749,In_1037,In_2577);
or U1750 (N_1750,N_229,N_752);
xnor U1751 (N_1751,N_600,In_2191);
nand U1752 (N_1752,N_356,N_338);
xor U1753 (N_1753,In_989,In_883);
nand U1754 (N_1754,In_1295,N_624);
nand U1755 (N_1755,N_999,In_170);
nand U1756 (N_1756,In_831,N_140);
nor U1757 (N_1757,N_1193,N_838);
nor U1758 (N_1758,N_287,N_696);
or U1759 (N_1759,In_2362,N_983);
nand U1760 (N_1760,In_1762,In_860);
or U1761 (N_1761,In_795,In_2481);
nor U1762 (N_1762,In_223,N_926);
and U1763 (N_1763,N_947,In_48);
xnor U1764 (N_1764,In_2682,In_1105);
xor U1765 (N_1765,N_1034,In_1870);
and U1766 (N_1766,In_290,In_135);
and U1767 (N_1767,In_2201,In_2016);
nor U1768 (N_1768,In_611,In_63);
or U1769 (N_1769,In_2408,N_218);
nor U1770 (N_1770,N_646,N_957);
or U1771 (N_1771,N_4,In_2857);
or U1772 (N_1772,In_2840,In_255);
nand U1773 (N_1773,N_1093,N_784);
xor U1774 (N_1774,In_1212,N_890);
and U1775 (N_1775,N_680,N_636);
or U1776 (N_1776,N_325,N_903);
and U1777 (N_1777,In_2137,N_997);
or U1778 (N_1778,In_2615,N_631);
and U1779 (N_1779,In_929,In_2171);
xor U1780 (N_1780,N_224,In_2725);
nor U1781 (N_1781,N_349,N_1113);
nor U1782 (N_1782,In_1232,N_759);
nor U1783 (N_1783,N_466,In_618);
xor U1784 (N_1784,N_658,N_721);
or U1785 (N_1785,In_1349,N_637);
and U1786 (N_1786,N_1114,N_542);
and U1787 (N_1787,N_457,In_653);
nand U1788 (N_1788,In_83,In_2083);
xor U1789 (N_1789,N_653,N_1192);
nor U1790 (N_1790,N_1117,N_210);
xor U1791 (N_1791,N_940,N_1049);
nand U1792 (N_1792,In_1949,In_2662);
nand U1793 (N_1793,N_241,N_891);
nor U1794 (N_1794,N_1056,N_1170);
and U1795 (N_1795,In_1460,In_2770);
nand U1796 (N_1796,In_1784,In_758);
nand U1797 (N_1797,N_820,N_1039);
nand U1798 (N_1798,In_369,In_2830);
nand U1799 (N_1799,In_95,N_1128);
or U1800 (N_1800,In_1311,N_1446);
nor U1801 (N_1801,In_2826,N_1040);
xnor U1802 (N_1802,N_1723,N_1518);
xor U1803 (N_1803,N_1177,In_2173);
xor U1804 (N_1804,N_1231,N_1654);
and U1805 (N_1805,N_270,N_1648);
nand U1806 (N_1806,N_280,N_1398);
nand U1807 (N_1807,In_1143,N_501);
and U1808 (N_1808,In_1274,In_2336);
nand U1809 (N_1809,In_1485,N_48);
or U1810 (N_1810,N_1689,N_1526);
nor U1811 (N_1811,In_1113,N_470);
and U1812 (N_1812,In_596,N_477);
nor U1813 (N_1813,N_1343,N_1366);
nand U1814 (N_1814,N_827,N_1705);
xor U1815 (N_1815,N_1312,N_1625);
or U1816 (N_1816,N_1590,N_1523);
xor U1817 (N_1817,N_1609,N_1477);
nand U1818 (N_1818,In_1011,N_709);
nand U1819 (N_1819,In_562,N_191);
nand U1820 (N_1820,In_2049,N_1651);
or U1821 (N_1821,N_639,N_1618);
xnor U1822 (N_1822,N_1473,N_1588);
nor U1823 (N_1823,N_621,N_1021);
or U1824 (N_1824,In_2843,In_118);
nand U1825 (N_1825,N_1229,N_854);
xor U1826 (N_1826,N_533,N_1327);
nor U1827 (N_1827,N_780,N_1698);
and U1828 (N_1828,In_422,N_1574);
xnor U1829 (N_1829,N_1454,N_1707);
xnor U1830 (N_1830,In_1463,N_1345);
and U1831 (N_1831,N_1591,In_2115);
and U1832 (N_1832,N_1415,N_14);
or U1833 (N_1833,N_757,In_2780);
nand U1834 (N_1834,N_1778,In_1240);
nand U1835 (N_1835,N_1687,In_1756);
nand U1836 (N_1836,N_1764,In_510);
or U1837 (N_1837,N_1284,N_464);
or U1838 (N_1838,N_1350,N_1212);
nor U1839 (N_1839,N_1727,N_1674);
or U1840 (N_1840,In_1532,N_1369);
or U1841 (N_1841,N_972,N_523);
and U1842 (N_1842,N_1268,In_1466);
nand U1843 (N_1843,N_575,N_73);
nand U1844 (N_1844,N_1430,N_1391);
xnor U1845 (N_1845,In_2126,N_1455);
or U1846 (N_1846,N_1565,In_324);
nand U1847 (N_1847,N_856,N_1308);
nor U1848 (N_1848,N_1554,In_2141);
nor U1849 (N_1849,N_1216,N_563);
nand U1850 (N_1850,N_1213,In_102);
nand U1851 (N_1851,N_283,N_1669);
nor U1852 (N_1852,N_1600,N_657);
and U1853 (N_1853,N_1494,N_1384);
xor U1854 (N_1854,In_398,N_837);
xnor U1855 (N_1855,N_1346,N_1576);
or U1856 (N_1856,N_1630,In_2571);
and U1857 (N_1857,In_427,N_1639);
nor U1858 (N_1858,N_1797,N_754);
nand U1859 (N_1859,N_1278,N_1564);
nor U1860 (N_1860,In_783,N_1675);
nor U1861 (N_1861,In_1509,In_247);
and U1862 (N_1862,N_1791,N_1058);
or U1863 (N_1863,In_1881,N_1386);
and U1864 (N_1864,In_2187,N_1463);
and U1865 (N_1865,N_1143,N_1465);
nor U1866 (N_1866,In_502,In_2311);
xnor U1867 (N_1867,N_1380,N_1772);
or U1868 (N_1868,N_1251,N_1664);
nor U1869 (N_1869,N_1627,N_1724);
nand U1870 (N_1870,N_831,N_1298);
nand U1871 (N_1871,N_1241,In_2419);
nand U1872 (N_1872,N_169,N_1302);
nor U1873 (N_1873,N_1317,N_1045);
xor U1874 (N_1874,N_1718,In_377);
xnor U1875 (N_1875,N_1426,N_1410);
nor U1876 (N_1876,N_845,N_1156);
and U1877 (N_1877,In_976,N_1746);
nor U1878 (N_1878,N_1408,N_1014);
or U1879 (N_1879,N_1692,N_1349);
or U1880 (N_1880,In_395,N_1657);
nor U1881 (N_1881,N_1264,N_178);
nor U1882 (N_1882,N_1626,N_1183);
xnor U1883 (N_1883,N_1167,N_1555);
nand U1884 (N_1884,N_318,In_2297);
nand U1885 (N_1885,N_1782,N_1205);
or U1886 (N_1886,In_139,N_1645);
or U1887 (N_1887,N_1484,In_1821);
and U1888 (N_1888,N_1666,In_0);
or U1889 (N_1889,N_1047,N_1406);
and U1890 (N_1890,N_1320,N_1173);
nand U1891 (N_1891,N_1700,N_1684);
xnor U1892 (N_1892,N_1153,N_1291);
and U1893 (N_1893,N_1720,N_1572);
xor U1894 (N_1894,N_1530,N_1221);
nand U1895 (N_1895,N_1563,N_1003);
nand U1896 (N_1896,In_1391,N_1315);
and U1897 (N_1897,N_1510,N_1799);
nand U1898 (N_1898,N_1597,In_679);
or U1899 (N_1899,In_1666,N_102);
or U1900 (N_1900,N_1751,N_1239);
or U1901 (N_1901,In_2206,N_628);
or U1902 (N_1902,N_494,N_1339);
nand U1903 (N_1903,N_1631,N_1253);
and U1904 (N_1904,In_535,In_2985);
and U1905 (N_1905,N_1360,N_290);
nor U1906 (N_1906,N_1469,N_1295);
nand U1907 (N_1907,In_1546,In_1794);
or U1908 (N_1908,N_1636,N_1506);
xnor U1909 (N_1909,N_764,N_1100);
nor U1910 (N_1910,N_1441,In_1816);
xor U1911 (N_1911,N_266,N_1442);
xnor U1912 (N_1912,N_1558,N_986);
xnor U1913 (N_1913,N_949,N_1303);
nand U1914 (N_1914,N_1557,N_1712);
nor U1915 (N_1915,In_168,N_1616);
nand U1916 (N_1916,In_1149,N_1443);
nor U1917 (N_1917,In_2136,N_1235);
nand U1918 (N_1918,N_1580,N_1529);
or U1919 (N_1919,N_616,N_1353);
nor U1920 (N_1920,N_1491,N_928);
nand U1921 (N_1921,N_412,In_2743);
nor U1922 (N_1922,In_2707,N_1781);
xnor U1923 (N_1923,N_1656,In_708);
xnor U1924 (N_1924,N_1767,In_2961);
and U1925 (N_1925,In_453,In_2159);
or U1926 (N_1926,N_1261,N_40);
nor U1927 (N_1927,In_2021,In_644);
nand U1928 (N_1928,N_664,In_161);
nor U1929 (N_1929,N_1660,N_364);
and U1930 (N_1930,N_987,N_1123);
nor U1931 (N_1931,N_1532,N_1417);
xor U1932 (N_1932,N_1749,N_98);
nor U1933 (N_1933,N_1071,In_401);
and U1934 (N_1934,N_803,N_1610);
and U1935 (N_1935,N_366,N_1544);
nor U1936 (N_1936,N_330,In_1147);
nand U1937 (N_1937,N_1482,In_1980);
or U1938 (N_1938,N_1644,N_649);
xor U1939 (N_1939,N_1274,N_1503);
nor U1940 (N_1940,In_1127,N_1581);
nor U1941 (N_1941,N_1762,N_168);
nor U1942 (N_1942,N_1632,N_119);
nand U1943 (N_1943,N_451,N_1560);
or U1944 (N_1944,In_2251,In_1833);
or U1945 (N_1945,N_1328,N_1541);
nand U1946 (N_1946,N_1290,N_808);
nand U1947 (N_1947,In_2986,In_2689);
nor U1948 (N_1948,N_1445,N_678);
and U1949 (N_1949,N_1435,N_1351);
and U1950 (N_1950,In_1396,N_153);
and U1951 (N_1951,N_924,In_2965);
or U1952 (N_1952,N_1393,N_578);
and U1953 (N_1953,N_1138,N_454);
and U1954 (N_1954,N_758,N_793);
xor U1955 (N_1955,N_38,N_1691);
nor U1956 (N_1956,N_1524,In_730);
or U1957 (N_1957,N_1561,N_1628);
or U1958 (N_1958,N_371,In_1203);
and U1959 (N_1959,N_990,N_1200);
xnor U1960 (N_1960,N_76,N_760);
xnor U1961 (N_1961,N_1759,N_798);
nor U1962 (N_1962,In_2668,In_1824);
and U1963 (N_1963,N_1228,N_976);
nor U1964 (N_1964,N_823,N_213);
or U1965 (N_1965,N_10,In_2657);
xnor U1966 (N_1966,N_1259,N_1232);
nor U1967 (N_1967,N_866,In_2977);
or U1968 (N_1968,N_335,N_1275);
nand U1969 (N_1969,In_2569,N_1181);
xnor U1970 (N_1970,N_1450,N_1162);
nor U1971 (N_1971,N_324,N_1059);
or U1972 (N_1972,N_1358,N_304);
xor U1973 (N_1973,N_633,N_1622);
xor U1974 (N_1974,In_587,N_1104);
xor U1975 (N_1975,N_1008,N_1378);
or U1976 (N_1976,N_1354,N_1605);
or U1977 (N_1977,In_2499,N_1739);
xnor U1978 (N_1978,N_1407,In_2273);
or U1979 (N_1979,In_1071,N_1240);
xor U1980 (N_1980,N_619,N_1334);
nand U1981 (N_1981,In_158,N_1548);
or U1982 (N_1982,N_1571,In_763);
nor U1983 (N_1983,N_1699,In_1696);
or U1984 (N_1984,N_1783,N_1753);
xnor U1985 (N_1985,N_1055,N_848);
nor U1986 (N_1986,N_1531,In_2735);
nand U1987 (N_1987,In_1703,In_2919);
xnor U1988 (N_1988,N_1433,N_1313);
or U1989 (N_1989,In_2693,N_710);
nand U1990 (N_1990,N_1215,N_1775);
and U1991 (N_1991,N_1282,N_699);
and U1992 (N_1992,N_1245,N_1796);
and U1993 (N_1993,In_2680,N_1257);
nand U1994 (N_1994,N_1696,N_1270);
xnor U1995 (N_1995,N_1538,N_1757);
and U1996 (N_1996,N_1652,In_78);
nor U1997 (N_1997,In_815,N_996);
nor U1998 (N_1998,N_401,In_709);
and U1999 (N_1999,In_1114,N_1451);
or U2000 (N_2000,N_326,N_711);
nor U2001 (N_2001,N_1734,N_1731);
nor U2002 (N_2002,N_174,N_1383);
nor U2003 (N_2003,N_1583,In_696);
nor U2004 (N_2004,N_1462,N_1756);
or U2005 (N_2005,In_2055,In_1080);
and U2006 (N_2006,In_1150,N_828);
nand U2007 (N_2007,N_1311,N_1766);
xor U2008 (N_2008,N_1701,N_1080);
nand U2009 (N_2009,In_1481,N_1363);
or U2010 (N_2010,In_2761,In_1155);
xnor U2011 (N_2011,N_1508,N_1647);
xnor U2012 (N_2012,N_1516,N_327);
nor U2013 (N_2013,In_1777,In_788);
xor U2014 (N_2014,N_1695,N_1722);
and U2015 (N_2015,N_85,N_1122);
and U2016 (N_2016,N_791,N_1535);
and U2017 (N_2017,N_1403,In_2916);
and U2018 (N_2018,In_505,N_1287);
and U2019 (N_2019,N_1348,N_1649);
and U2020 (N_2020,N_994,N_880);
or U2021 (N_2021,N_1195,In_1907);
or U2022 (N_2022,In_1285,N_1394);
xor U2023 (N_2023,In_1079,In_2204);
nand U2024 (N_2024,N_1083,N_625);
nor U2025 (N_2025,N_1390,N_1533);
and U2026 (N_2026,N_1534,N_1422);
nand U2027 (N_2027,N_385,N_716);
nand U2028 (N_2028,N_1480,N_1146);
nor U2029 (N_2029,N_1062,In_501);
nor U2030 (N_2030,N_1305,In_2524);
and U2031 (N_2031,N_1211,N_922);
nand U2032 (N_2032,N_1567,N_1357);
or U2033 (N_2033,N_1721,N_1568);
nand U2034 (N_2034,N_1713,N_1151);
xor U2035 (N_2035,N_30,N_1769);
or U2036 (N_2036,N_1013,N_1643);
xnor U2037 (N_2037,N_1027,In_1092);
or U2038 (N_2038,N_902,N_1697);
and U2039 (N_2039,In_514,In_2143);
and U2040 (N_2040,N_1329,In_794);
nor U2041 (N_2041,N_1234,N_1355);
or U2042 (N_2042,N_1362,N_1220);
nand U2043 (N_2043,N_1111,N_1418);
nand U2044 (N_2044,N_1481,N_443);
xnor U2045 (N_2045,N_134,N_1594);
xnor U2046 (N_2046,N_683,N_1467);
and U2047 (N_2047,N_1401,N_1776);
nand U2048 (N_2048,N_1084,N_1488);
nor U2049 (N_2049,N_1742,In_2639);
nor U2050 (N_2050,N_1364,In_2875);
or U2051 (N_2051,N_1615,N_956);
or U2052 (N_2052,In_2245,N_1758);
nor U2053 (N_2053,In_2172,N_1780);
or U2054 (N_2054,N_1760,In_2879);
nor U2055 (N_2055,N_1326,N_1341);
nor U2056 (N_2056,N_1785,N_655);
nor U2057 (N_2057,N_1595,N_1164);
or U2058 (N_2058,In_917,In_2863);
and U2059 (N_2059,In_1456,N_1166);
and U2060 (N_2060,In_906,N_1405);
xnor U2061 (N_2061,N_905,N_1589);
and U2062 (N_2062,N_937,N_1793);
nor U2063 (N_2063,In_2153,N_1585);
nor U2064 (N_2064,N_1703,N_844);
and U2065 (N_2065,N_1202,N_1520);
xor U2066 (N_2066,In_2828,N_1543);
nor U2067 (N_2067,N_1297,In_2758);
nand U2068 (N_2068,N_1365,N_1267);
nand U2069 (N_2069,In_1354,N_1206);
or U2070 (N_2070,In_2435,N_1489);
and U2071 (N_2071,In_848,N_877);
or U2072 (N_2072,N_942,N_1009);
or U2073 (N_2073,In_1727,N_486);
and U2074 (N_2074,N_1269,N_834);
nand U2075 (N_2075,In_365,N_1310);
nor U2076 (N_2076,In_1188,N_675);
nand U2077 (N_2077,N_405,N_1225);
or U2078 (N_2078,In_425,N_1688);
and U2079 (N_2079,N_1659,N_1322);
and U2080 (N_2080,In_1897,N_1210);
nand U2081 (N_2081,N_1468,In_1685);
nor U2082 (N_2082,N_755,N_964);
or U2083 (N_2083,N_1256,N_1069);
and U2084 (N_2084,N_1740,In_469);
nand U2085 (N_2085,N_1500,N_1515);
nor U2086 (N_2086,N_1237,N_1280);
nand U2087 (N_2087,In_183,In_273);
nand U2088 (N_2088,N_1036,In_1010);
xor U2089 (N_2089,N_1573,In_2809);
nand U2090 (N_2090,N_1372,N_1301);
or U2091 (N_2091,N_1582,In_807);
nand U2092 (N_2092,N_1768,N_308);
nand U2093 (N_2093,N_1331,N_1175);
and U2094 (N_2094,N_1371,N_1736);
or U2095 (N_2095,In_2353,N_635);
xnor U2096 (N_2096,N_200,N_695);
or U2097 (N_2097,N_1788,In_1868);
or U2098 (N_2098,N_567,In_2686);
and U2099 (N_2099,N_1686,N_1620);
nor U2100 (N_2100,N_1677,N_1335);
nand U2101 (N_2101,In_698,In_211);
and U2102 (N_2102,In_2529,N_1725);
and U2103 (N_2103,In_1388,N_1710);
or U2104 (N_2104,N_1763,N_1294);
and U2105 (N_2105,N_1624,N_1528);
xor U2106 (N_2106,N_1356,In_1973);
xor U2107 (N_2107,N_1377,N_1293);
xor U2108 (N_2108,In_586,In_2359);
xnor U2109 (N_2109,N_1425,N_1337);
or U2110 (N_2110,In_1967,N_1409);
nand U2111 (N_2111,In_2938,N_943);
and U2112 (N_2112,In_2383,N_807);
or U2113 (N_2113,In_1991,N_1309);
xnor U2114 (N_2114,In_1093,N_1498);
nor U2115 (N_2115,N_506,N_1743);
nand U2116 (N_2116,N_1683,N_1227);
or U2117 (N_2117,N_1487,N_1741);
and U2118 (N_2118,In_771,N_1599);
or U2119 (N_2119,N_1411,In_330);
and U2120 (N_2120,In_960,N_1396);
xor U2121 (N_2121,N_1217,In_2403);
xnor U2122 (N_2122,In_1592,N_1545);
nand U2123 (N_2123,N_1733,In_2381);
nor U2124 (N_2124,N_1655,In_575);
xor U2125 (N_2125,In_82,N_1562);
nand U2126 (N_2126,N_1226,In_1340);
nand U2127 (N_2127,In_1612,N_1613);
and U2128 (N_2128,N_1476,N_607);
nand U2129 (N_2129,N_1431,In_766);
nor U2130 (N_2130,In_1494,N_515);
and U2131 (N_2131,N_1621,In_2015);
nand U2132 (N_2132,N_919,In_966);
or U2133 (N_2133,N_399,In_2732);
or U2134 (N_2134,In_2656,N_1457);
or U2135 (N_2135,N_1490,N_1499);
nand U2136 (N_2136,N_1133,N_1324);
nand U2137 (N_2137,N_1249,In_203);
xor U2138 (N_2138,N_1798,N_1051);
nor U2139 (N_2139,N_1109,N_1608);
nand U2140 (N_2140,N_1230,N_1629);
nor U2141 (N_2141,N_692,N_1316);
or U2142 (N_2142,N_1273,N_1464);
or U2143 (N_2143,N_1744,N_887);
and U2144 (N_2144,N_1244,N_1512);
nand U2145 (N_2145,In_1922,N_717);
nor U2146 (N_2146,N_1266,N_1436);
and U2147 (N_2147,N_1429,In_2954);
nor U2148 (N_2148,N_1134,In_400);
or U2149 (N_2149,N_1587,In_2205);
nand U2150 (N_2150,N_298,In_1755);
and U2151 (N_2151,N_1250,In_64);
nor U2152 (N_2152,N_1550,N_790);
nand U2153 (N_2153,In_2767,In_2420);
xor U2154 (N_2154,N_1392,N_1204);
nand U2155 (N_2155,N_1243,N_1761);
xor U2156 (N_2156,In_1584,In_1805);
nand U2157 (N_2157,N_1288,N_1501);
and U2158 (N_2158,N_504,N_1755);
xor U2159 (N_2159,N_1646,N_465);
xor U2160 (N_2160,N_694,N_245);
nand U2161 (N_2161,In_1389,N_1252);
nand U2162 (N_2162,N_1601,N_1460);
or U2163 (N_2163,N_1728,N_1527);
nor U2164 (N_2164,N_1385,N_1607);
nor U2165 (N_2165,N_1057,N_1285);
and U2166 (N_2166,N_1777,N_1502);
and U2167 (N_2167,N_1402,In_2337);
xnor U2168 (N_2168,In_2906,N_1258);
and U2169 (N_2169,In_2492,N_1726);
or U2170 (N_2170,N_1786,N_558);
or U2171 (N_2171,N_1779,In_2900);
nor U2172 (N_2172,N_389,N_1547);
and U2173 (N_2173,In_1862,N_1413);
xor U2174 (N_2174,N_1614,N_398);
nand U2175 (N_2175,In_2482,N_1276);
xor U2176 (N_2176,N_1399,In_1467);
nor U2177 (N_2177,In_592,N_1711);
and U2178 (N_2178,N_1787,N_1670);
nand U2179 (N_2179,N_1770,N_1611);
or U2180 (N_2180,N_686,N_125);
and U2181 (N_2181,N_1690,N_1794);
or U2182 (N_2182,In_1938,In_2951);
or U2183 (N_2183,In_645,N_1546);
or U2184 (N_2184,N_1373,In_1056);
nor U2185 (N_2185,In_2692,N_1139);
nor U2186 (N_2186,N_1419,N_1340);
nor U2187 (N_2187,N_343,N_1635);
and U2188 (N_2188,N_981,N_1246);
xor U2189 (N_2189,N_1077,N_1002);
nor U2190 (N_2190,N_1236,N_822);
xnor U2191 (N_2191,N_1172,In_1725);
nand U2192 (N_2192,N_777,In_1444);
nand U2193 (N_2193,In_748,N_1024);
or U2194 (N_2194,N_875,N_1072);
xor U2195 (N_2195,N_1709,N_1495);
nand U2196 (N_2196,In_268,N_1129);
or U2197 (N_2197,N_1159,In_1136);
nor U2198 (N_2198,N_1306,N_1199);
xnor U2199 (N_2199,N_1368,N_1592);
and U2200 (N_2200,N_83,N_1325);
nor U2201 (N_2201,N_995,N_1792);
or U2202 (N_2202,In_1958,N_1260);
nand U2203 (N_2203,In_1522,N_1388);
xnor U2204 (N_2204,N_1207,N_1549);
nand U2205 (N_2205,N_1479,N_1679);
and U2206 (N_2206,In_613,In_200);
and U2207 (N_2207,N_1729,N_1474);
nor U2208 (N_2208,N_1158,N_1745);
or U2209 (N_2209,N_1208,N_1662);
and U2210 (N_2210,N_1536,In_1473);
xor U2211 (N_2211,N_1182,N_460);
nor U2212 (N_2212,N_1539,N_1747);
nand U2213 (N_2213,In_2326,In_1310);
nand U2214 (N_2214,N_1540,N_749);
xnor U2215 (N_2215,In_864,N_1606);
and U2216 (N_2216,N_1444,N_1404);
or U2217 (N_2217,N_462,N_1420);
xnor U2218 (N_2218,In_2338,N_906);
or U2219 (N_2219,N_1586,N_1359);
nor U2220 (N_2220,N_110,N_1319);
xor U2221 (N_2221,N_1507,N_1642);
nand U2222 (N_2222,N_1185,N_913);
nand U2223 (N_2223,N_437,N_1314);
nor U2224 (N_2224,N_1719,N_1338);
or U2225 (N_2225,N_61,N_1209);
xnor U2226 (N_2226,N_1292,N_691);
nor U2227 (N_2227,In_2641,N_1593);
and U2228 (N_2228,In_1669,N_1453);
xor U2229 (N_2229,N_1485,N_1321);
and U2230 (N_2230,In_1229,N_886);
and U2231 (N_2231,In_2296,In_517);
or U2232 (N_2232,N_1638,N_1578);
nor U2233 (N_2233,In_1883,N_1559);
nor U2234 (N_2234,N_1222,In_2827);
xnor U2235 (N_2235,N_1738,N_1277);
nor U2236 (N_2236,In_455,N_839);
nand U2237 (N_2237,N_1784,N_1421);
xnor U2238 (N_2238,N_1566,N_1575);
nand U2239 (N_2239,In_1565,N_1569);
nor U2240 (N_2240,N_1716,N_1704);
nand U2241 (N_2241,N_510,N_573);
xor U2242 (N_2242,N_1344,N_1693);
or U2243 (N_2243,N_1412,N_1737);
or U2244 (N_2244,N_1434,N_1505);
or U2245 (N_2245,N_1437,N_548);
nor U2246 (N_2246,In_1472,In_750);
nor U2247 (N_2247,In_1359,N_1428);
and U2248 (N_2248,N_1459,N_139);
xor U2249 (N_2249,N_929,In_1511);
nand U2250 (N_2250,In_2940,In_2666);
xnor U2251 (N_2251,N_23,In_279);
xor U2252 (N_2252,N_1511,N_768);
and U2253 (N_2253,N_1323,N_1203);
nor U2254 (N_2254,N_1281,In_2821);
nand U2255 (N_2255,N_1735,N_1714);
xnor U2256 (N_2256,N_1265,In_1986);
and U2257 (N_2257,N_1382,In_1307);
nor U2258 (N_2258,N_1336,N_1577);
nand U2259 (N_2259,N_1414,N_612);
and U2260 (N_2260,In_2896,In_1152);
nor U2261 (N_2261,In_1443,N_348);
and U2262 (N_2262,In_1889,N_702);
or U2263 (N_2263,N_1078,In_1581);
nor U2264 (N_2264,N_1748,N_703);
or U2265 (N_2265,N_1765,N_1771);
xor U2266 (N_2266,In_2669,N_1774);
and U2267 (N_2267,In_953,In_2667);
and U2268 (N_2268,N_1079,In_466);
nor U2269 (N_2269,N_1486,N_1397);
or U2270 (N_2270,N_1090,In_1734);
xnor U2271 (N_2271,In_2256,N_1283);
xor U2272 (N_2272,N_221,N_620);
or U2273 (N_2273,N_1717,N_1438);
or U2274 (N_2274,N_238,N_933);
xnor U2275 (N_2275,N_1286,N_1579);
xor U2276 (N_2276,In_700,N_930);
xor U2277 (N_2277,N_1376,N_622);
xnor U2278 (N_2278,N_1663,N_1634);
nand U2279 (N_2279,In_2372,N_984);
and U2280 (N_2280,In_1198,N_1478);
xor U2281 (N_2281,In_1975,N_1423);
nor U2282 (N_2282,N_1458,N_1330);
xor U2283 (N_2283,N_1296,N_1497);
or U2284 (N_2284,N_1026,In_578);
or U2285 (N_2285,In_1707,N_1000);
and U2286 (N_2286,N_1299,N_1472);
nand U2287 (N_2287,N_518,In_342);
and U2288 (N_2288,N_1461,In_664);
xnor U2289 (N_2289,N_1233,N_1790);
or U2290 (N_2290,N_1247,In_2526);
nand U2291 (N_2291,N_1271,N_106);
xor U2292 (N_2292,N_1730,N_1750);
nand U2293 (N_2293,N_1342,In_487);
or U2294 (N_2294,In_1271,N_1676);
nor U2295 (N_2295,N_1381,In_412);
nor U2296 (N_2296,N_580,N_1440);
nand U2297 (N_2297,In_2106,N_1367);
and U2298 (N_2298,In_190,N_1370);
xnor U2299 (N_2299,N_1653,In_798);
nand U2300 (N_2300,N_901,N_1706);
and U2301 (N_2301,N_1773,N_1623);
and U2302 (N_2302,N_1619,N_1604);
or U2303 (N_2303,N_128,N_1682);
or U2304 (N_2304,In_2844,N_923);
nand U2305 (N_2305,N_1242,N_1552);
nor U2306 (N_2306,N_701,In_760);
xnor U2307 (N_2307,N_55,N_1361);
nand U2308 (N_2308,N_1439,N_728);
and U2309 (N_2309,In_2255,N_1395);
xor U2310 (N_2310,In_1519,N_795);
nand U2311 (N_2311,N_1752,N_1374);
and U2312 (N_2312,In_1128,N_1424);
nor U2313 (N_2313,N_697,N_656);
xnor U2314 (N_2314,N_872,In_182);
nor U2315 (N_2315,N_1224,N_1658);
and U2316 (N_2316,N_1633,In_1664);
xor U2317 (N_2317,In_631,N_1254);
nand U2318 (N_2318,In_2448,N_1678);
and U2319 (N_2319,N_1466,In_1459);
nand U2320 (N_2320,N_1214,N_1304);
nand U2321 (N_2321,N_1496,N_1456);
xor U2322 (N_2322,N_660,N_785);
or U2323 (N_2323,N_1671,N_1279);
xor U2324 (N_2324,N_1262,N_1517);
or U2325 (N_2325,N_1617,N_282);
nor U2326 (N_2326,N_1612,N_1665);
xnor U2327 (N_2327,N_1514,N_1272);
and U2328 (N_2328,N_1504,N_1641);
xor U2329 (N_2329,In_2511,N_969);
xnor U2330 (N_2330,In_1896,N_541);
or U2331 (N_2331,N_1219,N_1672);
and U2332 (N_2332,N_1556,N_606);
and U2333 (N_2333,In_804,N_1332);
or U2334 (N_2334,N_829,In_2708);
xnor U2335 (N_2335,N_1513,N_1789);
xor U2336 (N_2336,N_329,In_1400);
nor U2337 (N_2337,In_293,N_295);
nor U2338 (N_2338,In_227,In_1292);
and U2339 (N_2339,N_1448,In_1266);
nor U2340 (N_2340,N_316,In_2103);
nand U2341 (N_2341,N_676,N_1475);
and U2342 (N_2342,N_1432,In_635);
nor U2343 (N_2343,N_1300,N_1525);
and U2344 (N_2344,N_1673,N_1307);
nand U2345 (N_2345,N_1188,N_907);
nor U2346 (N_2346,N_1318,In_34);
and U2347 (N_2347,N_1640,N_303);
nand U2348 (N_2348,In_1799,N_350);
nand U2349 (N_2349,N_1570,N_1650);
or U2350 (N_2350,N_1387,N_1449);
xor U2351 (N_2351,N_1521,N_931);
or U2352 (N_2352,N_1352,N_769);
nand U2353 (N_2353,N_1427,N_1702);
or U2354 (N_2354,N_1795,N_1333);
xnor U2355 (N_2355,In_309,N_671);
xnor U2356 (N_2356,N_1667,N_610);
or U2357 (N_2357,N_1680,In_2034);
nand U2358 (N_2358,N_1248,N_1732);
nor U2359 (N_2359,N_24,N_1542);
xor U2360 (N_2360,N_991,In_129);
and U2361 (N_2361,N_1685,N_706);
nand U2362 (N_2362,In_2352,N_190);
xor U2363 (N_2363,N_313,N_1602);
nor U2364 (N_2364,N_1694,N_781);
nor U2365 (N_2365,N_1010,N_1483);
nand U2366 (N_2366,N_1596,In_317);
xor U2367 (N_2367,N_1637,N_954);
and U2368 (N_2368,In_2600,N_1121);
nand U2369 (N_2369,N_1092,N_508);
or U2370 (N_2370,In_1191,N_1186);
xnor U2371 (N_2371,N_1519,N_1452);
xor U2372 (N_2372,N_1681,N_1551);
nor U2373 (N_2373,N_771,N_1553);
xor U2374 (N_2374,N_1668,In_1495);
xnor U2375 (N_2375,N_1754,N_1603);
and U2376 (N_2376,N_1509,N_1218);
xor U2377 (N_2377,In_495,N_1708);
or U2378 (N_2378,In_2955,N_1584);
or U2379 (N_2379,In_2581,N_1492);
and U2380 (N_2380,In_31,In_35);
and U2381 (N_2381,In_834,N_1471);
nand U2382 (N_2382,N_1537,N_1598);
xor U2383 (N_2383,N_1470,N_1223);
xor U2384 (N_2384,In_704,In_2366);
nand U2385 (N_2385,N_1347,N_1715);
and U2386 (N_2386,N_651,In_1013);
nand U2387 (N_2387,N_1178,N_1661);
xnor U2388 (N_2388,N_1238,In_2644);
xnor U2389 (N_2389,In_1505,N_1263);
and U2390 (N_2390,N_1007,N_1255);
xor U2391 (N_2391,N_672,N_1389);
nand U2392 (N_2392,N_1289,N_1400);
nor U2393 (N_2393,N_623,N_1447);
and U2394 (N_2394,N_1493,N_1416);
xor U2395 (N_2395,N_801,N_1375);
or U2396 (N_2396,N_1379,N_483);
nand U2397 (N_2397,N_1005,In_2717);
nor U2398 (N_2398,N_1201,N_1522);
nand U2399 (N_2399,N_816,N_779);
and U2400 (N_2400,N_2185,N_1963);
xnor U2401 (N_2401,N_2382,N_2242);
or U2402 (N_2402,N_2330,N_1886);
nor U2403 (N_2403,N_2328,N_2055);
xnor U2404 (N_2404,N_2008,N_2016);
or U2405 (N_2405,N_1976,N_2210);
xor U2406 (N_2406,N_2356,N_2072);
nor U2407 (N_2407,N_2252,N_2331);
nor U2408 (N_2408,N_1940,N_2158);
and U2409 (N_2409,N_2159,N_1884);
nor U2410 (N_2410,N_2013,N_1866);
nand U2411 (N_2411,N_1856,N_2049);
nor U2412 (N_2412,N_2094,N_2146);
or U2413 (N_2413,N_2370,N_2206);
nor U2414 (N_2414,N_2324,N_2241);
and U2415 (N_2415,N_2209,N_2216);
and U2416 (N_2416,N_2188,N_2364);
nand U2417 (N_2417,N_1986,N_1810);
or U2418 (N_2418,N_2132,N_1898);
nand U2419 (N_2419,N_2000,N_2021);
and U2420 (N_2420,N_1918,N_2231);
nor U2421 (N_2421,N_2335,N_2054);
and U2422 (N_2422,N_2139,N_2040);
and U2423 (N_2423,N_2162,N_1897);
nand U2424 (N_2424,N_1818,N_2230);
and U2425 (N_2425,N_2124,N_1958);
nor U2426 (N_2426,N_2184,N_1851);
xnor U2427 (N_2427,N_2226,N_2204);
nor U2428 (N_2428,N_1823,N_2061);
or U2429 (N_2429,N_2372,N_1902);
and U2430 (N_2430,N_1879,N_1802);
xnor U2431 (N_2431,N_1867,N_2155);
nor U2432 (N_2432,N_1999,N_2213);
nand U2433 (N_2433,N_2379,N_2098);
nand U2434 (N_2434,N_1968,N_1832);
nor U2435 (N_2435,N_2083,N_2174);
nand U2436 (N_2436,N_2366,N_2079);
or U2437 (N_2437,N_2329,N_2220);
and U2438 (N_2438,N_1801,N_1939);
nor U2439 (N_2439,N_2352,N_2048);
nand U2440 (N_2440,N_1907,N_2166);
or U2441 (N_2441,N_2243,N_1847);
nor U2442 (N_2442,N_2194,N_1857);
nand U2443 (N_2443,N_1949,N_2229);
xnor U2444 (N_2444,N_1874,N_2388);
nor U2445 (N_2445,N_2398,N_1901);
or U2446 (N_2446,N_2037,N_2293);
nor U2447 (N_2447,N_1890,N_2284);
xor U2448 (N_2448,N_2347,N_1861);
or U2449 (N_2449,N_2270,N_2369);
nor U2450 (N_2450,N_1824,N_2300);
and U2451 (N_2451,N_1883,N_2039);
nand U2452 (N_2452,N_2030,N_1915);
nor U2453 (N_2453,N_2365,N_2333);
nor U2454 (N_2454,N_2336,N_1880);
nor U2455 (N_2455,N_1869,N_2321);
and U2456 (N_2456,N_2149,N_1973);
nor U2457 (N_2457,N_2113,N_1935);
xor U2458 (N_2458,N_2097,N_2190);
xnor U2459 (N_2459,N_2322,N_2395);
and U2460 (N_2460,N_2310,N_2092);
nor U2461 (N_2461,N_2325,N_2114);
nor U2462 (N_2462,N_2259,N_2161);
xor U2463 (N_2463,N_2110,N_1909);
xnor U2464 (N_2464,N_1912,N_2002);
xnor U2465 (N_2465,N_2170,N_1905);
nor U2466 (N_2466,N_1971,N_2362);
or U2467 (N_2467,N_1925,N_1894);
nor U2468 (N_2468,N_1955,N_2386);
nand U2469 (N_2469,N_2085,N_2253);
nor U2470 (N_2470,N_2060,N_2344);
nand U2471 (N_2471,N_1953,N_2053);
or U2472 (N_2472,N_1829,N_2116);
xnor U2473 (N_2473,N_2112,N_2311);
xor U2474 (N_2474,N_2232,N_1814);
xnor U2475 (N_2475,N_2339,N_2211);
and U2476 (N_2476,N_2378,N_1854);
nand U2477 (N_2477,N_2014,N_2165);
or U2478 (N_2478,N_1889,N_1822);
nand U2479 (N_2479,N_1908,N_2125);
nor U2480 (N_2480,N_2069,N_2004);
and U2481 (N_2481,N_2217,N_2141);
or U2482 (N_2482,N_2237,N_1828);
xor U2483 (N_2483,N_1930,N_2154);
or U2484 (N_2484,N_2323,N_2240);
and U2485 (N_2485,N_1931,N_1806);
or U2486 (N_2486,N_2319,N_1938);
nand U2487 (N_2487,N_1950,N_2262);
and U2488 (N_2488,N_2168,N_2306);
xor U2489 (N_2489,N_2108,N_1805);
nand U2490 (N_2490,N_1967,N_2144);
nor U2491 (N_2491,N_2373,N_2163);
nand U2492 (N_2492,N_1970,N_2056);
xnor U2493 (N_2493,N_1995,N_2160);
nor U2494 (N_2494,N_2145,N_2228);
or U2495 (N_2495,N_2394,N_2153);
xor U2496 (N_2496,N_1816,N_1996);
and U2497 (N_2497,N_2371,N_2143);
or U2498 (N_2498,N_2199,N_2317);
nor U2499 (N_2499,N_2374,N_2025);
nand U2500 (N_2500,N_2381,N_2179);
nor U2501 (N_2501,N_1927,N_2015);
xor U2502 (N_2502,N_2073,N_2218);
nor U2503 (N_2503,N_2245,N_2180);
or U2504 (N_2504,N_2338,N_2182);
or U2505 (N_2505,N_2051,N_2193);
nand U2506 (N_2506,N_1809,N_2361);
or U2507 (N_2507,N_1992,N_2164);
or U2508 (N_2508,N_2298,N_2263);
or U2509 (N_2509,N_1990,N_2349);
and U2510 (N_2510,N_2266,N_2119);
and U2511 (N_2511,N_1961,N_2215);
xor U2512 (N_2512,N_1933,N_1957);
xnor U2513 (N_2513,N_1875,N_1969);
or U2514 (N_2514,N_2157,N_2063);
xnor U2515 (N_2515,N_1960,N_2387);
nand U2516 (N_2516,N_2358,N_2254);
nand U2517 (N_2517,N_1952,N_2178);
nor U2518 (N_2518,N_1800,N_1864);
nand U2519 (N_2519,N_1946,N_1920);
or U2520 (N_2520,N_1972,N_1951);
or U2521 (N_2521,N_1873,N_2299);
nor U2522 (N_2522,N_2359,N_1811);
or U2523 (N_2523,N_2286,N_2267);
and U2524 (N_2524,N_2005,N_2341);
or U2525 (N_2525,N_2375,N_2227);
nor U2526 (N_2526,N_1845,N_2316);
nor U2527 (N_2527,N_2289,N_2033);
and U2528 (N_2528,N_1819,N_2308);
nand U2529 (N_2529,N_1899,N_2214);
xor U2530 (N_2530,N_2089,N_1944);
xor U2531 (N_2531,N_2244,N_2208);
xor U2532 (N_2532,N_1876,N_2007);
and U2533 (N_2533,N_2292,N_2312);
nor U2534 (N_2534,N_2389,N_2172);
nor U2535 (N_2535,N_2082,N_2340);
nand U2536 (N_2536,N_2169,N_1947);
xor U2537 (N_2537,N_1964,N_1965);
and U2538 (N_2538,N_2280,N_1923);
nor U2539 (N_2539,N_1903,N_2318);
nor U2540 (N_2540,N_1836,N_1926);
nand U2541 (N_2541,N_1917,N_1937);
xnor U2542 (N_2542,N_2360,N_1862);
nand U2543 (N_2543,N_1888,N_1895);
and U2544 (N_2544,N_2044,N_2304);
xor U2545 (N_2545,N_1981,N_1859);
and U2546 (N_2546,N_1842,N_2295);
and U2547 (N_2547,N_2135,N_2057);
and U2548 (N_2548,N_2128,N_2062);
and U2549 (N_2549,N_2121,N_1870);
nor U2550 (N_2550,N_2393,N_2224);
or U2551 (N_2551,N_1966,N_2314);
xor U2552 (N_2552,N_2122,N_2065);
nor U2553 (N_2553,N_1919,N_2384);
and U2554 (N_2554,N_1941,N_2042);
nand U2555 (N_2555,N_1831,N_2271);
and U2556 (N_2556,N_1932,N_2096);
xor U2557 (N_2557,N_1913,N_2134);
nor U2558 (N_2558,N_2029,N_1987);
and U2559 (N_2559,N_2258,N_2235);
xnor U2560 (N_2560,N_2084,N_2222);
nand U2561 (N_2561,N_2183,N_2203);
xor U2562 (N_2562,N_1844,N_2131);
nand U2563 (N_2563,N_2246,N_1893);
and U2564 (N_2564,N_2100,N_2117);
nand U2565 (N_2565,N_2315,N_2207);
nand U2566 (N_2566,N_2279,N_2093);
xnor U2567 (N_2567,N_2177,N_2027);
and U2568 (N_2568,N_2105,N_1858);
or U2569 (N_2569,N_2195,N_2291);
and U2570 (N_2570,N_2354,N_2107);
and U2571 (N_2571,N_2080,N_1882);
nand U2572 (N_2572,N_1834,N_1827);
nor U2573 (N_2573,N_1983,N_2303);
nor U2574 (N_2574,N_2281,N_2038);
xnor U2575 (N_2575,N_1812,N_1978);
or U2576 (N_2576,N_2337,N_2350);
and U2577 (N_2577,N_2377,N_1942);
and U2578 (N_2578,N_2041,N_2301);
nand U2579 (N_2579,N_2383,N_1954);
or U2580 (N_2580,N_2277,N_2020);
nand U2581 (N_2581,N_1928,N_1840);
nand U2582 (N_2582,N_1849,N_2320);
or U2583 (N_2583,N_2081,N_2272);
nor U2584 (N_2584,N_2353,N_2091);
xnor U2585 (N_2585,N_1807,N_1904);
or U2586 (N_2586,N_1977,N_2102);
and U2587 (N_2587,N_2196,N_2302);
nor U2588 (N_2588,N_2181,N_1962);
nor U2589 (N_2589,N_2390,N_2111);
nor U2590 (N_2590,N_2123,N_2028);
xnor U2591 (N_2591,N_2247,N_2238);
nand U2592 (N_2592,N_1887,N_2059);
nand U2593 (N_2593,N_1852,N_2137);
nor U2594 (N_2594,N_2261,N_2225);
nor U2595 (N_2595,N_2251,N_1825);
and U2596 (N_2596,N_2087,N_2250);
xnor U2597 (N_2597,N_1860,N_2011);
or U2598 (N_2598,N_1877,N_2288);
nor U2599 (N_2599,N_1921,N_2066);
xnor U2600 (N_2600,N_1998,N_2086);
or U2601 (N_2601,N_2043,N_1959);
nand U2602 (N_2602,N_2396,N_1804);
and U2603 (N_2603,N_2076,N_2070);
xor U2604 (N_2604,N_2067,N_2290);
xnor U2605 (N_2605,N_1929,N_2392);
or U2606 (N_2606,N_2221,N_2283);
nand U2607 (N_2607,N_2176,N_1843);
or U2608 (N_2608,N_2009,N_1846);
or U2609 (N_2609,N_2255,N_1922);
xnor U2610 (N_2610,N_2088,N_2150);
nand U2611 (N_2611,N_1821,N_2294);
or U2612 (N_2612,N_2142,N_1863);
and U2613 (N_2613,N_1994,N_2265);
nand U2614 (N_2614,N_2327,N_1980);
or U2615 (N_2615,N_2257,N_2189);
nand U2616 (N_2616,N_1817,N_2064);
nor U2617 (N_2617,N_2234,N_2380);
xnor U2618 (N_2618,N_2367,N_1853);
nand U2619 (N_2619,N_2017,N_2212);
or U2620 (N_2620,N_2010,N_2200);
nor U2621 (N_2621,N_2223,N_1914);
or U2622 (N_2622,N_2268,N_2045);
or U2623 (N_2623,N_2077,N_2036);
nor U2624 (N_2624,N_2363,N_1868);
or U2625 (N_2625,N_2342,N_2032);
xor U2626 (N_2626,N_1872,N_2173);
and U2627 (N_2627,N_2239,N_1891);
and U2628 (N_2628,N_1885,N_1984);
nor U2629 (N_2629,N_1815,N_2355);
nor U2630 (N_2630,N_2034,N_2026);
or U2631 (N_2631,N_2198,N_1979);
or U2632 (N_2632,N_1803,N_2136);
and U2633 (N_2633,N_1943,N_1906);
xor U2634 (N_2634,N_2348,N_2071);
or U2635 (N_2635,N_1936,N_1826);
nor U2636 (N_2636,N_1896,N_2171);
xor U2637 (N_2637,N_2275,N_2106);
xnor U2638 (N_2638,N_1991,N_2095);
or U2639 (N_2639,N_2126,N_1881);
or U2640 (N_2640,N_2249,N_1871);
nor U2641 (N_2641,N_2385,N_1830);
or U2642 (N_2642,N_1974,N_2006);
and U2643 (N_2643,N_2287,N_2151);
or U2644 (N_2644,N_2023,N_1865);
nand U2645 (N_2645,N_2343,N_2129);
and U2646 (N_2646,N_2309,N_2031);
xor U2647 (N_2647,N_2264,N_2376);
or U2648 (N_2648,N_2269,N_2047);
and U2649 (N_2649,N_2167,N_1997);
xnor U2650 (N_2650,N_2022,N_2068);
and U2651 (N_2651,N_2175,N_2186);
nand U2652 (N_2652,N_2140,N_2296);
and U2653 (N_2653,N_2205,N_2313);
nor U2654 (N_2654,N_2187,N_2156);
nand U2655 (N_2655,N_2297,N_1813);
nor U2656 (N_2656,N_2192,N_1808);
and U2657 (N_2657,N_1833,N_2219);
nand U2658 (N_2658,N_2019,N_1838);
nand U2659 (N_2659,N_2197,N_2326);
and U2660 (N_2660,N_2202,N_2101);
or U2661 (N_2661,N_2191,N_2050);
or U2662 (N_2662,N_2001,N_1855);
xnor U2663 (N_2663,N_2201,N_2274);
nand U2664 (N_2664,N_2305,N_1956);
xor U2665 (N_2665,N_1989,N_1892);
nor U2666 (N_2666,N_2248,N_2332);
xnor U2667 (N_2667,N_2256,N_1934);
nor U2668 (N_2668,N_2236,N_2120);
and U2669 (N_2669,N_1878,N_1839);
xor U2670 (N_2670,N_1985,N_2046);
or U2671 (N_2671,N_2115,N_2285);
and U2672 (N_2672,N_2109,N_2334);
nand U2673 (N_2673,N_1850,N_1982);
xor U2674 (N_2674,N_2133,N_2130);
nand U2675 (N_2675,N_2018,N_1848);
nor U2676 (N_2676,N_2307,N_2346);
and U2677 (N_2677,N_1900,N_1910);
xor U2678 (N_2678,N_2391,N_2078);
nand U2679 (N_2679,N_2003,N_2090);
nor U2680 (N_2680,N_2278,N_2152);
xor U2681 (N_2681,N_2099,N_1820);
and U2682 (N_2682,N_1835,N_2345);
nor U2683 (N_2683,N_1837,N_2368);
xnor U2684 (N_2684,N_2276,N_2233);
or U2685 (N_2685,N_1993,N_1945);
nor U2686 (N_2686,N_1975,N_2035);
nor U2687 (N_2687,N_2024,N_1916);
or U2688 (N_2688,N_2399,N_2052);
nor U2689 (N_2689,N_1924,N_2104);
and U2690 (N_2690,N_2074,N_2127);
nor U2691 (N_2691,N_2357,N_2273);
xor U2692 (N_2692,N_1841,N_2138);
nor U2693 (N_2693,N_2012,N_2058);
nand U2694 (N_2694,N_2148,N_2282);
and U2695 (N_2695,N_2351,N_1911);
xor U2696 (N_2696,N_2147,N_2118);
nand U2697 (N_2697,N_1948,N_2103);
xnor U2698 (N_2698,N_2397,N_2075);
and U2699 (N_2699,N_1988,N_2260);
nand U2700 (N_2700,N_2016,N_1884);
and U2701 (N_2701,N_1988,N_1832);
xnor U2702 (N_2702,N_1985,N_1949);
nor U2703 (N_2703,N_1851,N_2301);
and U2704 (N_2704,N_1926,N_2361);
and U2705 (N_2705,N_1966,N_2084);
nor U2706 (N_2706,N_2193,N_2281);
nand U2707 (N_2707,N_2150,N_2064);
nor U2708 (N_2708,N_1975,N_2330);
and U2709 (N_2709,N_1827,N_2165);
xnor U2710 (N_2710,N_2033,N_2348);
nand U2711 (N_2711,N_2292,N_2340);
xnor U2712 (N_2712,N_1918,N_2307);
or U2713 (N_2713,N_1822,N_2218);
nor U2714 (N_2714,N_1802,N_2179);
nor U2715 (N_2715,N_2268,N_1858);
nor U2716 (N_2716,N_2107,N_2102);
nand U2717 (N_2717,N_2136,N_2025);
xor U2718 (N_2718,N_2345,N_2201);
or U2719 (N_2719,N_2309,N_2375);
or U2720 (N_2720,N_2113,N_2108);
nor U2721 (N_2721,N_2310,N_1909);
and U2722 (N_2722,N_1912,N_2396);
nor U2723 (N_2723,N_2260,N_1807);
or U2724 (N_2724,N_2118,N_1980);
nand U2725 (N_2725,N_1970,N_2280);
xnor U2726 (N_2726,N_2133,N_1992);
and U2727 (N_2727,N_2261,N_1896);
nor U2728 (N_2728,N_1934,N_2308);
or U2729 (N_2729,N_2325,N_2223);
nor U2730 (N_2730,N_2116,N_2033);
nand U2731 (N_2731,N_2397,N_2172);
nor U2732 (N_2732,N_2047,N_1883);
or U2733 (N_2733,N_2162,N_1850);
nor U2734 (N_2734,N_2131,N_2286);
nor U2735 (N_2735,N_1857,N_1932);
and U2736 (N_2736,N_2297,N_1992);
xnor U2737 (N_2737,N_2251,N_1877);
nand U2738 (N_2738,N_1896,N_2268);
nand U2739 (N_2739,N_2311,N_1853);
xnor U2740 (N_2740,N_1881,N_2305);
and U2741 (N_2741,N_1977,N_2195);
xnor U2742 (N_2742,N_2039,N_2395);
xnor U2743 (N_2743,N_2299,N_1944);
nor U2744 (N_2744,N_2220,N_2085);
and U2745 (N_2745,N_1932,N_2199);
or U2746 (N_2746,N_2284,N_2298);
xor U2747 (N_2747,N_2330,N_2026);
and U2748 (N_2748,N_2294,N_2161);
nand U2749 (N_2749,N_2318,N_2256);
or U2750 (N_2750,N_1837,N_2049);
nor U2751 (N_2751,N_1940,N_1935);
nand U2752 (N_2752,N_2323,N_1811);
xor U2753 (N_2753,N_2153,N_1856);
and U2754 (N_2754,N_2351,N_1902);
or U2755 (N_2755,N_2340,N_2122);
nand U2756 (N_2756,N_2251,N_2043);
or U2757 (N_2757,N_2062,N_2211);
nand U2758 (N_2758,N_2139,N_1826);
nor U2759 (N_2759,N_1930,N_2095);
xor U2760 (N_2760,N_1964,N_1974);
nor U2761 (N_2761,N_2270,N_1993);
xnor U2762 (N_2762,N_1950,N_2091);
or U2763 (N_2763,N_2304,N_2137);
nand U2764 (N_2764,N_1971,N_2364);
and U2765 (N_2765,N_2027,N_2216);
xnor U2766 (N_2766,N_2082,N_2282);
xor U2767 (N_2767,N_2211,N_2006);
nand U2768 (N_2768,N_2109,N_2370);
nand U2769 (N_2769,N_1909,N_1983);
or U2770 (N_2770,N_2048,N_2219);
and U2771 (N_2771,N_2262,N_2152);
nand U2772 (N_2772,N_2107,N_2158);
nor U2773 (N_2773,N_2327,N_2165);
or U2774 (N_2774,N_1864,N_2013);
or U2775 (N_2775,N_1838,N_2117);
xor U2776 (N_2776,N_2260,N_2120);
nor U2777 (N_2777,N_2250,N_2197);
xor U2778 (N_2778,N_2114,N_2000);
and U2779 (N_2779,N_1830,N_1911);
nand U2780 (N_2780,N_2162,N_2212);
and U2781 (N_2781,N_2007,N_1829);
nand U2782 (N_2782,N_2247,N_2054);
nand U2783 (N_2783,N_2208,N_2065);
xor U2784 (N_2784,N_1924,N_2197);
xor U2785 (N_2785,N_1835,N_2232);
nor U2786 (N_2786,N_2321,N_2088);
nand U2787 (N_2787,N_2174,N_1935);
or U2788 (N_2788,N_2328,N_1914);
nand U2789 (N_2789,N_1884,N_1865);
nor U2790 (N_2790,N_2057,N_2126);
nor U2791 (N_2791,N_2002,N_2073);
xnor U2792 (N_2792,N_2066,N_1963);
nand U2793 (N_2793,N_2131,N_1880);
xnor U2794 (N_2794,N_1860,N_2186);
nand U2795 (N_2795,N_2374,N_2337);
and U2796 (N_2796,N_2285,N_2099);
and U2797 (N_2797,N_2128,N_2113);
or U2798 (N_2798,N_2273,N_1826);
or U2799 (N_2799,N_2265,N_2166);
xor U2800 (N_2800,N_2093,N_2069);
nor U2801 (N_2801,N_2053,N_2067);
xor U2802 (N_2802,N_1869,N_1952);
nor U2803 (N_2803,N_2244,N_2387);
nand U2804 (N_2804,N_2213,N_1871);
or U2805 (N_2805,N_2068,N_2258);
xor U2806 (N_2806,N_2328,N_2224);
and U2807 (N_2807,N_1867,N_2304);
or U2808 (N_2808,N_1880,N_2353);
nor U2809 (N_2809,N_2145,N_2156);
xnor U2810 (N_2810,N_2054,N_2377);
and U2811 (N_2811,N_2074,N_1918);
nor U2812 (N_2812,N_2043,N_2052);
nand U2813 (N_2813,N_1922,N_2310);
xor U2814 (N_2814,N_2112,N_2261);
nand U2815 (N_2815,N_2044,N_1804);
nand U2816 (N_2816,N_2058,N_1977);
xor U2817 (N_2817,N_1810,N_2168);
xor U2818 (N_2818,N_2082,N_2371);
or U2819 (N_2819,N_2021,N_2140);
and U2820 (N_2820,N_2201,N_2351);
or U2821 (N_2821,N_2060,N_2252);
or U2822 (N_2822,N_1840,N_2264);
nor U2823 (N_2823,N_1872,N_2349);
nand U2824 (N_2824,N_2189,N_2224);
xnor U2825 (N_2825,N_2004,N_1992);
and U2826 (N_2826,N_2380,N_2194);
nor U2827 (N_2827,N_2034,N_1829);
and U2828 (N_2828,N_2095,N_2215);
or U2829 (N_2829,N_2345,N_2136);
xnor U2830 (N_2830,N_1931,N_2129);
or U2831 (N_2831,N_2170,N_2004);
nor U2832 (N_2832,N_2055,N_2357);
xnor U2833 (N_2833,N_2201,N_2299);
nor U2834 (N_2834,N_2293,N_2147);
nand U2835 (N_2835,N_1996,N_1802);
nor U2836 (N_2836,N_1858,N_2229);
nor U2837 (N_2837,N_1886,N_1977);
and U2838 (N_2838,N_2266,N_2234);
nand U2839 (N_2839,N_2335,N_2030);
nand U2840 (N_2840,N_1892,N_2000);
and U2841 (N_2841,N_1806,N_1997);
nor U2842 (N_2842,N_2011,N_1859);
xor U2843 (N_2843,N_2043,N_2374);
and U2844 (N_2844,N_1961,N_2064);
xnor U2845 (N_2845,N_1955,N_1993);
nor U2846 (N_2846,N_1896,N_2301);
and U2847 (N_2847,N_2210,N_2100);
nand U2848 (N_2848,N_2149,N_2089);
xnor U2849 (N_2849,N_2337,N_2108);
xnor U2850 (N_2850,N_1933,N_2069);
xnor U2851 (N_2851,N_2138,N_1847);
xnor U2852 (N_2852,N_2329,N_1882);
nor U2853 (N_2853,N_2232,N_1999);
nor U2854 (N_2854,N_2227,N_2136);
nor U2855 (N_2855,N_1838,N_2376);
nand U2856 (N_2856,N_1889,N_1882);
xor U2857 (N_2857,N_2101,N_1889);
and U2858 (N_2858,N_1854,N_2208);
and U2859 (N_2859,N_1944,N_1967);
nand U2860 (N_2860,N_2361,N_2181);
and U2861 (N_2861,N_1914,N_1944);
and U2862 (N_2862,N_2255,N_1884);
nor U2863 (N_2863,N_2138,N_2080);
nor U2864 (N_2864,N_2157,N_2264);
or U2865 (N_2865,N_2363,N_2090);
or U2866 (N_2866,N_2279,N_2008);
and U2867 (N_2867,N_2330,N_2379);
nand U2868 (N_2868,N_2173,N_1964);
and U2869 (N_2869,N_2309,N_2242);
or U2870 (N_2870,N_2372,N_2117);
and U2871 (N_2871,N_2225,N_2354);
or U2872 (N_2872,N_1853,N_2219);
and U2873 (N_2873,N_2267,N_2125);
and U2874 (N_2874,N_2026,N_1941);
and U2875 (N_2875,N_2355,N_2173);
nor U2876 (N_2876,N_2117,N_1827);
and U2877 (N_2877,N_1873,N_1968);
nor U2878 (N_2878,N_1846,N_2387);
nor U2879 (N_2879,N_2183,N_2091);
or U2880 (N_2880,N_1960,N_1986);
nand U2881 (N_2881,N_1833,N_2142);
nand U2882 (N_2882,N_1925,N_2038);
and U2883 (N_2883,N_2032,N_2013);
xnor U2884 (N_2884,N_2113,N_2393);
nand U2885 (N_2885,N_1829,N_2390);
xnor U2886 (N_2886,N_2031,N_2335);
nor U2887 (N_2887,N_2028,N_1887);
and U2888 (N_2888,N_2364,N_1937);
and U2889 (N_2889,N_2213,N_2299);
and U2890 (N_2890,N_1997,N_1975);
and U2891 (N_2891,N_1806,N_2330);
xor U2892 (N_2892,N_2058,N_2253);
or U2893 (N_2893,N_2233,N_2116);
xnor U2894 (N_2894,N_1921,N_2161);
nand U2895 (N_2895,N_2357,N_1879);
nand U2896 (N_2896,N_2003,N_1852);
or U2897 (N_2897,N_1913,N_2024);
xor U2898 (N_2898,N_2280,N_1948);
xnor U2899 (N_2899,N_2095,N_1860);
and U2900 (N_2900,N_1934,N_1999);
or U2901 (N_2901,N_1889,N_1814);
or U2902 (N_2902,N_1919,N_1908);
or U2903 (N_2903,N_2083,N_2377);
nand U2904 (N_2904,N_2291,N_1978);
and U2905 (N_2905,N_2222,N_1950);
nor U2906 (N_2906,N_2169,N_1964);
xor U2907 (N_2907,N_2369,N_2077);
nand U2908 (N_2908,N_2165,N_2283);
nor U2909 (N_2909,N_2129,N_2186);
nand U2910 (N_2910,N_2141,N_2349);
or U2911 (N_2911,N_1838,N_2311);
xor U2912 (N_2912,N_2214,N_2129);
nand U2913 (N_2913,N_2356,N_2232);
or U2914 (N_2914,N_1993,N_2028);
nor U2915 (N_2915,N_2158,N_2175);
nor U2916 (N_2916,N_2060,N_2336);
xor U2917 (N_2917,N_2146,N_1998);
nor U2918 (N_2918,N_2392,N_1844);
nor U2919 (N_2919,N_2293,N_1853);
and U2920 (N_2920,N_1834,N_1961);
nand U2921 (N_2921,N_2296,N_2370);
xnor U2922 (N_2922,N_2148,N_2178);
nand U2923 (N_2923,N_2353,N_2285);
or U2924 (N_2924,N_1845,N_1997);
nand U2925 (N_2925,N_2294,N_2304);
xnor U2926 (N_2926,N_1822,N_2094);
or U2927 (N_2927,N_2275,N_2064);
xnor U2928 (N_2928,N_2016,N_2148);
xnor U2929 (N_2929,N_2181,N_2309);
xor U2930 (N_2930,N_1808,N_2256);
and U2931 (N_2931,N_2113,N_2065);
and U2932 (N_2932,N_2373,N_2278);
and U2933 (N_2933,N_1960,N_2263);
or U2934 (N_2934,N_2273,N_2274);
xor U2935 (N_2935,N_2049,N_1950);
xnor U2936 (N_2936,N_1955,N_2280);
or U2937 (N_2937,N_2103,N_2247);
xnor U2938 (N_2938,N_1823,N_2119);
and U2939 (N_2939,N_2237,N_2390);
and U2940 (N_2940,N_2301,N_2051);
or U2941 (N_2941,N_1914,N_1880);
xnor U2942 (N_2942,N_2355,N_1820);
nor U2943 (N_2943,N_1835,N_2222);
and U2944 (N_2944,N_2341,N_2033);
and U2945 (N_2945,N_2172,N_2393);
or U2946 (N_2946,N_1962,N_2169);
xnor U2947 (N_2947,N_2346,N_1981);
or U2948 (N_2948,N_1949,N_2019);
xor U2949 (N_2949,N_2040,N_1998);
and U2950 (N_2950,N_1846,N_2105);
or U2951 (N_2951,N_2221,N_2280);
nor U2952 (N_2952,N_2235,N_2033);
nand U2953 (N_2953,N_2242,N_1831);
and U2954 (N_2954,N_2055,N_2232);
nor U2955 (N_2955,N_2371,N_2029);
nand U2956 (N_2956,N_2304,N_1942);
and U2957 (N_2957,N_1942,N_2227);
and U2958 (N_2958,N_1884,N_1969);
xor U2959 (N_2959,N_2304,N_1891);
nor U2960 (N_2960,N_2035,N_1932);
xor U2961 (N_2961,N_2274,N_2045);
nand U2962 (N_2962,N_2251,N_2342);
or U2963 (N_2963,N_1808,N_2341);
or U2964 (N_2964,N_2137,N_2168);
nand U2965 (N_2965,N_2339,N_1910);
nor U2966 (N_2966,N_1949,N_2224);
and U2967 (N_2967,N_2354,N_2104);
or U2968 (N_2968,N_2156,N_1907);
nand U2969 (N_2969,N_1878,N_2059);
nand U2970 (N_2970,N_1946,N_2001);
xnor U2971 (N_2971,N_1910,N_2331);
xnor U2972 (N_2972,N_2032,N_2228);
nand U2973 (N_2973,N_2336,N_1912);
nor U2974 (N_2974,N_2044,N_2390);
xor U2975 (N_2975,N_2193,N_1921);
xor U2976 (N_2976,N_1837,N_2037);
xor U2977 (N_2977,N_2147,N_2050);
xor U2978 (N_2978,N_1920,N_2309);
xnor U2979 (N_2979,N_2244,N_1906);
xnor U2980 (N_2980,N_1888,N_1950);
xnor U2981 (N_2981,N_2358,N_2395);
nand U2982 (N_2982,N_1982,N_2183);
nor U2983 (N_2983,N_1840,N_2124);
and U2984 (N_2984,N_2105,N_2371);
and U2985 (N_2985,N_2327,N_2292);
and U2986 (N_2986,N_2217,N_1931);
or U2987 (N_2987,N_2196,N_2089);
nor U2988 (N_2988,N_2187,N_2123);
xor U2989 (N_2989,N_1827,N_2309);
nand U2990 (N_2990,N_1801,N_1896);
nand U2991 (N_2991,N_2359,N_1943);
nor U2992 (N_2992,N_1871,N_2339);
nand U2993 (N_2993,N_2255,N_2126);
nor U2994 (N_2994,N_2177,N_1920);
and U2995 (N_2995,N_2240,N_1935);
nor U2996 (N_2996,N_2144,N_2156);
or U2997 (N_2997,N_2318,N_1806);
nor U2998 (N_2998,N_1994,N_2105);
nand U2999 (N_2999,N_1948,N_1919);
and U3000 (N_3000,N_2653,N_2517);
nand U3001 (N_3001,N_2847,N_2532);
or U3002 (N_3002,N_2470,N_2900);
and U3003 (N_3003,N_2560,N_2666);
xor U3004 (N_3004,N_2541,N_2652);
or U3005 (N_3005,N_2467,N_2672);
nor U3006 (N_3006,N_2529,N_2704);
nor U3007 (N_3007,N_2970,N_2542);
nand U3008 (N_3008,N_2926,N_2886);
or U3009 (N_3009,N_2911,N_2875);
or U3010 (N_3010,N_2526,N_2505);
and U3011 (N_3011,N_2414,N_2726);
nor U3012 (N_3012,N_2942,N_2769);
nand U3013 (N_3013,N_2421,N_2494);
and U3014 (N_3014,N_2638,N_2691);
nor U3015 (N_3015,N_2885,N_2924);
nand U3016 (N_3016,N_2496,N_2798);
or U3017 (N_3017,N_2448,N_2751);
and U3018 (N_3018,N_2462,N_2565);
nor U3019 (N_3019,N_2760,N_2641);
and U3020 (N_3020,N_2405,N_2774);
or U3021 (N_3021,N_2734,N_2409);
or U3022 (N_3022,N_2819,N_2733);
and U3023 (N_3023,N_2568,N_2827);
or U3024 (N_3024,N_2739,N_2537);
nand U3025 (N_3025,N_2658,N_2834);
xor U3026 (N_3026,N_2512,N_2592);
xnor U3027 (N_3027,N_2964,N_2628);
or U3028 (N_3028,N_2502,N_2497);
and U3029 (N_3029,N_2780,N_2707);
nand U3030 (N_3030,N_2689,N_2775);
and U3031 (N_3031,N_2941,N_2822);
xor U3032 (N_3032,N_2711,N_2404);
xor U3033 (N_3033,N_2966,N_2511);
xor U3034 (N_3034,N_2755,N_2665);
nor U3035 (N_3035,N_2837,N_2443);
nand U3036 (N_3036,N_2651,N_2572);
or U3037 (N_3037,N_2730,N_2823);
xor U3038 (N_3038,N_2573,N_2852);
nor U3039 (N_3039,N_2934,N_2598);
nor U3040 (N_3040,N_2850,N_2981);
xor U3041 (N_3041,N_2872,N_2668);
and U3042 (N_3042,N_2682,N_2998);
or U3043 (N_3043,N_2862,N_2810);
and U3044 (N_3044,N_2548,N_2701);
or U3045 (N_3045,N_2622,N_2463);
xor U3046 (N_3046,N_2519,N_2438);
xor U3047 (N_3047,N_2887,N_2508);
nor U3048 (N_3048,N_2932,N_2670);
nor U3049 (N_3049,N_2960,N_2783);
nor U3050 (N_3050,N_2562,N_2506);
or U3051 (N_3051,N_2680,N_2871);
or U3052 (N_3052,N_2864,N_2476);
nor U3053 (N_3053,N_2640,N_2851);
nand U3054 (N_3054,N_2855,N_2967);
nand U3055 (N_3055,N_2993,N_2940);
or U3056 (N_3056,N_2831,N_2644);
nor U3057 (N_3057,N_2841,N_2796);
xnor U3058 (N_3058,N_2646,N_2988);
xor U3059 (N_3059,N_2430,N_2453);
or U3060 (N_3060,N_2824,N_2481);
nand U3061 (N_3061,N_2913,N_2809);
nand U3062 (N_3062,N_2659,N_2759);
or U3063 (N_3063,N_2999,N_2907);
nor U3064 (N_3064,N_2893,N_2863);
nand U3065 (N_3065,N_2884,N_2579);
xor U3066 (N_3066,N_2575,N_2498);
nand U3067 (N_3067,N_2718,N_2627);
nand U3068 (N_3068,N_2571,N_2762);
and U3069 (N_3069,N_2844,N_2996);
xor U3070 (N_3070,N_2814,N_2800);
nand U3071 (N_3071,N_2958,N_2539);
and U3072 (N_3072,N_2793,N_2766);
nand U3073 (N_3073,N_2499,N_2738);
xor U3074 (N_3074,N_2770,N_2699);
or U3075 (N_3075,N_2521,N_2475);
and U3076 (N_3076,N_2696,N_2802);
nand U3077 (N_3077,N_2559,N_2528);
and U3078 (N_3078,N_2585,N_2564);
and U3079 (N_3079,N_2626,N_2853);
or U3080 (N_3080,N_2583,N_2683);
nand U3081 (N_3081,N_2771,N_2749);
xnor U3082 (N_3082,N_2801,N_2637);
nor U3083 (N_3083,N_2747,N_2619);
and U3084 (N_3084,N_2763,N_2931);
and U3085 (N_3085,N_2446,N_2576);
nor U3086 (N_3086,N_2980,N_2879);
nand U3087 (N_3087,N_2451,N_2845);
or U3088 (N_3088,N_2631,N_2472);
xnor U3089 (N_3089,N_2563,N_2434);
xor U3090 (N_3090,N_2957,N_2412);
or U3091 (N_3091,N_2577,N_2588);
xnor U3092 (N_3092,N_2946,N_2503);
nand U3093 (N_3093,N_2890,N_2977);
or U3094 (N_3094,N_2849,N_2950);
or U3095 (N_3095,N_2587,N_2752);
nand U3096 (N_3096,N_2488,N_2584);
nor U3097 (N_3097,N_2660,N_2433);
or U3098 (N_3098,N_2961,N_2553);
xor U3099 (N_3099,N_2790,N_2440);
nor U3100 (N_3100,N_2925,N_2617);
nand U3101 (N_3101,N_2838,N_2840);
xnor U3102 (N_3102,N_2504,N_2877);
xor U3103 (N_3103,N_2558,N_2469);
xnor U3104 (N_3104,N_2507,N_2540);
xor U3105 (N_3105,N_2929,N_2791);
or U3106 (N_3106,N_2768,N_2570);
or U3107 (N_3107,N_2663,N_2818);
nor U3108 (N_3108,N_2500,N_2524);
xor U3109 (N_3109,N_2935,N_2543);
or U3110 (N_3110,N_2685,N_2690);
xor U3111 (N_3111,N_2968,N_2686);
xnor U3112 (N_3112,N_2899,N_2654);
xor U3113 (N_3113,N_2447,N_2535);
or U3114 (N_3114,N_2664,N_2482);
or U3115 (N_3115,N_2590,N_2677);
or U3116 (N_3116,N_2867,N_2994);
nor U3117 (N_3117,N_2544,N_2675);
nor U3118 (N_3118,N_2779,N_2902);
nor U3119 (N_3119,N_2483,N_2567);
xor U3120 (N_3120,N_2797,N_2905);
nand U3121 (N_3121,N_2546,N_2510);
nand U3122 (N_3122,N_2746,N_2489);
and U3123 (N_3123,N_2908,N_2557);
xnor U3124 (N_3124,N_2611,N_2735);
or U3125 (N_3125,N_2410,N_2625);
nor U3126 (N_3126,N_2679,N_2761);
and U3127 (N_3127,N_2623,N_2894);
and U3128 (N_3128,N_2439,N_2432);
or U3129 (N_3129,N_2477,N_2426);
or U3130 (N_3130,N_2669,N_2785);
nor U3131 (N_3131,N_2811,N_2678);
or U3132 (N_3132,N_2878,N_2431);
nor U3133 (N_3133,N_2953,N_2804);
xnor U3134 (N_3134,N_2859,N_2748);
nor U3135 (N_3135,N_2826,N_2985);
xor U3136 (N_3136,N_2815,N_2468);
nor U3137 (N_3137,N_2842,N_2717);
nand U3138 (N_3138,N_2525,N_2832);
nand U3139 (N_3139,N_2792,N_2866);
xor U3140 (N_3140,N_2634,N_2416);
xnor U3141 (N_3141,N_2778,N_2982);
and U3142 (N_3142,N_2989,N_2501);
or U3143 (N_3143,N_2916,N_2984);
nand U3144 (N_3144,N_2662,N_2991);
or U3145 (N_3145,N_2473,N_2649);
or U3146 (N_3146,N_2424,N_2784);
and U3147 (N_3147,N_2895,N_2605);
nand U3148 (N_3148,N_2955,N_2400);
xnor U3149 (N_3149,N_2962,N_2808);
and U3150 (N_3150,N_2522,N_2693);
nand U3151 (N_3151,N_2930,N_2445);
nand U3152 (N_3152,N_2765,N_2645);
nand U3153 (N_3153,N_2464,N_2956);
or U3154 (N_3154,N_2868,N_2594);
nor U3155 (N_3155,N_2614,N_2731);
nand U3156 (N_3156,N_2408,N_2455);
nor U3157 (N_3157,N_2648,N_2624);
and U3158 (N_3158,N_2580,N_2732);
nor U3159 (N_3159,N_2604,N_2436);
nand U3160 (N_3160,N_2465,N_2610);
or U3161 (N_3161,N_2657,N_2466);
nand U3162 (N_3162,N_2882,N_2402);
nor U3163 (N_3163,N_2856,N_2552);
and U3164 (N_3164,N_2520,N_2596);
nand U3165 (N_3165,N_2478,N_2773);
xnor U3166 (N_3166,N_2609,N_2835);
or U3167 (N_3167,N_2607,N_2971);
and U3168 (N_3168,N_2694,N_2873);
or U3169 (N_3169,N_2937,N_2741);
and U3170 (N_3170,N_2423,N_2406);
nor U3171 (N_3171,N_2758,N_2710);
nor U3172 (N_3172,N_2549,N_2582);
nor U3173 (N_3173,N_2700,N_2724);
or U3174 (N_3174,N_2684,N_2817);
and U3175 (N_3175,N_2547,N_2865);
xnor U3176 (N_3176,N_2742,N_2716);
or U3177 (N_3177,N_2939,N_2715);
and U3178 (N_3178,N_2427,N_2720);
and U3179 (N_3179,N_2471,N_2639);
nor U3180 (N_3180,N_2597,N_2903);
xor U3181 (N_3181,N_2554,N_2487);
or U3182 (N_3182,N_2754,N_2947);
nand U3183 (N_3183,N_2881,N_2990);
xnor U3184 (N_3184,N_2566,N_2921);
nor U3185 (N_3185,N_2417,N_2750);
nor U3186 (N_3186,N_2603,N_2945);
xor U3187 (N_3187,N_2538,N_2721);
nor U3188 (N_3188,N_2556,N_2972);
or U3189 (N_3189,N_2987,N_2983);
nand U3190 (N_3190,N_2671,N_2459);
nand U3191 (N_3191,N_2629,N_2632);
xnor U3192 (N_3192,N_2836,N_2601);
xnor U3193 (N_3193,N_2788,N_2687);
nor U3194 (N_3194,N_2725,N_2712);
nor U3195 (N_3195,N_2674,N_2608);
nand U3196 (N_3196,N_2723,N_2805);
and U3197 (N_3197,N_2457,N_2647);
and U3198 (N_3198,N_2456,N_2949);
xnor U3199 (N_3199,N_2753,N_2697);
nand U3200 (N_3200,N_2764,N_2550);
or U3201 (N_3201,N_2413,N_2479);
xor U3202 (N_3202,N_2437,N_2706);
and U3203 (N_3203,N_2860,N_2736);
nor U3204 (N_3204,N_2667,N_2782);
and U3205 (N_3205,N_2491,N_2643);
xnor U3206 (N_3206,N_2727,N_2534);
or U3207 (N_3207,N_2708,N_2460);
nor U3208 (N_3208,N_2767,N_2454);
or U3209 (N_3209,N_2812,N_2883);
xor U3210 (N_3210,N_2719,N_2613);
or U3211 (N_3211,N_2411,N_2442);
or U3212 (N_3212,N_2591,N_2915);
xor U3213 (N_3213,N_2909,N_2839);
xnor U3214 (N_3214,N_2642,N_2918);
nor U3215 (N_3215,N_2485,N_2518);
and U3216 (N_3216,N_2650,N_2786);
xnor U3217 (N_3217,N_2870,N_2936);
xor U3218 (N_3218,N_2880,N_2904);
nand U3219 (N_3219,N_2618,N_2745);
nor U3220 (N_3220,N_2515,N_2969);
nand U3221 (N_3221,N_2843,N_2449);
nor U3222 (N_3222,N_2531,N_2419);
or U3223 (N_3223,N_2495,N_2656);
and U3224 (N_3224,N_2729,N_2910);
or U3225 (N_3225,N_2551,N_2612);
and U3226 (N_3226,N_2403,N_2420);
or U3227 (N_3227,N_2787,N_2901);
nor U3228 (N_3228,N_2702,N_2829);
or U3229 (N_3229,N_2965,N_2995);
and U3230 (N_3230,N_2897,N_2533);
and U3231 (N_3231,N_2777,N_2536);
or U3232 (N_3232,N_2795,N_2976);
or U3233 (N_3233,N_2820,N_2615);
or U3234 (N_3234,N_2513,N_2794);
or U3235 (N_3235,N_2441,N_2586);
or U3236 (N_3236,N_2401,N_2630);
and U3237 (N_3237,N_2688,N_2616);
nand U3238 (N_3238,N_2407,N_2772);
and U3239 (N_3239,N_2633,N_2889);
or U3240 (N_3240,N_2673,N_2492);
or U3241 (N_3241,N_2914,N_2606);
nor U3242 (N_3242,N_2593,N_2555);
nor U3243 (N_3243,N_2861,N_2516);
nand U3244 (N_3244,N_2833,N_2858);
xnor U3245 (N_3245,N_2963,N_2561);
nand U3246 (N_3246,N_2922,N_2480);
or U3247 (N_3247,N_2923,N_2952);
nand U3248 (N_3248,N_2461,N_2635);
or U3249 (N_3249,N_2944,N_2444);
nand U3250 (N_3250,N_2415,N_2602);
nand U3251 (N_3251,N_2545,N_2425);
nand U3252 (N_3252,N_2891,N_2848);
nor U3253 (N_3253,N_2530,N_2744);
or U3254 (N_3254,N_2789,N_2943);
nand U3255 (N_3255,N_2509,N_2493);
nand U3256 (N_3256,N_2830,N_2484);
and U3257 (N_3257,N_2722,N_2661);
or U3258 (N_3258,N_2756,N_2986);
nand U3259 (N_3259,N_2927,N_2523);
nor U3260 (N_3260,N_2874,N_2813);
xnor U3261 (N_3261,N_2450,N_2973);
xor U3262 (N_3262,N_2428,N_2692);
nor U3263 (N_3263,N_2620,N_2954);
and U3264 (N_3264,N_2806,N_2574);
nor U3265 (N_3265,N_2709,N_2698);
and U3266 (N_3266,N_2974,N_2828);
xnor U3267 (N_3267,N_2992,N_2490);
and U3268 (N_3268,N_2912,N_2599);
xor U3269 (N_3269,N_2920,N_2418);
xnor U3270 (N_3270,N_2919,N_2892);
nand U3271 (N_3271,N_2527,N_2825);
nand U3272 (N_3272,N_2979,N_2600);
nand U3273 (N_3273,N_2799,N_2743);
nor U3274 (N_3274,N_2846,N_2803);
and U3275 (N_3275,N_2997,N_2776);
xor U3276 (N_3276,N_2898,N_2636);
nand U3277 (N_3277,N_2728,N_2933);
or U3278 (N_3278,N_2695,N_2581);
nor U3279 (N_3279,N_2435,N_2681);
and U3280 (N_3280,N_2959,N_2703);
nand U3281 (N_3281,N_2757,N_2906);
xor U3282 (N_3282,N_2713,N_2705);
or U3283 (N_3283,N_2737,N_2429);
nor U3284 (N_3284,N_2821,N_2569);
nand U3285 (N_3285,N_2486,N_2595);
or U3286 (N_3286,N_2807,N_2951);
nor U3287 (N_3287,N_2676,N_2816);
and U3288 (N_3288,N_2928,N_2458);
xor U3289 (N_3289,N_2857,N_2896);
and U3290 (N_3290,N_2948,N_2781);
xnor U3291 (N_3291,N_2655,N_2854);
and U3292 (N_3292,N_2888,N_2578);
nor U3293 (N_3293,N_2740,N_2876);
nor U3294 (N_3294,N_2452,N_2422);
nand U3295 (N_3295,N_2978,N_2869);
or U3296 (N_3296,N_2514,N_2714);
or U3297 (N_3297,N_2589,N_2917);
xor U3298 (N_3298,N_2975,N_2938);
or U3299 (N_3299,N_2474,N_2621);
nand U3300 (N_3300,N_2602,N_2976);
nand U3301 (N_3301,N_2959,N_2605);
xnor U3302 (N_3302,N_2422,N_2638);
nand U3303 (N_3303,N_2943,N_2509);
nor U3304 (N_3304,N_2806,N_2721);
nor U3305 (N_3305,N_2857,N_2642);
or U3306 (N_3306,N_2642,N_2592);
nand U3307 (N_3307,N_2847,N_2472);
nor U3308 (N_3308,N_2625,N_2597);
xnor U3309 (N_3309,N_2444,N_2578);
or U3310 (N_3310,N_2693,N_2910);
nand U3311 (N_3311,N_2940,N_2724);
nor U3312 (N_3312,N_2457,N_2461);
nand U3313 (N_3313,N_2499,N_2904);
or U3314 (N_3314,N_2699,N_2454);
nor U3315 (N_3315,N_2512,N_2483);
xnor U3316 (N_3316,N_2791,N_2910);
nor U3317 (N_3317,N_2456,N_2652);
nand U3318 (N_3318,N_2489,N_2881);
nor U3319 (N_3319,N_2765,N_2518);
and U3320 (N_3320,N_2450,N_2802);
or U3321 (N_3321,N_2948,N_2910);
nor U3322 (N_3322,N_2688,N_2629);
or U3323 (N_3323,N_2822,N_2927);
nand U3324 (N_3324,N_2833,N_2768);
nand U3325 (N_3325,N_2442,N_2515);
nand U3326 (N_3326,N_2873,N_2747);
nor U3327 (N_3327,N_2936,N_2959);
xnor U3328 (N_3328,N_2503,N_2524);
nand U3329 (N_3329,N_2643,N_2530);
xor U3330 (N_3330,N_2761,N_2480);
and U3331 (N_3331,N_2428,N_2541);
and U3332 (N_3332,N_2650,N_2558);
and U3333 (N_3333,N_2690,N_2867);
nor U3334 (N_3334,N_2862,N_2775);
and U3335 (N_3335,N_2699,N_2999);
and U3336 (N_3336,N_2652,N_2481);
nor U3337 (N_3337,N_2818,N_2584);
or U3338 (N_3338,N_2885,N_2721);
nor U3339 (N_3339,N_2998,N_2609);
nor U3340 (N_3340,N_2838,N_2763);
and U3341 (N_3341,N_2634,N_2922);
and U3342 (N_3342,N_2821,N_2923);
or U3343 (N_3343,N_2606,N_2650);
and U3344 (N_3344,N_2697,N_2436);
nor U3345 (N_3345,N_2618,N_2641);
and U3346 (N_3346,N_2415,N_2657);
or U3347 (N_3347,N_2822,N_2414);
nand U3348 (N_3348,N_2612,N_2615);
and U3349 (N_3349,N_2661,N_2846);
and U3350 (N_3350,N_2794,N_2419);
or U3351 (N_3351,N_2794,N_2535);
xor U3352 (N_3352,N_2423,N_2926);
or U3353 (N_3353,N_2546,N_2999);
nand U3354 (N_3354,N_2902,N_2918);
or U3355 (N_3355,N_2420,N_2433);
and U3356 (N_3356,N_2704,N_2642);
nor U3357 (N_3357,N_2604,N_2939);
and U3358 (N_3358,N_2847,N_2435);
xnor U3359 (N_3359,N_2642,N_2561);
xnor U3360 (N_3360,N_2985,N_2572);
and U3361 (N_3361,N_2858,N_2991);
nor U3362 (N_3362,N_2906,N_2832);
or U3363 (N_3363,N_2751,N_2497);
or U3364 (N_3364,N_2676,N_2638);
nand U3365 (N_3365,N_2977,N_2589);
and U3366 (N_3366,N_2470,N_2694);
or U3367 (N_3367,N_2644,N_2635);
nor U3368 (N_3368,N_2586,N_2778);
or U3369 (N_3369,N_2953,N_2590);
or U3370 (N_3370,N_2598,N_2591);
and U3371 (N_3371,N_2933,N_2542);
xnor U3372 (N_3372,N_2424,N_2780);
nor U3373 (N_3373,N_2592,N_2457);
xor U3374 (N_3374,N_2863,N_2809);
xnor U3375 (N_3375,N_2452,N_2911);
nor U3376 (N_3376,N_2629,N_2652);
or U3377 (N_3377,N_2857,N_2736);
and U3378 (N_3378,N_2989,N_2613);
nor U3379 (N_3379,N_2959,N_2911);
or U3380 (N_3380,N_2587,N_2971);
or U3381 (N_3381,N_2635,N_2826);
and U3382 (N_3382,N_2484,N_2654);
or U3383 (N_3383,N_2783,N_2464);
xnor U3384 (N_3384,N_2494,N_2449);
xnor U3385 (N_3385,N_2653,N_2891);
xnor U3386 (N_3386,N_2441,N_2699);
nand U3387 (N_3387,N_2898,N_2515);
nor U3388 (N_3388,N_2682,N_2438);
nand U3389 (N_3389,N_2925,N_2847);
or U3390 (N_3390,N_2628,N_2703);
or U3391 (N_3391,N_2962,N_2584);
nand U3392 (N_3392,N_2689,N_2489);
xor U3393 (N_3393,N_2975,N_2708);
and U3394 (N_3394,N_2445,N_2500);
and U3395 (N_3395,N_2498,N_2455);
or U3396 (N_3396,N_2578,N_2985);
and U3397 (N_3397,N_2729,N_2552);
xor U3398 (N_3398,N_2730,N_2523);
nand U3399 (N_3399,N_2892,N_2785);
nor U3400 (N_3400,N_2579,N_2507);
xor U3401 (N_3401,N_2854,N_2431);
xor U3402 (N_3402,N_2648,N_2799);
nand U3403 (N_3403,N_2929,N_2786);
or U3404 (N_3404,N_2540,N_2942);
or U3405 (N_3405,N_2935,N_2815);
nand U3406 (N_3406,N_2514,N_2978);
nand U3407 (N_3407,N_2970,N_2704);
nand U3408 (N_3408,N_2575,N_2557);
or U3409 (N_3409,N_2859,N_2404);
or U3410 (N_3410,N_2864,N_2993);
nand U3411 (N_3411,N_2836,N_2569);
and U3412 (N_3412,N_2479,N_2498);
or U3413 (N_3413,N_2913,N_2732);
nor U3414 (N_3414,N_2814,N_2607);
xor U3415 (N_3415,N_2420,N_2874);
xor U3416 (N_3416,N_2870,N_2498);
xor U3417 (N_3417,N_2597,N_2417);
nand U3418 (N_3418,N_2653,N_2970);
xor U3419 (N_3419,N_2770,N_2468);
or U3420 (N_3420,N_2803,N_2753);
nand U3421 (N_3421,N_2819,N_2511);
nand U3422 (N_3422,N_2578,N_2820);
or U3423 (N_3423,N_2682,N_2875);
nor U3424 (N_3424,N_2726,N_2418);
and U3425 (N_3425,N_2435,N_2461);
nand U3426 (N_3426,N_2582,N_2471);
xnor U3427 (N_3427,N_2689,N_2739);
and U3428 (N_3428,N_2690,N_2457);
xnor U3429 (N_3429,N_2415,N_2849);
and U3430 (N_3430,N_2504,N_2422);
and U3431 (N_3431,N_2940,N_2413);
nor U3432 (N_3432,N_2400,N_2587);
xnor U3433 (N_3433,N_2788,N_2882);
xor U3434 (N_3434,N_2923,N_2998);
nand U3435 (N_3435,N_2455,N_2502);
or U3436 (N_3436,N_2915,N_2653);
nor U3437 (N_3437,N_2597,N_2982);
nor U3438 (N_3438,N_2585,N_2419);
xnor U3439 (N_3439,N_2509,N_2565);
xnor U3440 (N_3440,N_2886,N_2709);
nor U3441 (N_3441,N_2584,N_2587);
nand U3442 (N_3442,N_2470,N_2569);
xnor U3443 (N_3443,N_2749,N_2711);
nand U3444 (N_3444,N_2778,N_2575);
nand U3445 (N_3445,N_2488,N_2756);
xnor U3446 (N_3446,N_2612,N_2889);
xnor U3447 (N_3447,N_2913,N_2878);
and U3448 (N_3448,N_2658,N_2955);
xnor U3449 (N_3449,N_2590,N_2469);
nand U3450 (N_3450,N_2506,N_2703);
and U3451 (N_3451,N_2984,N_2810);
and U3452 (N_3452,N_2654,N_2702);
or U3453 (N_3453,N_2544,N_2809);
or U3454 (N_3454,N_2541,N_2715);
nand U3455 (N_3455,N_2880,N_2579);
or U3456 (N_3456,N_2915,N_2713);
or U3457 (N_3457,N_2519,N_2469);
nor U3458 (N_3458,N_2859,N_2945);
xor U3459 (N_3459,N_2612,N_2706);
nand U3460 (N_3460,N_2860,N_2990);
nand U3461 (N_3461,N_2587,N_2541);
and U3462 (N_3462,N_2431,N_2791);
nand U3463 (N_3463,N_2421,N_2417);
nand U3464 (N_3464,N_2995,N_2968);
and U3465 (N_3465,N_2515,N_2847);
or U3466 (N_3466,N_2835,N_2717);
and U3467 (N_3467,N_2479,N_2408);
and U3468 (N_3468,N_2979,N_2464);
and U3469 (N_3469,N_2871,N_2627);
nor U3470 (N_3470,N_2504,N_2945);
and U3471 (N_3471,N_2465,N_2510);
xnor U3472 (N_3472,N_2941,N_2447);
and U3473 (N_3473,N_2429,N_2577);
and U3474 (N_3474,N_2796,N_2726);
nor U3475 (N_3475,N_2900,N_2926);
nor U3476 (N_3476,N_2891,N_2839);
and U3477 (N_3477,N_2909,N_2934);
nor U3478 (N_3478,N_2838,N_2424);
nor U3479 (N_3479,N_2653,N_2570);
or U3480 (N_3480,N_2798,N_2851);
or U3481 (N_3481,N_2900,N_2859);
xor U3482 (N_3482,N_2438,N_2540);
or U3483 (N_3483,N_2461,N_2904);
xnor U3484 (N_3484,N_2473,N_2489);
xor U3485 (N_3485,N_2404,N_2402);
nand U3486 (N_3486,N_2664,N_2827);
xor U3487 (N_3487,N_2568,N_2678);
nor U3488 (N_3488,N_2518,N_2593);
or U3489 (N_3489,N_2590,N_2436);
xor U3490 (N_3490,N_2663,N_2975);
nand U3491 (N_3491,N_2920,N_2545);
xnor U3492 (N_3492,N_2425,N_2424);
or U3493 (N_3493,N_2785,N_2849);
xnor U3494 (N_3494,N_2711,N_2585);
nor U3495 (N_3495,N_2738,N_2955);
nand U3496 (N_3496,N_2651,N_2458);
nor U3497 (N_3497,N_2863,N_2643);
or U3498 (N_3498,N_2829,N_2738);
nand U3499 (N_3499,N_2520,N_2531);
and U3500 (N_3500,N_2934,N_2569);
and U3501 (N_3501,N_2551,N_2415);
or U3502 (N_3502,N_2685,N_2930);
xnor U3503 (N_3503,N_2535,N_2924);
and U3504 (N_3504,N_2892,N_2505);
xor U3505 (N_3505,N_2493,N_2595);
nor U3506 (N_3506,N_2575,N_2701);
xor U3507 (N_3507,N_2471,N_2653);
nand U3508 (N_3508,N_2681,N_2465);
and U3509 (N_3509,N_2907,N_2493);
xnor U3510 (N_3510,N_2836,N_2503);
or U3511 (N_3511,N_2431,N_2955);
nand U3512 (N_3512,N_2458,N_2539);
and U3513 (N_3513,N_2908,N_2662);
nor U3514 (N_3514,N_2825,N_2470);
and U3515 (N_3515,N_2624,N_2592);
and U3516 (N_3516,N_2589,N_2960);
or U3517 (N_3517,N_2962,N_2433);
xor U3518 (N_3518,N_2613,N_2528);
and U3519 (N_3519,N_2637,N_2665);
and U3520 (N_3520,N_2694,N_2681);
nand U3521 (N_3521,N_2826,N_2690);
nor U3522 (N_3522,N_2824,N_2685);
nand U3523 (N_3523,N_2626,N_2942);
xor U3524 (N_3524,N_2596,N_2589);
nor U3525 (N_3525,N_2648,N_2584);
and U3526 (N_3526,N_2580,N_2647);
nor U3527 (N_3527,N_2555,N_2646);
nor U3528 (N_3528,N_2748,N_2554);
or U3529 (N_3529,N_2923,N_2613);
or U3530 (N_3530,N_2743,N_2705);
xor U3531 (N_3531,N_2636,N_2718);
and U3532 (N_3532,N_2588,N_2584);
nor U3533 (N_3533,N_2726,N_2758);
nand U3534 (N_3534,N_2579,N_2487);
xnor U3535 (N_3535,N_2814,N_2605);
nor U3536 (N_3536,N_2724,N_2410);
xnor U3537 (N_3537,N_2754,N_2849);
and U3538 (N_3538,N_2631,N_2766);
or U3539 (N_3539,N_2719,N_2938);
and U3540 (N_3540,N_2543,N_2835);
or U3541 (N_3541,N_2860,N_2666);
or U3542 (N_3542,N_2859,N_2403);
nand U3543 (N_3543,N_2784,N_2850);
xnor U3544 (N_3544,N_2646,N_2911);
nand U3545 (N_3545,N_2727,N_2968);
nand U3546 (N_3546,N_2732,N_2763);
or U3547 (N_3547,N_2627,N_2507);
nor U3548 (N_3548,N_2585,N_2940);
nand U3549 (N_3549,N_2528,N_2416);
and U3550 (N_3550,N_2670,N_2726);
nor U3551 (N_3551,N_2484,N_2829);
xor U3552 (N_3552,N_2547,N_2414);
xnor U3553 (N_3553,N_2672,N_2770);
nand U3554 (N_3554,N_2924,N_2969);
and U3555 (N_3555,N_2818,N_2940);
or U3556 (N_3556,N_2785,N_2584);
nor U3557 (N_3557,N_2774,N_2973);
nand U3558 (N_3558,N_2522,N_2469);
xor U3559 (N_3559,N_2497,N_2901);
or U3560 (N_3560,N_2491,N_2718);
or U3561 (N_3561,N_2866,N_2735);
and U3562 (N_3562,N_2471,N_2844);
xnor U3563 (N_3563,N_2737,N_2802);
and U3564 (N_3564,N_2966,N_2510);
nand U3565 (N_3565,N_2444,N_2930);
or U3566 (N_3566,N_2678,N_2947);
or U3567 (N_3567,N_2412,N_2529);
or U3568 (N_3568,N_2651,N_2889);
or U3569 (N_3569,N_2842,N_2494);
nor U3570 (N_3570,N_2799,N_2437);
or U3571 (N_3571,N_2906,N_2632);
nand U3572 (N_3572,N_2415,N_2887);
and U3573 (N_3573,N_2670,N_2415);
and U3574 (N_3574,N_2516,N_2487);
xnor U3575 (N_3575,N_2920,N_2516);
xor U3576 (N_3576,N_2603,N_2495);
nand U3577 (N_3577,N_2720,N_2925);
nor U3578 (N_3578,N_2863,N_2936);
nor U3579 (N_3579,N_2488,N_2990);
xnor U3580 (N_3580,N_2537,N_2892);
or U3581 (N_3581,N_2971,N_2784);
and U3582 (N_3582,N_2646,N_2562);
or U3583 (N_3583,N_2433,N_2481);
nand U3584 (N_3584,N_2985,N_2919);
or U3585 (N_3585,N_2800,N_2480);
nor U3586 (N_3586,N_2985,N_2628);
xor U3587 (N_3587,N_2965,N_2409);
and U3588 (N_3588,N_2813,N_2899);
nand U3589 (N_3589,N_2603,N_2565);
xor U3590 (N_3590,N_2864,N_2672);
nand U3591 (N_3591,N_2494,N_2502);
nand U3592 (N_3592,N_2694,N_2718);
and U3593 (N_3593,N_2720,N_2982);
xor U3594 (N_3594,N_2922,N_2521);
xnor U3595 (N_3595,N_2932,N_2665);
or U3596 (N_3596,N_2802,N_2663);
or U3597 (N_3597,N_2957,N_2704);
and U3598 (N_3598,N_2834,N_2503);
or U3599 (N_3599,N_2792,N_2688);
and U3600 (N_3600,N_3307,N_3253);
nand U3601 (N_3601,N_3022,N_3296);
xnor U3602 (N_3602,N_3548,N_3153);
nor U3603 (N_3603,N_3254,N_3097);
and U3604 (N_3604,N_3553,N_3147);
xnor U3605 (N_3605,N_3394,N_3032);
xnor U3606 (N_3606,N_3229,N_3322);
and U3607 (N_3607,N_3277,N_3351);
nand U3608 (N_3608,N_3256,N_3034);
nand U3609 (N_3609,N_3067,N_3243);
and U3610 (N_3610,N_3207,N_3534);
and U3611 (N_3611,N_3455,N_3055);
nand U3612 (N_3612,N_3048,N_3154);
nor U3613 (N_3613,N_3536,N_3279);
nand U3614 (N_3614,N_3598,N_3135);
and U3615 (N_3615,N_3327,N_3571);
nor U3616 (N_3616,N_3562,N_3462);
and U3617 (N_3617,N_3070,N_3266);
or U3618 (N_3618,N_3306,N_3194);
xor U3619 (N_3619,N_3555,N_3586);
and U3620 (N_3620,N_3384,N_3165);
nand U3621 (N_3621,N_3596,N_3551);
nor U3622 (N_3622,N_3374,N_3131);
xnor U3623 (N_3623,N_3486,N_3017);
or U3624 (N_3624,N_3525,N_3444);
and U3625 (N_3625,N_3281,N_3578);
and U3626 (N_3626,N_3508,N_3356);
nor U3627 (N_3627,N_3523,N_3205);
xnor U3628 (N_3628,N_3181,N_3357);
or U3629 (N_3629,N_3474,N_3469);
and U3630 (N_3630,N_3128,N_3101);
nand U3631 (N_3631,N_3299,N_3366);
or U3632 (N_3632,N_3113,N_3592);
nor U3633 (N_3633,N_3099,N_3115);
nor U3634 (N_3634,N_3259,N_3533);
xnor U3635 (N_3635,N_3236,N_3359);
xnor U3636 (N_3636,N_3352,N_3290);
nor U3637 (N_3637,N_3163,N_3188);
or U3638 (N_3638,N_3164,N_3583);
or U3639 (N_3639,N_3334,N_3513);
nand U3640 (N_3640,N_3541,N_3521);
nand U3641 (N_3641,N_3363,N_3439);
nor U3642 (N_3642,N_3544,N_3192);
nor U3643 (N_3643,N_3071,N_3265);
or U3644 (N_3644,N_3104,N_3076);
or U3645 (N_3645,N_3517,N_3196);
or U3646 (N_3646,N_3567,N_3464);
nor U3647 (N_3647,N_3200,N_3214);
nor U3648 (N_3648,N_3020,N_3354);
and U3649 (N_3649,N_3095,N_3509);
xnor U3650 (N_3650,N_3287,N_3230);
nor U3651 (N_3651,N_3162,N_3410);
nor U3652 (N_3652,N_3011,N_3185);
xor U3653 (N_3653,N_3554,N_3589);
or U3654 (N_3654,N_3199,N_3002);
and U3655 (N_3655,N_3221,N_3402);
nand U3656 (N_3656,N_3244,N_3240);
or U3657 (N_3657,N_3062,N_3143);
or U3658 (N_3658,N_3460,N_3297);
and U3659 (N_3659,N_3547,N_3431);
or U3660 (N_3660,N_3543,N_3072);
or U3661 (N_3661,N_3187,N_3039);
nand U3662 (N_3662,N_3408,N_3052);
and U3663 (N_3663,N_3272,N_3390);
or U3664 (N_3664,N_3376,N_3325);
or U3665 (N_3665,N_3186,N_3159);
and U3666 (N_3666,N_3137,N_3506);
nand U3667 (N_3667,N_3420,N_3545);
nor U3668 (N_3668,N_3251,N_3443);
xor U3669 (N_3669,N_3475,N_3549);
or U3670 (N_3670,N_3057,N_3546);
nand U3671 (N_3671,N_3247,N_3177);
and U3672 (N_3672,N_3078,N_3249);
or U3673 (N_3673,N_3255,N_3489);
nand U3674 (N_3674,N_3063,N_3428);
xor U3675 (N_3675,N_3216,N_3454);
xnor U3676 (N_3676,N_3447,N_3211);
nor U3677 (N_3677,N_3528,N_3274);
nor U3678 (N_3678,N_3465,N_3360);
xor U3679 (N_3679,N_3395,N_3479);
and U3680 (N_3680,N_3416,N_3463);
and U3681 (N_3681,N_3233,N_3422);
nor U3682 (N_3682,N_3096,N_3145);
nor U3683 (N_3683,N_3350,N_3576);
or U3684 (N_3684,N_3250,N_3550);
xnor U3685 (N_3685,N_3396,N_3347);
nand U3686 (N_3686,N_3314,N_3086);
nor U3687 (N_3687,N_3556,N_3468);
nand U3688 (N_3688,N_3488,N_3049);
nand U3689 (N_3689,N_3507,N_3239);
xor U3690 (N_3690,N_3029,N_3263);
nand U3691 (N_3691,N_3497,N_3080);
or U3692 (N_3692,N_3111,N_3203);
nor U3693 (N_3693,N_3579,N_3175);
nand U3694 (N_3694,N_3433,N_3313);
xor U3695 (N_3695,N_3245,N_3529);
nand U3696 (N_3696,N_3380,N_3105);
nor U3697 (N_3697,N_3599,N_3167);
xnor U3698 (N_3698,N_3225,N_3491);
nand U3699 (N_3699,N_3574,N_3157);
and U3700 (N_3700,N_3499,N_3150);
xnor U3701 (N_3701,N_3492,N_3442);
and U3702 (N_3702,N_3471,N_3064);
nand U3703 (N_3703,N_3127,N_3120);
xnor U3704 (N_3704,N_3090,N_3558);
or U3705 (N_3705,N_3031,N_3432);
xnor U3706 (N_3706,N_3224,N_3344);
or U3707 (N_3707,N_3172,N_3461);
xor U3708 (N_3708,N_3594,N_3386);
or U3709 (N_3709,N_3414,N_3392);
or U3710 (N_3710,N_3066,N_3282);
nand U3711 (N_3711,N_3368,N_3398);
xor U3712 (N_3712,N_3595,N_3341);
nand U3713 (N_3713,N_3208,N_3301);
and U3714 (N_3714,N_3478,N_3114);
nor U3715 (N_3715,N_3160,N_3535);
xor U3716 (N_3716,N_3530,N_3424);
xor U3717 (N_3717,N_3019,N_3449);
xor U3718 (N_3718,N_3112,N_3005);
and U3719 (N_3719,N_3570,N_3563);
and U3720 (N_3720,N_3093,N_3219);
nor U3721 (N_3721,N_3531,N_3401);
or U3722 (N_3722,N_3580,N_3082);
nand U3723 (N_3723,N_3081,N_3210);
nand U3724 (N_3724,N_3333,N_3271);
nor U3725 (N_3725,N_3527,N_3045);
and U3726 (N_3726,N_3448,N_3496);
xor U3727 (N_3727,N_3425,N_3267);
nor U3728 (N_3728,N_3413,N_3260);
xnor U3729 (N_3729,N_3537,N_3291);
nor U3730 (N_3730,N_3283,N_3107);
or U3731 (N_3731,N_3053,N_3015);
nor U3732 (N_3732,N_3332,N_3407);
or U3733 (N_3733,N_3252,N_3298);
or U3734 (N_3734,N_3047,N_3557);
nor U3735 (N_3735,N_3126,N_3069);
and U3736 (N_3736,N_3269,N_3142);
and U3737 (N_3737,N_3280,N_3387);
nand U3738 (N_3738,N_3309,N_3326);
and U3739 (N_3739,N_3445,N_3370);
or U3740 (N_3740,N_3028,N_3430);
nor U3741 (N_3741,N_3305,N_3382);
nand U3742 (N_3742,N_3423,N_3593);
nor U3743 (N_3743,N_3084,N_3399);
nor U3744 (N_3744,N_3321,N_3241);
nand U3745 (N_3745,N_3343,N_3151);
or U3746 (N_3746,N_3450,N_3195);
or U3747 (N_3747,N_3110,N_3480);
xor U3748 (N_3748,N_3191,N_3237);
nand U3749 (N_3749,N_3311,N_3060);
nand U3750 (N_3750,N_3419,N_3268);
and U3751 (N_3751,N_3565,N_3117);
xor U3752 (N_3752,N_3409,N_3498);
and U3753 (N_3753,N_3597,N_3122);
nand U3754 (N_3754,N_3415,N_3456);
or U3755 (N_3755,N_3582,N_3246);
nor U3756 (N_3756,N_3133,N_3295);
and U3757 (N_3757,N_3505,N_3440);
and U3758 (N_3758,N_3013,N_3234);
or U3759 (N_3759,N_3170,N_3391);
nand U3760 (N_3760,N_3323,N_3161);
and U3761 (N_3761,N_3538,N_3361);
nand U3762 (N_3762,N_3083,N_3477);
and U3763 (N_3763,N_3318,N_3152);
or U3764 (N_3764,N_3232,N_3103);
nor U3765 (N_3765,N_3476,N_3575);
xnor U3766 (N_3766,N_3218,N_3058);
xnor U3767 (N_3767,N_3148,N_3339);
nor U3768 (N_3768,N_3085,N_3516);
and U3769 (N_3769,N_3446,N_3046);
and U3770 (N_3770,N_3552,N_3591);
nand U3771 (N_3771,N_3176,N_3198);
nand U3772 (N_3772,N_3174,N_3515);
and U3773 (N_3773,N_3504,N_3033);
or U3774 (N_3774,N_3317,N_3561);
or U3775 (N_3775,N_3000,N_3136);
and U3776 (N_3776,N_3123,N_3532);
nor U3777 (N_3777,N_3018,N_3308);
xnor U3778 (N_3778,N_3212,N_3572);
nor U3779 (N_3779,N_3539,N_3238);
or U3780 (N_3780,N_3473,N_3560);
nand U3781 (N_3781,N_3519,N_3209);
nand U3782 (N_3782,N_3411,N_3190);
xor U3783 (N_3783,N_3073,N_3215);
nor U3784 (N_3784,N_3466,N_3088);
nand U3785 (N_3785,N_3038,N_3044);
nand U3786 (N_3786,N_3526,N_3264);
nor U3787 (N_3787,N_3118,N_3119);
nand U3788 (N_3788,N_3220,N_3418);
nand U3789 (N_3789,N_3248,N_3522);
or U3790 (N_3790,N_3481,N_3483);
nand U3791 (N_3791,N_3369,N_3008);
nor U3792 (N_3792,N_3092,N_3336);
nor U3793 (N_3793,N_3180,N_3429);
xor U3794 (N_3794,N_3041,N_3169);
nand U3795 (N_3795,N_3358,N_3542);
nand U3796 (N_3796,N_3009,N_3012);
nor U3797 (N_3797,N_3102,N_3559);
and U3798 (N_3798,N_3487,N_3304);
and U3799 (N_3799,N_3108,N_3146);
and U3800 (N_3800,N_3050,N_3184);
nor U3801 (N_3801,N_3065,N_3337);
nor U3802 (N_3802,N_3079,N_3043);
nor U3803 (N_3803,N_3149,N_3024);
or U3804 (N_3804,N_3292,N_3213);
and U3805 (N_3805,N_3087,N_3524);
nor U3806 (N_3806,N_3089,N_3338);
nand U3807 (N_3807,N_3312,N_3302);
or U3808 (N_3808,N_3438,N_3129);
or U3809 (N_3809,N_3204,N_3061);
or U3810 (N_3810,N_3023,N_3124);
nor U3811 (N_3811,N_3231,N_3502);
nor U3812 (N_3812,N_3435,N_3331);
nand U3813 (N_3813,N_3493,N_3346);
nor U3814 (N_3814,N_3141,N_3270);
or U3815 (N_3815,N_3156,N_3179);
xor U3816 (N_3816,N_3182,N_3319);
nor U3817 (N_3817,N_3037,N_3566);
and U3818 (N_3818,N_3470,N_3377);
nand U3819 (N_3819,N_3495,N_3364);
and U3820 (N_3820,N_3510,N_3345);
xor U3821 (N_3821,N_3193,N_3383);
and U3822 (N_3822,N_3016,N_3036);
and U3823 (N_3823,N_3042,N_3168);
nor U3824 (N_3824,N_3132,N_3257);
xnor U3825 (N_3825,N_3276,N_3371);
nand U3826 (N_3826,N_3511,N_3348);
or U3827 (N_3827,N_3501,N_3140);
or U3828 (N_3828,N_3125,N_3166);
nand U3829 (N_3829,N_3378,N_3242);
or U3830 (N_3830,N_3590,N_3278);
or U3831 (N_3831,N_3288,N_3421);
nor U3832 (N_3832,N_3417,N_3584);
xor U3833 (N_3833,N_3155,N_3379);
nor U3834 (N_3834,N_3006,N_3385);
and U3835 (N_3835,N_3294,N_3403);
xnor U3836 (N_3836,N_3007,N_3010);
and U3837 (N_3837,N_3217,N_3286);
xnor U3838 (N_3838,N_3427,N_3482);
nor U3839 (N_3839,N_3353,N_3178);
nand U3840 (N_3840,N_3030,N_3365);
nand U3841 (N_3841,N_3512,N_3316);
nor U3842 (N_3842,N_3300,N_3585);
and U3843 (N_3843,N_3404,N_3349);
nand U3844 (N_3844,N_3173,N_3228);
xor U3845 (N_3845,N_3202,N_3235);
nor U3846 (N_3846,N_3400,N_3441);
nor U3847 (N_3847,N_3144,N_3275);
nand U3848 (N_3848,N_3289,N_3340);
nand U3849 (N_3849,N_3106,N_3503);
and U3850 (N_3850,N_3035,N_3197);
or U3851 (N_3851,N_3569,N_3201);
and U3852 (N_3852,N_3226,N_3273);
and U3853 (N_3853,N_3452,N_3458);
xor U3854 (N_3854,N_3406,N_3121);
or U3855 (N_3855,N_3587,N_3183);
xor U3856 (N_3856,N_3320,N_3303);
nor U3857 (N_3857,N_3074,N_3258);
xor U3858 (N_3858,N_3014,N_3222);
nand U3859 (N_3859,N_3094,N_3116);
or U3860 (N_3860,N_3130,N_3310);
nor U3861 (N_3861,N_3059,N_3342);
nand U3862 (N_3862,N_3001,N_3520);
nor U3863 (N_3863,N_3581,N_3540);
and U3864 (N_3864,N_3171,N_3472);
xnor U3865 (N_3865,N_3223,N_3573);
xor U3866 (N_3866,N_3285,N_3004);
and U3867 (N_3867,N_3451,N_3412);
or U3868 (N_3868,N_3397,N_3098);
nand U3869 (N_3869,N_3324,N_3027);
nand U3870 (N_3870,N_3091,N_3025);
or U3871 (N_3871,N_3056,N_3158);
nand U3872 (N_3872,N_3484,N_3075);
nand U3873 (N_3873,N_3588,N_3329);
xnor U3874 (N_3874,N_3315,N_3330);
and U3875 (N_3875,N_3189,N_3453);
nand U3876 (N_3876,N_3467,N_3393);
and U3877 (N_3877,N_3284,N_3054);
nor U3878 (N_3878,N_3293,N_3262);
xnor U3879 (N_3879,N_3138,N_3500);
and U3880 (N_3880,N_3003,N_3051);
nand U3881 (N_3881,N_3100,N_3434);
nand U3882 (N_3882,N_3068,N_3426);
and U3883 (N_3883,N_3373,N_3485);
nor U3884 (N_3884,N_3490,N_3261);
and U3885 (N_3885,N_3437,N_3040);
xor U3886 (N_3886,N_3568,N_3139);
and U3887 (N_3887,N_3134,N_3457);
or U3888 (N_3888,N_3436,N_3381);
nand U3889 (N_3889,N_3375,N_3227);
xnor U3890 (N_3890,N_3514,N_3518);
or U3891 (N_3891,N_3459,N_3362);
and U3892 (N_3892,N_3494,N_3335);
nor U3893 (N_3893,N_3328,N_3388);
nor U3894 (N_3894,N_3026,N_3564);
nor U3895 (N_3895,N_3577,N_3109);
nor U3896 (N_3896,N_3206,N_3372);
xor U3897 (N_3897,N_3367,N_3389);
nor U3898 (N_3898,N_3021,N_3355);
xor U3899 (N_3899,N_3405,N_3077);
or U3900 (N_3900,N_3197,N_3185);
nand U3901 (N_3901,N_3284,N_3128);
or U3902 (N_3902,N_3458,N_3188);
xnor U3903 (N_3903,N_3164,N_3336);
or U3904 (N_3904,N_3218,N_3489);
nor U3905 (N_3905,N_3160,N_3190);
xnor U3906 (N_3906,N_3021,N_3191);
xor U3907 (N_3907,N_3559,N_3409);
nor U3908 (N_3908,N_3047,N_3373);
and U3909 (N_3909,N_3367,N_3465);
nand U3910 (N_3910,N_3081,N_3190);
nor U3911 (N_3911,N_3177,N_3046);
nand U3912 (N_3912,N_3576,N_3435);
xnor U3913 (N_3913,N_3587,N_3353);
nand U3914 (N_3914,N_3400,N_3040);
xor U3915 (N_3915,N_3498,N_3193);
xor U3916 (N_3916,N_3597,N_3250);
xnor U3917 (N_3917,N_3361,N_3031);
nand U3918 (N_3918,N_3428,N_3348);
or U3919 (N_3919,N_3271,N_3263);
xnor U3920 (N_3920,N_3262,N_3032);
or U3921 (N_3921,N_3092,N_3381);
and U3922 (N_3922,N_3500,N_3077);
xnor U3923 (N_3923,N_3105,N_3455);
or U3924 (N_3924,N_3562,N_3286);
xnor U3925 (N_3925,N_3114,N_3503);
or U3926 (N_3926,N_3456,N_3082);
nand U3927 (N_3927,N_3222,N_3575);
and U3928 (N_3928,N_3205,N_3115);
and U3929 (N_3929,N_3122,N_3504);
and U3930 (N_3930,N_3502,N_3538);
and U3931 (N_3931,N_3526,N_3140);
xor U3932 (N_3932,N_3565,N_3150);
and U3933 (N_3933,N_3359,N_3184);
nand U3934 (N_3934,N_3515,N_3115);
nor U3935 (N_3935,N_3583,N_3368);
and U3936 (N_3936,N_3427,N_3195);
xor U3937 (N_3937,N_3108,N_3476);
or U3938 (N_3938,N_3098,N_3373);
and U3939 (N_3939,N_3130,N_3008);
nand U3940 (N_3940,N_3583,N_3226);
nand U3941 (N_3941,N_3086,N_3541);
xnor U3942 (N_3942,N_3308,N_3233);
nor U3943 (N_3943,N_3395,N_3065);
or U3944 (N_3944,N_3048,N_3066);
or U3945 (N_3945,N_3097,N_3101);
nand U3946 (N_3946,N_3411,N_3410);
nor U3947 (N_3947,N_3152,N_3524);
and U3948 (N_3948,N_3279,N_3494);
nand U3949 (N_3949,N_3004,N_3346);
xor U3950 (N_3950,N_3003,N_3580);
nor U3951 (N_3951,N_3380,N_3486);
nor U3952 (N_3952,N_3204,N_3039);
xnor U3953 (N_3953,N_3061,N_3433);
nor U3954 (N_3954,N_3175,N_3576);
nand U3955 (N_3955,N_3008,N_3290);
or U3956 (N_3956,N_3381,N_3251);
or U3957 (N_3957,N_3597,N_3229);
xnor U3958 (N_3958,N_3532,N_3313);
or U3959 (N_3959,N_3268,N_3467);
xnor U3960 (N_3960,N_3335,N_3104);
or U3961 (N_3961,N_3344,N_3211);
nand U3962 (N_3962,N_3459,N_3395);
nand U3963 (N_3963,N_3489,N_3270);
nor U3964 (N_3964,N_3008,N_3528);
nor U3965 (N_3965,N_3251,N_3301);
and U3966 (N_3966,N_3295,N_3026);
and U3967 (N_3967,N_3061,N_3409);
and U3968 (N_3968,N_3242,N_3124);
xor U3969 (N_3969,N_3172,N_3454);
xnor U3970 (N_3970,N_3222,N_3414);
nand U3971 (N_3971,N_3135,N_3087);
nor U3972 (N_3972,N_3102,N_3488);
xor U3973 (N_3973,N_3460,N_3521);
or U3974 (N_3974,N_3420,N_3180);
or U3975 (N_3975,N_3323,N_3535);
nand U3976 (N_3976,N_3183,N_3505);
or U3977 (N_3977,N_3256,N_3445);
xnor U3978 (N_3978,N_3065,N_3042);
or U3979 (N_3979,N_3169,N_3428);
nor U3980 (N_3980,N_3298,N_3175);
nand U3981 (N_3981,N_3100,N_3346);
and U3982 (N_3982,N_3593,N_3333);
nor U3983 (N_3983,N_3062,N_3077);
xnor U3984 (N_3984,N_3121,N_3589);
xnor U3985 (N_3985,N_3012,N_3490);
and U3986 (N_3986,N_3350,N_3502);
and U3987 (N_3987,N_3453,N_3076);
nor U3988 (N_3988,N_3448,N_3348);
or U3989 (N_3989,N_3360,N_3278);
or U3990 (N_3990,N_3186,N_3257);
xor U3991 (N_3991,N_3591,N_3260);
nand U3992 (N_3992,N_3261,N_3464);
xnor U3993 (N_3993,N_3305,N_3332);
nor U3994 (N_3994,N_3585,N_3052);
xor U3995 (N_3995,N_3302,N_3280);
or U3996 (N_3996,N_3362,N_3437);
nand U3997 (N_3997,N_3488,N_3190);
xnor U3998 (N_3998,N_3304,N_3517);
xor U3999 (N_3999,N_3418,N_3131);
xnor U4000 (N_4000,N_3288,N_3568);
nand U4001 (N_4001,N_3046,N_3315);
or U4002 (N_4002,N_3083,N_3346);
and U4003 (N_4003,N_3210,N_3200);
nor U4004 (N_4004,N_3349,N_3172);
xnor U4005 (N_4005,N_3205,N_3099);
nor U4006 (N_4006,N_3233,N_3077);
xnor U4007 (N_4007,N_3148,N_3085);
and U4008 (N_4008,N_3524,N_3574);
nor U4009 (N_4009,N_3431,N_3094);
xor U4010 (N_4010,N_3350,N_3320);
nand U4011 (N_4011,N_3328,N_3378);
and U4012 (N_4012,N_3495,N_3036);
or U4013 (N_4013,N_3082,N_3379);
or U4014 (N_4014,N_3254,N_3127);
nand U4015 (N_4015,N_3090,N_3011);
nand U4016 (N_4016,N_3557,N_3526);
and U4017 (N_4017,N_3084,N_3236);
nor U4018 (N_4018,N_3430,N_3147);
nand U4019 (N_4019,N_3152,N_3296);
or U4020 (N_4020,N_3009,N_3353);
nand U4021 (N_4021,N_3587,N_3196);
xor U4022 (N_4022,N_3285,N_3044);
and U4023 (N_4023,N_3318,N_3483);
or U4024 (N_4024,N_3278,N_3211);
and U4025 (N_4025,N_3175,N_3363);
nand U4026 (N_4026,N_3187,N_3277);
nand U4027 (N_4027,N_3524,N_3310);
xnor U4028 (N_4028,N_3335,N_3333);
and U4029 (N_4029,N_3373,N_3394);
xnor U4030 (N_4030,N_3582,N_3511);
nor U4031 (N_4031,N_3466,N_3297);
and U4032 (N_4032,N_3280,N_3411);
xor U4033 (N_4033,N_3175,N_3567);
xor U4034 (N_4034,N_3388,N_3268);
and U4035 (N_4035,N_3077,N_3001);
and U4036 (N_4036,N_3135,N_3203);
nor U4037 (N_4037,N_3496,N_3573);
nor U4038 (N_4038,N_3153,N_3150);
nand U4039 (N_4039,N_3003,N_3322);
and U4040 (N_4040,N_3504,N_3403);
nand U4041 (N_4041,N_3084,N_3199);
nor U4042 (N_4042,N_3201,N_3557);
nand U4043 (N_4043,N_3318,N_3296);
or U4044 (N_4044,N_3300,N_3370);
xor U4045 (N_4045,N_3156,N_3083);
nor U4046 (N_4046,N_3572,N_3171);
nor U4047 (N_4047,N_3037,N_3562);
and U4048 (N_4048,N_3219,N_3043);
nor U4049 (N_4049,N_3025,N_3371);
nor U4050 (N_4050,N_3213,N_3135);
nor U4051 (N_4051,N_3529,N_3078);
nor U4052 (N_4052,N_3057,N_3348);
xnor U4053 (N_4053,N_3231,N_3331);
xnor U4054 (N_4054,N_3422,N_3238);
nor U4055 (N_4055,N_3397,N_3001);
nand U4056 (N_4056,N_3434,N_3547);
nor U4057 (N_4057,N_3342,N_3023);
and U4058 (N_4058,N_3480,N_3066);
xor U4059 (N_4059,N_3408,N_3021);
and U4060 (N_4060,N_3408,N_3041);
or U4061 (N_4061,N_3035,N_3555);
xnor U4062 (N_4062,N_3287,N_3448);
and U4063 (N_4063,N_3347,N_3158);
or U4064 (N_4064,N_3352,N_3361);
nand U4065 (N_4065,N_3298,N_3465);
and U4066 (N_4066,N_3409,N_3287);
or U4067 (N_4067,N_3435,N_3226);
nand U4068 (N_4068,N_3225,N_3278);
nor U4069 (N_4069,N_3229,N_3410);
nor U4070 (N_4070,N_3351,N_3125);
xnor U4071 (N_4071,N_3297,N_3427);
xor U4072 (N_4072,N_3176,N_3266);
nor U4073 (N_4073,N_3447,N_3291);
xor U4074 (N_4074,N_3294,N_3474);
nand U4075 (N_4075,N_3444,N_3587);
or U4076 (N_4076,N_3457,N_3012);
nand U4077 (N_4077,N_3355,N_3315);
or U4078 (N_4078,N_3035,N_3060);
nand U4079 (N_4079,N_3466,N_3280);
or U4080 (N_4080,N_3386,N_3080);
xnor U4081 (N_4081,N_3406,N_3405);
or U4082 (N_4082,N_3580,N_3467);
nor U4083 (N_4083,N_3583,N_3089);
nor U4084 (N_4084,N_3319,N_3300);
nand U4085 (N_4085,N_3245,N_3334);
xnor U4086 (N_4086,N_3081,N_3304);
or U4087 (N_4087,N_3242,N_3472);
and U4088 (N_4088,N_3175,N_3510);
or U4089 (N_4089,N_3330,N_3483);
xor U4090 (N_4090,N_3208,N_3074);
nand U4091 (N_4091,N_3205,N_3089);
nor U4092 (N_4092,N_3114,N_3558);
nor U4093 (N_4093,N_3452,N_3333);
xnor U4094 (N_4094,N_3138,N_3368);
nand U4095 (N_4095,N_3400,N_3340);
nand U4096 (N_4096,N_3249,N_3388);
nor U4097 (N_4097,N_3128,N_3270);
nand U4098 (N_4098,N_3330,N_3148);
or U4099 (N_4099,N_3200,N_3265);
nor U4100 (N_4100,N_3375,N_3286);
nor U4101 (N_4101,N_3424,N_3545);
and U4102 (N_4102,N_3016,N_3590);
xor U4103 (N_4103,N_3469,N_3535);
nand U4104 (N_4104,N_3569,N_3546);
or U4105 (N_4105,N_3155,N_3498);
nand U4106 (N_4106,N_3420,N_3221);
nor U4107 (N_4107,N_3304,N_3327);
nand U4108 (N_4108,N_3144,N_3495);
and U4109 (N_4109,N_3206,N_3061);
and U4110 (N_4110,N_3020,N_3528);
or U4111 (N_4111,N_3481,N_3401);
nor U4112 (N_4112,N_3330,N_3425);
or U4113 (N_4113,N_3554,N_3213);
and U4114 (N_4114,N_3380,N_3344);
nand U4115 (N_4115,N_3019,N_3432);
nor U4116 (N_4116,N_3094,N_3125);
and U4117 (N_4117,N_3112,N_3539);
xor U4118 (N_4118,N_3108,N_3092);
and U4119 (N_4119,N_3256,N_3203);
nor U4120 (N_4120,N_3145,N_3253);
nor U4121 (N_4121,N_3410,N_3110);
or U4122 (N_4122,N_3470,N_3368);
or U4123 (N_4123,N_3016,N_3346);
xor U4124 (N_4124,N_3115,N_3261);
nor U4125 (N_4125,N_3020,N_3039);
nor U4126 (N_4126,N_3260,N_3142);
nor U4127 (N_4127,N_3265,N_3154);
and U4128 (N_4128,N_3567,N_3024);
or U4129 (N_4129,N_3534,N_3373);
and U4130 (N_4130,N_3244,N_3154);
nor U4131 (N_4131,N_3092,N_3444);
nand U4132 (N_4132,N_3580,N_3055);
and U4133 (N_4133,N_3542,N_3225);
nand U4134 (N_4134,N_3049,N_3156);
and U4135 (N_4135,N_3549,N_3224);
nand U4136 (N_4136,N_3523,N_3195);
or U4137 (N_4137,N_3138,N_3306);
nor U4138 (N_4138,N_3067,N_3131);
nor U4139 (N_4139,N_3413,N_3363);
xnor U4140 (N_4140,N_3013,N_3275);
and U4141 (N_4141,N_3094,N_3184);
nand U4142 (N_4142,N_3332,N_3284);
and U4143 (N_4143,N_3362,N_3267);
xnor U4144 (N_4144,N_3320,N_3417);
and U4145 (N_4145,N_3415,N_3455);
nand U4146 (N_4146,N_3243,N_3498);
nand U4147 (N_4147,N_3301,N_3253);
nor U4148 (N_4148,N_3451,N_3016);
nand U4149 (N_4149,N_3444,N_3300);
nor U4150 (N_4150,N_3087,N_3293);
xnor U4151 (N_4151,N_3336,N_3444);
and U4152 (N_4152,N_3576,N_3331);
or U4153 (N_4153,N_3055,N_3097);
and U4154 (N_4154,N_3202,N_3281);
nand U4155 (N_4155,N_3000,N_3187);
and U4156 (N_4156,N_3364,N_3424);
and U4157 (N_4157,N_3386,N_3042);
nand U4158 (N_4158,N_3309,N_3025);
or U4159 (N_4159,N_3278,N_3174);
nor U4160 (N_4160,N_3414,N_3365);
nor U4161 (N_4161,N_3539,N_3394);
and U4162 (N_4162,N_3530,N_3248);
and U4163 (N_4163,N_3316,N_3356);
xnor U4164 (N_4164,N_3127,N_3292);
or U4165 (N_4165,N_3581,N_3064);
xnor U4166 (N_4166,N_3515,N_3477);
nor U4167 (N_4167,N_3451,N_3527);
nand U4168 (N_4168,N_3105,N_3576);
xnor U4169 (N_4169,N_3193,N_3073);
nand U4170 (N_4170,N_3488,N_3005);
xnor U4171 (N_4171,N_3234,N_3564);
and U4172 (N_4172,N_3557,N_3149);
and U4173 (N_4173,N_3356,N_3433);
or U4174 (N_4174,N_3589,N_3113);
or U4175 (N_4175,N_3260,N_3321);
nor U4176 (N_4176,N_3211,N_3402);
or U4177 (N_4177,N_3121,N_3320);
and U4178 (N_4178,N_3017,N_3364);
nand U4179 (N_4179,N_3168,N_3023);
or U4180 (N_4180,N_3582,N_3128);
xnor U4181 (N_4181,N_3186,N_3516);
xor U4182 (N_4182,N_3297,N_3451);
and U4183 (N_4183,N_3056,N_3439);
and U4184 (N_4184,N_3063,N_3569);
and U4185 (N_4185,N_3143,N_3012);
nor U4186 (N_4186,N_3107,N_3457);
nand U4187 (N_4187,N_3256,N_3101);
xor U4188 (N_4188,N_3383,N_3390);
nand U4189 (N_4189,N_3369,N_3462);
nand U4190 (N_4190,N_3483,N_3540);
nor U4191 (N_4191,N_3112,N_3145);
nor U4192 (N_4192,N_3500,N_3090);
nor U4193 (N_4193,N_3158,N_3502);
or U4194 (N_4194,N_3336,N_3152);
nand U4195 (N_4195,N_3534,N_3354);
nor U4196 (N_4196,N_3290,N_3257);
nor U4197 (N_4197,N_3110,N_3271);
and U4198 (N_4198,N_3009,N_3369);
or U4199 (N_4199,N_3126,N_3325);
nor U4200 (N_4200,N_4025,N_4040);
nor U4201 (N_4201,N_3835,N_4139);
nand U4202 (N_4202,N_4169,N_3745);
xor U4203 (N_4203,N_3830,N_4074);
and U4204 (N_4204,N_3717,N_3767);
nand U4205 (N_4205,N_3740,N_4160);
and U4206 (N_4206,N_3960,N_4177);
nor U4207 (N_4207,N_3875,N_4056);
or U4208 (N_4208,N_4149,N_4179);
and U4209 (N_4209,N_3999,N_3618);
xnor U4210 (N_4210,N_3696,N_3751);
and U4211 (N_4211,N_3866,N_3724);
nor U4212 (N_4212,N_3954,N_4109);
nor U4213 (N_4213,N_3733,N_3632);
or U4214 (N_4214,N_3901,N_3915);
nor U4215 (N_4215,N_3821,N_3814);
and U4216 (N_4216,N_4112,N_3837);
or U4217 (N_4217,N_3785,N_3721);
nand U4218 (N_4218,N_4061,N_3601);
nor U4219 (N_4219,N_3797,N_3886);
xnor U4220 (N_4220,N_4104,N_3738);
and U4221 (N_4221,N_3896,N_4119);
and U4222 (N_4222,N_3925,N_3661);
nor U4223 (N_4223,N_3776,N_3613);
xnor U4224 (N_4224,N_3929,N_4063);
and U4225 (N_4225,N_3774,N_3640);
and U4226 (N_4226,N_3863,N_3719);
nand U4227 (N_4227,N_3757,N_4143);
nand U4228 (N_4228,N_4062,N_4133);
nand U4229 (N_4229,N_3827,N_3743);
nor U4230 (N_4230,N_3968,N_4186);
nand U4231 (N_4231,N_3769,N_3622);
nand U4232 (N_4232,N_4069,N_3957);
and U4233 (N_4233,N_3869,N_3753);
nor U4234 (N_4234,N_4092,N_3800);
nand U4235 (N_4235,N_4097,N_4084);
xnor U4236 (N_4236,N_4090,N_3679);
or U4237 (N_4237,N_4171,N_3903);
nor U4238 (N_4238,N_3712,N_3950);
and U4239 (N_4239,N_3955,N_3644);
xor U4240 (N_4240,N_3958,N_3994);
and U4241 (N_4241,N_4137,N_3676);
nor U4242 (N_4242,N_3732,N_4048);
or U4243 (N_4243,N_4014,N_4141);
or U4244 (N_4244,N_3692,N_3672);
or U4245 (N_4245,N_3897,N_3841);
nor U4246 (N_4246,N_3844,N_4181);
and U4247 (N_4247,N_3707,N_3665);
xor U4248 (N_4248,N_4106,N_3984);
xnor U4249 (N_4249,N_4178,N_4180);
nor U4250 (N_4250,N_4036,N_3891);
xnor U4251 (N_4251,N_3972,N_3671);
and U4252 (N_4252,N_4124,N_4033);
or U4253 (N_4253,N_3937,N_3723);
nand U4254 (N_4254,N_4013,N_4130);
or U4255 (N_4255,N_3771,N_4002);
and U4256 (N_4256,N_3762,N_4020);
and U4257 (N_4257,N_3736,N_4005);
nor U4258 (N_4258,N_3857,N_3605);
or U4259 (N_4259,N_3853,N_4072);
nand U4260 (N_4260,N_3971,N_3910);
and U4261 (N_4261,N_3847,N_4093);
and U4262 (N_4262,N_3775,N_3782);
and U4263 (N_4263,N_3790,N_3610);
xor U4264 (N_4264,N_3674,N_3786);
xor U4265 (N_4265,N_4032,N_3703);
and U4266 (N_4266,N_3858,N_3684);
nand U4267 (N_4267,N_3811,N_3970);
nor U4268 (N_4268,N_4144,N_3749);
nand U4269 (N_4269,N_4155,N_3752);
nor U4270 (N_4270,N_3695,N_3870);
nand U4271 (N_4271,N_3728,N_3691);
and U4272 (N_4272,N_4159,N_3667);
nor U4273 (N_4273,N_4135,N_3626);
nand U4274 (N_4274,N_3655,N_3849);
xor U4275 (N_4275,N_3922,N_4111);
or U4276 (N_4276,N_3935,N_3900);
and U4277 (N_4277,N_4076,N_3996);
xor U4278 (N_4278,N_3959,N_4000);
or U4279 (N_4279,N_4082,N_3680);
and U4280 (N_4280,N_3746,N_3889);
nor U4281 (N_4281,N_3808,N_3973);
nor U4282 (N_4282,N_3852,N_3697);
nand U4283 (N_4283,N_3908,N_3899);
or U4284 (N_4284,N_3948,N_4163);
or U4285 (N_4285,N_4140,N_4016);
or U4286 (N_4286,N_3986,N_3780);
nand U4287 (N_4287,N_3918,N_3832);
nor U4288 (N_4288,N_3739,N_3798);
nor U4289 (N_4289,N_3768,N_3947);
nand U4290 (N_4290,N_3998,N_3962);
and U4291 (N_4291,N_3704,N_3627);
nor U4292 (N_4292,N_3611,N_4158);
nor U4293 (N_4293,N_3628,N_3887);
nor U4294 (N_4294,N_3823,N_3839);
nor U4295 (N_4295,N_3854,N_3729);
or U4296 (N_4296,N_3845,N_3735);
xnor U4297 (N_4297,N_3687,N_4151);
xor U4298 (N_4298,N_3609,N_4129);
xor U4299 (N_4299,N_4191,N_3754);
xnor U4300 (N_4300,N_3834,N_4168);
xor U4301 (N_4301,N_3791,N_3734);
and U4302 (N_4302,N_4037,N_4156);
or U4303 (N_4303,N_3690,N_4096);
and U4304 (N_4304,N_4075,N_4022);
and U4305 (N_4305,N_3942,N_3931);
nand U4306 (N_4306,N_3612,N_4049);
and U4307 (N_4307,N_4136,N_4194);
xor U4308 (N_4308,N_3877,N_3822);
nand U4309 (N_4309,N_3843,N_3944);
or U4310 (N_4310,N_3916,N_3964);
nor U4311 (N_4311,N_4054,N_3792);
and U4312 (N_4312,N_4028,N_4043);
nand U4313 (N_4313,N_3698,N_3961);
xnor U4314 (N_4314,N_4021,N_3934);
nor U4315 (N_4315,N_3895,N_4019);
xnor U4316 (N_4316,N_3643,N_3985);
and U4317 (N_4317,N_3975,N_3726);
and U4318 (N_4318,N_3921,N_3783);
xor U4319 (N_4319,N_3639,N_3670);
nor U4320 (N_4320,N_3794,N_3705);
nand U4321 (N_4321,N_4058,N_3906);
or U4322 (N_4322,N_4121,N_4101);
nor U4323 (N_4323,N_3763,N_4070);
nand U4324 (N_4324,N_3744,N_3608);
nand U4325 (N_4325,N_4031,N_3702);
nand U4326 (N_4326,N_4066,N_3815);
nand U4327 (N_4327,N_3989,N_3966);
nand U4328 (N_4328,N_3936,N_4175);
xor U4329 (N_4329,N_3983,N_3820);
nand U4330 (N_4330,N_3646,N_4107);
xnor U4331 (N_4331,N_4118,N_3997);
nand U4332 (N_4332,N_4162,N_3758);
and U4333 (N_4333,N_4077,N_3663);
or U4334 (N_4334,N_3805,N_3833);
xnor U4335 (N_4335,N_4166,N_4017);
and U4336 (N_4336,N_3913,N_4164);
and U4337 (N_4337,N_3750,N_3842);
nand U4338 (N_4338,N_3779,N_3812);
xnor U4339 (N_4339,N_3658,N_4195);
or U4340 (N_4340,N_3874,N_4035);
xnor U4341 (N_4341,N_3810,N_4059);
xor U4342 (N_4342,N_3720,N_3642);
or U4343 (N_4343,N_3713,N_3930);
xnor U4344 (N_4344,N_4198,N_3772);
xor U4345 (N_4345,N_4192,N_3988);
nor U4346 (N_4346,N_3657,N_3796);
or U4347 (N_4347,N_3678,N_4081);
or U4348 (N_4348,N_3991,N_3864);
xor U4349 (N_4349,N_4008,N_3876);
nor U4350 (N_4350,N_3621,N_3880);
nand U4351 (N_4351,N_3619,N_4038);
nand U4352 (N_4352,N_3607,N_4188);
and U4353 (N_4353,N_3755,N_3664);
nor U4354 (N_4354,N_3917,N_3836);
or U4355 (N_4355,N_4123,N_3855);
xor U4356 (N_4356,N_4095,N_4086);
nand U4357 (N_4357,N_4170,N_4091);
or U4358 (N_4358,N_3699,N_3969);
xnor U4359 (N_4359,N_3708,N_3795);
nand U4360 (N_4360,N_3629,N_3993);
xnor U4361 (N_4361,N_3635,N_3606);
xnor U4362 (N_4362,N_4146,N_3881);
or U4363 (N_4363,N_3741,N_3920);
and U4364 (N_4364,N_3883,N_3894);
nand U4365 (N_4365,N_3617,N_3828);
nand U4366 (N_4366,N_3825,N_4065);
xor U4367 (N_4367,N_4055,N_3689);
nor U4368 (N_4368,N_3788,N_3807);
xor U4369 (N_4369,N_3760,N_4190);
nor U4370 (N_4370,N_4087,N_4060);
xnor U4371 (N_4371,N_3904,N_4183);
nor U4372 (N_4372,N_3861,N_4006);
nor U4373 (N_4373,N_3649,N_3681);
or U4374 (N_4374,N_3818,N_3761);
xnor U4375 (N_4375,N_3784,N_3919);
xor U4376 (N_4376,N_3995,N_3848);
nor U4377 (N_4377,N_4100,N_3846);
or U4378 (N_4378,N_3816,N_3871);
xnor U4379 (N_4379,N_3953,N_3789);
nand U4380 (N_4380,N_3980,N_3778);
nor U4381 (N_4381,N_3802,N_4080);
nand U4382 (N_4382,N_4173,N_4128);
or U4383 (N_4383,N_3781,N_3927);
nor U4384 (N_4384,N_4126,N_4131);
or U4385 (N_4385,N_4051,N_4157);
nand U4386 (N_4386,N_4122,N_3716);
nor U4387 (N_4387,N_3614,N_3987);
nor U4388 (N_4388,N_4068,N_4161);
or U4389 (N_4389,N_4153,N_3799);
or U4390 (N_4390,N_3648,N_3709);
and U4391 (N_4391,N_3867,N_3653);
nor U4392 (N_4392,N_4120,N_4125);
and U4393 (N_4393,N_3890,N_3694);
xor U4394 (N_4394,N_3773,N_3862);
and U4395 (N_4395,N_3838,N_3911);
and U4396 (N_4396,N_3748,N_4067);
or U4397 (N_4397,N_3706,N_4046);
nor U4398 (N_4398,N_3888,N_4113);
nand U4399 (N_4399,N_3727,N_3637);
xor U4400 (N_4400,N_4148,N_3764);
nor U4401 (N_4401,N_4057,N_4024);
xnor U4402 (N_4402,N_3662,N_4071);
nor U4403 (N_4403,N_3647,N_4199);
nand U4404 (N_4404,N_4172,N_3759);
and U4405 (N_4405,N_4083,N_3860);
xor U4406 (N_4406,N_3616,N_3809);
xor U4407 (N_4407,N_4154,N_3868);
and U4408 (N_4408,N_3685,N_4174);
or U4409 (N_4409,N_4009,N_3976);
or U4410 (N_4410,N_3878,N_4018);
and U4411 (N_4411,N_3872,N_3829);
nand U4412 (N_4412,N_4189,N_3656);
nand U4413 (N_4413,N_3912,N_3625);
xnor U4414 (N_4414,N_3892,N_3824);
nor U4415 (N_4415,N_3949,N_3683);
nor U4416 (N_4416,N_4114,N_3806);
xnor U4417 (N_4417,N_4150,N_4027);
xnor U4418 (N_4418,N_3873,N_3715);
or U4419 (N_4419,N_4089,N_4039);
or U4420 (N_4420,N_3893,N_3659);
and U4421 (N_4421,N_4102,N_3725);
and U4422 (N_4422,N_3951,N_4176);
nor U4423 (N_4423,N_3851,N_3940);
and U4424 (N_4424,N_3840,N_3965);
and U4425 (N_4425,N_3700,N_3787);
and U4426 (N_4426,N_4004,N_3882);
or U4427 (N_4427,N_4015,N_3933);
nor U4428 (N_4428,N_3850,N_3979);
or U4429 (N_4429,N_3620,N_4108);
xor U4430 (N_4430,N_4034,N_4132);
and U4431 (N_4431,N_4110,N_3722);
nand U4432 (N_4432,N_3943,N_3765);
xor U4433 (N_4433,N_3660,N_3926);
or U4434 (N_4434,N_3652,N_3928);
or U4435 (N_4435,N_4115,N_4094);
or U4436 (N_4436,N_4073,N_3615);
nor U4437 (N_4437,N_4029,N_3819);
nand U4438 (N_4438,N_3756,N_3666);
and U4439 (N_4439,N_3938,N_4023);
nor U4440 (N_4440,N_4117,N_4187);
nor U4441 (N_4441,N_4138,N_3677);
and U4442 (N_4442,N_3711,N_4003);
nor U4443 (N_4443,N_4085,N_4182);
or U4444 (N_4444,N_3766,N_3956);
xor U4445 (N_4445,N_4052,N_4142);
xor U4446 (N_4446,N_3793,N_4050);
or U4447 (N_4447,N_4001,N_4165);
xor U4448 (N_4448,N_4064,N_3826);
xnor U4449 (N_4449,N_3604,N_3701);
nor U4450 (N_4450,N_3638,N_3777);
nand U4451 (N_4451,N_3714,N_3817);
and U4452 (N_4452,N_4041,N_3630);
nor U4453 (N_4453,N_3693,N_3932);
and U4454 (N_4454,N_4011,N_3742);
and U4455 (N_4455,N_4134,N_3982);
nor U4456 (N_4456,N_4185,N_3902);
nor U4457 (N_4457,N_3686,N_3600);
xor U4458 (N_4458,N_3668,N_3654);
xor U4459 (N_4459,N_3946,N_3945);
nor U4460 (N_4460,N_3804,N_3624);
or U4461 (N_4461,N_3633,N_3905);
or U4462 (N_4462,N_4053,N_3885);
or U4463 (N_4463,N_3641,N_4152);
or U4464 (N_4464,N_3770,N_4088);
xnor U4465 (N_4465,N_3924,N_3831);
nand U4466 (N_4466,N_3631,N_3813);
nand U4467 (N_4467,N_3651,N_3688);
nor U4468 (N_4468,N_3923,N_3675);
or U4469 (N_4469,N_4105,N_3737);
nor U4470 (N_4470,N_4098,N_3673);
and U4471 (N_4471,N_3710,N_3731);
and U4472 (N_4472,N_4026,N_3939);
or U4473 (N_4473,N_3603,N_4042);
nand U4474 (N_4474,N_3682,N_3992);
or U4475 (N_4475,N_4145,N_4007);
xor U4476 (N_4476,N_4044,N_3718);
nor U4477 (N_4477,N_4196,N_4099);
nand U4478 (N_4478,N_4012,N_4116);
nor U4479 (N_4479,N_3859,N_3803);
and U4480 (N_4480,N_3636,N_3884);
xor U4481 (N_4481,N_4030,N_4103);
xor U4482 (N_4482,N_4127,N_3879);
or U4483 (N_4483,N_3963,N_4167);
and U4484 (N_4484,N_3967,N_3669);
and U4485 (N_4485,N_4193,N_3909);
xnor U4486 (N_4486,N_3645,N_3856);
nand U4487 (N_4487,N_3977,N_4078);
or U4488 (N_4488,N_3952,N_3978);
xor U4489 (N_4489,N_3634,N_3898);
nand U4490 (N_4490,N_3907,N_3990);
nand U4491 (N_4491,N_4010,N_4047);
nor U4492 (N_4492,N_4147,N_3941);
and U4493 (N_4493,N_3602,N_4197);
nor U4494 (N_4494,N_3650,N_4184);
and U4495 (N_4495,N_3865,N_3747);
xor U4496 (N_4496,N_3623,N_3801);
nand U4497 (N_4497,N_3730,N_4045);
xnor U4498 (N_4498,N_3914,N_3974);
or U4499 (N_4499,N_4079,N_3981);
nand U4500 (N_4500,N_3937,N_3674);
or U4501 (N_4501,N_3809,N_4113);
nand U4502 (N_4502,N_3951,N_3601);
nand U4503 (N_4503,N_3978,N_4098);
xnor U4504 (N_4504,N_4090,N_4157);
nor U4505 (N_4505,N_3810,N_4145);
nor U4506 (N_4506,N_3640,N_4112);
nand U4507 (N_4507,N_3734,N_4142);
nor U4508 (N_4508,N_3674,N_3934);
and U4509 (N_4509,N_3707,N_4146);
nand U4510 (N_4510,N_4107,N_3866);
and U4511 (N_4511,N_3980,N_3615);
xor U4512 (N_4512,N_4112,N_3873);
xor U4513 (N_4513,N_3933,N_3944);
nand U4514 (N_4514,N_3744,N_3904);
and U4515 (N_4515,N_3914,N_3858);
xnor U4516 (N_4516,N_3855,N_4174);
nand U4517 (N_4517,N_3773,N_3846);
nor U4518 (N_4518,N_3613,N_3638);
nand U4519 (N_4519,N_3902,N_3882);
xnor U4520 (N_4520,N_3679,N_3755);
nand U4521 (N_4521,N_4164,N_3750);
nand U4522 (N_4522,N_3758,N_3711);
xor U4523 (N_4523,N_3960,N_3849);
xnor U4524 (N_4524,N_3944,N_3754);
xnor U4525 (N_4525,N_3915,N_3780);
nand U4526 (N_4526,N_3932,N_3681);
xnor U4527 (N_4527,N_3832,N_3767);
xnor U4528 (N_4528,N_3749,N_3868);
and U4529 (N_4529,N_3996,N_4085);
nor U4530 (N_4530,N_4113,N_3654);
nor U4531 (N_4531,N_4166,N_3726);
nand U4532 (N_4532,N_4121,N_3969);
or U4533 (N_4533,N_4045,N_3658);
and U4534 (N_4534,N_3638,N_4013);
nand U4535 (N_4535,N_3665,N_4010);
nand U4536 (N_4536,N_3757,N_3747);
nor U4537 (N_4537,N_4007,N_3956);
nor U4538 (N_4538,N_4074,N_3763);
nand U4539 (N_4539,N_3735,N_3743);
or U4540 (N_4540,N_3985,N_3923);
nand U4541 (N_4541,N_3999,N_3798);
and U4542 (N_4542,N_3714,N_3721);
or U4543 (N_4543,N_3816,N_3712);
and U4544 (N_4544,N_4197,N_3932);
or U4545 (N_4545,N_3995,N_4078);
nand U4546 (N_4546,N_3980,N_3814);
and U4547 (N_4547,N_4039,N_3690);
xnor U4548 (N_4548,N_4018,N_3903);
or U4549 (N_4549,N_3903,N_3638);
nand U4550 (N_4550,N_4149,N_3632);
nor U4551 (N_4551,N_4049,N_3972);
and U4552 (N_4552,N_4052,N_3999);
xor U4553 (N_4553,N_3604,N_3826);
nor U4554 (N_4554,N_3996,N_3613);
nor U4555 (N_4555,N_4125,N_4051);
nor U4556 (N_4556,N_3771,N_3652);
nand U4557 (N_4557,N_3768,N_3825);
nor U4558 (N_4558,N_3961,N_4195);
nor U4559 (N_4559,N_3818,N_3826);
or U4560 (N_4560,N_3643,N_3999);
nand U4561 (N_4561,N_3754,N_3889);
xor U4562 (N_4562,N_3875,N_3609);
and U4563 (N_4563,N_3891,N_3632);
xnor U4564 (N_4564,N_3807,N_3976);
xnor U4565 (N_4565,N_4003,N_3679);
nor U4566 (N_4566,N_3989,N_3685);
nor U4567 (N_4567,N_3820,N_3655);
and U4568 (N_4568,N_3684,N_3982);
xnor U4569 (N_4569,N_3675,N_3871);
and U4570 (N_4570,N_3971,N_3636);
nor U4571 (N_4571,N_3768,N_3954);
or U4572 (N_4572,N_3644,N_4120);
xor U4573 (N_4573,N_3877,N_3814);
and U4574 (N_4574,N_4187,N_3665);
xor U4575 (N_4575,N_4002,N_3886);
nand U4576 (N_4576,N_4176,N_3759);
xor U4577 (N_4577,N_4118,N_4084);
xnor U4578 (N_4578,N_3954,N_3905);
xor U4579 (N_4579,N_4008,N_4109);
or U4580 (N_4580,N_3993,N_3833);
xnor U4581 (N_4581,N_3875,N_3674);
and U4582 (N_4582,N_3759,N_3926);
nor U4583 (N_4583,N_3903,N_3769);
xnor U4584 (N_4584,N_4186,N_3919);
nand U4585 (N_4585,N_3821,N_4192);
nor U4586 (N_4586,N_4071,N_3721);
and U4587 (N_4587,N_3957,N_3931);
nor U4588 (N_4588,N_3619,N_3691);
nand U4589 (N_4589,N_3947,N_4196);
nor U4590 (N_4590,N_4197,N_3611);
nor U4591 (N_4591,N_4049,N_3664);
xnor U4592 (N_4592,N_4085,N_4007);
xnor U4593 (N_4593,N_4048,N_4044);
nand U4594 (N_4594,N_3989,N_4144);
xnor U4595 (N_4595,N_3641,N_3694);
xor U4596 (N_4596,N_3809,N_3640);
nor U4597 (N_4597,N_3809,N_4036);
or U4598 (N_4598,N_4070,N_3651);
nor U4599 (N_4599,N_3825,N_3864);
and U4600 (N_4600,N_3919,N_3757);
nor U4601 (N_4601,N_4019,N_3915);
xor U4602 (N_4602,N_4004,N_4085);
nand U4603 (N_4603,N_3655,N_3840);
nand U4604 (N_4604,N_3978,N_3773);
nand U4605 (N_4605,N_3681,N_3692);
and U4606 (N_4606,N_3725,N_4187);
and U4607 (N_4607,N_4155,N_3884);
or U4608 (N_4608,N_3639,N_4131);
and U4609 (N_4609,N_3675,N_4018);
xnor U4610 (N_4610,N_3774,N_3951);
or U4611 (N_4611,N_3963,N_3882);
and U4612 (N_4612,N_3938,N_4182);
nor U4613 (N_4613,N_4046,N_3907);
nor U4614 (N_4614,N_3758,N_3935);
and U4615 (N_4615,N_4167,N_3925);
xor U4616 (N_4616,N_3798,N_4123);
or U4617 (N_4617,N_3672,N_3681);
nand U4618 (N_4618,N_4058,N_3676);
or U4619 (N_4619,N_4153,N_3606);
nor U4620 (N_4620,N_3684,N_4062);
nand U4621 (N_4621,N_3806,N_4025);
xor U4622 (N_4622,N_3789,N_4198);
nand U4623 (N_4623,N_3802,N_3866);
or U4624 (N_4624,N_3976,N_3603);
xnor U4625 (N_4625,N_3666,N_4130);
or U4626 (N_4626,N_3997,N_4065);
xor U4627 (N_4627,N_4179,N_3625);
xor U4628 (N_4628,N_3720,N_4154);
nor U4629 (N_4629,N_3707,N_3640);
nor U4630 (N_4630,N_3727,N_4014);
and U4631 (N_4631,N_3631,N_3945);
xor U4632 (N_4632,N_4071,N_4014);
and U4633 (N_4633,N_3983,N_3687);
and U4634 (N_4634,N_3731,N_4153);
xor U4635 (N_4635,N_4069,N_4041);
xnor U4636 (N_4636,N_3795,N_3631);
and U4637 (N_4637,N_3938,N_4106);
xnor U4638 (N_4638,N_3864,N_4173);
nor U4639 (N_4639,N_3748,N_4035);
and U4640 (N_4640,N_3800,N_4138);
and U4641 (N_4641,N_4169,N_4101);
nand U4642 (N_4642,N_3788,N_3653);
nand U4643 (N_4643,N_4072,N_4104);
or U4644 (N_4644,N_3723,N_3671);
xnor U4645 (N_4645,N_3910,N_3899);
nand U4646 (N_4646,N_4198,N_3668);
nor U4647 (N_4647,N_3896,N_3999);
and U4648 (N_4648,N_3690,N_3869);
xnor U4649 (N_4649,N_3800,N_3809);
and U4650 (N_4650,N_4059,N_3721);
and U4651 (N_4651,N_3910,N_3921);
nor U4652 (N_4652,N_3657,N_3716);
nand U4653 (N_4653,N_3680,N_3949);
or U4654 (N_4654,N_3952,N_3610);
nand U4655 (N_4655,N_3980,N_3639);
and U4656 (N_4656,N_4100,N_3849);
or U4657 (N_4657,N_4171,N_4074);
nand U4658 (N_4658,N_3635,N_3970);
and U4659 (N_4659,N_3838,N_4073);
and U4660 (N_4660,N_3946,N_4087);
xnor U4661 (N_4661,N_4195,N_3968);
nor U4662 (N_4662,N_3916,N_4060);
and U4663 (N_4663,N_3662,N_4148);
and U4664 (N_4664,N_4018,N_3749);
and U4665 (N_4665,N_4187,N_4063);
or U4666 (N_4666,N_4194,N_3953);
nand U4667 (N_4667,N_4070,N_3938);
nor U4668 (N_4668,N_3697,N_4117);
and U4669 (N_4669,N_4021,N_3962);
or U4670 (N_4670,N_3775,N_3958);
nor U4671 (N_4671,N_4028,N_4134);
and U4672 (N_4672,N_3974,N_3648);
and U4673 (N_4673,N_3639,N_3721);
and U4674 (N_4674,N_4094,N_3815);
or U4675 (N_4675,N_4085,N_3933);
and U4676 (N_4676,N_3984,N_3781);
xnor U4677 (N_4677,N_3655,N_3737);
and U4678 (N_4678,N_3935,N_3796);
and U4679 (N_4679,N_3647,N_3833);
xor U4680 (N_4680,N_3901,N_3611);
xor U4681 (N_4681,N_3908,N_3837);
or U4682 (N_4682,N_3625,N_3934);
nand U4683 (N_4683,N_4112,N_4065);
and U4684 (N_4684,N_4122,N_3811);
nand U4685 (N_4685,N_3620,N_3780);
nor U4686 (N_4686,N_4165,N_4029);
or U4687 (N_4687,N_3964,N_3845);
or U4688 (N_4688,N_4077,N_4084);
nor U4689 (N_4689,N_3859,N_3861);
nor U4690 (N_4690,N_3928,N_4117);
xor U4691 (N_4691,N_3693,N_3636);
xor U4692 (N_4692,N_3772,N_4185);
nor U4693 (N_4693,N_3877,N_4194);
nor U4694 (N_4694,N_3620,N_4163);
nor U4695 (N_4695,N_3751,N_3722);
xnor U4696 (N_4696,N_3859,N_3696);
nor U4697 (N_4697,N_3606,N_3646);
and U4698 (N_4698,N_4196,N_4177);
nand U4699 (N_4699,N_3959,N_3616);
and U4700 (N_4700,N_3725,N_4018);
or U4701 (N_4701,N_3646,N_3986);
and U4702 (N_4702,N_3711,N_3776);
xnor U4703 (N_4703,N_3715,N_4148);
nand U4704 (N_4704,N_4037,N_3840);
and U4705 (N_4705,N_4137,N_3886);
and U4706 (N_4706,N_3600,N_3651);
or U4707 (N_4707,N_3888,N_4187);
nor U4708 (N_4708,N_4004,N_4009);
or U4709 (N_4709,N_3862,N_3905);
and U4710 (N_4710,N_3674,N_3913);
xnor U4711 (N_4711,N_3936,N_3702);
nand U4712 (N_4712,N_4190,N_4105);
nand U4713 (N_4713,N_4043,N_4025);
and U4714 (N_4714,N_3704,N_3943);
and U4715 (N_4715,N_3616,N_4109);
xnor U4716 (N_4716,N_4120,N_4061);
and U4717 (N_4717,N_3671,N_4044);
or U4718 (N_4718,N_3986,N_3785);
nand U4719 (N_4719,N_3635,N_3955);
nand U4720 (N_4720,N_3896,N_3841);
xnor U4721 (N_4721,N_3712,N_3800);
xor U4722 (N_4722,N_4179,N_4050);
nor U4723 (N_4723,N_3857,N_3656);
nand U4724 (N_4724,N_3975,N_3648);
nor U4725 (N_4725,N_4048,N_3761);
xor U4726 (N_4726,N_4016,N_3772);
xor U4727 (N_4727,N_4070,N_4192);
nand U4728 (N_4728,N_4063,N_3772);
or U4729 (N_4729,N_3611,N_4172);
and U4730 (N_4730,N_3837,N_3696);
nand U4731 (N_4731,N_3959,N_4169);
nor U4732 (N_4732,N_4131,N_3981);
nor U4733 (N_4733,N_3626,N_3654);
xor U4734 (N_4734,N_3775,N_3818);
nor U4735 (N_4735,N_3782,N_3994);
or U4736 (N_4736,N_3894,N_3851);
or U4737 (N_4737,N_3932,N_3676);
nand U4738 (N_4738,N_4026,N_3919);
xor U4739 (N_4739,N_4036,N_3892);
or U4740 (N_4740,N_3999,N_4193);
and U4741 (N_4741,N_4068,N_3754);
or U4742 (N_4742,N_4035,N_3652);
xnor U4743 (N_4743,N_3738,N_3894);
nand U4744 (N_4744,N_4006,N_3802);
or U4745 (N_4745,N_3899,N_4196);
and U4746 (N_4746,N_3743,N_4084);
nand U4747 (N_4747,N_4056,N_3767);
nand U4748 (N_4748,N_4123,N_3998);
nor U4749 (N_4749,N_4015,N_4162);
or U4750 (N_4750,N_3706,N_3647);
or U4751 (N_4751,N_3798,N_4074);
nand U4752 (N_4752,N_3905,N_4046);
nand U4753 (N_4753,N_3766,N_3913);
or U4754 (N_4754,N_3666,N_4182);
xnor U4755 (N_4755,N_3723,N_3835);
or U4756 (N_4756,N_3975,N_3854);
xor U4757 (N_4757,N_3667,N_4154);
or U4758 (N_4758,N_3993,N_4066);
nand U4759 (N_4759,N_3835,N_3742);
nand U4760 (N_4760,N_3910,N_3929);
or U4761 (N_4761,N_3762,N_4143);
nand U4762 (N_4762,N_3681,N_4049);
xnor U4763 (N_4763,N_3669,N_3775);
nor U4764 (N_4764,N_3723,N_3748);
nor U4765 (N_4765,N_3799,N_3665);
nor U4766 (N_4766,N_3918,N_3931);
nor U4767 (N_4767,N_4161,N_3663);
and U4768 (N_4768,N_3931,N_4090);
nand U4769 (N_4769,N_3754,N_3689);
and U4770 (N_4770,N_3729,N_3697);
or U4771 (N_4771,N_3747,N_3666);
and U4772 (N_4772,N_3704,N_3948);
nor U4773 (N_4773,N_3791,N_3605);
and U4774 (N_4774,N_4026,N_3648);
xnor U4775 (N_4775,N_4159,N_3822);
nand U4776 (N_4776,N_3755,N_4017);
nor U4777 (N_4777,N_4111,N_3742);
and U4778 (N_4778,N_3909,N_4029);
and U4779 (N_4779,N_3630,N_3613);
nor U4780 (N_4780,N_4012,N_3855);
nor U4781 (N_4781,N_4065,N_3888);
nand U4782 (N_4782,N_3814,N_4114);
nor U4783 (N_4783,N_3973,N_4032);
and U4784 (N_4784,N_3693,N_3606);
xor U4785 (N_4785,N_3694,N_3730);
or U4786 (N_4786,N_3637,N_3710);
and U4787 (N_4787,N_4058,N_3722);
xor U4788 (N_4788,N_4071,N_3773);
xor U4789 (N_4789,N_3694,N_3939);
or U4790 (N_4790,N_4087,N_4052);
and U4791 (N_4791,N_3881,N_3919);
nor U4792 (N_4792,N_3983,N_3851);
and U4793 (N_4793,N_4132,N_4148);
and U4794 (N_4794,N_3760,N_3939);
and U4795 (N_4795,N_4148,N_3875);
nor U4796 (N_4796,N_4112,N_4022);
nor U4797 (N_4797,N_3718,N_3801);
nand U4798 (N_4798,N_4038,N_3649);
and U4799 (N_4799,N_4118,N_4039);
or U4800 (N_4800,N_4405,N_4520);
and U4801 (N_4801,N_4463,N_4652);
nor U4802 (N_4802,N_4395,N_4765);
or U4803 (N_4803,N_4289,N_4202);
or U4804 (N_4804,N_4692,N_4348);
xnor U4805 (N_4805,N_4790,N_4283);
or U4806 (N_4806,N_4236,N_4775);
nor U4807 (N_4807,N_4732,N_4339);
or U4808 (N_4808,N_4642,N_4325);
and U4809 (N_4809,N_4713,N_4263);
and U4810 (N_4810,N_4678,N_4551);
and U4811 (N_4811,N_4311,N_4739);
and U4812 (N_4812,N_4382,N_4402);
and U4813 (N_4813,N_4350,N_4466);
xor U4814 (N_4814,N_4323,N_4303);
nand U4815 (N_4815,N_4343,N_4735);
and U4816 (N_4816,N_4674,N_4508);
xnor U4817 (N_4817,N_4287,N_4273);
nor U4818 (N_4818,N_4414,N_4637);
xnor U4819 (N_4819,N_4379,N_4515);
nor U4820 (N_4820,N_4269,N_4421);
nand U4821 (N_4821,N_4424,N_4258);
nor U4822 (N_4822,N_4592,N_4222);
and U4823 (N_4823,N_4399,N_4749);
and U4824 (N_4824,N_4530,N_4361);
nand U4825 (N_4825,N_4358,N_4235);
nor U4826 (N_4826,N_4568,N_4294);
nand U4827 (N_4827,N_4688,N_4791);
and U4828 (N_4828,N_4524,N_4355);
or U4829 (N_4829,N_4366,N_4367);
or U4830 (N_4830,N_4302,N_4543);
nor U4831 (N_4831,N_4368,N_4268);
nor U4832 (N_4832,N_4756,N_4649);
xor U4833 (N_4833,N_4225,N_4449);
nand U4834 (N_4834,N_4696,N_4702);
xor U4835 (N_4835,N_4359,N_4341);
nor U4836 (N_4836,N_4392,N_4489);
xor U4837 (N_4837,N_4754,N_4586);
nand U4838 (N_4838,N_4608,N_4207);
xnor U4839 (N_4839,N_4614,N_4787);
xor U4840 (N_4840,N_4576,N_4386);
nor U4841 (N_4841,N_4435,N_4306);
and U4842 (N_4842,N_4577,N_4601);
and U4843 (N_4843,N_4354,N_4476);
xor U4844 (N_4844,N_4253,N_4540);
or U4845 (N_4845,N_4347,N_4553);
nor U4846 (N_4846,N_4535,N_4590);
nor U4847 (N_4847,N_4635,N_4747);
xnor U4848 (N_4848,N_4293,N_4667);
and U4849 (N_4849,N_4768,N_4479);
or U4850 (N_4850,N_4763,N_4709);
and U4851 (N_4851,N_4338,N_4730);
xor U4852 (N_4852,N_4721,N_4511);
xor U4853 (N_4853,N_4216,N_4701);
nand U4854 (N_4854,N_4682,N_4661);
nor U4855 (N_4855,N_4671,N_4658);
xnor U4856 (N_4856,N_4407,N_4206);
and U4857 (N_4857,N_4377,N_4786);
nor U4858 (N_4858,N_4760,N_4457);
nand U4859 (N_4859,N_4251,N_4740);
nor U4860 (N_4860,N_4643,N_4536);
nand U4861 (N_4861,N_4229,N_4334);
and U4862 (N_4862,N_4617,N_4444);
nor U4863 (N_4863,N_4410,N_4409);
xor U4864 (N_4864,N_4728,N_4537);
nand U4865 (N_4865,N_4404,N_4364);
or U4866 (N_4866,N_4591,N_4381);
and U4867 (N_4867,N_4324,N_4753);
or U4868 (N_4868,N_4498,N_4423);
and U4869 (N_4869,N_4369,N_4308);
or U4870 (N_4870,N_4351,N_4391);
xnor U4871 (N_4871,N_4356,N_4558);
nor U4872 (N_4872,N_4525,N_4434);
nor U4873 (N_4873,N_4610,N_4644);
or U4874 (N_4874,N_4388,N_4442);
or U4875 (N_4875,N_4741,N_4342);
or U4876 (N_4876,N_4465,N_4772);
or U4877 (N_4877,N_4401,N_4398);
nand U4878 (N_4878,N_4594,N_4651);
and U4879 (N_4879,N_4598,N_4440);
nand U4880 (N_4880,N_4439,N_4403);
nand U4881 (N_4881,N_4267,N_4552);
nor U4882 (N_4882,N_4290,N_4452);
and U4883 (N_4883,N_4657,N_4722);
xnor U4884 (N_4884,N_4687,N_4570);
nand U4885 (N_4885,N_4231,N_4481);
nor U4886 (N_4886,N_4213,N_4510);
xor U4887 (N_4887,N_4228,N_4232);
nand U4888 (N_4888,N_4602,N_4256);
or U4889 (N_4889,N_4646,N_4224);
xor U4890 (N_4890,N_4613,N_4242);
and U4891 (N_4891,N_4501,N_4729);
nor U4892 (N_4892,N_4545,N_4738);
nand U4893 (N_4893,N_4281,N_4420);
nand U4894 (N_4894,N_4217,N_4270);
or U4895 (N_4895,N_4566,N_4719);
or U4896 (N_4896,N_4549,N_4779);
xor U4897 (N_4897,N_4335,N_4499);
xor U4898 (N_4898,N_4711,N_4632);
and U4899 (N_4899,N_4707,N_4731);
nand U4900 (N_4900,N_4668,N_4527);
nor U4901 (N_4901,N_4659,N_4685);
or U4902 (N_4902,N_4264,N_4700);
or U4903 (N_4903,N_4336,N_4579);
nor U4904 (N_4904,N_4633,N_4265);
nand U4905 (N_4905,N_4726,N_4546);
nand U4906 (N_4906,N_4288,N_4681);
nand U4907 (N_4907,N_4345,N_4517);
and U4908 (N_4908,N_4660,N_4636);
nand U4909 (N_4909,N_4641,N_4611);
xnor U4910 (N_4910,N_4725,N_4218);
nor U4911 (N_4911,N_4792,N_4389);
or U4912 (N_4912,N_4246,N_4794);
nand U4913 (N_4913,N_4259,N_4477);
nand U4914 (N_4914,N_4745,N_4438);
xnor U4915 (N_4915,N_4560,N_4375);
nor U4916 (N_4916,N_4291,N_4203);
nand U4917 (N_4917,N_4322,N_4419);
and U4918 (N_4918,N_4349,N_4561);
or U4919 (N_4919,N_4495,N_4677);
and U4920 (N_4920,N_4390,N_4471);
xor U4921 (N_4921,N_4654,N_4534);
or U4922 (N_4922,N_4468,N_4784);
xnor U4923 (N_4923,N_4565,N_4569);
nand U4924 (N_4924,N_4396,N_4506);
and U4925 (N_4925,N_4788,N_4310);
nand U4926 (N_4926,N_4631,N_4214);
and U4927 (N_4927,N_4362,N_4412);
or U4928 (N_4928,N_4781,N_4331);
xor U4929 (N_4929,N_4445,N_4239);
or U4930 (N_4930,N_4514,N_4669);
xor U4931 (N_4931,N_4778,N_4428);
or U4932 (N_4932,N_4215,N_4647);
or U4933 (N_4933,N_4201,N_4758);
or U4934 (N_4934,N_4597,N_4799);
xnor U4935 (N_4935,N_4704,N_4662);
or U4936 (N_4936,N_4777,N_4714);
nor U4937 (N_4937,N_4575,N_4665);
or U4938 (N_4938,N_4639,N_4245);
or U4939 (N_4939,N_4488,N_4309);
nand U4940 (N_4940,N_4249,N_4528);
xor U4941 (N_4941,N_4526,N_4757);
nor U4942 (N_4942,N_4493,N_4307);
nand U4943 (N_4943,N_4798,N_4482);
and U4944 (N_4944,N_4562,N_4544);
and U4945 (N_4945,N_4504,N_4764);
nor U4946 (N_4946,N_4266,N_4491);
and U4947 (N_4947,N_4538,N_4451);
and U4948 (N_4948,N_4762,N_4630);
xor U4949 (N_4949,N_4789,N_4250);
and U4950 (N_4950,N_4378,N_4512);
nor U4951 (N_4951,N_4619,N_4433);
and U4952 (N_4952,N_4581,N_4718);
or U4953 (N_4953,N_4326,N_4737);
and U4954 (N_4954,N_4208,N_4582);
or U4955 (N_4955,N_4400,N_4712);
nor U4956 (N_4956,N_4509,N_4521);
nor U4957 (N_4957,N_4475,N_4455);
nand U4958 (N_4958,N_4411,N_4584);
and U4959 (N_4959,N_4505,N_4675);
nand U4960 (N_4960,N_4564,N_4387);
xnor U4961 (N_4961,N_4680,N_4279);
or U4962 (N_4962,N_4304,N_4703);
nand U4963 (N_4963,N_4317,N_4609);
and U4964 (N_4964,N_4430,N_4244);
nand U4965 (N_4965,N_4664,N_4241);
and U4966 (N_4966,N_4585,N_4769);
nand U4967 (N_4967,N_4766,N_4376);
and U4968 (N_4968,N_4697,N_4285);
or U4969 (N_4969,N_4655,N_4415);
or U4970 (N_4970,N_4484,N_4456);
and U4971 (N_4971,N_4698,N_4596);
xnor U4972 (N_4972,N_4605,N_4629);
nand U4973 (N_4973,N_4638,N_4461);
and U4974 (N_4974,N_4313,N_4588);
nor U4975 (N_4975,N_4785,N_4767);
and U4976 (N_4976,N_4248,N_4300);
and U4977 (N_4977,N_4755,N_4532);
nand U4978 (N_4978,N_4469,N_4417);
and U4979 (N_4979,N_4223,N_4542);
nor U4980 (N_4980,N_4612,N_4292);
nor U4981 (N_4981,N_4319,N_4274);
nand U4982 (N_4982,N_4723,N_4221);
xnor U4983 (N_4983,N_4370,N_4238);
or U4984 (N_4984,N_4793,N_4426);
xor U4985 (N_4985,N_4599,N_4795);
xor U4986 (N_4986,N_4478,N_4406);
or U4987 (N_4987,N_4333,N_4272);
xnor U4988 (N_4988,N_4571,N_4262);
and U4989 (N_4989,N_4446,N_4607);
or U4990 (N_4990,N_4284,N_4673);
or U4991 (N_4991,N_4578,N_4550);
nand U4992 (N_4992,N_4640,N_4497);
xor U4993 (N_4993,N_4751,N_4559);
or U4994 (N_4994,N_4353,N_4796);
xor U4995 (N_4995,N_4337,N_4486);
and U4996 (N_4996,N_4458,N_4467);
nand U4997 (N_4997,N_4204,N_4243);
xor U4998 (N_4998,N_4371,N_4299);
nand U4999 (N_4999,N_4522,N_4254);
nor U5000 (N_5000,N_4320,N_4234);
nand U5001 (N_5001,N_4332,N_4684);
and U5002 (N_5002,N_4305,N_4328);
or U5003 (N_5003,N_4770,N_4523);
nand U5004 (N_5004,N_4715,N_4352);
and U5005 (N_5005,N_4750,N_4459);
xnor U5006 (N_5006,N_4694,N_4436);
or U5007 (N_5007,N_4220,N_4443);
and U5008 (N_5008,N_4454,N_4393);
xnor U5009 (N_5009,N_4625,N_4472);
xnor U5010 (N_5010,N_4418,N_4260);
nand U5011 (N_5011,N_4209,N_4595);
nand U5012 (N_5012,N_4394,N_4450);
nor U5013 (N_5013,N_4464,N_4716);
nand U5014 (N_5014,N_4622,N_4363);
nand U5015 (N_5015,N_4518,N_4318);
and U5016 (N_5016,N_4425,N_4623);
nor U5017 (N_5017,N_4727,N_4494);
and U5018 (N_5018,N_4429,N_4330);
and U5019 (N_5019,N_4645,N_4321);
nor U5020 (N_5020,N_4621,N_4314);
or U5021 (N_5021,N_4567,N_4460);
and U5022 (N_5022,N_4689,N_4780);
or U5023 (N_5023,N_4298,N_4485);
and U5024 (N_5024,N_4663,N_4365);
nor U5025 (N_5025,N_4483,N_4554);
nand U5026 (N_5026,N_4670,N_4547);
and U5027 (N_5027,N_4474,N_4748);
and U5028 (N_5028,N_4502,N_4280);
or U5029 (N_5029,N_4492,N_4416);
or U5030 (N_5030,N_4752,N_4490);
and U5031 (N_5031,N_4529,N_4556);
nand U5032 (N_5032,N_4533,N_4771);
or U5033 (N_5033,N_4230,N_4301);
and U5034 (N_5034,N_4620,N_4373);
and U5035 (N_5035,N_4503,N_4587);
or U5036 (N_5036,N_4276,N_4385);
nand U5037 (N_5037,N_4761,N_4212);
nor U5038 (N_5038,N_4346,N_4743);
or U5039 (N_5039,N_4679,N_4672);
nand U5040 (N_5040,N_4531,N_4782);
or U5041 (N_5041,N_4516,N_4210);
and U5042 (N_5042,N_4773,N_4408);
or U5043 (N_5043,N_4742,N_4448);
and U5044 (N_5044,N_4686,N_4634);
nor U5045 (N_5045,N_4774,N_4470);
xnor U5046 (N_5046,N_4589,N_4447);
or U5047 (N_5047,N_4344,N_4295);
and U5048 (N_5048,N_4296,N_4710);
and U5049 (N_5049,N_4252,N_4275);
xnor U5050 (N_5050,N_4437,N_4383);
nor U5051 (N_5051,N_4441,N_4695);
nand U5052 (N_5052,N_4312,N_4211);
xor U5053 (N_5053,N_4724,N_4422);
and U5054 (N_5054,N_4776,N_4573);
nand U5055 (N_5055,N_4271,N_4513);
nor U5056 (N_5056,N_4257,N_4255);
and U5057 (N_5057,N_4519,N_4380);
nor U5058 (N_5058,N_4563,N_4432);
nor U5059 (N_5059,N_4604,N_4615);
nor U5060 (N_5060,N_4316,N_4539);
nor U5061 (N_5061,N_4720,N_4360);
xnor U5062 (N_5062,N_4431,N_4580);
nand U5063 (N_5063,N_4693,N_4487);
and U5064 (N_5064,N_4227,N_4744);
and U5065 (N_5065,N_4627,N_4691);
and U5066 (N_5066,N_4708,N_4548);
and U5067 (N_5067,N_4648,N_4297);
or U5068 (N_5068,N_4783,N_4606);
or U5069 (N_5069,N_4219,N_4600);
and U5070 (N_5070,N_4374,N_4247);
or U5071 (N_5071,N_4372,N_4656);
nand U5072 (N_5072,N_4237,N_4699);
nor U5073 (N_5073,N_4496,N_4357);
nand U5074 (N_5074,N_4500,N_4593);
nand U5075 (N_5075,N_4583,N_4555);
or U5076 (N_5076,N_4233,N_4480);
or U5077 (N_5077,N_4616,N_4462);
nor U5078 (N_5078,N_4666,N_4572);
nor U5079 (N_5079,N_4340,N_4413);
nor U5080 (N_5080,N_4286,N_4278);
xor U5081 (N_5081,N_4650,N_4734);
xor U5082 (N_5082,N_4733,N_4603);
and U5083 (N_5083,N_4706,N_4473);
and U5084 (N_5084,N_4507,N_4746);
xor U5085 (N_5085,N_4226,N_4277);
and U5086 (N_5086,N_4329,N_4427);
xnor U5087 (N_5087,N_4574,N_4541);
or U5088 (N_5088,N_4315,N_4200);
nor U5089 (N_5089,N_4557,N_4736);
xnor U5090 (N_5090,N_4384,N_4453);
or U5091 (N_5091,N_4261,N_4676);
nand U5092 (N_5092,N_4628,N_4759);
and U5093 (N_5093,N_4683,N_4717);
and U5094 (N_5094,N_4205,N_4282);
or U5095 (N_5095,N_4240,N_4705);
xor U5096 (N_5096,N_4626,N_4327);
xor U5097 (N_5097,N_4618,N_4397);
and U5098 (N_5098,N_4690,N_4653);
nor U5099 (N_5099,N_4624,N_4797);
or U5100 (N_5100,N_4265,N_4469);
or U5101 (N_5101,N_4630,N_4665);
and U5102 (N_5102,N_4469,N_4654);
nand U5103 (N_5103,N_4342,N_4604);
xnor U5104 (N_5104,N_4495,N_4519);
nor U5105 (N_5105,N_4589,N_4384);
nor U5106 (N_5106,N_4276,N_4792);
nand U5107 (N_5107,N_4725,N_4698);
xor U5108 (N_5108,N_4401,N_4446);
xor U5109 (N_5109,N_4357,N_4245);
and U5110 (N_5110,N_4246,N_4686);
or U5111 (N_5111,N_4436,N_4337);
xor U5112 (N_5112,N_4268,N_4346);
nand U5113 (N_5113,N_4207,N_4638);
xor U5114 (N_5114,N_4238,N_4342);
xnor U5115 (N_5115,N_4208,N_4241);
nor U5116 (N_5116,N_4656,N_4581);
and U5117 (N_5117,N_4477,N_4298);
and U5118 (N_5118,N_4588,N_4555);
or U5119 (N_5119,N_4747,N_4545);
and U5120 (N_5120,N_4794,N_4443);
or U5121 (N_5121,N_4422,N_4397);
nor U5122 (N_5122,N_4510,N_4527);
nand U5123 (N_5123,N_4739,N_4363);
nor U5124 (N_5124,N_4626,N_4725);
or U5125 (N_5125,N_4623,N_4358);
or U5126 (N_5126,N_4660,N_4491);
xnor U5127 (N_5127,N_4248,N_4596);
xor U5128 (N_5128,N_4715,N_4627);
and U5129 (N_5129,N_4572,N_4343);
or U5130 (N_5130,N_4321,N_4552);
and U5131 (N_5131,N_4417,N_4699);
xor U5132 (N_5132,N_4406,N_4448);
and U5133 (N_5133,N_4652,N_4599);
and U5134 (N_5134,N_4330,N_4314);
and U5135 (N_5135,N_4644,N_4377);
nor U5136 (N_5136,N_4635,N_4492);
nor U5137 (N_5137,N_4711,N_4755);
nor U5138 (N_5138,N_4377,N_4352);
or U5139 (N_5139,N_4205,N_4517);
nor U5140 (N_5140,N_4484,N_4690);
nor U5141 (N_5141,N_4460,N_4528);
and U5142 (N_5142,N_4546,N_4458);
and U5143 (N_5143,N_4722,N_4387);
nor U5144 (N_5144,N_4381,N_4693);
nand U5145 (N_5145,N_4780,N_4744);
xor U5146 (N_5146,N_4514,N_4539);
nand U5147 (N_5147,N_4320,N_4266);
nor U5148 (N_5148,N_4786,N_4645);
xnor U5149 (N_5149,N_4227,N_4265);
xnor U5150 (N_5150,N_4759,N_4603);
nor U5151 (N_5151,N_4796,N_4512);
xnor U5152 (N_5152,N_4767,N_4372);
nand U5153 (N_5153,N_4310,N_4613);
and U5154 (N_5154,N_4723,N_4352);
nor U5155 (N_5155,N_4363,N_4394);
or U5156 (N_5156,N_4566,N_4483);
nand U5157 (N_5157,N_4797,N_4501);
nand U5158 (N_5158,N_4612,N_4249);
and U5159 (N_5159,N_4640,N_4756);
xnor U5160 (N_5160,N_4246,N_4202);
nor U5161 (N_5161,N_4201,N_4678);
xnor U5162 (N_5162,N_4316,N_4238);
or U5163 (N_5163,N_4779,N_4604);
or U5164 (N_5164,N_4764,N_4347);
nand U5165 (N_5165,N_4645,N_4526);
or U5166 (N_5166,N_4599,N_4317);
and U5167 (N_5167,N_4727,N_4409);
and U5168 (N_5168,N_4229,N_4266);
nor U5169 (N_5169,N_4588,N_4396);
nor U5170 (N_5170,N_4404,N_4403);
xor U5171 (N_5171,N_4743,N_4764);
xnor U5172 (N_5172,N_4499,N_4542);
or U5173 (N_5173,N_4587,N_4396);
nor U5174 (N_5174,N_4577,N_4302);
or U5175 (N_5175,N_4246,N_4785);
and U5176 (N_5176,N_4656,N_4715);
nand U5177 (N_5177,N_4783,N_4380);
and U5178 (N_5178,N_4385,N_4626);
or U5179 (N_5179,N_4569,N_4395);
nand U5180 (N_5180,N_4466,N_4615);
and U5181 (N_5181,N_4542,N_4679);
nor U5182 (N_5182,N_4545,N_4447);
nor U5183 (N_5183,N_4565,N_4589);
xor U5184 (N_5184,N_4631,N_4675);
or U5185 (N_5185,N_4505,N_4338);
or U5186 (N_5186,N_4271,N_4371);
xor U5187 (N_5187,N_4225,N_4579);
xor U5188 (N_5188,N_4232,N_4233);
and U5189 (N_5189,N_4625,N_4382);
nor U5190 (N_5190,N_4713,N_4768);
and U5191 (N_5191,N_4423,N_4511);
nor U5192 (N_5192,N_4617,N_4791);
nand U5193 (N_5193,N_4768,N_4769);
nand U5194 (N_5194,N_4422,N_4572);
nor U5195 (N_5195,N_4624,N_4564);
nand U5196 (N_5196,N_4220,N_4654);
or U5197 (N_5197,N_4336,N_4325);
nand U5198 (N_5198,N_4528,N_4751);
xnor U5199 (N_5199,N_4381,N_4264);
or U5200 (N_5200,N_4512,N_4763);
and U5201 (N_5201,N_4780,N_4676);
nor U5202 (N_5202,N_4415,N_4335);
xnor U5203 (N_5203,N_4367,N_4717);
or U5204 (N_5204,N_4547,N_4385);
and U5205 (N_5205,N_4236,N_4281);
xor U5206 (N_5206,N_4472,N_4540);
xnor U5207 (N_5207,N_4394,N_4523);
or U5208 (N_5208,N_4201,N_4542);
or U5209 (N_5209,N_4322,N_4674);
and U5210 (N_5210,N_4555,N_4306);
or U5211 (N_5211,N_4746,N_4491);
and U5212 (N_5212,N_4629,N_4529);
xnor U5213 (N_5213,N_4379,N_4254);
nand U5214 (N_5214,N_4386,N_4486);
nand U5215 (N_5215,N_4545,N_4676);
or U5216 (N_5216,N_4403,N_4591);
nor U5217 (N_5217,N_4334,N_4391);
and U5218 (N_5218,N_4297,N_4594);
nand U5219 (N_5219,N_4387,N_4277);
or U5220 (N_5220,N_4715,N_4471);
and U5221 (N_5221,N_4574,N_4393);
and U5222 (N_5222,N_4290,N_4569);
nand U5223 (N_5223,N_4696,N_4378);
nand U5224 (N_5224,N_4384,N_4708);
and U5225 (N_5225,N_4679,N_4516);
nand U5226 (N_5226,N_4799,N_4782);
xnor U5227 (N_5227,N_4423,N_4636);
nor U5228 (N_5228,N_4236,N_4531);
or U5229 (N_5229,N_4444,N_4732);
xnor U5230 (N_5230,N_4386,N_4414);
and U5231 (N_5231,N_4639,N_4376);
and U5232 (N_5232,N_4325,N_4439);
xnor U5233 (N_5233,N_4414,N_4631);
xnor U5234 (N_5234,N_4541,N_4370);
nor U5235 (N_5235,N_4220,N_4555);
and U5236 (N_5236,N_4213,N_4440);
nor U5237 (N_5237,N_4446,N_4533);
nand U5238 (N_5238,N_4362,N_4434);
and U5239 (N_5239,N_4287,N_4700);
xor U5240 (N_5240,N_4226,N_4672);
or U5241 (N_5241,N_4323,N_4486);
and U5242 (N_5242,N_4419,N_4382);
nand U5243 (N_5243,N_4581,N_4327);
xor U5244 (N_5244,N_4437,N_4300);
xnor U5245 (N_5245,N_4434,N_4329);
nor U5246 (N_5246,N_4651,N_4540);
xor U5247 (N_5247,N_4718,N_4453);
or U5248 (N_5248,N_4363,N_4249);
nand U5249 (N_5249,N_4451,N_4670);
nor U5250 (N_5250,N_4641,N_4627);
nor U5251 (N_5251,N_4314,N_4264);
or U5252 (N_5252,N_4715,N_4356);
nand U5253 (N_5253,N_4378,N_4357);
or U5254 (N_5254,N_4224,N_4406);
and U5255 (N_5255,N_4473,N_4781);
or U5256 (N_5256,N_4722,N_4611);
or U5257 (N_5257,N_4689,N_4531);
nor U5258 (N_5258,N_4704,N_4532);
and U5259 (N_5259,N_4349,N_4421);
nor U5260 (N_5260,N_4219,N_4780);
xnor U5261 (N_5261,N_4242,N_4655);
xnor U5262 (N_5262,N_4641,N_4657);
nor U5263 (N_5263,N_4726,N_4625);
nand U5264 (N_5264,N_4400,N_4693);
or U5265 (N_5265,N_4332,N_4486);
xnor U5266 (N_5266,N_4565,N_4347);
nor U5267 (N_5267,N_4586,N_4497);
nand U5268 (N_5268,N_4470,N_4300);
xor U5269 (N_5269,N_4651,N_4306);
or U5270 (N_5270,N_4770,N_4533);
nor U5271 (N_5271,N_4744,N_4596);
and U5272 (N_5272,N_4703,N_4254);
or U5273 (N_5273,N_4625,N_4580);
xor U5274 (N_5274,N_4546,N_4218);
nor U5275 (N_5275,N_4281,N_4489);
nand U5276 (N_5276,N_4607,N_4782);
xnor U5277 (N_5277,N_4561,N_4754);
xor U5278 (N_5278,N_4454,N_4528);
nand U5279 (N_5279,N_4273,N_4494);
nor U5280 (N_5280,N_4434,N_4560);
and U5281 (N_5281,N_4333,N_4211);
xor U5282 (N_5282,N_4287,N_4796);
and U5283 (N_5283,N_4423,N_4435);
or U5284 (N_5284,N_4488,N_4215);
nor U5285 (N_5285,N_4200,N_4705);
and U5286 (N_5286,N_4647,N_4744);
or U5287 (N_5287,N_4440,N_4353);
nor U5288 (N_5288,N_4582,N_4237);
nor U5289 (N_5289,N_4509,N_4758);
xnor U5290 (N_5290,N_4657,N_4690);
or U5291 (N_5291,N_4635,N_4336);
xnor U5292 (N_5292,N_4525,N_4429);
or U5293 (N_5293,N_4369,N_4212);
nand U5294 (N_5294,N_4280,N_4430);
or U5295 (N_5295,N_4631,N_4415);
xor U5296 (N_5296,N_4476,N_4727);
nor U5297 (N_5297,N_4473,N_4389);
xor U5298 (N_5298,N_4607,N_4747);
and U5299 (N_5299,N_4456,N_4217);
or U5300 (N_5300,N_4204,N_4712);
nor U5301 (N_5301,N_4429,N_4292);
nand U5302 (N_5302,N_4615,N_4439);
xor U5303 (N_5303,N_4265,N_4736);
and U5304 (N_5304,N_4330,N_4210);
nand U5305 (N_5305,N_4413,N_4234);
nand U5306 (N_5306,N_4513,N_4567);
xnor U5307 (N_5307,N_4449,N_4650);
or U5308 (N_5308,N_4322,N_4581);
xnor U5309 (N_5309,N_4792,N_4682);
xor U5310 (N_5310,N_4789,N_4338);
and U5311 (N_5311,N_4282,N_4207);
nand U5312 (N_5312,N_4525,N_4780);
or U5313 (N_5313,N_4721,N_4712);
and U5314 (N_5314,N_4532,N_4402);
xor U5315 (N_5315,N_4752,N_4323);
nor U5316 (N_5316,N_4553,N_4676);
and U5317 (N_5317,N_4642,N_4439);
xor U5318 (N_5318,N_4401,N_4696);
xnor U5319 (N_5319,N_4241,N_4755);
nor U5320 (N_5320,N_4364,N_4788);
nand U5321 (N_5321,N_4751,N_4277);
nand U5322 (N_5322,N_4211,N_4228);
and U5323 (N_5323,N_4676,N_4771);
or U5324 (N_5324,N_4284,N_4540);
nor U5325 (N_5325,N_4449,N_4215);
nor U5326 (N_5326,N_4605,N_4727);
nand U5327 (N_5327,N_4201,N_4341);
nand U5328 (N_5328,N_4337,N_4610);
or U5329 (N_5329,N_4711,N_4319);
or U5330 (N_5330,N_4292,N_4530);
nand U5331 (N_5331,N_4775,N_4699);
nor U5332 (N_5332,N_4342,N_4748);
nor U5333 (N_5333,N_4418,N_4384);
or U5334 (N_5334,N_4366,N_4680);
or U5335 (N_5335,N_4768,N_4636);
and U5336 (N_5336,N_4308,N_4474);
nor U5337 (N_5337,N_4528,N_4742);
nor U5338 (N_5338,N_4486,N_4465);
and U5339 (N_5339,N_4683,N_4439);
xnor U5340 (N_5340,N_4404,N_4236);
nand U5341 (N_5341,N_4701,N_4259);
xnor U5342 (N_5342,N_4429,N_4205);
and U5343 (N_5343,N_4310,N_4512);
nor U5344 (N_5344,N_4734,N_4591);
or U5345 (N_5345,N_4694,N_4368);
nor U5346 (N_5346,N_4496,N_4432);
or U5347 (N_5347,N_4449,N_4366);
nand U5348 (N_5348,N_4317,N_4351);
or U5349 (N_5349,N_4599,N_4399);
nor U5350 (N_5350,N_4238,N_4308);
xor U5351 (N_5351,N_4431,N_4244);
or U5352 (N_5352,N_4395,N_4302);
xor U5353 (N_5353,N_4576,N_4262);
xnor U5354 (N_5354,N_4388,N_4431);
and U5355 (N_5355,N_4592,N_4605);
and U5356 (N_5356,N_4307,N_4434);
or U5357 (N_5357,N_4281,N_4425);
xnor U5358 (N_5358,N_4218,N_4689);
or U5359 (N_5359,N_4305,N_4416);
or U5360 (N_5360,N_4274,N_4388);
xor U5361 (N_5361,N_4696,N_4338);
xor U5362 (N_5362,N_4396,N_4524);
and U5363 (N_5363,N_4524,N_4230);
xor U5364 (N_5364,N_4253,N_4441);
xor U5365 (N_5365,N_4494,N_4459);
nor U5366 (N_5366,N_4403,N_4251);
or U5367 (N_5367,N_4646,N_4623);
and U5368 (N_5368,N_4402,N_4386);
xnor U5369 (N_5369,N_4243,N_4322);
and U5370 (N_5370,N_4417,N_4384);
nand U5371 (N_5371,N_4476,N_4794);
or U5372 (N_5372,N_4282,N_4333);
or U5373 (N_5373,N_4403,N_4280);
or U5374 (N_5374,N_4469,N_4585);
or U5375 (N_5375,N_4698,N_4319);
or U5376 (N_5376,N_4432,N_4654);
nand U5377 (N_5377,N_4373,N_4702);
nand U5378 (N_5378,N_4231,N_4409);
or U5379 (N_5379,N_4358,N_4303);
nor U5380 (N_5380,N_4451,N_4216);
or U5381 (N_5381,N_4729,N_4347);
and U5382 (N_5382,N_4279,N_4578);
nor U5383 (N_5383,N_4698,N_4324);
nand U5384 (N_5384,N_4776,N_4793);
nor U5385 (N_5385,N_4212,N_4662);
or U5386 (N_5386,N_4363,N_4621);
and U5387 (N_5387,N_4724,N_4659);
nand U5388 (N_5388,N_4614,N_4411);
or U5389 (N_5389,N_4475,N_4457);
and U5390 (N_5390,N_4566,N_4438);
xor U5391 (N_5391,N_4479,N_4413);
nor U5392 (N_5392,N_4599,N_4593);
nor U5393 (N_5393,N_4311,N_4246);
xor U5394 (N_5394,N_4306,N_4364);
nor U5395 (N_5395,N_4600,N_4623);
and U5396 (N_5396,N_4601,N_4737);
xor U5397 (N_5397,N_4288,N_4519);
nand U5398 (N_5398,N_4673,N_4522);
nor U5399 (N_5399,N_4606,N_4664);
and U5400 (N_5400,N_5397,N_5283);
nand U5401 (N_5401,N_5256,N_4914);
and U5402 (N_5402,N_4851,N_4963);
and U5403 (N_5403,N_4975,N_5238);
xor U5404 (N_5404,N_4823,N_4961);
xnor U5405 (N_5405,N_5157,N_5240);
xnor U5406 (N_5406,N_5188,N_5323);
nor U5407 (N_5407,N_5230,N_4840);
nor U5408 (N_5408,N_5395,N_5115);
nand U5409 (N_5409,N_5264,N_5312);
xnor U5410 (N_5410,N_4866,N_4938);
and U5411 (N_5411,N_5385,N_5314);
and U5412 (N_5412,N_5338,N_5216);
or U5413 (N_5413,N_5033,N_4803);
nor U5414 (N_5414,N_5164,N_4815);
or U5415 (N_5415,N_5378,N_5326);
nor U5416 (N_5416,N_4971,N_5398);
xor U5417 (N_5417,N_5151,N_4877);
nor U5418 (N_5418,N_5104,N_5041);
or U5419 (N_5419,N_5122,N_5340);
nand U5420 (N_5420,N_5137,N_5106);
nor U5421 (N_5421,N_4974,N_5308);
and U5422 (N_5422,N_4891,N_5381);
and U5423 (N_5423,N_5224,N_5059);
nor U5424 (N_5424,N_4928,N_5310);
and U5425 (N_5425,N_4944,N_4842);
and U5426 (N_5426,N_5274,N_4824);
nor U5427 (N_5427,N_5003,N_5026);
nor U5428 (N_5428,N_5217,N_4935);
nor U5429 (N_5429,N_5210,N_5013);
and U5430 (N_5430,N_4850,N_4822);
and U5431 (N_5431,N_5253,N_5111);
or U5432 (N_5432,N_5054,N_4896);
xnor U5433 (N_5433,N_5155,N_5218);
nor U5434 (N_5434,N_5249,N_4899);
nand U5435 (N_5435,N_5040,N_4876);
or U5436 (N_5436,N_5108,N_4986);
xnor U5437 (N_5437,N_5291,N_4806);
and U5438 (N_5438,N_5025,N_5069);
nand U5439 (N_5439,N_5051,N_5192);
nor U5440 (N_5440,N_4884,N_5229);
or U5441 (N_5441,N_5296,N_5076);
nand U5442 (N_5442,N_5214,N_4981);
nand U5443 (N_5443,N_4933,N_5209);
nand U5444 (N_5444,N_5363,N_5067);
or U5445 (N_5445,N_5023,N_5097);
nand U5446 (N_5446,N_5128,N_4959);
and U5447 (N_5447,N_4925,N_4998);
nor U5448 (N_5448,N_4911,N_5208);
nor U5449 (N_5449,N_5081,N_5182);
nand U5450 (N_5450,N_5130,N_5147);
nand U5451 (N_5451,N_5101,N_4912);
and U5452 (N_5452,N_5096,N_5358);
and U5453 (N_5453,N_5311,N_5317);
nor U5454 (N_5454,N_5005,N_5204);
or U5455 (N_5455,N_5201,N_5021);
and U5456 (N_5456,N_4859,N_5272);
xor U5457 (N_5457,N_4839,N_5258);
nor U5458 (N_5458,N_4955,N_4980);
and U5459 (N_5459,N_5043,N_5347);
or U5460 (N_5460,N_5337,N_5309);
nand U5461 (N_5461,N_4906,N_5391);
and U5462 (N_5462,N_5191,N_5367);
xnor U5463 (N_5463,N_5083,N_4816);
and U5464 (N_5464,N_5279,N_4894);
nor U5465 (N_5465,N_5116,N_5286);
nand U5466 (N_5466,N_5292,N_4807);
or U5467 (N_5467,N_5047,N_5284);
nor U5468 (N_5468,N_5354,N_5222);
xnor U5469 (N_5469,N_4885,N_4875);
or U5470 (N_5470,N_5046,N_5380);
nand U5471 (N_5471,N_5223,N_5185);
and U5472 (N_5472,N_4953,N_4869);
nor U5473 (N_5473,N_4872,N_5012);
xnor U5474 (N_5474,N_5149,N_4878);
and U5475 (N_5475,N_4956,N_5074);
and U5476 (N_5476,N_5095,N_5319);
or U5477 (N_5477,N_5144,N_4874);
or U5478 (N_5478,N_5320,N_5241);
nand U5479 (N_5479,N_5390,N_5060);
nor U5480 (N_5480,N_4804,N_5017);
or U5481 (N_5481,N_5287,N_5334);
nor U5482 (N_5482,N_5177,N_5031);
nor U5483 (N_5483,N_5163,N_5330);
nor U5484 (N_5484,N_4942,N_5190);
xor U5485 (N_5485,N_5350,N_5120);
or U5486 (N_5486,N_4965,N_5316);
xnor U5487 (N_5487,N_5091,N_4819);
nand U5488 (N_5488,N_4836,N_5006);
nand U5489 (N_5489,N_4898,N_4856);
xor U5490 (N_5490,N_4987,N_5393);
xnor U5491 (N_5491,N_5133,N_4920);
nor U5492 (N_5492,N_5198,N_4949);
xnor U5493 (N_5493,N_5343,N_5353);
and U5494 (N_5494,N_5269,N_4993);
nand U5495 (N_5495,N_5299,N_5225);
xor U5496 (N_5496,N_4957,N_5084);
and U5497 (N_5497,N_5268,N_5065);
and U5498 (N_5498,N_5288,N_4926);
nor U5499 (N_5499,N_5129,N_4910);
nor U5500 (N_5500,N_4948,N_4905);
or U5501 (N_5501,N_5034,N_4946);
and U5502 (N_5502,N_5359,N_4958);
xnor U5503 (N_5503,N_5261,N_4814);
and U5504 (N_5504,N_4923,N_5127);
and U5505 (N_5505,N_5200,N_4863);
nor U5506 (N_5506,N_4999,N_5145);
or U5507 (N_5507,N_5165,N_5121);
or U5508 (N_5508,N_5117,N_5019);
and U5509 (N_5509,N_4817,N_5082);
nand U5510 (N_5510,N_5114,N_5064);
nand U5511 (N_5511,N_5068,N_5180);
nor U5512 (N_5512,N_5248,N_5161);
nand U5513 (N_5513,N_5220,N_5212);
and U5514 (N_5514,N_5061,N_5105);
and U5515 (N_5515,N_4805,N_5260);
nand U5516 (N_5516,N_5125,N_4812);
and U5517 (N_5517,N_5360,N_5331);
nand U5518 (N_5518,N_4883,N_4900);
or U5519 (N_5519,N_4827,N_5370);
nor U5520 (N_5520,N_5294,N_5044);
or U5521 (N_5521,N_4849,N_5307);
or U5522 (N_5522,N_5318,N_5004);
nor U5523 (N_5523,N_5183,N_5276);
or U5524 (N_5524,N_5138,N_5369);
and U5525 (N_5525,N_5265,N_4967);
nor U5526 (N_5526,N_4855,N_4882);
and U5527 (N_5527,N_5078,N_5071);
and U5528 (N_5528,N_5001,N_5364);
and U5529 (N_5529,N_5328,N_5139);
xnor U5530 (N_5530,N_4813,N_4844);
nand U5531 (N_5531,N_5346,N_5199);
xor U5532 (N_5532,N_5196,N_5304);
nor U5533 (N_5533,N_4909,N_5245);
nand U5534 (N_5534,N_5302,N_5169);
xnor U5535 (N_5535,N_5152,N_5072);
nor U5536 (N_5536,N_5186,N_5285);
xnor U5537 (N_5537,N_5366,N_5235);
xor U5538 (N_5538,N_5202,N_4830);
and U5539 (N_5539,N_5184,N_4831);
or U5540 (N_5540,N_4893,N_5211);
nand U5541 (N_5541,N_5301,N_5087);
and U5542 (N_5542,N_5227,N_5056);
xnor U5543 (N_5543,N_4892,N_4964);
nand U5544 (N_5544,N_4835,N_4908);
nor U5545 (N_5545,N_5039,N_5322);
nand U5546 (N_5546,N_5016,N_4801);
and U5547 (N_5547,N_4983,N_5313);
nor U5548 (N_5548,N_4862,N_5252);
xor U5549 (N_5549,N_5049,N_5244);
nor U5550 (N_5550,N_4913,N_5389);
and U5551 (N_5551,N_4989,N_5329);
xor U5552 (N_5552,N_5228,N_5085);
nand U5553 (N_5553,N_4922,N_5058);
nand U5554 (N_5554,N_5374,N_5305);
xnor U5555 (N_5555,N_5112,N_4848);
or U5556 (N_5556,N_5386,N_5148);
nand U5557 (N_5557,N_5221,N_5153);
or U5558 (N_5558,N_5070,N_5159);
nand U5559 (N_5559,N_5266,N_5052);
nor U5560 (N_5560,N_5189,N_5270);
nand U5561 (N_5561,N_5242,N_5042);
nor U5562 (N_5562,N_4834,N_5348);
nor U5563 (N_5563,N_5048,N_5349);
nor U5564 (N_5564,N_5140,N_4943);
nand U5565 (N_5565,N_4837,N_5156);
xnor U5566 (N_5566,N_5394,N_5088);
and U5567 (N_5567,N_5193,N_4995);
xnor U5568 (N_5568,N_5336,N_5321);
and U5569 (N_5569,N_5123,N_5361);
xor U5570 (N_5570,N_5045,N_4847);
xor U5571 (N_5571,N_5035,N_4952);
and U5572 (N_5572,N_4843,N_4857);
nor U5573 (N_5573,N_5022,N_5073);
xnor U5574 (N_5574,N_5267,N_5344);
xor U5575 (N_5575,N_5110,N_5194);
and U5576 (N_5576,N_5057,N_5126);
or U5577 (N_5577,N_5357,N_4841);
nand U5578 (N_5578,N_5089,N_5351);
nand U5579 (N_5579,N_5100,N_4968);
and U5580 (N_5580,N_5327,N_5018);
nor U5581 (N_5581,N_5113,N_5333);
xor U5582 (N_5582,N_4941,N_5086);
or U5583 (N_5583,N_5280,N_5203);
and U5584 (N_5584,N_4915,N_5055);
and U5585 (N_5585,N_5154,N_4939);
xnor U5586 (N_5586,N_5399,N_5251);
xor U5587 (N_5587,N_5124,N_5118);
xor U5588 (N_5588,N_5011,N_5195);
xnor U5589 (N_5589,N_5226,N_5102);
xnor U5590 (N_5590,N_4954,N_5368);
or U5591 (N_5591,N_5372,N_5332);
or U5592 (N_5592,N_5298,N_4861);
nor U5593 (N_5593,N_4916,N_5080);
or U5594 (N_5594,N_4996,N_5092);
nand U5595 (N_5595,N_5170,N_5342);
or U5596 (N_5596,N_5315,N_4972);
or U5597 (N_5597,N_4997,N_5219);
nor U5598 (N_5598,N_5277,N_4890);
nand U5599 (N_5599,N_5303,N_5243);
xor U5600 (N_5600,N_4810,N_5231);
or U5601 (N_5601,N_5234,N_5027);
nand U5602 (N_5602,N_4991,N_5098);
and U5603 (N_5603,N_5030,N_4846);
nand U5604 (N_5604,N_5236,N_4870);
and U5605 (N_5605,N_5099,N_4930);
nor U5606 (N_5606,N_4918,N_4802);
xnor U5607 (N_5607,N_5373,N_5206);
nor U5608 (N_5608,N_4969,N_5167);
and U5609 (N_5609,N_4931,N_4904);
or U5610 (N_5610,N_5352,N_5050);
xnor U5611 (N_5611,N_4828,N_5014);
or U5612 (N_5612,N_5171,N_5246);
xor U5613 (N_5613,N_4858,N_4808);
nand U5614 (N_5614,N_5355,N_5362);
nor U5615 (N_5615,N_4825,N_5392);
nor U5616 (N_5616,N_4826,N_4902);
and U5617 (N_5617,N_5281,N_5396);
or U5618 (N_5618,N_4907,N_5207);
nand U5619 (N_5619,N_5384,N_4984);
nand U5620 (N_5620,N_4994,N_5379);
or U5621 (N_5621,N_5371,N_5375);
xnor U5622 (N_5622,N_5103,N_5077);
nand U5623 (N_5623,N_5306,N_5365);
or U5624 (N_5624,N_4962,N_4937);
or U5625 (N_5625,N_4881,N_5295);
or U5626 (N_5626,N_5007,N_5213);
nand U5627 (N_5627,N_5008,N_4887);
or U5628 (N_5628,N_5020,N_5377);
nor U5629 (N_5629,N_5166,N_5187);
nor U5630 (N_5630,N_5160,N_4888);
nand U5631 (N_5631,N_5037,N_5024);
nor U5632 (N_5632,N_5002,N_5174);
nand U5633 (N_5633,N_5109,N_4927);
nand U5634 (N_5634,N_5290,N_5289);
nand U5635 (N_5635,N_5255,N_4979);
xnor U5636 (N_5636,N_4845,N_5131);
nand U5637 (N_5637,N_5247,N_5143);
or U5638 (N_5638,N_4929,N_4990);
nand U5639 (N_5639,N_4970,N_4889);
nor U5640 (N_5640,N_5000,N_5339);
nand U5641 (N_5641,N_4879,N_5173);
nor U5642 (N_5642,N_4940,N_5036);
xnor U5643 (N_5643,N_4978,N_5356);
and U5644 (N_5644,N_4934,N_4901);
nor U5645 (N_5645,N_5293,N_5066);
and U5646 (N_5646,N_5029,N_5239);
or U5647 (N_5647,N_4820,N_5090);
or U5648 (N_5648,N_5172,N_5383);
xor U5649 (N_5649,N_5038,N_4977);
and U5650 (N_5650,N_5134,N_5032);
xor U5651 (N_5651,N_5009,N_4895);
or U5652 (N_5652,N_5162,N_5262);
nand U5653 (N_5653,N_4982,N_5345);
and U5654 (N_5654,N_5063,N_5028);
nor U5655 (N_5655,N_4903,N_4821);
nand U5656 (N_5656,N_5175,N_4829);
or U5657 (N_5657,N_4880,N_4973);
or U5658 (N_5658,N_5250,N_4854);
nor U5659 (N_5659,N_4852,N_5179);
or U5660 (N_5660,N_5136,N_4868);
xnor U5661 (N_5661,N_5168,N_5335);
xnor U5662 (N_5662,N_4811,N_4921);
and U5663 (N_5663,N_4924,N_5094);
nor U5664 (N_5664,N_5237,N_4919);
nand U5665 (N_5665,N_5278,N_5275);
nor U5666 (N_5666,N_5178,N_4932);
and U5667 (N_5667,N_5387,N_5300);
and U5668 (N_5668,N_5146,N_5382);
nand U5669 (N_5669,N_5135,N_5197);
and U5670 (N_5670,N_4897,N_4966);
nor U5671 (N_5671,N_4867,N_4985);
xor U5672 (N_5672,N_5150,N_4950);
and U5673 (N_5673,N_5325,N_5254);
or U5674 (N_5674,N_4988,N_4864);
nor U5675 (N_5675,N_4800,N_5341);
and U5676 (N_5676,N_5257,N_5324);
xor U5677 (N_5677,N_5233,N_5158);
or U5678 (N_5678,N_5093,N_4947);
or U5679 (N_5679,N_5053,N_5132);
nand U5680 (N_5680,N_4886,N_5107);
nor U5681 (N_5681,N_5388,N_4832);
nor U5682 (N_5682,N_4838,N_5215);
nand U5683 (N_5683,N_4860,N_5075);
and U5684 (N_5684,N_5232,N_4992);
or U5685 (N_5685,N_5271,N_4871);
and U5686 (N_5686,N_5141,N_5079);
nor U5687 (N_5687,N_4865,N_5142);
and U5688 (N_5688,N_5273,N_4853);
nand U5689 (N_5689,N_5010,N_4833);
xor U5690 (N_5690,N_5119,N_4917);
nor U5691 (N_5691,N_5376,N_5062);
or U5692 (N_5692,N_4945,N_5015);
nor U5693 (N_5693,N_5263,N_5282);
or U5694 (N_5694,N_5297,N_4951);
nor U5695 (N_5695,N_4960,N_5205);
xnor U5696 (N_5696,N_5176,N_5181);
nor U5697 (N_5697,N_4818,N_4976);
nor U5698 (N_5698,N_4873,N_4809);
xnor U5699 (N_5699,N_5259,N_4936);
or U5700 (N_5700,N_5284,N_5281);
and U5701 (N_5701,N_4987,N_4916);
or U5702 (N_5702,N_4944,N_5185);
xnor U5703 (N_5703,N_5329,N_5332);
nor U5704 (N_5704,N_4860,N_5301);
xor U5705 (N_5705,N_5195,N_4895);
nand U5706 (N_5706,N_4826,N_5282);
xor U5707 (N_5707,N_5380,N_5193);
xor U5708 (N_5708,N_4959,N_5197);
and U5709 (N_5709,N_5005,N_5002);
or U5710 (N_5710,N_5099,N_4801);
and U5711 (N_5711,N_4896,N_4988);
or U5712 (N_5712,N_4923,N_4971);
nor U5713 (N_5713,N_4983,N_5159);
or U5714 (N_5714,N_5122,N_5039);
and U5715 (N_5715,N_5245,N_5248);
xor U5716 (N_5716,N_5238,N_5399);
nor U5717 (N_5717,N_5307,N_4914);
and U5718 (N_5718,N_5157,N_5271);
nor U5719 (N_5719,N_4941,N_4858);
nor U5720 (N_5720,N_5019,N_4987);
nor U5721 (N_5721,N_5338,N_5282);
nor U5722 (N_5722,N_5215,N_5062);
nand U5723 (N_5723,N_5339,N_5019);
or U5724 (N_5724,N_5327,N_5164);
xor U5725 (N_5725,N_5140,N_5365);
or U5726 (N_5726,N_5317,N_5186);
xor U5727 (N_5727,N_4981,N_4926);
nor U5728 (N_5728,N_5381,N_5303);
nand U5729 (N_5729,N_4861,N_5399);
nand U5730 (N_5730,N_5379,N_5389);
and U5731 (N_5731,N_5306,N_5057);
nor U5732 (N_5732,N_5144,N_5390);
or U5733 (N_5733,N_5390,N_5066);
or U5734 (N_5734,N_5355,N_4872);
nand U5735 (N_5735,N_5128,N_4912);
xor U5736 (N_5736,N_5166,N_5056);
or U5737 (N_5737,N_5159,N_5057);
and U5738 (N_5738,N_5215,N_5325);
nand U5739 (N_5739,N_4943,N_5160);
nor U5740 (N_5740,N_4886,N_5067);
nor U5741 (N_5741,N_5351,N_4893);
or U5742 (N_5742,N_4920,N_5146);
nand U5743 (N_5743,N_4847,N_4851);
nand U5744 (N_5744,N_5389,N_5090);
xnor U5745 (N_5745,N_4972,N_5325);
nor U5746 (N_5746,N_5281,N_5296);
nor U5747 (N_5747,N_5046,N_5388);
xnor U5748 (N_5748,N_4986,N_5172);
and U5749 (N_5749,N_4926,N_5028);
xor U5750 (N_5750,N_4963,N_4848);
nor U5751 (N_5751,N_4996,N_5312);
or U5752 (N_5752,N_5310,N_4840);
xor U5753 (N_5753,N_4898,N_5111);
xor U5754 (N_5754,N_5364,N_5291);
nor U5755 (N_5755,N_5063,N_5223);
nor U5756 (N_5756,N_5292,N_5214);
xnor U5757 (N_5757,N_5035,N_5276);
nor U5758 (N_5758,N_4834,N_4953);
or U5759 (N_5759,N_4963,N_5039);
nor U5760 (N_5760,N_4813,N_5141);
nand U5761 (N_5761,N_4836,N_5360);
nor U5762 (N_5762,N_5214,N_5124);
or U5763 (N_5763,N_4815,N_5063);
or U5764 (N_5764,N_4901,N_4912);
nand U5765 (N_5765,N_5353,N_5208);
xnor U5766 (N_5766,N_4962,N_5218);
nor U5767 (N_5767,N_5288,N_4952);
nand U5768 (N_5768,N_5266,N_5065);
nand U5769 (N_5769,N_5120,N_5119);
xor U5770 (N_5770,N_4996,N_4870);
nand U5771 (N_5771,N_5283,N_5371);
xnor U5772 (N_5772,N_5144,N_5161);
xnor U5773 (N_5773,N_5096,N_4901);
xor U5774 (N_5774,N_4990,N_5105);
xnor U5775 (N_5775,N_4983,N_5353);
and U5776 (N_5776,N_4870,N_5058);
or U5777 (N_5777,N_5230,N_5306);
xor U5778 (N_5778,N_5158,N_4972);
or U5779 (N_5779,N_5192,N_5304);
nor U5780 (N_5780,N_5065,N_5244);
nand U5781 (N_5781,N_5203,N_5309);
or U5782 (N_5782,N_5262,N_4984);
or U5783 (N_5783,N_5005,N_4837);
xor U5784 (N_5784,N_5025,N_5175);
xnor U5785 (N_5785,N_5063,N_5195);
nor U5786 (N_5786,N_4849,N_4976);
and U5787 (N_5787,N_5359,N_5157);
or U5788 (N_5788,N_4800,N_4879);
nand U5789 (N_5789,N_5145,N_5363);
xnor U5790 (N_5790,N_5240,N_5396);
or U5791 (N_5791,N_4854,N_4821);
and U5792 (N_5792,N_4858,N_4804);
and U5793 (N_5793,N_5008,N_5160);
xnor U5794 (N_5794,N_5398,N_4854);
xnor U5795 (N_5795,N_4845,N_5162);
nand U5796 (N_5796,N_4871,N_5192);
nand U5797 (N_5797,N_5373,N_4920);
and U5798 (N_5798,N_4912,N_4824);
and U5799 (N_5799,N_4991,N_5012);
xor U5800 (N_5800,N_4857,N_5364);
xnor U5801 (N_5801,N_4908,N_4981);
nand U5802 (N_5802,N_5316,N_5092);
nand U5803 (N_5803,N_5081,N_5388);
xnor U5804 (N_5804,N_4908,N_5245);
and U5805 (N_5805,N_5179,N_4989);
nand U5806 (N_5806,N_4834,N_5184);
nor U5807 (N_5807,N_4881,N_5366);
or U5808 (N_5808,N_5211,N_5084);
or U5809 (N_5809,N_4980,N_5134);
xnor U5810 (N_5810,N_5367,N_5371);
nand U5811 (N_5811,N_5296,N_5316);
or U5812 (N_5812,N_4834,N_5222);
and U5813 (N_5813,N_4878,N_4960);
and U5814 (N_5814,N_4861,N_4919);
xnor U5815 (N_5815,N_5104,N_5380);
and U5816 (N_5816,N_5374,N_4806);
and U5817 (N_5817,N_5301,N_5256);
or U5818 (N_5818,N_4943,N_5392);
and U5819 (N_5819,N_4963,N_4817);
or U5820 (N_5820,N_4850,N_4919);
nor U5821 (N_5821,N_4966,N_5146);
or U5822 (N_5822,N_4872,N_5236);
and U5823 (N_5823,N_4826,N_4814);
nand U5824 (N_5824,N_4962,N_5244);
xor U5825 (N_5825,N_5298,N_5024);
xor U5826 (N_5826,N_5168,N_5344);
or U5827 (N_5827,N_5353,N_5001);
xor U5828 (N_5828,N_4986,N_5192);
xnor U5829 (N_5829,N_4930,N_4918);
and U5830 (N_5830,N_5392,N_4829);
xnor U5831 (N_5831,N_5254,N_5290);
xnor U5832 (N_5832,N_4966,N_5170);
nand U5833 (N_5833,N_5134,N_5181);
or U5834 (N_5834,N_5033,N_4901);
xor U5835 (N_5835,N_4891,N_5211);
nor U5836 (N_5836,N_5206,N_5389);
nor U5837 (N_5837,N_4860,N_5310);
xor U5838 (N_5838,N_4945,N_5233);
nor U5839 (N_5839,N_5291,N_5084);
nor U5840 (N_5840,N_4800,N_5023);
or U5841 (N_5841,N_4851,N_4864);
nand U5842 (N_5842,N_5284,N_5333);
nand U5843 (N_5843,N_5055,N_5309);
nor U5844 (N_5844,N_4872,N_5352);
or U5845 (N_5845,N_4852,N_4919);
and U5846 (N_5846,N_5152,N_5268);
or U5847 (N_5847,N_4952,N_5387);
xor U5848 (N_5848,N_5092,N_4914);
nand U5849 (N_5849,N_5074,N_4895);
nor U5850 (N_5850,N_5032,N_5347);
and U5851 (N_5851,N_5195,N_5169);
nand U5852 (N_5852,N_4987,N_4993);
nand U5853 (N_5853,N_5019,N_5113);
and U5854 (N_5854,N_5246,N_5158);
and U5855 (N_5855,N_5000,N_4869);
nor U5856 (N_5856,N_5011,N_4901);
nor U5857 (N_5857,N_5330,N_5303);
nor U5858 (N_5858,N_5236,N_5260);
and U5859 (N_5859,N_5034,N_4926);
nor U5860 (N_5860,N_5041,N_5105);
and U5861 (N_5861,N_5177,N_5011);
xnor U5862 (N_5862,N_4925,N_4959);
or U5863 (N_5863,N_4992,N_5014);
and U5864 (N_5864,N_5232,N_4960);
nor U5865 (N_5865,N_4928,N_5222);
nor U5866 (N_5866,N_5278,N_5197);
and U5867 (N_5867,N_4960,N_5000);
or U5868 (N_5868,N_5072,N_5130);
nand U5869 (N_5869,N_5170,N_4833);
and U5870 (N_5870,N_4835,N_5289);
nor U5871 (N_5871,N_5262,N_5391);
nor U5872 (N_5872,N_4848,N_4883);
nor U5873 (N_5873,N_5216,N_5247);
or U5874 (N_5874,N_5165,N_5088);
xor U5875 (N_5875,N_4918,N_4973);
nand U5876 (N_5876,N_5091,N_5074);
and U5877 (N_5877,N_4847,N_5329);
xor U5878 (N_5878,N_4949,N_5265);
nand U5879 (N_5879,N_5211,N_4868);
and U5880 (N_5880,N_4866,N_5236);
xnor U5881 (N_5881,N_5362,N_5344);
nor U5882 (N_5882,N_5199,N_5045);
xnor U5883 (N_5883,N_4892,N_5175);
and U5884 (N_5884,N_4971,N_5393);
or U5885 (N_5885,N_4920,N_5256);
nand U5886 (N_5886,N_4862,N_4887);
xor U5887 (N_5887,N_4907,N_5246);
nand U5888 (N_5888,N_5114,N_4829);
or U5889 (N_5889,N_4917,N_5276);
nor U5890 (N_5890,N_4929,N_5264);
xnor U5891 (N_5891,N_5276,N_5389);
nand U5892 (N_5892,N_4876,N_5054);
and U5893 (N_5893,N_5052,N_5011);
nor U5894 (N_5894,N_5079,N_5137);
and U5895 (N_5895,N_5176,N_5239);
or U5896 (N_5896,N_5241,N_4979);
and U5897 (N_5897,N_4953,N_4924);
or U5898 (N_5898,N_5084,N_5041);
xor U5899 (N_5899,N_5029,N_5317);
nor U5900 (N_5900,N_4908,N_4887);
xnor U5901 (N_5901,N_5358,N_5074);
or U5902 (N_5902,N_5380,N_5269);
nor U5903 (N_5903,N_5067,N_5175);
nand U5904 (N_5904,N_4862,N_5232);
xnor U5905 (N_5905,N_5370,N_5063);
nand U5906 (N_5906,N_4836,N_4978);
nand U5907 (N_5907,N_4952,N_5355);
or U5908 (N_5908,N_5227,N_5073);
nor U5909 (N_5909,N_4967,N_5339);
xor U5910 (N_5910,N_5369,N_5310);
xor U5911 (N_5911,N_4849,N_5164);
xor U5912 (N_5912,N_5107,N_4894);
nor U5913 (N_5913,N_5180,N_4984);
and U5914 (N_5914,N_5310,N_5028);
nor U5915 (N_5915,N_5213,N_5155);
nor U5916 (N_5916,N_5301,N_4800);
nand U5917 (N_5917,N_4920,N_4806);
xor U5918 (N_5918,N_4926,N_5012);
and U5919 (N_5919,N_5361,N_5204);
or U5920 (N_5920,N_4883,N_4919);
nand U5921 (N_5921,N_4854,N_4866);
and U5922 (N_5922,N_4924,N_5228);
xnor U5923 (N_5923,N_4949,N_4922);
and U5924 (N_5924,N_5265,N_5381);
xnor U5925 (N_5925,N_5193,N_5366);
and U5926 (N_5926,N_5137,N_5152);
and U5927 (N_5927,N_5238,N_5310);
nor U5928 (N_5928,N_4847,N_5068);
nand U5929 (N_5929,N_4959,N_4905);
and U5930 (N_5930,N_4986,N_5297);
nand U5931 (N_5931,N_5344,N_5185);
nor U5932 (N_5932,N_4916,N_5011);
or U5933 (N_5933,N_5190,N_4881);
and U5934 (N_5934,N_5317,N_4865);
xor U5935 (N_5935,N_5318,N_5131);
nand U5936 (N_5936,N_5301,N_5214);
or U5937 (N_5937,N_5285,N_5176);
or U5938 (N_5938,N_5325,N_5241);
and U5939 (N_5939,N_4903,N_5261);
xor U5940 (N_5940,N_4990,N_5210);
and U5941 (N_5941,N_5358,N_4990);
nor U5942 (N_5942,N_5124,N_4912);
or U5943 (N_5943,N_5321,N_5295);
nor U5944 (N_5944,N_5071,N_4949);
nand U5945 (N_5945,N_4909,N_5011);
nand U5946 (N_5946,N_5371,N_5184);
and U5947 (N_5947,N_5282,N_4810);
and U5948 (N_5948,N_5230,N_5369);
nor U5949 (N_5949,N_5105,N_5216);
and U5950 (N_5950,N_5076,N_5172);
nand U5951 (N_5951,N_5299,N_4977);
and U5952 (N_5952,N_5365,N_5127);
and U5953 (N_5953,N_4999,N_5187);
and U5954 (N_5954,N_4934,N_4933);
nor U5955 (N_5955,N_5020,N_5364);
nor U5956 (N_5956,N_5396,N_5200);
and U5957 (N_5957,N_5175,N_4875);
nor U5958 (N_5958,N_5231,N_4979);
or U5959 (N_5959,N_4917,N_5198);
or U5960 (N_5960,N_5397,N_5341);
or U5961 (N_5961,N_5379,N_4926);
nor U5962 (N_5962,N_4943,N_4903);
xnor U5963 (N_5963,N_5320,N_4975);
nor U5964 (N_5964,N_5267,N_5308);
xor U5965 (N_5965,N_5289,N_4893);
nand U5966 (N_5966,N_5350,N_5265);
nand U5967 (N_5967,N_4858,N_4933);
or U5968 (N_5968,N_5297,N_5222);
nand U5969 (N_5969,N_4924,N_5046);
xor U5970 (N_5970,N_5162,N_4945);
nor U5971 (N_5971,N_4866,N_4971);
or U5972 (N_5972,N_5225,N_4920);
or U5973 (N_5973,N_5381,N_4914);
nor U5974 (N_5974,N_4995,N_5252);
nor U5975 (N_5975,N_5291,N_5005);
nor U5976 (N_5976,N_5019,N_5043);
xnor U5977 (N_5977,N_4995,N_4924);
nand U5978 (N_5978,N_4882,N_5093);
nor U5979 (N_5979,N_4955,N_4834);
and U5980 (N_5980,N_5346,N_5012);
xor U5981 (N_5981,N_5022,N_4995);
nor U5982 (N_5982,N_4888,N_4952);
nand U5983 (N_5983,N_4823,N_5047);
nand U5984 (N_5984,N_5384,N_5034);
and U5985 (N_5985,N_5049,N_5276);
and U5986 (N_5986,N_4951,N_4849);
nor U5987 (N_5987,N_4895,N_5393);
nor U5988 (N_5988,N_5278,N_5369);
nor U5989 (N_5989,N_5326,N_5046);
xnor U5990 (N_5990,N_4827,N_5181);
nand U5991 (N_5991,N_4865,N_5319);
nor U5992 (N_5992,N_5273,N_5141);
or U5993 (N_5993,N_5177,N_5061);
xor U5994 (N_5994,N_4917,N_4841);
nand U5995 (N_5995,N_5076,N_5357);
or U5996 (N_5996,N_5121,N_5351);
or U5997 (N_5997,N_4871,N_5308);
and U5998 (N_5998,N_5178,N_5326);
or U5999 (N_5999,N_4975,N_5062);
nor U6000 (N_6000,N_5775,N_5727);
nor U6001 (N_6001,N_5876,N_5797);
and U6002 (N_6002,N_5894,N_5459);
and U6003 (N_6003,N_5549,N_5930);
and U6004 (N_6004,N_5823,N_5936);
or U6005 (N_6005,N_5713,N_5481);
nor U6006 (N_6006,N_5550,N_5914);
xor U6007 (N_6007,N_5557,N_5642);
and U6008 (N_6008,N_5430,N_5898);
xnor U6009 (N_6009,N_5856,N_5610);
nand U6010 (N_6010,N_5933,N_5434);
and U6011 (N_6011,N_5998,N_5540);
or U6012 (N_6012,N_5616,N_5491);
and U6013 (N_6013,N_5615,N_5660);
nor U6014 (N_6014,N_5868,N_5818);
nor U6015 (N_6015,N_5408,N_5804);
nand U6016 (N_6016,N_5544,N_5625);
and U6017 (N_6017,N_5563,N_5714);
nor U6018 (N_6018,N_5975,N_5709);
and U6019 (N_6019,N_5631,N_5955);
or U6020 (N_6020,N_5893,N_5529);
nand U6021 (N_6021,N_5826,N_5979);
nor U6022 (N_6022,N_5520,N_5497);
and U6023 (N_6023,N_5514,N_5897);
xor U6024 (N_6024,N_5668,N_5632);
and U6025 (N_6025,N_5724,N_5847);
or U6026 (N_6026,N_5865,N_5451);
nor U6027 (N_6027,N_5947,N_5988);
nor U6028 (N_6028,N_5944,N_5609);
xnor U6029 (N_6029,N_5411,N_5462);
or U6030 (N_6030,N_5417,N_5526);
nand U6031 (N_6031,N_5982,N_5743);
nand U6032 (N_6032,N_5488,N_5728);
and U6033 (N_6033,N_5414,N_5949);
and U6034 (N_6034,N_5519,N_5703);
or U6035 (N_6035,N_5870,N_5644);
or U6036 (N_6036,N_5901,N_5404);
xor U6037 (N_6037,N_5959,N_5424);
nor U6038 (N_6038,N_5731,N_5630);
or U6039 (N_6039,N_5512,N_5957);
xor U6040 (N_6040,N_5696,N_5891);
nor U6041 (N_6041,N_5694,N_5822);
nand U6042 (N_6042,N_5857,N_5538);
nor U6043 (N_6043,N_5581,N_5806);
nand U6044 (N_6044,N_5556,N_5785);
xor U6045 (N_6045,N_5887,N_5968);
xor U6046 (N_6046,N_5686,N_5587);
nor U6047 (N_6047,N_5405,N_5541);
and U6048 (N_6048,N_5889,N_5861);
and U6049 (N_6049,N_5457,N_5720);
nand U6050 (N_6050,N_5839,N_5428);
nand U6051 (N_6051,N_5678,N_5531);
nand U6052 (N_6052,N_5721,N_5612);
and U6053 (N_6053,N_5426,N_5712);
nor U6054 (N_6054,N_5594,N_5987);
xor U6055 (N_6055,N_5869,N_5432);
xor U6056 (N_6056,N_5677,N_5474);
xor U6057 (N_6057,N_5814,N_5588);
nand U6058 (N_6058,N_5567,N_5729);
and U6059 (N_6059,N_5995,N_5535);
nor U6060 (N_6060,N_5811,N_5664);
nand U6061 (N_6061,N_5726,N_5485);
or U6062 (N_6062,N_5855,N_5776);
xnor U6063 (N_6063,N_5722,N_5621);
xnor U6064 (N_6064,N_5412,N_5977);
xnor U6065 (N_6065,N_5504,N_5848);
xnor U6066 (N_6066,N_5659,N_5693);
xor U6067 (N_6067,N_5939,N_5748);
nor U6068 (N_6068,N_5964,N_5971);
xnor U6069 (N_6069,N_5913,N_5884);
nor U6070 (N_6070,N_5812,N_5701);
nor U6071 (N_6071,N_5871,N_5527);
and U6072 (N_6072,N_5699,N_5681);
nand U6073 (N_6073,N_5738,N_5761);
or U6074 (N_6074,N_5445,N_5685);
xor U6075 (N_6075,N_5917,N_5999);
xor U6076 (N_6076,N_5885,N_5986);
nand U6077 (N_6077,N_5436,N_5505);
nand U6078 (N_6078,N_5570,N_5970);
or U6079 (N_6079,N_5888,N_5499);
xor U6080 (N_6080,N_5771,N_5768);
nand U6081 (N_6081,N_5458,N_5990);
nand U6082 (N_6082,N_5569,N_5716);
xnor U6083 (N_6083,N_5607,N_5628);
nand U6084 (N_6084,N_5576,N_5415);
nand U6085 (N_6085,N_5506,N_5786);
or U6086 (N_6086,N_5912,N_5866);
or U6087 (N_6087,N_5633,N_5854);
or U6088 (N_6088,N_5695,N_5765);
or U6089 (N_6089,N_5962,N_5820);
nor U6090 (N_6090,N_5552,N_5928);
nand U6091 (N_6091,N_5915,N_5573);
nor U6092 (N_6092,N_5600,N_5444);
nor U6093 (N_6093,N_5440,N_5403);
and U6094 (N_6094,N_5952,N_5683);
nor U6095 (N_6095,N_5762,N_5788);
xnor U6096 (N_6096,N_5908,N_5793);
nand U6097 (N_6097,N_5770,N_5781);
or U6098 (N_6098,N_5754,N_5568);
or U6099 (N_6099,N_5443,N_5503);
nand U6100 (N_6100,N_5649,N_5844);
nor U6101 (N_6101,N_5425,N_5476);
xor U6102 (N_6102,N_5456,N_5680);
and U6103 (N_6103,N_5983,N_5654);
and U6104 (N_6104,N_5923,N_5718);
or U6105 (N_6105,N_5803,N_5500);
xnor U6106 (N_6106,N_5467,N_5602);
xor U6107 (N_6107,N_5522,N_5437);
nor U6108 (N_6108,N_5449,N_5619);
or U6109 (N_6109,N_5640,N_5493);
nand U6110 (N_6110,N_5438,N_5838);
nor U6111 (N_6111,N_5574,N_5782);
or U6112 (N_6112,N_5816,N_5571);
xor U6113 (N_6113,N_5954,N_5455);
xnor U6114 (N_6114,N_5945,N_5672);
xnor U6115 (N_6115,N_5673,N_5702);
nor U6116 (N_6116,N_5706,N_5966);
and U6117 (N_6117,N_5518,N_5978);
xnor U6118 (N_6118,N_5652,N_5852);
xor U6119 (N_6119,N_5882,N_5583);
nand U6120 (N_6120,N_5691,N_5539);
or U6121 (N_6121,N_5963,N_5523);
or U6122 (N_6122,N_5584,N_5472);
nor U6123 (N_6123,N_5943,N_5779);
nor U6124 (N_6124,N_5647,N_5525);
nor U6125 (N_6125,N_5495,N_5953);
and U6126 (N_6126,N_5745,N_5688);
nand U6127 (N_6127,N_5725,N_5601);
nand U6128 (N_6128,N_5554,N_5605);
nand U6129 (N_6129,N_5471,N_5409);
nand U6130 (N_6130,N_5850,N_5624);
nor U6131 (N_6131,N_5591,N_5623);
or U6132 (N_6132,N_5749,N_5629);
and U6133 (N_6133,N_5760,N_5617);
nor U6134 (N_6134,N_5817,N_5419);
and U6135 (N_6135,N_5662,N_5980);
and U6136 (N_6136,N_5635,N_5807);
xnor U6137 (N_6137,N_5956,N_5646);
nor U6138 (N_6138,N_5704,N_5469);
or U6139 (N_6139,N_5634,N_5763);
or U6140 (N_6140,N_5942,N_5547);
and U6141 (N_6141,N_5972,N_5698);
nor U6142 (N_6142,N_5585,N_5994);
nor U6143 (N_6143,N_5833,N_5902);
and U6144 (N_6144,N_5466,N_5840);
nor U6145 (N_6145,N_5513,N_5796);
nor U6146 (N_6146,N_5932,N_5593);
nand U6147 (N_6147,N_5827,N_5965);
or U6148 (N_6148,N_5739,N_5477);
nand U6149 (N_6149,N_5951,N_5551);
and U6150 (N_6150,N_5730,N_5516);
xor U6151 (N_6151,N_5922,N_5692);
and U6152 (N_6152,N_5684,N_5489);
and U6153 (N_6153,N_5774,N_5639);
nand U6154 (N_6154,N_5663,N_5929);
nor U6155 (N_6155,N_5864,N_5446);
and U6156 (N_6156,N_5809,N_5690);
or U6157 (N_6157,N_5881,N_5498);
nand U6158 (N_6158,N_5508,N_5441);
nand U6159 (N_6159,N_5764,N_5517);
nand U6160 (N_6160,N_5572,N_5845);
nand U6161 (N_6161,N_5883,N_5920);
nor U6162 (N_6162,N_5784,N_5697);
nor U6163 (N_6163,N_5967,N_5973);
and U6164 (N_6164,N_5808,N_5849);
xor U6165 (N_6165,N_5528,N_5736);
nor U6166 (N_6166,N_5789,N_5905);
xor U6167 (N_6167,N_5627,N_5879);
and U6168 (N_6168,N_5530,N_5859);
xor U6169 (N_6169,N_5741,N_5465);
nand U6170 (N_6170,N_5643,N_5565);
and U6171 (N_6171,N_5661,N_5750);
xnor U6172 (N_6172,N_5470,N_5769);
or U6173 (N_6173,N_5658,N_5834);
or U6174 (N_6174,N_5874,N_5431);
nand U6175 (N_6175,N_5911,N_5402);
nor U6176 (N_6176,N_5766,N_5903);
nor U6177 (N_6177,N_5580,N_5447);
nor U6178 (N_6178,N_5596,N_5909);
or U6179 (N_6179,N_5991,N_5984);
nand U6180 (N_6180,N_5524,N_5558);
nand U6181 (N_6181,N_5759,N_5961);
or U6182 (N_6182,N_5960,N_5401);
or U6183 (N_6183,N_5723,N_5710);
and U6184 (N_6184,N_5496,N_5510);
nor U6185 (N_6185,N_5480,N_5910);
xnor U6186 (N_6186,N_5611,N_5618);
or U6187 (N_6187,N_5622,N_5794);
or U6188 (N_6188,N_5439,N_5821);
xnor U6189 (N_6189,N_5561,N_5407);
nor U6190 (N_6190,N_5482,N_5740);
xnor U6191 (N_6191,N_5800,N_5641);
or U6192 (N_6192,N_5705,N_5532);
and U6193 (N_6193,N_5413,N_5416);
nor U6194 (N_6194,N_5502,N_5919);
and U6195 (N_6195,N_5464,N_5478);
nand U6196 (N_6196,N_5599,N_5867);
nand U6197 (N_6197,N_5545,N_5756);
and U6198 (N_6198,N_5492,N_5435);
nor U6199 (N_6199,N_5548,N_5707);
or U6200 (N_6200,N_5579,N_5442);
xor U6201 (N_6201,N_5974,N_5597);
and U6202 (N_6202,N_5461,N_5626);
nand U6203 (N_6203,N_5700,N_5935);
and U6204 (N_6204,N_5976,N_5787);
or U6205 (N_6205,N_5598,N_5757);
and U6206 (N_6206,N_5946,N_5484);
nand U6207 (N_6207,N_5735,N_5555);
and U6208 (N_6208,N_5655,N_5872);
xor U6209 (N_6209,N_5711,N_5483);
nand U6210 (N_6210,N_5753,N_5589);
nand U6211 (N_6211,N_5777,N_5613);
or U6212 (N_6212,N_5851,N_5981);
or U6213 (N_6213,N_5875,N_5904);
nand U6214 (N_6214,N_5537,N_5604);
nand U6215 (N_6215,N_5858,N_5533);
or U6216 (N_6216,N_5906,N_5501);
nor U6217 (N_6217,N_5479,N_5665);
nand U6218 (N_6218,N_5810,N_5860);
and U6219 (N_6219,N_5824,N_5669);
xor U6220 (N_6220,N_5452,N_5507);
and U6221 (N_6221,N_5836,N_5896);
xor U6222 (N_6222,N_5400,N_5798);
nor U6223 (N_6223,N_5772,N_5575);
or U6224 (N_6224,N_5924,N_5890);
nand U6225 (N_6225,N_5801,N_5941);
and U6226 (N_6226,N_5423,N_5795);
nor U6227 (N_6227,N_5521,N_5468);
and U6228 (N_6228,N_5819,N_5752);
nand U6229 (N_6229,N_5969,N_5937);
nor U6230 (N_6230,N_5899,N_5670);
nand U6231 (N_6231,N_5767,N_5751);
xnor U6232 (N_6232,N_5674,N_5606);
and U6233 (N_6233,N_5862,N_5755);
nor U6234 (N_6234,N_5689,N_5564);
and U6235 (N_6235,N_5940,N_5733);
xor U6236 (N_6236,N_5657,N_5559);
nor U6237 (N_6237,N_5825,N_5802);
xor U6238 (N_6238,N_5985,N_5427);
and U6239 (N_6239,N_5715,N_5475);
or U6240 (N_6240,N_5679,N_5832);
nand U6241 (N_6241,N_5487,N_5746);
nor U6242 (N_6242,N_5546,N_5420);
nand U6243 (N_6243,N_5791,N_5511);
or U6244 (N_6244,N_5648,N_5878);
or U6245 (N_6245,N_5595,N_5747);
and U6246 (N_6246,N_5590,N_5543);
and U6247 (N_6247,N_5422,N_5656);
and U6248 (N_6248,N_5542,N_5676);
nand U6249 (N_6249,N_5638,N_5926);
nand U6250 (N_6250,N_5418,N_5553);
xnor U6251 (N_6251,N_5742,N_5592);
nor U6252 (N_6252,N_5830,N_5433);
nand U6253 (N_6253,N_5509,N_5562);
nor U6254 (N_6254,N_5645,N_5454);
or U6255 (N_6255,N_5829,N_5846);
nand U6256 (N_6256,N_5892,N_5992);
or U6257 (N_6257,N_5837,N_5925);
nand U6258 (N_6258,N_5637,N_5675);
nand U6259 (N_6259,N_5636,N_5620);
or U6260 (N_6260,N_5880,N_5841);
and U6261 (N_6261,N_5448,N_5603);
and U6262 (N_6262,N_5515,N_5993);
and U6263 (N_6263,N_5717,N_5877);
or U6264 (N_6264,N_5900,N_5842);
xor U6265 (N_6265,N_5799,N_5758);
xnor U6266 (N_6266,N_5429,N_5790);
or U6267 (N_6267,N_5780,N_5734);
or U6268 (N_6268,N_5931,N_5792);
or U6269 (N_6269,N_5421,N_5608);
nor U6270 (N_6270,N_5460,N_5744);
and U6271 (N_6271,N_5996,N_5843);
nor U6272 (N_6272,N_5907,N_5566);
nand U6273 (N_6273,N_5719,N_5687);
nor U6274 (N_6274,N_5671,N_5582);
xnor U6275 (N_6275,N_5450,N_5886);
nor U6276 (N_6276,N_5948,N_5653);
nor U6277 (N_6277,N_5813,N_5831);
and U6278 (N_6278,N_5938,N_5578);
or U6279 (N_6279,N_5486,N_5453);
xnor U6280 (N_6280,N_5835,N_5805);
or U6281 (N_6281,N_5682,N_5473);
or U6282 (N_6282,N_5895,N_5614);
xor U6283 (N_6283,N_5783,N_5958);
xor U6284 (N_6284,N_5927,N_5490);
and U6285 (N_6285,N_5410,N_5406);
nor U6286 (N_6286,N_5921,N_5773);
and U6287 (N_6287,N_5560,N_5916);
nand U6288 (N_6288,N_5651,N_5494);
xnor U6289 (N_6289,N_5667,N_5997);
and U6290 (N_6290,N_5650,N_5534);
or U6291 (N_6291,N_5815,N_5863);
or U6292 (N_6292,N_5732,N_5463);
and U6293 (N_6293,N_5778,N_5853);
xnor U6294 (N_6294,N_5918,N_5577);
or U6295 (N_6295,N_5737,N_5989);
and U6296 (N_6296,N_5708,N_5828);
nand U6297 (N_6297,N_5666,N_5873);
and U6298 (N_6298,N_5586,N_5934);
or U6299 (N_6299,N_5536,N_5950);
xnor U6300 (N_6300,N_5522,N_5866);
xor U6301 (N_6301,N_5754,N_5448);
nor U6302 (N_6302,N_5747,N_5521);
or U6303 (N_6303,N_5569,N_5861);
nor U6304 (N_6304,N_5490,N_5938);
nand U6305 (N_6305,N_5916,N_5428);
xnor U6306 (N_6306,N_5713,N_5981);
xnor U6307 (N_6307,N_5669,N_5705);
and U6308 (N_6308,N_5599,N_5603);
xnor U6309 (N_6309,N_5702,N_5590);
and U6310 (N_6310,N_5564,N_5616);
xnor U6311 (N_6311,N_5673,N_5417);
nand U6312 (N_6312,N_5621,N_5672);
and U6313 (N_6313,N_5987,N_5962);
xor U6314 (N_6314,N_5645,N_5610);
or U6315 (N_6315,N_5686,N_5699);
nor U6316 (N_6316,N_5743,N_5681);
and U6317 (N_6317,N_5622,N_5482);
or U6318 (N_6318,N_5641,N_5608);
xor U6319 (N_6319,N_5985,N_5817);
and U6320 (N_6320,N_5455,N_5850);
or U6321 (N_6321,N_5428,N_5887);
or U6322 (N_6322,N_5767,N_5858);
and U6323 (N_6323,N_5936,N_5488);
and U6324 (N_6324,N_5590,N_5524);
and U6325 (N_6325,N_5551,N_5895);
xnor U6326 (N_6326,N_5604,N_5842);
and U6327 (N_6327,N_5933,N_5762);
nand U6328 (N_6328,N_5620,N_5435);
nor U6329 (N_6329,N_5685,N_5607);
nor U6330 (N_6330,N_5805,N_5648);
or U6331 (N_6331,N_5938,N_5730);
nand U6332 (N_6332,N_5745,N_5837);
xnor U6333 (N_6333,N_5530,N_5693);
nor U6334 (N_6334,N_5704,N_5656);
xor U6335 (N_6335,N_5839,N_5638);
and U6336 (N_6336,N_5708,N_5639);
and U6337 (N_6337,N_5799,N_5947);
or U6338 (N_6338,N_5679,N_5553);
nor U6339 (N_6339,N_5500,N_5404);
and U6340 (N_6340,N_5824,N_5647);
nand U6341 (N_6341,N_5748,N_5831);
nand U6342 (N_6342,N_5653,N_5605);
and U6343 (N_6343,N_5527,N_5573);
xnor U6344 (N_6344,N_5574,N_5478);
nor U6345 (N_6345,N_5520,N_5823);
and U6346 (N_6346,N_5808,N_5788);
and U6347 (N_6347,N_5767,N_5502);
xnor U6348 (N_6348,N_5777,N_5767);
and U6349 (N_6349,N_5830,N_5605);
or U6350 (N_6350,N_5509,N_5608);
nand U6351 (N_6351,N_5576,N_5648);
and U6352 (N_6352,N_5434,N_5961);
and U6353 (N_6353,N_5675,N_5563);
xnor U6354 (N_6354,N_5818,N_5608);
nor U6355 (N_6355,N_5781,N_5687);
nand U6356 (N_6356,N_5739,N_5845);
nand U6357 (N_6357,N_5659,N_5704);
nor U6358 (N_6358,N_5925,N_5554);
and U6359 (N_6359,N_5599,N_5962);
xnor U6360 (N_6360,N_5681,N_5572);
xor U6361 (N_6361,N_5865,N_5935);
or U6362 (N_6362,N_5828,N_5518);
and U6363 (N_6363,N_5516,N_5822);
or U6364 (N_6364,N_5689,N_5873);
xnor U6365 (N_6365,N_5920,N_5689);
nand U6366 (N_6366,N_5505,N_5500);
xnor U6367 (N_6367,N_5513,N_5510);
nand U6368 (N_6368,N_5468,N_5420);
xor U6369 (N_6369,N_5780,N_5746);
xor U6370 (N_6370,N_5989,N_5924);
xnor U6371 (N_6371,N_5673,N_5839);
or U6372 (N_6372,N_5810,N_5421);
or U6373 (N_6373,N_5686,N_5798);
xnor U6374 (N_6374,N_5956,N_5832);
nand U6375 (N_6375,N_5710,N_5684);
nor U6376 (N_6376,N_5492,N_5524);
nand U6377 (N_6377,N_5886,N_5741);
or U6378 (N_6378,N_5546,N_5464);
and U6379 (N_6379,N_5527,N_5817);
xor U6380 (N_6380,N_5808,N_5812);
nor U6381 (N_6381,N_5471,N_5438);
or U6382 (N_6382,N_5925,N_5902);
xor U6383 (N_6383,N_5745,N_5900);
xor U6384 (N_6384,N_5555,N_5664);
nand U6385 (N_6385,N_5884,N_5509);
xnor U6386 (N_6386,N_5460,N_5404);
and U6387 (N_6387,N_5972,N_5772);
xor U6388 (N_6388,N_5885,N_5468);
nor U6389 (N_6389,N_5552,N_5733);
nand U6390 (N_6390,N_5847,N_5412);
nand U6391 (N_6391,N_5830,N_5921);
xor U6392 (N_6392,N_5967,N_5970);
xor U6393 (N_6393,N_5503,N_5551);
nand U6394 (N_6394,N_5959,N_5544);
or U6395 (N_6395,N_5537,N_5958);
nand U6396 (N_6396,N_5498,N_5412);
nor U6397 (N_6397,N_5714,N_5482);
and U6398 (N_6398,N_5421,N_5663);
and U6399 (N_6399,N_5689,N_5695);
xor U6400 (N_6400,N_5881,N_5524);
or U6401 (N_6401,N_5667,N_5783);
and U6402 (N_6402,N_5658,N_5921);
xnor U6403 (N_6403,N_5590,N_5947);
or U6404 (N_6404,N_5507,N_5669);
xor U6405 (N_6405,N_5792,N_5496);
xnor U6406 (N_6406,N_5740,N_5679);
nand U6407 (N_6407,N_5489,N_5659);
and U6408 (N_6408,N_5985,N_5734);
nor U6409 (N_6409,N_5566,N_5790);
and U6410 (N_6410,N_5435,N_5922);
nor U6411 (N_6411,N_5577,N_5511);
and U6412 (N_6412,N_5746,N_5692);
nand U6413 (N_6413,N_5672,N_5820);
and U6414 (N_6414,N_5883,N_5957);
xor U6415 (N_6415,N_5990,N_5857);
xor U6416 (N_6416,N_5633,N_5891);
and U6417 (N_6417,N_5438,N_5675);
xnor U6418 (N_6418,N_5928,N_5508);
nand U6419 (N_6419,N_5990,N_5709);
and U6420 (N_6420,N_5868,N_5751);
or U6421 (N_6421,N_5648,N_5928);
xnor U6422 (N_6422,N_5711,N_5762);
or U6423 (N_6423,N_5845,N_5603);
nand U6424 (N_6424,N_5780,N_5788);
xnor U6425 (N_6425,N_5435,N_5872);
or U6426 (N_6426,N_5912,N_5531);
and U6427 (N_6427,N_5762,N_5710);
xnor U6428 (N_6428,N_5441,N_5875);
xnor U6429 (N_6429,N_5799,N_5587);
nor U6430 (N_6430,N_5436,N_5661);
or U6431 (N_6431,N_5871,N_5581);
and U6432 (N_6432,N_5472,N_5827);
or U6433 (N_6433,N_5462,N_5985);
and U6434 (N_6434,N_5497,N_5453);
and U6435 (N_6435,N_5481,N_5766);
nand U6436 (N_6436,N_5705,N_5988);
xor U6437 (N_6437,N_5482,N_5657);
nand U6438 (N_6438,N_5877,N_5570);
nand U6439 (N_6439,N_5559,N_5440);
xnor U6440 (N_6440,N_5857,N_5667);
nor U6441 (N_6441,N_5853,N_5447);
or U6442 (N_6442,N_5580,N_5603);
nor U6443 (N_6443,N_5741,N_5799);
and U6444 (N_6444,N_5676,N_5947);
or U6445 (N_6445,N_5749,N_5683);
nand U6446 (N_6446,N_5697,N_5779);
xor U6447 (N_6447,N_5612,N_5581);
nand U6448 (N_6448,N_5929,N_5975);
nor U6449 (N_6449,N_5951,N_5446);
and U6450 (N_6450,N_5909,N_5593);
and U6451 (N_6451,N_5833,N_5442);
or U6452 (N_6452,N_5577,N_5864);
and U6453 (N_6453,N_5463,N_5988);
and U6454 (N_6454,N_5937,N_5555);
nor U6455 (N_6455,N_5718,N_5815);
and U6456 (N_6456,N_5604,N_5711);
xnor U6457 (N_6457,N_5996,N_5701);
or U6458 (N_6458,N_5732,N_5447);
nor U6459 (N_6459,N_5569,N_5785);
and U6460 (N_6460,N_5878,N_5570);
nor U6461 (N_6461,N_5866,N_5642);
nand U6462 (N_6462,N_5993,N_5760);
xnor U6463 (N_6463,N_5581,N_5604);
and U6464 (N_6464,N_5403,N_5856);
xor U6465 (N_6465,N_5462,N_5465);
or U6466 (N_6466,N_5895,N_5482);
xnor U6467 (N_6467,N_5419,N_5416);
or U6468 (N_6468,N_5597,N_5706);
nand U6469 (N_6469,N_5840,N_5570);
nand U6470 (N_6470,N_5954,N_5407);
nor U6471 (N_6471,N_5908,N_5570);
and U6472 (N_6472,N_5507,N_5731);
or U6473 (N_6473,N_5838,N_5769);
or U6474 (N_6474,N_5856,N_5955);
or U6475 (N_6475,N_5616,N_5610);
xnor U6476 (N_6476,N_5965,N_5400);
or U6477 (N_6477,N_5674,N_5509);
nand U6478 (N_6478,N_5773,N_5642);
nor U6479 (N_6479,N_5407,N_5433);
nor U6480 (N_6480,N_5680,N_5552);
xnor U6481 (N_6481,N_5609,N_5629);
xnor U6482 (N_6482,N_5562,N_5527);
and U6483 (N_6483,N_5559,N_5428);
and U6484 (N_6484,N_5652,N_5884);
nor U6485 (N_6485,N_5952,N_5925);
nand U6486 (N_6486,N_5488,N_5508);
or U6487 (N_6487,N_5987,N_5877);
xor U6488 (N_6488,N_5824,N_5481);
nand U6489 (N_6489,N_5524,N_5688);
and U6490 (N_6490,N_5640,N_5977);
or U6491 (N_6491,N_5829,N_5784);
and U6492 (N_6492,N_5866,N_5617);
nand U6493 (N_6493,N_5753,N_5856);
xor U6494 (N_6494,N_5576,N_5405);
nand U6495 (N_6495,N_5884,N_5922);
nand U6496 (N_6496,N_5609,N_5986);
nor U6497 (N_6497,N_5719,N_5838);
nor U6498 (N_6498,N_5888,N_5737);
nand U6499 (N_6499,N_5590,N_5455);
and U6500 (N_6500,N_5574,N_5909);
nand U6501 (N_6501,N_5432,N_5959);
or U6502 (N_6502,N_5947,N_5954);
nand U6503 (N_6503,N_5888,N_5742);
and U6504 (N_6504,N_5915,N_5866);
and U6505 (N_6505,N_5555,N_5915);
or U6506 (N_6506,N_5907,N_5520);
and U6507 (N_6507,N_5727,N_5648);
or U6508 (N_6508,N_5536,N_5971);
or U6509 (N_6509,N_5560,N_5535);
nand U6510 (N_6510,N_5687,N_5892);
or U6511 (N_6511,N_5515,N_5773);
xnor U6512 (N_6512,N_5698,N_5610);
or U6513 (N_6513,N_5624,N_5996);
nand U6514 (N_6514,N_5523,N_5909);
nor U6515 (N_6515,N_5834,N_5778);
nor U6516 (N_6516,N_5486,N_5427);
nand U6517 (N_6517,N_5845,N_5732);
and U6518 (N_6518,N_5604,N_5681);
and U6519 (N_6519,N_5810,N_5922);
nor U6520 (N_6520,N_5567,N_5604);
and U6521 (N_6521,N_5489,N_5539);
nand U6522 (N_6522,N_5419,N_5800);
nor U6523 (N_6523,N_5680,N_5907);
and U6524 (N_6524,N_5660,N_5781);
nor U6525 (N_6525,N_5929,N_5448);
or U6526 (N_6526,N_5588,N_5887);
nor U6527 (N_6527,N_5723,N_5979);
nand U6528 (N_6528,N_5469,N_5975);
or U6529 (N_6529,N_5568,N_5984);
xor U6530 (N_6530,N_5616,N_5924);
or U6531 (N_6531,N_5558,N_5840);
and U6532 (N_6532,N_5422,N_5565);
and U6533 (N_6533,N_5510,N_5689);
or U6534 (N_6534,N_5616,N_5999);
and U6535 (N_6535,N_5974,N_5502);
or U6536 (N_6536,N_5985,N_5990);
nand U6537 (N_6537,N_5706,N_5411);
nor U6538 (N_6538,N_5948,N_5672);
xor U6539 (N_6539,N_5956,N_5622);
or U6540 (N_6540,N_5697,N_5685);
xnor U6541 (N_6541,N_5728,N_5589);
nor U6542 (N_6542,N_5998,N_5906);
nand U6543 (N_6543,N_5512,N_5976);
and U6544 (N_6544,N_5450,N_5423);
xor U6545 (N_6545,N_5507,N_5465);
and U6546 (N_6546,N_5853,N_5857);
nor U6547 (N_6547,N_5810,N_5429);
and U6548 (N_6548,N_5958,N_5852);
nor U6549 (N_6549,N_5964,N_5887);
nand U6550 (N_6550,N_5449,N_5853);
or U6551 (N_6551,N_5697,N_5431);
and U6552 (N_6552,N_5642,N_5964);
and U6553 (N_6553,N_5497,N_5586);
and U6554 (N_6554,N_5977,N_5567);
nor U6555 (N_6555,N_5864,N_5812);
and U6556 (N_6556,N_5576,N_5406);
nand U6557 (N_6557,N_5649,N_5570);
or U6558 (N_6558,N_5486,N_5811);
xor U6559 (N_6559,N_5499,N_5428);
or U6560 (N_6560,N_5912,N_5739);
xor U6561 (N_6561,N_5666,N_5928);
and U6562 (N_6562,N_5521,N_5508);
and U6563 (N_6563,N_5878,N_5474);
nand U6564 (N_6564,N_5548,N_5770);
or U6565 (N_6565,N_5650,N_5674);
nand U6566 (N_6566,N_5922,N_5888);
nor U6567 (N_6567,N_5580,N_5987);
nor U6568 (N_6568,N_5824,N_5720);
or U6569 (N_6569,N_5581,N_5467);
nor U6570 (N_6570,N_5727,N_5949);
xor U6571 (N_6571,N_5687,N_5794);
or U6572 (N_6572,N_5751,N_5521);
or U6573 (N_6573,N_5887,N_5454);
or U6574 (N_6574,N_5452,N_5550);
nor U6575 (N_6575,N_5701,N_5674);
nand U6576 (N_6576,N_5931,N_5698);
and U6577 (N_6577,N_5596,N_5881);
or U6578 (N_6578,N_5522,N_5655);
nand U6579 (N_6579,N_5630,N_5793);
xnor U6580 (N_6580,N_5846,N_5989);
and U6581 (N_6581,N_5897,N_5425);
nand U6582 (N_6582,N_5785,N_5631);
and U6583 (N_6583,N_5976,N_5486);
nand U6584 (N_6584,N_5478,N_5618);
nand U6585 (N_6585,N_5566,N_5982);
nand U6586 (N_6586,N_5661,N_5420);
and U6587 (N_6587,N_5792,N_5630);
and U6588 (N_6588,N_5958,N_5441);
nand U6589 (N_6589,N_5952,N_5432);
xnor U6590 (N_6590,N_5721,N_5648);
and U6591 (N_6591,N_5603,N_5954);
or U6592 (N_6592,N_5835,N_5419);
or U6593 (N_6593,N_5760,N_5630);
or U6594 (N_6594,N_5579,N_5722);
nor U6595 (N_6595,N_5931,N_5502);
or U6596 (N_6596,N_5989,N_5674);
nor U6597 (N_6597,N_5618,N_5743);
or U6598 (N_6598,N_5979,N_5818);
nand U6599 (N_6599,N_5763,N_5707);
nor U6600 (N_6600,N_6549,N_6532);
xnor U6601 (N_6601,N_6081,N_6238);
nor U6602 (N_6602,N_6257,N_6239);
xnor U6603 (N_6603,N_6444,N_6358);
nor U6604 (N_6604,N_6561,N_6158);
nand U6605 (N_6605,N_6297,N_6077);
or U6606 (N_6606,N_6362,N_6062);
nor U6607 (N_6607,N_6125,N_6118);
xnor U6608 (N_6608,N_6567,N_6051);
or U6609 (N_6609,N_6533,N_6226);
nor U6610 (N_6610,N_6520,N_6582);
and U6611 (N_6611,N_6080,N_6043);
xor U6612 (N_6612,N_6550,N_6577);
xor U6613 (N_6613,N_6527,N_6281);
nor U6614 (N_6614,N_6050,N_6468);
or U6615 (N_6615,N_6015,N_6588);
and U6616 (N_6616,N_6345,N_6013);
or U6617 (N_6617,N_6544,N_6303);
nand U6618 (N_6618,N_6055,N_6083);
and U6619 (N_6619,N_6480,N_6515);
or U6620 (N_6620,N_6518,N_6485);
nor U6621 (N_6621,N_6207,N_6131);
nor U6622 (N_6622,N_6006,N_6137);
xnor U6623 (N_6623,N_6348,N_6499);
nand U6624 (N_6624,N_6531,N_6314);
nor U6625 (N_6625,N_6156,N_6133);
xor U6626 (N_6626,N_6203,N_6318);
nor U6627 (N_6627,N_6211,N_6412);
nand U6628 (N_6628,N_6074,N_6579);
xor U6629 (N_6629,N_6047,N_6166);
and U6630 (N_6630,N_6424,N_6105);
nor U6631 (N_6631,N_6396,N_6108);
xor U6632 (N_6632,N_6383,N_6065);
nor U6633 (N_6633,N_6415,N_6583);
and U6634 (N_6634,N_6299,N_6143);
nand U6635 (N_6635,N_6017,N_6256);
xor U6636 (N_6636,N_6357,N_6491);
and U6637 (N_6637,N_6023,N_6472);
nand U6638 (N_6638,N_6097,N_6088);
and U6639 (N_6639,N_6402,N_6474);
xor U6640 (N_6640,N_6384,N_6179);
or U6641 (N_6641,N_6274,N_6553);
nor U6642 (N_6642,N_6150,N_6269);
nor U6643 (N_6643,N_6420,N_6599);
and U6644 (N_6644,N_6315,N_6511);
and U6645 (N_6645,N_6115,N_6288);
or U6646 (N_6646,N_6285,N_6102);
and U6647 (N_6647,N_6103,N_6305);
nand U6648 (N_6648,N_6221,N_6490);
nand U6649 (N_6649,N_6507,N_6425);
and U6650 (N_6650,N_6178,N_6236);
nand U6651 (N_6651,N_6439,N_6573);
and U6652 (N_6652,N_6564,N_6366);
and U6653 (N_6653,N_6482,N_6460);
nor U6654 (N_6654,N_6145,N_6165);
nand U6655 (N_6655,N_6325,N_6087);
or U6656 (N_6656,N_6370,N_6494);
or U6657 (N_6657,N_6250,N_6227);
nand U6658 (N_6658,N_6379,N_6521);
or U6659 (N_6659,N_6168,N_6546);
nor U6660 (N_6660,N_6073,N_6302);
nand U6661 (N_6661,N_6427,N_6175);
xnor U6662 (N_6662,N_6308,N_6502);
or U6663 (N_6663,N_6008,N_6413);
nor U6664 (N_6664,N_6049,N_6408);
nand U6665 (N_6665,N_6240,N_6428);
nor U6666 (N_6666,N_6246,N_6421);
or U6667 (N_6667,N_6078,N_6068);
and U6668 (N_6668,N_6445,N_6566);
nor U6669 (N_6669,N_6394,N_6371);
and U6670 (N_6670,N_6096,N_6481);
nor U6671 (N_6671,N_6067,N_6182);
xnor U6672 (N_6672,N_6104,N_6254);
or U6673 (N_6673,N_6132,N_6558);
and U6674 (N_6674,N_6094,N_6066);
or U6675 (N_6675,N_6127,N_6032);
nand U6676 (N_6676,N_6595,N_6506);
nor U6677 (N_6677,N_6570,N_6330);
xor U6678 (N_6678,N_6433,N_6181);
nand U6679 (N_6679,N_6119,N_6009);
nand U6680 (N_6680,N_6149,N_6448);
and U6681 (N_6681,N_6557,N_6545);
xnor U6682 (N_6682,N_6327,N_6026);
xor U6683 (N_6683,N_6587,N_6466);
nand U6684 (N_6684,N_6031,N_6296);
nand U6685 (N_6685,N_6192,N_6385);
nor U6686 (N_6686,N_6117,N_6113);
nor U6687 (N_6687,N_6069,N_6033);
and U6688 (N_6688,N_6241,N_6523);
xnor U6689 (N_6689,N_6027,N_6162);
or U6690 (N_6690,N_6317,N_6524);
or U6691 (N_6691,N_6138,N_6501);
xor U6692 (N_6692,N_6283,N_6110);
xnor U6693 (N_6693,N_6224,N_6216);
nor U6694 (N_6694,N_6537,N_6002);
or U6695 (N_6695,N_6007,N_6148);
nor U6696 (N_6696,N_6029,N_6407);
or U6697 (N_6697,N_6134,N_6041);
nand U6698 (N_6698,N_6436,N_6070);
nand U6699 (N_6699,N_6359,N_6497);
and U6700 (N_6700,N_6522,N_6024);
or U6701 (N_6701,N_6293,N_6266);
or U6702 (N_6702,N_6021,N_6289);
and U6703 (N_6703,N_6393,N_6405);
or U6704 (N_6704,N_6441,N_6326);
xnor U6705 (N_6705,N_6160,N_6157);
or U6706 (N_6706,N_6112,N_6596);
nand U6707 (N_6707,N_6306,N_6300);
xor U6708 (N_6708,N_6556,N_6082);
and U6709 (N_6709,N_6416,N_6386);
nand U6710 (N_6710,N_6279,N_6276);
nor U6711 (N_6711,N_6053,N_6543);
or U6712 (N_6712,N_6225,N_6153);
nor U6713 (N_6713,N_6352,N_6331);
nand U6714 (N_6714,N_6169,N_6126);
xor U6715 (N_6715,N_6061,N_6085);
or U6716 (N_6716,N_6171,N_6205);
nand U6717 (N_6717,N_6229,N_6349);
and U6718 (N_6718,N_6204,N_6064);
nor U6719 (N_6719,N_6429,N_6014);
xor U6720 (N_6720,N_6406,N_6139);
and U6721 (N_6721,N_6091,N_6350);
nor U6722 (N_6722,N_6530,N_6307);
nor U6723 (N_6723,N_6128,N_6399);
xor U6724 (N_6724,N_6534,N_6419);
xor U6725 (N_6725,N_6493,N_6059);
or U6726 (N_6726,N_6397,N_6278);
nand U6727 (N_6727,N_6377,N_6388);
and U6728 (N_6728,N_6255,N_6417);
nor U6729 (N_6729,N_6206,N_6010);
and U6730 (N_6730,N_6090,N_6547);
and U6731 (N_6731,N_6319,N_6184);
or U6732 (N_6732,N_6526,N_6598);
nand U6733 (N_6733,N_6343,N_6016);
and U6734 (N_6734,N_6589,N_6500);
xnor U6735 (N_6735,N_6146,N_6242);
xor U6736 (N_6736,N_6540,N_6000);
nor U6737 (N_6737,N_6249,N_6484);
and U6738 (N_6738,N_6247,N_6590);
xor U6739 (N_6739,N_6323,N_6195);
nand U6740 (N_6740,N_6322,N_6341);
nand U6741 (N_6741,N_6199,N_6310);
nor U6742 (N_6742,N_6382,N_6245);
nand U6743 (N_6743,N_6372,N_6464);
and U6744 (N_6744,N_6344,N_6025);
nor U6745 (N_6745,N_6487,N_6580);
and U6746 (N_6746,N_6235,N_6368);
xor U6747 (N_6747,N_6332,N_6333);
or U6748 (N_6748,N_6347,N_6196);
or U6749 (N_6749,N_6107,N_6152);
xor U6750 (N_6750,N_6003,N_6334);
or U6751 (N_6751,N_6124,N_6035);
nor U6752 (N_6752,N_6495,N_6155);
xnor U6753 (N_6753,N_6271,N_6282);
nand U6754 (N_6754,N_6198,N_6563);
xor U6755 (N_6755,N_6046,N_6095);
nor U6756 (N_6756,N_6018,N_6565);
or U6757 (N_6757,N_6400,N_6311);
nor U6758 (N_6758,N_6304,N_6581);
and U6759 (N_6759,N_6447,N_6508);
xnor U6760 (N_6760,N_6454,N_6346);
nand U6761 (N_6761,N_6479,N_6079);
nand U6762 (N_6762,N_6172,N_6121);
nand U6763 (N_6763,N_6355,N_6164);
and U6764 (N_6764,N_6571,N_6111);
nand U6765 (N_6765,N_6093,N_6551);
and U6766 (N_6766,N_6180,N_6173);
nor U6767 (N_6767,N_6071,N_6012);
xnor U6768 (N_6768,N_6361,N_6202);
nor U6769 (N_6769,N_6159,N_6360);
or U6770 (N_6770,N_6489,N_6513);
and U6771 (N_6771,N_6471,N_6151);
nand U6772 (N_6772,N_6450,N_6324);
and U6773 (N_6773,N_6130,N_6259);
nand U6774 (N_6774,N_6176,N_6404);
nor U6775 (N_6775,N_6432,N_6042);
or U6776 (N_6776,N_6273,N_6292);
nor U6777 (N_6777,N_6552,N_6340);
and U6778 (N_6778,N_6272,N_6434);
and U6779 (N_6779,N_6336,N_6232);
nand U6780 (N_6780,N_6234,N_6048);
and U6781 (N_6781,N_6554,N_6418);
or U6782 (N_6782,N_6536,N_6456);
xor U6783 (N_6783,N_6034,N_6437);
nand U6784 (N_6784,N_6389,N_6395);
nand U6785 (N_6785,N_6270,N_6170);
xnor U6786 (N_6786,N_6298,N_6209);
nor U6787 (N_6787,N_6378,N_6541);
and U6788 (N_6788,N_6076,N_6542);
xnor U6789 (N_6789,N_6123,N_6509);
nand U6790 (N_6790,N_6516,N_6309);
and U6791 (N_6791,N_6375,N_6351);
or U6792 (N_6792,N_6183,N_6228);
xor U6793 (N_6793,N_6089,N_6387);
and U6794 (N_6794,N_6560,N_6578);
xnor U6795 (N_6795,N_6422,N_6510);
nand U6796 (N_6796,N_6072,N_6496);
nor U6797 (N_6797,N_6056,N_6030);
and U6798 (N_6798,N_6392,N_6449);
xor U6799 (N_6799,N_6328,N_6457);
and U6800 (N_6800,N_6440,N_6265);
or U6801 (N_6801,N_6020,N_6286);
nor U6802 (N_6802,N_6201,N_6106);
and U6803 (N_6803,N_6261,N_6186);
nor U6804 (N_6804,N_6248,N_6568);
nor U6805 (N_6805,N_6597,N_6353);
or U6806 (N_6806,N_6364,N_6409);
xor U6807 (N_6807,N_6218,N_6092);
nand U6808 (N_6808,N_6462,N_6354);
xor U6809 (N_6809,N_6519,N_6280);
nor U6810 (N_6810,N_6461,N_6197);
xnor U6811 (N_6811,N_6222,N_6045);
and U6812 (N_6812,N_6086,N_6562);
or U6813 (N_6813,N_6463,N_6215);
xor U6814 (N_6814,N_6109,N_6430);
or U6815 (N_6815,N_6057,N_6038);
nand U6816 (N_6816,N_6189,N_6483);
nor U6817 (N_6817,N_6054,N_6473);
nand U6818 (N_6818,N_6210,N_6217);
xnor U6819 (N_6819,N_6529,N_6264);
xnor U6820 (N_6820,N_6174,N_6548);
nand U6821 (N_6821,N_6337,N_6141);
xnor U6822 (N_6822,N_6019,N_6426);
nand U6823 (N_6823,N_6122,N_6154);
and U6824 (N_6824,N_6576,N_6135);
nand U6825 (N_6825,N_6028,N_6287);
nor U6826 (N_6826,N_6190,N_6039);
nand U6827 (N_6827,N_6260,N_6188);
nand U6828 (N_6828,N_6277,N_6244);
nand U6829 (N_6829,N_6301,N_6313);
nor U6830 (N_6830,N_6044,N_6321);
and U6831 (N_6831,N_6574,N_6446);
and U6832 (N_6832,N_6163,N_6114);
xor U6833 (N_6833,N_6147,N_6099);
nand U6834 (N_6834,N_6380,N_6267);
and U6835 (N_6835,N_6252,N_6136);
nor U6836 (N_6836,N_6098,N_6312);
and U6837 (N_6837,N_6390,N_6528);
xnor U6838 (N_6838,N_6435,N_6478);
or U6839 (N_6839,N_6329,N_6492);
xnor U6840 (N_6840,N_6220,N_6129);
nor U6841 (N_6841,N_6052,N_6120);
and U6842 (N_6842,N_6284,N_6453);
nor U6843 (N_6843,N_6438,N_6243);
nor U6844 (N_6844,N_6410,N_6559);
xor U6845 (N_6845,N_6374,N_6208);
nand U6846 (N_6846,N_6213,N_6339);
nor U6847 (N_6847,N_6177,N_6381);
or U6848 (N_6848,N_6477,N_6036);
xor U6849 (N_6849,N_6452,N_6594);
nand U6850 (N_6850,N_6037,N_6475);
and U6851 (N_6851,N_6369,N_6116);
xor U6852 (N_6852,N_6465,N_6467);
and U6853 (N_6853,N_6367,N_6411);
or U6854 (N_6854,N_6291,N_6191);
nor U6855 (N_6855,N_6470,N_6363);
xor U6856 (N_6856,N_6223,N_6486);
nor U6857 (N_6857,N_6338,N_6365);
nand U6858 (N_6858,N_6263,N_6185);
nor U6859 (N_6859,N_6488,N_6101);
and U6860 (N_6860,N_6525,N_6512);
xor U6861 (N_6861,N_6194,N_6401);
nand U6862 (N_6862,N_6219,N_6262);
and U6863 (N_6863,N_6161,N_6100);
and U6864 (N_6864,N_6193,N_6212);
and U6865 (N_6865,N_6144,N_6398);
or U6866 (N_6866,N_6373,N_6140);
nor U6867 (N_6867,N_6505,N_6233);
or U6868 (N_6868,N_6004,N_6214);
nor U6869 (N_6869,N_6569,N_6455);
xnor U6870 (N_6870,N_6538,N_6476);
or U6871 (N_6871,N_6356,N_6459);
or U6872 (N_6872,N_6504,N_6335);
nor U6873 (N_6873,N_6230,N_6058);
nor U6874 (N_6874,N_6258,N_6294);
and U6875 (N_6875,N_6142,N_6584);
xor U6876 (N_6876,N_6503,N_6592);
nand U6877 (N_6877,N_6011,N_6231);
or U6878 (N_6878,N_6040,N_6320);
nand U6879 (N_6879,N_6585,N_6575);
nor U6880 (N_6880,N_6458,N_6084);
or U6881 (N_6881,N_6414,N_6555);
nand U6882 (N_6882,N_6268,N_6075);
nor U6883 (N_6883,N_6275,N_6517);
and U6884 (N_6884,N_6539,N_6443);
or U6885 (N_6885,N_6001,N_6403);
or U6886 (N_6886,N_6022,N_6237);
xnor U6887 (N_6887,N_6005,N_6342);
xor U6888 (N_6888,N_6200,N_6063);
xor U6889 (N_6889,N_6451,N_6431);
nand U6890 (N_6890,N_6060,N_6391);
or U6891 (N_6891,N_6498,N_6316);
and U6892 (N_6892,N_6187,N_6572);
xor U6893 (N_6893,N_6295,N_6376);
xnor U6894 (N_6894,N_6253,N_6593);
nand U6895 (N_6895,N_6535,N_6514);
nand U6896 (N_6896,N_6251,N_6423);
or U6897 (N_6897,N_6591,N_6167);
xnor U6898 (N_6898,N_6290,N_6586);
and U6899 (N_6899,N_6469,N_6442);
nand U6900 (N_6900,N_6153,N_6133);
and U6901 (N_6901,N_6536,N_6323);
nand U6902 (N_6902,N_6099,N_6454);
xnor U6903 (N_6903,N_6437,N_6394);
or U6904 (N_6904,N_6329,N_6502);
nor U6905 (N_6905,N_6563,N_6249);
and U6906 (N_6906,N_6585,N_6318);
and U6907 (N_6907,N_6464,N_6200);
and U6908 (N_6908,N_6395,N_6327);
nor U6909 (N_6909,N_6565,N_6439);
nor U6910 (N_6910,N_6485,N_6365);
xor U6911 (N_6911,N_6303,N_6140);
and U6912 (N_6912,N_6518,N_6506);
xor U6913 (N_6913,N_6256,N_6567);
nand U6914 (N_6914,N_6212,N_6355);
nor U6915 (N_6915,N_6048,N_6095);
xor U6916 (N_6916,N_6475,N_6595);
xor U6917 (N_6917,N_6086,N_6539);
xor U6918 (N_6918,N_6007,N_6070);
xnor U6919 (N_6919,N_6101,N_6182);
and U6920 (N_6920,N_6392,N_6332);
nand U6921 (N_6921,N_6029,N_6181);
nor U6922 (N_6922,N_6226,N_6545);
or U6923 (N_6923,N_6196,N_6033);
nor U6924 (N_6924,N_6385,N_6447);
and U6925 (N_6925,N_6345,N_6363);
and U6926 (N_6926,N_6217,N_6487);
and U6927 (N_6927,N_6565,N_6083);
and U6928 (N_6928,N_6537,N_6011);
and U6929 (N_6929,N_6306,N_6521);
nor U6930 (N_6930,N_6061,N_6183);
nor U6931 (N_6931,N_6538,N_6045);
nand U6932 (N_6932,N_6463,N_6181);
nor U6933 (N_6933,N_6237,N_6231);
nor U6934 (N_6934,N_6325,N_6467);
and U6935 (N_6935,N_6077,N_6331);
or U6936 (N_6936,N_6153,N_6151);
nor U6937 (N_6937,N_6215,N_6041);
nor U6938 (N_6938,N_6134,N_6396);
nor U6939 (N_6939,N_6465,N_6362);
and U6940 (N_6940,N_6134,N_6306);
or U6941 (N_6941,N_6265,N_6518);
xor U6942 (N_6942,N_6412,N_6472);
xor U6943 (N_6943,N_6507,N_6141);
xnor U6944 (N_6944,N_6470,N_6453);
xnor U6945 (N_6945,N_6048,N_6360);
and U6946 (N_6946,N_6500,N_6511);
or U6947 (N_6947,N_6097,N_6421);
and U6948 (N_6948,N_6288,N_6193);
nor U6949 (N_6949,N_6363,N_6357);
nor U6950 (N_6950,N_6348,N_6458);
nor U6951 (N_6951,N_6267,N_6373);
xor U6952 (N_6952,N_6172,N_6380);
nor U6953 (N_6953,N_6049,N_6307);
nand U6954 (N_6954,N_6292,N_6480);
and U6955 (N_6955,N_6079,N_6250);
nor U6956 (N_6956,N_6479,N_6214);
and U6957 (N_6957,N_6310,N_6053);
or U6958 (N_6958,N_6164,N_6566);
nor U6959 (N_6959,N_6190,N_6005);
or U6960 (N_6960,N_6440,N_6092);
or U6961 (N_6961,N_6552,N_6010);
or U6962 (N_6962,N_6017,N_6271);
nor U6963 (N_6963,N_6118,N_6577);
nand U6964 (N_6964,N_6596,N_6278);
or U6965 (N_6965,N_6021,N_6422);
or U6966 (N_6966,N_6151,N_6562);
and U6967 (N_6967,N_6087,N_6079);
nor U6968 (N_6968,N_6590,N_6331);
or U6969 (N_6969,N_6215,N_6092);
xor U6970 (N_6970,N_6367,N_6388);
xnor U6971 (N_6971,N_6456,N_6090);
nor U6972 (N_6972,N_6079,N_6364);
nand U6973 (N_6973,N_6473,N_6288);
xnor U6974 (N_6974,N_6164,N_6528);
or U6975 (N_6975,N_6096,N_6082);
xnor U6976 (N_6976,N_6433,N_6582);
xor U6977 (N_6977,N_6014,N_6178);
and U6978 (N_6978,N_6310,N_6509);
or U6979 (N_6979,N_6141,N_6240);
nand U6980 (N_6980,N_6127,N_6599);
or U6981 (N_6981,N_6078,N_6251);
xor U6982 (N_6982,N_6363,N_6278);
nor U6983 (N_6983,N_6545,N_6523);
or U6984 (N_6984,N_6191,N_6520);
xor U6985 (N_6985,N_6056,N_6401);
xnor U6986 (N_6986,N_6158,N_6415);
nand U6987 (N_6987,N_6490,N_6204);
xnor U6988 (N_6988,N_6182,N_6217);
nand U6989 (N_6989,N_6534,N_6526);
and U6990 (N_6990,N_6096,N_6121);
nor U6991 (N_6991,N_6085,N_6183);
nor U6992 (N_6992,N_6067,N_6020);
nand U6993 (N_6993,N_6443,N_6115);
and U6994 (N_6994,N_6369,N_6215);
nand U6995 (N_6995,N_6332,N_6406);
and U6996 (N_6996,N_6135,N_6061);
or U6997 (N_6997,N_6281,N_6027);
and U6998 (N_6998,N_6038,N_6141);
xnor U6999 (N_6999,N_6304,N_6283);
xor U7000 (N_7000,N_6594,N_6255);
xor U7001 (N_7001,N_6491,N_6548);
xor U7002 (N_7002,N_6132,N_6124);
xor U7003 (N_7003,N_6576,N_6398);
nand U7004 (N_7004,N_6569,N_6139);
nor U7005 (N_7005,N_6249,N_6103);
xnor U7006 (N_7006,N_6579,N_6355);
and U7007 (N_7007,N_6471,N_6069);
or U7008 (N_7008,N_6237,N_6316);
nor U7009 (N_7009,N_6369,N_6134);
nor U7010 (N_7010,N_6016,N_6396);
and U7011 (N_7011,N_6180,N_6190);
xor U7012 (N_7012,N_6032,N_6174);
nand U7013 (N_7013,N_6460,N_6391);
xnor U7014 (N_7014,N_6291,N_6219);
nand U7015 (N_7015,N_6252,N_6536);
nand U7016 (N_7016,N_6110,N_6367);
nor U7017 (N_7017,N_6519,N_6130);
nand U7018 (N_7018,N_6353,N_6287);
xnor U7019 (N_7019,N_6575,N_6052);
nand U7020 (N_7020,N_6256,N_6351);
and U7021 (N_7021,N_6295,N_6357);
xnor U7022 (N_7022,N_6488,N_6175);
nor U7023 (N_7023,N_6198,N_6163);
nand U7024 (N_7024,N_6504,N_6034);
and U7025 (N_7025,N_6235,N_6593);
or U7026 (N_7026,N_6514,N_6504);
nand U7027 (N_7027,N_6411,N_6343);
and U7028 (N_7028,N_6550,N_6067);
or U7029 (N_7029,N_6277,N_6101);
or U7030 (N_7030,N_6452,N_6283);
and U7031 (N_7031,N_6413,N_6486);
and U7032 (N_7032,N_6428,N_6209);
nand U7033 (N_7033,N_6214,N_6379);
nand U7034 (N_7034,N_6212,N_6259);
xor U7035 (N_7035,N_6047,N_6515);
or U7036 (N_7036,N_6397,N_6506);
nand U7037 (N_7037,N_6263,N_6497);
xor U7038 (N_7038,N_6278,N_6048);
nor U7039 (N_7039,N_6493,N_6136);
and U7040 (N_7040,N_6548,N_6486);
nor U7041 (N_7041,N_6258,N_6516);
xor U7042 (N_7042,N_6204,N_6148);
nor U7043 (N_7043,N_6057,N_6159);
or U7044 (N_7044,N_6551,N_6283);
and U7045 (N_7045,N_6188,N_6167);
nand U7046 (N_7046,N_6158,N_6305);
and U7047 (N_7047,N_6105,N_6415);
nor U7048 (N_7048,N_6469,N_6330);
nand U7049 (N_7049,N_6425,N_6297);
or U7050 (N_7050,N_6485,N_6133);
nor U7051 (N_7051,N_6352,N_6418);
nand U7052 (N_7052,N_6528,N_6264);
and U7053 (N_7053,N_6278,N_6432);
nor U7054 (N_7054,N_6024,N_6147);
nor U7055 (N_7055,N_6046,N_6563);
nand U7056 (N_7056,N_6058,N_6286);
and U7057 (N_7057,N_6099,N_6033);
xnor U7058 (N_7058,N_6267,N_6463);
nand U7059 (N_7059,N_6110,N_6148);
nand U7060 (N_7060,N_6369,N_6230);
xnor U7061 (N_7061,N_6440,N_6146);
and U7062 (N_7062,N_6045,N_6556);
and U7063 (N_7063,N_6276,N_6572);
nand U7064 (N_7064,N_6284,N_6442);
and U7065 (N_7065,N_6559,N_6094);
nand U7066 (N_7066,N_6413,N_6350);
or U7067 (N_7067,N_6133,N_6050);
nor U7068 (N_7068,N_6297,N_6079);
nor U7069 (N_7069,N_6369,N_6407);
xor U7070 (N_7070,N_6356,N_6496);
xnor U7071 (N_7071,N_6208,N_6562);
and U7072 (N_7072,N_6282,N_6404);
xor U7073 (N_7073,N_6400,N_6166);
and U7074 (N_7074,N_6333,N_6394);
xnor U7075 (N_7075,N_6408,N_6142);
nand U7076 (N_7076,N_6476,N_6193);
nor U7077 (N_7077,N_6094,N_6394);
nor U7078 (N_7078,N_6544,N_6169);
nand U7079 (N_7079,N_6183,N_6117);
and U7080 (N_7080,N_6488,N_6104);
and U7081 (N_7081,N_6274,N_6063);
nand U7082 (N_7082,N_6305,N_6437);
nand U7083 (N_7083,N_6491,N_6280);
nand U7084 (N_7084,N_6567,N_6420);
and U7085 (N_7085,N_6200,N_6581);
nand U7086 (N_7086,N_6385,N_6305);
nand U7087 (N_7087,N_6472,N_6499);
nor U7088 (N_7088,N_6214,N_6216);
and U7089 (N_7089,N_6386,N_6168);
xor U7090 (N_7090,N_6006,N_6211);
or U7091 (N_7091,N_6540,N_6010);
or U7092 (N_7092,N_6282,N_6114);
xor U7093 (N_7093,N_6244,N_6021);
nor U7094 (N_7094,N_6385,N_6536);
xor U7095 (N_7095,N_6109,N_6389);
nor U7096 (N_7096,N_6366,N_6133);
or U7097 (N_7097,N_6080,N_6273);
and U7098 (N_7098,N_6514,N_6560);
xnor U7099 (N_7099,N_6368,N_6510);
and U7100 (N_7100,N_6223,N_6195);
or U7101 (N_7101,N_6019,N_6298);
nor U7102 (N_7102,N_6078,N_6583);
or U7103 (N_7103,N_6164,N_6284);
nor U7104 (N_7104,N_6109,N_6221);
and U7105 (N_7105,N_6498,N_6561);
nor U7106 (N_7106,N_6598,N_6095);
xor U7107 (N_7107,N_6014,N_6316);
nand U7108 (N_7108,N_6310,N_6152);
nor U7109 (N_7109,N_6386,N_6098);
and U7110 (N_7110,N_6478,N_6076);
nand U7111 (N_7111,N_6115,N_6305);
or U7112 (N_7112,N_6350,N_6394);
xnor U7113 (N_7113,N_6289,N_6166);
xnor U7114 (N_7114,N_6531,N_6523);
nand U7115 (N_7115,N_6459,N_6095);
nor U7116 (N_7116,N_6030,N_6457);
nand U7117 (N_7117,N_6348,N_6153);
or U7118 (N_7118,N_6551,N_6452);
xor U7119 (N_7119,N_6495,N_6166);
xor U7120 (N_7120,N_6061,N_6164);
and U7121 (N_7121,N_6040,N_6238);
and U7122 (N_7122,N_6194,N_6132);
or U7123 (N_7123,N_6596,N_6234);
nand U7124 (N_7124,N_6141,N_6477);
xnor U7125 (N_7125,N_6279,N_6246);
or U7126 (N_7126,N_6560,N_6111);
and U7127 (N_7127,N_6023,N_6017);
xor U7128 (N_7128,N_6451,N_6401);
and U7129 (N_7129,N_6287,N_6572);
xor U7130 (N_7130,N_6140,N_6108);
nand U7131 (N_7131,N_6400,N_6030);
nor U7132 (N_7132,N_6383,N_6009);
nor U7133 (N_7133,N_6112,N_6296);
nor U7134 (N_7134,N_6545,N_6400);
xnor U7135 (N_7135,N_6254,N_6506);
nor U7136 (N_7136,N_6457,N_6458);
or U7137 (N_7137,N_6518,N_6284);
xor U7138 (N_7138,N_6225,N_6576);
nor U7139 (N_7139,N_6568,N_6015);
xor U7140 (N_7140,N_6357,N_6463);
and U7141 (N_7141,N_6063,N_6289);
nor U7142 (N_7142,N_6329,N_6477);
xnor U7143 (N_7143,N_6277,N_6135);
and U7144 (N_7144,N_6183,N_6127);
or U7145 (N_7145,N_6375,N_6128);
nor U7146 (N_7146,N_6295,N_6511);
nor U7147 (N_7147,N_6071,N_6291);
and U7148 (N_7148,N_6161,N_6303);
nor U7149 (N_7149,N_6190,N_6554);
nor U7150 (N_7150,N_6115,N_6005);
and U7151 (N_7151,N_6478,N_6216);
nor U7152 (N_7152,N_6224,N_6241);
nor U7153 (N_7153,N_6000,N_6093);
nor U7154 (N_7154,N_6025,N_6125);
nor U7155 (N_7155,N_6276,N_6024);
nor U7156 (N_7156,N_6559,N_6103);
xnor U7157 (N_7157,N_6574,N_6068);
nor U7158 (N_7158,N_6504,N_6498);
nand U7159 (N_7159,N_6544,N_6219);
nor U7160 (N_7160,N_6164,N_6250);
nand U7161 (N_7161,N_6091,N_6533);
and U7162 (N_7162,N_6243,N_6102);
xnor U7163 (N_7163,N_6336,N_6037);
and U7164 (N_7164,N_6442,N_6164);
or U7165 (N_7165,N_6382,N_6527);
xnor U7166 (N_7166,N_6356,N_6365);
or U7167 (N_7167,N_6166,N_6220);
nand U7168 (N_7168,N_6129,N_6462);
nor U7169 (N_7169,N_6372,N_6470);
xnor U7170 (N_7170,N_6517,N_6401);
xor U7171 (N_7171,N_6199,N_6436);
nor U7172 (N_7172,N_6435,N_6057);
xnor U7173 (N_7173,N_6130,N_6340);
nor U7174 (N_7174,N_6437,N_6428);
nand U7175 (N_7175,N_6052,N_6507);
xnor U7176 (N_7176,N_6318,N_6178);
xor U7177 (N_7177,N_6445,N_6448);
xor U7178 (N_7178,N_6310,N_6565);
nor U7179 (N_7179,N_6473,N_6461);
or U7180 (N_7180,N_6414,N_6089);
and U7181 (N_7181,N_6254,N_6542);
xnor U7182 (N_7182,N_6337,N_6117);
nor U7183 (N_7183,N_6071,N_6459);
nand U7184 (N_7184,N_6134,N_6521);
nor U7185 (N_7185,N_6414,N_6452);
nand U7186 (N_7186,N_6114,N_6536);
nor U7187 (N_7187,N_6006,N_6450);
or U7188 (N_7188,N_6451,N_6257);
and U7189 (N_7189,N_6562,N_6057);
nand U7190 (N_7190,N_6113,N_6222);
nand U7191 (N_7191,N_6244,N_6174);
or U7192 (N_7192,N_6394,N_6530);
nand U7193 (N_7193,N_6309,N_6142);
and U7194 (N_7194,N_6023,N_6564);
or U7195 (N_7195,N_6400,N_6355);
nor U7196 (N_7196,N_6019,N_6335);
and U7197 (N_7197,N_6549,N_6307);
and U7198 (N_7198,N_6551,N_6561);
nor U7199 (N_7199,N_6267,N_6114);
and U7200 (N_7200,N_7131,N_6985);
xor U7201 (N_7201,N_7191,N_6864);
nand U7202 (N_7202,N_6746,N_7162);
nand U7203 (N_7203,N_6900,N_7183);
and U7204 (N_7204,N_7198,N_7072);
or U7205 (N_7205,N_7089,N_6618);
nand U7206 (N_7206,N_7019,N_7090);
nand U7207 (N_7207,N_6696,N_7181);
and U7208 (N_7208,N_7071,N_6806);
nor U7209 (N_7209,N_6736,N_6994);
xor U7210 (N_7210,N_6666,N_6804);
nor U7211 (N_7211,N_7151,N_6945);
or U7212 (N_7212,N_6642,N_7176);
xnor U7213 (N_7213,N_6831,N_7032);
nand U7214 (N_7214,N_6606,N_6894);
and U7215 (N_7215,N_6796,N_6936);
xor U7216 (N_7216,N_6929,N_6837);
and U7217 (N_7217,N_6940,N_6949);
nand U7218 (N_7218,N_7016,N_7056);
and U7219 (N_7219,N_6996,N_6926);
nand U7220 (N_7220,N_6798,N_7004);
nand U7221 (N_7221,N_6711,N_6893);
nor U7222 (N_7222,N_6899,N_7036);
xnor U7223 (N_7223,N_6610,N_7129);
xnor U7224 (N_7224,N_6978,N_7160);
and U7225 (N_7225,N_6673,N_7159);
xnor U7226 (N_7226,N_6629,N_7174);
or U7227 (N_7227,N_7078,N_6719);
and U7228 (N_7228,N_7155,N_7063);
nand U7229 (N_7229,N_7165,N_6924);
xnor U7230 (N_7230,N_6875,N_6975);
xnor U7231 (N_7231,N_6625,N_6971);
xnor U7232 (N_7232,N_6939,N_6944);
xnor U7233 (N_7233,N_7178,N_6675);
xor U7234 (N_7234,N_6664,N_7021);
xor U7235 (N_7235,N_7088,N_7055);
xor U7236 (N_7236,N_7137,N_6777);
nor U7237 (N_7237,N_6890,N_6833);
or U7238 (N_7238,N_7041,N_7157);
and U7239 (N_7239,N_6750,N_6813);
nor U7240 (N_7240,N_6923,N_6827);
nor U7241 (N_7241,N_6756,N_6644);
and U7242 (N_7242,N_7018,N_6886);
nand U7243 (N_7243,N_6704,N_6879);
nand U7244 (N_7244,N_6948,N_6716);
nor U7245 (N_7245,N_6974,N_6999);
or U7246 (N_7246,N_6650,N_6737);
xnor U7247 (N_7247,N_6843,N_6674);
and U7248 (N_7248,N_6793,N_6612);
nor U7249 (N_7249,N_6748,N_7135);
nand U7250 (N_7250,N_7096,N_6742);
xnor U7251 (N_7251,N_7081,N_6867);
and U7252 (N_7252,N_6845,N_6706);
xor U7253 (N_7253,N_7054,N_6604);
or U7254 (N_7254,N_6920,N_6931);
nand U7255 (N_7255,N_7128,N_6934);
xnor U7256 (N_7256,N_7104,N_6714);
xor U7257 (N_7257,N_6871,N_6907);
nor U7258 (N_7258,N_6614,N_7122);
xnor U7259 (N_7259,N_6679,N_6768);
and U7260 (N_7260,N_6870,N_6951);
xnor U7261 (N_7261,N_6849,N_6701);
nand U7262 (N_7262,N_6671,N_7001);
nor U7263 (N_7263,N_6782,N_6964);
nor U7264 (N_7264,N_7098,N_6757);
xor U7265 (N_7265,N_6992,N_7051);
nor U7266 (N_7266,N_6744,N_7103);
nand U7267 (N_7267,N_6928,N_6662);
xor U7268 (N_7268,N_6892,N_6660);
xor U7269 (N_7269,N_6914,N_6967);
or U7270 (N_7270,N_6669,N_6904);
nor U7271 (N_7271,N_6895,N_6630);
and U7272 (N_7272,N_6691,N_6766);
nor U7273 (N_7273,N_6814,N_7085);
or U7274 (N_7274,N_7044,N_6993);
and U7275 (N_7275,N_6792,N_6620);
and U7276 (N_7276,N_6815,N_7168);
nand U7277 (N_7277,N_6910,N_6688);
xnor U7278 (N_7278,N_7076,N_6811);
nor U7279 (N_7279,N_6623,N_6784);
nand U7280 (N_7280,N_7121,N_6639);
or U7281 (N_7281,N_7086,N_6822);
xor U7282 (N_7282,N_6876,N_6624);
or U7283 (N_7283,N_6755,N_6626);
and U7284 (N_7284,N_7099,N_6621);
xor U7285 (N_7285,N_6690,N_7070);
or U7286 (N_7286,N_6887,N_7068);
and U7287 (N_7287,N_7040,N_6725);
and U7288 (N_7288,N_6972,N_6764);
xor U7289 (N_7289,N_7023,N_6747);
or U7290 (N_7290,N_6754,N_6687);
and U7291 (N_7291,N_6726,N_6645);
nand U7292 (N_7292,N_6856,N_6941);
nand U7293 (N_7293,N_7043,N_6731);
and U7294 (N_7294,N_7013,N_6617);
nor U7295 (N_7295,N_6769,N_6773);
xor U7296 (N_7296,N_6795,N_7146);
and U7297 (N_7297,N_6667,N_6863);
nor U7298 (N_7298,N_7189,N_6678);
nand U7299 (N_7299,N_6836,N_6647);
or U7300 (N_7300,N_6869,N_6676);
nand U7301 (N_7301,N_7152,N_6693);
xor U7302 (N_7302,N_6987,N_6763);
or U7303 (N_7303,N_6976,N_7075);
nand U7304 (N_7304,N_6959,N_7084);
and U7305 (N_7305,N_6800,N_7091);
nand U7306 (N_7306,N_6823,N_7062);
nor U7307 (N_7307,N_6973,N_6981);
nor U7308 (N_7308,N_7053,N_6741);
and U7309 (N_7309,N_6652,N_7161);
nor U7310 (N_7310,N_6700,N_7130);
and U7311 (N_7311,N_7117,N_6712);
and U7312 (N_7312,N_6860,N_6616);
nand U7313 (N_7313,N_6848,N_6685);
and U7314 (N_7314,N_6600,N_6854);
xnor U7315 (N_7315,N_6670,N_7185);
xnor U7316 (N_7316,N_6838,N_7102);
xnor U7317 (N_7317,N_6668,N_7143);
nor U7318 (N_7318,N_6657,N_6765);
nor U7319 (N_7319,N_6615,N_7074);
and U7320 (N_7320,N_6906,N_6969);
and U7321 (N_7321,N_6634,N_6966);
nor U7322 (N_7322,N_6715,N_7124);
xor U7323 (N_7323,N_7197,N_7120);
and U7324 (N_7324,N_6780,N_7000);
and U7325 (N_7325,N_6607,N_6859);
or U7326 (N_7326,N_6637,N_6775);
nand U7327 (N_7327,N_6631,N_6877);
nor U7328 (N_7328,N_6774,N_6901);
nor U7329 (N_7329,N_6720,N_6891);
nand U7330 (N_7330,N_6705,N_7025);
nand U7331 (N_7331,N_6850,N_7042);
nor U7332 (N_7332,N_6922,N_7035);
nand U7333 (N_7333,N_6788,N_6828);
or U7334 (N_7334,N_7047,N_7182);
nor U7335 (N_7335,N_7037,N_7186);
and U7336 (N_7336,N_7140,N_7148);
nor U7337 (N_7337,N_6692,N_6703);
nand U7338 (N_7338,N_6799,N_7127);
xnor U7339 (N_7339,N_6842,N_6724);
and U7340 (N_7340,N_7125,N_6957);
and U7341 (N_7341,N_6912,N_6970);
xor U7342 (N_7342,N_6932,N_7010);
and U7343 (N_7343,N_7144,N_6861);
and U7344 (N_7344,N_6834,N_6878);
or U7345 (N_7345,N_6884,N_7009);
xnor U7346 (N_7346,N_7111,N_7106);
and U7347 (N_7347,N_6846,N_7003);
or U7348 (N_7348,N_6649,N_6968);
nor U7349 (N_7349,N_6762,N_6873);
and U7350 (N_7350,N_7017,N_7110);
xor U7351 (N_7351,N_6802,N_6732);
or U7352 (N_7352,N_6868,N_7058);
nor U7353 (N_7353,N_6640,N_6979);
nor U7354 (N_7354,N_7187,N_6633);
nand U7355 (N_7355,N_6882,N_7164);
and U7356 (N_7356,N_7060,N_6865);
and U7357 (N_7357,N_6611,N_6829);
or U7358 (N_7358,N_7142,N_6880);
nor U7359 (N_7359,N_6699,N_7177);
and U7360 (N_7360,N_7015,N_6897);
or U7361 (N_7361,N_7093,N_7138);
nor U7362 (N_7362,N_6952,N_6761);
xor U7363 (N_7363,N_6803,N_6980);
and U7364 (N_7364,N_7119,N_6816);
or U7365 (N_7365,N_7145,N_6619);
xnor U7366 (N_7366,N_7107,N_7079);
and U7367 (N_7367,N_7011,N_6779);
xor U7368 (N_7368,N_7172,N_6909);
and U7369 (N_7369,N_6840,N_7034);
and U7370 (N_7370,N_6648,N_6658);
xnor U7371 (N_7371,N_7014,N_6622);
or U7372 (N_7372,N_7059,N_6603);
and U7373 (N_7373,N_6790,N_7067);
nand U7374 (N_7374,N_6998,N_7024);
nand U7375 (N_7375,N_6821,N_6960);
xnor U7376 (N_7376,N_7083,N_6916);
nand U7377 (N_7377,N_6628,N_6740);
nand U7378 (N_7378,N_6760,N_6683);
xnor U7379 (N_7379,N_6776,N_6759);
xnor U7380 (N_7380,N_6733,N_6807);
nor U7381 (N_7381,N_7190,N_6862);
or U7382 (N_7382,N_7154,N_6866);
nor U7383 (N_7383,N_6778,N_7194);
nor U7384 (N_7384,N_7101,N_6983);
nor U7385 (N_7385,N_6995,N_6723);
nand U7386 (N_7386,N_7109,N_6955);
and U7387 (N_7387,N_6694,N_6824);
and U7388 (N_7388,N_6810,N_6632);
nor U7389 (N_7389,N_6708,N_7147);
xnor U7390 (N_7390,N_6682,N_6908);
nor U7391 (N_7391,N_6707,N_7087);
nor U7392 (N_7392,N_7126,N_6681);
xnor U7393 (N_7393,N_6989,N_7180);
nor U7394 (N_7394,N_7082,N_6772);
nand U7395 (N_7395,N_6977,N_6935);
or U7396 (N_7396,N_7045,N_7171);
xnor U7397 (N_7397,N_6727,N_7193);
xnor U7398 (N_7398,N_7153,N_6677);
nand U7399 (N_7399,N_6832,N_7114);
and U7400 (N_7400,N_7112,N_6656);
xnor U7401 (N_7401,N_6709,N_7195);
xnor U7402 (N_7402,N_6697,N_6913);
xor U7403 (N_7403,N_7052,N_7169);
and U7404 (N_7404,N_7095,N_6608);
and U7405 (N_7405,N_6686,N_7057);
xor U7406 (N_7406,N_6787,N_6605);
and U7407 (N_7407,N_7100,N_7158);
or U7408 (N_7408,N_6627,N_7026);
and U7409 (N_7409,N_7134,N_6735);
and U7410 (N_7410,N_7027,N_6954);
or U7411 (N_7411,N_7139,N_7028);
nand U7412 (N_7412,N_7033,N_6874);
or U7413 (N_7413,N_7179,N_6881);
and U7414 (N_7414,N_6830,N_7192);
nor U7415 (N_7415,N_6729,N_6857);
and U7416 (N_7416,N_6918,N_6930);
or U7417 (N_7417,N_6942,N_6958);
xnor U7418 (N_7418,N_6752,N_6982);
or U7419 (N_7419,N_7065,N_7029);
and U7420 (N_7420,N_7066,N_6641);
or U7421 (N_7421,N_6767,N_7039);
nand U7422 (N_7422,N_7048,N_7108);
nand U7423 (N_7423,N_7156,N_6730);
xor U7424 (N_7424,N_6927,N_7097);
nand U7425 (N_7425,N_6783,N_6943);
and U7426 (N_7426,N_6638,N_6825);
or U7427 (N_7427,N_6808,N_6990);
or U7428 (N_7428,N_6885,N_6728);
nand U7429 (N_7429,N_7030,N_7163);
xor U7430 (N_7430,N_6841,N_7116);
and U7431 (N_7431,N_6911,N_6710);
nand U7432 (N_7432,N_7002,N_7199);
xnor U7433 (N_7433,N_7005,N_6722);
nor U7434 (N_7434,N_6739,N_6684);
nand U7435 (N_7435,N_7049,N_7077);
or U7436 (N_7436,N_6801,N_6791);
nor U7437 (N_7437,N_7012,N_6771);
or U7438 (N_7438,N_6902,N_6663);
and U7439 (N_7439,N_6986,N_6937);
nand U7440 (N_7440,N_6809,N_7118);
and U7441 (N_7441,N_7080,N_6855);
or U7442 (N_7442,N_6672,N_7136);
nand U7443 (N_7443,N_6609,N_6839);
xnor U7444 (N_7444,N_6938,N_7022);
xor U7445 (N_7445,N_6898,N_6786);
nand U7446 (N_7446,N_6915,N_6858);
xor U7447 (N_7447,N_6853,N_6651);
xor U7448 (N_7448,N_6933,N_7061);
or U7449 (N_7449,N_6770,N_7031);
or U7450 (N_7450,N_6646,N_6602);
or U7451 (N_7451,N_6655,N_7167);
nand U7452 (N_7452,N_6794,N_6785);
or U7453 (N_7453,N_7105,N_6956);
nor U7454 (N_7454,N_6665,N_6889);
nor U7455 (N_7455,N_6601,N_7149);
and U7456 (N_7456,N_6718,N_6872);
nand U7457 (N_7457,N_6888,N_6851);
and U7458 (N_7458,N_6820,N_6961);
nor U7459 (N_7459,N_6689,N_7020);
nand U7460 (N_7460,N_7123,N_6988);
and U7461 (N_7461,N_7133,N_7069);
or U7462 (N_7462,N_6698,N_6984);
nor U7463 (N_7463,N_7038,N_6852);
nand U7464 (N_7464,N_6734,N_6738);
nand U7465 (N_7465,N_6947,N_6844);
nor U7466 (N_7466,N_6817,N_7150);
and U7467 (N_7467,N_6653,N_6745);
nand U7468 (N_7468,N_6805,N_7196);
xor U7469 (N_7469,N_7170,N_7008);
and U7470 (N_7470,N_6643,N_6917);
xor U7471 (N_7471,N_7166,N_7132);
xor U7472 (N_7472,N_6654,N_6753);
nor U7473 (N_7473,N_6758,N_6905);
nor U7474 (N_7474,N_6812,N_6695);
nand U7475 (N_7475,N_7050,N_7113);
nand U7476 (N_7476,N_7092,N_7073);
or U7477 (N_7477,N_6721,N_6636);
nor U7478 (N_7478,N_6883,N_6896);
or U7479 (N_7479,N_6835,N_6789);
nor U7480 (N_7480,N_6903,N_6826);
or U7481 (N_7481,N_6659,N_6921);
nor U7482 (N_7482,N_6991,N_7007);
nor U7483 (N_7483,N_6749,N_6661);
or U7484 (N_7484,N_6847,N_6925);
nor U7485 (N_7485,N_6702,N_6743);
nand U7486 (N_7486,N_7141,N_6797);
xor U7487 (N_7487,N_6751,N_7173);
nand U7488 (N_7488,N_6950,N_7184);
or U7489 (N_7489,N_7175,N_6819);
nand U7490 (N_7490,N_6997,N_6713);
nand U7491 (N_7491,N_6946,N_6680);
nor U7492 (N_7492,N_7115,N_6613);
and U7493 (N_7493,N_6963,N_6818);
and U7494 (N_7494,N_6635,N_6953);
nor U7495 (N_7495,N_6781,N_7094);
or U7496 (N_7496,N_6717,N_7006);
nor U7497 (N_7497,N_6965,N_7046);
nor U7498 (N_7498,N_7188,N_6962);
and U7499 (N_7499,N_7064,N_6919);
or U7500 (N_7500,N_6931,N_6939);
xnor U7501 (N_7501,N_6954,N_6838);
or U7502 (N_7502,N_6915,N_6983);
or U7503 (N_7503,N_6663,N_6722);
and U7504 (N_7504,N_6698,N_6682);
xnor U7505 (N_7505,N_7181,N_6742);
nor U7506 (N_7506,N_7030,N_7003);
and U7507 (N_7507,N_6873,N_7074);
xnor U7508 (N_7508,N_7113,N_6671);
or U7509 (N_7509,N_6728,N_6840);
or U7510 (N_7510,N_6662,N_7181);
xnor U7511 (N_7511,N_6929,N_6875);
nor U7512 (N_7512,N_6977,N_7072);
nor U7513 (N_7513,N_7059,N_6637);
and U7514 (N_7514,N_7169,N_6883);
or U7515 (N_7515,N_6776,N_6639);
or U7516 (N_7516,N_7179,N_6862);
and U7517 (N_7517,N_7066,N_6703);
nand U7518 (N_7518,N_6729,N_6695);
or U7519 (N_7519,N_6697,N_7011);
xnor U7520 (N_7520,N_6838,N_6782);
nor U7521 (N_7521,N_7144,N_6883);
or U7522 (N_7522,N_6880,N_7021);
nand U7523 (N_7523,N_6790,N_7082);
nor U7524 (N_7524,N_6641,N_7024);
xnor U7525 (N_7525,N_7018,N_6600);
nand U7526 (N_7526,N_7012,N_7162);
nor U7527 (N_7527,N_6791,N_6974);
xnor U7528 (N_7528,N_7129,N_7041);
or U7529 (N_7529,N_6958,N_7119);
nand U7530 (N_7530,N_6926,N_6652);
nand U7531 (N_7531,N_7044,N_7104);
xnor U7532 (N_7532,N_6855,N_7142);
nand U7533 (N_7533,N_6855,N_7106);
nand U7534 (N_7534,N_6658,N_6799);
nand U7535 (N_7535,N_6955,N_6642);
xnor U7536 (N_7536,N_7012,N_6819);
and U7537 (N_7537,N_6600,N_6753);
xnor U7538 (N_7538,N_6985,N_7182);
xnor U7539 (N_7539,N_7028,N_6689);
and U7540 (N_7540,N_6920,N_7111);
nor U7541 (N_7541,N_6886,N_7077);
and U7542 (N_7542,N_6688,N_6622);
xor U7543 (N_7543,N_7095,N_6775);
or U7544 (N_7544,N_6894,N_6987);
or U7545 (N_7545,N_6790,N_6848);
xnor U7546 (N_7546,N_6709,N_6827);
and U7547 (N_7547,N_6953,N_7146);
or U7548 (N_7548,N_7143,N_7132);
and U7549 (N_7549,N_6983,N_6754);
or U7550 (N_7550,N_6916,N_6665);
xor U7551 (N_7551,N_7023,N_7115);
and U7552 (N_7552,N_6819,N_7068);
and U7553 (N_7553,N_7085,N_6826);
nand U7554 (N_7554,N_6773,N_6929);
nand U7555 (N_7555,N_6702,N_6987);
nor U7556 (N_7556,N_7107,N_6761);
or U7557 (N_7557,N_6611,N_6963);
or U7558 (N_7558,N_6859,N_7076);
or U7559 (N_7559,N_6767,N_7152);
nor U7560 (N_7560,N_6665,N_6606);
or U7561 (N_7561,N_6807,N_6631);
xor U7562 (N_7562,N_7049,N_6869);
and U7563 (N_7563,N_6679,N_6802);
or U7564 (N_7564,N_6834,N_7123);
nand U7565 (N_7565,N_6803,N_7174);
nand U7566 (N_7566,N_6699,N_6803);
nor U7567 (N_7567,N_7184,N_7029);
nand U7568 (N_7568,N_6876,N_6804);
or U7569 (N_7569,N_6829,N_7131);
nand U7570 (N_7570,N_6639,N_6688);
and U7571 (N_7571,N_6855,N_6955);
and U7572 (N_7572,N_7184,N_6622);
and U7573 (N_7573,N_6923,N_6887);
xnor U7574 (N_7574,N_7026,N_6979);
nand U7575 (N_7575,N_6634,N_6889);
nor U7576 (N_7576,N_7113,N_7098);
or U7577 (N_7577,N_6824,N_6629);
or U7578 (N_7578,N_7034,N_6893);
or U7579 (N_7579,N_6659,N_6600);
xnor U7580 (N_7580,N_6934,N_6601);
nand U7581 (N_7581,N_6808,N_6938);
xor U7582 (N_7582,N_7169,N_7093);
nor U7583 (N_7583,N_7047,N_6969);
xor U7584 (N_7584,N_6856,N_7056);
nand U7585 (N_7585,N_6740,N_7061);
xnor U7586 (N_7586,N_6654,N_7118);
nand U7587 (N_7587,N_6726,N_7056);
or U7588 (N_7588,N_6891,N_6758);
nor U7589 (N_7589,N_6795,N_6766);
nand U7590 (N_7590,N_7096,N_7175);
nor U7591 (N_7591,N_6932,N_6692);
nand U7592 (N_7592,N_7153,N_6969);
and U7593 (N_7593,N_7142,N_6942);
nand U7594 (N_7594,N_6916,N_6896);
or U7595 (N_7595,N_7082,N_6825);
xor U7596 (N_7596,N_6967,N_6872);
nor U7597 (N_7597,N_6718,N_7089);
xor U7598 (N_7598,N_7197,N_7094);
or U7599 (N_7599,N_7148,N_7172);
nor U7600 (N_7600,N_6603,N_7156);
nor U7601 (N_7601,N_6862,N_6688);
and U7602 (N_7602,N_6633,N_7069);
and U7603 (N_7603,N_6970,N_6681);
nand U7604 (N_7604,N_6673,N_6668);
nand U7605 (N_7605,N_6855,N_6643);
nor U7606 (N_7606,N_6680,N_6983);
nand U7607 (N_7607,N_6927,N_6966);
and U7608 (N_7608,N_6750,N_6883);
nand U7609 (N_7609,N_6766,N_6986);
and U7610 (N_7610,N_6772,N_7180);
and U7611 (N_7611,N_6853,N_7031);
nand U7612 (N_7612,N_6826,N_6794);
or U7613 (N_7613,N_7125,N_6825);
or U7614 (N_7614,N_6817,N_6727);
nor U7615 (N_7615,N_6741,N_7030);
nor U7616 (N_7616,N_7154,N_7179);
nand U7617 (N_7617,N_7014,N_6874);
or U7618 (N_7618,N_6872,N_6865);
and U7619 (N_7619,N_6951,N_6999);
xor U7620 (N_7620,N_6786,N_6944);
and U7621 (N_7621,N_7109,N_6787);
and U7622 (N_7622,N_6857,N_7096);
nand U7623 (N_7623,N_7085,N_7087);
xnor U7624 (N_7624,N_7022,N_7145);
or U7625 (N_7625,N_7119,N_6721);
nor U7626 (N_7626,N_6995,N_7035);
nand U7627 (N_7627,N_6947,N_6662);
and U7628 (N_7628,N_6963,N_6823);
or U7629 (N_7629,N_6853,N_7028);
or U7630 (N_7630,N_6987,N_6789);
nor U7631 (N_7631,N_6786,N_6781);
and U7632 (N_7632,N_6661,N_7130);
nor U7633 (N_7633,N_7027,N_6783);
nor U7634 (N_7634,N_6890,N_6612);
and U7635 (N_7635,N_6746,N_7007);
nor U7636 (N_7636,N_6987,N_6881);
nand U7637 (N_7637,N_6752,N_6755);
xnor U7638 (N_7638,N_7108,N_6843);
nor U7639 (N_7639,N_7102,N_7132);
and U7640 (N_7640,N_6840,N_6926);
nand U7641 (N_7641,N_6942,N_6793);
xor U7642 (N_7642,N_7018,N_6865);
or U7643 (N_7643,N_7182,N_6704);
nor U7644 (N_7644,N_7184,N_7137);
nor U7645 (N_7645,N_6927,N_7143);
or U7646 (N_7646,N_7140,N_7150);
and U7647 (N_7647,N_7043,N_6953);
nor U7648 (N_7648,N_6842,N_6746);
or U7649 (N_7649,N_6736,N_6831);
or U7650 (N_7650,N_6647,N_6873);
and U7651 (N_7651,N_7198,N_6846);
nor U7652 (N_7652,N_6910,N_7061);
nor U7653 (N_7653,N_6998,N_6794);
nor U7654 (N_7654,N_6880,N_6976);
xnor U7655 (N_7655,N_7167,N_6610);
xnor U7656 (N_7656,N_7136,N_6624);
and U7657 (N_7657,N_7105,N_6942);
or U7658 (N_7658,N_7180,N_7132);
nor U7659 (N_7659,N_7195,N_7161);
nand U7660 (N_7660,N_6849,N_7010);
nor U7661 (N_7661,N_6659,N_7075);
nor U7662 (N_7662,N_6919,N_7124);
nor U7663 (N_7663,N_6717,N_7167);
or U7664 (N_7664,N_6752,N_6694);
xnor U7665 (N_7665,N_6913,N_7012);
nand U7666 (N_7666,N_6696,N_6645);
and U7667 (N_7667,N_6851,N_7134);
or U7668 (N_7668,N_6930,N_6968);
nor U7669 (N_7669,N_7034,N_7142);
xnor U7670 (N_7670,N_6731,N_6946);
nand U7671 (N_7671,N_7017,N_6614);
xnor U7672 (N_7672,N_6691,N_6888);
xor U7673 (N_7673,N_7082,N_6736);
or U7674 (N_7674,N_7077,N_7093);
or U7675 (N_7675,N_7024,N_7065);
xnor U7676 (N_7676,N_7107,N_6762);
nor U7677 (N_7677,N_6843,N_7156);
or U7678 (N_7678,N_6845,N_7080);
nor U7679 (N_7679,N_7133,N_6687);
and U7680 (N_7680,N_6762,N_6704);
xnor U7681 (N_7681,N_6775,N_7071);
xnor U7682 (N_7682,N_6752,N_6833);
nor U7683 (N_7683,N_6868,N_7165);
or U7684 (N_7684,N_6601,N_6709);
xor U7685 (N_7685,N_6846,N_6923);
xor U7686 (N_7686,N_6851,N_6741);
xnor U7687 (N_7687,N_6792,N_6710);
nand U7688 (N_7688,N_7116,N_6877);
or U7689 (N_7689,N_7042,N_7105);
nand U7690 (N_7690,N_6654,N_7001);
nand U7691 (N_7691,N_6783,N_7155);
and U7692 (N_7692,N_7026,N_6965);
or U7693 (N_7693,N_7173,N_6756);
nand U7694 (N_7694,N_7164,N_6898);
and U7695 (N_7695,N_7163,N_6642);
xor U7696 (N_7696,N_7104,N_6605);
xnor U7697 (N_7697,N_6862,N_6993);
nor U7698 (N_7698,N_7012,N_7141);
nand U7699 (N_7699,N_6675,N_6952);
and U7700 (N_7700,N_6774,N_6618);
nor U7701 (N_7701,N_7021,N_6688);
or U7702 (N_7702,N_6968,N_6742);
and U7703 (N_7703,N_7155,N_6776);
nor U7704 (N_7704,N_7191,N_6660);
or U7705 (N_7705,N_6787,N_7098);
and U7706 (N_7706,N_6759,N_7036);
or U7707 (N_7707,N_6992,N_7021);
nor U7708 (N_7708,N_6961,N_6647);
nor U7709 (N_7709,N_6907,N_6987);
nor U7710 (N_7710,N_7121,N_7006);
and U7711 (N_7711,N_7045,N_6728);
and U7712 (N_7712,N_7047,N_6632);
nor U7713 (N_7713,N_6951,N_6819);
and U7714 (N_7714,N_7005,N_6639);
and U7715 (N_7715,N_7060,N_6665);
xor U7716 (N_7716,N_6657,N_6679);
and U7717 (N_7717,N_7145,N_6867);
xnor U7718 (N_7718,N_6603,N_7032);
xnor U7719 (N_7719,N_6938,N_7085);
or U7720 (N_7720,N_7046,N_6966);
or U7721 (N_7721,N_7109,N_7188);
nor U7722 (N_7722,N_6690,N_6842);
nor U7723 (N_7723,N_7030,N_7076);
nand U7724 (N_7724,N_6810,N_6613);
xor U7725 (N_7725,N_6801,N_6968);
and U7726 (N_7726,N_6628,N_6897);
and U7727 (N_7727,N_6898,N_7079);
nor U7728 (N_7728,N_6690,N_6874);
nor U7729 (N_7729,N_7085,N_6740);
or U7730 (N_7730,N_7178,N_6976);
nor U7731 (N_7731,N_7066,N_7037);
xor U7732 (N_7732,N_6810,N_6673);
nand U7733 (N_7733,N_6888,N_6749);
or U7734 (N_7734,N_6655,N_6972);
nor U7735 (N_7735,N_7172,N_6688);
nor U7736 (N_7736,N_7046,N_6754);
and U7737 (N_7737,N_6716,N_6680);
nand U7738 (N_7738,N_7172,N_7051);
nand U7739 (N_7739,N_6884,N_6740);
and U7740 (N_7740,N_6885,N_6749);
nand U7741 (N_7741,N_6626,N_6758);
nor U7742 (N_7742,N_6758,N_6634);
nor U7743 (N_7743,N_6610,N_6675);
nor U7744 (N_7744,N_6615,N_7104);
or U7745 (N_7745,N_6797,N_6891);
nand U7746 (N_7746,N_7115,N_6814);
or U7747 (N_7747,N_7162,N_6747);
or U7748 (N_7748,N_6825,N_7076);
and U7749 (N_7749,N_7019,N_6817);
and U7750 (N_7750,N_6861,N_7045);
xnor U7751 (N_7751,N_6767,N_7033);
nand U7752 (N_7752,N_6620,N_6982);
and U7753 (N_7753,N_7137,N_7097);
nand U7754 (N_7754,N_6778,N_6840);
nor U7755 (N_7755,N_7188,N_7040);
or U7756 (N_7756,N_6805,N_6734);
or U7757 (N_7757,N_6738,N_6815);
nor U7758 (N_7758,N_6986,N_7139);
and U7759 (N_7759,N_6642,N_7027);
nand U7760 (N_7760,N_6827,N_6996);
nor U7761 (N_7761,N_6855,N_6900);
and U7762 (N_7762,N_6881,N_6638);
or U7763 (N_7763,N_6940,N_6751);
xor U7764 (N_7764,N_6954,N_6963);
and U7765 (N_7765,N_6746,N_6890);
xor U7766 (N_7766,N_7036,N_7021);
or U7767 (N_7767,N_6953,N_6828);
nor U7768 (N_7768,N_6906,N_7141);
or U7769 (N_7769,N_7127,N_6989);
nor U7770 (N_7770,N_7033,N_6625);
xor U7771 (N_7771,N_6630,N_6887);
nor U7772 (N_7772,N_6757,N_6802);
xnor U7773 (N_7773,N_6845,N_6983);
nor U7774 (N_7774,N_7084,N_6678);
nor U7775 (N_7775,N_6930,N_6804);
nand U7776 (N_7776,N_7021,N_6713);
nor U7777 (N_7777,N_6782,N_7179);
or U7778 (N_7778,N_6874,N_6652);
nor U7779 (N_7779,N_6686,N_6667);
xor U7780 (N_7780,N_7018,N_6753);
or U7781 (N_7781,N_6734,N_6712);
or U7782 (N_7782,N_7116,N_7157);
and U7783 (N_7783,N_6810,N_6941);
and U7784 (N_7784,N_6702,N_6718);
nand U7785 (N_7785,N_7090,N_6777);
nor U7786 (N_7786,N_6875,N_6928);
or U7787 (N_7787,N_6892,N_7075);
nor U7788 (N_7788,N_7048,N_6970);
nand U7789 (N_7789,N_6770,N_6977);
or U7790 (N_7790,N_6920,N_6902);
or U7791 (N_7791,N_6628,N_6914);
nand U7792 (N_7792,N_7155,N_7136);
xnor U7793 (N_7793,N_6766,N_6952);
nor U7794 (N_7794,N_6877,N_6601);
xor U7795 (N_7795,N_6983,N_6957);
or U7796 (N_7796,N_6817,N_6655);
nand U7797 (N_7797,N_6635,N_6863);
nor U7798 (N_7798,N_6874,N_6806);
or U7799 (N_7799,N_6928,N_6641);
xnor U7800 (N_7800,N_7463,N_7406);
xor U7801 (N_7801,N_7695,N_7632);
nand U7802 (N_7802,N_7210,N_7236);
nor U7803 (N_7803,N_7470,N_7542);
nor U7804 (N_7804,N_7601,N_7397);
nor U7805 (N_7805,N_7453,N_7574);
or U7806 (N_7806,N_7740,N_7402);
or U7807 (N_7807,N_7264,N_7640);
or U7808 (N_7808,N_7338,N_7727);
xor U7809 (N_7809,N_7459,N_7745);
nor U7810 (N_7810,N_7238,N_7228);
nand U7811 (N_7811,N_7723,N_7529);
nor U7812 (N_7812,N_7625,N_7431);
xor U7813 (N_7813,N_7499,N_7478);
nor U7814 (N_7814,N_7505,N_7708);
and U7815 (N_7815,N_7462,N_7337);
or U7816 (N_7816,N_7648,N_7317);
and U7817 (N_7817,N_7654,N_7369);
or U7818 (N_7818,N_7293,N_7415);
or U7819 (N_7819,N_7646,N_7536);
nor U7820 (N_7820,N_7231,N_7675);
or U7821 (N_7821,N_7700,N_7329);
nand U7822 (N_7822,N_7628,N_7656);
nand U7823 (N_7823,N_7241,N_7440);
or U7824 (N_7824,N_7750,N_7299);
and U7825 (N_7825,N_7331,N_7558);
xnor U7826 (N_7826,N_7732,N_7355);
nand U7827 (N_7827,N_7497,N_7667);
nor U7828 (N_7828,N_7596,N_7328);
xor U7829 (N_7829,N_7682,N_7502);
nor U7830 (N_7830,N_7491,N_7658);
xnor U7831 (N_7831,N_7666,N_7799);
xnor U7832 (N_7832,N_7468,N_7334);
xor U7833 (N_7833,N_7278,N_7318);
xnor U7834 (N_7834,N_7594,N_7220);
nand U7835 (N_7835,N_7399,N_7386);
nor U7836 (N_7836,N_7736,N_7751);
nand U7837 (N_7837,N_7509,N_7520);
and U7838 (N_7838,N_7531,N_7635);
and U7839 (N_7839,N_7325,N_7322);
nor U7840 (N_7840,N_7511,N_7642);
or U7841 (N_7841,N_7668,N_7219);
nor U7842 (N_7842,N_7370,N_7395);
nand U7843 (N_7843,N_7275,N_7435);
xor U7844 (N_7844,N_7631,N_7758);
nor U7845 (N_7845,N_7494,N_7607);
or U7846 (N_7846,N_7523,N_7327);
and U7847 (N_7847,N_7394,N_7772);
nand U7848 (N_7848,N_7434,N_7613);
or U7849 (N_7849,N_7634,N_7411);
nand U7850 (N_7850,N_7788,N_7243);
nand U7851 (N_7851,N_7721,N_7230);
nor U7852 (N_7852,N_7484,N_7771);
nor U7853 (N_7853,N_7584,N_7432);
nand U7854 (N_7854,N_7202,N_7291);
xor U7855 (N_7855,N_7316,N_7547);
xor U7856 (N_7856,N_7240,N_7333);
nand U7857 (N_7857,N_7413,N_7624);
or U7858 (N_7858,N_7617,N_7223);
or U7859 (N_7859,N_7754,N_7731);
and U7860 (N_7860,N_7604,N_7599);
xor U7861 (N_7861,N_7266,N_7218);
and U7862 (N_7862,N_7460,N_7650);
nor U7863 (N_7863,N_7439,N_7757);
nand U7864 (N_7864,N_7621,N_7438);
and U7865 (N_7865,N_7669,N_7208);
nor U7866 (N_7866,N_7543,N_7225);
nand U7867 (N_7867,N_7618,N_7786);
or U7868 (N_7868,N_7797,N_7749);
and U7869 (N_7869,N_7733,N_7390);
nor U7870 (N_7870,N_7388,N_7703);
xnor U7871 (N_7871,N_7451,N_7510);
xnor U7872 (N_7872,N_7200,N_7546);
or U7873 (N_7873,N_7756,N_7472);
or U7874 (N_7874,N_7789,N_7259);
nor U7875 (N_7875,N_7466,N_7437);
xnor U7876 (N_7876,N_7215,N_7473);
xnor U7877 (N_7877,N_7591,N_7715);
xnor U7878 (N_7878,N_7759,N_7252);
or U7879 (N_7879,N_7354,N_7344);
nor U7880 (N_7880,N_7777,N_7479);
or U7881 (N_7881,N_7237,N_7716);
or U7882 (N_7882,N_7516,N_7670);
or U7883 (N_7883,N_7792,N_7647);
and U7884 (N_7884,N_7524,N_7576);
or U7885 (N_7885,N_7515,N_7739);
and U7886 (N_7886,N_7489,N_7442);
nand U7887 (N_7887,N_7573,N_7704);
xor U7888 (N_7888,N_7677,N_7540);
xnor U7889 (N_7889,N_7368,N_7269);
nor U7890 (N_7890,N_7420,N_7261);
nor U7891 (N_7891,N_7360,N_7744);
nor U7892 (N_7892,N_7229,N_7752);
xor U7893 (N_7893,N_7726,N_7679);
nand U7894 (N_7894,N_7506,N_7492);
nor U7895 (N_7895,N_7551,N_7633);
nand U7896 (N_7896,N_7405,N_7201);
and U7897 (N_7897,N_7698,N_7794);
or U7898 (N_7898,N_7712,N_7701);
or U7899 (N_7899,N_7268,N_7209);
nor U7900 (N_7900,N_7519,N_7717);
or U7901 (N_7901,N_7769,N_7359);
xnor U7902 (N_7902,N_7694,N_7778);
nand U7903 (N_7903,N_7298,N_7475);
nor U7904 (N_7904,N_7396,N_7222);
nor U7905 (N_7905,N_7637,N_7764);
nor U7906 (N_7906,N_7553,N_7244);
xnor U7907 (N_7907,N_7587,N_7284);
nor U7908 (N_7908,N_7755,N_7371);
or U7909 (N_7909,N_7517,N_7471);
or U7910 (N_7910,N_7363,N_7671);
nor U7911 (N_7911,N_7699,N_7581);
nand U7912 (N_7912,N_7748,N_7426);
or U7913 (N_7913,N_7643,N_7720);
nor U7914 (N_7914,N_7400,N_7541);
nand U7915 (N_7915,N_7290,N_7382);
xor U7916 (N_7916,N_7614,N_7560);
nand U7917 (N_7917,N_7710,N_7310);
nor U7918 (N_7918,N_7486,N_7341);
or U7919 (N_7919,N_7320,N_7790);
nor U7920 (N_7920,N_7455,N_7256);
nor U7921 (N_7921,N_7255,N_7697);
xor U7922 (N_7922,N_7728,N_7645);
and U7923 (N_7923,N_7212,N_7305);
or U7924 (N_7924,N_7608,N_7566);
or U7925 (N_7925,N_7401,N_7738);
nor U7926 (N_7926,N_7730,N_7452);
and U7927 (N_7927,N_7387,N_7655);
xnor U7928 (N_7928,N_7336,N_7367);
and U7929 (N_7929,N_7485,N_7545);
or U7930 (N_7930,N_7454,N_7270);
and U7931 (N_7931,N_7765,N_7693);
xnor U7932 (N_7932,N_7358,N_7595);
and U7933 (N_7933,N_7301,N_7557);
and U7934 (N_7934,N_7476,N_7441);
nor U7935 (N_7935,N_7678,N_7257);
xor U7936 (N_7936,N_7323,N_7611);
xnor U7937 (N_7937,N_7664,N_7378);
xor U7938 (N_7938,N_7652,N_7709);
xnor U7939 (N_7939,N_7606,N_7641);
and U7940 (N_7940,N_7603,N_7780);
nor U7941 (N_7941,N_7307,N_7629);
nand U7942 (N_7942,N_7674,N_7304);
xor U7943 (N_7943,N_7429,N_7271);
or U7944 (N_7944,N_7550,N_7768);
xor U7945 (N_7945,N_7782,N_7385);
and U7946 (N_7946,N_7292,N_7684);
or U7947 (N_7947,N_7559,N_7315);
xnor U7948 (N_7948,N_7504,N_7422);
or U7949 (N_7949,N_7663,N_7722);
nor U7950 (N_7950,N_7417,N_7586);
nor U7951 (N_7951,N_7242,N_7619);
xnor U7952 (N_7952,N_7622,N_7450);
nand U7953 (N_7953,N_7501,N_7224);
and U7954 (N_7954,N_7262,N_7552);
nand U7955 (N_7955,N_7620,N_7421);
and U7956 (N_7956,N_7449,N_7213);
nand U7957 (N_7957,N_7391,N_7308);
xnor U7958 (N_7958,N_7577,N_7623);
xor U7959 (N_7959,N_7234,N_7312);
nor U7960 (N_7960,N_7430,N_7376);
and U7961 (N_7961,N_7570,N_7447);
and U7962 (N_7962,N_7522,N_7313);
nand U7963 (N_7963,N_7326,N_7549);
nand U7964 (N_7964,N_7735,N_7251);
xor U7965 (N_7965,N_7711,N_7427);
nor U7966 (N_7966,N_7548,N_7537);
xor U7967 (N_7967,N_7295,N_7773);
and U7968 (N_7968,N_7458,N_7375);
or U7969 (N_7969,N_7356,N_7630);
nor U7970 (N_7970,N_7366,N_7448);
and U7971 (N_7971,N_7474,N_7638);
or U7972 (N_7972,N_7766,N_7512);
nor U7973 (N_7973,N_7571,N_7791);
nand U7974 (N_7974,N_7651,N_7636);
xnor U7975 (N_7975,N_7514,N_7719);
nand U7976 (N_7976,N_7232,N_7477);
and U7977 (N_7977,N_7518,N_7418);
or U7978 (N_7978,N_7206,N_7364);
and U7979 (N_7979,N_7776,N_7702);
and U7980 (N_7980,N_7384,N_7374);
and U7981 (N_7981,N_7469,N_7285);
xor U7982 (N_7982,N_7443,N_7688);
nand U7983 (N_7983,N_7562,N_7775);
nand U7984 (N_7984,N_7569,N_7428);
and U7985 (N_7985,N_7361,N_7741);
nand U7986 (N_7986,N_7277,N_7692);
or U7987 (N_7987,N_7221,N_7207);
nor U7988 (N_7988,N_7260,N_7481);
xor U7989 (N_7989,N_7249,N_7345);
or U7990 (N_7990,N_7561,N_7350);
xnor U7991 (N_7991,N_7467,N_7311);
or U7992 (N_7992,N_7480,N_7464);
nand U7993 (N_7993,N_7381,N_7565);
or U7994 (N_7994,N_7572,N_7774);
and U7995 (N_7995,N_7233,N_7690);
nand U7996 (N_7996,N_7211,N_7347);
xor U7997 (N_7997,N_7302,N_7245);
xnor U7998 (N_7998,N_7393,N_7685);
or U7999 (N_7999,N_7383,N_7456);
or U8000 (N_8000,N_7483,N_7767);
xnor U8001 (N_8001,N_7681,N_7487);
xnor U8002 (N_8002,N_7598,N_7534);
or U8003 (N_8003,N_7410,N_7653);
and U8004 (N_8004,N_7226,N_7407);
xor U8005 (N_8005,N_7753,N_7339);
nand U8006 (N_8006,N_7253,N_7273);
or U8007 (N_8007,N_7609,N_7589);
xnor U8008 (N_8008,N_7508,N_7414);
and U8009 (N_8009,N_7762,N_7525);
and U8010 (N_8010,N_7662,N_7672);
nand U8011 (N_8011,N_7309,N_7575);
nand U8012 (N_8012,N_7644,N_7507);
xnor U8013 (N_8013,N_7258,N_7239);
nand U8014 (N_8014,N_7707,N_7433);
or U8015 (N_8015,N_7335,N_7683);
xnor U8016 (N_8016,N_7661,N_7539);
and U8017 (N_8017,N_7343,N_7659);
and U8018 (N_8018,N_7392,N_7482);
nand U8019 (N_8019,N_7580,N_7365);
xor U8020 (N_8020,N_7747,N_7706);
nor U8021 (N_8021,N_7605,N_7600);
and U8022 (N_8022,N_7556,N_7665);
or U8023 (N_8023,N_7362,N_7530);
or U8024 (N_8024,N_7490,N_7352);
or U8025 (N_8025,N_7657,N_7289);
xor U8026 (N_8026,N_7349,N_7314);
xnor U8027 (N_8027,N_7513,N_7423);
nand U8028 (N_8028,N_7235,N_7616);
or U8029 (N_8029,N_7424,N_7532);
and U8030 (N_8030,N_7203,N_7602);
and U8031 (N_8031,N_7660,N_7582);
nand U8032 (N_8032,N_7725,N_7588);
xnor U8033 (N_8033,N_7265,N_7246);
nand U8034 (N_8034,N_7680,N_7793);
nand U8035 (N_8035,N_7673,N_7743);
nor U8036 (N_8036,N_7425,N_7446);
nor U8037 (N_8037,N_7639,N_7610);
xor U8038 (N_8038,N_7296,N_7798);
or U8039 (N_8039,N_7205,N_7272);
nand U8040 (N_8040,N_7612,N_7729);
and U8041 (N_8041,N_7297,N_7714);
nor U8042 (N_8042,N_7332,N_7718);
or U8043 (N_8043,N_7250,N_7528);
and U8044 (N_8044,N_7585,N_7465);
and U8045 (N_8045,N_7445,N_7404);
xor U8046 (N_8046,N_7286,N_7303);
or U8047 (N_8047,N_7409,N_7597);
nand U8048 (N_8048,N_7294,N_7526);
xor U8049 (N_8049,N_7554,N_7444);
nand U8050 (N_8050,N_7324,N_7500);
and U8051 (N_8051,N_7351,N_7330);
nand U8052 (N_8052,N_7649,N_7691);
nor U8053 (N_8053,N_7676,N_7254);
and U8054 (N_8054,N_7306,N_7274);
xnor U8055 (N_8055,N_7263,N_7593);
xnor U8056 (N_8056,N_7783,N_7533);
and U8057 (N_8057,N_7781,N_7346);
xnor U8058 (N_8058,N_7555,N_7578);
xnor U8059 (N_8059,N_7267,N_7283);
xnor U8060 (N_8060,N_7784,N_7590);
xnor U8061 (N_8061,N_7770,N_7615);
nor U8062 (N_8062,N_7389,N_7568);
nor U8063 (N_8063,N_7742,N_7288);
xor U8064 (N_8064,N_7538,N_7503);
nand U8065 (N_8065,N_7282,N_7353);
and U8066 (N_8066,N_7705,N_7281);
and U8067 (N_8067,N_7247,N_7687);
and U8068 (N_8068,N_7348,N_7498);
xor U8069 (N_8069,N_7300,N_7217);
xor U8070 (N_8070,N_7248,N_7544);
nor U8071 (N_8071,N_7535,N_7342);
or U8072 (N_8072,N_7795,N_7592);
and U8073 (N_8073,N_7280,N_7321);
nor U8074 (N_8074,N_7493,N_7457);
nor U8075 (N_8075,N_7746,N_7287);
and U8076 (N_8076,N_7357,N_7214);
xor U8077 (N_8077,N_7496,N_7567);
or U8078 (N_8078,N_7488,N_7319);
or U8079 (N_8079,N_7521,N_7216);
xnor U8080 (N_8080,N_7761,N_7563);
or U8081 (N_8081,N_7403,N_7379);
or U8082 (N_8082,N_7279,N_7373);
nand U8083 (N_8083,N_7527,N_7398);
xor U8084 (N_8084,N_7734,N_7416);
nand U8085 (N_8085,N_7696,N_7626);
and U8086 (N_8086,N_7380,N_7419);
or U8087 (N_8087,N_7564,N_7412);
and U8088 (N_8088,N_7796,N_7724);
and U8089 (N_8089,N_7461,N_7686);
xor U8090 (N_8090,N_7787,N_7785);
or U8091 (N_8091,N_7583,N_7779);
and U8092 (N_8092,N_7204,N_7627);
nand U8093 (N_8093,N_7276,N_7760);
or U8094 (N_8094,N_7340,N_7713);
and U8095 (N_8095,N_7737,N_7436);
nor U8096 (N_8096,N_7763,N_7227);
and U8097 (N_8097,N_7372,N_7689);
nor U8098 (N_8098,N_7408,N_7495);
nor U8099 (N_8099,N_7579,N_7377);
or U8100 (N_8100,N_7477,N_7404);
nand U8101 (N_8101,N_7545,N_7389);
or U8102 (N_8102,N_7793,N_7535);
or U8103 (N_8103,N_7638,N_7352);
and U8104 (N_8104,N_7417,N_7763);
xor U8105 (N_8105,N_7787,N_7416);
nand U8106 (N_8106,N_7586,N_7255);
nand U8107 (N_8107,N_7460,N_7611);
nand U8108 (N_8108,N_7611,N_7648);
xor U8109 (N_8109,N_7591,N_7358);
nand U8110 (N_8110,N_7335,N_7501);
nor U8111 (N_8111,N_7656,N_7705);
nor U8112 (N_8112,N_7495,N_7355);
and U8113 (N_8113,N_7591,N_7401);
or U8114 (N_8114,N_7573,N_7744);
or U8115 (N_8115,N_7544,N_7288);
nand U8116 (N_8116,N_7232,N_7294);
or U8117 (N_8117,N_7238,N_7370);
or U8118 (N_8118,N_7745,N_7215);
nor U8119 (N_8119,N_7590,N_7212);
and U8120 (N_8120,N_7294,N_7424);
nor U8121 (N_8121,N_7519,N_7421);
nor U8122 (N_8122,N_7566,N_7219);
nand U8123 (N_8123,N_7706,N_7437);
nand U8124 (N_8124,N_7554,N_7515);
and U8125 (N_8125,N_7682,N_7394);
xor U8126 (N_8126,N_7214,N_7796);
nor U8127 (N_8127,N_7447,N_7317);
and U8128 (N_8128,N_7462,N_7663);
nor U8129 (N_8129,N_7668,N_7277);
and U8130 (N_8130,N_7447,N_7607);
or U8131 (N_8131,N_7667,N_7730);
nand U8132 (N_8132,N_7369,N_7474);
and U8133 (N_8133,N_7572,N_7428);
nor U8134 (N_8134,N_7382,N_7433);
and U8135 (N_8135,N_7270,N_7696);
and U8136 (N_8136,N_7725,N_7234);
or U8137 (N_8137,N_7501,N_7650);
xor U8138 (N_8138,N_7263,N_7502);
nand U8139 (N_8139,N_7619,N_7461);
nand U8140 (N_8140,N_7379,N_7788);
nor U8141 (N_8141,N_7641,N_7629);
xnor U8142 (N_8142,N_7212,N_7414);
xnor U8143 (N_8143,N_7380,N_7703);
or U8144 (N_8144,N_7763,N_7496);
nand U8145 (N_8145,N_7252,N_7406);
or U8146 (N_8146,N_7363,N_7709);
nand U8147 (N_8147,N_7337,N_7583);
xnor U8148 (N_8148,N_7298,N_7440);
nor U8149 (N_8149,N_7776,N_7272);
nand U8150 (N_8150,N_7626,N_7649);
or U8151 (N_8151,N_7335,N_7793);
or U8152 (N_8152,N_7732,N_7675);
nand U8153 (N_8153,N_7213,N_7479);
or U8154 (N_8154,N_7754,N_7725);
nand U8155 (N_8155,N_7485,N_7715);
xor U8156 (N_8156,N_7574,N_7704);
nand U8157 (N_8157,N_7265,N_7469);
or U8158 (N_8158,N_7531,N_7668);
xnor U8159 (N_8159,N_7352,N_7468);
and U8160 (N_8160,N_7527,N_7712);
or U8161 (N_8161,N_7611,N_7741);
xnor U8162 (N_8162,N_7758,N_7302);
and U8163 (N_8163,N_7666,N_7747);
xnor U8164 (N_8164,N_7239,N_7311);
xnor U8165 (N_8165,N_7235,N_7318);
nor U8166 (N_8166,N_7592,N_7340);
and U8167 (N_8167,N_7604,N_7298);
or U8168 (N_8168,N_7578,N_7699);
nor U8169 (N_8169,N_7418,N_7770);
xor U8170 (N_8170,N_7388,N_7722);
nand U8171 (N_8171,N_7751,N_7454);
or U8172 (N_8172,N_7747,N_7248);
nor U8173 (N_8173,N_7375,N_7765);
xor U8174 (N_8174,N_7619,N_7378);
xnor U8175 (N_8175,N_7796,N_7283);
nor U8176 (N_8176,N_7538,N_7508);
nor U8177 (N_8177,N_7229,N_7566);
xnor U8178 (N_8178,N_7296,N_7655);
xnor U8179 (N_8179,N_7636,N_7711);
and U8180 (N_8180,N_7212,N_7556);
or U8181 (N_8181,N_7418,N_7491);
nand U8182 (N_8182,N_7422,N_7627);
or U8183 (N_8183,N_7295,N_7607);
and U8184 (N_8184,N_7778,N_7370);
xnor U8185 (N_8185,N_7650,N_7585);
or U8186 (N_8186,N_7349,N_7556);
nand U8187 (N_8187,N_7553,N_7310);
and U8188 (N_8188,N_7540,N_7773);
nand U8189 (N_8189,N_7711,N_7489);
nor U8190 (N_8190,N_7432,N_7283);
xor U8191 (N_8191,N_7238,N_7799);
or U8192 (N_8192,N_7600,N_7354);
or U8193 (N_8193,N_7696,N_7764);
or U8194 (N_8194,N_7698,N_7527);
nand U8195 (N_8195,N_7467,N_7251);
nand U8196 (N_8196,N_7408,N_7433);
nor U8197 (N_8197,N_7684,N_7578);
nor U8198 (N_8198,N_7318,N_7216);
nand U8199 (N_8199,N_7553,N_7267);
and U8200 (N_8200,N_7497,N_7624);
nand U8201 (N_8201,N_7591,N_7548);
and U8202 (N_8202,N_7364,N_7548);
or U8203 (N_8203,N_7427,N_7441);
and U8204 (N_8204,N_7329,N_7798);
nand U8205 (N_8205,N_7371,N_7721);
xnor U8206 (N_8206,N_7425,N_7666);
and U8207 (N_8207,N_7519,N_7300);
xor U8208 (N_8208,N_7246,N_7224);
xor U8209 (N_8209,N_7717,N_7772);
nor U8210 (N_8210,N_7293,N_7266);
nor U8211 (N_8211,N_7536,N_7501);
nor U8212 (N_8212,N_7780,N_7580);
nor U8213 (N_8213,N_7233,N_7483);
xor U8214 (N_8214,N_7429,N_7502);
xnor U8215 (N_8215,N_7395,N_7302);
or U8216 (N_8216,N_7785,N_7467);
or U8217 (N_8217,N_7597,N_7515);
nand U8218 (N_8218,N_7674,N_7417);
and U8219 (N_8219,N_7753,N_7411);
nor U8220 (N_8220,N_7492,N_7411);
and U8221 (N_8221,N_7751,N_7236);
nand U8222 (N_8222,N_7738,N_7243);
nand U8223 (N_8223,N_7440,N_7588);
and U8224 (N_8224,N_7591,N_7488);
nor U8225 (N_8225,N_7798,N_7209);
nand U8226 (N_8226,N_7479,N_7517);
or U8227 (N_8227,N_7318,N_7759);
and U8228 (N_8228,N_7507,N_7628);
nand U8229 (N_8229,N_7353,N_7400);
and U8230 (N_8230,N_7565,N_7369);
xor U8231 (N_8231,N_7572,N_7532);
and U8232 (N_8232,N_7710,N_7370);
nand U8233 (N_8233,N_7364,N_7355);
or U8234 (N_8234,N_7379,N_7715);
xor U8235 (N_8235,N_7248,N_7242);
and U8236 (N_8236,N_7259,N_7748);
xnor U8237 (N_8237,N_7710,N_7726);
or U8238 (N_8238,N_7263,N_7798);
or U8239 (N_8239,N_7521,N_7562);
nand U8240 (N_8240,N_7626,N_7740);
nand U8241 (N_8241,N_7257,N_7647);
xnor U8242 (N_8242,N_7754,N_7690);
nor U8243 (N_8243,N_7330,N_7365);
nand U8244 (N_8244,N_7315,N_7310);
and U8245 (N_8245,N_7478,N_7743);
nor U8246 (N_8246,N_7242,N_7204);
nand U8247 (N_8247,N_7710,N_7224);
nor U8248 (N_8248,N_7712,N_7314);
and U8249 (N_8249,N_7512,N_7321);
nor U8250 (N_8250,N_7343,N_7386);
or U8251 (N_8251,N_7783,N_7320);
nand U8252 (N_8252,N_7632,N_7278);
and U8253 (N_8253,N_7781,N_7585);
or U8254 (N_8254,N_7506,N_7706);
or U8255 (N_8255,N_7616,N_7443);
nand U8256 (N_8256,N_7371,N_7301);
or U8257 (N_8257,N_7265,N_7639);
nor U8258 (N_8258,N_7646,N_7732);
and U8259 (N_8259,N_7232,N_7773);
xnor U8260 (N_8260,N_7305,N_7760);
or U8261 (N_8261,N_7421,N_7707);
and U8262 (N_8262,N_7685,N_7291);
xor U8263 (N_8263,N_7636,N_7206);
nor U8264 (N_8264,N_7537,N_7586);
and U8265 (N_8265,N_7539,N_7556);
nand U8266 (N_8266,N_7663,N_7733);
xnor U8267 (N_8267,N_7355,N_7453);
xnor U8268 (N_8268,N_7614,N_7457);
and U8269 (N_8269,N_7720,N_7244);
and U8270 (N_8270,N_7293,N_7760);
and U8271 (N_8271,N_7644,N_7208);
nor U8272 (N_8272,N_7356,N_7534);
xnor U8273 (N_8273,N_7395,N_7748);
xor U8274 (N_8274,N_7625,N_7691);
nor U8275 (N_8275,N_7344,N_7460);
xnor U8276 (N_8276,N_7455,N_7467);
nor U8277 (N_8277,N_7221,N_7607);
nand U8278 (N_8278,N_7260,N_7728);
or U8279 (N_8279,N_7537,N_7631);
nand U8280 (N_8280,N_7471,N_7337);
nor U8281 (N_8281,N_7611,N_7257);
nor U8282 (N_8282,N_7595,N_7532);
or U8283 (N_8283,N_7594,N_7583);
or U8284 (N_8284,N_7482,N_7479);
xnor U8285 (N_8285,N_7214,N_7696);
and U8286 (N_8286,N_7794,N_7508);
and U8287 (N_8287,N_7348,N_7306);
or U8288 (N_8288,N_7635,N_7577);
nor U8289 (N_8289,N_7402,N_7349);
or U8290 (N_8290,N_7768,N_7527);
xor U8291 (N_8291,N_7427,N_7370);
and U8292 (N_8292,N_7485,N_7416);
and U8293 (N_8293,N_7292,N_7481);
and U8294 (N_8294,N_7671,N_7254);
or U8295 (N_8295,N_7219,N_7533);
xor U8296 (N_8296,N_7523,N_7322);
nor U8297 (N_8297,N_7229,N_7693);
nand U8298 (N_8298,N_7562,N_7731);
and U8299 (N_8299,N_7629,N_7343);
nor U8300 (N_8300,N_7681,N_7636);
xor U8301 (N_8301,N_7409,N_7712);
nor U8302 (N_8302,N_7680,N_7396);
nand U8303 (N_8303,N_7779,N_7421);
nor U8304 (N_8304,N_7282,N_7792);
xnor U8305 (N_8305,N_7526,N_7365);
nand U8306 (N_8306,N_7429,N_7667);
nand U8307 (N_8307,N_7409,N_7630);
xor U8308 (N_8308,N_7769,N_7412);
xor U8309 (N_8309,N_7213,N_7343);
nor U8310 (N_8310,N_7530,N_7418);
or U8311 (N_8311,N_7707,N_7790);
xor U8312 (N_8312,N_7215,N_7676);
xor U8313 (N_8313,N_7746,N_7728);
xnor U8314 (N_8314,N_7594,N_7634);
nor U8315 (N_8315,N_7309,N_7529);
or U8316 (N_8316,N_7251,N_7232);
or U8317 (N_8317,N_7213,N_7361);
nor U8318 (N_8318,N_7257,N_7435);
xor U8319 (N_8319,N_7482,N_7620);
or U8320 (N_8320,N_7512,N_7477);
nor U8321 (N_8321,N_7601,N_7610);
nor U8322 (N_8322,N_7273,N_7483);
and U8323 (N_8323,N_7293,N_7745);
nor U8324 (N_8324,N_7668,N_7593);
nor U8325 (N_8325,N_7557,N_7575);
and U8326 (N_8326,N_7234,N_7744);
or U8327 (N_8327,N_7604,N_7730);
and U8328 (N_8328,N_7391,N_7434);
xor U8329 (N_8329,N_7495,N_7687);
or U8330 (N_8330,N_7532,N_7207);
and U8331 (N_8331,N_7581,N_7768);
nand U8332 (N_8332,N_7211,N_7622);
xnor U8333 (N_8333,N_7466,N_7223);
or U8334 (N_8334,N_7417,N_7660);
or U8335 (N_8335,N_7728,N_7668);
and U8336 (N_8336,N_7682,N_7791);
nand U8337 (N_8337,N_7701,N_7568);
xnor U8338 (N_8338,N_7652,N_7442);
nor U8339 (N_8339,N_7671,N_7529);
or U8340 (N_8340,N_7559,N_7669);
xnor U8341 (N_8341,N_7434,N_7555);
nor U8342 (N_8342,N_7753,N_7478);
nand U8343 (N_8343,N_7567,N_7288);
and U8344 (N_8344,N_7298,N_7717);
and U8345 (N_8345,N_7367,N_7266);
and U8346 (N_8346,N_7350,N_7201);
or U8347 (N_8347,N_7639,N_7672);
or U8348 (N_8348,N_7703,N_7543);
nor U8349 (N_8349,N_7444,N_7631);
nor U8350 (N_8350,N_7287,N_7255);
or U8351 (N_8351,N_7342,N_7597);
xor U8352 (N_8352,N_7665,N_7286);
and U8353 (N_8353,N_7579,N_7786);
or U8354 (N_8354,N_7767,N_7419);
nor U8355 (N_8355,N_7619,N_7458);
and U8356 (N_8356,N_7363,N_7668);
xor U8357 (N_8357,N_7725,N_7512);
nor U8358 (N_8358,N_7287,N_7321);
nor U8359 (N_8359,N_7723,N_7616);
or U8360 (N_8360,N_7539,N_7475);
nor U8361 (N_8361,N_7603,N_7268);
nor U8362 (N_8362,N_7649,N_7792);
or U8363 (N_8363,N_7441,N_7389);
and U8364 (N_8364,N_7514,N_7247);
or U8365 (N_8365,N_7452,N_7369);
and U8366 (N_8366,N_7554,N_7350);
nor U8367 (N_8367,N_7560,N_7393);
or U8368 (N_8368,N_7321,N_7687);
or U8369 (N_8369,N_7265,N_7508);
xnor U8370 (N_8370,N_7358,N_7516);
nor U8371 (N_8371,N_7482,N_7687);
nand U8372 (N_8372,N_7520,N_7645);
or U8373 (N_8373,N_7637,N_7765);
xnor U8374 (N_8374,N_7392,N_7377);
xnor U8375 (N_8375,N_7536,N_7390);
nand U8376 (N_8376,N_7242,N_7634);
nand U8377 (N_8377,N_7326,N_7603);
and U8378 (N_8378,N_7784,N_7691);
or U8379 (N_8379,N_7378,N_7387);
xor U8380 (N_8380,N_7290,N_7635);
and U8381 (N_8381,N_7547,N_7211);
nand U8382 (N_8382,N_7263,N_7787);
nand U8383 (N_8383,N_7227,N_7772);
nand U8384 (N_8384,N_7284,N_7469);
or U8385 (N_8385,N_7276,N_7315);
nand U8386 (N_8386,N_7599,N_7586);
xnor U8387 (N_8387,N_7360,N_7267);
nand U8388 (N_8388,N_7489,N_7493);
xor U8389 (N_8389,N_7501,N_7546);
nor U8390 (N_8390,N_7485,N_7677);
nand U8391 (N_8391,N_7477,N_7671);
nand U8392 (N_8392,N_7683,N_7671);
or U8393 (N_8393,N_7307,N_7397);
nand U8394 (N_8394,N_7200,N_7341);
or U8395 (N_8395,N_7413,N_7630);
nand U8396 (N_8396,N_7237,N_7728);
nor U8397 (N_8397,N_7517,N_7214);
nand U8398 (N_8398,N_7603,N_7418);
nand U8399 (N_8399,N_7515,N_7566);
nor U8400 (N_8400,N_8307,N_7922);
nand U8401 (N_8401,N_7818,N_8198);
nor U8402 (N_8402,N_8295,N_8303);
or U8403 (N_8403,N_7825,N_8048);
and U8404 (N_8404,N_8069,N_7841);
nand U8405 (N_8405,N_8175,N_8078);
nor U8406 (N_8406,N_8352,N_8002);
nor U8407 (N_8407,N_8353,N_8298);
or U8408 (N_8408,N_8237,N_7964);
and U8409 (N_8409,N_8221,N_8385);
and U8410 (N_8410,N_8266,N_8196);
nor U8411 (N_8411,N_8128,N_8022);
or U8412 (N_8412,N_8099,N_8308);
and U8413 (N_8413,N_7835,N_8034);
nand U8414 (N_8414,N_7819,N_8315);
or U8415 (N_8415,N_8351,N_7847);
or U8416 (N_8416,N_8077,N_8043);
nor U8417 (N_8417,N_8359,N_8019);
nand U8418 (N_8418,N_7966,N_7807);
nor U8419 (N_8419,N_8345,N_8324);
and U8420 (N_8420,N_8013,N_7815);
nand U8421 (N_8421,N_8326,N_8086);
nor U8422 (N_8422,N_8375,N_7896);
xor U8423 (N_8423,N_8286,N_8178);
xnor U8424 (N_8424,N_8316,N_7809);
nand U8425 (N_8425,N_7906,N_8261);
or U8426 (N_8426,N_8249,N_8393);
or U8427 (N_8427,N_7822,N_8103);
nor U8428 (N_8428,N_8183,N_8205);
nor U8429 (N_8429,N_7853,N_8160);
nor U8430 (N_8430,N_8235,N_7907);
and U8431 (N_8431,N_8081,N_8039);
xor U8432 (N_8432,N_8306,N_7942);
or U8433 (N_8433,N_7990,N_8123);
nor U8434 (N_8434,N_8159,N_7876);
nor U8435 (N_8435,N_8384,N_8096);
or U8436 (N_8436,N_8149,N_8387);
nand U8437 (N_8437,N_7851,N_8218);
or U8438 (N_8438,N_8255,N_8113);
nor U8439 (N_8439,N_8390,N_7960);
and U8440 (N_8440,N_8024,N_8314);
nand U8441 (N_8441,N_7892,N_7806);
or U8442 (N_8442,N_8190,N_8110);
or U8443 (N_8443,N_8341,N_8246);
xnor U8444 (N_8444,N_8343,N_8289);
nand U8445 (N_8445,N_8256,N_7840);
nor U8446 (N_8446,N_8272,N_7808);
and U8447 (N_8447,N_7885,N_7828);
nor U8448 (N_8448,N_7869,N_7925);
and U8449 (N_8449,N_8346,N_8092);
xor U8450 (N_8450,N_8365,N_7977);
or U8451 (N_8451,N_7895,N_8065);
xor U8452 (N_8452,N_8072,N_8154);
nor U8453 (N_8453,N_8373,N_7918);
xor U8454 (N_8454,N_8150,N_8049);
or U8455 (N_8455,N_8056,N_7926);
nor U8456 (N_8456,N_8283,N_8066);
and U8457 (N_8457,N_7951,N_8233);
nor U8458 (N_8458,N_8085,N_8126);
or U8459 (N_8459,N_7865,N_8177);
nor U8460 (N_8460,N_8001,N_8089);
or U8461 (N_8461,N_7888,N_8293);
and U8462 (N_8462,N_8100,N_7909);
and U8463 (N_8463,N_8282,N_8216);
or U8464 (N_8464,N_8259,N_8379);
xnor U8465 (N_8465,N_8260,N_8084);
xnor U8466 (N_8466,N_8142,N_8374);
and U8467 (N_8467,N_8036,N_7810);
xnor U8468 (N_8468,N_7861,N_8309);
xor U8469 (N_8469,N_8277,N_7991);
and U8470 (N_8470,N_7967,N_7912);
or U8471 (N_8471,N_7893,N_7843);
xnor U8472 (N_8472,N_7997,N_8355);
or U8473 (N_8473,N_8264,N_8120);
xnor U8474 (N_8474,N_7911,N_8111);
xor U8475 (N_8475,N_7954,N_8155);
nand U8476 (N_8476,N_7987,N_8076);
nand U8477 (N_8477,N_7894,N_8370);
and U8478 (N_8478,N_8396,N_8145);
nor U8479 (N_8479,N_7812,N_7972);
xnor U8480 (N_8480,N_7996,N_7953);
or U8481 (N_8481,N_7859,N_8224);
xnor U8482 (N_8482,N_8029,N_8129);
xor U8483 (N_8483,N_8340,N_8025);
and U8484 (N_8484,N_8281,N_7927);
nand U8485 (N_8485,N_7978,N_8347);
xnor U8486 (N_8486,N_8189,N_7962);
nand U8487 (N_8487,N_8187,N_7916);
nand U8488 (N_8488,N_8135,N_8262);
nor U8489 (N_8489,N_8248,N_8383);
xor U8490 (N_8490,N_7948,N_8210);
or U8491 (N_8491,N_8234,N_8124);
xor U8492 (N_8492,N_8033,N_8222);
and U8493 (N_8493,N_8180,N_8334);
nor U8494 (N_8494,N_8068,N_8392);
or U8495 (N_8495,N_7880,N_8213);
nand U8496 (N_8496,N_8220,N_8217);
xor U8497 (N_8497,N_8284,N_8391);
xnor U8498 (N_8498,N_7946,N_8348);
nand U8499 (N_8499,N_8073,N_7921);
and U8500 (N_8500,N_8018,N_8325);
nor U8501 (N_8501,N_8361,N_8055);
nor U8502 (N_8502,N_7844,N_7868);
nor U8503 (N_8503,N_8265,N_8020);
or U8504 (N_8504,N_7845,N_8227);
nor U8505 (N_8505,N_8014,N_7802);
xnor U8506 (N_8506,N_8226,N_8063);
nand U8507 (N_8507,N_8143,N_7804);
nand U8508 (N_8508,N_8389,N_8125);
xnor U8509 (N_8509,N_7905,N_7832);
nand U8510 (N_8510,N_8269,N_7849);
and U8511 (N_8511,N_7898,N_8268);
nor U8512 (N_8512,N_8026,N_8007);
nor U8513 (N_8513,N_8208,N_8134);
or U8514 (N_8514,N_8109,N_7831);
and U8515 (N_8515,N_8161,N_8206);
nand U8516 (N_8516,N_7930,N_8299);
nand U8517 (N_8517,N_7834,N_8045);
xor U8518 (N_8518,N_7856,N_8288);
or U8519 (N_8519,N_8236,N_8164);
or U8520 (N_8520,N_7877,N_7854);
nor U8521 (N_8521,N_7914,N_8053);
nor U8522 (N_8522,N_8075,N_8057);
nor U8523 (N_8523,N_8214,N_7986);
nor U8524 (N_8524,N_7936,N_8193);
xnor U8525 (N_8525,N_7910,N_7857);
and U8526 (N_8526,N_8332,N_7801);
xor U8527 (N_8527,N_8093,N_8195);
and U8528 (N_8528,N_7993,N_7873);
nor U8529 (N_8529,N_7943,N_7886);
and U8530 (N_8530,N_7855,N_7814);
and U8531 (N_8531,N_7870,N_7933);
xnor U8532 (N_8532,N_7823,N_7887);
and U8533 (N_8533,N_8207,N_7864);
and U8534 (N_8534,N_7929,N_7908);
and U8535 (N_8535,N_8165,N_7891);
and U8536 (N_8536,N_8238,N_8139);
and U8537 (N_8537,N_8215,N_7924);
or U8538 (N_8538,N_8015,N_7989);
or U8539 (N_8539,N_7973,N_8058);
nand U8540 (N_8540,N_8270,N_8098);
or U8541 (N_8541,N_8245,N_8241);
nand U8542 (N_8542,N_8380,N_8037);
or U8543 (N_8543,N_7837,N_8051);
and U8544 (N_8544,N_8292,N_7836);
or U8545 (N_8545,N_8356,N_7913);
xor U8546 (N_8546,N_8127,N_8382);
or U8547 (N_8547,N_7867,N_8192);
or U8548 (N_8548,N_8080,N_8223);
and U8549 (N_8549,N_8074,N_8367);
and U8550 (N_8550,N_8267,N_7866);
nor U8551 (N_8551,N_8354,N_8004);
xnor U8552 (N_8552,N_7850,N_8225);
nor U8553 (N_8553,N_7902,N_8122);
xor U8554 (N_8554,N_8318,N_8242);
and U8555 (N_8555,N_7949,N_8174);
nor U8556 (N_8556,N_8179,N_8000);
nand U8557 (N_8557,N_8357,N_8202);
xnor U8558 (N_8558,N_7963,N_8204);
nor U8559 (N_8559,N_8031,N_7934);
and U8560 (N_8560,N_7992,N_8230);
and U8561 (N_8561,N_8136,N_7899);
and U8562 (N_8562,N_8251,N_8319);
nand U8563 (N_8563,N_8144,N_8006);
nand U8564 (N_8564,N_8366,N_7875);
nand U8565 (N_8565,N_8027,N_8231);
or U8566 (N_8566,N_8138,N_8276);
or U8567 (N_8567,N_7862,N_7939);
nand U8568 (N_8568,N_8108,N_8083);
nor U8569 (N_8569,N_7879,N_8331);
or U8570 (N_8570,N_8378,N_8082);
and U8571 (N_8571,N_8200,N_8012);
nor U8572 (N_8572,N_8046,N_7817);
or U8573 (N_8573,N_8239,N_8054);
nor U8574 (N_8574,N_8335,N_8350);
nor U8575 (N_8575,N_8003,N_8243);
or U8576 (N_8576,N_8016,N_8317);
nand U8577 (N_8577,N_8030,N_7999);
or U8578 (N_8578,N_7816,N_8360);
nor U8579 (N_8579,N_7821,N_8398);
xnor U8580 (N_8580,N_8040,N_8369);
and U8581 (N_8581,N_8185,N_8171);
or U8582 (N_8582,N_7863,N_7998);
nand U8583 (N_8583,N_8130,N_7931);
nor U8584 (N_8584,N_7995,N_8302);
nor U8585 (N_8585,N_7874,N_8064);
nand U8586 (N_8586,N_8168,N_8010);
xnor U8587 (N_8587,N_8313,N_7965);
nor U8588 (N_8588,N_8312,N_7935);
xor U8589 (N_8589,N_8199,N_8156);
nand U8590 (N_8590,N_8011,N_8140);
nand U8591 (N_8591,N_8062,N_7915);
and U8592 (N_8592,N_8333,N_8087);
and U8593 (N_8593,N_8059,N_8381);
and U8594 (N_8594,N_8050,N_7852);
nor U8595 (N_8595,N_8052,N_7824);
nand U8596 (N_8596,N_8151,N_7839);
nor U8597 (N_8597,N_8349,N_7803);
or U8598 (N_8598,N_8273,N_8327);
or U8599 (N_8599,N_7950,N_8368);
nor U8600 (N_8600,N_8336,N_8364);
nor U8601 (N_8601,N_7890,N_8290);
nor U8602 (N_8602,N_8294,N_8329);
xnor U8603 (N_8603,N_8363,N_7955);
nor U8604 (N_8604,N_8097,N_7884);
nand U8605 (N_8605,N_7872,N_7826);
and U8606 (N_8606,N_8395,N_8131);
and U8607 (N_8607,N_7820,N_7979);
or U8608 (N_8608,N_8115,N_8009);
and U8609 (N_8609,N_8291,N_8170);
nand U8610 (N_8610,N_8148,N_8061);
xor U8611 (N_8611,N_7968,N_8119);
xor U8612 (N_8612,N_8163,N_8219);
and U8613 (N_8613,N_8152,N_8362);
nand U8614 (N_8614,N_7944,N_7846);
and U8615 (N_8615,N_8181,N_8188);
or U8616 (N_8616,N_7938,N_8176);
and U8617 (N_8617,N_8047,N_8280);
nor U8618 (N_8618,N_8132,N_8250);
and U8619 (N_8619,N_8301,N_8133);
and U8620 (N_8620,N_8141,N_8028);
nand U8621 (N_8621,N_8310,N_8274);
or U8622 (N_8622,N_8258,N_8229);
nand U8623 (N_8623,N_8147,N_7903);
nand U8624 (N_8624,N_8090,N_8008);
nand U8625 (N_8625,N_8167,N_8311);
nand U8626 (N_8626,N_8182,N_8067);
and U8627 (N_8627,N_7830,N_7994);
or U8628 (N_8628,N_7842,N_8337);
nand U8629 (N_8629,N_8263,N_7860);
nand U8630 (N_8630,N_8186,N_8376);
or U8631 (N_8631,N_8116,N_8191);
and U8632 (N_8632,N_7848,N_7988);
or U8633 (N_8633,N_7920,N_8254);
xor U8634 (N_8634,N_8112,N_7829);
and U8635 (N_8635,N_7959,N_8240);
xor U8636 (N_8636,N_8173,N_7981);
xnor U8637 (N_8637,N_7974,N_8095);
xnor U8638 (N_8638,N_8114,N_8257);
nand U8639 (N_8639,N_7901,N_7945);
and U8640 (N_8640,N_7969,N_8275);
nor U8641 (N_8641,N_7941,N_8285);
nor U8642 (N_8642,N_7919,N_8107);
nor U8643 (N_8643,N_8042,N_8371);
and U8644 (N_8644,N_8005,N_8194);
nor U8645 (N_8645,N_8228,N_7878);
nor U8646 (N_8646,N_8287,N_8158);
or U8647 (N_8647,N_7937,N_8017);
or U8648 (N_8648,N_8023,N_7975);
and U8649 (N_8649,N_7940,N_8358);
and U8650 (N_8650,N_8021,N_8338);
xor U8651 (N_8651,N_8044,N_8088);
xnor U8652 (N_8652,N_8106,N_8328);
nand U8653 (N_8653,N_8038,N_7917);
nand U8654 (N_8654,N_7984,N_8397);
nand U8655 (N_8655,N_8094,N_8102);
xor U8656 (N_8656,N_8322,N_8394);
and U8657 (N_8657,N_8157,N_8169);
and U8658 (N_8658,N_7947,N_8344);
nor U8659 (N_8659,N_8279,N_8079);
and U8660 (N_8660,N_7883,N_7800);
nand U8661 (N_8661,N_7889,N_7858);
and U8662 (N_8662,N_7985,N_8304);
nand U8663 (N_8663,N_8247,N_7813);
or U8664 (N_8664,N_8137,N_7805);
xnor U8665 (N_8665,N_7980,N_8071);
nand U8666 (N_8666,N_7956,N_8118);
nand U8667 (N_8667,N_8297,N_8342);
or U8668 (N_8668,N_8323,N_8339);
nor U8669 (N_8669,N_7833,N_8032);
and U8670 (N_8670,N_8211,N_8166);
xor U8671 (N_8671,N_7957,N_7958);
or U8672 (N_8672,N_8146,N_8117);
nand U8673 (N_8673,N_8212,N_7976);
or U8674 (N_8674,N_8399,N_7923);
nand U8675 (N_8675,N_8105,N_8296);
xnor U8676 (N_8676,N_7971,N_8244);
nand U8677 (N_8677,N_8041,N_8104);
and U8678 (N_8678,N_7900,N_7881);
xor U8679 (N_8679,N_8197,N_8184);
nor U8680 (N_8680,N_7827,N_7811);
or U8681 (N_8681,N_8203,N_8330);
or U8682 (N_8682,N_7961,N_7897);
nand U8683 (N_8683,N_7871,N_7882);
or U8684 (N_8684,N_8060,N_8091);
nand U8685 (N_8685,N_8278,N_7932);
and U8686 (N_8686,N_7982,N_8172);
nand U8687 (N_8687,N_8201,N_8271);
xor U8688 (N_8688,N_8300,N_8320);
nor U8689 (N_8689,N_8035,N_8070);
or U8690 (N_8690,N_7983,N_8253);
nor U8691 (N_8691,N_8153,N_8372);
xor U8692 (N_8692,N_8209,N_7838);
or U8693 (N_8693,N_8252,N_8121);
or U8694 (N_8694,N_8321,N_8162);
nor U8695 (N_8695,N_7970,N_8388);
and U8696 (N_8696,N_8305,N_7928);
nor U8697 (N_8697,N_8386,N_7904);
nor U8698 (N_8698,N_8377,N_8101);
nand U8699 (N_8699,N_8232,N_7952);
nor U8700 (N_8700,N_8382,N_8040);
nand U8701 (N_8701,N_8047,N_8397);
nand U8702 (N_8702,N_7950,N_7802);
nand U8703 (N_8703,N_8033,N_7956);
nand U8704 (N_8704,N_7873,N_8092);
or U8705 (N_8705,N_7987,N_7949);
or U8706 (N_8706,N_7930,N_7899);
nor U8707 (N_8707,N_7934,N_8125);
or U8708 (N_8708,N_7829,N_8146);
and U8709 (N_8709,N_7803,N_7807);
nor U8710 (N_8710,N_8248,N_7812);
nand U8711 (N_8711,N_7829,N_8076);
xnor U8712 (N_8712,N_8191,N_8390);
or U8713 (N_8713,N_8009,N_8226);
nand U8714 (N_8714,N_8076,N_8043);
nand U8715 (N_8715,N_7891,N_8216);
and U8716 (N_8716,N_8021,N_8090);
nand U8717 (N_8717,N_7999,N_8094);
nand U8718 (N_8718,N_8329,N_8006);
xor U8719 (N_8719,N_8370,N_8201);
xor U8720 (N_8720,N_8378,N_7811);
nand U8721 (N_8721,N_8240,N_7951);
xor U8722 (N_8722,N_7861,N_7921);
or U8723 (N_8723,N_8341,N_7932);
and U8724 (N_8724,N_8136,N_8311);
xnor U8725 (N_8725,N_7988,N_7853);
and U8726 (N_8726,N_7889,N_8183);
nor U8727 (N_8727,N_8282,N_8032);
nor U8728 (N_8728,N_8281,N_7853);
xnor U8729 (N_8729,N_7839,N_8251);
nor U8730 (N_8730,N_8313,N_8310);
nand U8731 (N_8731,N_8228,N_8082);
xor U8732 (N_8732,N_8236,N_8087);
and U8733 (N_8733,N_8075,N_8160);
and U8734 (N_8734,N_8109,N_7801);
or U8735 (N_8735,N_8183,N_8258);
xnor U8736 (N_8736,N_8300,N_8016);
nand U8737 (N_8737,N_8313,N_8393);
xor U8738 (N_8738,N_8305,N_8066);
nand U8739 (N_8739,N_8342,N_8077);
or U8740 (N_8740,N_7925,N_7909);
or U8741 (N_8741,N_8207,N_8215);
nor U8742 (N_8742,N_8197,N_8239);
nand U8743 (N_8743,N_8040,N_8094);
nor U8744 (N_8744,N_8338,N_8126);
or U8745 (N_8745,N_8140,N_8112);
nor U8746 (N_8746,N_8148,N_8166);
xnor U8747 (N_8747,N_8255,N_8346);
nor U8748 (N_8748,N_8208,N_8320);
and U8749 (N_8749,N_8001,N_8235);
and U8750 (N_8750,N_7893,N_7821);
or U8751 (N_8751,N_8399,N_7884);
xnor U8752 (N_8752,N_8039,N_7982);
xnor U8753 (N_8753,N_8141,N_8327);
or U8754 (N_8754,N_8319,N_8140);
xor U8755 (N_8755,N_7895,N_8054);
nand U8756 (N_8756,N_7987,N_8252);
or U8757 (N_8757,N_8133,N_7933);
and U8758 (N_8758,N_8001,N_7891);
nand U8759 (N_8759,N_7926,N_8140);
xnor U8760 (N_8760,N_7865,N_8280);
nor U8761 (N_8761,N_8092,N_8315);
xor U8762 (N_8762,N_8383,N_7918);
nand U8763 (N_8763,N_8293,N_8303);
and U8764 (N_8764,N_8218,N_7849);
nor U8765 (N_8765,N_7978,N_8142);
xnor U8766 (N_8766,N_8292,N_8104);
nand U8767 (N_8767,N_8345,N_7885);
nor U8768 (N_8768,N_8025,N_8261);
and U8769 (N_8769,N_8038,N_8156);
nor U8770 (N_8770,N_7974,N_8002);
xor U8771 (N_8771,N_8373,N_8123);
xnor U8772 (N_8772,N_7991,N_8330);
xor U8773 (N_8773,N_8116,N_7824);
nand U8774 (N_8774,N_8149,N_8131);
nand U8775 (N_8775,N_8351,N_8278);
nand U8776 (N_8776,N_7813,N_7892);
or U8777 (N_8777,N_8155,N_7911);
nor U8778 (N_8778,N_8024,N_8166);
nor U8779 (N_8779,N_7801,N_8199);
or U8780 (N_8780,N_8156,N_8274);
or U8781 (N_8781,N_8154,N_7986);
or U8782 (N_8782,N_8213,N_7871);
and U8783 (N_8783,N_7850,N_7838);
nor U8784 (N_8784,N_8267,N_8380);
or U8785 (N_8785,N_8390,N_8031);
and U8786 (N_8786,N_8023,N_8380);
and U8787 (N_8787,N_7987,N_7804);
nand U8788 (N_8788,N_7990,N_8347);
or U8789 (N_8789,N_7864,N_8116);
xnor U8790 (N_8790,N_7911,N_8092);
nand U8791 (N_8791,N_7835,N_7818);
xnor U8792 (N_8792,N_8345,N_7840);
nor U8793 (N_8793,N_7994,N_7849);
and U8794 (N_8794,N_7808,N_8122);
or U8795 (N_8795,N_8189,N_8206);
xor U8796 (N_8796,N_8186,N_8112);
and U8797 (N_8797,N_7882,N_7872);
and U8798 (N_8798,N_8012,N_8044);
nor U8799 (N_8799,N_7848,N_8119);
or U8800 (N_8800,N_8163,N_8079);
nand U8801 (N_8801,N_7986,N_8189);
nand U8802 (N_8802,N_8040,N_8330);
or U8803 (N_8803,N_7810,N_8035);
and U8804 (N_8804,N_7844,N_7900);
nor U8805 (N_8805,N_8229,N_7880);
xnor U8806 (N_8806,N_8010,N_8042);
and U8807 (N_8807,N_8062,N_7833);
and U8808 (N_8808,N_7901,N_7845);
or U8809 (N_8809,N_7837,N_8178);
and U8810 (N_8810,N_8080,N_8081);
xor U8811 (N_8811,N_8395,N_8336);
and U8812 (N_8812,N_7991,N_8226);
or U8813 (N_8813,N_8171,N_7897);
nand U8814 (N_8814,N_7896,N_8173);
nor U8815 (N_8815,N_8357,N_8250);
and U8816 (N_8816,N_7817,N_8079);
or U8817 (N_8817,N_7919,N_8271);
nor U8818 (N_8818,N_8089,N_7947);
or U8819 (N_8819,N_8250,N_8359);
and U8820 (N_8820,N_8179,N_8321);
nand U8821 (N_8821,N_8188,N_7831);
and U8822 (N_8822,N_8397,N_8162);
xnor U8823 (N_8823,N_8218,N_8300);
or U8824 (N_8824,N_7851,N_8338);
nor U8825 (N_8825,N_8224,N_7953);
or U8826 (N_8826,N_8122,N_8323);
nand U8827 (N_8827,N_8208,N_8389);
xor U8828 (N_8828,N_7808,N_7867);
and U8829 (N_8829,N_8351,N_8133);
and U8830 (N_8830,N_8013,N_8061);
and U8831 (N_8831,N_8103,N_7934);
xor U8832 (N_8832,N_8194,N_8315);
or U8833 (N_8833,N_7836,N_8356);
xor U8834 (N_8834,N_7981,N_8151);
nor U8835 (N_8835,N_8224,N_7984);
nor U8836 (N_8836,N_8354,N_7830);
and U8837 (N_8837,N_8155,N_8211);
xnor U8838 (N_8838,N_7935,N_8127);
nand U8839 (N_8839,N_8052,N_8083);
xnor U8840 (N_8840,N_8297,N_8341);
xor U8841 (N_8841,N_8140,N_7990);
xnor U8842 (N_8842,N_8150,N_7863);
or U8843 (N_8843,N_8352,N_7873);
and U8844 (N_8844,N_8159,N_7860);
xnor U8845 (N_8845,N_8193,N_8027);
xor U8846 (N_8846,N_8357,N_7909);
xor U8847 (N_8847,N_8224,N_8226);
and U8848 (N_8848,N_7844,N_8322);
nor U8849 (N_8849,N_8021,N_7948);
and U8850 (N_8850,N_8090,N_7943);
xor U8851 (N_8851,N_8319,N_7929);
nand U8852 (N_8852,N_7825,N_8387);
nor U8853 (N_8853,N_8332,N_8290);
nand U8854 (N_8854,N_8050,N_8366);
xnor U8855 (N_8855,N_8052,N_8257);
or U8856 (N_8856,N_7889,N_8297);
xor U8857 (N_8857,N_8203,N_7910);
and U8858 (N_8858,N_7924,N_8394);
nor U8859 (N_8859,N_7974,N_8380);
or U8860 (N_8860,N_7959,N_8229);
nor U8861 (N_8861,N_8038,N_8061);
nand U8862 (N_8862,N_8225,N_7988);
or U8863 (N_8863,N_8061,N_8067);
nor U8864 (N_8864,N_8022,N_8191);
nor U8865 (N_8865,N_7942,N_8356);
or U8866 (N_8866,N_8292,N_8093);
nand U8867 (N_8867,N_7930,N_8024);
and U8868 (N_8868,N_7947,N_7977);
and U8869 (N_8869,N_8359,N_7957);
nor U8870 (N_8870,N_8390,N_8102);
xnor U8871 (N_8871,N_8030,N_8120);
or U8872 (N_8872,N_8393,N_7885);
or U8873 (N_8873,N_8056,N_8161);
nand U8874 (N_8874,N_8159,N_8190);
nand U8875 (N_8875,N_8163,N_8059);
nand U8876 (N_8876,N_8285,N_8148);
xnor U8877 (N_8877,N_8017,N_7931);
xor U8878 (N_8878,N_7900,N_8314);
nand U8879 (N_8879,N_8376,N_8024);
and U8880 (N_8880,N_8060,N_8270);
nor U8881 (N_8881,N_8323,N_8105);
nor U8882 (N_8882,N_8190,N_7965);
nor U8883 (N_8883,N_8238,N_8261);
xnor U8884 (N_8884,N_7830,N_8288);
and U8885 (N_8885,N_8300,N_7866);
or U8886 (N_8886,N_7867,N_7971);
nor U8887 (N_8887,N_7996,N_8248);
xor U8888 (N_8888,N_8065,N_7880);
nor U8889 (N_8889,N_8152,N_8291);
xnor U8890 (N_8890,N_7933,N_7986);
nor U8891 (N_8891,N_8009,N_7996);
nor U8892 (N_8892,N_7942,N_8188);
nor U8893 (N_8893,N_7812,N_8138);
xnor U8894 (N_8894,N_7960,N_8367);
or U8895 (N_8895,N_8224,N_7850);
nand U8896 (N_8896,N_8142,N_7897);
and U8897 (N_8897,N_8183,N_7956);
nor U8898 (N_8898,N_8266,N_8088);
and U8899 (N_8899,N_8145,N_7928);
nor U8900 (N_8900,N_7880,N_7877);
xor U8901 (N_8901,N_8338,N_8251);
xnor U8902 (N_8902,N_8033,N_7982);
and U8903 (N_8903,N_8117,N_8341);
nor U8904 (N_8904,N_8149,N_7988);
and U8905 (N_8905,N_8394,N_8132);
nand U8906 (N_8906,N_7854,N_7846);
or U8907 (N_8907,N_8268,N_8178);
nand U8908 (N_8908,N_8172,N_8145);
nand U8909 (N_8909,N_8044,N_7884);
or U8910 (N_8910,N_8229,N_7914);
and U8911 (N_8911,N_8195,N_8096);
and U8912 (N_8912,N_8105,N_7888);
nand U8913 (N_8913,N_8154,N_8269);
and U8914 (N_8914,N_8192,N_7961);
nand U8915 (N_8915,N_7845,N_8376);
and U8916 (N_8916,N_8028,N_7832);
and U8917 (N_8917,N_8215,N_8023);
nor U8918 (N_8918,N_8248,N_7845);
nand U8919 (N_8919,N_7893,N_8111);
and U8920 (N_8920,N_8235,N_7803);
xnor U8921 (N_8921,N_7861,N_7890);
and U8922 (N_8922,N_8266,N_7801);
nand U8923 (N_8923,N_8068,N_7826);
and U8924 (N_8924,N_8112,N_8178);
nand U8925 (N_8925,N_8129,N_7870);
nand U8926 (N_8926,N_8047,N_7948);
nand U8927 (N_8927,N_8024,N_8254);
nand U8928 (N_8928,N_7959,N_8231);
nand U8929 (N_8929,N_8333,N_8051);
and U8930 (N_8930,N_8332,N_8001);
nor U8931 (N_8931,N_8077,N_8141);
nor U8932 (N_8932,N_7987,N_8111);
nand U8933 (N_8933,N_8348,N_8283);
or U8934 (N_8934,N_8055,N_8316);
xnor U8935 (N_8935,N_8093,N_8343);
and U8936 (N_8936,N_8171,N_8082);
nand U8937 (N_8937,N_8324,N_8268);
or U8938 (N_8938,N_8355,N_8257);
xnor U8939 (N_8939,N_7925,N_8132);
xor U8940 (N_8940,N_8195,N_8049);
nand U8941 (N_8941,N_8268,N_8208);
nand U8942 (N_8942,N_8237,N_8229);
xnor U8943 (N_8943,N_8024,N_8312);
or U8944 (N_8944,N_8330,N_8156);
or U8945 (N_8945,N_8153,N_8071);
or U8946 (N_8946,N_7903,N_8047);
nor U8947 (N_8947,N_8004,N_8161);
and U8948 (N_8948,N_8071,N_8148);
and U8949 (N_8949,N_7816,N_8246);
or U8950 (N_8950,N_8120,N_8313);
and U8951 (N_8951,N_8343,N_8102);
xnor U8952 (N_8952,N_8342,N_8233);
and U8953 (N_8953,N_7986,N_8296);
nand U8954 (N_8954,N_8114,N_8100);
and U8955 (N_8955,N_8004,N_8397);
xnor U8956 (N_8956,N_7821,N_8335);
nand U8957 (N_8957,N_8357,N_7810);
or U8958 (N_8958,N_8025,N_8127);
and U8959 (N_8959,N_7880,N_7911);
xnor U8960 (N_8960,N_8211,N_8054);
nand U8961 (N_8961,N_8136,N_8379);
and U8962 (N_8962,N_7870,N_7894);
or U8963 (N_8963,N_8169,N_8351);
xor U8964 (N_8964,N_7994,N_8019);
nor U8965 (N_8965,N_8087,N_8100);
and U8966 (N_8966,N_8046,N_8252);
and U8967 (N_8967,N_8157,N_8147);
and U8968 (N_8968,N_7825,N_7873);
and U8969 (N_8969,N_7842,N_7995);
and U8970 (N_8970,N_8129,N_8296);
and U8971 (N_8971,N_8134,N_8041);
and U8972 (N_8972,N_8344,N_8221);
nand U8973 (N_8973,N_8025,N_8078);
and U8974 (N_8974,N_7906,N_8124);
nand U8975 (N_8975,N_8115,N_8068);
or U8976 (N_8976,N_7851,N_8359);
nor U8977 (N_8977,N_8125,N_8023);
or U8978 (N_8978,N_8168,N_7882);
xor U8979 (N_8979,N_8325,N_7896);
xnor U8980 (N_8980,N_8183,N_8249);
xnor U8981 (N_8981,N_7991,N_8286);
xor U8982 (N_8982,N_7841,N_8039);
and U8983 (N_8983,N_8341,N_7806);
and U8984 (N_8984,N_8021,N_8056);
nor U8985 (N_8985,N_8165,N_8212);
nor U8986 (N_8986,N_8359,N_7994);
or U8987 (N_8987,N_8069,N_8189);
and U8988 (N_8988,N_7801,N_7820);
and U8989 (N_8989,N_7970,N_8333);
nor U8990 (N_8990,N_8013,N_7974);
nor U8991 (N_8991,N_7991,N_8018);
xnor U8992 (N_8992,N_7844,N_8381);
or U8993 (N_8993,N_7939,N_7904);
nor U8994 (N_8994,N_8336,N_7908);
or U8995 (N_8995,N_8069,N_8007);
nor U8996 (N_8996,N_8335,N_7928);
or U8997 (N_8997,N_8213,N_8247);
nand U8998 (N_8998,N_8378,N_8021);
xnor U8999 (N_8999,N_7856,N_7925);
nor U9000 (N_9000,N_8413,N_8991);
nor U9001 (N_9001,N_8512,N_8587);
xnor U9002 (N_9002,N_8656,N_8667);
xor U9003 (N_9003,N_8535,N_8657);
nand U9004 (N_9004,N_8670,N_8415);
xor U9005 (N_9005,N_8430,N_8631);
nand U9006 (N_9006,N_8938,N_8486);
nand U9007 (N_9007,N_8465,N_8993);
and U9008 (N_9008,N_8899,N_8922);
xor U9009 (N_9009,N_8969,N_8616);
nor U9010 (N_9010,N_8572,N_8680);
or U9011 (N_9011,N_8596,N_8927);
nand U9012 (N_9012,N_8685,N_8487);
nand U9013 (N_9013,N_8763,N_8982);
or U9014 (N_9014,N_8962,N_8751);
nor U9015 (N_9015,N_8480,N_8752);
xnor U9016 (N_9016,N_8466,N_8437);
and U9017 (N_9017,N_8771,N_8961);
nor U9018 (N_9018,N_8711,N_8633);
nor U9019 (N_9019,N_8707,N_8626);
xnor U9020 (N_9020,N_8440,N_8674);
or U9021 (N_9021,N_8689,N_8839);
nand U9022 (N_9022,N_8911,N_8948);
nand U9023 (N_9023,N_8936,N_8560);
nand U9024 (N_9024,N_8421,N_8873);
or U9025 (N_9025,N_8518,N_8985);
xor U9026 (N_9026,N_8973,N_8640);
xor U9027 (N_9027,N_8916,N_8741);
xnor U9028 (N_9028,N_8809,N_8409);
xor U9029 (N_9029,N_8800,N_8979);
or U9030 (N_9030,N_8713,N_8438);
xnor U9031 (N_9031,N_8792,N_8723);
and U9032 (N_9032,N_8468,N_8523);
and U9033 (N_9033,N_8412,N_8545);
or U9034 (N_9034,N_8567,N_8872);
nor U9035 (N_9035,N_8450,N_8914);
and U9036 (N_9036,N_8658,N_8416);
and U9037 (N_9037,N_8770,N_8506);
nand U9038 (N_9038,N_8490,N_8503);
xnor U9039 (N_9039,N_8819,N_8576);
nand U9040 (N_9040,N_8875,N_8732);
xnor U9041 (N_9041,N_8470,N_8403);
or U9042 (N_9042,N_8501,N_8853);
or U9043 (N_9043,N_8758,N_8821);
xnor U9044 (N_9044,N_8692,N_8897);
xnor U9045 (N_9045,N_8739,N_8900);
or U9046 (N_9046,N_8942,N_8447);
or U9047 (N_9047,N_8791,N_8434);
or U9048 (N_9048,N_8599,N_8600);
xnor U9049 (N_9049,N_8983,N_8887);
and U9050 (N_9050,N_8925,N_8426);
or U9051 (N_9051,N_8433,N_8749);
or U9052 (N_9052,N_8917,N_8786);
nand U9053 (N_9053,N_8902,N_8418);
nand U9054 (N_9054,N_8452,N_8830);
or U9055 (N_9055,N_8642,N_8762);
nor U9056 (N_9056,N_8919,N_8414);
xnor U9057 (N_9057,N_8638,N_8442);
or U9058 (N_9058,N_8605,N_8530);
nand U9059 (N_9059,N_8876,N_8775);
xnor U9060 (N_9060,N_8457,N_8851);
nand U9061 (N_9061,N_8767,N_8491);
and U9062 (N_9062,N_8498,N_8539);
nand U9063 (N_9063,N_8582,N_8548);
nor U9064 (N_9064,N_8987,N_8878);
and U9065 (N_9065,N_8536,N_8688);
and U9066 (N_9066,N_8428,N_8419);
xnor U9067 (N_9067,N_8628,N_8533);
and U9068 (N_9068,N_8779,N_8402);
xor U9069 (N_9069,N_8777,N_8731);
nand U9070 (N_9070,N_8697,N_8829);
or U9071 (N_9071,N_8773,N_8882);
and U9072 (N_9072,N_8635,N_8462);
xor U9073 (N_9073,N_8508,N_8888);
nor U9074 (N_9074,N_8684,N_8890);
and U9075 (N_9075,N_8977,N_8643);
xnor U9076 (N_9076,N_8496,N_8517);
nor U9077 (N_9077,N_8672,N_8666);
nor U9078 (N_9078,N_8696,N_8592);
xor U9079 (N_9079,N_8422,N_8504);
and U9080 (N_9080,N_8717,N_8528);
or U9081 (N_9081,N_8476,N_8444);
or U9082 (N_9082,N_8677,N_8669);
or U9083 (N_9083,N_8651,N_8509);
xor U9084 (N_9084,N_8510,N_8683);
xor U9085 (N_9085,N_8482,N_8744);
nand U9086 (N_9086,N_8427,N_8710);
xnor U9087 (N_9087,N_8789,N_8924);
xnor U9088 (N_9088,N_8860,N_8694);
nand U9089 (N_9089,N_8755,N_8443);
and U9090 (N_9090,N_8661,N_8594);
and U9091 (N_9091,N_8960,N_8893);
nor U9092 (N_9092,N_8701,N_8810);
and U9093 (N_9093,N_8928,N_8679);
nand U9094 (N_9094,N_8579,N_8995);
or U9095 (N_9095,N_8400,N_8782);
and U9096 (N_9096,N_8757,N_8654);
nor U9097 (N_9097,N_8593,N_8514);
and U9098 (N_9098,N_8774,N_8542);
and U9099 (N_9099,N_8602,N_8889);
and U9100 (N_9100,N_8996,N_8648);
or U9101 (N_9101,N_8502,N_8735);
nor U9102 (N_9102,N_8583,N_8479);
and U9103 (N_9103,N_8745,N_8954);
or U9104 (N_9104,N_8841,N_8458);
and U9105 (N_9105,N_8705,N_8531);
and U9106 (N_9106,N_8994,N_8891);
xor U9107 (N_9107,N_8702,N_8526);
xnor U9108 (N_9108,N_8904,N_8975);
xnor U9109 (N_9109,N_8984,N_8577);
or U9110 (N_9110,N_8788,N_8483);
nor U9111 (N_9111,N_8898,N_8424);
and U9112 (N_9112,N_8877,N_8801);
nand U9113 (N_9113,N_8551,N_8737);
or U9114 (N_9114,N_8456,N_8691);
and U9115 (N_9115,N_8401,N_8718);
nor U9116 (N_9116,N_8842,N_8929);
nor U9117 (N_9117,N_8838,N_8624);
and U9118 (N_9118,N_8817,N_8974);
nor U9119 (N_9119,N_8949,N_8441);
or U9120 (N_9120,N_8429,N_8915);
or U9121 (N_9121,N_8734,N_8497);
xnor U9122 (N_9122,N_8549,N_8460);
xor U9123 (N_9123,N_8586,N_8826);
and U9124 (N_9124,N_8719,N_8469);
nor U9125 (N_9125,N_8619,N_8472);
nor U9126 (N_9126,N_8761,N_8404);
xor U9127 (N_9127,N_8935,N_8566);
nor U9128 (N_9128,N_8556,N_8453);
and U9129 (N_9129,N_8562,N_8866);
nor U9130 (N_9130,N_8471,N_8781);
or U9131 (N_9131,N_8709,N_8668);
xnor U9132 (N_9132,N_8495,N_8724);
or U9133 (N_9133,N_8417,N_8959);
xnor U9134 (N_9134,N_8952,N_8563);
nand U9135 (N_9135,N_8541,N_8647);
or U9136 (N_9136,N_8499,N_8478);
nand U9137 (N_9137,N_8520,N_8843);
xnor U9138 (N_9138,N_8609,N_8910);
nand U9139 (N_9139,N_8507,N_8653);
xor U9140 (N_9140,N_8815,N_8715);
xnor U9141 (N_9141,N_8997,N_8513);
nand U9142 (N_9142,N_8604,N_8601);
xor U9143 (N_9143,N_8550,N_8448);
nand U9144 (N_9144,N_8760,N_8931);
xnor U9145 (N_9145,N_8884,N_8671);
or U9146 (N_9146,N_8637,N_8958);
nor U9147 (N_9147,N_8909,N_8613);
nor U9148 (N_9148,N_8611,N_8913);
or U9149 (N_9149,N_8607,N_8743);
or U9150 (N_9150,N_8708,N_8742);
or U9151 (N_9151,N_8690,N_8765);
and U9152 (N_9152,N_8716,N_8967);
or U9153 (N_9153,N_8639,N_8617);
nand U9154 (N_9154,N_8733,N_8858);
nor U9155 (N_9155,N_8759,N_8591);
nand U9156 (N_9156,N_8516,N_8880);
xnor U9157 (N_9157,N_8461,N_8540);
nor U9158 (N_9158,N_8662,N_8620);
nand U9159 (N_9159,N_8769,N_8570);
or U9160 (N_9160,N_8901,N_8941);
nor U9161 (N_9161,N_8831,N_8807);
xor U9162 (N_9162,N_8699,N_8874);
and U9163 (N_9163,N_8822,N_8706);
nand U9164 (N_9164,N_8747,N_8623);
nor U9165 (N_9165,N_8976,N_8603);
xnor U9166 (N_9166,N_8663,N_8870);
xor U9167 (N_9167,N_8787,N_8748);
nor U9168 (N_9168,N_8721,N_8998);
or U9169 (N_9169,N_8864,N_8722);
nand U9170 (N_9170,N_8802,N_8956);
nand U9171 (N_9171,N_8565,N_8795);
and U9172 (N_9172,N_8678,N_8580);
nor U9173 (N_9173,N_8978,N_8793);
or U9174 (N_9174,N_8686,N_8855);
xor U9175 (N_9175,N_8644,N_8695);
or U9176 (N_9176,N_8538,N_8459);
xor U9177 (N_9177,N_8406,N_8756);
or U9178 (N_9178,N_8848,N_8753);
and U9179 (N_9179,N_8981,N_8816);
xnor U9180 (N_9180,N_8687,N_8559);
nor U9181 (N_9181,N_8629,N_8896);
nor U9182 (N_9182,N_8595,N_8423);
or U9183 (N_9183,N_8488,N_8812);
or U9184 (N_9184,N_8803,N_8589);
nor U9185 (N_9185,N_8828,N_8971);
or U9186 (N_9186,N_8546,N_8923);
xor U9187 (N_9187,N_8703,N_8989);
or U9188 (N_9188,N_8473,N_8966);
or U9189 (N_9189,N_8554,N_8411);
nor U9190 (N_9190,N_8581,N_8664);
xor U9191 (N_9191,N_8799,N_8537);
or U9192 (N_9192,N_8934,N_8933);
nor U9193 (N_9193,N_8944,N_8578);
or U9194 (N_9194,N_8432,N_8521);
and U9195 (N_9195,N_8818,N_8854);
nor U9196 (N_9196,N_8436,N_8811);
xnor U9197 (N_9197,N_8806,N_8634);
nand U9198 (N_9198,N_8790,N_8920);
or U9199 (N_9199,N_8772,N_8867);
or U9200 (N_9200,N_8840,N_8868);
and U9201 (N_9201,N_8797,N_8492);
xor U9202 (N_9202,N_8764,N_8879);
xnor U9203 (N_9203,N_8435,N_8675);
or U9204 (N_9204,N_8992,N_8704);
nand U9205 (N_9205,N_8439,N_8885);
xnor U9206 (N_9206,N_8814,N_8836);
or U9207 (N_9207,N_8676,N_8474);
nand U9208 (N_9208,N_8606,N_8859);
xnor U9209 (N_9209,N_8446,N_8780);
nor U9210 (N_9210,N_8588,N_8646);
nor U9211 (N_9211,N_8532,N_8527);
nor U9212 (N_9212,N_8543,N_8905);
or U9213 (N_9213,N_8481,N_8522);
xnor U9214 (N_9214,N_8571,N_8895);
xor U9215 (N_9215,N_8844,N_8950);
xor U9216 (N_9216,N_8608,N_8903);
xor U9217 (N_9217,N_8740,N_8846);
and U9218 (N_9218,N_8988,N_8585);
or U9219 (N_9219,N_8652,N_8785);
or U9220 (N_9220,N_8776,N_8798);
and U9221 (N_9221,N_8625,N_8477);
nor U9222 (N_9222,N_8636,N_8832);
or U9223 (N_9223,N_8912,N_8784);
and U9224 (N_9224,N_8932,N_8597);
or U9225 (N_9225,N_8622,N_8746);
and U9226 (N_9226,N_8660,N_8693);
or U9227 (N_9227,N_8930,N_8804);
nor U9228 (N_9228,N_8455,N_8632);
or U9229 (N_9229,N_8584,N_8943);
nor U9230 (N_9230,N_8552,N_8738);
xnor U9231 (N_9231,N_8500,N_8407);
nor U9232 (N_9232,N_8894,N_8778);
and U9233 (N_9233,N_8980,N_8820);
or U9234 (N_9234,N_8869,N_8673);
xor U9235 (N_9235,N_8610,N_8965);
nor U9236 (N_9236,N_8529,N_8856);
or U9237 (N_9237,N_8852,N_8445);
nand U9238 (N_9238,N_8926,N_8698);
nand U9239 (N_9239,N_8999,N_8865);
nor U9240 (N_9240,N_8768,N_8525);
or U9241 (N_9241,N_8964,N_8425);
and U9242 (N_9242,N_8645,N_8655);
nor U9243 (N_9243,N_8957,N_8485);
xnor U9244 (N_9244,N_8939,N_8649);
nor U9245 (N_9245,N_8547,N_8863);
or U9246 (N_9246,N_8464,N_8544);
or U9247 (N_9247,N_8754,N_8682);
and U9248 (N_9248,N_8847,N_8727);
xnor U9249 (N_9249,N_8730,N_8451);
nand U9250 (N_9250,N_8835,N_8720);
and U9251 (N_9251,N_8849,N_8953);
xor U9252 (N_9252,N_8630,N_8845);
or U9253 (N_9253,N_8805,N_8568);
and U9254 (N_9254,N_8505,N_8918);
xnor U9255 (N_9255,N_8850,N_8986);
and U9256 (N_9256,N_8946,N_8665);
nand U9257 (N_9257,N_8834,N_8725);
or U9258 (N_9258,N_8883,N_8467);
or U9259 (N_9259,N_8534,N_8825);
nand U9260 (N_9260,N_8621,N_8783);
nand U9261 (N_9261,N_8921,N_8558);
or U9262 (N_9262,N_8574,N_8493);
or U9263 (N_9263,N_8614,N_8555);
and U9264 (N_9264,N_8951,N_8886);
and U9265 (N_9265,N_8736,N_8837);
xnor U9266 (N_9266,N_8519,N_8972);
or U9267 (N_9267,N_8553,N_8908);
xor U9268 (N_9268,N_8612,N_8454);
and U9269 (N_9269,N_8489,N_8557);
and U9270 (N_9270,N_8650,N_8405);
xor U9271 (N_9271,N_8449,N_8431);
nor U9272 (N_9272,N_8641,N_8766);
or U9273 (N_9273,N_8824,N_8420);
nand U9274 (N_9274,N_8871,N_8861);
xnor U9275 (N_9275,N_8714,N_8906);
and U9276 (N_9276,N_8794,N_8726);
or U9277 (N_9277,N_8808,N_8881);
and U9278 (N_9278,N_8627,N_8590);
and U9279 (N_9279,N_8700,N_8515);
nor U9280 (N_9280,N_8729,N_8750);
nor U9281 (N_9281,N_8892,N_8564);
and U9282 (N_9282,N_8408,N_8561);
nand U9283 (N_9283,N_8796,N_8659);
xor U9284 (N_9284,N_8618,N_8573);
nand U9285 (N_9285,N_8990,N_8823);
and U9286 (N_9286,N_8575,N_8598);
nor U9287 (N_9287,N_8569,N_8712);
or U9288 (N_9288,N_8857,N_8475);
and U9289 (N_9289,N_8511,N_8955);
nand U9290 (N_9290,N_8827,N_8937);
and U9291 (N_9291,N_8940,N_8833);
nand U9292 (N_9292,N_8968,N_8963);
nand U9293 (N_9293,N_8862,N_8410);
nor U9294 (N_9294,N_8524,N_8907);
xnor U9295 (N_9295,N_8484,N_8463);
and U9296 (N_9296,N_8494,N_8945);
nor U9297 (N_9297,N_8728,N_8970);
nor U9298 (N_9298,N_8813,N_8615);
nor U9299 (N_9299,N_8681,N_8947);
nor U9300 (N_9300,N_8701,N_8505);
and U9301 (N_9301,N_8955,N_8499);
and U9302 (N_9302,N_8711,N_8902);
nor U9303 (N_9303,N_8940,N_8869);
nor U9304 (N_9304,N_8657,N_8727);
xnor U9305 (N_9305,N_8947,N_8889);
nand U9306 (N_9306,N_8671,N_8831);
xor U9307 (N_9307,N_8634,N_8981);
or U9308 (N_9308,N_8872,N_8805);
nand U9309 (N_9309,N_8613,N_8701);
and U9310 (N_9310,N_8775,N_8538);
nor U9311 (N_9311,N_8845,N_8673);
or U9312 (N_9312,N_8431,N_8504);
or U9313 (N_9313,N_8988,N_8753);
nand U9314 (N_9314,N_8629,N_8446);
and U9315 (N_9315,N_8724,N_8899);
or U9316 (N_9316,N_8544,N_8469);
nor U9317 (N_9317,N_8826,N_8590);
xnor U9318 (N_9318,N_8447,N_8719);
xnor U9319 (N_9319,N_8535,N_8940);
and U9320 (N_9320,N_8492,N_8980);
and U9321 (N_9321,N_8751,N_8639);
or U9322 (N_9322,N_8554,N_8645);
or U9323 (N_9323,N_8833,N_8443);
nand U9324 (N_9324,N_8991,N_8974);
xnor U9325 (N_9325,N_8901,N_8742);
and U9326 (N_9326,N_8818,N_8699);
nor U9327 (N_9327,N_8756,N_8859);
or U9328 (N_9328,N_8567,N_8986);
and U9329 (N_9329,N_8411,N_8481);
xnor U9330 (N_9330,N_8403,N_8449);
and U9331 (N_9331,N_8870,N_8649);
nand U9332 (N_9332,N_8987,N_8651);
nor U9333 (N_9333,N_8978,N_8878);
or U9334 (N_9334,N_8909,N_8492);
xnor U9335 (N_9335,N_8876,N_8565);
nor U9336 (N_9336,N_8660,N_8903);
nor U9337 (N_9337,N_8879,N_8555);
and U9338 (N_9338,N_8450,N_8966);
nand U9339 (N_9339,N_8439,N_8550);
xnor U9340 (N_9340,N_8999,N_8534);
nor U9341 (N_9341,N_8985,N_8593);
xor U9342 (N_9342,N_8886,N_8575);
nor U9343 (N_9343,N_8415,N_8449);
nor U9344 (N_9344,N_8552,N_8976);
or U9345 (N_9345,N_8964,N_8749);
nand U9346 (N_9346,N_8895,N_8442);
nand U9347 (N_9347,N_8884,N_8909);
nor U9348 (N_9348,N_8468,N_8577);
xor U9349 (N_9349,N_8897,N_8412);
nor U9350 (N_9350,N_8456,N_8424);
and U9351 (N_9351,N_8948,N_8533);
and U9352 (N_9352,N_8769,N_8449);
or U9353 (N_9353,N_8975,N_8964);
xor U9354 (N_9354,N_8422,N_8915);
nor U9355 (N_9355,N_8748,N_8960);
nor U9356 (N_9356,N_8634,N_8628);
nand U9357 (N_9357,N_8867,N_8420);
xnor U9358 (N_9358,N_8743,N_8490);
or U9359 (N_9359,N_8917,N_8558);
and U9360 (N_9360,N_8851,N_8749);
nor U9361 (N_9361,N_8671,N_8574);
xnor U9362 (N_9362,N_8529,N_8705);
nor U9363 (N_9363,N_8650,N_8579);
nand U9364 (N_9364,N_8865,N_8716);
and U9365 (N_9365,N_8681,N_8996);
xnor U9366 (N_9366,N_8901,N_8651);
nand U9367 (N_9367,N_8833,N_8449);
xor U9368 (N_9368,N_8831,N_8703);
or U9369 (N_9369,N_8856,N_8661);
and U9370 (N_9370,N_8629,N_8729);
nor U9371 (N_9371,N_8483,N_8892);
nand U9372 (N_9372,N_8410,N_8848);
or U9373 (N_9373,N_8740,N_8595);
nor U9374 (N_9374,N_8705,N_8458);
nand U9375 (N_9375,N_8870,N_8967);
or U9376 (N_9376,N_8841,N_8640);
nand U9377 (N_9377,N_8930,N_8883);
nor U9378 (N_9378,N_8878,N_8816);
xor U9379 (N_9379,N_8409,N_8834);
nand U9380 (N_9380,N_8582,N_8623);
or U9381 (N_9381,N_8470,N_8555);
xor U9382 (N_9382,N_8559,N_8809);
or U9383 (N_9383,N_8923,N_8763);
or U9384 (N_9384,N_8772,N_8925);
or U9385 (N_9385,N_8572,N_8784);
xor U9386 (N_9386,N_8996,N_8909);
nor U9387 (N_9387,N_8920,N_8891);
xnor U9388 (N_9388,N_8614,N_8881);
nand U9389 (N_9389,N_8485,N_8537);
and U9390 (N_9390,N_8548,N_8588);
and U9391 (N_9391,N_8612,N_8560);
nor U9392 (N_9392,N_8965,N_8413);
and U9393 (N_9393,N_8905,N_8767);
nand U9394 (N_9394,N_8633,N_8789);
nor U9395 (N_9395,N_8648,N_8851);
and U9396 (N_9396,N_8602,N_8677);
nor U9397 (N_9397,N_8442,N_8569);
and U9398 (N_9398,N_8429,N_8411);
and U9399 (N_9399,N_8725,N_8534);
nand U9400 (N_9400,N_8451,N_8961);
nand U9401 (N_9401,N_8571,N_8749);
or U9402 (N_9402,N_8602,N_8834);
or U9403 (N_9403,N_8586,N_8963);
xor U9404 (N_9404,N_8957,N_8541);
or U9405 (N_9405,N_8452,N_8568);
nand U9406 (N_9406,N_8815,N_8631);
nand U9407 (N_9407,N_8991,N_8736);
or U9408 (N_9408,N_8808,N_8467);
or U9409 (N_9409,N_8841,N_8723);
and U9410 (N_9410,N_8587,N_8936);
or U9411 (N_9411,N_8885,N_8402);
and U9412 (N_9412,N_8637,N_8466);
nand U9413 (N_9413,N_8762,N_8989);
and U9414 (N_9414,N_8649,N_8942);
or U9415 (N_9415,N_8580,N_8579);
or U9416 (N_9416,N_8983,N_8455);
and U9417 (N_9417,N_8427,N_8659);
nand U9418 (N_9418,N_8489,N_8972);
nand U9419 (N_9419,N_8931,N_8458);
nand U9420 (N_9420,N_8483,N_8982);
or U9421 (N_9421,N_8490,N_8558);
or U9422 (N_9422,N_8493,N_8809);
nand U9423 (N_9423,N_8409,N_8716);
or U9424 (N_9424,N_8839,N_8871);
or U9425 (N_9425,N_8416,N_8487);
nand U9426 (N_9426,N_8662,N_8900);
nor U9427 (N_9427,N_8908,N_8519);
xnor U9428 (N_9428,N_8849,N_8848);
nand U9429 (N_9429,N_8564,N_8702);
nand U9430 (N_9430,N_8926,N_8984);
nor U9431 (N_9431,N_8848,N_8953);
nand U9432 (N_9432,N_8650,N_8597);
nor U9433 (N_9433,N_8548,N_8516);
and U9434 (N_9434,N_8505,N_8616);
or U9435 (N_9435,N_8638,N_8830);
xnor U9436 (N_9436,N_8565,N_8460);
or U9437 (N_9437,N_8737,N_8469);
xnor U9438 (N_9438,N_8772,N_8828);
nand U9439 (N_9439,N_8619,N_8728);
nor U9440 (N_9440,N_8696,N_8873);
and U9441 (N_9441,N_8797,N_8534);
nand U9442 (N_9442,N_8475,N_8438);
or U9443 (N_9443,N_8580,N_8726);
xor U9444 (N_9444,N_8538,N_8577);
and U9445 (N_9445,N_8444,N_8856);
or U9446 (N_9446,N_8449,N_8615);
nand U9447 (N_9447,N_8777,N_8432);
nor U9448 (N_9448,N_8477,N_8755);
or U9449 (N_9449,N_8546,N_8640);
and U9450 (N_9450,N_8785,N_8813);
xor U9451 (N_9451,N_8791,N_8907);
and U9452 (N_9452,N_8496,N_8405);
xor U9453 (N_9453,N_8958,N_8532);
nor U9454 (N_9454,N_8539,N_8456);
xor U9455 (N_9455,N_8717,N_8684);
or U9456 (N_9456,N_8625,N_8774);
or U9457 (N_9457,N_8999,N_8851);
xnor U9458 (N_9458,N_8922,N_8426);
xor U9459 (N_9459,N_8982,N_8526);
or U9460 (N_9460,N_8660,N_8872);
xor U9461 (N_9461,N_8701,N_8506);
or U9462 (N_9462,N_8839,N_8693);
and U9463 (N_9463,N_8497,N_8755);
xor U9464 (N_9464,N_8603,N_8697);
nor U9465 (N_9465,N_8926,N_8651);
nor U9466 (N_9466,N_8987,N_8917);
and U9467 (N_9467,N_8422,N_8478);
and U9468 (N_9468,N_8857,N_8809);
nand U9469 (N_9469,N_8492,N_8659);
nor U9470 (N_9470,N_8729,N_8818);
nand U9471 (N_9471,N_8524,N_8776);
xnor U9472 (N_9472,N_8798,N_8545);
and U9473 (N_9473,N_8862,N_8921);
and U9474 (N_9474,N_8911,N_8671);
or U9475 (N_9475,N_8599,N_8578);
xnor U9476 (N_9476,N_8889,N_8840);
nor U9477 (N_9477,N_8976,N_8929);
xnor U9478 (N_9478,N_8645,N_8761);
or U9479 (N_9479,N_8784,N_8881);
nor U9480 (N_9480,N_8582,N_8760);
and U9481 (N_9481,N_8828,N_8604);
xnor U9482 (N_9482,N_8760,N_8875);
or U9483 (N_9483,N_8759,N_8644);
nor U9484 (N_9484,N_8776,N_8633);
xor U9485 (N_9485,N_8963,N_8565);
nor U9486 (N_9486,N_8881,N_8791);
nand U9487 (N_9487,N_8754,N_8616);
nand U9488 (N_9488,N_8742,N_8445);
or U9489 (N_9489,N_8897,N_8991);
nand U9490 (N_9490,N_8962,N_8427);
nor U9491 (N_9491,N_8738,N_8785);
nand U9492 (N_9492,N_8703,N_8515);
nor U9493 (N_9493,N_8940,N_8721);
xnor U9494 (N_9494,N_8663,N_8486);
nor U9495 (N_9495,N_8511,N_8875);
xnor U9496 (N_9496,N_8484,N_8938);
or U9497 (N_9497,N_8717,N_8581);
xnor U9498 (N_9498,N_8504,N_8768);
xor U9499 (N_9499,N_8883,N_8446);
and U9500 (N_9500,N_8920,N_8938);
xor U9501 (N_9501,N_8471,N_8671);
nor U9502 (N_9502,N_8904,N_8947);
or U9503 (N_9503,N_8571,N_8670);
and U9504 (N_9504,N_8870,N_8450);
nor U9505 (N_9505,N_8764,N_8720);
nand U9506 (N_9506,N_8852,N_8455);
and U9507 (N_9507,N_8579,N_8712);
nand U9508 (N_9508,N_8668,N_8889);
nor U9509 (N_9509,N_8645,N_8837);
or U9510 (N_9510,N_8910,N_8990);
and U9511 (N_9511,N_8600,N_8475);
xnor U9512 (N_9512,N_8786,N_8444);
and U9513 (N_9513,N_8800,N_8714);
xnor U9514 (N_9514,N_8999,N_8448);
xnor U9515 (N_9515,N_8527,N_8569);
nor U9516 (N_9516,N_8978,N_8885);
and U9517 (N_9517,N_8633,N_8959);
or U9518 (N_9518,N_8860,N_8503);
and U9519 (N_9519,N_8965,N_8745);
or U9520 (N_9520,N_8537,N_8732);
nand U9521 (N_9521,N_8544,N_8749);
xor U9522 (N_9522,N_8837,N_8840);
nand U9523 (N_9523,N_8769,N_8488);
or U9524 (N_9524,N_8665,N_8694);
nor U9525 (N_9525,N_8718,N_8711);
nor U9526 (N_9526,N_8701,N_8963);
nand U9527 (N_9527,N_8788,N_8446);
xor U9528 (N_9528,N_8737,N_8928);
nand U9529 (N_9529,N_8762,N_8563);
nand U9530 (N_9530,N_8955,N_8444);
nand U9531 (N_9531,N_8605,N_8432);
nor U9532 (N_9532,N_8411,N_8787);
or U9533 (N_9533,N_8536,N_8663);
nor U9534 (N_9534,N_8518,N_8473);
nand U9535 (N_9535,N_8695,N_8743);
and U9536 (N_9536,N_8817,N_8755);
nand U9537 (N_9537,N_8970,N_8475);
nor U9538 (N_9538,N_8504,N_8612);
xnor U9539 (N_9539,N_8921,N_8595);
nor U9540 (N_9540,N_8886,N_8839);
xor U9541 (N_9541,N_8922,N_8680);
nor U9542 (N_9542,N_8951,N_8787);
nor U9543 (N_9543,N_8898,N_8624);
nand U9544 (N_9544,N_8878,N_8625);
nand U9545 (N_9545,N_8482,N_8767);
and U9546 (N_9546,N_8480,N_8800);
nand U9547 (N_9547,N_8501,N_8992);
and U9548 (N_9548,N_8828,N_8485);
or U9549 (N_9549,N_8503,N_8612);
and U9550 (N_9550,N_8798,N_8739);
and U9551 (N_9551,N_8670,N_8652);
xnor U9552 (N_9552,N_8952,N_8596);
nor U9553 (N_9553,N_8574,N_8801);
and U9554 (N_9554,N_8960,N_8935);
nor U9555 (N_9555,N_8639,N_8472);
or U9556 (N_9556,N_8946,N_8472);
or U9557 (N_9557,N_8580,N_8411);
and U9558 (N_9558,N_8713,N_8927);
xnor U9559 (N_9559,N_8793,N_8768);
nand U9560 (N_9560,N_8528,N_8614);
xnor U9561 (N_9561,N_8739,N_8914);
and U9562 (N_9562,N_8777,N_8413);
or U9563 (N_9563,N_8412,N_8457);
and U9564 (N_9564,N_8968,N_8581);
xor U9565 (N_9565,N_8650,N_8843);
xor U9566 (N_9566,N_8886,N_8897);
nor U9567 (N_9567,N_8558,N_8430);
and U9568 (N_9568,N_8965,N_8568);
or U9569 (N_9569,N_8902,N_8871);
nor U9570 (N_9570,N_8635,N_8549);
nand U9571 (N_9571,N_8862,N_8560);
nand U9572 (N_9572,N_8738,N_8860);
or U9573 (N_9573,N_8526,N_8560);
and U9574 (N_9574,N_8589,N_8724);
nor U9575 (N_9575,N_8580,N_8991);
nor U9576 (N_9576,N_8487,N_8833);
nor U9577 (N_9577,N_8835,N_8523);
nand U9578 (N_9578,N_8863,N_8655);
xor U9579 (N_9579,N_8967,N_8510);
and U9580 (N_9580,N_8501,N_8951);
nor U9581 (N_9581,N_8956,N_8514);
nor U9582 (N_9582,N_8760,N_8822);
and U9583 (N_9583,N_8452,N_8997);
and U9584 (N_9584,N_8812,N_8874);
or U9585 (N_9585,N_8790,N_8621);
nand U9586 (N_9586,N_8955,N_8950);
xor U9587 (N_9587,N_8798,N_8405);
and U9588 (N_9588,N_8991,N_8440);
nand U9589 (N_9589,N_8918,N_8917);
nor U9590 (N_9590,N_8487,N_8808);
or U9591 (N_9591,N_8865,N_8948);
or U9592 (N_9592,N_8458,N_8860);
or U9593 (N_9593,N_8806,N_8854);
xor U9594 (N_9594,N_8428,N_8719);
nor U9595 (N_9595,N_8566,N_8575);
or U9596 (N_9596,N_8879,N_8638);
nand U9597 (N_9597,N_8763,N_8442);
or U9598 (N_9598,N_8665,N_8763);
nor U9599 (N_9599,N_8854,N_8495);
xnor U9600 (N_9600,N_9514,N_9261);
nor U9601 (N_9601,N_9215,N_9035);
nor U9602 (N_9602,N_9445,N_9135);
xor U9603 (N_9603,N_9573,N_9475);
xnor U9604 (N_9604,N_9022,N_9458);
nor U9605 (N_9605,N_9108,N_9251);
nor U9606 (N_9606,N_9304,N_9248);
nor U9607 (N_9607,N_9176,N_9542);
nand U9608 (N_9608,N_9509,N_9260);
or U9609 (N_9609,N_9243,N_9400);
nor U9610 (N_9610,N_9173,N_9491);
nor U9611 (N_9611,N_9012,N_9128);
nand U9612 (N_9612,N_9229,N_9536);
nor U9613 (N_9613,N_9537,N_9231);
and U9614 (N_9614,N_9444,N_9218);
and U9615 (N_9615,N_9438,N_9446);
nor U9616 (N_9616,N_9133,N_9538);
xor U9617 (N_9617,N_9184,N_9004);
nand U9618 (N_9618,N_9158,N_9385);
nor U9619 (N_9619,N_9157,N_9289);
xor U9620 (N_9620,N_9512,N_9520);
xnor U9621 (N_9621,N_9118,N_9353);
nand U9622 (N_9622,N_9003,N_9410);
and U9623 (N_9623,N_9511,N_9120);
and U9624 (N_9624,N_9437,N_9268);
nand U9625 (N_9625,N_9486,N_9221);
xor U9626 (N_9626,N_9171,N_9416);
nand U9627 (N_9627,N_9083,N_9593);
nor U9628 (N_9628,N_9266,N_9162);
nor U9629 (N_9629,N_9153,N_9467);
nand U9630 (N_9630,N_9571,N_9292);
nor U9631 (N_9631,N_9170,N_9177);
nor U9632 (N_9632,N_9129,N_9156);
and U9633 (N_9633,N_9354,N_9039);
nor U9634 (N_9634,N_9345,N_9332);
or U9635 (N_9635,N_9453,N_9029);
and U9636 (N_9636,N_9360,N_9502);
nor U9637 (N_9637,N_9252,N_9399);
xnor U9638 (N_9638,N_9471,N_9355);
nand U9639 (N_9639,N_9054,N_9186);
nor U9640 (N_9640,N_9234,N_9559);
or U9641 (N_9641,N_9506,N_9008);
and U9642 (N_9642,N_9359,N_9487);
and U9643 (N_9643,N_9504,N_9331);
or U9644 (N_9644,N_9356,N_9315);
xor U9645 (N_9645,N_9040,N_9267);
nor U9646 (N_9646,N_9305,N_9216);
nor U9647 (N_9647,N_9097,N_9044);
nand U9648 (N_9648,N_9508,N_9322);
nand U9649 (N_9649,N_9139,N_9333);
xnor U9650 (N_9650,N_9344,N_9068);
nand U9651 (N_9651,N_9207,N_9577);
nand U9652 (N_9652,N_9277,N_9262);
nand U9653 (N_9653,N_9440,N_9518);
xnor U9654 (N_9654,N_9589,N_9429);
and U9655 (N_9655,N_9343,N_9179);
or U9656 (N_9656,N_9510,N_9507);
and U9657 (N_9657,N_9116,N_9235);
nand U9658 (N_9658,N_9154,N_9222);
or U9659 (N_9659,N_9528,N_9288);
or U9660 (N_9660,N_9395,N_9285);
xor U9661 (N_9661,N_9055,N_9497);
nor U9662 (N_9662,N_9013,N_9271);
nor U9663 (N_9663,N_9411,N_9143);
nor U9664 (N_9664,N_9185,N_9392);
nand U9665 (N_9665,N_9591,N_9048);
xnor U9666 (N_9666,N_9334,N_9459);
and U9667 (N_9667,N_9279,N_9505);
nor U9668 (N_9668,N_9152,N_9311);
xor U9669 (N_9669,N_9325,N_9161);
xor U9670 (N_9670,N_9069,N_9348);
nor U9671 (N_9671,N_9023,N_9052);
nand U9672 (N_9672,N_9485,N_9275);
nand U9673 (N_9673,N_9586,N_9599);
or U9674 (N_9674,N_9066,N_9316);
nand U9675 (N_9675,N_9419,N_9373);
nor U9676 (N_9676,N_9532,N_9233);
and U9677 (N_9677,N_9553,N_9451);
and U9678 (N_9678,N_9383,N_9530);
and U9679 (N_9679,N_9110,N_9232);
or U9680 (N_9680,N_9436,N_9025);
and U9681 (N_9681,N_9115,N_9195);
or U9682 (N_9682,N_9551,N_9366);
xnor U9683 (N_9683,N_9312,N_9210);
nor U9684 (N_9684,N_9494,N_9093);
and U9685 (N_9685,N_9405,N_9310);
and U9686 (N_9686,N_9567,N_9001);
nor U9687 (N_9687,N_9295,N_9396);
nand U9688 (N_9688,N_9421,N_9202);
and U9689 (N_9689,N_9543,N_9018);
nor U9690 (N_9690,N_9302,N_9595);
nor U9691 (N_9691,N_9237,N_9560);
and U9692 (N_9692,N_9597,N_9282);
nor U9693 (N_9693,N_9501,N_9492);
or U9694 (N_9694,N_9377,N_9422);
xor U9695 (N_9695,N_9474,N_9329);
or U9696 (N_9696,N_9079,N_9071);
nand U9697 (N_9697,N_9273,N_9375);
nor U9698 (N_9698,N_9030,N_9199);
and U9699 (N_9699,N_9107,N_9140);
nor U9700 (N_9700,N_9317,N_9020);
xor U9701 (N_9701,N_9546,N_9070);
nand U9702 (N_9702,N_9136,N_9059);
nand U9703 (N_9703,N_9481,N_9413);
nand U9704 (N_9704,N_9596,N_9406);
and U9705 (N_9705,N_9371,N_9089);
nor U9706 (N_9706,N_9211,N_9298);
xor U9707 (N_9707,N_9009,N_9137);
nor U9708 (N_9708,N_9341,N_9016);
nand U9709 (N_9709,N_9010,N_9205);
and U9710 (N_9710,N_9223,N_9165);
or U9711 (N_9711,N_9263,N_9208);
xor U9712 (N_9712,N_9303,N_9477);
nand U9713 (N_9713,N_9535,N_9101);
or U9714 (N_9714,N_9236,N_9258);
xor U9715 (N_9715,N_9082,N_9283);
nor U9716 (N_9716,N_9549,N_9558);
nand U9717 (N_9717,N_9014,N_9043);
or U9718 (N_9718,N_9342,N_9575);
nand U9719 (N_9719,N_9121,N_9239);
xnor U9720 (N_9720,N_9397,N_9418);
nand U9721 (N_9721,N_9047,N_9037);
and U9722 (N_9722,N_9188,N_9313);
nand U9723 (N_9723,N_9281,N_9570);
nor U9724 (N_9724,N_9449,N_9072);
xor U9725 (N_9725,N_9306,N_9556);
nand U9726 (N_9726,N_9452,N_9041);
or U9727 (N_9727,N_9096,N_9147);
nor U9728 (N_9728,N_9105,N_9130);
or U9729 (N_9729,N_9579,N_9112);
and U9730 (N_9730,N_9021,N_9454);
or U9731 (N_9731,N_9381,N_9276);
and U9732 (N_9732,N_9301,N_9146);
nor U9733 (N_9733,N_9455,N_9533);
and U9734 (N_9734,N_9376,N_9339);
and U9735 (N_9735,N_9077,N_9521);
or U9736 (N_9736,N_9462,N_9201);
or U9737 (N_9737,N_9431,N_9094);
or U9738 (N_9738,N_9075,N_9464);
and U9739 (N_9739,N_9326,N_9212);
nor U9740 (N_9740,N_9240,N_9046);
and U9741 (N_9741,N_9131,N_9402);
xnor U9742 (N_9742,N_9517,N_9204);
xor U9743 (N_9743,N_9117,N_9472);
or U9744 (N_9744,N_9414,N_9337);
xnor U9745 (N_9745,N_9545,N_9141);
or U9746 (N_9746,N_9335,N_9578);
xor U9747 (N_9747,N_9124,N_9550);
or U9748 (N_9748,N_9382,N_9104);
or U9749 (N_9749,N_9358,N_9006);
nand U9750 (N_9750,N_9374,N_9324);
nand U9751 (N_9751,N_9238,N_9582);
nand U9752 (N_9752,N_9461,N_9319);
and U9753 (N_9753,N_9127,N_9328);
nor U9754 (N_9754,N_9209,N_9388);
nand U9755 (N_9755,N_9194,N_9450);
xnor U9756 (N_9756,N_9142,N_9480);
or U9757 (N_9757,N_9432,N_9198);
xor U9758 (N_9758,N_9484,N_9086);
and U9759 (N_9759,N_9144,N_9123);
and U9760 (N_9760,N_9109,N_9529);
nor U9761 (N_9761,N_9569,N_9524);
xor U9762 (N_9762,N_9338,N_9368);
and U9763 (N_9763,N_9206,N_9420);
xnor U9764 (N_9764,N_9428,N_9193);
nand U9765 (N_9765,N_9378,N_9245);
or U9766 (N_9766,N_9076,N_9554);
nor U9767 (N_9767,N_9056,N_9191);
xnor U9768 (N_9768,N_9427,N_9466);
nor U9769 (N_9769,N_9351,N_9469);
nand U9770 (N_9770,N_9389,N_9005);
or U9771 (N_9771,N_9213,N_9293);
and U9772 (N_9772,N_9307,N_9473);
and U9773 (N_9773,N_9439,N_9095);
and U9774 (N_9774,N_9196,N_9024);
nand U9775 (N_9775,N_9443,N_9036);
nand U9776 (N_9776,N_9042,N_9442);
or U9777 (N_9777,N_9557,N_9253);
or U9778 (N_9778,N_9098,N_9150);
or U9779 (N_9779,N_9028,N_9574);
nand U9780 (N_9780,N_9585,N_9387);
or U9781 (N_9781,N_9594,N_9519);
and U9782 (N_9782,N_9011,N_9361);
xor U9783 (N_9783,N_9463,N_9214);
and U9784 (N_9784,N_9224,N_9490);
and U9785 (N_9785,N_9327,N_9081);
or U9786 (N_9786,N_9180,N_9203);
nor U9787 (N_9787,N_9246,N_9478);
xnor U9788 (N_9788,N_9496,N_9049);
or U9789 (N_9789,N_9085,N_9132);
and U9790 (N_9790,N_9017,N_9190);
or U9791 (N_9791,N_9155,N_9225);
or U9792 (N_9792,N_9363,N_9365);
nor U9793 (N_9793,N_9590,N_9217);
nor U9794 (N_9794,N_9457,N_9178);
xor U9795 (N_9795,N_9031,N_9483);
and U9796 (N_9796,N_9045,N_9362);
nand U9797 (N_9797,N_9027,N_9000);
and U9798 (N_9798,N_9380,N_9297);
nand U9799 (N_9799,N_9227,N_9254);
or U9800 (N_9800,N_9134,N_9526);
nand U9801 (N_9801,N_9495,N_9168);
or U9802 (N_9802,N_9482,N_9367);
nand U9803 (N_9803,N_9565,N_9548);
and U9804 (N_9804,N_9181,N_9465);
and U9805 (N_9805,N_9057,N_9330);
and U9806 (N_9806,N_9113,N_9425);
nand U9807 (N_9807,N_9119,N_9357);
and U9808 (N_9808,N_9552,N_9230);
xnor U9809 (N_9809,N_9084,N_9448);
xor U9810 (N_9810,N_9051,N_9489);
nor U9811 (N_9811,N_9417,N_9587);
nand U9812 (N_9812,N_9200,N_9349);
and U9813 (N_9813,N_9265,N_9287);
or U9814 (N_9814,N_9149,N_9340);
nor U9815 (N_9815,N_9291,N_9159);
xnor U9816 (N_9816,N_9401,N_9308);
or U9817 (N_9817,N_9269,N_9092);
nor U9818 (N_9818,N_9409,N_9412);
or U9819 (N_9819,N_9309,N_9106);
xnor U9820 (N_9820,N_9540,N_9228);
nor U9821 (N_9821,N_9568,N_9584);
nand U9822 (N_9822,N_9192,N_9102);
nand U9823 (N_9823,N_9061,N_9278);
nand U9824 (N_9824,N_9296,N_9167);
or U9825 (N_9825,N_9053,N_9323);
xnor U9826 (N_9826,N_9257,N_9272);
xnor U9827 (N_9827,N_9062,N_9280);
nand U9828 (N_9828,N_9415,N_9270);
nor U9829 (N_9829,N_9122,N_9468);
nor U9830 (N_9830,N_9347,N_9197);
nor U9831 (N_9831,N_9247,N_9534);
or U9832 (N_9832,N_9423,N_9060);
nand U9833 (N_9833,N_9088,N_9390);
and U9834 (N_9834,N_9434,N_9433);
nor U9835 (N_9835,N_9516,N_9090);
nand U9836 (N_9836,N_9346,N_9050);
or U9837 (N_9837,N_9493,N_9065);
or U9838 (N_9838,N_9407,N_9539);
or U9839 (N_9839,N_9476,N_9163);
nand U9840 (N_9840,N_9259,N_9099);
nand U9841 (N_9841,N_9138,N_9370);
nand U9842 (N_9842,N_9002,N_9404);
xnor U9843 (N_9843,N_9256,N_9561);
or U9844 (N_9844,N_9126,N_9441);
nand U9845 (N_9845,N_9034,N_9320);
or U9846 (N_9846,N_9074,N_9350);
nor U9847 (N_9847,N_9015,N_9581);
or U9848 (N_9848,N_9125,N_9284);
xnor U9849 (N_9849,N_9576,N_9073);
xnor U9850 (N_9850,N_9588,N_9114);
and U9851 (N_9851,N_9364,N_9562);
xor U9852 (N_9852,N_9166,N_9372);
or U9853 (N_9853,N_9564,N_9523);
and U9854 (N_9854,N_9032,N_9274);
and U9855 (N_9855,N_9583,N_9183);
xnor U9856 (N_9856,N_9299,N_9544);
or U9857 (N_9857,N_9541,N_9498);
or U9858 (N_9858,N_9531,N_9182);
nand U9859 (N_9859,N_9386,N_9063);
nor U9860 (N_9860,N_9169,N_9525);
nand U9861 (N_9861,N_9408,N_9007);
and U9862 (N_9862,N_9087,N_9566);
xor U9863 (N_9863,N_9067,N_9488);
or U9864 (N_9864,N_9189,N_9435);
or U9865 (N_9865,N_9187,N_9160);
and U9866 (N_9866,N_9290,N_9175);
nand U9867 (N_9867,N_9555,N_9352);
xor U9868 (N_9868,N_9148,N_9580);
xor U9869 (N_9869,N_9255,N_9151);
nor U9870 (N_9870,N_9522,N_9447);
or U9871 (N_9871,N_9294,N_9430);
or U9872 (N_9872,N_9563,N_9172);
and U9873 (N_9873,N_9572,N_9091);
nor U9874 (N_9874,N_9164,N_9424);
nor U9875 (N_9875,N_9527,N_9379);
xor U9876 (N_9876,N_9300,N_9145);
nor U9877 (N_9877,N_9515,N_9314);
nor U9878 (N_9878,N_9391,N_9503);
nor U9879 (N_9879,N_9242,N_9321);
xnor U9880 (N_9880,N_9369,N_9460);
and U9881 (N_9881,N_9264,N_9033);
nor U9882 (N_9882,N_9038,N_9547);
xnor U9883 (N_9883,N_9219,N_9384);
and U9884 (N_9884,N_9479,N_9286);
xnor U9885 (N_9885,N_9111,N_9174);
or U9886 (N_9886,N_9249,N_9336);
or U9887 (N_9887,N_9220,N_9241);
nand U9888 (N_9888,N_9078,N_9403);
nand U9889 (N_9889,N_9244,N_9318);
or U9890 (N_9890,N_9499,N_9250);
nand U9891 (N_9891,N_9058,N_9500);
and U9892 (N_9892,N_9100,N_9103);
and U9893 (N_9893,N_9064,N_9456);
or U9894 (N_9894,N_9470,N_9513);
xor U9895 (N_9895,N_9026,N_9394);
or U9896 (N_9896,N_9426,N_9080);
nor U9897 (N_9897,N_9592,N_9226);
xor U9898 (N_9898,N_9398,N_9598);
xor U9899 (N_9899,N_9393,N_9019);
nand U9900 (N_9900,N_9146,N_9508);
nor U9901 (N_9901,N_9024,N_9348);
and U9902 (N_9902,N_9122,N_9156);
and U9903 (N_9903,N_9472,N_9146);
nor U9904 (N_9904,N_9140,N_9367);
nor U9905 (N_9905,N_9019,N_9348);
or U9906 (N_9906,N_9011,N_9425);
nand U9907 (N_9907,N_9450,N_9083);
xor U9908 (N_9908,N_9400,N_9030);
nand U9909 (N_9909,N_9547,N_9391);
xor U9910 (N_9910,N_9346,N_9254);
nand U9911 (N_9911,N_9252,N_9419);
nor U9912 (N_9912,N_9027,N_9332);
and U9913 (N_9913,N_9561,N_9123);
nand U9914 (N_9914,N_9296,N_9364);
nor U9915 (N_9915,N_9242,N_9519);
and U9916 (N_9916,N_9432,N_9148);
nand U9917 (N_9917,N_9471,N_9121);
or U9918 (N_9918,N_9469,N_9171);
and U9919 (N_9919,N_9588,N_9098);
nand U9920 (N_9920,N_9260,N_9501);
nand U9921 (N_9921,N_9027,N_9531);
nor U9922 (N_9922,N_9571,N_9106);
nand U9923 (N_9923,N_9379,N_9556);
and U9924 (N_9924,N_9369,N_9033);
nor U9925 (N_9925,N_9572,N_9285);
nor U9926 (N_9926,N_9184,N_9501);
and U9927 (N_9927,N_9037,N_9301);
nor U9928 (N_9928,N_9097,N_9563);
nand U9929 (N_9929,N_9527,N_9534);
xor U9930 (N_9930,N_9305,N_9150);
nor U9931 (N_9931,N_9214,N_9376);
xor U9932 (N_9932,N_9425,N_9124);
nand U9933 (N_9933,N_9512,N_9503);
and U9934 (N_9934,N_9277,N_9458);
xnor U9935 (N_9935,N_9123,N_9169);
nand U9936 (N_9936,N_9543,N_9457);
nand U9937 (N_9937,N_9290,N_9041);
nand U9938 (N_9938,N_9101,N_9326);
xor U9939 (N_9939,N_9190,N_9253);
xor U9940 (N_9940,N_9490,N_9104);
or U9941 (N_9941,N_9522,N_9256);
nor U9942 (N_9942,N_9494,N_9144);
nand U9943 (N_9943,N_9366,N_9545);
nor U9944 (N_9944,N_9246,N_9311);
nor U9945 (N_9945,N_9368,N_9559);
nor U9946 (N_9946,N_9467,N_9057);
or U9947 (N_9947,N_9374,N_9032);
nor U9948 (N_9948,N_9139,N_9284);
and U9949 (N_9949,N_9181,N_9132);
nand U9950 (N_9950,N_9067,N_9143);
or U9951 (N_9951,N_9329,N_9224);
xor U9952 (N_9952,N_9140,N_9269);
nor U9953 (N_9953,N_9472,N_9173);
nand U9954 (N_9954,N_9580,N_9123);
nand U9955 (N_9955,N_9570,N_9145);
xor U9956 (N_9956,N_9114,N_9243);
nor U9957 (N_9957,N_9349,N_9177);
or U9958 (N_9958,N_9431,N_9136);
and U9959 (N_9959,N_9581,N_9034);
and U9960 (N_9960,N_9199,N_9372);
nand U9961 (N_9961,N_9287,N_9052);
nor U9962 (N_9962,N_9212,N_9173);
and U9963 (N_9963,N_9308,N_9559);
and U9964 (N_9964,N_9337,N_9552);
and U9965 (N_9965,N_9128,N_9161);
nand U9966 (N_9966,N_9028,N_9532);
nor U9967 (N_9967,N_9269,N_9370);
nor U9968 (N_9968,N_9223,N_9355);
nand U9969 (N_9969,N_9100,N_9525);
nand U9970 (N_9970,N_9441,N_9058);
and U9971 (N_9971,N_9387,N_9298);
nor U9972 (N_9972,N_9344,N_9304);
and U9973 (N_9973,N_9088,N_9179);
or U9974 (N_9974,N_9467,N_9061);
and U9975 (N_9975,N_9401,N_9411);
or U9976 (N_9976,N_9134,N_9447);
xnor U9977 (N_9977,N_9082,N_9238);
xor U9978 (N_9978,N_9505,N_9022);
or U9979 (N_9979,N_9288,N_9072);
and U9980 (N_9980,N_9279,N_9417);
nor U9981 (N_9981,N_9090,N_9535);
nand U9982 (N_9982,N_9111,N_9171);
nor U9983 (N_9983,N_9291,N_9150);
nor U9984 (N_9984,N_9149,N_9121);
nand U9985 (N_9985,N_9333,N_9072);
xor U9986 (N_9986,N_9417,N_9132);
nand U9987 (N_9987,N_9098,N_9587);
xnor U9988 (N_9988,N_9267,N_9280);
nand U9989 (N_9989,N_9195,N_9367);
nand U9990 (N_9990,N_9480,N_9070);
and U9991 (N_9991,N_9217,N_9136);
xnor U9992 (N_9992,N_9120,N_9037);
nand U9993 (N_9993,N_9080,N_9323);
xnor U9994 (N_9994,N_9544,N_9520);
nand U9995 (N_9995,N_9010,N_9536);
or U9996 (N_9996,N_9173,N_9559);
or U9997 (N_9997,N_9530,N_9126);
nand U9998 (N_9998,N_9237,N_9185);
nor U9999 (N_9999,N_9390,N_9191);
nor U10000 (N_10000,N_9403,N_9446);
or U10001 (N_10001,N_9460,N_9185);
or U10002 (N_10002,N_9007,N_9252);
or U10003 (N_10003,N_9082,N_9568);
nor U10004 (N_10004,N_9331,N_9176);
nor U10005 (N_10005,N_9324,N_9575);
nand U10006 (N_10006,N_9003,N_9271);
or U10007 (N_10007,N_9235,N_9041);
and U10008 (N_10008,N_9461,N_9450);
nand U10009 (N_10009,N_9377,N_9426);
nor U10010 (N_10010,N_9138,N_9212);
xor U10011 (N_10011,N_9007,N_9020);
or U10012 (N_10012,N_9582,N_9376);
nand U10013 (N_10013,N_9539,N_9324);
and U10014 (N_10014,N_9389,N_9188);
nor U10015 (N_10015,N_9292,N_9099);
nor U10016 (N_10016,N_9130,N_9092);
nand U10017 (N_10017,N_9209,N_9404);
and U10018 (N_10018,N_9117,N_9295);
and U10019 (N_10019,N_9089,N_9540);
nand U10020 (N_10020,N_9042,N_9295);
nor U10021 (N_10021,N_9538,N_9526);
or U10022 (N_10022,N_9069,N_9514);
xor U10023 (N_10023,N_9562,N_9115);
or U10024 (N_10024,N_9231,N_9508);
xor U10025 (N_10025,N_9507,N_9431);
nand U10026 (N_10026,N_9208,N_9438);
nor U10027 (N_10027,N_9557,N_9121);
nand U10028 (N_10028,N_9322,N_9506);
or U10029 (N_10029,N_9149,N_9206);
and U10030 (N_10030,N_9572,N_9551);
xor U10031 (N_10031,N_9322,N_9373);
nor U10032 (N_10032,N_9311,N_9300);
nand U10033 (N_10033,N_9561,N_9223);
xor U10034 (N_10034,N_9115,N_9323);
nor U10035 (N_10035,N_9373,N_9580);
xnor U10036 (N_10036,N_9300,N_9180);
nand U10037 (N_10037,N_9218,N_9071);
and U10038 (N_10038,N_9551,N_9257);
nor U10039 (N_10039,N_9016,N_9271);
and U10040 (N_10040,N_9502,N_9228);
and U10041 (N_10041,N_9455,N_9244);
or U10042 (N_10042,N_9017,N_9476);
and U10043 (N_10043,N_9026,N_9368);
nor U10044 (N_10044,N_9153,N_9196);
nor U10045 (N_10045,N_9055,N_9201);
and U10046 (N_10046,N_9342,N_9597);
nand U10047 (N_10047,N_9276,N_9137);
nand U10048 (N_10048,N_9207,N_9336);
and U10049 (N_10049,N_9454,N_9077);
nor U10050 (N_10050,N_9075,N_9306);
or U10051 (N_10051,N_9424,N_9504);
nor U10052 (N_10052,N_9534,N_9280);
xor U10053 (N_10053,N_9548,N_9116);
nor U10054 (N_10054,N_9008,N_9259);
nor U10055 (N_10055,N_9114,N_9327);
nand U10056 (N_10056,N_9452,N_9130);
xor U10057 (N_10057,N_9273,N_9042);
or U10058 (N_10058,N_9543,N_9166);
nand U10059 (N_10059,N_9184,N_9012);
nor U10060 (N_10060,N_9054,N_9480);
nor U10061 (N_10061,N_9316,N_9006);
xnor U10062 (N_10062,N_9399,N_9008);
xor U10063 (N_10063,N_9558,N_9518);
nand U10064 (N_10064,N_9119,N_9434);
or U10065 (N_10065,N_9135,N_9270);
nor U10066 (N_10066,N_9416,N_9551);
xor U10067 (N_10067,N_9570,N_9531);
nand U10068 (N_10068,N_9452,N_9405);
xnor U10069 (N_10069,N_9414,N_9515);
nor U10070 (N_10070,N_9050,N_9357);
xor U10071 (N_10071,N_9033,N_9336);
nand U10072 (N_10072,N_9376,N_9348);
nand U10073 (N_10073,N_9474,N_9094);
nand U10074 (N_10074,N_9076,N_9462);
nor U10075 (N_10075,N_9531,N_9473);
and U10076 (N_10076,N_9239,N_9302);
nor U10077 (N_10077,N_9230,N_9524);
nand U10078 (N_10078,N_9562,N_9134);
and U10079 (N_10079,N_9566,N_9221);
and U10080 (N_10080,N_9425,N_9060);
xnor U10081 (N_10081,N_9103,N_9005);
nand U10082 (N_10082,N_9048,N_9282);
and U10083 (N_10083,N_9085,N_9310);
or U10084 (N_10084,N_9232,N_9323);
nand U10085 (N_10085,N_9423,N_9159);
and U10086 (N_10086,N_9095,N_9570);
nor U10087 (N_10087,N_9401,N_9300);
xor U10088 (N_10088,N_9531,N_9215);
xnor U10089 (N_10089,N_9545,N_9276);
or U10090 (N_10090,N_9107,N_9057);
nor U10091 (N_10091,N_9253,N_9008);
and U10092 (N_10092,N_9462,N_9347);
or U10093 (N_10093,N_9543,N_9328);
xnor U10094 (N_10094,N_9512,N_9436);
and U10095 (N_10095,N_9088,N_9035);
nand U10096 (N_10096,N_9308,N_9579);
nand U10097 (N_10097,N_9378,N_9246);
or U10098 (N_10098,N_9044,N_9324);
or U10099 (N_10099,N_9189,N_9267);
nand U10100 (N_10100,N_9456,N_9429);
nand U10101 (N_10101,N_9516,N_9483);
nor U10102 (N_10102,N_9414,N_9202);
or U10103 (N_10103,N_9494,N_9099);
nand U10104 (N_10104,N_9117,N_9176);
xor U10105 (N_10105,N_9533,N_9110);
xor U10106 (N_10106,N_9065,N_9494);
nand U10107 (N_10107,N_9365,N_9595);
or U10108 (N_10108,N_9053,N_9449);
nor U10109 (N_10109,N_9129,N_9136);
nor U10110 (N_10110,N_9053,N_9244);
nand U10111 (N_10111,N_9066,N_9362);
and U10112 (N_10112,N_9594,N_9571);
nor U10113 (N_10113,N_9098,N_9580);
or U10114 (N_10114,N_9136,N_9593);
or U10115 (N_10115,N_9279,N_9154);
or U10116 (N_10116,N_9339,N_9210);
and U10117 (N_10117,N_9257,N_9156);
or U10118 (N_10118,N_9533,N_9566);
nor U10119 (N_10119,N_9480,N_9161);
and U10120 (N_10120,N_9486,N_9180);
nor U10121 (N_10121,N_9031,N_9211);
xnor U10122 (N_10122,N_9389,N_9425);
and U10123 (N_10123,N_9276,N_9108);
nor U10124 (N_10124,N_9164,N_9379);
nand U10125 (N_10125,N_9585,N_9013);
or U10126 (N_10126,N_9148,N_9187);
nor U10127 (N_10127,N_9529,N_9020);
xor U10128 (N_10128,N_9449,N_9330);
or U10129 (N_10129,N_9194,N_9441);
nor U10130 (N_10130,N_9333,N_9101);
xor U10131 (N_10131,N_9097,N_9597);
nor U10132 (N_10132,N_9001,N_9513);
and U10133 (N_10133,N_9304,N_9404);
nand U10134 (N_10134,N_9554,N_9283);
nor U10135 (N_10135,N_9117,N_9411);
or U10136 (N_10136,N_9057,N_9128);
and U10137 (N_10137,N_9362,N_9109);
nand U10138 (N_10138,N_9333,N_9350);
nand U10139 (N_10139,N_9445,N_9589);
nand U10140 (N_10140,N_9384,N_9466);
or U10141 (N_10141,N_9413,N_9337);
and U10142 (N_10142,N_9460,N_9550);
nand U10143 (N_10143,N_9076,N_9327);
nor U10144 (N_10144,N_9248,N_9393);
or U10145 (N_10145,N_9505,N_9065);
and U10146 (N_10146,N_9255,N_9541);
or U10147 (N_10147,N_9402,N_9516);
nor U10148 (N_10148,N_9544,N_9150);
nand U10149 (N_10149,N_9158,N_9116);
xnor U10150 (N_10150,N_9404,N_9456);
and U10151 (N_10151,N_9420,N_9048);
and U10152 (N_10152,N_9457,N_9504);
nor U10153 (N_10153,N_9083,N_9059);
and U10154 (N_10154,N_9308,N_9304);
and U10155 (N_10155,N_9432,N_9204);
or U10156 (N_10156,N_9196,N_9201);
or U10157 (N_10157,N_9477,N_9261);
nand U10158 (N_10158,N_9280,N_9195);
or U10159 (N_10159,N_9347,N_9200);
nor U10160 (N_10160,N_9237,N_9328);
nor U10161 (N_10161,N_9101,N_9348);
nand U10162 (N_10162,N_9328,N_9440);
xnor U10163 (N_10163,N_9587,N_9585);
and U10164 (N_10164,N_9080,N_9550);
nor U10165 (N_10165,N_9441,N_9546);
nand U10166 (N_10166,N_9535,N_9450);
and U10167 (N_10167,N_9298,N_9246);
and U10168 (N_10168,N_9595,N_9540);
and U10169 (N_10169,N_9388,N_9495);
and U10170 (N_10170,N_9309,N_9161);
nor U10171 (N_10171,N_9294,N_9453);
xor U10172 (N_10172,N_9503,N_9035);
and U10173 (N_10173,N_9453,N_9159);
xnor U10174 (N_10174,N_9496,N_9030);
nor U10175 (N_10175,N_9261,N_9517);
and U10176 (N_10176,N_9473,N_9288);
and U10177 (N_10177,N_9046,N_9234);
and U10178 (N_10178,N_9310,N_9089);
nor U10179 (N_10179,N_9216,N_9346);
nand U10180 (N_10180,N_9445,N_9370);
nor U10181 (N_10181,N_9570,N_9519);
xnor U10182 (N_10182,N_9329,N_9451);
xor U10183 (N_10183,N_9440,N_9456);
xor U10184 (N_10184,N_9173,N_9571);
nor U10185 (N_10185,N_9338,N_9476);
nor U10186 (N_10186,N_9177,N_9475);
nand U10187 (N_10187,N_9394,N_9287);
nor U10188 (N_10188,N_9271,N_9417);
nand U10189 (N_10189,N_9233,N_9063);
nand U10190 (N_10190,N_9515,N_9535);
or U10191 (N_10191,N_9332,N_9409);
nand U10192 (N_10192,N_9032,N_9598);
nor U10193 (N_10193,N_9251,N_9163);
xor U10194 (N_10194,N_9211,N_9076);
or U10195 (N_10195,N_9550,N_9202);
and U10196 (N_10196,N_9202,N_9167);
and U10197 (N_10197,N_9144,N_9431);
nand U10198 (N_10198,N_9276,N_9284);
xnor U10199 (N_10199,N_9088,N_9037);
xnor U10200 (N_10200,N_10079,N_10129);
and U10201 (N_10201,N_9801,N_10103);
or U10202 (N_10202,N_10154,N_10075);
nor U10203 (N_10203,N_9779,N_10110);
xnor U10204 (N_10204,N_9617,N_10160);
xnor U10205 (N_10205,N_9997,N_9657);
xnor U10206 (N_10206,N_9712,N_9842);
xor U10207 (N_10207,N_10050,N_9609);
nand U10208 (N_10208,N_9631,N_9690);
nand U10209 (N_10209,N_9839,N_9887);
nor U10210 (N_10210,N_9820,N_10109);
and U10211 (N_10211,N_9787,N_10010);
nor U10212 (N_10212,N_9770,N_9974);
or U10213 (N_10213,N_10062,N_9760);
nor U10214 (N_10214,N_9727,N_10053);
or U10215 (N_10215,N_9741,N_10040);
and U10216 (N_10216,N_9722,N_9841);
nor U10217 (N_10217,N_9908,N_9999);
nand U10218 (N_10218,N_9715,N_9894);
or U10219 (N_10219,N_9647,N_9638);
nand U10220 (N_10220,N_9896,N_9828);
or U10221 (N_10221,N_10164,N_9680);
nand U10222 (N_10222,N_10004,N_10174);
xor U10223 (N_10223,N_10074,N_9718);
nand U10224 (N_10224,N_9853,N_10030);
xnor U10225 (N_10225,N_9642,N_9866);
or U10226 (N_10226,N_9794,N_9859);
and U10227 (N_10227,N_10149,N_9624);
nand U10228 (N_10228,N_10019,N_10131);
xnor U10229 (N_10229,N_10167,N_9869);
xnor U10230 (N_10230,N_9704,N_9683);
nand U10231 (N_10231,N_10108,N_9792);
xor U10232 (N_10232,N_9876,N_10195);
nand U10233 (N_10233,N_9943,N_9755);
nor U10234 (N_10234,N_9873,N_9738);
and U10235 (N_10235,N_9714,N_10151);
or U10236 (N_10236,N_9976,N_9996);
nor U10237 (N_10237,N_9815,N_9716);
nand U10238 (N_10238,N_9605,N_9721);
or U10239 (N_10239,N_9856,N_9670);
or U10240 (N_10240,N_10033,N_9667);
xnor U10241 (N_10241,N_9602,N_10141);
nand U10242 (N_10242,N_10139,N_9658);
and U10243 (N_10243,N_9991,N_9753);
or U10244 (N_10244,N_9942,N_10014);
nand U10245 (N_10245,N_10048,N_9860);
or U10246 (N_10246,N_10076,N_10112);
and U10247 (N_10247,N_9745,N_9799);
and U10248 (N_10248,N_10016,N_10156);
and U10249 (N_10249,N_9899,N_9987);
xor U10250 (N_10250,N_10182,N_9838);
nand U10251 (N_10251,N_10184,N_9634);
nor U10252 (N_10252,N_9886,N_10021);
xor U10253 (N_10253,N_9699,N_9954);
xor U10254 (N_10254,N_10080,N_10022);
or U10255 (N_10255,N_9622,N_10063);
nand U10256 (N_10256,N_10084,N_9831);
xnor U10257 (N_10257,N_9728,N_9880);
nand U10258 (N_10258,N_9879,N_10122);
or U10259 (N_10259,N_9808,N_9855);
or U10260 (N_10260,N_9928,N_9772);
xnor U10261 (N_10261,N_9972,N_9965);
or U10262 (N_10262,N_10024,N_9837);
nand U10263 (N_10263,N_9906,N_9726);
or U10264 (N_10264,N_9958,N_9751);
xnor U10265 (N_10265,N_9893,N_9659);
and U10266 (N_10266,N_10013,N_9615);
or U10267 (N_10267,N_10070,N_9688);
nor U10268 (N_10268,N_9871,N_10178);
xnor U10269 (N_10269,N_9710,N_9775);
or U10270 (N_10270,N_9832,N_9867);
or U10271 (N_10271,N_10100,N_9700);
or U10272 (N_10272,N_9730,N_9884);
xnor U10273 (N_10273,N_9606,N_9697);
or U10274 (N_10274,N_9931,N_9790);
xnor U10275 (N_10275,N_9907,N_9858);
nor U10276 (N_10276,N_9628,N_10085);
nor U10277 (N_10277,N_10197,N_9824);
nor U10278 (N_10278,N_9817,N_9619);
and U10279 (N_10279,N_10196,N_9982);
xor U10280 (N_10280,N_9909,N_10126);
nor U10281 (N_10281,N_9696,N_10009);
nand U10282 (N_10282,N_10017,N_9960);
or U10283 (N_10283,N_9949,N_9917);
nand U10284 (N_10284,N_10169,N_10157);
or U10285 (N_10285,N_9735,N_9967);
or U10286 (N_10286,N_9635,N_9849);
nor U10287 (N_10287,N_9800,N_10065);
nand U10288 (N_10288,N_9885,N_10003);
nor U10289 (N_10289,N_9834,N_10115);
or U10290 (N_10290,N_10092,N_9707);
and U10291 (N_10291,N_9663,N_9633);
xnor U10292 (N_10292,N_10029,N_9846);
and U10293 (N_10293,N_9969,N_9782);
nand U10294 (N_10294,N_9698,N_9951);
nand U10295 (N_10295,N_9980,N_9694);
xor U10296 (N_10296,N_10034,N_9780);
or U10297 (N_10297,N_9924,N_10026);
or U10298 (N_10298,N_9665,N_9798);
or U10299 (N_10299,N_9840,N_9978);
nand U10300 (N_10300,N_10189,N_10027);
nand U10301 (N_10301,N_9881,N_10068);
nand U10302 (N_10302,N_10000,N_9851);
xor U10303 (N_10303,N_10138,N_10199);
nor U10304 (N_10304,N_9783,N_10105);
nor U10305 (N_10305,N_9705,N_9636);
and U10306 (N_10306,N_9927,N_10173);
or U10307 (N_10307,N_10163,N_9903);
and U10308 (N_10308,N_10037,N_9744);
nand U10309 (N_10309,N_9850,N_9898);
nor U10310 (N_10310,N_9795,N_9711);
nand U10311 (N_10311,N_10159,N_9891);
nand U10312 (N_10312,N_10175,N_10165);
and U10313 (N_10313,N_9904,N_9748);
and U10314 (N_10314,N_9649,N_9607);
nand U10315 (N_10315,N_9754,N_9797);
or U10316 (N_10316,N_9939,N_9702);
or U10317 (N_10317,N_9673,N_10134);
nor U10318 (N_10318,N_9764,N_10020);
nand U10319 (N_10319,N_9901,N_10036);
nand U10320 (N_10320,N_10166,N_9731);
nand U10321 (N_10321,N_9910,N_10116);
or U10322 (N_10322,N_9825,N_9981);
nor U10323 (N_10323,N_9938,N_9740);
nor U10324 (N_10324,N_9778,N_9814);
or U10325 (N_10325,N_9749,N_9941);
or U10326 (N_10326,N_10125,N_9957);
xor U10327 (N_10327,N_10140,N_9864);
and U10328 (N_10328,N_10055,N_10054);
xor U10329 (N_10329,N_10176,N_9785);
nand U10330 (N_10330,N_9979,N_9672);
nor U10331 (N_10331,N_10090,N_10077);
xor U10332 (N_10332,N_9933,N_9805);
and U10333 (N_10333,N_9713,N_9720);
xnor U10334 (N_10334,N_9630,N_9878);
and U10335 (N_10335,N_9791,N_9668);
nor U10336 (N_10336,N_9693,N_10011);
xor U10337 (N_10337,N_9925,N_9905);
nand U10338 (N_10338,N_9811,N_9623);
nand U10339 (N_10339,N_9664,N_10143);
nor U10340 (N_10340,N_9948,N_9747);
or U10341 (N_10341,N_9883,N_10046);
nor U10342 (N_10342,N_9882,N_10051);
nand U10343 (N_10343,N_9998,N_9926);
and U10344 (N_10344,N_9626,N_9956);
and U10345 (N_10345,N_9955,N_10114);
and U10346 (N_10346,N_9613,N_9645);
nand U10347 (N_10347,N_9810,N_9776);
xor U10348 (N_10348,N_10191,N_10007);
xor U10349 (N_10349,N_9816,N_10128);
and U10350 (N_10350,N_10018,N_9788);
or U10351 (N_10351,N_9639,N_9681);
and U10352 (N_10352,N_9889,N_9802);
nand U10353 (N_10353,N_9654,N_9687);
xnor U10354 (N_10354,N_9734,N_9603);
or U10355 (N_10355,N_9874,N_10072);
and U10356 (N_10356,N_9652,N_9915);
and U10357 (N_10357,N_10015,N_9641);
nand U10358 (N_10358,N_10111,N_10031);
xor U10359 (N_10359,N_9923,N_9861);
nand U10360 (N_10360,N_10104,N_9868);
nor U10361 (N_10361,N_9691,N_10177);
or U10362 (N_10362,N_9935,N_10047);
and U10363 (N_10363,N_9608,N_10168);
nor U10364 (N_10364,N_9822,N_10142);
and U10365 (N_10365,N_9766,N_9872);
or U10366 (N_10366,N_9723,N_10102);
or U10367 (N_10367,N_10064,N_10137);
or U10368 (N_10368,N_9632,N_9675);
and U10369 (N_10369,N_9806,N_9655);
nand U10370 (N_10370,N_9769,N_10190);
nor U10371 (N_10371,N_10059,N_9701);
xnor U10372 (N_10372,N_9719,N_9643);
nand U10373 (N_10373,N_10098,N_10198);
nor U10374 (N_10374,N_10005,N_10023);
or U10375 (N_10375,N_9685,N_9934);
nand U10376 (N_10376,N_9804,N_10188);
xor U10377 (N_10377,N_9945,N_9848);
nor U10378 (N_10378,N_9875,N_9765);
and U10379 (N_10379,N_10094,N_9692);
nor U10380 (N_10380,N_9821,N_9758);
nand U10381 (N_10381,N_10086,N_9729);
xnor U10382 (N_10382,N_9950,N_9988);
xnor U10383 (N_10383,N_9600,N_9959);
xor U10384 (N_10384,N_9920,N_9992);
or U10385 (N_10385,N_9812,N_9819);
nor U10386 (N_10386,N_10130,N_9739);
or U10387 (N_10387,N_9971,N_9995);
nand U10388 (N_10388,N_9737,N_9897);
nor U10389 (N_10389,N_9611,N_10161);
nor U10390 (N_10390,N_9621,N_9977);
nor U10391 (N_10391,N_10193,N_9768);
nor U10392 (N_10392,N_9852,N_9830);
nand U10393 (N_10393,N_9646,N_9777);
xor U10394 (N_10394,N_10043,N_10186);
or U10395 (N_10395,N_10192,N_9627);
nor U10396 (N_10396,N_9984,N_9743);
and U10397 (N_10397,N_10042,N_10069);
or U10398 (N_10398,N_9914,N_9733);
xnor U10399 (N_10399,N_10106,N_10136);
and U10400 (N_10400,N_10038,N_9650);
nor U10401 (N_10401,N_10071,N_9989);
xnor U10402 (N_10402,N_9676,N_9836);
or U10403 (N_10403,N_10060,N_10119);
xnor U10404 (N_10404,N_10025,N_9807);
xor U10405 (N_10405,N_9656,N_9862);
or U10406 (N_10406,N_10185,N_9932);
nand U10407 (N_10407,N_10127,N_10133);
nor U10408 (N_10408,N_9786,N_9666);
nand U10409 (N_10409,N_10170,N_9990);
nor U10410 (N_10410,N_9604,N_9781);
nand U10411 (N_10411,N_9684,N_9661);
nor U10412 (N_10412,N_9847,N_9662);
xnor U10413 (N_10413,N_10172,N_10179);
nand U10414 (N_10414,N_10162,N_9946);
xor U10415 (N_10415,N_9809,N_10183);
nand U10416 (N_10416,N_10120,N_10044);
nand U10417 (N_10417,N_9703,N_10082);
and U10418 (N_10418,N_10008,N_9618);
or U10419 (N_10419,N_9913,N_9625);
and U10420 (N_10420,N_10073,N_10095);
or U10421 (N_10421,N_9961,N_10132);
xnor U10422 (N_10422,N_9784,N_9826);
nand U10423 (N_10423,N_10001,N_9877);
nand U10424 (N_10424,N_9612,N_9963);
xor U10425 (N_10425,N_9911,N_9912);
nor U10426 (N_10426,N_10093,N_9944);
and U10427 (N_10427,N_9763,N_9922);
and U10428 (N_10428,N_9660,N_10089);
and U10429 (N_10429,N_9671,N_9742);
and U10430 (N_10430,N_9900,N_9892);
nor U10431 (N_10431,N_9863,N_9921);
or U10432 (N_10432,N_9844,N_9601);
nor U10433 (N_10433,N_9833,N_9796);
and U10434 (N_10434,N_9610,N_9724);
and U10435 (N_10435,N_10056,N_9653);
or U10436 (N_10436,N_10087,N_9962);
xor U10437 (N_10437,N_9964,N_10123);
xnor U10438 (N_10438,N_10153,N_9679);
and U10439 (N_10439,N_9973,N_9870);
or U10440 (N_10440,N_9857,N_9829);
and U10441 (N_10441,N_9651,N_10187);
and U10442 (N_10442,N_10045,N_10107);
and U10443 (N_10443,N_9970,N_10152);
nand U10444 (N_10444,N_9890,N_10099);
nand U10445 (N_10445,N_9953,N_9637);
nor U10446 (N_10446,N_10028,N_10083);
and U10447 (N_10447,N_10121,N_9678);
or U10448 (N_10448,N_9916,N_9752);
nor U10449 (N_10449,N_10118,N_10158);
xnor U10450 (N_10450,N_9640,N_10006);
xor U10451 (N_10451,N_10147,N_10148);
xor U10452 (N_10452,N_9708,N_9736);
or U10453 (N_10453,N_9682,N_9929);
nand U10454 (N_10454,N_9746,N_9648);
or U10455 (N_10455,N_10171,N_9975);
nor U10456 (N_10456,N_9620,N_10058);
xor U10457 (N_10457,N_9614,N_9669);
or U10458 (N_10458,N_9725,N_10144);
nor U10459 (N_10459,N_9843,N_9644);
nand U10460 (N_10460,N_9757,N_9709);
nor U10461 (N_10461,N_10041,N_10081);
or U10462 (N_10462,N_9823,N_9674);
nand U10463 (N_10463,N_9968,N_9994);
nor U10464 (N_10464,N_10002,N_10155);
xor U10465 (N_10465,N_10067,N_10096);
nor U10466 (N_10466,N_10135,N_10146);
or U10467 (N_10467,N_9952,N_9983);
or U10468 (N_10468,N_9818,N_10012);
xor U10469 (N_10469,N_9918,N_9732);
and U10470 (N_10470,N_9761,N_10049);
or U10471 (N_10471,N_9888,N_10066);
and U10472 (N_10472,N_10057,N_10088);
nand U10473 (N_10473,N_9793,N_9827);
nand U10474 (N_10474,N_9774,N_9937);
or U10475 (N_10475,N_9756,N_9773);
or U10476 (N_10476,N_9986,N_9940);
nand U10477 (N_10477,N_9919,N_9686);
and U10478 (N_10478,N_9677,N_10117);
or U10479 (N_10479,N_9689,N_9803);
xnor U10480 (N_10480,N_9966,N_10035);
and U10481 (N_10481,N_10101,N_10061);
nand U10482 (N_10482,N_9629,N_9767);
nor U10483 (N_10483,N_10113,N_9902);
nand U10484 (N_10484,N_10181,N_10194);
and U10485 (N_10485,N_9695,N_10124);
xor U10486 (N_10486,N_9835,N_9750);
or U10487 (N_10487,N_9813,N_9616);
xnor U10488 (N_10488,N_10180,N_9854);
and U10489 (N_10489,N_9865,N_9993);
xnor U10490 (N_10490,N_9985,N_9706);
xnor U10491 (N_10491,N_10091,N_9717);
nor U10492 (N_10492,N_9845,N_9759);
nand U10493 (N_10493,N_10145,N_10052);
nor U10494 (N_10494,N_9771,N_10078);
or U10495 (N_10495,N_9947,N_10097);
xnor U10496 (N_10496,N_10150,N_10039);
xnor U10497 (N_10497,N_9895,N_9936);
xnor U10498 (N_10498,N_9789,N_9930);
or U10499 (N_10499,N_10032,N_9762);
nand U10500 (N_10500,N_9979,N_9882);
and U10501 (N_10501,N_9686,N_9697);
xor U10502 (N_10502,N_9918,N_10033);
and U10503 (N_10503,N_9623,N_9642);
nand U10504 (N_10504,N_10161,N_9755);
or U10505 (N_10505,N_9685,N_9766);
nand U10506 (N_10506,N_10145,N_10120);
or U10507 (N_10507,N_9719,N_10190);
nand U10508 (N_10508,N_9957,N_9689);
nor U10509 (N_10509,N_9844,N_9767);
nand U10510 (N_10510,N_9625,N_9641);
xnor U10511 (N_10511,N_10095,N_9650);
and U10512 (N_10512,N_10052,N_10034);
xor U10513 (N_10513,N_9878,N_9827);
nand U10514 (N_10514,N_9777,N_10021);
nand U10515 (N_10515,N_10113,N_9925);
and U10516 (N_10516,N_10036,N_9869);
and U10517 (N_10517,N_10092,N_9623);
or U10518 (N_10518,N_9661,N_10036);
xor U10519 (N_10519,N_9942,N_9717);
and U10520 (N_10520,N_9840,N_9828);
or U10521 (N_10521,N_9751,N_9790);
or U10522 (N_10522,N_9915,N_9823);
xor U10523 (N_10523,N_9884,N_9687);
and U10524 (N_10524,N_9601,N_9859);
or U10525 (N_10525,N_10099,N_9785);
xor U10526 (N_10526,N_9847,N_9948);
nand U10527 (N_10527,N_10022,N_9801);
xnor U10528 (N_10528,N_9984,N_9865);
and U10529 (N_10529,N_9856,N_9809);
xnor U10530 (N_10530,N_9695,N_9871);
and U10531 (N_10531,N_9629,N_9910);
nor U10532 (N_10532,N_9948,N_9754);
and U10533 (N_10533,N_9741,N_10014);
xnor U10534 (N_10534,N_10168,N_9930);
xor U10535 (N_10535,N_9689,N_10061);
nor U10536 (N_10536,N_10021,N_9716);
nor U10537 (N_10537,N_9729,N_9743);
nand U10538 (N_10538,N_9635,N_9746);
and U10539 (N_10539,N_9765,N_10113);
and U10540 (N_10540,N_10001,N_9909);
or U10541 (N_10541,N_9693,N_9646);
or U10542 (N_10542,N_9861,N_9730);
nor U10543 (N_10543,N_9613,N_10092);
and U10544 (N_10544,N_9605,N_9872);
nand U10545 (N_10545,N_10052,N_9709);
nand U10546 (N_10546,N_9880,N_9925);
and U10547 (N_10547,N_9676,N_9886);
or U10548 (N_10548,N_9912,N_9874);
nor U10549 (N_10549,N_10152,N_9939);
nand U10550 (N_10550,N_9669,N_9926);
nor U10551 (N_10551,N_9641,N_10056);
and U10552 (N_10552,N_10064,N_10176);
and U10553 (N_10553,N_10087,N_9744);
nor U10554 (N_10554,N_9933,N_9800);
or U10555 (N_10555,N_10078,N_9643);
xor U10556 (N_10556,N_10154,N_9817);
nand U10557 (N_10557,N_9865,N_9670);
nand U10558 (N_10558,N_9628,N_10162);
nor U10559 (N_10559,N_9722,N_9743);
nor U10560 (N_10560,N_9762,N_10017);
and U10561 (N_10561,N_10111,N_9860);
nand U10562 (N_10562,N_9822,N_9973);
and U10563 (N_10563,N_9945,N_9609);
nor U10564 (N_10564,N_9894,N_9827);
nor U10565 (N_10565,N_10182,N_9909);
nor U10566 (N_10566,N_9621,N_9644);
and U10567 (N_10567,N_9769,N_9917);
nor U10568 (N_10568,N_10064,N_10035);
nor U10569 (N_10569,N_9667,N_9844);
xnor U10570 (N_10570,N_10032,N_9856);
xor U10571 (N_10571,N_9897,N_9814);
xnor U10572 (N_10572,N_9656,N_9820);
nor U10573 (N_10573,N_9747,N_9602);
or U10574 (N_10574,N_9985,N_9714);
nand U10575 (N_10575,N_9821,N_9997);
nor U10576 (N_10576,N_9677,N_9880);
nor U10577 (N_10577,N_9930,N_9795);
or U10578 (N_10578,N_9714,N_10056);
or U10579 (N_10579,N_9860,N_9686);
xnor U10580 (N_10580,N_9901,N_9772);
xnor U10581 (N_10581,N_9884,N_9608);
nor U10582 (N_10582,N_9860,N_10137);
nand U10583 (N_10583,N_9687,N_9608);
nor U10584 (N_10584,N_9766,N_10011);
and U10585 (N_10585,N_9959,N_10032);
and U10586 (N_10586,N_9767,N_9794);
and U10587 (N_10587,N_10040,N_9825);
and U10588 (N_10588,N_9614,N_10080);
and U10589 (N_10589,N_9834,N_9949);
or U10590 (N_10590,N_9919,N_9877);
xnor U10591 (N_10591,N_9882,N_9711);
nand U10592 (N_10592,N_9825,N_9728);
nand U10593 (N_10593,N_9716,N_10196);
xor U10594 (N_10594,N_9958,N_10046);
nand U10595 (N_10595,N_9725,N_9978);
xnor U10596 (N_10596,N_10080,N_9847);
and U10597 (N_10597,N_9867,N_9847);
nor U10598 (N_10598,N_9897,N_10033);
nor U10599 (N_10599,N_10131,N_9730);
xor U10600 (N_10600,N_9943,N_10041);
or U10601 (N_10601,N_9628,N_9712);
and U10602 (N_10602,N_10074,N_9701);
and U10603 (N_10603,N_10080,N_9874);
and U10604 (N_10604,N_9753,N_10143);
and U10605 (N_10605,N_9610,N_9746);
or U10606 (N_10606,N_10109,N_9657);
and U10607 (N_10607,N_9712,N_9757);
and U10608 (N_10608,N_10119,N_9798);
nand U10609 (N_10609,N_9664,N_9651);
nand U10610 (N_10610,N_9717,N_9883);
nand U10611 (N_10611,N_9987,N_10118);
nand U10612 (N_10612,N_10019,N_9603);
nor U10613 (N_10613,N_9683,N_9928);
nor U10614 (N_10614,N_9962,N_9694);
xnor U10615 (N_10615,N_9913,N_9916);
xnor U10616 (N_10616,N_9868,N_9753);
or U10617 (N_10617,N_10176,N_9620);
xnor U10618 (N_10618,N_9692,N_10055);
or U10619 (N_10619,N_10039,N_9960);
and U10620 (N_10620,N_10051,N_9748);
xor U10621 (N_10621,N_9667,N_10197);
nor U10622 (N_10622,N_9874,N_9823);
and U10623 (N_10623,N_9857,N_9936);
or U10624 (N_10624,N_9989,N_9951);
xnor U10625 (N_10625,N_10064,N_9990);
or U10626 (N_10626,N_10165,N_9946);
nor U10627 (N_10627,N_9780,N_10159);
xnor U10628 (N_10628,N_10131,N_9714);
xor U10629 (N_10629,N_9917,N_10049);
and U10630 (N_10630,N_10043,N_9809);
nor U10631 (N_10631,N_10183,N_10085);
and U10632 (N_10632,N_9689,N_10062);
xnor U10633 (N_10633,N_9641,N_9994);
nor U10634 (N_10634,N_9774,N_9994);
nor U10635 (N_10635,N_9996,N_9874);
nand U10636 (N_10636,N_10085,N_9631);
nor U10637 (N_10637,N_10144,N_9903);
and U10638 (N_10638,N_9904,N_10035);
or U10639 (N_10639,N_10171,N_10054);
and U10640 (N_10640,N_9635,N_9741);
and U10641 (N_10641,N_10081,N_9695);
xnor U10642 (N_10642,N_9700,N_9973);
nor U10643 (N_10643,N_10154,N_9819);
xnor U10644 (N_10644,N_9879,N_9964);
nand U10645 (N_10645,N_10170,N_9822);
nor U10646 (N_10646,N_9799,N_9962);
nor U10647 (N_10647,N_9723,N_9863);
or U10648 (N_10648,N_10142,N_9855);
nand U10649 (N_10649,N_9814,N_9981);
and U10650 (N_10650,N_9931,N_9829);
and U10651 (N_10651,N_9913,N_9847);
nor U10652 (N_10652,N_9984,N_9644);
nor U10653 (N_10653,N_9978,N_9830);
xnor U10654 (N_10654,N_9640,N_9701);
or U10655 (N_10655,N_9823,N_9816);
nor U10656 (N_10656,N_9789,N_10147);
or U10657 (N_10657,N_9657,N_9717);
nand U10658 (N_10658,N_9709,N_9633);
and U10659 (N_10659,N_9628,N_9766);
nor U10660 (N_10660,N_9996,N_9746);
or U10661 (N_10661,N_9875,N_9626);
xor U10662 (N_10662,N_9849,N_9862);
xnor U10663 (N_10663,N_9970,N_10002);
nor U10664 (N_10664,N_9756,N_9799);
nand U10665 (N_10665,N_9922,N_10035);
nand U10666 (N_10666,N_10002,N_10114);
nor U10667 (N_10667,N_10180,N_9907);
nand U10668 (N_10668,N_9927,N_9713);
nand U10669 (N_10669,N_10199,N_10189);
nor U10670 (N_10670,N_9865,N_9960);
nand U10671 (N_10671,N_9882,N_10127);
or U10672 (N_10672,N_9708,N_9804);
and U10673 (N_10673,N_9944,N_9720);
and U10674 (N_10674,N_10036,N_9946);
nor U10675 (N_10675,N_9808,N_9844);
nand U10676 (N_10676,N_9676,N_9644);
or U10677 (N_10677,N_9989,N_9973);
nand U10678 (N_10678,N_10140,N_9911);
xor U10679 (N_10679,N_10072,N_10009);
xor U10680 (N_10680,N_9646,N_9965);
nor U10681 (N_10681,N_10124,N_9896);
nand U10682 (N_10682,N_9871,N_9917);
and U10683 (N_10683,N_9734,N_10170);
nand U10684 (N_10684,N_9734,N_9617);
nor U10685 (N_10685,N_9839,N_10139);
or U10686 (N_10686,N_9694,N_10087);
and U10687 (N_10687,N_9853,N_9843);
or U10688 (N_10688,N_9663,N_10006);
nor U10689 (N_10689,N_9966,N_10074);
and U10690 (N_10690,N_9687,N_9753);
nand U10691 (N_10691,N_10072,N_9709);
and U10692 (N_10692,N_9743,N_9755);
xnor U10693 (N_10693,N_9848,N_9994);
or U10694 (N_10694,N_10119,N_9628);
and U10695 (N_10695,N_9614,N_10037);
nand U10696 (N_10696,N_9767,N_9713);
nand U10697 (N_10697,N_10125,N_9996);
nand U10698 (N_10698,N_9849,N_9763);
nor U10699 (N_10699,N_9750,N_9864);
and U10700 (N_10700,N_10197,N_10178);
xnor U10701 (N_10701,N_9868,N_9827);
nor U10702 (N_10702,N_9963,N_9889);
nand U10703 (N_10703,N_10091,N_10161);
nor U10704 (N_10704,N_9854,N_10023);
nand U10705 (N_10705,N_9974,N_9988);
and U10706 (N_10706,N_9736,N_9797);
xor U10707 (N_10707,N_9746,N_9919);
xor U10708 (N_10708,N_9977,N_9741);
xnor U10709 (N_10709,N_10067,N_9987);
xor U10710 (N_10710,N_9976,N_9809);
nand U10711 (N_10711,N_9785,N_10145);
and U10712 (N_10712,N_9962,N_9727);
xnor U10713 (N_10713,N_10173,N_10055);
nand U10714 (N_10714,N_9676,N_9652);
and U10715 (N_10715,N_9648,N_9991);
nor U10716 (N_10716,N_10143,N_9915);
or U10717 (N_10717,N_9742,N_9859);
and U10718 (N_10718,N_9670,N_9951);
or U10719 (N_10719,N_10080,N_9961);
xor U10720 (N_10720,N_10162,N_9929);
nor U10721 (N_10721,N_9711,N_9743);
or U10722 (N_10722,N_9972,N_9636);
xor U10723 (N_10723,N_10093,N_10126);
or U10724 (N_10724,N_9654,N_9891);
nor U10725 (N_10725,N_9867,N_10096);
and U10726 (N_10726,N_9708,N_10015);
nand U10727 (N_10727,N_10150,N_9770);
and U10728 (N_10728,N_10020,N_9769);
nor U10729 (N_10729,N_9782,N_10133);
nand U10730 (N_10730,N_10138,N_9837);
or U10731 (N_10731,N_9842,N_9856);
nand U10732 (N_10732,N_9861,N_9943);
and U10733 (N_10733,N_9626,N_9671);
or U10734 (N_10734,N_10010,N_9680);
nor U10735 (N_10735,N_9856,N_9649);
and U10736 (N_10736,N_10006,N_9706);
nor U10737 (N_10737,N_10030,N_9655);
or U10738 (N_10738,N_9627,N_10144);
nand U10739 (N_10739,N_9917,N_9733);
nand U10740 (N_10740,N_9982,N_10079);
nand U10741 (N_10741,N_10182,N_10006);
nand U10742 (N_10742,N_9848,N_10094);
and U10743 (N_10743,N_9919,N_9663);
nand U10744 (N_10744,N_9824,N_10006);
nand U10745 (N_10745,N_9981,N_9989);
nand U10746 (N_10746,N_9641,N_10174);
nor U10747 (N_10747,N_9797,N_9934);
nor U10748 (N_10748,N_9696,N_10185);
and U10749 (N_10749,N_9647,N_9978);
and U10750 (N_10750,N_9717,N_9993);
nor U10751 (N_10751,N_9774,N_9757);
or U10752 (N_10752,N_9727,N_9641);
and U10753 (N_10753,N_9845,N_10150);
or U10754 (N_10754,N_9664,N_10082);
nor U10755 (N_10755,N_10123,N_9673);
and U10756 (N_10756,N_9939,N_9933);
and U10757 (N_10757,N_9745,N_9985);
xor U10758 (N_10758,N_9992,N_9853);
or U10759 (N_10759,N_9630,N_9663);
or U10760 (N_10760,N_9767,N_9663);
or U10761 (N_10761,N_9864,N_9645);
nand U10762 (N_10762,N_9867,N_9623);
or U10763 (N_10763,N_9753,N_9817);
or U10764 (N_10764,N_9918,N_9924);
xor U10765 (N_10765,N_9992,N_9892);
xor U10766 (N_10766,N_9738,N_9764);
nand U10767 (N_10767,N_9895,N_9702);
nor U10768 (N_10768,N_9967,N_10156);
and U10769 (N_10769,N_10139,N_9893);
and U10770 (N_10770,N_9831,N_9908);
or U10771 (N_10771,N_9609,N_9643);
xor U10772 (N_10772,N_9631,N_9893);
xor U10773 (N_10773,N_10179,N_9707);
nand U10774 (N_10774,N_9864,N_9857);
and U10775 (N_10775,N_9866,N_10108);
and U10776 (N_10776,N_10186,N_10019);
xnor U10777 (N_10777,N_9951,N_10097);
or U10778 (N_10778,N_9709,N_9705);
xnor U10779 (N_10779,N_9679,N_9819);
xnor U10780 (N_10780,N_9627,N_9819);
and U10781 (N_10781,N_9803,N_10198);
xnor U10782 (N_10782,N_9671,N_9927);
or U10783 (N_10783,N_10185,N_9884);
nor U10784 (N_10784,N_9716,N_9751);
xnor U10785 (N_10785,N_9649,N_9842);
nand U10786 (N_10786,N_9835,N_9847);
nand U10787 (N_10787,N_9911,N_9888);
nand U10788 (N_10788,N_9678,N_9934);
nor U10789 (N_10789,N_9806,N_10025);
nand U10790 (N_10790,N_9751,N_10063);
or U10791 (N_10791,N_10050,N_9625);
or U10792 (N_10792,N_10045,N_9769);
and U10793 (N_10793,N_9810,N_9876);
and U10794 (N_10794,N_9905,N_9614);
nor U10795 (N_10795,N_9770,N_9964);
xnor U10796 (N_10796,N_9745,N_10164);
nand U10797 (N_10797,N_9662,N_10133);
nor U10798 (N_10798,N_9855,N_9725);
nand U10799 (N_10799,N_9801,N_9912);
nor U10800 (N_10800,N_10674,N_10229);
nand U10801 (N_10801,N_10424,N_10636);
and U10802 (N_10802,N_10604,N_10351);
and U10803 (N_10803,N_10336,N_10312);
nand U10804 (N_10804,N_10301,N_10614);
nand U10805 (N_10805,N_10585,N_10234);
and U10806 (N_10806,N_10331,N_10399);
and U10807 (N_10807,N_10349,N_10577);
nand U10808 (N_10808,N_10204,N_10439);
xor U10809 (N_10809,N_10630,N_10392);
xor U10810 (N_10810,N_10406,N_10690);
and U10811 (N_10811,N_10703,N_10322);
nor U10812 (N_10812,N_10563,N_10381);
or U10813 (N_10813,N_10654,N_10669);
nor U10814 (N_10814,N_10490,N_10318);
nand U10815 (N_10815,N_10309,N_10771);
nor U10816 (N_10816,N_10347,N_10208);
or U10817 (N_10817,N_10428,N_10691);
or U10818 (N_10818,N_10230,N_10698);
or U10819 (N_10819,N_10238,N_10214);
and U10820 (N_10820,N_10602,N_10376);
and U10821 (N_10821,N_10702,N_10274);
or U10822 (N_10822,N_10427,N_10773);
or U10823 (N_10823,N_10549,N_10500);
and U10824 (N_10824,N_10725,N_10753);
xnor U10825 (N_10825,N_10611,N_10780);
xnor U10826 (N_10826,N_10641,N_10571);
nand U10827 (N_10827,N_10603,N_10592);
xor U10828 (N_10828,N_10705,N_10419);
or U10829 (N_10829,N_10250,N_10546);
xor U10830 (N_10830,N_10390,N_10438);
nand U10831 (N_10831,N_10482,N_10334);
and U10832 (N_10832,N_10432,N_10648);
or U10833 (N_10833,N_10774,N_10403);
xnor U10834 (N_10834,N_10662,N_10615);
and U10835 (N_10835,N_10413,N_10610);
nor U10836 (N_10836,N_10668,N_10499);
nand U10837 (N_10837,N_10562,N_10223);
and U10838 (N_10838,N_10665,N_10260);
nor U10839 (N_10839,N_10405,N_10433);
nor U10840 (N_10840,N_10617,N_10586);
and U10841 (N_10841,N_10782,N_10242);
xnor U10842 (N_10842,N_10781,N_10741);
or U10843 (N_10843,N_10512,N_10310);
nor U10844 (N_10844,N_10776,N_10326);
nor U10845 (N_10845,N_10538,N_10294);
and U10846 (N_10846,N_10593,N_10319);
xor U10847 (N_10847,N_10777,N_10708);
nand U10848 (N_10848,N_10332,N_10409);
nor U10849 (N_10849,N_10706,N_10494);
nor U10850 (N_10850,N_10479,N_10335);
or U10851 (N_10851,N_10219,N_10755);
nand U10852 (N_10852,N_10385,N_10793);
xor U10853 (N_10853,N_10685,N_10532);
nand U10854 (N_10854,N_10232,N_10244);
or U10855 (N_10855,N_10442,N_10431);
nand U10856 (N_10856,N_10564,N_10302);
nand U10857 (N_10857,N_10278,N_10465);
xnor U10858 (N_10858,N_10368,N_10270);
nor U10859 (N_10859,N_10537,N_10251);
or U10860 (N_10860,N_10487,N_10201);
and U10861 (N_10861,N_10306,N_10621);
nor U10862 (N_10862,N_10695,N_10797);
nor U10863 (N_10863,N_10280,N_10700);
nand U10864 (N_10864,N_10366,N_10638);
xnor U10865 (N_10865,N_10361,N_10449);
and U10866 (N_10866,N_10380,N_10600);
or U10867 (N_10867,N_10440,N_10647);
nor U10868 (N_10868,N_10475,N_10474);
and U10869 (N_10869,N_10383,N_10358);
nor U10870 (N_10870,N_10519,N_10325);
or U10871 (N_10871,N_10649,N_10285);
and U10872 (N_10872,N_10227,N_10724);
or U10873 (N_10873,N_10580,N_10572);
or U10874 (N_10874,N_10411,N_10425);
or U10875 (N_10875,N_10561,N_10575);
or U10876 (N_10876,N_10501,N_10412);
and U10877 (N_10877,N_10275,N_10209);
or U10878 (N_10878,N_10417,N_10407);
xnor U10879 (N_10879,N_10779,N_10359);
nor U10880 (N_10880,N_10692,N_10434);
nand U10881 (N_10881,N_10517,N_10357);
or U10882 (N_10882,N_10697,N_10770);
xor U10883 (N_10883,N_10548,N_10203);
and U10884 (N_10884,N_10582,N_10544);
nor U10885 (N_10885,N_10416,N_10245);
or U10886 (N_10886,N_10282,N_10554);
nor U10887 (N_10887,N_10748,N_10418);
nand U10888 (N_10888,N_10423,N_10622);
xor U10889 (N_10889,N_10645,N_10590);
xor U10890 (N_10890,N_10353,N_10402);
or U10891 (N_10891,N_10284,N_10505);
and U10892 (N_10892,N_10369,N_10657);
nor U10893 (N_10893,N_10217,N_10296);
nor U10894 (N_10894,N_10791,N_10675);
xnor U10895 (N_10895,N_10429,N_10218);
xor U10896 (N_10896,N_10459,N_10528);
or U10897 (N_10897,N_10364,N_10252);
or U10898 (N_10898,N_10283,N_10723);
nor U10899 (N_10899,N_10660,N_10502);
nand U10900 (N_10900,N_10785,N_10467);
xor U10901 (N_10901,N_10206,N_10664);
xnor U10902 (N_10902,N_10255,N_10268);
nand U10903 (N_10903,N_10768,N_10569);
or U10904 (N_10904,N_10624,N_10410);
or U10905 (N_10905,N_10315,N_10720);
or U10906 (N_10906,N_10279,N_10488);
nor U10907 (N_10907,N_10277,N_10536);
nand U10908 (N_10908,N_10518,N_10680);
nand U10909 (N_10909,N_10395,N_10643);
or U10910 (N_10910,N_10452,N_10495);
and U10911 (N_10911,N_10430,N_10540);
nand U10912 (N_10912,N_10609,N_10455);
nor U10913 (N_10913,N_10738,N_10655);
or U10914 (N_10914,N_10701,N_10749);
nand U10915 (N_10915,N_10507,N_10769);
nand U10916 (N_10916,N_10631,N_10300);
and U10917 (N_10917,N_10530,N_10524);
or U10918 (N_10918,N_10513,N_10795);
xnor U10919 (N_10919,N_10717,N_10496);
xnor U10920 (N_10920,N_10265,N_10595);
nand U10921 (N_10921,N_10462,N_10486);
or U10922 (N_10922,N_10707,N_10320);
and U10923 (N_10923,N_10772,N_10667);
and U10924 (N_10924,N_10420,N_10736);
xor U10925 (N_10925,N_10313,N_10286);
or U10926 (N_10926,N_10216,N_10225);
or U10927 (N_10927,N_10751,N_10639);
nand U10928 (N_10928,N_10343,N_10401);
nor U10929 (N_10929,N_10323,N_10775);
xor U10930 (N_10930,N_10450,N_10453);
nor U10931 (N_10931,N_10759,N_10307);
or U10932 (N_10932,N_10345,N_10354);
or U10933 (N_10933,N_10632,N_10527);
xnor U10934 (N_10934,N_10523,N_10210);
or U10935 (N_10935,N_10644,N_10635);
nor U10936 (N_10936,N_10626,N_10333);
nand U10937 (N_10937,N_10295,N_10314);
xnor U10938 (N_10938,N_10202,N_10766);
and U10939 (N_10939,N_10257,N_10739);
or U10940 (N_10940,N_10704,N_10559);
nor U10941 (N_10941,N_10716,N_10346);
and U10942 (N_10942,N_10422,N_10509);
xnor U10943 (N_10943,N_10786,N_10447);
nor U10944 (N_10944,N_10292,N_10408);
and U10945 (N_10945,N_10484,N_10634);
and U10946 (N_10946,N_10340,N_10398);
nor U10947 (N_10947,N_10344,N_10226);
or U10948 (N_10948,N_10689,N_10756);
and U10949 (N_10949,N_10616,N_10220);
xnor U10950 (N_10950,N_10460,N_10762);
nor U10951 (N_10951,N_10221,N_10784);
nor U10952 (N_10952,N_10355,N_10480);
nor U10953 (N_10953,N_10783,N_10625);
and U10954 (N_10954,N_10367,N_10683);
and U10955 (N_10955,N_10397,N_10646);
or U10956 (N_10956,N_10686,N_10393);
xor U10957 (N_10957,N_10448,N_10678);
xor U10958 (N_10958,N_10497,N_10763);
nor U10959 (N_10959,N_10729,N_10477);
xnor U10960 (N_10960,N_10466,N_10799);
nand U10961 (N_10961,N_10248,N_10446);
xnor U10962 (N_10962,N_10663,N_10525);
and U10963 (N_10963,N_10271,N_10652);
and U10964 (N_10964,N_10761,N_10363);
nand U10965 (N_10965,N_10568,N_10712);
or U10966 (N_10966,N_10566,N_10608);
xor U10967 (N_10967,N_10718,N_10299);
and U10968 (N_10968,N_10200,N_10461);
and U10969 (N_10969,N_10579,N_10677);
nand U10970 (N_10970,N_10338,N_10317);
or U10971 (N_10971,N_10740,N_10514);
nand U10972 (N_10972,N_10574,N_10583);
or U10973 (N_10973,N_10289,N_10327);
xor U10974 (N_10974,N_10629,N_10670);
nor U10975 (N_10975,N_10236,N_10732);
or U10976 (N_10976,N_10263,N_10515);
nor U10977 (N_10977,N_10730,N_10735);
or U10978 (N_10978,N_10231,N_10253);
nand U10979 (N_10979,N_10481,N_10650);
and U10980 (N_10980,N_10444,N_10478);
nor U10981 (N_10981,N_10587,N_10553);
or U10982 (N_10982,N_10305,N_10699);
and U10983 (N_10983,N_10371,N_10387);
nand U10984 (N_10984,N_10261,N_10721);
xnor U10985 (N_10985,N_10436,N_10688);
and U10986 (N_10986,N_10653,N_10356);
nor U10987 (N_10987,N_10339,N_10471);
xor U10988 (N_10988,N_10522,N_10605);
and U10989 (N_10989,N_10764,N_10237);
nand U10990 (N_10990,N_10443,N_10370);
xor U10991 (N_10991,N_10687,N_10570);
or U10992 (N_10992,N_10394,N_10329);
or U10993 (N_10993,N_10728,N_10567);
and U10994 (N_10994,N_10599,N_10656);
nor U10995 (N_10995,N_10281,N_10754);
nor U10996 (N_10996,N_10640,N_10789);
and U10997 (N_10997,N_10388,N_10521);
xnor U10998 (N_10998,N_10758,N_10722);
xnor U10999 (N_10999,N_10249,N_10352);
or U11000 (N_11000,N_10287,N_10273);
nor U11001 (N_11001,N_10426,N_10489);
and U11002 (N_11002,N_10374,N_10328);
xor U11003 (N_11003,N_10246,N_10205);
xor U11004 (N_11004,N_10606,N_10619);
and U11005 (N_11005,N_10276,N_10247);
or U11006 (N_11006,N_10743,N_10298);
and U11007 (N_11007,N_10472,N_10671);
and U11008 (N_11008,N_10457,N_10711);
xor U11009 (N_11009,N_10547,N_10742);
xor U11010 (N_11010,N_10552,N_10324);
nand U11011 (N_11011,N_10551,N_10458);
or U11012 (N_11012,N_10601,N_10607);
or U11013 (N_11013,N_10360,N_10672);
xor U11014 (N_11014,N_10321,N_10588);
or U11015 (N_11015,N_10222,N_10212);
or U11016 (N_11016,N_10215,N_10498);
nand U11017 (N_11017,N_10391,N_10384);
or U11018 (N_11018,N_10684,N_10414);
nand U11019 (N_11019,N_10239,N_10794);
or U11020 (N_11020,N_10241,N_10233);
nor U11021 (N_11021,N_10679,N_10709);
xor U11022 (N_11022,N_10262,N_10661);
nor U11023 (N_11023,N_10737,N_10375);
or U11024 (N_11024,N_10485,N_10578);
xnor U11025 (N_11025,N_10362,N_10539);
and U11026 (N_11026,N_10682,N_10435);
nand U11027 (N_11027,N_10290,N_10581);
and U11028 (N_11028,N_10437,N_10267);
nand U11029 (N_11029,N_10589,N_10594);
nor U11030 (N_11030,N_10787,N_10348);
nor U11031 (N_11031,N_10788,N_10681);
nand U11032 (N_11032,N_10464,N_10765);
nor U11033 (N_11033,N_10243,N_10731);
nor U11034 (N_11034,N_10757,N_10710);
xor U11035 (N_11035,N_10303,N_10213);
xor U11036 (N_11036,N_10400,N_10269);
and U11037 (N_11037,N_10372,N_10228);
or U11038 (N_11038,N_10713,N_10637);
or U11039 (N_11039,N_10342,N_10476);
xnor U11040 (N_11040,N_10456,N_10311);
or U11041 (N_11041,N_10365,N_10560);
nor U11042 (N_11042,N_10613,N_10516);
and U11043 (N_11043,N_10378,N_10373);
or U11044 (N_11044,N_10760,N_10535);
nand U11045 (N_11045,N_10316,N_10386);
or U11046 (N_11046,N_10337,N_10767);
and U11047 (N_11047,N_10473,N_10506);
and U11048 (N_11048,N_10792,N_10543);
and U11049 (N_11049,N_10676,N_10441);
xnor U11050 (N_11050,N_10520,N_10240);
xor U11051 (N_11051,N_10483,N_10211);
and U11052 (N_11052,N_10673,N_10341);
and U11053 (N_11053,N_10529,N_10235);
nor U11054 (N_11054,N_10291,N_10573);
xor U11055 (N_11055,N_10207,N_10726);
and U11056 (N_11056,N_10531,N_10597);
nand U11057 (N_11057,N_10790,N_10747);
and U11058 (N_11058,N_10715,N_10224);
and U11059 (N_11059,N_10469,N_10350);
or U11060 (N_11060,N_10468,N_10598);
nor U11061 (N_11061,N_10454,N_10744);
or U11062 (N_11062,N_10382,N_10451);
or U11063 (N_11063,N_10693,N_10259);
or U11064 (N_11064,N_10445,N_10666);
and U11065 (N_11065,N_10557,N_10746);
nand U11066 (N_11066,N_10752,N_10493);
nand U11067 (N_11067,N_10623,N_10297);
xnor U11068 (N_11068,N_10526,N_10555);
xor U11069 (N_11069,N_10511,N_10542);
or U11070 (N_11070,N_10389,N_10658);
or U11071 (N_11071,N_10492,N_10258);
nand U11072 (N_11072,N_10659,N_10651);
nand U11073 (N_11073,N_10696,N_10508);
or U11074 (N_11074,N_10558,N_10541);
or U11075 (N_11075,N_10491,N_10596);
nand U11076 (N_11076,N_10304,N_10404);
xnor U11077 (N_11077,N_10620,N_10510);
or U11078 (N_11078,N_10503,N_10714);
or U11079 (N_11079,N_10627,N_10533);
or U11080 (N_11080,N_10470,N_10798);
nand U11081 (N_11081,N_10534,N_10550);
nor U11082 (N_11082,N_10633,N_10377);
nor U11083 (N_11083,N_10778,N_10330);
or U11084 (N_11084,N_10628,N_10565);
or U11085 (N_11085,N_10545,N_10254);
xor U11086 (N_11086,N_10308,N_10734);
nand U11087 (N_11087,N_10256,N_10421);
or U11088 (N_11088,N_10745,N_10796);
xnor U11089 (N_11089,N_10288,N_10719);
nor U11090 (N_11090,N_10556,N_10463);
xor U11091 (N_11091,N_10264,N_10694);
nor U11092 (N_11092,N_10396,N_10379);
nor U11093 (N_11093,N_10415,N_10272);
nor U11094 (N_11094,N_10727,N_10750);
and U11095 (N_11095,N_10642,N_10584);
nor U11096 (N_11096,N_10612,N_10266);
nand U11097 (N_11097,N_10504,N_10733);
nor U11098 (N_11098,N_10576,N_10591);
nor U11099 (N_11099,N_10293,N_10618);
and U11100 (N_11100,N_10425,N_10281);
xor U11101 (N_11101,N_10363,N_10258);
or U11102 (N_11102,N_10392,N_10471);
nand U11103 (N_11103,N_10695,N_10321);
nand U11104 (N_11104,N_10271,N_10626);
or U11105 (N_11105,N_10555,N_10411);
nor U11106 (N_11106,N_10765,N_10338);
and U11107 (N_11107,N_10709,N_10730);
or U11108 (N_11108,N_10292,N_10226);
nand U11109 (N_11109,N_10469,N_10407);
or U11110 (N_11110,N_10376,N_10499);
nand U11111 (N_11111,N_10308,N_10274);
and U11112 (N_11112,N_10408,N_10361);
and U11113 (N_11113,N_10461,N_10245);
and U11114 (N_11114,N_10571,N_10598);
nor U11115 (N_11115,N_10383,N_10487);
xnor U11116 (N_11116,N_10361,N_10247);
nor U11117 (N_11117,N_10249,N_10294);
nand U11118 (N_11118,N_10500,N_10444);
nor U11119 (N_11119,N_10221,N_10662);
xor U11120 (N_11120,N_10605,N_10665);
and U11121 (N_11121,N_10546,N_10600);
xnor U11122 (N_11122,N_10610,N_10793);
nand U11123 (N_11123,N_10662,N_10440);
and U11124 (N_11124,N_10656,N_10259);
and U11125 (N_11125,N_10344,N_10293);
or U11126 (N_11126,N_10312,N_10387);
or U11127 (N_11127,N_10388,N_10561);
nand U11128 (N_11128,N_10240,N_10628);
xnor U11129 (N_11129,N_10306,N_10469);
and U11130 (N_11130,N_10645,N_10693);
or U11131 (N_11131,N_10499,N_10341);
nor U11132 (N_11132,N_10508,N_10639);
nor U11133 (N_11133,N_10302,N_10608);
or U11134 (N_11134,N_10410,N_10451);
and U11135 (N_11135,N_10359,N_10722);
nor U11136 (N_11136,N_10337,N_10562);
nor U11137 (N_11137,N_10339,N_10489);
or U11138 (N_11138,N_10281,N_10578);
and U11139 (N_11139,N_10757,N_10287);
or U11140 (N_11140,N_10202,N_10643);
or U11141 (N_11141,N_10402,N_10252);
xnor U11142 (N_11142,N_10577,N_10709);
nor U11143 (N_11143,N_10746,N_10662);
xor U11144 (N_11144,N_10249,N_10322);
and U11145 (N_11145,N_10699,N_10609);
nor U11146 (N_11146,N_10628,N_10763);
nor U11147 (N_11147,N_10414,N_10762);
xnor U11148 (N_11148,N_10640,N_10393);
and U11149 (N_11149,N_10267,N_10441);
nand U11150 (N_11150,N_10265,N_10362);
nand U11151 (N_11151,N_10429,N_10686);
and U11152 (N_11152,N_10454,N_10771);
nand U11153 (N_11153,N_10558,N_10467);
and U11154 (N_11154,N_10728,N_10534);
nand U11155 (N_11155,N_10790,N_10709);
nand U11156 (N_11156,N_10294,N_10229);
nand U11157 (N_11157,N_10200,N_10335);
nor U11158 (N_11158,N_10517,N_10748);
xor U11159 (N_11159,N_10510,N_10286);
nand U11160 (N_11160,N_10577,N_10699);
or U11161 (N_11161,N_10270,N_10434);
nand U11162 (N_11162,N_10682,N_10717);
or U11163 (N_11163,N_10465,N_10785);
or U11164 (N_11164,N_10754,N_10721);
xnor U11165 (N_11165,N_10426,N_10245);
xnor U11166 (N_11166,N_10416,N_10660);
or U11167 (N_11167,N_10220,N_10642);
and U11168 (N_11168,N_10572,N_10203);
nor U11169 (N_11169,N_10256,N_10732);
or U11170 (N_11170,N_10243,N_10217);
nand U11171 (N_11171,N_10246,N_10754);
and U11172 (N_11172,N_10414,N_10264);
xor U11173 (N_11173,N_10218,N_10460);
and U11174 (N_11174,N_10720,N_10213);
or U11175 (N_11175,N_10230,N_10758);
nor U11176 (N_11176,N_10636,N_10752);
nand U11177 (N_11177,N_10508,N_10598);
nor U11178 (N_11178,N_10448,N_10337);
nor U11179 (N_11179,N_10250,N_10243);
and U11180 (N_11180,N_10582,N_10490);
nor U11181 (N_11181,N_10238,N_10642);
nor U11182 (N_11182,N_10357,N_10789);
and U11183 (N_11183,N_10665,N_10738);
nor U11184 (N_11184,N_10751,N_10416);
xor U11185 (N_11185,N_10576,N_10316);
or U11186 (N_11186,N_10526,N_10553);
nand U11187 (N_11187,N_10660,N_10539);
nand U11188 (N_11188,N_10652,N_10333);
and U11189 (N_11189,N_10736,N_10691);
or U11190 (N_11190,N_10585,N_10648);
nand U11191 (N_11191,N_10480,N_10564);
or U11192 (N_11192,N_10690,N_10241);
or U11193 (N_11193,N_10347,N_10784);
nand U11194 (N_11194,N_10550,N_10689);
nor U11195 (N_11195,N_10447,N_10226);
nand U11196 (N_11196,N_10370,N_10492);
or U11197 (N_11197,N_10666,N_10237);
nand U11198 (N_11198,N_10756,N_10566);
nand U11199 (N_11199,N_10679,N_10400);
xor U11200 (N_11200,N_10441,N_10594);
xnor U11201 (N_11201,N_10495,N_10227);
and U11202 (N_11202,N_10462,N_10524);
or U11203 (N_11203,N_10491,N_10492);
or U11204 (N_11204,N_10236,N_10753);
and U11205 (N_11205,N_10271,N_10587);
xnor U11206 (N_11206,N_10781,N_10277);
nand U11207 (N_11207,N_10423,N_10440);
nand U11208 (N_11208,N_10348,N_10521);
or U11209 (N_11209,N_10514,N_10257);
and U11210 (N_11210,N_10510,N_10454);
nor U11211 (N_11211,N_10309,N_10512);
nand U11212 (N_11212,N_10645,N_10650);
nor U11213 (N_11213,N_10676,N_10589);
nand U11214 (N_11214,N_10209,N_10744);
and U11215 (N_11215,N_10419,N_10788);
xor U11216 (N_11216,N_10621,N_10522);
nor U11217 (N_11217,N_10621,N_10355);
nor U11218 (N_11218,N_10240,N_10254);
nor U11219 (N_11219,N_10480,N_10747);
nor U11220 (N_11220,N_10488,N_10237);
or U11221 (N_11221,N_10734,N_10313);
xnor U11222 (N_11222,N_10428,N_10513);
nor U11223 (N_11223,N_10348,N_10319);
xor U11224 (N_11224,N_10384,N_10485);
nor U11225 (N_11225,N_10688,N_10773);
xnor U11226 (N_11226,N_10418,N_10769);
xor U11227 (N_11227,N_10550,N_10219);
xnor U11228 (N_11228,N_10782,N_10307);
and U11229 (N_11229,N_10276,N_10436);
nor U11230 (N_11230,N_10330,N_10793);
nor U11231 (N_11231,N_10320,N_10686);
nor U11232 (N_11232,N_10265,N_10428);
or U11233 (N_11233,N_10774,N_10413);
and U11234 (N_11234,N_10655,N_10639);
nor U11235 (N_11235,N_10396,N_10294);
xnor U11236 (N_11236,N_10527,N_10250);
and U11237 (N_11237,N_10796,N_10224);
nand U11238 (N_11238,N_10469,N_10771);
xor U11239 (N_11239,N_10368,N_10718);
xnor U11240 (N_11240,N_10288,N_10507);
and U11241 (N_11241,N_10425,N_10732);
and U11242 (N_11242,N_10379,N_10697);
nand U11243 (N_11243,N_10721,N_10585);
and U11244 (N_11244,N_10413,N_10209);
nand U11245 (N_11245,N_10619,N_10362);
nand U11246 (N_11246,N_10528,N_10557);
nor U11247 (N_11247,N_10652,N_10306);
nand U11248 (N_11248,N_10292,N_10484);
and U11249 (N_11249,N_10513,N_10450);
xnor U11250 (N_11250,N_10303,N_10670);
and U11251 (N_11251,N_10593,N_10391);
and U11252 (N_11252,N_10717,N_10396);
nand U11253 (N_11253,N_10626,N_10679);
nand U11254 (N_11254,N_10522,N_10537);
nor U11255 (N_11255,N_10668,N_10795);
and U11256 (N_11256,N_10788,N_10536);
xor U11257 (N_11257,N_10474,N_10372);
nor U11258 (N_11258,N_10651,N_10556);
xnor U11259 (N_11259,N_10504,N_10234);
nand U11260 (N_11260,N_10725,N_10390);
nor U11261 (N_11261,N_10765,N_10788);
or U11262 (N_11262,N_10463,N_10301);
nor U11263 (N_11263,N_10689,N_10671);
nand U11264 (N_11264,N_10618,N_10369);
nor U11265 (N_11265,N_10207,N_10520);
xor U11266 (N_11266,N_10666,N_10716);
and U11267 (N_11267,N_10642,N_10624);
nand U11268 (N_11268,N_10309,N_10701);
nand U11269 (N_11269,N_10679,N_10515);
nand U11270 (N_11270,N_10622,N_10511);
nand U11271 (N_11271,N_10461,N_10787);
and U11272 (N_11272,N_10420,N_10761);
nand U11273 (N_11273,N_10590,N_10272);
xor U11274 (N_11274,N_10284,N_10625);
or U11275 (N_11275,N_10608,N_10481);
nand U11276 (N_11276,N_10737,N_10229);
xnor U11277 (N_11277,N_10265,N_10677);
xnor U11278 (N_11278,N_10241,N_10649);
xor U11279 (N_11279,N_10687,N_10574);
xor U11280 (N_11280,N_10706,N_10230);
and U11281 (N_11281,N_10597,N_10624);
or U11282 (N_11282,N_10659,N_10691);
nand U11283 (N_11283,N_10485,N_10730);
nand U11284 (N_11284,N_10687,N_10598);
nor U11285 (N_11285,N_10441,N_10544);
or U11286 (N_11286,N_10665,N_10488);
or U11287 (N_11287,N_10680,N_10797);
xor U11288 (N_11288,N_10393,N_10402);
nor U11289 (N_11289,N_10477,N_10603);
xor U11290 (N_11290,N_10322,N_10401);
or U11291 (N_11291,N_10478,N_10487);
nand U11292 (N_11292,N_10562,N_10373);
or U11293 (N_11293,N_10645,N_10746);
xor U11294 (N_11294,N_10362,N_10239);
nor U11295 (N_11295,N_10630,N_10687);
and U11296 (N_11296,N_10362,N_10368);
nor U11297 (N_11297,N_10733,N_10709);
or U11298 (N_11298,N_10771,N_10205);
xnor U11299 (N_11299,N_10728,N_10278);
nand U11300 (N_11300,N_10411,N_10484);
xnor U11301 (N_11301,N_10308,N_10298);
or U11302 (N_11302,N_10376,N_10269);
and U11303 (N_11303,N_10290,N_10316);
nand U11304 (N_11304,N_10570,N_10711);
xor U11305 (N_11305,N_10289,N_10434);
xor U11306 (N_11306,N_10730,N_10409);
nand U11307 (N_11307,N_10639,N_10225);
or U11308 (N_11308,N_10201,N_10503);
nand U11309 (N_11309,N_10630,N_10201);
xor U11310 (N_11310,N_10771,N_10556);
nand U11311 (N_11311,N_10497,N_10399);
or U11312 (N_11312,N_10734,N_10244);
nor U11313 (N_11313,N_10462,N_10771);
nor U11314 (N_11314,N_10326,N_10355);
nand U11315 (N_11315,N_10325,N_10639);
or U11316 (N_11316,N_10301,N_10724);
and U11317 (N_11317,N_10470,N_10301);
xnor U11318 (N_11318,N_10751,N_10449);
nor U11319 (N_11319,N_10722,N_10463);
nand U11320 (N_11320,N_10653,N_10526);
nor U11321 (N_11321,N_10485,N_10256);
nand U11322 (N_11322,N_10502,N_10370);
xor U11323 (N_11323,N_10637,N_10722);
xnor U11324 (N_11324,N_10749,N_10527);
and U11325 (N_11325,N_10699,N_10649);
nor U11326 (N_11326,N_10306,N_10232);
and U11327 (N_11327,N_10484,N_10579);
nor U11328 (N_11328,N_10333,N_10207);
and U11329 (N_11329,N_10316,N_10602);
nand U11330 (N_11330,N_10279,N_10227);
and U11331 (N_11331,N_10405,N_10496);
and U11332 (N_11332,N_10214,N_10267);
and U11333 (N_11333,N_10454,N_10417);
xnor U11334 (N_11334,N_10384,N_10366);
nand U11335 (N_11335,N_10701,N_10397);
and U11336 (N_11336,N_10482,N_10218);
and U11337 (N_11337,N_10430,N_10573);
nand U11338 (N_11338,N_10459,N_10476);
and U11339 (N_11339,N_10254,N_10484);
nand U11340 (N_11340,N_10612,N_10446);
nand U11341 (N_11341,N_10643,N_10663);
nor U11342 (N_11342,N_10664,N_10344);
nor U11343 (N_11343,N_10726,N_10277);
nor U11344 (N_11344,N_10262,N_10403);
and U11345 (N_11345,N_10502,N_10493);
nand U11346 (N_11346,N_10706,N_10235);
nand U11347 (N_11347,N_10281,N_10601);
nand U11348 (N_11348,N_10686,N_10617);
and U11349 (N_11349,N_10646,N_10656);
xnor U11350 (N_11350,N_10313,N_10407);
nand U11351 (N_11351,N_10350,N_10479);
or U11352 (N_11352,N_10541,N_10273);
or U11353 (N_11353,N_10485,N_10337);
and U11354 (N_11354,N_10751,N_10284);
xnor U11355 (N_11355,N_10497,N_10377);
or U11356 (N_11356,N_10480,N_10248);
nand U11357 (N_11357,N_10257,N_10799);
xor U11358 (N_11358,N_10345,N_10779);
nor U11359 (N_11359,N_10222,N_10463);
nor U11360 (N_11360,N_10698,N_10414);
nor U11361 (N_11361,N_10472,N_10741);
and U11362 (N_11362,N_10420,N_10539);
xnor U11363 (N_11363,N_10772,N_10704);
xor U11364 (N_11364,N_10405,N_10463);
and U11365 (N_11365,N_10431,N_10295);
nand U11366 (N_11366,N_10578,N_10796);
xor U11367 (N_11367,N_10368,N_10587);
xnor U11368 (N_11368,N_10282,N_10671);
xnor U11369 (N_11369,N_10637,N_10373);
or U11370 (N_11370,N_10401,N_10371);
xor U11371 (N_11371,N_10577,N_10754);
xor U11372 (N_11372,N_10775,N_10598);
xnor U11373 (N_11373,N_10490,N_10527);
nor U11374 (N_11374,N_10483,N_10393);
nor U11375 (N_11375,N_10259,N_10447);
nor U11376 (N_11376,N_10318,N_10767);
and U11377 (N_11377,N_10201,N_10710);
and U11378 (N_11378,N_10673,N_10242);
or U11379 (N_11379,N_10381,N_10218);
nand U11380 (N_11380,N_10729,N_10431);
or U11381 (N_11381,N_10515,N_10370);
or U11382 (N_11382,N_10421,N_10448);
or U11383 (N_11383,N_10267,N_10411);
nor U11384 (N_11384,N_10363,N_10721);
nand U11385 (N_11385,N_10703,N_10394);
nor U11386 (N_11386,N_10730,N_10411);
nand U11387 (N_11387,N_10443,N_10454);
xor U11388 (N_11388,N_10584,N_10649);
nor U11389 (N_11389,N_10321,N_10551);
nand U11390 (N_11390,N_10256,N_10778);
nor U11391 (N_11391,N_10712,N_10335);
and U11392 (N_11392,N_10476,N_10739);
nor U11393 (N_11393,N_10733,N_10783);
nand U11394 (N_11394,N_10360,N_10798);
nor U11395 (N_11395,N_10579,N_10589);
xor U11396 (N_11396,N_10750,N_10352);
nand U11397 (N_11397,N_10571,N_10283);
xor U11398 (N_11398,N_10495,N_10599);
xor U11399 (N_11399,N_10390,N_10217);
nand U11400 (N_11400,N_10830,N_10846);
xnor U11401 (N_11401,N_11368,N_10872);
nand U11402 (N_11402,N_11360,N_10861);
nand U11403 (N_11403,N_10842,N_11310);
or U11404 (N_11404,N_11388,N_11023);
or U11405 (N_11405,N_10913,N_11155);
and U11406 (N_11406,N_11312,N_10994);
and U11407 (N_11407,N_10865,N_11358);
nor U11408 (N_11408,N_11392,N_10945);
or U11409 (N_11409,N_11100,N_11379);
or U11410 (N_11410,N_10902,N_10895);
nor U11411 (N_11411,N_10996,N_11139);
xor U11412 (N_11412,N_11119,N_10826);
xor U11413 (N_11413,N_11134,N_11026);
nor U11414 (N_11414,N_10901,N_11185);
nor U11415 (N_11415,N_10951,N_11210);
nand U11416 (N_11416,N_10900,N_11265);
nand U11417 (N_11417,N_11326,N_11107);
nor U11418 (N_11418,N_11094,N_11218);
or U11419 (N_11419,N_11200,N_11315);
xnor U11420 (N_11420,N_11151,N_11266);
nand U11421 (N_11421,N_11005,N_10934);
xnor U11422 (N_11422,N_11015,N_10899);
nand U11423 (N_11423,N_11330,N_11150);
and U11424 (N_11424,N_11278,N_11209);
xor U11425 (N_11425,N_11165,N_11334);
xnor U11426 (N_11426,N_11186,N_11140);
xnor U11427 (N_11427,N_10952,N_11357);
xor U11428 (N_11428,N_10877,N_11125);
nand U11429 (N_11429,N_10985,N_11008);
nor U11430 (N_11430,N_11036,N_11286);
or U11431 (N_11431,N_11304,N_11093);
nand U11432 (N_11432,N_11257,N_11145);
nand U11433 (N_11433,N_11007,N_11154);
and U11434 (N_11434,N_11160,N_11287);
nor U11435 (N_11435,N_11375,N_11045);
or U11436 (N_11436,N_10839,N_11296);
xnor U11437 (N_11437,N_11307,N_10936);
nor U11438 (N_11438,N_10813,N_11173);
or U11439 (N_11439,N_11110,N_11213);
and U11440 (N_11440,N_10954,N_11269);
or U11441 (N_11441,N_11124,N_11108);
or U11442 (N_11442,N_11159,N_11277);
nand U11443 (N_11443,N_11120,N_11298);
nor U11444 (N_11444,N_11224,N_10818);
and U11445 (N_11445,N_11313,N_11196);
and U11446 (N_11446,N_11002,N_11361);
nand U11447 (N_11447,N_10930,N_11299);
nor U11448 (N_11448,N_11342,N_11053);
nor U11449 (N_11449,N_11086,N_11148);
nor U11450 (N_11450,N_10935,N_10843);
xor U11451 (N_11451,N_11212,N_11291);
xor U11452 (N_11452,N_10948,N_11144);
nand U11453 (N_11453,N_11081,N_11314);
nand U11454 (N_11454,N_11275,N_11395);
xor U11455 (N_11455,N_11131,N_11038);
xnor U11456 (N_11456,N_10822,N_10941);
nor U11457 (N_11457,N_10836,N_10938);
nor U11458 (N_11458,N_11063,N_11169);
xnor U11459 (N_11459,N_11013,N_11208);
and U11460 (N_11460,N_11092,N_10897);
xnor U11461 (N_11461,N_11306,N_10880);
xor U11462 (N_11462,N_11260,N_11198);
nor U11463 (N_11463,N_11029,N_10926);
or U11464 (N_11464,N_10851,N_11399);
nor U11465 (N_11465,N_10875,N_11164);
and U11466 (N_11466,N_11338,N_10881);
and U11467 (N_11467,N_11153,N_11389);
nor U11468 (N_11468,N_10959,N_11237);
xnor U11469 (N_11469,N_11295,N_10835);
xor U11470 (N_11470,N_11365,N_10983);
nor U11471 (N_11471,N_11281,N_10847);
and U11472 (N_11472,N_10873,N_11128);
xor U11473 (N_11473,N_11270,N_10982);
nand U11474 (N_11474,N_10924,N_11121);
and U11475 (N_11475,N_11006,N_10838);
and U11476 (N_11476,N_10907,N_11157);
or U11477 (N_11477,N_10988,N_10834);
and U11478 (N_11478,N_10810,N_11207);
nor U11479 (N_11479,N_11308,N_11137);
nand U11480 (N_11480,N_11058,N_10801);
nand U11481 (N_11481,N_11079,N_11027);
xor U11482 (N_11482,N_10968,N_10989);
and U11483 (N_11483,N_10979,N_11283);
nand U11484 (N_11484,N_11359,N_11259);
nand U11485 (N_11485,N_11227,N_11180);
and U11486 (N_11486,N_10944,N_10874);
xnor U11487 (N_11487,N_11397,N_11251);
nor U11488 (N_11488,N_11245,N_11043);
or U11489 (N_11489,N_11122,N_10870);
and U11490 (N_11490,N_10990,N_10860);
xor U11491 (N_11491,N_11235,N_11143);
nor U11492 (N_11492,N_10817,N_11345);
nor U11493 (N_11493,N_10933,N_11132);
and U11494 (N_11494,N_11332,N_11320);
xnor U11495 (N_11495,N_11255,N_11221);
and U11496 (N_11496,N_11367,N_11273);
and U11497 (N_11497,N_11206,N_11177);
xor U11498 (N_11498,N_11019,N_10960);
xor U11499 (N_11499,N_11030,N_11138);
xor U11500 (N_11500,N_10950,N_10845);
xor U11501 (N_11501,N_11352,N_10962);
nand U11502 (N_11502,N_11187,N_10921);
and U11503 (N_11503,N_10858,N_11032);
and U11504 (N_11504,N_10920,N_10925);
and U11505 (N_11505,N_10850,N_10819);
and U11506 (N_11506,N_11335,N_11271);
nand U11507 (N_11507,N_10854,N_10906);
nand U11508 (N_11508,N_11040,N_11072);
or U11509 (N_11509,N_11055,N_10882);
nand U11510 (N_11510,N_11396,N_11267);
or U11511 (N_11511,N_11398,N_11238);
nor U11512 (N_11512,N_11189,N_11303);
and U11513 (N_11513,N_11370,N_11195);
nor U11514 (N_11514,N_11044,N_11323);
nand U11515 (N_11515,N_10943,N_11056);
or U11516 (N_11516,N_11112,N_11118);
xor U11517 (N_11517,N_11067,N_11321);
or U11518 (N_11518,N_10997,N_11162);
nand U11519 (N_11519,N_11356,N_11022);
or U11520 (N_11520,N_11188,N_10947);
xnor U11521 (N_11521,N_11147,N_11347);
or U11522 (N_11522,N_11109,N_11101);
or U11523 (N_11523,N_11116,N_10905);
nand U11524 (N_11524,N_10909,N_11129);
and U11525 (N_11525,N_11016,N_11024);
nand U11526 (N_11526,N_11025,N_11219);
nor U11527 (N_11527,N_10912,N_11082);
or U11528 (N_11528,N_10859,N_10977);
xnor U11529 (N_11529,N_11127,N_11300);
or U11530 (N_11530,N_11102,N_10857);
nand U11531 (N_11531,N_10837,N_10987);
nor U11532 (N_11532,N_11037,N_11111);
nand U11533 (N_11533,N_10804,N_11062);
or U11534 (N_11534,N_11009,N_11241);
nand U11535 (N_11535,N_10896,N_10879);
nor U11536 (N_11536,N_11010,N_11204);
or U11537 (N_11537,N_11211,N_11123);
xor U11538 (N_11538,N_10863,N_10803);
nor U11539 (N_11539,N_10946,N_11105);
nor U11540 (N_11540,N_10972,N_10832);
nor U11541 (N_11541,N_11136,N_11194);
or U11542 (N_11542,N_11066,N_10829);
or U11543 (N_11543,N_11353,N_11325);
nand U11544 (N_11544,N_10973,N_10908);
xor U11545 (N_11545,N_10931,N_11231);
nand U11546 (N_11546,N_11004,N_10998);
or U11547 (N_11547,N_11234,N_11228);
nand U11548 (N_11548,N_11135,N_11167);
or U11549 (N_11549,N_11191,N_10961);
nor U11550 (N_11550,N_10999,N_11034);
and U11551 (N_11551,N_11190,N_10868);
nand U11552 (N_11552,N_11028,N_11099);
and U11553 (N_11553,N_11371,N_11233);
nor U11554 (N_11554,N_11252,N_11331);
and U11555 (N_11555,N_11214,N_11236);
and U11556 (N_11556,N_11372,N_11051);
nand U11557 (N_11557,N_11011,N_10911);
and U11558 (N_11558,N_11272,N_11052);
nor U11559 (N_11559,N_11288,N_11130);
nor U11560 (N_11560,N_11279,N_11316);
nand U11561 (N_11561,N_11250,N_11166);
and U11562 (N_11562,N_11184,N_10984);
nand U11563 (N_11563,N_11098,N_11373);
and U11564 (N_11564,N_11017,N_11362);
xnor U11565 (N_11565,N_10993,N_11341);
and U11566 (N_11566,N_11317,N_10958);
or U11567 (N_11567,N_10891,N_10883);
or U11568 (N_11568,N_10964,N_11083);
xor U11569 (N_11569,N_11355,N_11337);
or U11570 (N_11570,N_11378,N_10853);
and U11571 (N_11571,N_10808,N_11264);
nor U11572 (N_11572,N_11369,N_11163);
or U11573 (N_11573,N_11292,N_10806);
nor U11574 (N_11574,N_10923,N_10840);
nor U11575 (N_11575,N_11168,N_11174);
xnor U11576 (N_11576,N_11046,N_10919);
and U11577 (N_11577,N_10825,N_11088);
xor U11578 (N_11578,N_11350,N_11178);
nand U11579 (N_11579,N_11229,N_10816);
xnor U11580 (N_11580,N_10886,N_11071);
xor U11581 (N_11581,N_11202,N_11181);
xnor U11582 (N_11582,N_10820,N_10956);
nor U11583 (N_11583,N_11285,N_10831);
and U11584 (N_11584,N_10890,N_10855);
xnor U11585 (N_11585,N_11376,N_11087);
nor U11586 (N_11586,N_11170,N_11289);
xnor U11587 (N_11587,N_10889,N_10824);
and U11588 (N_11588,N_10927,N_10975);
xor U11589 (N_11589,N_10986,N_10957);
xnor U11590 (N_11590,N_10915,N_11047);
or U11591 (N_11591,N_10884,N_11329);
and U11592 (N_11592,N_11203,N_11319);
or U11593 (N_11593,N_11197,N_10992);
xnor U11594 (N_11594,N_11077,N_10841);
xor U11595 (N_11595,N_11089,N_11220);
nand U11596 (N_11596,N_11050,N_11156);
or U11597 (N_11597,N_10876,N_10869);
nand U11598 (N_11598,N_11363,N_11284);
or U11599 (N_11599,N_11183,N_11280);
or U11600 (N_11600,N_11254,N_10966);
and U11601 (N_11601,N_10910,N_11258);
nand U11602 (N_11602,N_11274,N_11247);
xor U11603 (N_11603,N_11018,N_10981);
or U11604 (N_11604,N_10805,N_10821);
or U11605 (N_11605,N_11049,N_11104);
xnor U11606 (N_11606,N_10965,N_10862);
or U11607 (N_11607,N_10828,N_11061);
or U11608 (N_11608,N_11276,N_10812);
nand U11609 (N_11609,N_11327,N_11161);
xnor U11610 (N_11610,N_11382,N_11085);
nor U11611 (N_11611,N_11354,N_11377);
nand U11612 (N_11612,N_11078,N_11126);
nand U11613 (N_11613,N_10974,N_11390);
nor U11614 (N_11614,N_10833,N_11106);
xor U11615 (N_11615,N_10811,N_11175);
or U11616 (N_11616,N_10849,N_11311);
nor U11617 (N_11617,N_11346,N_10814);
nand U11618 (N_11618,N_11232,N_11387);
xnor U11619 (N_11619,N_10940,N_11033);
and U11620 (N_11620,N_10887,N_10976);
or U11621 (N_11621,N_10929,N_10823);
nand U11622 (N_11622,N_11074,N_10971);
xor U11623 (N_11623,N_11158,N_11243);
and U11624 (N_11624,N_11351,N_11301);
xnor U11625 (N_11625,N_10893,N_10937);
xnor U11626 (N_11626,N_11305,N_11048);
xnor U11627 (N_11627,N_10809,N_11262);
nand U11628 (N_11628,N_11248,N_11263);
xnor U11629 (N_11629,N_11394,N_11075);
or U11630 (N_11630,N_11364,N_11001);
nand U11631 (N_11631,N_10942,N_10867);
nor U11632 (N_11632,N_11201,N_10827);
nand U11633 (N_11633,N_11282,N_11293);
and U11634 (N_11634,N_11095,N_11070);
nand U11635 (N_11635,N_11290,N_10866);
nand U11636 (N_11636,N_10967,N_11176);
nand U11637 (N_11637,N_11393,N_11065);
and U11638 (N_11638,N_11091,N_11012);
nor U11639 (N_11639,N_10894,N_11041);
nor U11640 (N_11640,N_11223,N_10922);
nor U11641 (N_11641,N_10848,N_11205);
and U11642 (N_11642,N_10949,N_11343);
nor U11643 (N_11643,N_10970,N_10917);
nand U11644 (N_11644,N_11193,N_11242);
and U11645 (N_11645,N_10991,N_11171);
or U11646 (N_11646,N_10916,N_11297);
xnor U11647 (N_11647,N_11383,N_10802);
nor U11648 (N_11648,N_11172,N_11039);
xnor U11649 (N_11649,N_11152,N_10885);
nor U11650 (N_11650,N_11114,N_11080);
and U11651 (N_11651,N_11344,N_11217);
xnor U11652 (N_11652,N_10864,N_11021);
nand U11653 (N_11653,N_11386,N_10878);
and U11654 (N_11654,N_11249,N_10969);
nand U11655 (N_11655,N_11042,N_11380);
nor U11656 (N_11656,N_11035,N_11142);
nand U11657 (N_11657,N_11216,N_11057);
nand U11658 (N_11658,N_11336,N_11141);
xor U11659 (N_11659,N_10800,N_10939);
and U11660 (N_11660,N_10844,N_10856);
nor U11661 (N_11661,N_11090,N_10898);
nand U11662 (N_11662,N_11000,N_11084);
or U11663 (N_11663,N_11003,N_10904);
or U11664 (N_11664,N_11302,N_11097);
nand U11665 (N_11665,N_11239,N_11391);
or U11666 (N_11666,N_11349,N_11261);
xor U11667 (N_11667,N_11069,N_10871);
nand U11668 (N_11668,N_11240,N_11348);
nor U11669 (N_11669,N_10980,N_11381);
nand U11670 (N_11670,N_11182,N_11096);
or U11671 (N_11671,N_11230,N_10978);
xor U11672 (N_11672,N_11215,N_11059);
xor U11673 (N_11673,N_11385,N_11064);
nand U11674 (N_11674,N_11244,N_11225);
nor U11675 (N_11675,N_11073,N_11149);
nand U11676 (N_11676,N_10892,N_11339);
nand U11677 (N_11677,N_11020,N_10995);
xor U11678 (N_11678,N_11199,N_10928);
nand U11679 (N_11679,N_11294,N_10953);
and U11680 (N_11680,N_11268,N_11333);
nand U11681 (N_11681,N_11226,N_11115);
xnor U11682 (N_11682,N_11374,N_11179);
xnor U11683 (N_11683,N_10955,N_11076);
xor U11684 (N_11684,N_11309,N_11256);
or U11685 (N_11685,N_11014,N_11068);
xor U11686 (N_11686,N_11324,N_10807);
xnor U11687 (N_11687,N_10963,N_10903);
or U11688 (N_11688,N_11133,N_10815);
xor U11689 (N_11689,N_10914,N_10918);
nand U11690 (N_11690,N_11246,N_11054);
nor U11691 (N_11691,N_10852,N_11031);
xor U11692 (N_11692,N_11103,N_11340);
and U11693 (N_11693,N_11253,N_11060);
nand U11694 (N_11694,N_11117,N_11384);
nand U11695 (N_11695,N_11328,N_11318);
nand U11696 (N_11696,N_11322,N_11192);
xor U11697 (N_11697,N_11113,N_10888);
xnor U11698 (N_11698,N_10932,N_11146);
xor U11699 (N_11699,N_11222,N_11366);
or U11700 (N_11700,N_11101,N_11117);
or U11701 (N_11701,N_10821,N_11157);
and U11702 (N_11702,N_10973,N_11381);
nand U11703 (N_11703,N_10900,N_10941);
nand U11704 (N_11704,N_10914,N_11219);
or U11705 (N_11705,N_11078,N_10946);
nand U11706 (N_11706,N_11301,N_10813);
and U11707 (N_11707,N_11232,N_11014);
or U11708 (N_11708,N_11160,N_11321);
nor U11709 (N_11709,N_11057,N_10966);
nor U11710 (N_11710,N_10857,N_10828);
or U11711 (N_11711,N_11330,N_10974);
and U11712 (N_11712,N_11217,N_11286);
and U11713 (N_11713,N_11009,N_10897);
or U11714 (N_11714,N_11284,N_11382);
or U11715 (N_11715,N_11381,N_11310);
or U11716 (N_11716,N_11006,N_11082);
and U11717 (N_11717,N_10845,N_11261);
or U11718 (N_11718,N_11247,N_11136);
nand U11719 (N_11719,N_11231,N_11001);
and U11720 (N_11720,N_10881,N_11314);
nand U11721 (N_11721,N_10935,N_11310);
and U11722 (N_11722,N_10911,N_11036);
nand U11723 (N_11723,N_11121,N_11302);
and U11724 (N_11724,N_11141,N_11262);
xnor U11725 (N_11725,N_11080,N_10885);
or U11726 (N_11726,N_10808,N_10882);
xnor U11727 (N_11727,N_10825,N_11308);
and U11728 (N_11728,N_11305,N_10917);
and U11729 (N_11729,N_11124,N_11217);
nand U11730 (N_11730,N_11059,N_11301);
and U11731 (N_11731,N_11040,N_10929);
nor U11732 (N_11732,N_11038,N_11299);
and U11733 (N_11733,N_10987,N_10886);
nor U11734 (N_11734,N_11048,N_10905);
and U11735 (N_11735,N_11305,N_10872);
xnor U11736 (N_11736,N_11266,N_11223);
xor U11737 (N_11737,N_10915,N_11359);
and U11738 (N_11738,N_11368,N_11327);
and U11739 (N_11739,N_11037,N_11121);
xor U11740 (N_11740,N_10811,N_11009);
nand U11741 (N_11741,N_11148,N_10902);
and U11742 (N_11742,N_11367,N_11329);
nor U11743 (N_11743,N_11062,N_11365);
nand U11744 (N_11744,N_11007,N_11141);
and U11745 (N_11745,N_11110,N_10903);
or U11746 (N_11746,N_10977,N_11125);
nor U11747 (N_11747,N_11013,N_11133);
and U11748 (N_11748,N_11266,N_11225);
nand U11749 (N_11749,N_11170,N_10990);
or U11750 (N_11750,N_11249,N_11271);
and U11751 (N_11751,N_11013,N_11246);
xnor U11752 (N_11752,N_11162,N_10897);
or U11753 (N_11753,N_11253,N_10938);
nor U11754 (N_11754,N_11032,N_11359);
nand U11755 (N_11755,N_10840,N_10904);
nand U11756 (N_11756,N_11131,N_11037);
and U11757 (N_11757,N_11257,N_11268);
and U11758 (N_11758,N_11383,N_11371);
or U11759 (N_11759,N_10814,N_11149);
and U11760 (N_11760,N_10954,N_11035);
and U11761 (N_11761,N_11150,N_11193);
and U11762 (N_11762,N_11275,N_10915);
and U11763 (N_11763,N_11079,N_11033);
nor U11764 (N_11764,N_11214,N_10928);
nand U11765 (N_11765,N_11071,N_11204);
and U11766 (N_11766,N_10853,N_11169);
nand U11767 (N_11767,N_11170,N_11381);
or U11768 (N_11768,N_11265,N_11134);
xor U11769 (N_11769,N_10940,N_11083);
or U11770 (N_11770,N_10873,N_11114);
nor U11771 (N_11771,N_10905,N_10801);
or U11772 (N_11772,N_10975,N_10940);
or U11773 (N_11773,N_10995,N_11155);
xor U11774 (N_11774,N_10914,N_11109);
xnor U11775 (N_11775,N_11369,N_11307);
nor U11776 (N_11776,N_11151,N_10999);
nor U11777 (N_11777,N_11286,N_11227);
and U11778 (N_11778,N_11256,N_11003);
nor U11779 (N_11779,N_11167,N_11009);
nand U11780 (N_11780,N_11279,N_11148);
or U11781 (N_11781,N_11068,N_11011);
nor U11782 (N_11782,N_11262,N_10917);
xnor U11783 (N_11783,N_10921,N_11387);
and U11784 (N_11784,N_11133,N_11372);
nand U11785 (N_11785,N_11393,N_11043);
nor U11786 (N_11786,N_11368,N_11197);
xnor U11787 (N_11787,N_10816,N_10919);
or U11788 (N_11788,N_10816,N_11034);
and U11789 (N_11789,N_10959,N_10858);
nand U11790 (N_11790,N_11173,N_10843);
nand U11791 (N_11791,N_11036,N_11216);
and U11792 (N_11792,N_10877,N_11102);
nor U11793 (N_11793,N_10855,N_11021);
and U11794 (N_11794,N_10816,N_11298);
xnor U11795 (N_11795,N_11222,N_11288);
or U11796 (N_11796,N_10999,N_10914);
nand U11797 (N_11797,N_10861,N_11231);
nand U11798 (N_11798,N_11092,N_11008);
nor U11799 (N_11799,N_11169,N_10995);
nand U11800 (N_11800,N_11355,N_10961);
nand U11801 (N_11801,N_10930,N_11258);
nand U11802 (N_11802,N_10848,N_10834);
or U11803 (N_11803,N_10886,N_11139);
nand U11804 (N_11804,N_10804,N_11389);
nor U11805 (N_11805,N_11394,N_11162);
nor U11806 (N_11806,N_10903,N_11089);
nand U11807 (N_11807,N_11015,N_11273);
xnor U11808 (N_11808,N_10952,N_10850);
nor U11809 (N_11809,N_11346,N_11344);
nor U11810 (N_11810,N_11190,N_11221);
nand U11811 (N_11811,N_11265,N_11173);
nand U11812 (N_11812,N_11099,N_11111);
xnor U11813 (N_11813,N_11328,N_11268);
nand U11814 (N_11814,N_10930,N_10847);
nand U11815 (N_11815,N_11199,N_11210);
and U11816 (N_11816,N_11200,N_11149);
nand U11817 (N_11817,N_11115,N_11160);
nand U11818 (N_11818,N_11234,N_11314);
and U11819 (N_11819,N_10950,N_11041);
and U11820 (N_11820,N_10968,N_11337);
and U11821 (N_11821,N_11212,N_10875);
nor U11822 (N_11822,N_10989,N_11188);
xor U11823 (N_11823,N_10976,N_11242);
xnor U11824 (N_11824,N_10968,N_11156);
nor U11825 (N_11825,N_11327,N_11057);
xnor U11826 (N_11826,N_10904,N_10857);
nor U11827 (N_11827,N_11341,N_10834);
nand U11828 (N_11828,N_10938,N_11111);
nand U11829 (N_11829,N_11044,N_11342);
or U11830 (N_11830,N_11102,N_11109);
and U11831 (N_11831,N_10968,N_11109);
or U11832 (N_11832,N_10965,N_11009);
and U11833 (N_11833,N_11159,N_11241);
or U11834 (N_11834,N_10945,N_11056);
nand U11835 (N_11835,N_11319,N_11130);
xnor U11836 (N_11836,N_10808,N_10950);
xnor U11837 (N_11837,N_11134,N_11025);
nand U11838 (N_11838,N_10930,N_11063);
and U11839 (N_11839,N_10814,N_10891);
nor U11840 (N_11840,N_11042,N_10935);
and U11841 (N_11841,N_11131,N_10801);
nor U11842 (N_11842,N_11159,N_11278);
and U11843 (N_11843,N_11270,N_10814);
and U11844 (N_11844,N_10829,N_10927);
and U11845 (N_11845,N_10829,N_11076);
xnor U11846 (N_11846,N_11347,N_11067);
nand U11847 (N_11847,N_10867,N_11006);
or U11848 (N_11848,N_10884,N_11021);
nand U11849 (N_11849,N_11059,N_11315);
or U11850 (N_11850,N_11340,N_11283);
or U11851 (N_11851,N_10902,N_11306);
or U11852 (N_11852,N_11006,N_11055);
nand U11853 (N_11853,N_11280,N_10884);
xnor U11854 (N_11854,N_11270,N_11238);
nand U11855 (N_11855,N_11334,N_11271);
nor U11856 (N_11856,N_10961,N_10986);
nor U11857 (N_11857,N_10964,N_10963);
or U11858 (N_11858,N_11183,N_11056);
xnor U11859 (N_11859,N_11088,N_10933);
nor U11860 (N_11860,N_11028,N_11391);
xor U11861 (N_11861,N_11241,N_10815);
nand U11862 (N_11862,N_11319,N_11079);
xor U11863 (N_11863,N_11053,N_11349);
and U11864 (N_11864,N_10869,N_10981);
nand U11865 (N_11865,N_11104,N_11088);
nand U11866 (N_11866,N_10910,N_10900);
nor U11867 (N_11867,N_10946,N_11166);
and U11868 (N_11868,N_11302,N_10878);
xor U11869 (N_11869,N_11040,N_11392);
nor U11870 (N_11870,N_11003,N_11377);
or U11871 (N_11871,N_10924,N_11055);
nor U11872 (N_11872,N_11203,N_11247);
or U11873 (N_11873,N_10839,N_10810);
nand U11874 (N_11874,N_10975,N_11196);
nor U11875 (N_11875,N_10808,N_11087);
xnor U11876 (N_11876,N_10917,N_11356);
nor U11877 (N_11877,N_11009,N_11121);
nor U11878 (N_11878,N_10820,N_11354);
nor U11879 (N_11879,N_10951,N_11093);
xor U11880 (N_11880,N_11134,N_11230);
nor U11881 (N_11881,N_11112,N_11151);
nor U11882 (N_11882,N_10928,N_11238);
nand U11883 (N_11883,N_10974,N_11085);
or U11884 (N_11884,N_11338,N_11154);
or U11885 (N_11885,N_11154,N_11145);
xor U11886 (N_11886,N_10832,N_11057);
nor U11887 (N_11887,N_11298,N_10925);
or U11888 (N_11888,N_10819,N_11054);
and U11889 (N_11889,N_10874,N_11175);
or U11890 (N_11890,N_10939,N_10964);
nor U11891 (N_11891,N_11346,N_11063);
nand U11892 (N_11892,N_11334,N_11261);
and U11893 (N_11893,N_11202,N_10978);
and U11894 (N_11894,N_10894,N_11269);
xnor U11895 (N_11895,N_11230,N_11141);
xnor U11896 (N_11896,N_11260,N_10819);
or U11897 (N_11897,N_10972,N_11050);
nand U11898 (N_11898,N_11025,N_10807);
and U11899 (N_11899,N_11132,N_10876);
and U11900 (N_11900,N_11274,N_11318);
and U11901 (N_11901,N_10944,N_11183);
nor U11902 (N_11902,N_10882,N_11381);
nor U11903 (N_11903,N_10915,N_10846);
nor U11904 (N_11904,N_10980,N_10864);
nand U11905 (N_11905,N_11274,N_11039);
nor U11906 (N_11906,N_10884,N_10907);
or U11907 (N_11907,N_11200,N_11368);
or U11908 (N_11908,N_11086,N_10989);
nand U11909 (N_11909,N_10967,N_11328);
nor U11910 (N_11910,N_10964,N_11044);
nand U11911 (N_11911,N_11088,N_11099);
nor U11912 (N_11912,N_11006,N_11350);
xor U11913 (N_11913,N_10942,N_10959);
or U11914 (N_11914,N_10998,N_10856);
nor U11915 (N_11915,N_11216,N_11061);
nor U11916 (N_11916,N_10922,N_11040);
nor U11917 (N_11917,N_11350,N_11388);
xnor U11918 (N_11918,N_11254,N_11348);
xnor U11919 (N_11919,N_10812,N_11392);
nor U11920 (N_11920,N_11036,N_10861);
nor U11921 (N_11921,N_11398,N_11082);
and U11922 (N_11922,N_11243,N_11127);
nand U11923 (N_11923,N_11252,N_10983);
xnor U11924 (N_11924,N_10832,N_11225);
and U11925 (N_11925,N_10847,N_11146);
xnor U11926 (N_11926,N_10944,N_11110);
xor U11927 (N_11927,N_11227,N_11288);
nand U11928 (N_11928,N_11237,N_10844);
nand U11929 (N_11929,N_11088,N_11334);
and U11930 (N_11930,N_11164,N_11204);
nor U11931 (N_11931,N_11139,N_10979);
nand U11932 (N_11932,N_10850,N_10976);
xor U11933 (N_11933,N_11260,N_10924);
or U11934 (N_11934,N_11023,N_10869);
or U11935 (N_11935,N_11342,N_11048);
or U11936 (N_11936,N_11388,N_11276);
nand U11937 (N_11937,N_10972,N_10965);
or U11938 (N_11938,N_11106,N_10999);
or U11939 (N_11939,N_11063,N_11046);
and U11940 (N_11940,N_11299,N_10819);
nand U11941 (N_11941,N_11328,N_10959);
and U11942 (N_11942,N_10951,N_11329);
and U11943 (N_11943,N_11059,N_11174);
and U11944 (N_11944,N_11352,N_10846);
xor U11945 (N_11945,N_11338,N_11140);
and U11946 (N_11946,N_10995,N_11292);
nor U11947 (N_11947,N_10896,N_11267);
or U11948 (N_11948,N_10859,N_11252);
and U11949 (N_11949,N_11313,N_11176);
xor U11950 (N_11950,N_11106,N_11134);
xor U11951 (N_11951,N_11113,N_11118);
or U11952 (N_11952,N_10984,N_11313);
xor U11953 (N_11953,N_11135,N_11184);
xor U11954 (N_11954,N_11069,N_10824);
nand U11955 (N_11955,N_11157,N_11152);
nand U11956 (N_11956,N_11236,N_10969);
nor U11957 (N_11957,N_11316,N_10853);
nor U11958 (N_11958,N_11193,N_11022);
and U11959 (N_11959,N_11306,N_10849);
nand U11960 (N_11960,N_10980,N_11304);
and U11961 (N_11961,N_11256,N_11327);
nand U11962 (N_11962,N_11100,N_11019);
nand U11963 (N_11963,N_11270,N_10815);
nand U11964 (N_11964,N_11216,N_11264);
nor U11965 (N_11965,N_11303,N_11340);
xnor U11966 (N_11966,N_11071,N_11327);
nor U11967 (N_11967,N_10954,N_10810);
nor U11968 (N_11968,N_11255,N_10852);
xnor U11969 (N_11969,N_11113,N_10816);
nor U11970 (N_11970,N_11144,N_11309);
nand U11971 (N_11971,N_11199,N_10988);
xnor U11972 (N_11972,N_11172,N_10931);
nand U11973 (N_11973,N_10960,N_11204);
nand U11974 (N_11974,N_11032,N_11327);
and U11975 (N_11975,N_11236,N_10921);
or U11976 (N_11976,N_11223,N_10902);
xor U11977 (N_11977,N_11121,N_11284);
or U11978 (N_11978,N_11394,N_10980);
xor U11979 (N_11979,N_11145,N_11237);
xor U11980 (N_11980,N_10813,N_11321);
nand U11981 (N_11981,N_11350,N_11133);
or U11982 (N_11982,N_11011,N_11390);
nor U11983 (N_11983,N_11268,N_11378);
and U11984 (N_11984,N_10887,N_11167);
or U11985 (N_11985,N_11287,N_10820);
nor U11986 (N_11986,N_11171,N_11086);
nand U11987 (N_11987,N_11381,N_10843);
xor U11988 (N_11988,N_10995,N_11310);
nand U11989 (N_11989,N_11343,N_11103);
or U11990 (N_11990,N_10915,N_10879);
or U11991 (N_11991,N_11090,N_10807);
nand U11992 (N_11992,N_11205,N_10813);
xor U11993 (N_11993,N_11204,N_11130);
nor U11994 (N_11994,N_11246,N_11323);
xnor U11995 (N_11995,N_11029,N_10919);
and U11996 (N_11996,N_10891,N_10903);
nand U11997 (N_11997,N_10897,N_10942);
and U11998 (N_11998,N_11128,N_11090);
xor U11999 (N_11999,N_10861,N_11200);
and U12000 (N_12000,N_11710,N_11676);
or U12001 (N_12001,N_11974,N_11601);
nor U12002 (N_12002,N_11733,N_11589);
nand U12003 (N_12003,N_11923,N_11559);
or U12004 (N_12004,N_11585,N_11877);
or U12005 (N_12005,N_11813,N_11908);
xnor U12006 (N_12006,N_11883,N_11749);
nor U12007 (N_12007,N_11999,N_11555);
or U12008 (N_12008,N_11568,N_11567);
xor U12009 (N_12009,N_11497,N_11916);
xnor U12010 (N_12010,N_11899,N_11564);
nand U12011 (N_12011,N_11863,N_11487);
or U12012 (N_12012,N_11981,N_11469);
and U12013 (N_12013,N_11410,N_11951);
nand U12014 (N_12014,N_11884,N_11898);
xnor U12015 (N_12015,N_11722,N_11540);
nor U12016 (N_12016,N_11965,N_11505);
nand U12017 (N_12017,N_11569,N_11551);
nand U12018 (N_12018,N_11699,N_11897);
and U12019 (N_12019,N_11616,N_11962);
nor U12020 (N_12020,N_11546,N_11489);
nand U12021 (N_12021,N_11550,N_11707);
or U12022 (N_12022,N_11495,N_11641);
and U12023 (N_12023,N_11583,N_11693);
nand U12024 (N_12024,N_11642,N_11434);
and U12025 (N_12025,N_11956,N_11742);
nand U12026 (N_12026,N_11486,N_11932);
nor U12027 (N_12027,N_11724,N_11440);
and U12028 (N_12028,N_11781,N_11779);
or U12029 (N_12029,N_11826,N_11920);
xor U12030 (N_12030,N_11598,N_11459);
and U12031 (N_12031,N_11620,N_11480);
and U12032 (N_12032,N_11558,N_11772);
nor U12033 (N_12033,N_11905,N_11771);
nor U12034 (N_12034,N_11844,N_11514);
or U12035 (N_12035,N_11995,N_11515);
and U12036 (N_12036,N_11873,N_11457);
or U12037 (N_12037,N_11741,N_11802);
nor U12038 (N_12038,N_11785,N_11572);
and U12039 (N_12039,N_11869,N_11740);
nand U12040 (N_12040,N_11437,N_11491);
nor U12041 (N_12041,N_11453,N_11987);
nor U12042 (N_12042,N_11586,N_11580);
and U12043 (N_12043,N_11891,N_11937);
nand U12044 (N_12044,N_11870,N_11861);
and U12045 (N_12045,N_11958,N_11425);
nand U12046 (N_12046,N_11872,N_11827);
nor U12047 (N_12047,N_11684,N_11853);
nand U12048 (N_12048,N_11709,N_11788);
xor U12049 (N_12049,N_11618,N_11566);
nand U12050 (N_12050,N_11720,N_11747);
xor U12051 (N_12051,N_11454,N_11886);
xnor U12052 (N_12052,N_11815,N_11881);
nor U12053 (N_12053,N_11744,N_11966);
or U12054 (N_12054,N_11413,N_11824);
nor U12055 (N_12055,N_11483,N_11681);
and U12056 (N_12056,N_11573,N_11516);
xnor U12057 (N_12057,N_11603,N_11982);
nand U12058 (N_12058,N_11832,N_11766);
nand U12059 (N_12059,N_11426,N_11512);
or U12060 (N_12060,N_11474,N_11996);
nand U12061 (N_12061,N_11765,N_11810);
xor U12062 (N_12062,N_11860,N_11544);
xor U12063 (N_12063,N_11612,N_11754);
nand U12064 (N_12064,N_11675,N_11424);
or U12065 (N_12065,N_11432,N_11461);
xor U12066 (N_12066,N_11695,N_11809);
and U12067 (N_12067,N_11475,N_11455);
or U12068 (N_12068,N_11798,N_11614);
or U12069 (N_12069,N_11757,N_11721);
xnor U12070 (N_12070,N_11470,N_11677);
or U12071 (N_12071,N_11581,N_11975);
nor U12072 (N_12072,N_11760,N_11792);
nand U12073 (N_12073,N_11660,N_11683);
and U12074 (N_12074,N_11420,N_11859);
and U12075 (N_12075,N_11602,N_11935);
xor U12076 (N_12076,N_11793,N_11763);
xnor U12077 (N_12077,N_11423,N_11993);
and U12078 (N_12078,N_11851,N_11864);
or U12079 (N_12079,N_11625,N_11593);
and U12080 (N_12080,N_11629,N_11626);
or U12081 (N_12081,N_11630,N_11472);
and U12082 (N_12082,N_11926,N_11592);
and U12083 (N_12083,N_11452,N_11922);
xnor U12084 (N_12084,N_11431,N_11837);
and U12085 (N_12085,N_11727,N_11790);
or U12086 (N_12086,N_11704,N_11449);
xnor U12087 (N_12087,N_11825,N_11979);
nor U12088 (N_12088,N_11617,N_11686);
nand U12089 (N_12089,N_11823,N_11488);
nand U12090 (N_12090,N_11854,N_11415);
and U12091 (N_12091,N_11575,N_11600);
nor U12092 (N_12092,N_11541,N_11622);
and U12093 (N_12093,N_11715,N_11998);
nor U12094 (N_12094,N_11759,N_11441);
nor U12095 (N_12095,N_11403,N_11621);
nor U12096 (N_12096,N_11443,N_11820);
nor U12097 (N_12097,N_11698,N_11439);
nor U12098 (N_12098,N_11549,N_11914);
and U12099 (N_12099,N_11490,N_11682);
xor U12100 (N_12100,N_11588,N_11624);
xnor U12101 (N_12101,N_11756,N_11892);
and U12102 (N_12102,N_11828,N_11991);
and U12103 (N_12103,N_11796,N_11786);
nor U12104 (N_12104,N_11421,N_11503);
xor U12105 (N_12105,N_11963,N_11866);
nor U12106 (N_12106,N_11534,N_11697);
and U12107 (N_12107,N_11977,N_11604);
xor U12108 (N_12108,N_11918,N_11730);
or U12109 (N_12109,N_11731,N_11942);
or U12110 (N_12110,N_11755,N_11562);
xor U12111 (N_12111,N_11606,N_11406);
xnor U12112 (N_12112,N_11723,N_11670);
xor U12113 (N_12113,N_11578,N_11554);
xnor U12114 (N_12114,N_11738,N_11502);
xnor U12115 (N_12115,N_11875,N_11791);
nand U12116 (N_12116,N_11584,N_11808);
xnor U12117 (N_12117,N_11692,N_11985);
and U12118 (N_12118,N_11553,N_11811);
nor U12119 (N_12119,N_11649,N_11969);
nor U12120 (N_12120,N_11430,N_11753);
nor U12121 (N_12121,N_11735,N_11822);
nor U12122 (N_12122,N_11547,N_11419);
xor U12123 (N_12123,N_11978,N_11679);
nor U12124 (N_12124,N_11911,N_11463);
xnor U12125 (N_12125,N_11662,N_11961);
nand U12126 (N_12126,N_11527,N_11468);
or U12127 (N_12127,N_11532,N_11464);
nand U12128 (N_12128,N_11973,N_11764);
nand U12129 (N_12129,N_11852,N_11835);
and U12130 (N_12130,N_11451,N_11673);
and U12131 (N_12131,N_11513,N_11448);
nor U12132 (N_12132,N_11506,N_11518);
or U12133 (N_12133,N_11543,N_11739);
and U12134 (N_12134,N_11719,N_11849);
nand U12135 (N_12135,N_11680,N_11652);
and U12136 (N_12136,N_11640,N_11725);
or U12137 (N_12137,N_11526,N_11499);
and U12138 (N_12138,N_11609,N_11889);
nor U12139 (N_12139,N_11645,N_11557);
and U12140 (N_12140,N_11800,N_11646);
nand U12141 (N_12141,N_11501,N_11596);
nor U12142 (N_12142,N_11767,N_11623);
and U12143 (N_12143,N_11444,N_11632);
nor U12144 (N_12144,N_11666,N_11797);
nor U12145 (N_12145,N_11538,N_11433);
xnor U12146 (N_12146,N_11903,N_11819);
xnor U12147 (N_12147,N_11970,N_11874);
nand U12148 (N_12148,N_11561,N_11481);
and U12149 (N_12149,N_11591,N_11711);
or U12150 (N_12150,N_11988,N_11737);
nor U12151 (N_12151,N_11984,N_11768);
nand U12152 (N_12152,N_11647,N_11634);
nor U12153 (N_12153,N_11804,N_11436);
xnor U12154 (N_12154,N_11701,N_11934);
and U12155 (N_12155,N_11523,N_11530);
and U12156 (N_12156,N_11658,N_11599);
nor U12157 (N_12157,N_11967,N_11989);
xnor U12158 (N_12158,N_11460,N_11597);
nand U12159 (N_12159,N_11847,N_11947);
nand U12160 (N_12160,N_11894,N_11577);
xor U12161 (N_12161,N_11838,N_11845);
nor U12162 (N_12162,N_11980,N_11493);
and U12163 (N_12163,N_11776,N_11638);
and U12164 (N_12164,N_11840,N_11885);
and U12165 (N_12165,N_11478,N_11836);
nand U12166 (N_12166,N_11446,N_11972);
and U12167 (N_12167,N_11777,N_11643);
xnor U12168 (N_12168,N_11829,N_11705);
or U12169 (N_12169,N_11949,N_11528);
nand U12170 (N_12170,N_11678,N_11848);
and U12171 (N_12171,N_11450,N_11648);
xor U12172 (N_12172,N_11971,N_11445);
nor U12173 (N_12173,N_11834,N_11594);
xor U12174 (N_12174,N_11587,N_11990);
nand U12175 (N_12175,N_11465,N_11563);
nand U12176 (N_12176,N_11535,N_11539);
nand U12177 (N_12177,N_11611,N_11917);
nand U12178 (N_12178,N_11841,N_11896);
xnor U12179 (N_12179,N_11651,N_11613);
nor U12180 (N_12180,N_11782,N_11895);
xor U12181 (N_12181,N_11494,N_11628);
nand U12182 (N_12182,N_11936,N_11477);
nand U12183 (N_12183,N_11983,N_11830);
or U12184 (N_12184,N_11761,N_11952);
nand U12185 (N_12185,N_11924,N_11579);
or U12186 (N_12186,N_11882,N_11812);
nor U12187 (N_12187,N_11565,N_11750);
and U12188 (N_12188,N_11930,N_11479);
and U12189 (N_12189,N_11939,N_11659);
or U12190 (N_12190,N_11655,N_11462);
nand U12191 (N_12191,N_11644,N_11664);
or U12192 (N_12192,N_11703,N_11950);
nor U12193 (N_12193,N_11510,N_11411);
or U12194 (N_12194,N_11960,N_11954);
xnor U12195 (N_12195,N_11904,N_11504);
and U12196 (N_12196,N_11857,N_11780);
nor U12197 (N_12197,N_11574,N_11933);
or U12198 (N_12198,N_11878,N_11524);
xor U12199 (N_12199,N_11778,N_11787);
nor U12200 (N_12200,N_11856,N_11795);
and U12201 (N_12201,N_11615,N_11751);
nor U12202 (N_12202,N_11467,N_11672);
nand U12203 (N_12203,N_11605,N_11746);
or U12204 (N_12204,N_11729,N_11893);
or U12205 (N_12205,N_11633,N_11702);
nor U12206 (N_12206,N_11783,N_11656);
xor U12207 (N_12207,N_11485,N_11531);
nand U12208 (N_12208,N_11803,N_11748);
nor U12209 (N_12209,N_11818,N_11955);
nand U12210 (N_12210,N_11435,N_11831);
nand U12211 (N_12211,N_11608,N_11921);
nand U12212 (N_12212,N_11429,N_11508);
nor U12213 (N_12213,N_11769,N_11595);
xnor U12214 (N_12214,N_11520,N_11986);
xnor U12215 (N_12215,N_11850,N_11405);
nand U12216 (N_12216,N_11862,N_11519);
or U12217 (N_12217,N_11968,N_11401);
nor U12218 (N_12218,N_11789,N_11799);
xnor U12219 (N_12219,N_11694,N_11417);
nand U12220 (N_12220,N_11442,N_11957);
nor U12221 (N_12221,N_11758,N_11507);
and U12222 (N_12222,N_11627,N_11654);
and U12223 (N_12223,N_11521,N_11402);
nor U12224 (N_12224,N_11700,N_11696);
nand U12225 (N_12225,N_11533,N_11552);
or U12226 (N_12226,N_11471,N_11687);
xnor U12227 (N_12227,N_11713,N_11484);
nand U12228 (N_12228,N_11639,N_11428);
nor U12229 (N_12229,N_11888,N_11807);
and U12230 (N_12230,N_11691,N_11925);
nor U12231 (N_12231,N_11560,N_11964);
nor U12232 (N_12232,N_11665,N_11548);
and U12233 (N_12233,N_11941,N_11498);
nand U12234 (N_12234,N_11536,N_11846);
nand U12235 (N_12235,N_11653,N_11714);
and U12236 (N_12236,N_11466,N_11674);
nand U12237 (N_12237,N_11473,N_11931);
or U12238 (N_12238,N_11945,N_11953);
or U12239 (N_12239,N_11492,N_11938);
xnor U12240 (N_12240,N_11529,N_11948);
nand U12241 (N_12241,N_11805,N_11690);
nand U12242 (N_12242,N_11773,N_11631);
nand U12243 (N_12243,N_11912,N_11901);
or U12244 (N_12244,N_11910,N_11590);
or U12245 (N_12245,N_11671,N_11400);
xnor U12246 (N_12246,N_11661,N_11887);
or U12247 (N_12247,N_11814,N_11706);
xnor U12248 (N_12248,N_11794,N_11708);
nand U12249 (N_12249,N_11775,N_11556);
xor U12250 (N_12250,N_11865,N_11734);
xnor U12251 (N_12251,N_11716,N_11839);
or U12252 (N_12252,N_11517,N_11929);
xnor U12253 (N_12253,N_11992,N_11511);
and U12254 (N_12254,N_11855,N_11635);
xor U12255 (N_12255,N_11743,N_11582);
nor U12256 (N_12256,N_11416,N_11610);
nand U12257 (N_12257,N_11688,N_11427);
or U12258 (N_12258,N_11762,N_11657);
and U12259 (N_12259,N_11685,N_11907);
xor U12260 (N_12260,N_11959,N_11736);
nor U12261 (N_12261,N_11456,N_11571);
nand U12262 (N_12262,N_11928,N_11636);
nor U12263 (N_12263,N_11770,N_11919);
nand U12264 (N_12264,N_11717,N_11868);
nand U12265 (N_12265,N_11774,N_11496);
or U12266 (N_12266,N_11900,N_11407);
nand U12267 (N_12267,N_11458,N_11879);
and U12268 (N_12268,N_11669,N_11906);
or U12269 (N_12269,N_11576,N_11545);
xor U12270 (N_12270,N_11607,N_11732);
or U12271 (N_12271,N_11537,N_11806);
xor U12272 (N_12272,N_11525,N_11909);
xnor U12273 (N_12273,N_11689,N_11843);
nand U12274 (N_12274,N_11418,N_11902);
nor U12275 (N_12275,N_11943,N_11858);
nand U12276 (N_12276,N_11500,N_11976);
xor U12277 (N_12277,N_11667,N_11663);
nand U12278 (N_12278,N_11871,N_11570);
or U12279 (N_12279,N_11522,N_11509);
nand U12280 (N_12280,N_11997,N_11842);
and U12281 (N_12281,N_11409,N_11816);
or U12282 (N_12282,N_11817,N_11637);
nor U12283 (N_12283,N_11784,N_11482);
nor U12284 (N_12284,N_11726,N_11833);
nor U12285 (N_12285,N_11712,N_11821);
xor U12286 (N_12286,N_11745,N_11876);
nand U12287 (N_12287,N_11668,N_11867);
nand U12288 (N_12288,N_11408,N_11946);
or U12289 (N_12289,N_11927,N_11404);
nand U12290 (N_12290,N_11447,N_11915);
nand U12291 (N_12291,N_11438,N_11944);
nor U12292 (N_12292,N_11542,N_11422);
and U12293 (N_12293,N_11412,N_11801);
xnor U12294 (N_12294,N_11890,N_11650);
nand U12295 (N_12295,N_11752,N_11414);
or U12296 (N_12296,N_11940,N_11880);
nor U12297 (N_12297,N_11476,N_11718);
nor U12298 (N_12298,N_11728,N_11619);
and U12299 (N_12299,N_11913,N_11994);
xnor U12300 (N_12300,N_11621,N_11882);
nor U12301 (N_12301,N_11794,N_11795);
and U12302 (N_12302,N_11529,N_11821);
xor U12303 (N_12303,N_11736,N_11521);
and U12304 (N_12304,N_11500,N_11948);
or U12305 (N_12305,N_11692,N_11880);
nand U12306 (N_12306,N_11592,N_11430);
or U12307 (N_12307,N_11850,N_11911);
xor U12308 (N_12308,N_11721,N_11870);
nand U12309 (N_12309,N_11985,N_11992);
or U12310 (N_12310,N_11760,N_11958);
xnor U12311 (N_12311,N_11781,N_11575);
or U12312 (N_12312,N_11652,N_11738);
nor U12313 (N_12313,N_11574,N_11694);
xor U12314 (N_12314,N_11793,N_11830);
xor U12315 (N_12315,N_11424,N_11999);
nand U12316 (N_12316,N_11737,N_11552);
xor U12317 (N_12317,N_11640,N_11938);
nor U12318 (N_12318,N_11990,N_11775);
or U12319 (N_12319,N_11577,N_11759);
or U12320 (N_12320,N_11724,N_11880);
xor U12321 (N_12321,N_11984,N_11614);
xnor U12322 (N_12322,N_11417,N_11994);
or U12323 (N_12323,N_11578,N_11450);
nand U12324 (N_12324,N_11743,N_11929);
xnor U12325 (N_12325,N_11630,N_11868);
nor U12326 (N_12326,N_11449,N_11484);
nor U12327 (N_12327,N_11845,N_11676);
and U12328 (N_12328,N_11688,N_11794);
xnor U12329 (N_12329,N_11808,N_11966);
nand U12330 (N_12330,N_11685,N_11985);
nor U12331 (N_12331,N_11647,N_11753);
nor U12332 (N_12332,N_11432,N_11708);
or U12333 (N_12333,N_11466,N_11809);
nand U12334 (N_12334,N_11559,N_11669);
nand U12335 (N_12335,N_11493,N_11429);
xor U12336 (N_12336,N_11866,N_11674);
nand U12337 (N_12337,N_11626,N_11794);
xor U12338 (N_12338,N_11407,N_11541);
nor U12339 (N_12339,N_11610,N_11739);
nor U12340 (N_12340,N_11527,N_11771);
nand U12341 (N_12341,N_11754,N_11830);
or U12342 (N_12342,N_11807,N_11752);
xnor U12343 (N_12343,N_11449,N_11974);
nand U12344 (N_12344,N_11416,N_11783);
or U12345 (N_12345,N_11824,N_11605);
and U12346 (N_12346,N_11567,N_11770);
xnor U12347 (N_12347,N_11727,N_11704);
or U12348 (N_12348,N_11832,N_11636);
nor U12349 (N_12349,N_11816,N_11660);
and U12350 (N_12350,N_11423,N_11478);
nor U12351 (N_12351,N_11857,N_11730);
nor U12352 (N_12352,N_11545,N_11493);
and U12353 (N_12353,N_11881,N_11576);
nand U12354 (N_12354,N_11949,N_11903);
nand U12355 (N_12355,N_11670,N_11881);
and U12356 (N_12356,N_11601,N_11831);
nor U12357 (N_12357,N_11732,N_11452);
or U12358 (N_12358,N_11649,N_11446);
or U12359 (N_12359,N_11725,N_11785);
nor U12360 (N_12360,N_11812,N_11456);
nor U12361 (N_12361,N_11582,N_11904);
nand U12362 (N_12362,N_11489,N_11941);
and U12363 (N_12363,N_11429,N_11441);
nor U12364 (N_12364,N_11761,N_11515);
and U12365 (N_12365,N_11668,N_11989);
nand U12366 (N_12366,N_11983,N_11437);
nand U12367 (N_12367,N_11872,N_11530);
xnor U12368 (N_12368,N_11641,N_11581);
and U12369 (N_12369,N_11458,N_11824);
nand U12370 (N_12370,N_11600,N_11557);
and U12371 (N_12371,N_11432,N_11930);
nand U12372 (N_12372,N_11748,N_11508);
or U12373 (N_12373,N_11937,N_11569);
xor U12374 (N_12374,N_11539,N_11885);
and U12375 (N_12375,N_11794,N_11648);
nand U12376 (N_12376,N_11754,N_11978);
and U12377 (N_12377,N_11650,N_11412);
xnor U12378 (N_12378,N_11426,N_11891);
xor U12379 (N_12379,N_11848,N_11413);
xor U12380 (N_12380,N_11572,N_11717);
xor U12381 (N_12381,N_11955,N_11786);
nand U12382 (N_12382,N_11539,N_11915);
nor U12383 (N_12383,N_11704,N_11607);
or U12384 (N_12384,N_11646,N_11523);
nor U12385 (N_12385,N_11813,N_11791);
or U12386 (N_12386,N_11420,N_11886);
or U12387 (N_12387,N_11746,N_11775);
nand U12388 (N_12388,N_11653,N_11410);
or U12389 (N_12389,N_11827,N_11632);
nor U12390 (N_12390,N_11776,N_11601);
nand U12391 (N_12391,N_11705,N_11860);
and U12392 (N_12392,N_11664,N_11656);
and U12393 (N_12393,N_11721,N_11569);
and U12394 (N_12394,N_11666,N_11814);
nand U12395 (N_12395,N_11546,N_11793);
xor U12396 (N_12396,N_11762,N_11420);
nor U12397 (N_12397,N_11826,N_11839);
nand U12398 (N_12398,N_11776,N_11805);
nand U12399 (N_12399,N_11583,N_11644);
nand U12400 (N_12400,N_11705,N_11750);
nand U12401 (N_12401,N_11750,N_11980);
nor U12402 (N_12402,N_11529,N_11671);
nor U12403 (N_12403,N_11830,N_11995);
or U12404 (N_12404,N_11860,N_11563);
and U12405 (N_12405,N_11632,N_11494);
and U12406 (N_12406,N_11904,N_11518);
nand U12407 (N_12407,N_11867,N_11865);
nor U12408 (N_12408,N_11954,N_11577);
and U12409 (N_12409,N_11803,N_11400);
or U12410 (N_12410,N_11971,N_11843);
xor U12411 (N_12411,N_11735,N_11962);
or U12412 (N_12412,N_11419,N_11785);
and U12413 (N_12413,N_11716,N_11510);
nand U12414 (N_12414,N_11816,N_11794);
xor U12415 (N_12415,N_11792,N_11630);
and U12416 (N_12416,N_11613,N_11818);
or U12417 (N_12417,N_11556,N_11618);
nand U12418 (N_12418,N_11705,N_11876);
nor U12419 (N_12419,N_11639,N_11618);
and U12420 (N_12420,N_11705,N_11707);
nor U12421 (N_12421,N_11549,N_11578);
nor U12422 (N_12422,N_11470,N_11781);
xnor U12423 (N_12423,N_11671,N_11428);
xnor U12424 (N_12424,N_11905,N_11574);
nand U12425 (N_12425,N_11731,N_11474);
and U12426 (N_12426,N_11563,N_11549);
nor U12427 (N_12427,N_11713,N_11893);
nand U12428 (N_12428,N_11977,N_11575);
xor U12429 (N_12429,N_11421,N_11984);
xor U12430 (N_12430,N_11992,N_11659);
and U12431 (N_12431,N_11533,N_11971);
xnor U12432 (N_12432,N_11731,N_11409);
nand U12433 (N_12433,N_11424,N_11680);
xnor U12434 (N_12434,N_11531,N_11856);
xor U12435 (N_12435,N_11412,N_11509);
nand U12436 (N_12436,N_11847,N_11729);
and U12437 (N_12437,N_11974,N_11635);
xnor U12438 (N_12438,N_11907,N_11521);
nor U12439 (N_12439,N_11577,N_11825);
nor U12440 (N_12440,N_11994,N_11479);
or U12441 (N_12441,N_11688,N_11683);
and U12442 (N_12442,N_11493,N_11526);
or U12443 (N_12443,N_11663,N_11749);
and U12444 (N_12444,N_11924,N_11706);
nor U12445 (N_12445,N_11435,N_11424);
nor U12446 (N_12446,N_11638,N_11521);
and U12447 (N_12447,N_11986,N_11847);
nor U12448 (N_12448,N_11913,N_11659);
and U12449 (N_12449,N_11874,N_11938);
nor U12450 (N_12450,N_11928,N_11548);
nand U12451 (N_12451,N_11516,N_11926);
nor U12452 (N_12452,N_11962,N_11597);
xor U12453 (N_12453,N_11567,N_11731);
nor U12454 (N_12454,N_11871,N_11819);
nand U12455 (N_12455,N_11664,N_11900);
nor U12456 (N_12456,N_11572,N_11796);
nand U12457 (N_12457,N_11568,N_11714);
and U12458 (N_12458,N_11685,N_11519);
xnor U12459 (N_12459,N_11864,N_11462);
or U12460 (N_12460,N_11888,N_11566);
nand U12461 (N_12461,N_11478,N_11792);
nand U12462 (N_12462,N_11504,N_11626);
and U12463 (N_12463,N_11655,N_11698);
or U12464 (N_12464,N_11771,N_11595);
or U12465 (N_12465,N_11690,N_11804);
xnor U12466 (N_12466,N_11673,N_11972);
nand U12467 (N_12467,N_11467,N_11427);
nand U12468 (N_12468,N_11980,N_11873);
or U12469 (N_12469,N_11919,N_11796);
or U12470 (N_12470,N_11625,N_11960);
nand U12471 (N_12471,N_11586,N_11560);
or U12472 (N_12472,N_11885,N_11764);
nand U12473 (N_12473,N_11439,N_11492);
nand U12474 (N_12474,N_11527,N_11748);
or U12475 (N_12475,N_11801,N_11959);
or U12476 (N_12476,N_11484,N_11850);
or U12477 (N_12477,N_11865,N_11913);
nand U12478 (N_12478,N_11920,N_11913);
or U12479 (N_12479,N_11462,N_11488);
and U12480 (N_12480,N_11447,N_11638);
nor U12481 (N_12481,N_11685,N_11482);
and U12482 (N_12482,N_11617,N_11621);
or U12483 (N_12483,N_11496,N_11635);
xor U12484 (N_12484,N_11721,N_11565);
nand U12485 (N_12485,N_11508,N_11451);
nand U12486 (N_12486,N_11614,N_11474);
nand U12487 (N_12487,N_11934,N_11475);
or U12488 (N_12488,N_11759,N_11664);
xnor U12489 (N_12489,N_11411,N_11586);
and U12490 (N_12490,N_11406,N_11577);
and U12491 (N_12491,N_11956,N_11532);
xnor U12492 (N_12492,N_11527,N_11644);
and U12493 (N_12493,N_11777,N_11680);
xnor U12494 (N_12494,N_11620,N_11699);
nand U12495 (N_12495,N_11704,N_11443);
xor U12496 (N_12496,N_11444,N_11614);
or U12497 (N_12497,N_11524,N_11650);
or U12498 (N_12498,N_11601,N_11997);
xnor U12499 (N_12499,N_11675,N_11929);
and U12500 (N_12500,N_11774,N_11629);
nand U12501 (N_12501,N_11587,N_11498);
or U12502 (N_12502,N_11504,N_11538);
xnor U12503 (N_12503,N_11911,N_11647);
nor U12504 (N_12504,N_11484,N_11504);
xnor U12505 (N_12505,N_11542,N_11867);
nand U12506 (N_12506,N_11611,N_11817);
xor U12507 (N_12507,N_11760,N_11527);
or U12508 (N_12508,N_11616,N_11400);
and U12509 (N_12509,N_11891,N_11577);
xnor U12510 (N_12510,N_11686,N_11687);
nor U12511 (N_12511,N_11612,N_11446);
nor U12512 (N_12512,N_11452,N_11904);
xor U12513 (N_12513,N_11471,N_11526);
xor U12514 (N_12514,N_11554,N_11838);
xnor U12515 (N_12515,N_11872,N_11699);
nor U12516 (N_12516,N_11579,N_11522);
nand U12517 (N_12517,N_11420,N_11661);
and U12518 (N_12518,N_11579,N_11598);
and U12519 (N_12519,N_11696,N_11540);
nor U12520 (N_12520,N_11535,N_11529);
nand U12521 (N_12521,N_11812,N_11425);
nor U12522 (N_12522,N_11622,N_11487);
or U12523 (N_12523,N_11561,N_11885);
or U12524 (N_12524,N_11628,N_11995);
nand U12525 (N_12525,N_11551,N_11752);
nor U12526 (N_12526,N_11419,N_11960);
or U12527 (N_12527,N_11753,N_11789);
nor U12528 (N_12528,N_11808,N_11824);
and U12529 (N_12529,N_11924,N_11928);
xor U12530 (N_12530,N_11649,N_11893);
nor U12531 (N_12531,N_11896,N_11443);
and U12532 (N_12532,N_11728,N_11869);
nor U12533 (N_12533,N_11578,N_11459);
or U12534 (N_12534,N_11698,N_11948);
nor U12535 (N_12535,N_11748,N_11447);
and U12536 (N_12536,N_11906,N_11884);
or U12537 (N_12537,N_11545,N_11855);
nor U12538 (N_12538,N_11433,N_11479);
or U12539 (N_12539,N_11814,N_11687);
nand U12540 (N_12540,N_11929,N_11919);
or U12541 (N_12541,N_11926,N_11960);
nand U12542 (N_12542,N_11426,N_11787);
and U12543 (N_12543,N_11570,N_11461);
nor U12544 (N_12544,N_11436,N_11607);
nor U12545 (N_12545,N_11851,N_11419);
nand U12546 (N_12546,N_11404,N_11723);
nor U12547 (N_12547,N_11630,N_11713);
nand U12548 (N_12548,N_11683,N_11893);
and U12549 (N_12549,N_11760,N_11967);
nand U12550 (N_12550,N_11712,N_11466);
and U12551 (N_12551,N_11522,N_11685);
or U12552 (N_12552,N_11782,N_11427);
nand U12553 (N_12553,N_11695,N_11698);
nor U12554 (N_12554,N_11881,N_11750);
or U12555 (N_12555,N_11500,N_11701);
xnor U12556 (N_12556,N_11442,N_11999);
or U12557 (N_12557,N_11573,N_11817);
and U12558 (N_12558,N_11480,N_11845);
or U12559 (N_12559,N_11540,N_11607);
nand U12560 (N_12560,N_11780,N_11746);
and U12561 (N_12561,N_11708,N_11507);
and U12562 (N_12562,N_11747,N_11585);
nor U12563 (N_12563,N_11470,N_11430);
nand U12564 (N_12564,N_11455,N_11888);
or U12565 (N_12565,N_11557,N_11751);
xnor U12566 (N_12566,N_11408,N_11945);
nand U12567 (N_12567,N_11518,N_11423);
nand U12568 (N_12568,N_11961,N_11689);
xnor U12569 (N_12569,N_11753,N_11456);
nor U12570 (N_12570,N_11710,N_11643);
and U12571 (N_12571,N_11533,N_11892);
or U12572 (N_12572,N_11584,N_11599);
xor U12573 (N_12573,N_11694,N_11558);
nor U12574 (N_12574,N_11961,N_11639);
and U12575 (N_12575,N_11826,N_11457);
nand U12576 (N_12576,N_11517,N_11587);
or U12577 (N_12577,N_11918,N_11512);
and U12578 (N_12578,N_11404,N_11973);
or U12579 (N_12579,N_11405,N_11816);
nand U12580 (N_12580,N_11871,N_11707);
or U12581 (N_12581,N_11703,N_11529);
xor U12582 (N_12582,N_11839,N_11778);
xnor U12583 (N_12583,N_11877,N_11508);
or U12584 (N_12584,N_11956,N_11903);
nand U12585 (N_12585,N_11535,N_11892);
nand U12586 (N_12586,N_11490,N_11724);
nand U12587 (N_12587,N_11487,N_11915);
xor U12588 (N_12588,N_11766,N_11507);
nand U12589 (N_12589,N_11541,N_11487);
or U12590 (N_12590,N_11923,N_11837);
nor U12591 (N_12591,N_11637,N_11613);
xor U12592 (N_12592,N_11664,N_11734);
or U12593 (N_12593,N_11743,N_11408);
xnor U12594 (N_12594,N_11917,N_11994);
xnor U12595 (N_12595,N_11427,N_11643);
xnor U12596 (N_12596,N_11629,N_11540);
nor U12597 (N_12597,N_11942,N_11643);
or U12598 (N_12598,N_11751,N_11727);
and U12599 (N_12599,N_11941,N_11787);
xor U12600 (N_12600,N_12480,N_12089);
nor U12601 (N_12601,N_12194,N_12339);
or U12602 (N_12602,N_12126,N_12522);
xor U12603 (N_12603,N_12597,N_12416);
nor U12604 (N_12604,N_12375,N_12579);
nor U12605 (N_12605,N_12091,N_12190);
nor U12606 (N_12606,N_12499,N_12525);
nor U12607 (N_12607,N_12454,N_12340);
nand U12608 (N_12608,N_12311,N_12033);
or U12609 (N_12609,N_12288,N_12181);
nor U12610 (N_12610,N_12401,N_12108);
nand U12611 (N_12611,N_12254,N_12263);
and U12612 (N_12612,N_12364,N_12426);
or U12613 (N_12613,N_12028,N_12558);
nand U12614 (N_12614,N_12225,N_12088);
nor U12615 (N_12615,N_12574,N_12541);
and U12616 (N_12616,N_12468,N_12206);
nand U12617 (N_12617,N_12047,N_12144);
xnor U12618 (N_12618,N_12293,N_12436);
nand U12619 (N_12619,N_12590,N_12071);
and U12620 (N_12620,N_12596,N_12354);
xor U12621 (N_12621,N_12422,N_12081);
nand U12622 (N_12622,N_12456,N_12006);
or U12623 (N_12623,N_12017,N_12378);
and U12624 (N_12624,N_12157,N_12409);
and U12625 (N_12625,N_12418,N_12537);
nand U12626 (N_12626,N_12324,N_12387);
nand U12627 (N_12627,N_12166,N_12437);
nor U12628 (N_12628,N_12245,N_12272);
and U12629 (N_12629,N_12087,N_12327);
xnor U12630 (N_12630,N_12269,N_12459);
and U12631 (N_12631,N_12270,N_12304);
xor U12632 (N_12632,N_12209,N_12345);
nor U12633 (N_12633,N_12106,N_12149);
nand U12634 (N_12634,N_12344,N_12391);
nand U12635 (N_12635,N_12466,N_12580);
nand U12636 (N_12636,N_12576,N_12479);
or U12637 (N_12637,N_12425,N_12407);
xor U12638 (N_12638,N_12388,N_12299);
or U12639 (N_12639,N_12420,N_12187);
xnor U12640 (N_12640,N_12565,N_12271);
xor U12641 (N_12641,N_12408,N_12450);
or U12642 (N_12642,N_12261,N_12275);
nor U12643 (N_12643,N_12498,N_12569);
and U12644 (N_12644,N_12413,N_12204);
or U12645 (N_12645,N_12040,N_12584);
xnor U12646 (N_12646,N_12262,N_12423);
nand U12647 (N_12647,N_12533,N_12158);
nor U12648 (N_12648,N_12515,N_12382);
nor U12649 (N_12649,N_12504,N_12547);
and U12650 (N_12650,N_12022,N_12531);
and U12651 (N_12651,N_12010,N_12491);
nand U12652 (N_12652,N_12084,N_12430);
or U12653 (N_12653,N_12192,N_12027);
nor U12654 (N_12654,N_12312,N_12265);
xnor U12655 (N_12655,N_12247,N_12189);
nand U12656 (N_12656,N_12317,N_12036);
and U12657 (N_12657,N_12101,N_12119);
or U12658 (N_12658,N_12147,N_12449);
nor U12659 (N_12659,N_12346,N_12185);
and U12660 (N_12660,N_12357,N_12500);
xnor U12661 (N_12661,N_12411,N_12148);
or U12662 (N_12662,N_12109,N_12403);
or U12663 (N_12663,N_12062,N_12337);
nand U12664 (N_12664,N_12202,N_12285);
xnor U12665 (N_12665,N_12096,N_12046);
and U12666 (N_12666,N_12308,N_12322);
xor U12667 (N_12667,N_12287,N_12003);
nand U12668 (N_12668,N_12279,N_12412);
xor U12669 (N_12669,N_12004,N_12264);
nand U12670 (N_12670,N_12384,N_12439);
nand U12671 (N_12671,N_12208,N_12267);
and U12672 (N_12672,N_12325,N_12585);
xor U12673 (N_12673,N_12234,N_12593);
xnor U12674 (N_12674,N_12215,N_12122);
xor U12675 (N_12675,N_12059,N_12514);
nand U12676 (N_12676,N_12554,N_12484);
nor U12677 (N_12677,N_12009,N_12309);
and U12678 (N_12678,N_12421,N_12118);
nor U12679 (N_12679,N_12517,N_12107);
nor U12680 (N_12680,N_12534,N_12182);
or U12681 (N_12681,N_12055,N_12079);
nand U12682 (N_12682,N_12080,N_12443);
and U12683 (N_12683,N_12072,N_12550);
xor U12684 (N_12684,N_12535,N_12381);
nand U12685 (N_12685,N_12471,N_12496);
and U12686 (N_12686,N_12336,N_12217);
nand U12687 (N_12687,N_12048,N_12050);
and U12688 (N_12688,N_12394,N_12508);
nand U12689 (N_12689,N_12365,N_12486);
and U12690 (N_12690,N_12174,N_12244);
nor U12691 (N_12691,N_12298,N_12564);
nor U12692 (N_12692,N_12112,N_12528);
and U12693 (N_12693,N_12195,N_12350);
or U12694 (N_12694,N_12183,N_12125);
or U12695 (N_12695,N_12133,N_12044);
xnor U12696 (N_12696,N_12447,N_12197);
or U12697 (N_12697,N_12153,N_12014);
nand U12698 (N_12698,N_12054,N_12130);
and U12699 (N_12699,N_12131,N_12026);
and U12700 (N_12700,N_12025,N_12524);
nor U12701 (N_12701,N_12410,N_12239);
nand U12702 (N_12702,N_12376,N_12518);
nand U12703 (N_12703,N_12061,N_12495);
xor U12704 (N_12704,N_12116,N_12591);
nand U12705 (N_12705,N_12577,N_12374);
nor U12706 (N_12706,N_12427,N_12169);
nor U12707 (N_12707,N_12493,N_12257);
nand U12708 (N_12708,N_12224,N_12451);
nor U12709 (N_12709,N_12458,N_12137);
xnor U12710 (N_12710,N_12582,N_12276);
or U12711 (N_12711,N_12372,N_12064);
and U12712 (N_12712,N_12575,N_12561);
or U12713 (N_12713,N_12552,N_12445);
and U12714 (N_12714,N_12207,N_12502);
and U12715 (N_12715,N_12049,N_12328);
nand U12716 (N_12716,N_12083,N_12452);
nor U12717 (N_12717,N_12599,N_12310);
nand U12718 (N_12718,N_12377,N_12543);
and U12719 (N_12719,N_12492,N_12161);
xor U12720 (N_12720,N_12395,N_12373);
xnor U12721 (N_12721,N_12348,N_12295);
nor U12722 (N_12722,N_12203,N_12219);
or U12723 (N_12723,N_12453,N_12250);
nand U12724 (N_12724,N_12589,N_12464);
nand U12725 (N_12725,N_12164,N_12428);
and U12726 (N_12726,N_12542,N_12505);
or U12727 (N_12727,N_12594,N_12274);
xor U12728 (N_12728,N_12477,N_12159);
nand U12729 (N_12729,N_12513,N_12284);
and U12730 (N_12730,N_12082,N_12196);
nand U12731 (N_12731,N_12058,N_12380);
nor U12732 (N_12732,N_12503,N_12332);
nand U12733 (N_12733,N_12069,N_12165);
nand U12734 (N_12734,N_12231,N_12235);
or U12735 (N_12735,N_12487,N_12463);
nor U12736 (N_12736,N_12007,N_12562);
or U12737 (N_12737,N_12548,N_12056);
or U12738 (N_12738,N_12023,N_12000);
nand U12739 (N_12739,N_12156,N_12019);
nand U12740 (N_12740,N_12201,N_12352);
xnor U12741 (N_12741,N_12123,N_12511);
nor U12742 (N_12742,N_12090,N_12127);
xor U12743 (N_12743,N_12494,N_12462);
nor U12744 (N_12744,N_12470,N_12549);
or U12745 (N_12745,N_12038,N_12353);
or U12746 (N_12746,N_12286,N_12573);
nand U12747 (N_12747,N_12583,N_12297);
or U12748 (N_12748,N_12334,N_12446);
nor U12749 (N_12749,N_12538,N_12240);
nor U12750 (N_12750,N_12570,N_12444);
and U12751 (N_12751,N_12221,N_12251);
nand U12752 (N_12752,N_12306,N_12478);
and U12753 (N_12753,N_12301,N_12140);
and U12754 (N_12754,N_12143,N_12002);
nand U12755 (N_12755,N_12016,N_12232);
nand U12756 (N_12756,N_12103,N_12595);
nor U12757 (N_12757,N_12476,N_12555);
nand U12758 (N_12758,N_12361,N_12406);
and U12759 (N_12759,N_12544,N_12402);
nand U12760 (N_12760,N_12586,N_12483);
and U12761 (N_12761,N_12114,N_12441);
or U12762 (N_12762,N_12553,N_12282);
and U12763 (N_12763,N_12307,N_12199);
nor U12764 (N_12764,N_12005,N_12469);
nand U12765 (N_12765,N_12211,N_12434);
nand U12766 (N_12766,N_12085,N_12472);
xor U12767 (N_12767,N_12008,N_12588);
nand U12768 (N_12768,N_12256,N_12370);
nand U12769 (N_12769,N_12011,N_12142);
and U12770 (N_12770,N_12094,N_12145);
nor U12771 (N_12771,N_12121,N_12146);
xor U12772 (N_12772,N_12236,N_12179);
and U12773 (N_12773,N_12021,N_12516);
nand U12774 (N_12774,N_12155,N_12102);
xnor U12775 (N_12775,N_12135,N_12001);
or U12776 (N_12776,N_12519,N_12120);
xor U12777 (N_12777,N_12520,N_12316);
xor U12778 (N_12778,N_12031,N_12442);
xor U12779 (N_12779,N_12229,N_12419);
xor U12780 (N_12780,N_12020,N_12223);
and U12781 (N_12781,N_12034,N_12172);
or U12782 (N_12782,N_12546,N_12475);
nand U12783 (N_12783,N_12222,N_12030);
and U12784 (N_12784,N_12253,N_12536);
and U12785 (N_12785,N_12457,N_12060);
and U12786 (N_12786,N_12170,N_12053);
xor U12787 (N_12787,N_12323,N_12351);
or U12788 (N_12788,N_12291,N_12198);
or U12789 (N_12789,N_12249,N_12246);
nand U12790 (N_12790,N_12398,N_12512);
xor U12791 (N_12791,N_12448,N_12160);
or U12792 (N_12792,N_12433,N_12393);
nand U12793 (N_12793,N_12294,N_12404);
and U12794 (N_12794,N_12243,N_12313);
or U12795 (N_12795,N_12032,N_12128);
xnor U12796 (N_12796,N_12193,N_12220);
and U12797 (N_12797,N_12063,N_12191);
xor U12798 (N_12798,N_12134,N_12018);
nand U12799 (N_12799,N_12273,N_12474);
and U12800 (N_12800,N_12214,N_12563);
xor U12801 (N_12801,N_12440,N_12024);
nor U12802 (N_12802,N_12051,N_12176);
and U12803 (N_12803,N_12210,N_12216);
nor U12804 (N_12804,N_12093,N_12326);
nor U12805 (N_12805,N_12151,N_12242);
and U12806 (N_12806,N_12556,N_12540);
xor U12807 (N_12807,N_12358,N_12037);
xnor U12808 (N_12808,N_12226,N_12396);
nor U12809 (N_12809,N_12481,N_12111);
nand U12810 (N_12810,N_12200,N_12566);
xor U12811 (N_12811,N_12162,N_12074);
nand U12812 (N_12812,N_12237,N_12526);
nand U12813 (N_12813,N_12057,N_12171);
nor U12814 (N_12814,N_12073,N_12392);
and U12815 (N_12815,N_12539,N_12068);
nor U12816 (N_12816,N_12077,N_12330);
nand U12817 (N_12817,N_12259,N_12067);
or U12818 (N_12818,N_12424,N_12012);
nor U12819 (N_12819,N_12482,N_12414);
xor U12820 (N_12820,N_12296,N_12139);
xnor U12821 (N_12821,N_12371,N_12173);
or U12822 (N_12822,N_12429,N_12136);
nand U12823 (N_12823,N_12355,N_12399);
nand U12824 (N_12824,N_12129,N_12367);
or U12825 (N_12825,N_12241,N_12015);
and U12826 (N_12826,N_12100,N_12314);
xor U12827 (N_12827,N_12186,N_12417);
nor U12828 (N_12828,N_12248,N_12510);
or U12829 (N_12829,N_12485,N_12098);
nor U12830 (N_12830,N_12360,N_12213);
nor U12831 (N_12831,N_12013,N_12435);
or U12832 (N_12832,N_12343,N_12379);
or U12833 (N_12833,N_12230,N_12321);
and U12834 (N_12834,N_12559,N_12238);
xor U12835 (N_12835,N_12557,N_12105);
xnor U12836 (N_12836,N_12052,N_12258);
and U12837 (N_12837,N_12356,N_12507);
nor U12838 (N_12838,N_12347,N_12099);
nor U12839 (N_12839,N_12252,N_12141);
and U12840 (N_12840,N_12587,N_12029);
or U12841 (N_12841,N_12592,N_12042);
and U12842 (N_12842,N_12092,N_12043);
or U12843 (N_12843,N_12397,N_12305);
nor U12844 (N_12844,N_12461,N_12167);
nand U12845 (N_12845,N_12568,N_12473);
nor U12846 (N_12846,N_12152,N_12070);
nand U12847 (N_12847,N_12150,N_12460);
and U12848 (N_12848,N_12154,N_12104);
xnor U12849 (N_12849,N_12302,N_12349);
nor U12850 (N_12850,N_12551,N_12415);
nand U12851 (N_12851,N_12527,N_12389);
nand U12852 (N_12852,N_12228,N_12132);
nand U12853 (N_12853,N_12163,N_12385);
nand U12854 (N_12854,N_12039,N_12455);
and U12855 (N_12855,N_12075,N_12431);
and U12856 (N_12856,N_12233,N_12095);
nor U12857 (N_12857,N_12390,N_12366);
nor U12858 (N_12858,N_12278,N_12205);
xor U12859 (N_12859,N_12280,N_12490);
nor U12860 (N_12860,N_12489,N_12115);
xnor U12861 (N_12861,N_12110,N_12383);
and U12862 (N_12862,N_12260,N_12363);
and U12863 (N_12863,N_12086,N_12041);
or U12864 (N_12864,N_12465,N_12560);
and U12865 (N_12865,N_12318,N_12386);
and U12866 (N_12866,N_12177,N_12368);
xor U12867 (N_12867,N_12212,N_12497);
and U12868 (N_12868,N_12467,N_12117);
nand U12869 (N_12869,N_12078,N_12168);
nor U12870 (N_12870,N_12289,N_12124);
nand U12871 (N_12871,N_12175,N_12506);
nor U12872 (N_12872,N_12331,N_12341);
nand U12873 (N_12873,N_12438,N_12501);
or U12874 (N_12874,N_12342,N_12581);
and U12875 (N_12875,N_12400,N_12076);
or U12876 (N_12876,N_12292,N_12523);
and U12877 (N_12877,N_12578,N_12598);
or U12878 (N_12878,N_12320,N_12530);
xor U12879 (N_12879,N_12359,N_12255);
or U12880 (N_12880,N_12281,N_12283);
xnor U12881 (N_12881,N_12521,N_12571);
and U12882 (N_12882,N_12045,N_12333);
xnor U12883 (N_12883,N_12303,N_12178);
or U12884 (N_12884,N_12138,N_12509);
xnor U12885 (N_12885,N_12315,N_12268);
or U12886 (N_12886,N_12184,N_12290);
or U12887 (N_12887,N_12188,N_12532);
and U12888 (N_12888,N_12227,N_12572);
and U12889 (N_12889,N_12113,N_12300);
nor U12890 (N_12890,N_12035,N_12335);
nor U12891 (N_12891,N_12277,N_12405);
xor U12892 (N_12892,N_12529,N_12319);
or U12893 (N_12893,N_12065,N_12488);
nand U12894 (N_12894,N_12545,N_12180);
nand U12895 (N_12895,N_12266,N_12097);
and U12896 (N_12896,N_12432,N_12338);
or U12897 (N_12897,N_12329,N_12362);
and U12898 (N_12898,N_12369,N_12218);
and U12899 (N_12899,N_12066,N_12567);
and U12900 (N_12900,N_12216,N_12352);
nand U12901 (N_12901,N_12107,N_12071);
or U12902 (N_12902,N_12266,N_12545);
and U12903 (N_12903,N_12429,N_12196);
nor U12904 (N_12904,N_12485,N_12560);
xnor U12905 (N_12905,N_12184,N_12301);
nand U12906 (N_12906,N_12030,N_12376);
nand U12907 (N_12907,N_12410,N_12489);
and U12908 (N_12908,N_12288,N_12282);
nand U12909 (N_12909,N_12076,N_12437);
and U12910 (N_12910,N_12512,N_12149);
xor U12911 (N_12911,N_12472,N_12214);
nand U12912 (N_12912,N_12405,N_12149);
or U12913 (N_12913,N_12404,N_12438);
or U12914 (N_12914,N_12263,N_12043);
and U12915 (N_12915,N_12593,N_12469);
or U12916 (N_12916,N_12228,N_12202);
nor U12917 (N_12917,N_12557,N_12049);
nand U12918 (N_12918,N_12113,N_12384);
and U12919 (N_12919,N_12221,N_12327);
nor U12920 (N_12920,N_12549,N_12060);
nor U12921 (N_12921,N_12382,N_12334);
nor U12922 (N_12922,N_12054,N_12097);
xnor U12923 (N_12923,N_12247,N_12288);
or U12924 (N_12924,N_12187,N_12044);
xnor U12925 (N_12925,N_12205,N_12077);
and U12926 (N_12926,N_12553,N_12514);
or U12927 (N_12927,N_12166,N_12203);
and U12928 (N_12928,N_12261,N_12588);
and U12929 (N_12929,N_12168,N_12430);
nand U12930 (N_12930,N_12406,N_12502);
nand U12931 (N_12931,N_12596,N_12374);
or U12932 (N_12932,N_12537,N_12162);
xor U12933 (N_12933,N_12529,N_12472);
nor U12934 (N_12934,N_12490,N_12419);
xor U12935 (N_12935,N_12264,N_12109);
and U12936 (N_12936,N_12422,N_12192);
or U12937 (N_12937,N_12176,N_12587);
and U12938 (N_12938,N_12545,N_12017);
xnor U12939 (N_12939,N_12550,N_12242);
nand U12940 (N_12940,N_12177,N_12101);
and U12941 (N_12941,N_12096,N_12400);
and U12942 (N_12942,N_12032,N_12224);
or U12943 (N_12943,N_12014,N_12172);
and U12944 (N_12944,N_12399,N_12072);
or U12945 (N_12945,N_12477,N_12272);
or U12946 (N_12946,N_12393,N_12513);
nor U12947 (N_12947,N_12163,N_12508);
or U12948 (N_12948,N_12405,N_12301);
nand U12949 (N_12949,N_12232,N_12083);
nand U12950 (N_12950,N_12252,N_12378);
nand U12951 (N_12951,N_12280,N_12145);
xor U12952 (N_12952,N_12426,N_12261);
xnor U12953 (N_12953,N_12209,N_12024);
nor U12954 (N_12954,N_12464,N_12521);
xor U12955 (N_12955,N_12068,N_12377);
or U12956 (N_12956,N_12379,N_12435);
nand U12957 (N_12957,N_12495,N_12231);
or U12958 (N_12958,N_12063,N_12458);
nor U12959 (N_12959,N_12388,N_12533);
nor U12960 (N_12960,N_12270,N_12318);
and U12961 (N_12961,N_12415,N_12032);
xor U12962 (N_12962,N_12363,N_12257);
or U12963 (N_12963,N_12544,N_12048);
or U12964 (N_12964,N_12285,N_12572);
or U12965 (N_12965,N_12254,N_12180);
xnor U12966 (N_12966,N_12366,N_12010);
and U12967 (N_12967,N_12375,N_12066);
and U12968 (N_12968,N_12403,N_12287);
nor U12969 (N_12969,N_12551,N_12198);
xor U12970 (N_12970,N_12582,N_12205);
xor U12971 (N_12971,N_12554,N_12334);
or U12972 (N_12972,N_12445,N_12273);
nand U12973 (N_12973,N_12348,N_12210);
xnor U12974 (N_12974,N_12398,N_12390);
and U12975 (N_12975,N_12260,N_12494);
or U12976 (N_12976,N_12045,N_12054);
nand U12977 (N_12977,N_12011,N_12201);
xnor U12978 (N_12978,N_12254,N_12289);
and U12979 (N_12979,N_12411,N_12495);
nor U12980 (N_12980,N_12436,N_12526);
or U12981 (N_12981,N_12179,N_12049);
nand U12982 (N_12982,N_12284,N_12188);
and U12983 (N_12983,N_12255,N_12220);
nand U12984 (N_12984,N_12119,N_12417);
and U12985 (N_12985,N_12137,N_12481);
nand U12986 (N_12986,N_12205,N_12170);
xnor U12987 (N_12987,N_12540,N_12072);
nor U12988 (N_12988,N_12293,N_12493);
xor U12989 (N_12989,N_12596,N_12572);
xor U12990 (N_12990,N_12098,N_12160);
and U12991 (N_12991,N_12439,N_12351);
nand U12992 (N_12992,N_12147,N_12235);
nand U12993 (N_12993,N_12312,N_12288);
nand U12994 (N_12994,N_12323,N_12293);
xnor U12995 (N_12995,N_12393,N_12127);
or U12996 (N_12996,N_12484,N_12218);
xor U12997 (N_12997,N_12054,N_12452);
and U12998 (N_12998,N_12246,N_12302);
and U12999 (N_12999,N_12094,N_12168);
nand U13000 (N_13000,N_12556,N_12275);
nand U13001 (N_13001,N_12485,N_12235);
nor U13002 (N_13002,N_12161,N_12489);
or U13003 (N_13003,N_12018,N_12513);
and U13004 (N_13004,N_12143,N_12330);
or U13005 (N_13005,N_12457,N_12099);
or U13006 (N_13006,N_12107,N_12329);
xnor U13007 (N_13007,N_12562,N_12277);
and U13008 (N_13008,N_12410,N_12350);
nor U13009 (N_13009,N_12547,N_12591);
nor U13010 (N_13010,N_12361,N_12130);
or U13011 (N_13011,N_12370,N_12047);
xor U13012 (N_13012,N_12236,N_12162);
nand U13013 (N_13013,N_12574,N_12224);
or U13014 (N_13014,N_12450,N_12059);
xor U13015 (N_13015,N_12328,N_12249);
xnor U13016 (N_13016,N_12280,N_12304);
or U13017 (N_13017,N_12059,N_12035);
nand U13018 (N_13018,N_12133,N_12476);
or U13019 (N_13019,N_12581,N_12228);
or U13020 (N_13020,N_12161,N_12056);
or U13021 (N_13021,N_12244,N_12199);
xor U13022 (N_13022,N_12314,N_12518);
xor U13023 (N_13023,N_12316,N_12466);
or U13024 (N_13024,N_12095,N_12524);
nor U13025 (N_13025,N_12310,N_12345);
nor U13026 (N_13026,N_12283,N_12279);
nor U13027 (N_13027,N_12171,N_12058);
nor U13028 (N_13028,N_12513,N_12519);
xnor U13029 (N_13029,N_12367,N_12192);
nor U13030 (N_13030,N_12354,N_12309);
nor U13031 (N_13031,N_12058,N_12152);
nor U13032 (N_13032,N_12356,N_12302);
and U13033 (N_13033,N_12491,N_12247);
and U13034 (N_13034,N_12349,N_12199);
and U13035 (N_13035,N_12214,N_12456);
nand U13036 (N_13036,N_12015,N_12003);
xnor U13037 (N_13037,N_12316,N_12099);
or U13038 (N_13038,N_12091,N_12537);
nand U13039 (N_13039,N_12359,N_12288);
nand U13040 (N_13040,N_12548,N_12427);
xor U13041 (N_13041,N_12464,N_12152);
nor U13042 (N_13042,N_12547,N_12212);
and U13043 (N_13043,N_12067,N_12077);
xnor U13044 (N_13044,N_12343,N_12151);
and U13045 (N_13045,N_12469,N_12551);
and U13046 (N_13046,N_12335,N_12427);
xor U13047 (N_13047,N_12371,N_12523);
or U13048 (N_13048,N_12162,N_12268);
nand U13049 (N_13049,N_12555,N_12204);
and U13050 (N_13050,N_12427,N_12121);
or U13051 (N_13051,N_12141,N_12452);
xnor U13052 (N_13052,N_12551,N_12101);
nand U13053 (N_13053,N_12037,N_12072);
or U13054 (N_13054,N_12428,N_12396);
or U13055 (N_13055,N_12420,N_12578);
and U13056 (N_13056,N_12051,N_12376);
nor U13057 (N_13057,N_12410,N_12026);
xnor U13058 (N_13058,N_12214,N_12047);
nor U13059 (N_13059,N_12017,N_12226);
or U13060 (N_13060,N_12062,N_12108);
xnor U13061 (N_13061,N_12257,N_12052);
nand U13062 (N_13062,N_12349,N_12487);
xor U13063 (N_13063,N_12346,N_12448);
nand U13064 (N_13064,N_12014,N_12243);
nor U13065 (N_13065,N_12527,N_12348);
xnor U13066 (N_13066,N_12360,N_12284);
nor U13067 (N_13067,N_12331,N_12571);
xor U13068 (N_13068,N_12187,N_12493);
xnor U13069 (N_13069,N_12328,N_12136);
nand U13070 (N_13070,N_12371,N_12441);
xnor U13071 (N_13071,N_12277,N_12449);
or U13072 (N_13072,N_12322,N_12092);
xnor U13073 (N_13073,N_12280,N_12359);
nor U13074 (N_13074,N_12387,N_12074);
nor U13075 (N_13075,N_12304,N_12511);
nor U13076 (N_13076,N_12385,N_12454);
or U13077 (N_13077,N_12315,N_12205);
nand U13078 (N_13078,N_12558,N_12465);
nor U13079 (N_13079,N_12018,N_12173);
and U13080 (N_13080,N_12555,N_12446);
or U13081 (N_13081,N_12070,N_12229);
and U13082 (N_13082,N_12030,N_12112);
and U13083 (N_13083,N_12379,N_12118);
and U13084 (N_13084,N_12242,N_12387);
and U13085 (N_13085,N_12030,N_12484);
xnor U13086 (N_13086,N_12198,N_12146);
nor U13087 (N_13087,N_12343,N_12022);
nor U13088 (N_13088,N_12309,N_12327);
and U13089 (N_13089,N_12531,N_12529);
nor U13090 (N_13090,N_12252,N_12067);
nor U13091 (N_13091,N_12497,N_12575);
nor U13092 (N_13092,N_12316,N_12421);
nor U13093 (N_13093,N_12161,N_12138);
or U13094 (N_13094,N_12595,N_12296);
nand U13095 (N_13095,N_12456,N_12539);
or U13096 (N_13096,N_12347,N_12231);
nand U13097 (N_13097,N_12518,N_12386);
xnor U13098 (N_13098,N_12252,N_12383);
and U13099 (N_13099,N_12389,N_12555);
or U13100 (N_13100,N_12266,N_12140);
xor U13101 (N_13101,N_12294,N_12365);
nand U13102 (N_13102,N_12444,N_12490);
or U13103 (N_13103,N_12316,N_12394);
nand U13104 (N_13104,N_12323,N_12388);
nor U13105 (N_13105,N_12159,N_12037);
or U13106 (N_13106,N_12153,N_12010);
xor U13107 (N_13107,N_12272,N_12531);
nand U13108 (N_13108,N_12277,N_12430);
nor U13109 (N_13109,N_12424,N_12097);
and U13110 (N_13110,N_12283,N_12268);
nand U13111 (N_13111,N_12219,N_12037);
nor U13112 (N_13112,N_12361,N_12103);
and U13113 (N_13113,N_12459,N_12224);
nor U13114 (N_13114,N_12039,N_12154);
and U13115 (N_13115,N_12249,N_12345);
nand U13116 (N_13116,N_12500,N_12125);
nor U13117 (N_13117,N_12479,N_12227);
nand U13118 (N_13118,N_12158,N_12292);
xnor U13119 (N_13119,N_12114,N_12556);
xor U13120 (N_13120,N_12457,N_12070);
nor U13121 (N_13121,N_12161,N_12262);
or U13122 (N_13122,N_12258,N_12518);
nor U13123 (N_13123,N_12124,N_12078);
or U13124 (N_13124,N_12273,N_12230);
nand U13125 (N_13125,N_12150,N_12064);
xnor U13126 (N_13126,N_12079,N_12584);
nor U13127 (N_13127,N_12445,N_12014);
nor U13128 (N_13128,N_12284,N_12383);
or U13129 (N_13129,N_12318,N_12484);
nor U13130 (N_13130,N_12120,N_12442);
or U13131 (N_13131,N_12491,N_12023);
and U13132 (N_13132,N_12279,N_12323);
nand U13133 (N_13133,N_12456,N_12046);
nor U13134 (N_13134,N_12081,N_12569);
or U13135 (N_13135,N_12048,N_12453);
nor U13136 (N_13136,N_12282,N_12574);
nor U13137 (N_13137,N_12165,N_12273);
or U13138 (N_13138,N_12208,N_12570);
and U13139 (N_13139,N_12224,N_12158);
or U13140 (N_13140,N_12304,N_12053);
xor U13141 (N_13141,N_12378,N_12087);
xor U13142 (N_13142,N_12248,N_12538);
nand U13143 (N_13143,N_12180,N_12011);
or U13144 (N_13144,N_12064,N_12138);
xor U13145 (N_13145,N_12486,N_12269);
nor U13146 (N_13146,N_12115,N_12351);
and U13147 (N_13147,N_12425,N_12540);
xor U13148 (N_13148,N_12050,N_12098);
xor U13149 (N_13149,N_12501,N_12001);
or U13150 (N_13150,N_12182,N_12593);
nand U13151 (N_13151,N_12096,N_12071);
and U13152 (N_13152,N_12072,N_12520);
nor U13153 (N_13153,N_12228,N_12356);
and U13154 (N_13154,N_12280,N_12484);
and U13155 (N_13155,N_12084,N_12305);
xor U13156 (N_13156,N_12227,N_12355);
nand U13157 (N_13157,N_12541,N_12305);
nor U13158 (N_13158,N_12183,N_12034);
xor U13159 (N_13159,N_12169,N_12537);
nor U13160 (N_13160,N_12352,N_12168);
nor U13161 (N_13161,N_12352,N_12022);
or U13162 (N_13162,N_12386,N_12316);
xor U13163 (N_13163,N_12520,N_12508);
nor U13164 (N_13164,N_12594,N_12042);
and U13165 (N_13165,N_12094,N_12562);
or U13166 (N_13166,N_12244,N_12218);
or U13167 (N_13167,N_12020,N_12131);
nor U13168 (N_13168,N_12259,N_12556);
or U13169 (N_13169,N_12382,N_12518);
or U13170 (N_13170,N_12472,N_12255);
or U13171 (N_13171,N_12515,N_12595);
xnor U13172 (N_13172,N_12221,N_12574);
xor U13173 (N_13173,N_12546,N_12318);
and U13174 (N_13174,N_12355,N_12530);
and U13175 (N_13175,N_12258,N_12118);
nand U13176 (N_13176,N_12305,N_12144);
and U13177 (N_13177,N_12305,N_12228);
nor U13178 (N_13178,N_12077,N_12043);
nand U13179 (N_13179,N_12090,N_12101);
xnor U13180 (N_13180,N_12218,N_12537);
xor U13181 (N_13181,N_12088,N_12107);
nor U13182 (N_13182,N_12344,N_12093);
and U13183 (N_13183,N_12138,N_12154);
nand U13184 (N_13184,N_12111,N_12511);
or U13185 (N_13185,N_12243,N_12082);
xnor U13186 (N_13186,N_12034,N_12245);
xnor U13187 (N_13187,N_12280,N_12059);
and U13188 (N_13188,N_12179,N_12590);
xnor U13189 (N_13189,N_12000,N_12510);
or U13190 (N_13190,N_12165,N_12558);
or U13191 (N_13191,N_12582,N_12033);
and U13192 (N_13192,N_12229,N_12039);
and U13193 (N_13193,N_12580,N_12351);
or U13194 (N_13194,N_12562,N_12021);
nand U13195 (N_13195,N_12567,N_12309);
xnor U13196 (N_13196,N_12317,N_12587);
or U13197 (N_13197,N_12568,N_12341);
xor U13198 (N_13198,N_12171,N_12427);
and U13199 (N_13199,N_12186,N_12526);
or U13200 (N_13200,N_12763,N_13199);
nor U13201 (N_13201,N_12712,N_13037);
nand U13202 (N_13202,N_13141,N_13167);
nor U13203 (N_13203,N_13135,N_12833);
nand U13204 (N_13204,N_12629,N_13017);
and U13205 (N_13205,N_13022,N_12824);
and U13206 (N_13206,N_13002,N_13095);
or U13207 (N_13207,N_12776,N_12917);
or U13208 (N_13208,N_12849,N_13129);
or U13209 (N_13209,N_12721,N_12768);
nand U13210 (N_13210,N_13125,N_12656);
nor U13211 (N_13211,N_12739,N_13179);
and U13212 (N_13212,N_12627,N_13015);
or U13213 (N_13213,N_13120,N_13164);
or U13214 (N_13214,N_12910,N_13050);
or U13215 (N_13215,N_13126,N_13006);
xnor U13216 (N_13216,N_12643,N_12935);
xnor U13217 (N_13217,N_12693,N_12808);
or U13218 (N_13218,N_13137,N_13084);
xor U13219 (N_13219,N_12899,N_13012);
xor U13220 (N_13220,N_12773,N_13074);
xnor U13221 (N_13221,N_12796,N_12619);
nand U13222 (N_13222,N_12982,N_13131);
nand U13223 (N_13223,N_12992,N_12651);
nand U13224 (N_13224,N_13091,N_13182);
nor U13225 (N_13225,N_12702,N_12886);
nor U13226 (N_13226,N_12701,N_12969);
nand U13227 (N_13227,N_13175,N_12984);
and U13228 (N_13228,N_12914,N_13109);
nor U13229 (N_13229,N_12714,N_13134);
xnor U13230 (N_13230,N_12756,N_13078);
or U13231 (N_13231,N_12749,N_13088);
nand U13232 (N_13232,N_13083,N_12754);
nand U13233 (N_13233,N_12665,N_12755);
and U13234 (N_13234,N_12863,N_13154);
or U13235 (N_13235,N_13021,N_12858);
nor U13236 (N_13236,N_13193,N_13171);
or U13237 (N_13237,N_12669,N_12658);
nand U13238 (N_13238,N_12900,N_13068);
and U13239 (N_13239,N_12645,N_13052);
and U13240 (N_13240,N_12868,N_13044);
or U13241 (N_13241,N_12678,N_12624);
nor U13242 (N_13242,N_12946,N_12743);
nand U13243 (N_13243,N_12828,N_12662);
nor U13244 (N_13244,N_12862,N_12971);
nand U13245 (N_13245,N_13176,N_13198);
nor U13246 (N_13246,N_13183,N_12847);
and U13247 (N_13247,N_13145,N_12852);
nand U13248 (N_13248,N_12797,N_13048);
nor U13249 (N_13249,N_12883,N_12894);
and U13250 (N_13250,N_12961,N_13077);
and U13251 (N_13251,N_12944,N_12879);
nand U13252 (N_13252,N_12681,N_13026);
xor U13253 (N_13253,N_12890,N_13032);
or U13254 (N_13254,N_12696,N_12860);
nand U13255 (N_13255,N_12607,N_13113);
nand U13256 (N_13256,N_12973,N_12933);
nand U13257 (N_13257,N_12759,N_13055);
and U13258 (N_13258,N_12830,N_12789);
or U13259 (N_13259,N_12994,N_13073);
xnor U13260 (N_13260,N_13102,N_13023);
xor U13261 (N_13261,N_13180,N_12941);
nand U13262 (N_13262,N_12908,N_12778);
nand U13263 (N_13263,N_13003,N_12794);
nand U13264 (N_13264,N_13070,N_13172);
or U13265 (N_13265,N_13019,N_12955);
xnor U13266 (N_13266,N_13028,N_12659);
and U13267 (N_13267,N_12741,N_13049);
xor U13268 (N_13268,N_12764,N_12762);
and U13269 (N_13269,N_12806,N_13186);
nand U13270 (N_13270,N_13143,N_12803);
and U13271 (N_13271,N_13057,N_12939);
and U13272 (N_13272,N_13065,N_12731);
nor U13273 (N_13273,N_12630,N_13136);
and U13274 (N_13274,N_12734,N_12835);
xor U13275 (N_13275,N_12765,N_12811);
nand U13276 (N_13276,N_12725,N_12807);
xnor U13277 (N_13277,N_12628,N_13067);
xor U13278 (N_13278,N_13115,N_13086);
xor U13279 (N_13279,N_12817,N_12742);
nand U13280 (N_13280,N_12909,N_12747);
nand U13281 (N_13281,N_12716,N_12892);
and U13282 (N_13282,N_12898,N_13170);
nor U13283 (N_13283,N_13051,N_12885);
xor U13284 (N_13284,N_12815,N_13060);
nand U13285 (N_13285,N_12934,N_12613);
or U13286 (N_13286,N_13165,N_12928);
nand U13287 (N_13287,N_12987,N_12788);
xnor U13288 (N_13288,N_13150,N_13197);
xnor U13289 (N_13289,N_13079,N_12729);
nand U13290 (N_13290,N_12623,N_13168);
nor U13291 (N_13291,N_12834,N_12612);
or U13292 (N_13292,N_12728,N_13064);
xnor U13293 (N_13293,N_13119,N_13054);
xnor U13294 (N_13294,N_13082,N_12960);
and U13295 (N_13295,N_13033,N_12634);
or U13296 (N_13296,N_12947,N_12615);
nor U13297 (N_13297,N_12821,N_12942);
and U13298 (N_13298,N_13185,N_13100);
and U13299 (N_13299,N_12737,N_12748);
or U13300 (N_13300,N_12979,N_13076);
xnor U13301 (N_13301,N_12915,N_12779);
and U13302 (N_13302,N_13038,N_12666);
or U13303 (N_13303,N_12838,N_13138);
xnor U13304 (N_13304,N_13024,N_12745);
and U13305 (N_13305,N_12903,N_13005);
and U13306 (N_13306,N_12770,N_13035);
xnor U13307 (N_13307,N_12924,N_12854);
or U13308 (N_13308,N_12679,N_12641);
and U13309 (N_13309,N_13056,N_12784);
xnor U13310 (N_13310,N_12866,N_12724);
and U13311 (N_13311,N_12953,N_13151);
nand U13312 (N_13312,N_13045,N_12839);
or U13313 (N_13313,N_12962,N_12932);
xnor U13314 (N_13314,N_12600,N_13173);
nor U13315 (N_13315,N_13063,N_12649);
nand U13316 (N_13316,N_13146,N_13071);
and U13317 (N_13317,N_13001,N_12667);
and U13318 (N_13318,N_12676,N_12823);
nand U13319 (N_13319,N_12775,N_12790);
nand U13320 (N_13320,N_13130,N_12875);
nor U13321 (N_13321,N_12949,N_12738);
or U13322 (N_13322,N_12638,N_12786);
or U13323 (N_13323,N_12608,N_13110);
or U13324 (N_13324,N_12733,N_12744);
xnor U13325 (N_13325,N_12672,N_12753);
nand U13326 (N_13326,N_13192,N_13112);
and U13327 (N_13327,N_12675,N_12884);
xor U13328 (N_13328,N_12995,N_12606);
or U13329 (N_13329,N_12648,N_12818);
nand U13330 (N_13330,N_12795,N_13177);
nor U13331 (N_13331,N_12804,N_12881);
and U13332 (N_13332,N_12976,N_12967);
xor U13333 (N_13333,N_12893,N_12660);
or U13334 (N_13334,N_13020,N_13148);
nor U13335 (N_13335,N_12895,N_12652);
nor U13336 (N_13336,N_13030,N_12611);
and U13337 (N_13337,N_12950,N_13059);
nor U13338 (N_13338,N_12988,N_13178);
or U13339 (N_13339,N_12640,N_12601);
or U13340 (N_13340,N_13142,N_12926);
nor U13341 (N_13341,N_12814,N_12736);
or U13342 (N_13342,N_13097,N_12952);
or U13343 (N_13343,N_12816,N_13027);
or U13344 (N_13344,N_12896,N_12889);
nor U13345 (N_13345,N_12869,N_12902);
nor U13346 (N_13346,N_12717,N_12735);
or U13347 (N_13347,N_12713,N_12867);
nand U13348 (N_13348,N_12945,N_12621);
and U13349 (N_13349,N_13162,N_13195);
xnor U13350 (N_13350,N_13155,N_12777);
xor U13351 (N_13351,N_12657,N_13156);
and U13352 (N_13352,N_12810,N_13029);
xor U13353 (N_13353,N_13163,N_12752);
or U13354 (N_13354,N_13013,N_12906);
and U13355 (N_13355,N_12874,N_12951);
nand U13356 (N_13356,N_13169,N_13075);
nor U13357 (N_13357,N_12771,N_12691);
or U13358 (N_13358,N_13159,N_12793);
or U13359 (N_13359,N_12997,N_12699);
or U13360 (N_13360,N_12975,N_12663);
nand U13361 (N_13361,N_13016,N_12963);
and U13362 (N_13362,N_12977,N_13144);
or U13363 (N_13363,N_12706,N_13041);
and U13364 (N_13364,N_12792,N_12689);
nand U13365 (N_13365,N_12620,N_12943);
nor U13366 (N_13366,N_12826,N_13161);
and U13367 (N_13367,N_12639,N_13108);
and U13368 (N_13368,N_12974,N_12825);
nor U13369 (N_13369,N_12837,N_12798);
xor U13370 (N_13370,N_13105,N_13094);
and U13371 (N_13371,N_13062,N_12980);
or U13372 (N_13372,N_12888,N_13018);
nor U13373 (N_13373,N_13128,N_13087);
nor U13374 (N_13374,N_12829,N_12887);
and U13375 (N_13375,N_12602,N_12938);
and U13376 (N_13376,N_13009,N_13031);
and U13377 (N_13377,N_12993,N_12664);
or U13378 (N_13378,N_13188,N_12880);
nand U13379 (N_13379,N_13114,N_13010);
or U13380 (N_13380,N_12948,N_13149);
xnor U13381 (N_13381,N_12625,N_12840);
nand U13382 (N_13382,N_12637,N_12685);
nor U13383 (N_13383,N_12654,N_12855);
nor U13384 (N_13384,N_13085,N_13196);
xnor U13385 (N_13385,N_13080,N_12646);
nand U13386 (N_13386,N_13117,N_12616);
xor U13387 (N_13387,N_12700,N_12872);
xor U13388 (N_13388,N_12781,N_12760);
or U13389 (N_13389,N_13184,N_12626);
and U13390 (N_13390,N_12709,N_12986);
xor U13391 (N_13391,N_12972,N_12710);
nor U13392 (N_13392,N_13043,N_13174);
xnor U13393 (N_13393,N_13123,N_13111);
nor U13394 (N_13394,N_12920,N_12750);
nand U13395 (N_13395,N_12769,N_12871);
nand U13396 (N_13396,N_13157,N_12851);
nand U13397 (N_13397,N_12965,N_13092);
nor U13398 (N_13398,N_13190,N_12916);
nor U13399 (N_13399,N_12703,N_13191);
and U13400 (N_13400,N_12930,N_12682);
nor U13401 (N_13401,N_13158,N_12897);
and U13402 (N_13402,N_12846,N_12730);
nor U13403 (N_13403,N_13122,N_13121);
or U13404 (N_13404,N_12726,N_12878);
and U13405 (N_13405,N_12956,N_13046);
xor U13406 (N_13406,N_12873,N_13061);
or U13407 (N_13407,N_13132,N_12761);
nor U13408 (N_13408,N_13099,N_12882);
or U13409 (N_13409,N_12891,N_12683);
nor U13410 (N_13410,N_12800,N_12694);
xor U13411 (N_13411,N_12985,N_12931);
or U13412 (N_13412,N_12998,N_12991);
nand U13413 (N_13413,N_12785,N_12644);
nand U13414 (N_13414,N_12813,N_13053);
nand U13415 (N_13415,N_13004,N_12958);
and U13416 (N_13416,N_12751,N_12705);
nand U13417 (N_13417,N_12850,N_12957);
nand U13418 (N_13418,N_12604,N_12999);
or U13419 (N_13419,N_12836,N_12697);
nor U13420 (N_13420,N_12632,N_12722);
xor U13421 (N_13421,N_12708,N_12901);
nand U13422 (N_13422,N_12844,N_12853);
nand U13423 (N_13423,N_13040,N_12704);
nor U13424 (N_13424,N_12925,N_12772);
xnor U13425 (N_13425,N_12820,N_12688);
nor U13426 (N_13426,N_12653,N_12633);
xor U13427 (N_13427,N_13039,N_12695);
or U13428 (N_13428,N_13007,N_13011);
nor U13429 (N_13429,N_12981,N_12978);
xnor U13430 (N_13430,N_12740,N_12996);
xor U13431 (N_13431,N_12715,N_13090);
nor U13432 (N_13432,N_12922,N_12848);
xnor U13433 (N_13433,N_13034,N_12780);
xor U13434 (N_13434,N_12959,N_13036);
or U13435 (N_13435,N_12650,N_12610);
xnor U13436 (N_13436,N_13160,N_13098);
xor U13437 (N_13437,N_12918,N_12617);
nand U13438 (N_13438,N_12783,N_12870);
nand U13439 (N_13439,N_12727,N_12671);
nor U13440 (N_13440,N_12684,N_12711);
or U13441 (N_13441,N_12905,N_12904);
xnor U13442 (N_13442,N_12841,N_13042);
xnor U13443 (N_13443,N_12827,N_12865);
and U13444 (N_13444,N_12668,N_13058);
nand U13445 (N_13445,N_12655,N_12907);
nor U13446 (N_13446,N_13116,N_13093);
nor U13447 (N_13447,N_12647,N_12774);
and U13448 (N_13448,N_13118,N_12642);
nand U13449 (N_13449,N_12842,N_12856);
xor U13450 (N_13450,N_13124,N_12990);
and U13451 (N_13451,N_13025,N_12674);
or U13452 (N_13452,N_12609,N_13014);
nor U13453 (N_13453,N_13127,N_12636);
nor U13454 (N_13454,N_12677,N_12661);
or U13455 (N_13455,N_12845,N_12966);
xnor U13456 (N_13456,N_12603,N_12723);
xor U13457 (N_13457,N_12912,N_12970);
and U13458 (N_13458,N_12831,N_12767);
xor U13459 (N_13459,N_12968,N_13069);
and U13460 (N_13460,N_12859,N_13103);
nor U13461 (N_13461,N_12673,N_12635);
or U13462 (N_13462,N_12936,N_12718);
xnor U13463 (N_13463,N_12954,N_13152);
xor U13464 (N_13464,N_13081,N_12787);
xnor U13465 (N_13465,N_12937,N_13066);
and U13466 (N_13466,N_12799,N_12631);
nor U13467 (N_13467,N_12927,N_12670);
nor U13468 (N_13468,N_13106,N_13153);
or U13469 (N_13469,N_12812,N_12698);
nand U13470 (N_13470,N_12843,N_13140);
or U13471 (N_13471,N_12614,N_12618);
nand U13472 (N_13472,N_12921,N_12832);
or U13473 (N_13473,N_12746,N_12940);
nand U13474 (N_13474,N_12923,N_13072);
and U13475 (N_13475,N_12719,N_12876);
xor U13476 (N_13476,N_12864,N_13187);
xnor U13477 (N_13477,N_12707,N_12732);
and U13478 (N_13478,N_12622,N_13181);
or U13479 (N_13479,N_12692,N_13096);
and U13480 (N_13480,N_12802,N_13133);
nor U13481 (N_13481,N_13194,N_13189);
nand U13482 (N_13482,N_13089,N_12782);
nor U13483 (N_13483,N_12680,N_13008);
nand U13484 (N_13484,N_13101,N_13104);
and U13485 (N_13485,N_12822,N_12766);
xnor U13486 (N_13486,N_12757,N_12913);
or U13487 (N_13487,N_12805,N_12819);
and U13488 (N_13488,N_13139,N_12605);
and U13489 (N_13489,N_12791,N_12687);
nand U13490 (N_13490,N_13107,N_12989);
xor U13491 (N_13491,N_12929,N_12911);
xor U13492 (N_13492,N_12801,N_12861);
nor U13493 (N_13493,N_12877,N_12809);
nor U13494 (N_13494,N_12758,N_12983);
xor U13495 (N_13495,N_13147,N_12857);
and U13496 (N_13496,N_13000,N_12919);
and U13497 (N_13497,N_12720,N_13166);
and U13498 (N_13498,N_12964,N_12690);
or U13499 (N_13499,N_13047,N_12686);
nor U13500 (N_13500,N_12685,N_13122);
or U13501 (N_13501,N_13164,N_12943);
xnor U13502 (N_13502,N_12949,N_12618);
nand U13503 (N_13503,N_13093,N_12640);
nor U13504 (N_13504,N_12952,N_12817);
and U13505 (N_13505,N_12681,N_12667);
nor U13506 (N_13506,N_12719,N_12606);
and U13507 (N_13507,N_13175,N_13084);
and U13508 (N_13508,N_12954,N_12958);
nor U13509 (N_13509,N_12607,N_12761);
nor U13510 (N_13510,N_12762,N_13192);
or U13511 (N_13511,N_12783,N_13083);
nand U13512 (N_13512,N_12844,N_12799);
and U13513 (N_13513,N_12818,N_12807);
and U13514 (N_13514,N_13003,N_12679);
nand U13515 (N_13515,N_13094,N_12621);
nand U13516 (N_13516,N_13147,N_12606);
nand U13517 (N_13517,N_13124,N_13195);
nand U13518 (N_13518,N_12623,N_12695);
and U13519 (N_13519,N_12642,N_12670);
xnor U13520 (N_13520,N_12625,N_12933);
or U13521 (N_13521,N_13057,N_12607);
nor U13522 (N_13522,N_12910,N_12759);
nor U13523 (N_13523,N_13081,N_13184);
and U13524 (N_13524,N_12667,N_12998);
xor U13525 (N_13525,N_12788,N_12719);
nor U13526 (N_13526,N_12769,N_12921);
nor U13527 (N_13527,N_12632,N_12855);
or U13528 (N_13528,N_13006,N_13029);
or U13529 (N_13529,N_12948,N_12700);
or U13530 (N_13530,N_12796,N_13081);
xor U13531 (N_13531,N_13143,N_12703);
or U13532 (N_13532,N_13120,N_12666);
xnor U13533 (N_13533,N_12785,N_13167);
xor U13534 (N_13534,N_13137,N_13067);
and U13535 (N_13535,N_13059,N_12738);
xor U13536 (N_13536,N_12881,N_13197);
nand U13537 (N_13537,N_12832,N_12890);
and U13538 (N_13538,N_12806,N_13061);
and U13539 (N_13539,N_12670,N_12730);
nor U13540 (N_13540,N_12885,N_12700);
xor U13541 (N_13541,N_12951,N_13179);
nand U13542 (N_13542,N_13180,N_12919);
and U13543 (N_13543,N_13110,N_13048);
and U13544 (N_13544,N_12703,N_12966);
and U13545 (N_13545,N_12826,N_12796);
and U13546 (N_13546,N_12666,N_12672);
or U13547 (N_13547,N_12905,N_13122);
and U13548 (N_13548,N_13047,N_12988);
or U13549 (N_13549,N_12894,N_13049);
nor U13550 (N_13550,N_12782,N_12634);
nor U13551 (N_13551,N_12906,N_12733);
or U13552 (N_13552,N_12979,N_13161);
nor U13553 (N_13553,N_12635,N_12949);
xor U13554 (N_13554,N_12661,N_12999);
nor U13555 (N_13555,N_13066,N_12917);
nor U13556 (N_13556,N_12808,N_13180);
xnor U13557 (N_13557,N_13112,N_12830);
nand U13558 (N_13558,N_13103,N_13042);
and U13559 (N_13559,N_12795,N_12873);
xor U13560 (N_13560,N_12787,N_12650);
xor U13561 (N_13561,N_12885,N_13164);
xor U13562 (N_13562,N_13169,N_13182);
nor U13563 (N_13563,N_12654,N_12666);
nor U13564 (N_13564,N_13110,N_13187);
or U13565 (N_13565,N_13134,N_12994);
nand U13566 (N_13566,N_13100,N_12618);
xor U13567 (N_13567,N_12650,N_13009);
nor U13568 (N_13568,N_12969,N_12805);
or U13569 (N_13569,N_13061,N_13169);
xnor U13570 (N_13570,N_12864,N_13029);
and U13571 (N_13571,N_12878,N_12923);
xor U13572 (N_13572,N_12692,N_12696);
and U13573 (N_13573,N_12766,N_12907);
nor U13574 (N_13574,N_12753,N_13070);
xor U13575 (N_13575,N_13000,N_13150);
nor U13576 (N_13576,N_12802,N_12619);
nor U13577 (N_13577,N_12914,N_12975);
nor U13578 (N_13578,N_13100,N_12910);
nor U13579 (N_13579,N_12741,N_12939);
or U13580 (N_13580,N_12730,N_12739);
nand U13581 (N_13581,N_12912,N_12924);
nand U13582 (N_13582,N_13143,N_12682);
or U13583 (N_13583,N_12620,N_12926);
xnor U13584 (N_13584,N_13140,N_12665);
nand U13585 (N_13585,N_12645,N_13092);
or U13586 (N_13586,N_12711,N_12804);
nand U13587 (N_13587,N_12889,N_12847);
or U13588 (N_13588,N_12885,N_12842);
nor U13589 (N_13589,N_12843,N_12835);
xnor U13590 (N_13590,N_12840,N_13012);
and U13591 (N_13591,N_12600,N_13089);
nand U13592 (N_13592,N_12960,N_13010);
and U13593 (N_13593,N_12901,N_12604);
nor U13594 (N_13594,N_13186,N_13143);
nand U13595 (N_13595,N_12711,N_13122);
nor U13596 (N_13596,N_13129,N_12801);
nand U13597 (N_13597,N_13002,N_12688);
xor U13598 (N_13598,N_13106,N_12816);
xor U13599 (N_13599,N_12659,N_13174);
and U13600 (N_13600,N_12883,N_13078);
or U13601 (N_13601,N_12620,N_12744);
and U13602 (N_13602,N_13089,N_12820);
nand U13603 (N_13603,N_12765,N_12826);
or U13604 (N_13604,N_13141,N_12673);
nand U13605 (N_13605,N_12867,N_12964);
or U13606 (N_13606,N_12635,N_12907);
nor U13607 (N_13607,N_12755,N_12865);
xor U13608 (N_13608,N_12908,N_12947);
nand U13609 (N_13609,N_12704,N_12729);
nand U13610 (N_13610,N_12748,N_13113);
and U13611 (N_13611,N_13036,N_12702);
xor U13612 (N_13612,N_13129,N_13023);
or U13613 (N_13613,N_12958,N_12979);
nand U13614 (N_13614,N_13186,N_13137);
or U13615 (N_13615,N_13128,N_12893);
nand U13616 (N_13616,N_12879,N_13057);
nor U13617 (N_13617,N_12613,N_13193);
nand U13618 (N_13618,N_13110,N_12822);
and U13619 (N_13619,N_13117,N_13081);
xor U13620 (N_13620,N_12717,N_12894);
or U13621 (N_13621,N_12704,N_12895);
or U13622 (N_13622,N_12670,N_12717);
xnor U13623 (N_13623,N_12707,N_13193);
xnor U13624 (N_13624,N_13068,N_13172);
nand U13625 (N_13625,N_13004,N_13071);
nand U13626 (N_13626,N_12708,N_12819);
xnor U13627 (N_13627,N_13177,N_12966);
or U13628 (N_13628,N_12844,N_12819);
nand U13629 (N_13629,N_12699,N_13008);
nand U13630 (N_13630,N_12962,N_12809);
xor U13631 (N_13631,N_12648,N_12778);
nor U13632 (N_13632,N_12882,N_13182);
or U13633 (N_13633,N_13168,N_12973);
or U13634 (N_13634,N_13031,N_13115);
nand U13635 (N_13635,N_12657,N_13130);
and U13636 (N_13636,N_13114,N_13122);
nand U13637 (N_13637,N_12858,N_12699);
and U13638 (N_13638,N_12888,N_13146);
xnor U13639 (N_13639,N_12746,N_12603);
xor U13640 (N_13640,N_13098,N_12681);
xnor U13641 (N_13641,N_12698,N_13039);
or U13642 (N_13642,N_12793,N_12616);
nor U13643 (N_13643,N_12951,N_12890);
xnor U13644 (N_13644,N_12746,N_12727);
nand U13645 (N_13645,N_12882,N_13094);
and U13646 (N_13646,N_12989,N_12739);
nor U13647 (N_13647,N_12704,N_13091);
and U13648 (N_13648,N_12973,N_12741);
nor U13649 (N_13649,N_13092,N_12708);
or U13650 (N_13650,N_12656,N_12651);
nor U13651 (N_13651,N_12749,N_12890);
or U13652 (N_13652,N_13141,N_12867);
nand U13653 (N_13653,N_12888,N_13060);
nand U13654 (N_13654,N_12621,N_12618);
nand U13655 (N_13655,N_13071,N_12970);
nor U13656 (N_13656,N_12683,N_13094);
nand U13657 (N_13657,N_13092,N_12884);
xnor U13658 (N_13658,N_12625,N_12972);
or U13659 (N_13659,N_12711,N_12634);
or U13660 (N_13660,N_12615,N_13043);
nor U13661 (N_13661,N_13030,N_12972);
or U13662 (N_13662,N_12883,N_13194);
or U13663 (N_13663,N_13066,N_12682);
xnor U13664 (N_13664,N_12759,N_12896);
and U13665 (N_13665,N_13158,N_13021);
and U13666 (N_13666,N_12952,N_13042);
nand U13667 (N_13667,N_12658,N_12646);
or U13668 (N_13668,N_13193,N_12680);
xnor U13669 (N_13669,N_13072,N_12721);
xor U13670 (N_13670,N_12686,N_13102);
nor U13671 (N_13671,N_12975,N_12857);
and U13672 (N_13672,N_13059,N_12825);
or U13673 (N_13673,N_13083,N_12805);
nor U13674 (N_13674,N_13198,N_12756);
xnor U13675 (N_13675,N_12846,N_13103);
or U13676 (N_13676,N_12633,N_12877);
or U13677 (N_13677,N_12803,N_12960);
nand U13678 (N_13678,N_12634,N_12687);
nand U13679 (N_13679,N_12781,N_12812);
or U13680 (N_13680,N_12972,N_13046);
nor U13681 (N_13681,N_12629,N_12623);
nor U13682 (N_13682,N_12683,N_12694);
and U13683 (N_13683,N_13178,N_12762);
and U13684 (N_13684,N_12718,N_12839);
xor U13685 (N_13685,N_12758,N_12872);
nor U13686 (N_13686,N_13095,N_12840);
or U13687 (N_13687,N_12701,N_12831);
xnor U13688 (N_13688,N_12605,N_13007);
and U13689 (N_13689,N_13082,N_12682);
and U13690 (N_13690,N_13008,N_13123);
or U13691 (N_13691,N_13184,N_13125);
nand U13692 (N_13692,N_12886,N_12890);
or U13693 (N_13693,N_12796,N_13139);
or U13694 (N_13694,N_13080,N_12728);
nor U13695 (N_13695,N_12687,N_12819);
nand U13696 (N_13696,N_12981,N_12800);
nand U13697 (N_13697,N_12726,N_13134);
and U13698 (N_13698,N_12659,N_12938);
and U13699 (N_13699,N_12672,N_13180);
nand U13700 (N_13700,N_12919,N_12977);
and U13701 (N_13701,N_12623,N_12903);
and U13702 (N_13702,N_12721,N_12674);
and U13703 (N_13703,N_12910,N_13036);
and U13704 (N_13704,N_12705,N_12654);
or U13705 (N_13705,N_12650,N_13157);
xor U13706 (N_13706,N_12773,N_12871);
nand U13707 (N_13707,N_13178,N_12614);
or U13708 (N_13708,N_13162,N_12653);
nor U13709 (N_13709,N_12748,N_12723);
xnor U13710 (N_13710,N_13135,N_12854);
nor U13711 (N_13711,N_12717,N_12821);
nor U13712 (N_13712,N_12613,N_13169);
nand U13713 (N_13713,N_13127,N_12989);
nor U13714 (N_13714,N_13126,N_13029);
nand U13715 (N_13715,N_13087,N_13140);
nor U13716 (N_13716,N_12720,N_13163);
or U13717 (N_13717,N_13155,N_13098);
xor U13718 (N_13718,N_12633,N_13152);
or U13719 (N_13719,N_12836,N_12926);
and U13720 (N_13720,N_12766,N_12614);
and U13721 (N_13721,N_13024,N_12835);
nand U13722 (N_13722,N_13125,N_13004);
or U13723 (N_13723,N_12672,N_12852);
or U13724 (N_13724,N_12981,N_12731);
nor U13725 (N_13725,N_12866,N_13194);
nand U13726 (N_13726,N_12628,N_12642);
xnor U13727 (N_13727,N_12726,N_12919);
and U13728 (N_13728,N_12735,N_12967);
and U13729 (N_13729,N_12947,N_12932);
or U13730 (N_13730,N_13174,N_12670);
or U13731 (N_13731,N_12818,N_13190);
or U13732 (N_13732,N_13002,N_12693);
xor U13733 (N_13733,N_12846,N_12820);
nor U13734 (N_13734,N_13024,N_12838);
nor U13735 (N_13735,N_12953,N_12878);
or U13736 (N_13736,N_13192,N_12960);
or U13737 (N_13737,N_12931,N_12641);
and U13738 (N_13738,N_12811,N_12716);
xnor U13739 (N_13739,N_12924,N_12612);
nand U13740 (N_13740,N_12786,N_13043);
xor U13741 (N_13741,N_12828,N_12807);
and U13742 (N_13742,N_12921,N_13010);
nor U13743 (N_13743,N_12721,N_13103);
or U13744 (N_13744,N_12819,N_13172);
or U13745 (N_13745,N_12860,N_13146);
and U13746 (N_13746,N_12977,N_13174);
nor U13747 (N_13747,N_13194,N_12801);
xor U13748 (N_13748,N_13066,N_12767);
or U13749 (N_13749,N_13155,N_12685);
or U13750 (N_13750,N_12987,N_12606);
or U13751 (N_13751,N_12852,N_12623);
nor U13752 (N_13752,N_13047,N_12655);
or U13753 (N_13753,N_12851,N_13035);
xor U13754 (N_13754,N_12828,N_13012);
nand U13755 (N_13755,N_13079,N_13052);
nand U13756 (N_13756,N_12614,N_12885);
nor U13757 (N_13757,N_12658,N_13006);
or U13758 (N_13758,N_12651,N_13199);
and U13759 (N_13759,N_12609,N_12985);
and U13760 (N_13760,N_13169,N_13090);
xnor U13761 (N_13761,N_13192,N_13196);
nand U13762 (N_13762,N_13069,N_12744);
nand U13763 (N_13763,N_12807,N_12709);
nand U13764 (N_13764,N_12739,N_12674);
xnor U13765 (N_13765,N_12799,N_12930);
xnor U13766 (N_13766,N_12622,N_13126);
and U13767 (N_13767,N_12657,N_12718);
xnor U13768 (N_13768,N_13173,N_12918);
xnor U13769 (N_13769,N_12721,N_13169);
nand U13770 (N_13770,N_12910,N_12905);
or U13771 (N_13771,N_12951,N_13039);
xnor U13772 (N_13772,N_12902,N_12973);
nand U13773 (N_13773,N_12805,N_12608);
or U13774 (N_13774,N_13062,N_12606);
and U13775 (N_13775,N_12617,N_13063);
nor U13776 (N_13776,N_12671,N_12685);
xnor U13777 (N_13777,N_13150,N_13100);
or U13778 (N_13778,N_12616,N_13166);
xnor U13779 (N_13779,N_12668,N_12694);
xor U13780 (N_13780,N_12750,N_12612);
and U13781 (N_13781,N_12773,N_12748);
and U13782 (N_13782,N_12847,N_12833);
xor U13783 (N_13783,N_12733,N_12955);
nor U13784 (N_13784,N_13150,N_12899);
nand U13785 (N_13785,N_12919,N_13022);
xor U13786 (N_13786,N_13006,N_13133);
nor U13787 (N_13787,N_12850,N_12688);
or U13788 (N_13788,N_12891,N_12816);
or U13789 (N_13789,N_12770,N_13142);
and U13790 (N_13790,N_12825,N_12659);
or U13791 (N_13791,N_12863,N_13141);
or U13792 (N_13792,N_12682,N_12650);
nand U13793 (N_13793,N_12797,N_12833);
nor U13794 (N_13794,N_13155,N_13010);
and U13795 (N_13795,N_13176,N_12701);
nor U13796 (N_13796,N_12601,N_12860);
nor U13797 (N_13797,N_12724,N_12808);
or U13798 (N_13798,N_12716,N_13131);
and U13799 (N_13799,N_13095,N_13017);
xnor U13800 (N_13800,N_13415,N_13490);
or U13801 (N_13801,N_13506,N_13661);
xnor U13802 (N_13802,N_13410,N_13649);
and U13803 (N_13803,N_13309,N_13342);
xor U13804 (N_13804,N_13430,N_13634);
xnor U13805 (N_13805,N_13449,N_13717);
and U13806 (N_13806,N_13489,N_13285);
and U13807 (N_13807,N_13457,N_13647);
or U13808 (N_13808,N_13478,N_13334);
xnor U13809 (N_13809,N_13654,N_13364);
and U13810 (N_13810,N_13228,N_13480);
nand U13811 (N_13811,N_13281,N_13221);
and U13812 (N_13812,N_13709,N_13739);
and U13813 (N_13813,N_13770,N_13411);
nor U13814 (N_13814,N_13695,N_13249);
and U13815 (N_13815,N_13749,N_13635);
and U13816 (N_13816,N_13621,N_13322);
and U13817 (N_13817,N_13774,N_13338);
or U13818 (N_13818,N_13672,N_13656);
xnor U13819 (N_13819,N_13360,N_13768);
nand U13820 (N_13820,N_13252,N_13636);
or U13821 (N_13821,N_13556,N_13202);
nor U13822 (N_13822,N_13323,N_13355);
nor U13823 (N_13823,N_13592,N_13796);
and U13824 (N_13824,N_13623,N_13232);
and U13825 (N_13825,N_13353,N_13372);
and U13826 (N_13826,N_13555,N_13491);
xnor U13827 (N_13827,N_13648,N_13759);
or U13828 (N_13828,N_13629,N_13277);
xnor U13829 (N_13829,N_13744,N_13399);
or U13830 (N_13830,N_13312,N_13255);
or U13831 (N_13831,N_13513,N_13754);
or U13832 (N_13832,N_13423,N_13518);
nand U13833 (N_13833,N_13375,N_13791);
and U13834 (N_13834,N_13667,N_13406);
nor U13835 (N_13835,N_13272,N_13524);
nor U13836 (N_13836,N_13321,N_13225);
nand U13837 (N_13837,N_13377,N_13441);
or U13838 (N_13838,N_13563,N_13271);
and U13839 (N_13839,N_13533,N_13320);
and U13840 (N_13840,N_13397,N_13663);
and U13841 (N_13841,N_13664,N_13653);
nor U13842 (N_13842,N_13669,N_13628);
xnor U13843 (N_13843,N_13731,N_13409);
nor U13844 (N_13844,N_13729,N_13448);
and U13845 (N_13845,N_13598,N_13608);
nor U13846 (N_13846,N_13565,N_13504);
or U13847 (N_13847,N_13712,N_13226);
xnor U13848 (N_13848,N_13725,N_13660);
or U13849 (N_13849,N_13687,N_13436);
nor U13850 (N_13850,N_13548,N_13439);
nor U13851 (N_13851,N_13275,N_13203);
xor U13852 (N_13852,N_13704,N_13378);
nand U13853 (N_13853,N_13771,N_13218);
and U13854 (N_13854,N_13392,N_13696);
and U13855 (N_13855,N_13651,N_13760);
nor U13856 (N_13856,N_13434,N_13276);
and U13857 (N_13857,N_13568,N_13350);
nand U13858 (N_13858,N_13561,N_13476);
nor U13859 (N_13859,N_13456,N_13580);
nand U13860 (N_13860,N_13349,N_13671);
or U13861 (N_13861,N_13286,N_13597);
or U13862 (N_13862,N_13605,N_13590);
nand U13863 (N_13863,N_13753,N_13750);
nor U13864 (N_13864,N_13584,N_13694);
and U13865 (N_13865,N_13640,N_13677);
or U13866 (N_13866,N_13560,N_13201);
xor U13867 (N_13867,N_13740,N_13789);
or U13868 (N_13868,N_13401,N_13773);
xnor U13869 (N_13869,N_13359,N_13279);
nor U13870 (N_13870,N_13311,N_13784);
xnor U13871 (N_13871,N_13339,N_13497);
nor U13872 (N_13872,N_13413,N_13698);
or U13873 (N_13873,N_13777,N_13438);
and U13874 (N_13874,N_13668,N_13599);
and U13875 (N_13875,N_13676,N_13607);
nand U13876 (N_13876,N_13797,N_13588);
xor U13877 (N_13877,N_13317,N_13354);
and U13878 (N_13878,N_13546,N_13642);
nor U13879 (N_13879,N_13542,N_13270);
nand U13880 (N_13880,N_13529,N_13310);
or U13881 (N_13881,N_13540,N_13626);
or U13882 (N_13882,N_13673,N_13788);
nand U13883 (N_13883,N_13658,N_13313);
or U13884 (N_13884,N_13243,N_13303);
nor U13885 (N_13885,N_13785,N_13655);
xnor U13886 (N_13886,N_13421,N_13222);
xor U13887 (N_13887,N_13601,N_13500);
xor U13888 (N_13888,N_13611,N_13499);
xor U13889 (N_13889,N_13251,N_13559);
xnor U13890 (N_13890,N_13370,N_13408);
and U13891 (N_13891,N_13246,N_13319);
xor U13892 (N_13892,N_13324,N_13257);
and U13893 (N_13893,N_13643,N_13675);
or U13894 (N_13894,N_13470,N_13348);
nor U13895 (N_13895,N_13240,N_13236);
nand U13896 (N_13896,N_13767,N_13707);
and U13897 (N_13897,N_13520,N_13547);
nor U13898 (N_13898,N_13308,N_13267);
nand U13899 (N_13899,N_13213,N_13389);
nand U13900 (N_13900,N_13775,N_13443);
xor U13901 (N_13901,N_13570,N_13685);
nor U13902 (N_13902,N_13508,N_13437);
and U13903 (N_13903,N_13296,N_13790);
nor U13904 (N_13904,N_13525,N_13778);
or U13905 (N_13905,N_13371,N_13528);
and U13906 (N_13906,N_13289,N_13446);
nor U13907 (N_13907,N_13795,N_13216);
or U13908 (N_13908,N_13485,N_13517);
xnor U13909 (N_13909,N_13666,N_13404);
or U13910 (N_13910,N_13557,N_13301);
and U13911 (N_13911,N_13341,N_13724);
and U13912 (N_13912,N_13428,N_13644);
or U13913 (N_13913,N_13425,N_13328);
xor U13914 (N_13914,N_13776,N_13674);
nor U13915 (N_13915,N_13701,N_13210);
or U13916 (N_13916,N_13587,N_13535);
or U13917 (N_13917,N_13769,N_13764);
nor U13918 (N_13918,N_13234,N_13420);
xor U13919 (N_13919,N_13248,N_13365);
nand U13920 (N_13920,N_13783,N_13381);
xnor U13921 (N_13921,N_13288,N_13624);
nor U13922 (N_13922,N_13742,N_13702);
or U13923 (N_13923,N_13627,N_13385);
nand U13924 (N_13924,N_13299,N_13551);
or U13925 (N_13925,N_13575,N_13356);
xor U13926 (N_13926,N_13435,N_13250);
or U13927 (N_13927,N_13393,N_13733);
nor U13928 (N_13928,N_13606,N_13268);
xor U13929 (N_13929,N_13798,N_13610);
or U13930 (N_13930,N_13297,N_13625);
nand U13931 (N_13931,N_13569,N_13466);
xor U13932 (N_13932,N_13501,N_13464);
xor U13933 (N_13933,N_13207,N_13617);
and U13934 (N_13934,N_13532,N_13473);
nor U13935 (N_13935,N_13332,N_13427);
nor U13936 (N_13936,N_13206,N_13612);
xor U13937 (N_13937,N_13444,N_13429);
or U13938 (N_13938,N_13343,N_13209);
or U13939 (N_13939,N_13572,N_13762);
xnor U13940 (N_13940,N_13387,N_13755);
nand U13941 (N_13941,N_13614,N_13283);
nor U13942 (N_13942,N_13720,N_13550);
nor U13943 (N_13943,N_13521,N_13467);
nor U13944 (N_13944,N_13619,N_13458);
nand U13945 (N_13945,N_13689,N_13361);
nand U13946 (N_13946,N_13215,N_13505);
xnor U13947 (N_13947,N_13242,N_13477);
or U13948 (N_13948,N_13600,N_13552);
or U13949 (N_13949,N_13486,N_13287);
xnor U13950 (N_13950,N_13734,N_13541);
xor U13951 (N_13951,N_13578,N_13693);
or U13952 (N_13952,N_13418,N_13705);
xnor U13953 (N_13953,N_13722,N_13678);
nor U13954 (N_13954,N_13223,N_13493);
nor U13955 (N_13955,N_13442,N_13602);
nand U13956 (N_13956,N_13639,N_13238);
nand U13957 (N_13957,N_13307,N_13424);
and U13958 (N_13958,N_13522,N_13264);
xnor U13959 (N_13959,N_13609,N_13657);
xnor U13960 (N_13960,N_13692,N_13645);
or U13961 (N_13961,N_13659,N_13732);
and U13962 (N_13962,N_13567,N_13779);
xnor U13963 (N_13963,N_13214,N_13217);
xor U13964 (N_13964,N_13258,N_13670);
nor U13965 (N_13965,N_13380,N_13682);
nand U13966 (N_13966,N_13727,N_13719);
nor U13967 (N_13967,N_13579,N_13266);
or U13968 (N_13968,N_13752,N_13582);
xnor U13969 (N_13969,N_13262,N_13507);
or U13970 (N_13970,N_13453,N_13713);
or U13971 (N_13971,N_13412,N_13714);
and U13972 (N_13972,N_13756,N_13468);
or U13973 (N_13973,N_13703,N_13333);
nor U13974 (N_13974,N_13589,N_13683);
nand U13975 (N_13975,N_13315,N_13745);
and U13976 (N_13976,N_13260,N_13400);
or U13977 (N_13977,N_13405,N_13261);
xnor U13978 (N_13978,N_13259,N_13616);
or U13979 (N_13979,N_13498,N_13761);
or U13980 (N_13980,N_13204,N_13382);
xnor U13981 (N_13981,N_13794,N_13593);
and U13982 (N_13982,N_13273,N_13472);
nand U13983 (N_13983,N_13331,N_13562);
nor U13984 (N_13984,N_13454,N_13586);
nand U13985 (N_13985,N_13536,N_13509);
or U13986 (N_13986,N_13487,N_13245);
nor U13987 (N_13987,N_13736,N_13447);
and U13988 (N_13988,N_13316,N_13706);
and U13989 (N_13989,N_13269,N_13366);
or U13990 (N_13990,N_13554,N_13479);
nand U13991 (N_13991,N_13553,N_13481);
nor U13992 (N_13992,N_13633,N_13632);
nand U13993 (N_13993,N_13594,N_13743);
xor U13994 (N_13994,N_13716,N_13256);
or U13995 (N_13995,N_13646,N_13200);
nor U13996 (N_13996,N_13686,N_13576);
nand U13997 (N_13997,N_13780,N_13537);
and U13998 (N_13998,N_13335,N_13662);
nand U13999 (N_13999,N_13726,N_13715);
and U14000 (N_14000,N_13208,N_13205);
or U14001 (N_14001,N_13220,N_13314);
nand U14002 (N_14002,N_13294,N_13585);
nor U14003 (N_14003,N_13302,N_13679);
or U14004 (N_14004,N_13304,N_13337);
or U14005 (N_14005,N_13566,N_13402);
or U14006 (N_14006,N_13665,N_13363);
xnor U14007 (N_14007,N_13306,N_13748);
nand U14008 (N_14008,N_13298,N_13613);
and U14009 (N_14009,N_13708,N_13741);
or U14010 (N_14010,N_13539,N_13414);
nand U14011 (N_14011,N_13384,N_13792);
and U14012 (N_14012,N_13581,N_13545);
xor U14013 (N_14013,N_13326,N_13511);
or U14014 (N_14014,N_13786,N_13390);
and U14015 (N_14015,N_13765,N_13358);
nor U14016 (N_14016,N_13475,N_13227);
nand U14017 (N_14017,N_13422,N_13357);
or U14018 (N_14018,N_13515,N_13737);
and U14019 (N_14019,N_13431,N_13465);
xnor U14020 (N_14020,N_13318,N_13231);
xnor U14021 (N_14021,N_13224,N_13793);
and U14022 (N_14022,N_13688,N_13530);
xnor U14023 (N_14023,N_13351,N_13631);
or U14024 (N_14024,N_13280,N_13212);
xor U14025 (N_14025,N_13230,N_13253);
and U14026 (N_14026,N_13403,N_13379);
xnor U14027 (N_14027,N_13388,N_13690);
xor U14028 (N_14028,N_13305,N_13758);
xor U14029 (N_14029,N_13782,N_13700);
nand U14030 (N_14030,N_13416,N_13751);
nor U14031 (N_14031,N_13383,N_13757);
or U14032 (N_14032,N_13766,N_13650);
nand U14033 (N_14033,N_13325,N_13398);
xor U14034 (N_14034,N_13583,N_13235);
xor U14035 (N_14035,N_13461,N_13241);
xor U14036 (N_14036,N_13526,N_13352);
nand U14037 (N_14037,N_13391,N_13274);
and U14038 (N_14038,N_13503,N_13367);
nand U14039 (N_14039,N_13345,N_13284);
and U14040 (N_14040,N_13419,N_13211);
nor U14041 (N_14041,N_13394,N_13327);
and U14042 (N_14042,N_13718,N_13638);
nand U14043 (N_14043,N_13620,N_13492);
nand U14044 (N_14044,N_13482,N_13573);
nor U14045 (N_14045,N_13558,N_13455);
and U14046 (N_14046,N_13538,N_13219);
or U14047 (N_14047,N_13596,N_13329);
nand U14048 (N_14048,N_13738,N_13781);
or U14049 (N_14049,N_13293,N_13571);
xnor U14050 (N_14050,N_13374,N_13502);
or U14051 (N_14051,N_13747,N_13591);
or U14052 (N_14052,N_13799,N_13291);
or U14053 (N_14053,N_13637,N_13395);
or U14054 (N_14054,N_13344,N_13787);
nand U14055 (N_14055,N_13463,N_13721);
or U14056 (N_14056,N_13495,N_13233);
or U14057 (N_14057,N_13534,N_13254);
or U14058 (N_14058,N_13746,N_13452);
or U14059 (N_14059,N_13484,N_13462);
xnor U14060 (N_14060,N_13265,N_13723);
nor U14061 (N_14061,N_13451,N_13433);
or U14062 (N_14062,N_13330,N_13512);
or U14063 (N_14063,N_13516,N_13728);
xor U14064 (N_14064,N_13244,N_13603);
nand U14065 (N_14065,N_13369,N_13450);
nand U14066 (N_14066,N_13469,N_13630);
xor U14067 (N_14067,N_13460,N_13362);
nor U14068 (N_14068,N_13615,N_13595);
nor U14069 (N_14069,N_13510,N_13496);
nand U14070 (N_14070,N_13459,N_13549);
nor U14071 (N_14071,N_13735,N_13697);
or U14072 (N_14072,N_13229,N_13396);
and U14073 (N_14073,N_13523,N_13368);
nand U14074 (N_14074,N_13488,N_13622);
nor U14075 (N_14075,N_13263,N_13681);
nand U14076 (N_14076,N_13531,N_13292);
xor U14077 (N_14077,N_13426,N_13543);
nor U14078 (N_14078,N_13699,N_13684);
or U14079 (N_14079,N_13376,N_13247);
or U14080 (N_14080,N_13574,N_13346);
and U14081 (N_14081,N_13527,N_13483);
or U14082 (N_14082,N_13440,N_13386);
nor U14083 (N_14083,N_13577,N_13432);
or U14084 (N_14084,N_13730,N_13295);
nor U14085 (N_14085,N_13641,N_13544);
nor U14086 (N_14086,N_13471,N_13336);
and U14087 (N_14087,N_13494,N_13710);
nand U14088 (N_14088,N_13474,N_13680);
and U14089 (N_14089,N_13237,N_13278);
xor U14090 (N_14090,N_13239,N_13519);
nand U14091 (N_14091,N_13300,N_13340);
or U14092 (N_14092,N_13763,N_13711);
xor U14093 (N_14093,N_13407,N_13290);
nor U14094 (N_14094,N_13282,N_13604);
xor U14095 (N_14095,N_13373,N_13618);
or U14096 (N_14096,N_13514,N_13691);
xor U14097 (N_14097,N_13772,N_13652);
xnor U14098 (N_14098,N_13417,N_13564);
nand U14099 (N_14099,N_13347,N_13445);
nor U14100 (N_14100,N_13734,N_13394);
nor U14101 (N_14101,N_13359,N_13694);
and U14102 (N_14102,N_13268,N_13216);
and U14103 (N_14103,N_13574,N_13351);
and U14104 (N_14104,N_13764,N_13575);
xor U14105 (N_14105,N_13497,N_13547);
nor U14106 (N_14106,N_13689,N_13209);
and U14107 (N_14107,N_13504,N_13611);
xnor U14108 (N_14108,N_13232,N_13590);
nand U14109 (N_14109,N_13733,N_13453);
nand U14110 (N_14110,N_13446,N_13583);
or U14111 (N_14111,N_13461,N_13202);
or U14112 (N_14112,N_13343,N_13702);
xor U14113 (N_14113,N_13337,N_13316);
or U14114 (N_14114,N_13265,N_13497);
nand U14115 (N_14115,N_13712,N_13353);
nand U14116 (N_14116,N_13331,N_13226);
nor U14117 (N_14117,N_13399,N_13395);
xnor U14118 (N_14118,N_13324,N_13447);
nand U14119 (N_14119,N_13748,N_13639);
or U14120 (N_14120,N_13774,N_13247);
nor U14121 (N_14121,N_13788,N_13219);
or U14122 (N_14122,N_13317,N_13325);
nand U14123 (N_14123,N_13368,N_13421);
and U14124 (N_14124,N_13439,N_13398);
or U14125 (N_14125,N_13744,N_13356);
nand U14126 (N_14126,N_13713,N_13739);
and U14127 (N_14127,N_13741,N_13563);
xor U14128 (N_14128,N_13389,N_13408);
and U14129 (N_14129,N_13219,N_13548);
xnor U14130 (N_14130,N_13251,N_13596);
or U14131 (N_14131,N_13516,N_13285);
or U14132 (N_14132,N_13658,N_13720);
and U14133 (N_14133,N_13343,N_13618);
and U14134 (N_14134,N_13387,N_13200);
or U14135 (N_14135,N_13580,N_13559);
and U14136 (N_14136,N_13452,N_13625);
nor U14137 (N_14137,N_13263,N_13723);
or U14138 (N_14138,N_13780,N_13762);
nand U14139 (N_14139,N_13296,N_13789);
nor U14140 (N_14140,N_13536,N_13205);
or U14141 (N_14141,N_13562,N_13716);
and U14142 (N_14142,N_13208,N_13433);
or U14143 (N_14143,N_13200,N_13371);
xor U14144 (N_14144,N_13232,N_13349);
or U14145 (N_14145,N_13359,N_13434);
nand U14146 (N_14146,N_13579,N_13795);
xor U14147 (N_14147,N_13436,N_13476);
and U14148 (N_14148,N_13781,N_13540);
xor U14149 (N_14149,N_13491,N_13389);
xnor U14150 (N_14150,N_13212,N_13357);
nand U14151 (N_14151,N_13719,N_13601);
nand U14152 (N_14152,N_13569,N_13587);
nand U14153 (N_14153,N_13715,N_13490);
xnor U14154 (N_14154,N_13400,N_13627);
or U14155 (N_14155,N_13309,N_13684);
xor U14156 (N_14156,N_13446,N_13295);
nor U14157 (N_14157,N_13683,N_13371);
xnor U14158 (N_14158,N_13750,N_13632);
nand U14159 (N_14159,N_13308,N_13654);
and U14160 (N_14160,N_13771,N_13512);
and U14161 (N_14161,N_13542,N_13715);
nand U14162 (N_14162,N_13232,N_13543);
or U14163 (N_14163,N_13788,N_13534);
nor U14164 (N_14164,N_13398,N_13628);
and U14165 (N_14165,N_13389,N_13208);
nor U14166 (N_14166,N_13782,N_13721);
and U14167 (N_14167,N_13499,N_13561);
nand U14168 (N_14168,N_13204,N_13400);
and U14169 (N_14169,N_13648,N_13299);
or U14170 (N_14170,N_13658,N_13606);
and U14171 (N_14171,N_13738,N_13286);
nor U14172 (N_14172,N_13692,N_13764);
xor U14173 (N_14173,N_13302,N_13771);
xnor U14174 (N_14174,N_13733,N_13375);
nand U14175 (N_14175,N_13607,N_13704);
nor U14176 (N_14176,N_13720,N_13513);
and U14177 (N_14177,N_13282,N_13541);
nor U14178 (N_14178,N_13416,N_13517);
nand U14179 (N_14179,N_13504,N_13480);
nand U14180 (N_14180,N_13536,N_13549);
nor U14181 (N_14181,N_13557,N_13223);
nor U14182 (N_14182,N_13691,N_13710);
nor U14183 (N_14183,N_13423,N_13364);
nor U14184 (N_14184,N_13279,N_13353);
nor U14185 (N_14185,N_13787,N_13448);
nand U14186 (N_14186,N_13512,N_13796);
nor U14187 (N_14187,N_13228,N_13360);
xor U14188 (N_14188,N_13678,N_13326);
and U14189 (N_14189,N_13509,N_13236);
or U14190 (N_14190,N_13561,N_13473);
nand U14191 (N_14191,N_13646,N_13696);
or U14192 (N_14192,N_13731,N_13710);
nor U14193 (N_14193,N_13766,N_13786);
and U14194 (N_14194,N_13393,N_13452);
nand U14195 (N_14195,N_13484,N_13202);
xor U14196 (N_14196,N_13273,N_13721);
nor U14197 (N_14197,N_13270,N_13768);
xnor U14198 (N_14198,N_13713,N_13293);
xor U14199 (N_14199,N_13661,N_13740);
and U14200 (N_14200,N_13635,N_13538);
or U14201 (N_14201,N_13332,N_13690);
xor U14202 (N_14202,N_13723,N_13267);
nor U14203 (N_14203,N_13343,N_13337);
or U14204 (N_14204,N_13586,N_13564);
xor U14205 (N_14205,N_13504,N_13528);
or U14206 (N_14206,N_13741,N_13565);
xnor U14207 (N_14207,N_13316,N_13489);
and U14208 (N_14208,N_13231,N_13752);
nand U14209 (N_14209,N_13660,N_13743);
and U14210 (N_14210,N_13795,N_13390);
nand U14211 (N_14211,N_13556,N_13367);
nand U14212 (N_14212,N_13547,N_13515);
or U14213 (N_14213,N_13625,N_13745);
nand U14214 (N_14214,N_13585,N_13746);
nor U14215 (N_14215,N_13200,N_13311);
nand U14216 (N_14216,N_13302,N_13277);
or U14217 (N_14217,N_13291,N_13278);
xnor U14218 (N_14218,N_13737,N_13310);
nor U14219 (N_14219,N_13252,N_13248);
nand U14220 (N_14220,N_13404,N_13348);
and U14221 (N_14221,N_13435,N_13718);
or U14222 (N_14222,N_13417,N_13518);
xnor U14223 (N_14223,N_13297,N_13534);
nor U14224 (N_14224,N_13743,N_13338);
or U14225 (N_14225,N_13567,N_13782);
and U14226 (N_14226,N_13437,N_13556);
or U14227 (N_14227,N_13309,N_13759);
and U14228 (N_14228,N_13425,N_13781);
xor U14229 (N_14229,N_13229,N_13554);
or U14230 (N_14230,N_13728,N_13235);
and U14231 (N_14231,N_13392,N_13202);
and U14232 (N_14232,N_13637,N_13280);
xor U14233 (N_14233,N_13475,N_13212);
nand U14234 (N_14234,N_13427,N_13538);
or U14235 (N_14235,N_13550,N_13689);
nor U14236 (N_14236,N_13275,N_13491);
nor U14237 (N_14237,N_13473,N_13518);
xnor U14238 (N_14238,N_13268,N_13680);
or U14239 (N_14239,N_13364,N_13486);
and U14240 (N_14240,N_13580,N_13590);
nor U14241 (N_14241,N_13625,N_13596);
nor U14242 (N_14242,N_13373,N_13328);
xnor U14243 (N_14243,N_13702,N_13299);
and U14244 (N_14244,N_13700,N_13496);
and U14245 (N_14245,N_13394,N_13499);
or U14246 (N_14246,N_13309,N_13392);
nor U14247 (N_14247,N_13707,N_13690);
nor U14248 (N_14248,N_13334,N_13652);
and U14249 (N_14249,N_13677,N_13779);
and U14250 (N_14250,N_13459,N_13487);
and U14251 (N_14251,N_13400,N_13771);
and U14252 (N_14252,N_13459,N_13401);
or U14253 (N_14253,N_13491,N_13353);
xnor U14254 (N_14254,N_13409,N_13633);
nand U14255 (N_14255,N_13659,N_13777);
and U14256 (N_14256,N_13326,N_13680);
and U14257 (N_14257,N_13264,N_13613);
or U14258 (N_14258,N_13707,N_13337);
nand U14259 (N_14259,N_13308,N_13515);
nand U14260 (N_14260,N_13728,N_13532);
xor U14261 (N_14261,N_13541,N_13757);
nor U14262 (N_14262,N_13351,N_13525);
nor U14263 (N_14263,N_13513,N_13384);
nand U14264 (N_14264,N_13602,N_13326);
or U14265 (N_14265,N_13327,N_13406);
or U14266 (N_14266,N_13549,N_13448);
nand U14267 (N_14267,N_13763,N_13620);
or U14268 (N_14268,N_13560,N_13216);
xor U14269 (N_14269,N_13675,N_13588);
xnor U14270 (N_14270,N_13437,N_13654);
nor U14271 (N_14271,N_13623,N_13748);
xnor U14272 (N_14272,N_13276,N_13335);
and U14273 (N_14273,N_13723,N_13410);
nor U14274 (N_14274,N_13686,N_13698);
nor U14275 (N_14275,N_13302,N_13510);
and U14276 (N_14276,N_13573,N_13771);
xnor U14277 (N_14277,N_13498,N_13435);
or U14278 (N_14278,N_13448,N_13604);
nand U14279 (N_14279,N_13562,N_13774);
nand U14280 (N_14280,N_13237,N_13436);
nand U14281 (N_14281,N_13648,N_13745);
and U14282 (N_14282,N_13712,N_13436);
or U14283 (N_14283,N_13437,N_13308);
or U14284 (N_14284,N_13346,N_13335);
or U14285 (N_14285,N_13485,N_13293);
and U14286 (N_14286,N_13483,N_13322);
nand U14287 (N_14287,N_13271,N_13461);
nand U14288 (N_14288,N_13599,N_13610);
or U14289 (N_14289,N_13728,N_13315);
nor U14290 (N_14290,N_13477,N_13703);
and U14291 (N_14291,N_13690,N_13616);
nor U14292 (N_14292,N_13245,N_13428);
nor U14293 (N_14293,N_13626,N_13444);
and U14294 (N_14294,N_13347,N_13325);
or U14295 (N_14295,N_13631,N_13225);
nor U14296 (N_14296,N_13636,N_13677);
or U14297 (N_14297,N_13203,N_13776);
nand U14298 (N_14298,N_13398,N_13449);
or U14299 (N_14299,N_13404,N_13656);
and U14300 (N_14300,N_13314,N_13470);
and U14301 (N_14301,N_13432,N_13240);
or U14302 (N_14302,N_13328,N_13346);
and U14303 (N_14303,N_13581,N_13575);
or U14304 (N_14304,N_13457,N_13423);
or U14305 (N_14305,N_13522,N_13733);
and U14306 (N_14306,N_13245,N_13752);
or U14307 (N_14307,N_13545,N_13276);
xnor U14308 (N_14308,N_13509,N_13709);
or U14309 (N_14309,N_13488,N_13561);
xnor U14310 (N_14310,N_13421,N_13320);
xnor U14311 (N_14311,N_13552,N_13566);
xor U14312 (N_14312,N_13272,N_13751);
nor U14313 (N_14313,N_13507,N_13624);
or U14314 (N_14314,N_13552,N_13588);
or U14315 (N_14315,N_13664,N_13222);
or U14316 (N_14316,N_13600,N_13440);
and U14317 (N_14317,N_13403,N_13425);
nor U14318 (N_14318,N_13295,N_13640);
xnor U14319 (N_14319,N_13513,N_13582);
nor U14320 (N_14320,N_13634,N_13551);
and U14321 (N_14321,N_13510,N_13700);
xnor U14322 (N_14322,N_13315,N_13333);
or U14323 (N_14323,N_13252,N_13575);
and U14324 (N_14324,N_13494,N_13708);
xnor U14325 (N_14325,N_13712,N_13660);
or U14326 (N_14326,N_13546,N_13685);
nand U14327 (N_14327,N_13358,N_13592);
nor U14328 (N_14328,N_13320,N_13679);
and U14329 (N_14329,N_13485,N_13691);
and U14330 (N_14330,N_13317,N_13267);
nor U14331 (N_14331,N_13388,N_13294);
xnor U14332 (N_14332,N_13762,N_13537);
xor U14333 (N_14333,N_13516,N_13561);
nor U14334 (N_14334,N_13597,N_13225);
nand U14335 (N_14335,N_13590,N_13459);
or U14336 (N_14336,N_13516,N_13646);
or U14337 (N_14337,N_13386,N_13309);
and U14338 (N_14338,N_13700,N_13212);
and U14339 (N_14339,N_13676,N_13627);
or U14340 (N_14340,N_13613,N_13506);
or U14341 (N_14341,N_13448,N_13462);
nor U14342 (N_14342,N_13254,N_13712);
nand U14343 (N_14343,N_13587,N_13447);
or U14344 (N_14344,N_13705,N_13663);
and U14345 (N_14345,N_13704,N_13719);
and U14346 (N_14346,N_13681,N_13492);
nand U14347 (N_14347,N_13768,N_13207);
or U14348 (N_14348,N_13750,N_13511);
nand U14349 (N_14349,N_13588,N_13712);
nand U14350 (N_14350,N_13360,N_13490);
or U14351 (N_14351,N_13609,N_13246);
xor U14352 (N_14352,N_13683,N_13212);
and U14353 (N_14353,N_13747,N_13608);
and U14354 (N_14354,N_13389,N_13418);
nor U14355 (N_14355,N_13436,N_13489);
xnor U14356 (N_14356,N_13425,N_13363);
xnor U14357 (N_14357,N_13463,N_13708);
nor U14358 (N_14358,N_13255,N_13729);
nand U14359 (N_14359,N_13361,N_13546);
or U14360 (N_14360,N_13654,N_13248);
or U14361 (N_14361,N_13239,N_13306);
nand U14362 (N_14362,N_13501,N_13604);
or U14363 (N_14363,N_13529,N_13341);
nand U14364 (N_14364,N_13268,N_13355);
and U14365 (N_14365,N_13788,N_13718);
xor U14366 (N_14366,N_13433,N_13779);
xnor U14367 (N_14367,N_13321,N_13626);
nand U14368 (N_14368,N_13484,N_13294);
or U14369 (N_14369,N_13733,N_13588);
and U14370 (N_14370,N_13529,N_13214);
nor U14371 (N_14371,N_13685,N_13326);
xor U14372 (N_14372,N_13410,N_13280);
and U14373 (N_14373,N_13717,N_13518);
nand U14374 (N_14374,N_13233,N_13257);
xnor U14375 (N_14375,N_13452,N_13235);
nand U14376 (N_14376,N_13533,N_13571);
and U14377 (N_14377,N_13477,N_13248);
nand U14378 (N_14378,N_13425,N_13236);
and U14379 (N_14379,N_13221,N_13546);
or U14380 (N_14380,N_13291,N_13781);
and U14381 (N_14381,N_13296,N_13740);
or U14382 (N_14382,N_13599,N_13492);
and U14383 (N_14383,N_13216,N_13757);
and U14384 (N_14384,N_13777,N_13332);
nor U14385 (N_14385,N_13638,N_13538);
or U14386 (N_14386,N_13641,N_13475);
and U14387 (N_14387,N_13776,N_13531);
xor U14388 (N_14388,N_13361,N_13549);
nor U14389 (N_14389,N_13399,N_13543);
nor U14390 (N_14390,N_13422,N_13424);
or U14391 (N_14391,N_13386,N_13799);
nand U14392 (N_14392,N_13388,N_13562);
xor U14393 (N_14393,N_13245,N_13411);
nand U14394 (N_14394,N_13334,N_13592);
nor U14395 (N_14395,N_13359,N_13410);
nand U14396 (N_14396,N_13577,N_13310);
and U14397 (N_14397,N_13555,N_13345);
xnor U14398 (N_14398,N_13605,N_13334);
and U14399 (N_14399,N_13544,N_13747);
nand U14400 (N_14400,N_14314,N_14369);
nand U14401 (N_14401,N_14169,N_14221);
or U14402 (N_14402,N_13830,N_14237);
or U14403 (N_14403,N_14261,N_14062);
xnor U14404 (N_14404,N_13806,N_14027);
nor U14405 (N_14405,N_14194,N_13834);
and U14406 (N_14406,N_13882,N_14165);
nor U14407 (N_14407,N_13928,N_14344);
and U14408 (N_14408,N_14111,N_14322);
nor U14409 (N_14409,N_13943,N_14370);
xnor U14410 (N_14410,N_14351,N_14391);
and U14411 (N_14411,N_14039,N_14392);
nand U14412 (N_14412,N_14230,N_13946);
and U14413 (N_14413,N_14166,N_14247);
nand U14414 (N_14414,N_14206,N_14227);
nand U14415 (N_14415,N_13888,N_13923);
nor U14416 (N_14416,N_13853,N_13885);
and U14417 (N_14417,N_13974,N_13931);
nand U14418 (N_14418,N_14080,N_14071);
or U14419 (N_14419,N_14297,N_14362);
and U14420 (N_14420,N_14152,N_14063);
and U14421 (N_14421,N_14304,N_14271);
or U14422 (N_14422,N_14382,N_14375);
xor U14423 (N_14423,N_14002,N_14296);
xnor U14424 (N_14424,N_14018,N_14195);
and U14425 (N_14425,N_14270,N_14276);
nand U14426 (N_14426,N_14277,N_14098);
xnor U14427 (N_14427,N_13994,N_13881);
xor U14428 (N_14428,N_13933,N_14145);
or U14429 (N_14429,N_14100,N_14081);
or U14430 (N_14430,N_14174,N_14191);
nand U14431 (N_14431,N_14396,N_14015);
nand U14432 (N_14432,N_14102,N_14216);
and U14433 (N_14433,N_14170,N_14163);
nand U14434 (N_14434,N_14073,N_14265);
or U14435 (N_14435,N_14380,N_14243);
nand U14436 (N_14436,N_14184,N_14125);
or U14437 (N_14437,N_14017,N_14309);
xnor U14438 (N_14438,N_14006,N_14151);
and U14439 (N_14439,N_13847,N_14354);
or U14440 (N_14440,N_14346,N_13969);
and U14441 (N_14441,N_14058,N_14241);
xnor U14442 (N_14442,N_13808,N_13907);
or U14443 (N_14443,N_14156,N_14334);
nand U14444 (N_14444,N_14341,N_14105);
xnor U14445 (N_14445,N_14229,N_13859);
and U14446 (N_14446,N_13942,N_13915);
nor U14447 (N_14447,N_13843,N_14342);
and U14448 (N_14448,N_14025,N_14364);
or U14449 (N_14449,N_14262,N_13913);
or U14450 (N_14450,N_14150,N_14371);
nor U14451 (N_14451,N_14385,N_14088);
nand U14452 (N_14452,N_13944,N_14000);
nand U14453 (N_14453,N_14246,N_14070);
and U14454 (N_14454,N_14272,N_14094);
or U14455 (N_14455,N_14122,N_13892);
xnor U14456 (N_14456,N_13871,N_14175);
xor U14457 (N_14457,N_14007,N_14303);
xnor U14458 (N_14458,N_14257,N_13980);
and U14459 (N_14459,N_14263,N_13821);
nor U14460 (N_14460,N_14137,N_14008);
and U14461 (N_14461,N_14146,N_13864);
nor U14462 (N_14462,N_13873,N_13813);
nand U14463 (N_14463,N_13833,N_14386);
and U14464 (N_14464,N_13935,N_13901);
and U14465 (N_14465,N_13908,N_14235);
and U14466 (N_14466,N_14343,N_14160);
xor U14467 (N_14467,N_14238,N_13848);
xnor U14468 (N_14468,N_14057,N_14016);
xnor U14469 (N_14469,N_13890,N_14179);
nor U14470 (N_14470,N_14345,N_13809);
nand U14471 (N_14471,N_13953,N_14124);
and U14472 (N_14472,N_13920,N_13996);
nand U14473 (N_14473,N_14273,N_13875);
nor U14474 (N_14474,N_14110,N_14209);
nand U14475 (N_14475,N_13831,N_14089);
and U14476 (N_14476,N_13891,N_14168);
xor U14477 (N_14477,N_13984,N_14126);
nor U14478 (N_14478,N_14260,N_13869);
xnor U14479 (N_14479,N_14144,N_14042);
or U14480 (N_14480,N_14225,N_14255);
or U14481 (N_14481,N_14250,N_14210);
or U14482 (N_14482,N_14218,N_14035);
nand U14483 (N_14483,N_13826,N_13965);
nor U14484 (N_14484,N_13812,N_13835);
or U14485 (N_14485,N_13815,N_13878);
nand U14486 (N_14486,N_13949,N_14038);
nand U14487 (N_14487,N_14004,N_14101);
and U14488 (N_14488,N_13962,N_14056);
or U14489 (N_14489,N_13870,N_13865);
nand U14490 (N_14490,N_14041,N_14139);
nand U14491 (N_14491,N_14381,N_14248);
xor U14492 (N_14492,N_14350,N_13836);
xnor U14493 (N_14493,N_14307,N_14316);
and U14494 (N_14494,N_14352,N_14136);
or U14495 (N_14495,N_14109,N_14357);
or U14496 (N_14496,N_14368,N_14107);
nand U14497 (N_14497,N_13868,N_14065);
xnor U14498 (N_14498,N_14275,N_14298);
xnor U14499 (N_14499,N_14176,N_13905);
xor U14500 (N_14500,N_13818,N_14133);
nand U14501 (N_14501,N_13880,N_14361);
nor U14502 (N_14502,N_13898,N_14161);
or U14503 (N_14503,N_13958,N_13828);
nor U14504 (N_14504,N_14299,N_13840);
xor U14505 (N_14505,N_13910,N_14326);
or U14506 (N_14506,N_14045,N_14055);
nor U14507 (N_14507,N_14023,N_13927);
nand U14508 (N_14508,N_14116,N_14212);
nand U14509 (N_14509,N_14009,N_14164);
xor U14510 (N_14510,N_14249,N_13954);
nand U14511 (N_14511,N_13924,N_14205);
and U14512 (N_14512,N_14019,N_14214);
or U14513 (N_14513,N_14177,N_14220);
xor U14514 (N_14514,N_14189,N_14388);
or U14515 (N_14515,N_14037,N_14399);
nor U14516 (N_14516,N_14384,N_14284);
xnor U14517 (N_14517,N_14286,N_13981);
or U14518 (N_14518,N_14279,N_14213);
and U14519 (N_14519,N_14117,N_14372);
nand U14520 (N_14520,N_13998,N_14077);
nor U14521 (N_14521,N_13872,N_13976);
or U14522 (N_14522,N_14320,N_14092);
and U14523 (N_14523,N_14087,N_13919);
nand U14524 (N_14524,N_14099,N_13900);
xnor U14525 (N_14525,N_14329,N_14049);
or U14526 (N_14526,N_13992,N_14367);
and U14527 (N_14527,N_13961,N_14256);
or U14528 (N_14528,N_14069,N_14294);
nand U14529 (N_14529,N_14389,N_14028);
xor U14530 (N_14530,N_14252,N_13987);
or U14531 (N_14531,N_14112,N_13879);
and U14532 (N_14532,N_14202,N_14291);
and U14533 (N_14533,N_14026,N_13801);
xnor U14534 (N_14534,N_13916,N_14355);
nor U14535 (N_14535,N_14143,N_14233);
xor U14536 (N_14536,N_13862,N_13842);
or U14537 (N_14537,N_13999,N_14190);
xnor U14538 (N_14538,N_14197,N_14106);
or U14539 (N_14539,N_14387,N_13805);
or U14540 (N_14540,N_14050,N_14280);
and U14541 (N_14541,N_13811,N_14103);
and U14542 (N_14542,N_14236,N_13971);
nand U14543 (N_14543,N_14234,N_14231);
nand U14544 (N_14544,N_14390,N_14155);
and U14545 (N_14545,N_13968,N_13918);
and U14546 (N_14546,N_14223,N_13829);
and U14547 (N_14547,N_13963,N_14226);
nor U14548 (N_14548,N_14131,N_13903);
or U14549 (N_14549,N_14181,N_14118);
or U14550 (N_14550,N_14259,N_14091);
nand U14551 (N_14551,N_14158,N_13816);
and U14552 (N_14552,N_13964,N_14147);
nand U14553 (N_14553,N_14066,N_14365);
nand U14554 (N_14554,N_13948,N_13986);
nor U14555 (N_14555,N_14266,N_14132);
xnor U14556 (N_14556,N_13852,N_13912);
xor U14557 (N_14557,N_13938,N_14327);
nor U14558 (N_14558,N_14325,N_14353);
and U14559 (N_14559,N_14356,N_14185);
xnor U14560 (N_14560,N_13883,N_14032);
or U14561 (N_14561,N_13951,N_14217);
nand U14562 (N_14562,N_14306,N_14013);
xnor U14563 (N_14563,N_13950,N_14211);
or U14564 (N_14564,N_14075,N_14383);
or U14565 (N_14565,N_13988,N_13858);
or U14566 (N_14566,N_14059,N_14076);
xnor U14567 (N_14567,N_13838,N_14047);
and U14568 (N_14568,N_14173,N_14090);
and U14569 (N_14569,N_14064,N_14287);
nor U14570 (N_14570,N_14119,N_13997);
xnor U14571 (N_14571,N_13934,N_14321);
nand U14572 (N_14572,N_14104,N_13917);
or U14573 (N_14573,N_13937,N_14053);
nor U14574 (N_14574,N_14251,N_14203);
nand U14575 (N_14575,N_14258,N_13867);
nand U14576 (N_14576,N_13800,N_14061);
xor U14577 (N_14577,N_14254,N_14395);
nor U14578 (N_14578,N_13895,N_13952);
nor U14579 (N_14579,N_14378,N_13814);
or U14580 (N_14580,N_13921,N_14363);
nand U14581 (N_14581,N_13945,N_14011);
and U14582 (N_14582,N_14085,N_13967);
and U14583 (N_14583,N_14201,N_14127);
or U14584 (N_14584,N_14113,N_14030);
and U14585 (N_14585,N_14128,N_14242);
and U14586 (N_14586,N_13959,N_14347);
or U14587 (N_14587,N_14114,N_13832);
or U14588 (N_14588,N_14224,N_14290);
nand U14589 (N_14589,N_14359,N_14333);
nor U14590 (N_14590,N_14148,N_14003);
nand U14591 (N_14591,N_14328,N_14331);
and U14592 (N_14592,N_13925,N_14207);
and U14593 (N_14593,N_14052,N_13849);
or U14594 (N_14594,N_14302,N_13956);
xor U14595 (N_14595,N_14083,N_14278);
nand U14596 (N_14596,N_14348,N_13940);
nor U14597 (N_14597,N_14188,N_14068);
nand U14598 (N_14598,N_13807,N_13854);
and U14599 (N_14599,N_14204,N_13993);
and U14600 (N_14600,N_13896,N_13966);
nand U14601 (N_14601,N_14084,N_13886);
and U14602 (N_14602,N_14162,N_14196);
nor U14603 (N_14603,N_14308,N_13810);
nor U14604 (N_14604,N_14337,N_13979);
xnor U14605 (N_14605,N_14012,N_13941);
and U14606 (N_14606,N_14374,N_13893);
or U14607 (N_14607,N_14239,N_14274);
or U14608 (N_14608,N_14324,N_14373);
and U14609 (N_14609,N_13877,N_14393);
nor U14610 (N_14610,N_13902,N_14046);
and U14611 (N_14611,N_14159,N_14010);
nand U14612 (N_14612,N_13990,N_14043);
and U14613 (N_14613,N_14349,N_14072);
xnor U14614 (N_14614,N_13906,N_14339);
nor U14615 (N_14615,N_13823,N_13989);
and U14616 (N_14616,N_14033,N_14108);
and U14617 (N_14617,N_14022,N_14319);
xor U14618 (N_14618,N_13837,N_14282);
nor U14619 (N_14619,N_14269,N_14312);
xnor U14620 (N_14620,N_14215,N_13802);
or U14621 (N_14621,N_13889,N_14253);
nor U14622 (N_14622,N_14311,N_14074);
nand U14623 (N_14623,N_13922,N_14054);
nor U14624 (N_14624,N_14115,N_14288);
or U14625 (N_14625,N_14157,N_14335);
or U14626 (N_14626,N_13982,N_14153);
or U14627 (N_14627,N_14096,N_14040);
xnor U14628 (N_14628,N_14300,N_13856);
or U14629 (N_14629,N_14121,N_13972);
nor U14630 (N_14630,N_14198,N_13824);
or U14631 (N_14631,N_13904,N_14232);
nor U14632 (N_14632,N_14044,N_14142);
nor U14633 (N_14633,N_14244,N_13936);
nand U14634 (N_14634,N_13926,N_14219);
or U14635 (N_14635,N_13841,N_14289);
nand U14636 (N_14636,N_14167,N_13955);
and U14637 (N_14637,N_14292,N_14267);
or U14638 (N_14638,N_14377,N_14024);
or U14639 (N_14639,N_14134,N_14186);
xor U14640 (N_14640,N_13845,N_13839);
nand U14641 (N_14641,N_14171,N_13985);
xnor U14642 (N_14642,N_14285,N_14305);
or U14643 (N_14643,N_13855,N_13894);
nand U14644 (N_14644,N_13983,N_13975);
xor U14645 (N_14645,N_13914,N_14192);
nand U14646 (N_14646,N_14336,N_13887);
xnor U14647 (N_14647,N_14281,N_13825);
and U14648 (N_14648,N_14093,N_14268);
xnor U14649 (N_14649,N_13827,N_13897);
or U14650 (N_14650,N_14310,N_14293);
nor U14651 (N_14651,N_14180,N_13803);
nor U14652 (N_14652,N_14154,N_14001);
and U14653 (N_14653,N_13874,N_14240);
nor U14654 (N_14654,N_14138,N_14036);
nand U14655 (N_14655,N_14264,N_14301);
xnor U14656 (N_14656,N_14020,N_14172);
nand U14657 (N_14657,N_13973,N_14330);
nor U14658 (N_14658,N_14082,N_14141);
xor U14659 (N_14659,N_13939,N_13929);
and U14660 (N_14660,N_14318,N_14187);
xor U14661 (N_14661,N_13857,N_14048);
nor U14662 (N_14662,N_13930,N_14340);
or U14663 (N_14663,N_13911,N_14295);
or U14664 (N_14664,N_13861,N_14051);
or U14665 (N_14665,N_14313,N_14149);
or U14666 (N_14666,N_14358,N_13850);
and U14667 (N_14667,N_14135,N_14029);
and U14668 (N_14668,N_14182,N_14379);
nor U14669 (N_14669,N_14120,N_13884);
or U14670 (N_14670,N_14086,N_14222);
xnor U14671 (N_14671,N_14398,N_13846);
nor U14672 (N_14672,N_13899,N_13995);
nand U14673 (N_14673,N_13978,N_13909);
or U14674 (N_14674,N_13977,N_13991);
nor U14675 (N_14675,N_14376,N_14034);
and U14676 (N_14676,N_14394,N_14332);
xnor U14677 (N_14677,N_14067,N_14021);
or U14678 (N_14678,N_14208,N_14366);
or U14679 (N_14679,N_13820,N_13947);
and U14680 (N_14680,N_14031,N_14200);
nand U14681 (N_14681,N_14397,N_13866);
xor U14682 (N_14682,N_14338,N_14228);
nor U14683 (N_14683,N_13819,N_14199);
nor U14684 (N_14684,N_13970,N_14317);
nand U14685 (N_14685,N_13860,N_13932);
xnor U14686 (N_14686,N_14140,N_13957);
nand U14687 (N_14687,N_14060,N_14129);
or U14688 (N_14688,N_14315,N_14183);
or U14689 (N_14689,N_14078,N_13844);
nor U14690 (N_14690,N_13876,N_14178);
or U14691 (N_14691,N_14005,N_14130);
nand U14692 (N_14692,N_14193,N_14123);
and U14693 (N_14693,N_14360,N_13817);
nor U14694 (N_14694,N_14245,N_14095);
and U14695 (N_14695,N_14097,N_13822);
nand U14696 (N_14696,N_14283,N_14323);
nor U14697 (N_14697,N_13804,N_13851);
xor U14698 (N_14698,N_14079,N_14014);
nand U14699 (N_14699,N_13960,N_13863);
nor U14700 (N_14700,N_14007,N_13890);
and U14701 (N_14701,N_14359,N_14056);
xor U14702 (N_14702,N_13835,N_14082);
and U14703 (N_14703,N_14070,N_14167);
nand U14704 (N_14704,N_14391,N_13874);
xnor U14705 (N_14705,N_14164,N_14398);
xnor U14706 (N_14706,N_14061,N_14141);
xor U14707 (N_14707,N_13954,N_14204);
xnor U14708 (N_14708,N_14201,N_13929);
and U14709 (N_14709,N_13917,N_13826);
xor U14710 (N_14710,N_14191,N_13918);
xnor U14711 (N_14711,N_14211,N_14003);
and U14712 (N_14712,N_13878,N_14381);
nor U14713 (N_14713,N_13808,N_13865);
xnor U14714 (N_14714,N_14333,N_13936);
and U14715 (N_14715,N_14029,N_14018);
nor U14716 (N_14716,N_13893,N_14049);
xor U14717 (N_14717,N_14384,N_13850);
or U14718 (N_14718,N_14144,N_14318);
nor U14719 (N_14719,N_13997,N_14047);
and U14720 (N_14720,N_13928,N_14159);
nor U14721 (N_14721,N_13925,N_14040);
or U14722 (N_14722,N_14260,N_14043);
nor U14723 (N_14723,N_14097,N_14219);
nand U14724 (N_14724,N_13966,N_13993);
and U14725 (N_14725,N_14090,N_14150);
xor U14726 (N_14726,N_13881,N_14353);
nor U14727 (N_14727,N_14293,N_14183);
or U14728 (N_14728,N_14255,N_14215);
nor U14729 (N_14729,N_13930,N_13979);
xor U14730 (N_14730,N_14369,N_14185);
nor U14731 (N_14731,N_14044,N_14361);
or U14732 (N_14732,N_14120,N_14138);
nand U14733 (N_14733,N_13952,N_14124);
nand U14734 (N_14734,N_13867,N_14355);
xnor U14735 (N_14735,N_14157,N_13978);
and U14736 (N_14736,N_14355,N_14222);
xnor U14737 (N_14737,N_14220,N_13804);
nor U14738 (N_14738,N_14253,N_13844);
nor U14739 (N_14739,N_14221,N_13921);
nor U14740 (N_14740,N_14130,N_14184);
xnor U14741 (N_14741,N_14252,N_13921);
or U14742 (N_14742,N_14204,N_13941);
xor U14743 (N_14743,N_14049,N_14359);
nand U14744 (N_14744,N_14051,N_13920);
xnor U14745 (N_14745,N_14003,N_13898);
nor U14746 (N_14746,N_14092,N_13818);
or U14747 (N_14747,N_13862,N_14309);
nor U14748 (N_14748,N_13844,N_14226);
xnor U14749 (N_14749,N_14212,N_14214);
and U14750 (N_14750,N_14328,N_13802);
or U14751 (N_14751,N_13992,N_14083);
nor U14752 (N_14752,N_14347,N_14328);
or U14753 (N_14753,N_13917,N_14184);
nor U14754 (N_14754,N_14267,N_13865);
and U14755 (N_14755,N_14228,N_13822);
xnor U14756 (N_14756,N_14083,N_14336);
xnor U14757 (N_14757,N_14366,N_14111);
and U14758 (N_14758,N_14084,N_13843);
xor U14759 (N_14759,N_14349,N_13899);
and U14760 (N_14760,N_14330,N_13915);
xor U14761 (N_14761,N_14220,N_13920);
nand U14762 (N_14762,N_14313,N_13935);
nand U14763 (N_14763,N_14014,N_14335);
or U14764 (N_14764,N_14036,N_14217);
nor U14765 (N_14765,N_13973,N_14223);
nor U14766 (N_14766,N_14003,N_14057);
or U14767 (N_14767,N_13857,N_14078);
or U14768 (N_14768,N_13923,N_13862);
or U14769 (N_14769,N_14043,N_14024);
xor U14770 (N_14770,N_14395,N_14322);
and U14771 (N_14771,N_14285,N_13983);
or U14772 (N_14772,N_13967,N_14268);
or U14773 (N_14773,N_14091,N_14359);
nor U14774 (N_14774,N_13850,N_14260);
nand U14775 (N_14775,N_14263,N_14393);
nor U14776 (N_14776,N_13912,N_13997);
nor U14777 (N_14777,N_14232,N_13887);
xor U14778 (N_14778,N_14235,N_14118);
and U14779 (N_14779,N_14234,N_13838);
xor U14780 (N_14780,N_13879,N_14031);
or U14781 (N_14781,N_13809,N_14302);
nand U14782 (N_14782,N_13875,N_14340);
xnor U14783 (N_14783,N_14039,N_14170);
xor U14784 (N_14784,N_14081,N_14013);
nor U14785 (N_14785,N_14301,N_14344);
xor U14786 (N_14786,N_14288,N_14396);
nand U14787 (N_14787,N_13929,N_13902);
nand U14788 (N_14788,N_13992,N_14259);
xor U14789 (N_14789,N_13907,N_14235);
nand U14790 (N_14790,N_13804,N_14374);
or U14791 (N_14791,N_14178,N_14140);
xor U14792 (N_14792,N_13805,N_13861);
xor U14793 (N_14793,N_14058,N_14024);
nand U14794 (N_14794,N_14065,N_13953);
and U14795 (N_14795,N_14251,N_13852);
or U14796 (N_14796,N_14372,N_14381);
xnor U14797 (N_14797,N_14179,N_13941);
nor U14798 (N_14798,N_14009,N_14189);
xnor U14799 (N_14799,N_13974,N_13928);
xnor U14800 (N_14800,N_13992,N_14054);
and U14801 (N_14801,N_13818,N_14109);
nor U14802 (N_14802,N_14059,N_13995);
xnor U14803 (N_14803,N_14273,N_14180);
or U14804 (N_14804,N_14259,N_14053);
nor U14805 (N_14805,N_13815,N_14170);
nor U14806 (N_14806,N_14099,N_14287);
nor U14807 (N_14807,N_14181,N_14344);
nand U14808 (N_14808,N_13850,N_13895);
nor U14809 (N_14809,N_14172,N_13871);
or U14810 (N_14810,N_14348,N_14320);
and U14811 (N_14811,N_13837,N_14285);
nand U14812 (N_14812,N_14338,N_13948);
or U14813 (N_14813,N_14268,N_14099);
and U14814 (N_14814,N_14394,N_13818);
or U14815 (N_14815,N_14284,N_14147);
nand U14816 (N_14816,N_14249,N_14269);
nand U14817 (N_14817,N_13967,N_14187);
and U14818 (N_14818,N_13964,N_13953);
nor U14819 (N_14819,N_14057,N_14002);
or U14820 (N_14820,N_14264,N_14159);
and U14821 (N_14821,N_14328,N_14141);
nand U14822 (N_14822,N_13810,N_14326);
nor U14823 (N_14823,N_14000,N_14059);
xnor U14824 (N_14824,N_14253,N_13964);
or U14825 (N_14825,N_13895,N_14251);
nor U14826 (N_14826,N_13990,N_13931);
or U14827 (N_14827,N_14362,N_14076);
xor U14828 (N_14828,N_14105,N_14045);
xor U14829 (N_14829,N_13820,N_13933);
nor U14830 (N_14830,N_13928,N_14103);
xnor U14831 (N_14831,N_13903,N_14367);
nor U14832 (N_14832,N_13964,N_14351);
xnor U14833 (N_14833,N_14205,N_14102);
and U14834 (N_14834,N_13830,N_14136);
or U14835 (N_14835,N_14128,N_13815);
xor U14836 (N_14836,N_13913,N_14351);
or U14837 (N_14837,N_14174,N_14377);
and U14838 (N_14838,N_13883,N_14125);
and U14839 (N_14839,N_13900,N_13931);
nand U14840 (N_14840,N_13823,N_14386);
or U14841 (N_14841,N_13817,N_14307);
nor U14842 (N_14842,N_14004,N_14338);
nand U14843 (N_14843,N_13917,N_14308);
nor U14844 (N_14844,N_14169,N_14226);
and U14845 (N_14845,N_14062,N_14296);
and U14846 (N_14846,N_14118,N_14230);
or U14847 (N_14847,N_13857,N_14337);
nor U14848 (N_14848,N_13845,N_13876);
xnor U14849 (N_14849,N_13933,N_14002);
nor U14850 (N_14850,N_14089,N_13931);
and U14851 (N_14851,N_14141,N_13998);
xor U14852 (N_14852,N_13976,N_14148);
nor U14853 (N_14853,N_14352,N_14205);
or U14854 (N_14854,N_13900,N_14032);
xnor U14855 (N_14855,N_14020,N_14236);
and U14856 (N_14856,N_14078,N_13836);
nand U14857 (N_14857,N_13983,N_13989);
nand U14858 (N_14858,N_13939,N_14163);
xor U14859 (N_14859,N_14149,N_14245);
nand U14860 (N_14860,N_14167,N_13915);
nand U14861 (N_14861,N_13993,N_14321);
xor U14862 (N_14862,N_14183,N_14218);
and U14863 (N_14863,N_14122,N_14303);
and U14864 (N_14864,N_13818,N_14212);
nand U14865 (N_14865,N_14134,N_13805);
nor U14866 (N_14866,N_13862,N_13907);
nor U14867 (N_14867,N_13879,N_13935);
nand U14868 (N_14868,N_14097,N_13934);
xor U14869 (N_14869,N_13908,N_14101);
nand U14870 (N_14870,N_14257,N_13904);
nor U14871 (N_14871,N_14249,N_13991);
xor U14872 (N_14872,N_14056,N_13975);
xnor U14873 (N_14873,N_14214,N_14229);
and U14874 (N_14874,N_14358,N_13807);
or U14875 (N_14875,N_14340,N_14270);
xnor U14876 (N_14876,N_13844,N_14162);
and U14877 (N_14877,N_14223,N_14142);
nand U14878 (N_14878,N_14336,N_14094);
or U14879 (N_14879,N_14033,N_14329);
or U14880 (N_14880,N_14100,N_13977);
or U14881 (N_14881,N_14030,N_14088);
xnor U14882 (N_14882,N_14323,N_14059);
or U14883 (N_14883,N_14283,N_14131);
or U14884 (N_14884,N_14015,N_14388);
or U14885 (N_14885,N_13998,N_13988);
and U14886 (N_14886,N_13942,N_14392);
or U14887 (N_14887,N_14063,N_14236);
nor U14888 (N_14888,N_14120,N_14398);
and U14889 (N_14889,N_14056,N_13930);
nor U14890 (N_14890,N_13941,N_14143);
or U14891 (N_14891,N_13992,N_14072);
nor U14892 (N_14892,N_13941,N_14357);
or U14893 (N_14893,N_14052,N_13862);
and U14894 (N_14894,N_13849,N_14064);
or U14895 (N_14895,N_14196,N_13870);
and U14896 (N_14896,N_14168,N_14066);
nor U14897 (N_14897,N_14041,N_14098);
nand U14898 (N_14898,N_13809,N_14092);
nand U14899 (N_14899,N_14134,N_14335);
and U14900 (N_14900,N_13928,N_14151);
and U14901 (N_14901,N_13979,N_13927);
or U14902 (N_14902,N_14170,N_14350);
xnor U14903 (N_14903,N_13891,N_13938);
xnor U14904 (N_14904,N_13996,N_14066);
nand U14905 (N_14905,N_14113,N_13943);
nand U14906 (N_14906,N_14269,N_14262);
and U14907 (N_14907,N_14020,N_14251);
nor U14908 (N_14908,N_13934,N_14248);
xor U14909 (N_14909,N_14097,N_14060);
nor U14910 (N_14910,N_14312,N_13805);
xor U14911 (N_14911,N_13835,N_14087);
and U14912 (N_14912,N_14097,N_14019);
or U14913 (N_14913,N_13959,N_13897);
nor U14914 (N_14914,N_14391,N_14186);
xor U14915 (N_14915,N_14041,N_13917);
xnor U14916 (N_14916,N_14103,N_13964);
nand U14917 (N_14917,N_13980,N_14067);
and U14918 (N_14918,N_14195,N_14107);
and U14919 (N_14919,N_13902,N_14392);
nor U14920 (N_14920,N_14295,N_14162);
or U14921 (N_14921,N_13846,N_14354);
xnor U14922 (N_14922,N_14240,N_13984);
or U14923 (N_14923,N_14211,N_14226);
nor U14924 (N_14924,N_13836,N_14304);
and U14925 (N_14925,N_13864,N_13915);
nand U14926 (N_14926,N_13980,N_14124);
or U14927 (N_14927,N_14210,N_14220);
nand U14928 (N_14928,N_14120,N_14332);
nand U14929 (N_14929,N_14127,N_13976);
xor U14930 (N_14930,N_13967,N_14366);
nor U14931 (N_14931,N_13991,N_13874);
and U14932 (N_14932,N_13962,N_14139);
or U14933 (N_14933,N_14243,N_13983);
nand U14934 (N_14934,N_13998,N_13888);
xor U14935 (N_14935,N_14297,N_14327);
and U14936 (N_14936,N_14279,N_13880);
nor U14937 (N_14937,N_14062,N_14331);
or U14938 (N_14938,N_14310,N_13812);
or U14939 (N_14939,N_14063,N_14346);
and U14940 (N_14940,N_13880,N_14275);
xor U14941 (N_14941,N_14295,N_14276);
xor U14942 (N_14942,N_14278,N_14164);
or U14943 (N_14943,N_14052,N_13990);
nand U14944 (N_14944,N_14068,N_13803);
and U14945 (N_14945,N_14380,N_14078);
nor U14946 (N_14946,N_13972,N_13921);
xnor U14947 (N_14947,N_14076,N_13913);
nand U14948 (N_14948,N_13980,N_14288);
nand U14949 (N_14949,N_13816,N_14267);
nor U14950 (N_14950,N_13870,N_14072);
nor U14951 (N_14951,N_14178,N_13850);
or U14952 (N_14952,N_14215,N_13912);
nor U14953 (N_14953,N_14390,N_14288);
xor U14954 (N_14954,N_13860,N_13903);
nor U14955 (N_14955,N_14059,N_14126);
nor U14956 (N_14956,N_14162,N_13895);
and U14957 (N_14957,N_13826,N_14307);
or U14958 (N_14958,N_14050,N_14215);
nand U14959 (N_14959,N_14345,N_13876);
and U14960 (N_14960,N_14125,N_13953);
nor U14961 (N_14961,N_13951,N_14352);
nand U14962 (N_14962,N_13868,N_13834);
xnor U14963 (N_14963,N_14053,N_14301);
nand U14964 (N_14964,N_14192,N_14321);
nor U14965 (N_14965,N_14176,N_14052);
nand U14966 (N_14966,N_14366,N_14380);
and U14967 (N_14967,N_14245,N_14195);
or U14968 (N_14968,N_14090,N_13839);
or U14969 (N_14969,N_13883,N_14245);
xnor U14970 (N_14970,N_13935,N_14366);
or U14971 (N_14971,N_13945,N_14221);
nand U14972 (N_14972,N_14139,N_13943);
nor U14973 (N_14973,N_13811,N_13878);
and U14974 (N_14974,N_14111,N_13953);
xnor U14975 (N_14975,N_14282,N_14398);
and U14976 (N_14976,N_13832,N_14116);
xnor U14977 (N_14977,N_13894,N_14399);
or U14978 (N_14978,N_13807,N_14379);
nor U14979 (N_14979,N_14397,N_14086);
nand U14980 (N_14980,N_13842,N_13961);
nor U14981 (N_14981,N_14343,N_14214);
or U14982 (N_14982,N_14203,N_14243);
or U14983 (N_14983,N_14171,N_14168);
and U14984 (N_14984,N_14205,N_13987);
or U14985 (N_14985,N_13986,N_14297);
nor U14986 (N_14986,N_14013,N_14184);
nand U14987 (N_14987,N_14073,N_14205);
or U14988 (N_14988,N_14298,N_13862);
nand U14989 (N_14989,N_14022,N_14137);
nand U14990 (N_14990,N_14178,N_14393);
nand U14991 (N_14991,N_14056,N_14276);
or U14992 (N_14992,N_14118,N_14262);
xnor U14993 (N_14993,N_13965,N_14295);
and U14994 (N_14994,N_14117,N_14309);
nand U14995 (N_14995,N_14218,N_14311);
nand U14996 (N_14996,N_14072,N_13848);
and U14997 (N_14997,N_13923,N_14186);
nor U14998 (N_14998,N_14240,N_14367);
nand U14999 (N_14999,N_14215,N_13866);
or U15000 (N_15000,N_14449,N_14803);
nor U15001 (N_15001,N_14822,N_14664);
and U15002 (N_15002,N_14765,N_14855);
nor U15003 (N_15003,N_14938,N_14888);
nor U15004 (N_15004,N_14998,N_14617);
nor U15005 (N_15005,N_14984,N_14798);
and U15006 (N_15006,N_14643,N_14770);
or U15007 (N_15007,N_14440,N_14678);
nor U15008 (N_15008,N_14940,N_14553);
xor U15009 (N_15009,N_14808,N_14978);
xnor U15010 (N_15010,N_14972,N_14936);
or U15011 (N_15011,N_14407,N_14791);
xnor U15012 (N_15012,N_14996,N_14575);
nor U15013 (N_15013,N_14868,N_14467);
xnor U15014 (N_15014,N_14403,N_14797);
nand U15015 (N_15015,N_14919,N_14827);
nor U15016 (N_15016,N_14691,N_14559);
xnor U15017 (N_15017,N_14437,N_14489);
nand U15018 (N_15018,N_14739,N_14472);
xnor U15019 (N_15019,N_14762,N_14928);
or U15020 (N_15020,N_14433,N_14478);
xnor U15021 (N_15021,N_14723,N_14953);
nor U15022 (N_15022,N_14698,N_14991);
nor U15023 (N_15023,N_14790,N_14496);
nand U15024 (N_15024,N_14659,N_14952);
or U15025 (N_15025,N_14509,N_14893);
nor U15026 (N_15026,N_14572,N_14750);
or U15027 (N_15027,N_14732,N_14687);
nand U15028 (N_15028,N_14843,N_14986);
nor U15029 (N_15029,N_14767,N_14902);
or U15030 (N_15030,N_14474,N_14987);
nor U15031 (N_15031,N_14684,N_14892);
and U15032 (N_15032,N_14840,N_14673);
nor U15033 (N_15033,N_14849,N_14525);
nand U15034 (N_15034,N_14679,N_14645);
or U15035 (N_15035,N_14626,N_14547);
nor U15036 (N_15036,N_14568,N_14555);
and U15037 (N_15037,N_14900,N_14789);
nor U15038 (N_15038,N_14431,N_14445);
nor U15039 (N_15039,N_14700,N_14966);
xor U15040 (N_15040,N_14728,N_14704);
nor U15041 (N_15041,N_14740,N_14523);
and U15042 (N_15042,N_14794,N_14578);
nand U15043 (N_15043,N_14482,N_14420);
or U15044 (N_15044,N_14957,N_14557);
nor U15045 (N_15045,N_14944,N_14533);
xor U15046 (N_15046,N_14484,N_14453);
nor U15047 (N_15047,N_14622,N_14677);
xor U15048 (N_15048,N_14963,N_14712);
xnor U15049 (N_15049,N_14571,N_14722);
or U15050 (N_15050,N_14534,N_14701);
nor U15051 (N_15051,N_14899,N_14425);
nor U15052 (N_15052,N_14551,N_14585);
nor U15053 (N_15053,N_14414,N_14895);
nand U15054 (N_15054,N_14951,N_14869);
or U15055 (N_15055,N_14662,N_14683);
nand U15056 (N_15056,N_14707,N_14644);
nand U15057 (N_15057,N_14753,N_14625);
nand U15058 (N_15058,N_14427,N_14805);
nor U15059 (N_15059,N_14675,N_14799);
xor U15060 (N_15060,N_14587,N_14468);
or U15061 (N_15061,N_14956,N_14415);
xnor U15062 (N_15062,N_14490,N_14973);
and U15063 (N_15063,N_14458,N_14749);
nand U15064 (N_15064,N_14716,N_14635);
nor U15065 (N_15065,N_14937,N_14760);
and U15066 (N_15066,N_14444,N_14516);
nor U15067 (N_15067,N_14714,N_14878);
nand U15068 (N_15068,N_14579,N_14730);
xor U15069 (N_15069,N_14593,N_14428);
nor U15070 (N_15070,N_14844,N_14550);
nor U15071 (N_15071,N_14810,N_14495);
nor U15072 (N_15072,N_14763,N_14573);
nor U15073 (N_15073,N_14402,N_14649);
nor U15074 (N_15074,N_14608,N_14686);
and U15075 (N_15075,N_14564,N_14529);
and U15076 (N_15076,N_14945,N_14512);
xor U15077 (N_15077,N_14419,N_14884);
nand U15078 (N_15078,N_14904,N_14846);
nor U15079 (N_15079,N_14775,N_14929);
and U15080 (N_15080,N_14795,N_14618);
nor U15081 (N_15081,N_14503,N_14852);
nand U15082 (N_15082,N_14526,N_14779);
nand U15083 (N_15083,N_14964,N_14519);
xor U15084 (N_15084,N_14586,N_14657);
or U15085 (N_15085,N_14486,N_14909);
nor U15086 (N_15086,N_14977,N_14695);
and U15087 (N_15087,N_14736,N_14982);
and U15088 (N_15088,N_14432,N_14501);
and U15089 (N_15089,N_14784,N_14513);
nand U15090 (N_15090,N_14653,N_14514);
or U15091 (N_15091,N_14702,N_14850);
nor U15092 (N_15092,N_14515,N_14861);
xor U15093 (N_15093,N_14755,N_14439);
nor U15094 (N_15094,N_14706,N_14450);
and U15095 (N_15095,N_14821,N_14914);
nand U15096 (N_15096,N_14518,N_14989);
or U15097 (N_15097,N_14521,N_14621);
nand U15098 (N_15098,N_14615,N_14804);
xnor U15099 (N_15099,N_14668,N_14833);
nor U15100 (N_15100,N_14494,N_14674);
nor U15101 (N_15101,N_14891,N_14429);
xnor U15102 (N_15102,N_14567,N_14883);
or U15103 (N_15103,N_14435,N_14412);
nor U15104 (N_15104,N_14520,N_14746);
and U15105 (N_15105,N_14882,N_14713);
xnor U15106 (N_15106,N_14502,N_14807);
nand U15107 (N_15107,N_14866,N_14655);
nor U15108 (N_15108,N_14970,N_14639);
nand U15109 (N_15109,N_14881,N_14464);
nor U15110 (N_15110,N_14811,N_14661);
and U15111 (N_15111,N_14614,N_14967);
or U15112 (N_15112,N_14629,N_14766);
nand U15113 (N_15113,N_14491,N_14911);
and U15114 (N_15114,N_14461,N_14824);
nand U15115 (N_15115,N_14600,N_14851);
nor U15116 (N_15116,N_14934,N_14954);
and U15117 (N_15117,N_14656,N_14576);
or U15118 (N_15118,N_14873,N_14510);
nand U15119 (N_15119,N_14814,N_14566);
xor U15120 (N_15120,N_14733,N_14979);
or U15121 (N_15121,N_14499,N_14594);
nand U15122 (N_15122,N_14511,N_14837);
or U15123 (N_15123,N_14451,N_14436);
nand U15124 (N_15124,N_14917,N_14738);
xnor U15125 (N_15125,N_14829,N_14876);
and U15126 (N_15126,N_14652,N_14971);
or U15127 (N_15127,N_14492,N_14471);
nand U15128 (N_15128,N_14809,N_14853);
or U15129 (N_15129,N_14773,N_14935);
xnor U15130 (N_15130,N_14741,N_14806);
and U15131 (N_15131,N_14735,N_14574);
xor U15132 (N_15132,N_14719,N_14724);
nor U15133 (N_15133,N_14842,N_14565);
and U15134 (N_15134,N_14692,N_14693);
or U15135 (N_15135,N_14903,N_14825);
or U15136 (N_15136,N_14897,N_14624);
and U15137 (N_15137,N_14859,N_14898);
nand U15138 (N_15138,N_14581,N_14540);
and U15139 (N_15139,N_14932,N_14672);
and U15140 (N_15140,N_14705,N_14793);
or U15141 (N_15141,N_14430,N_14976);
and U15142 (N_15142,N_14930,N_14602);
or U15143 (N_15143,N_14856,N_14708);
nor U15144 (N_15144,N_14792,N_14950);
and U15145 (N_15145,N_14641,N_14820);
nand U15146 (N_15146,N_14865,N_14654);
nand U15147 (N_15147,N_14959,N_14623);
nand U15148 (N_15148,N_14682,N_14912);
nand U15149 (N_15149,N_14828,N_14737);
or U15150 (N_15150,N_14636,N_14549);
and U15151 (N_15151,N_14459,N_14637);
or U15152 (N_15152,N_14992,N_14696);
nand U15153 (N_15153,N_14670,N_14589);
and U15154 (N_15154,N_14962,N_14786);
nor U15155 (N_15155,N_14504,N_14556);
nand U15156 (N_15156,N_14596,N_14532);
xor U15157 (N_15157,N_14598,N_14465);
nor U15158 (N_15158,N_14812,N_14651);
nand U15159 (N_15159,N_14462,N_14665);
nor U15160 (N_15160,N_14421,N_14946);
nand U15161 (N_15161,N_14417,N_14631);
nand U15162 (N_15162,N_14539,N_14815);
xor U15163 (N_15163,N_14999,N_14880);
or U15164 (N_15164,N_14718,N_14839);
xnor U15165 (N_15165,N_14921,N_14648);
and U15166 (N_15166,N_14727,N_14569);
nand U15167 (N_15167,N_14703,N_14831);
xor U15168 (N_15168,N_14864,N_14841);
nand U15169 (N_15169,N_14500,N_14890);
and U15170 (N_15170,N_14874,N_14548);
nand U15171 (N_15171,N_14633,N_14942);
or U15172 (N_15172,N_14619,N_14601);
nand U15173 (N_15173,N_14894,N_14907);
nand U15174 (N_15174,N_14582,N_14993);
and U15175 (N_15175,N_14871,N_14506);
and U15176 (N_15176,N_14721,N_14910);
and U15177 (N_15177,N_14782,N_14801);
nor U15178 (N_15178,N_14463,N_14613);
xnor U15179 (N_15179,N_14546,N_14454);
or U15180 (N_15180,N_14406,N_14627);
and U15181 (N_15181,N_14667,N_14422);
and U15182 (N_15182,N_14413,N_14906);
and U15183 (N_15183,N_14642,N_14980);
or U15184 (N_15184,N_14689,N_14697);
xnor U15185 (N_15185,N_14616,N_14711);
or U15186 (N_15186,N_14537,N_14958);
or U15187 (N_15187,N_14400,N_14817);
or U15188 (N_15188,N_14694,N_14699);
xor U15189 (N_15189,N_14835,N_14922);
and U15190 (N_15190,N_14442,N_14452);
nand U15191 (N_15191,N_14778,N_14742);
nor U15192 (N_15192,N_14709,N_14577);
nor U15193 (N_15193,N_14836,N_14774);
and U15194 (N_15194,N_14542,N_14505);
and U15195 (N_15195,N_14558,N_14592);
nor U15196 (N_15196,N_14438,N_14983);
xnor U15197 (N_15197,N_14751,N_14923);
and U15198 (N_15198,N_14469,N_14638);
nand U15199 (N_15199,N_14776,N_14603);
and U15200 (N_15200,N_14780,N_14560);
and U15201 (N_15201,N_14816,N_14446);
and U15202 (N_15202,N_14720,N_14981);
nand U15203 (N_15203,N_14772,N_14787);
nor U15204 (N_15204,N_14796,N_14680);
xor U15205 (N_15205,N_14745,N_14920);
or U15206 (N_15206,N_14609,N_14524);
nand U15207 (N_15207,N_14771,N_14563);
nand U15208 (N_15208,N_14597,N_14676);
nand U15209 (N_15209,N_14470,N_14715);
and U15210 (N_15210,N_14990,N_14632);
xor U15211 (N_15211,N_14854,N_14498);
xnor U15212 (N_15212,N_14570,N_14647);
nor U15213 (N_15213,N_14456,N_14965);
nand U15214 (N_15214,N_14752,N_14931);
nand U15215 (N_15215,N_14493,N_14830);
or U15216 (N_15216,N_14819,N_14475);
nand U15217 (N_15217,N_14756,N_14480);
nor U15218 (N_15218,N_14630,N_14561);
nor U15219 (N_15219,N_14788,N_14848);
nor U15220 (N_15220,N_14584,N_14863);
xor U15221 (N_15221,N_14681,N_14860);
nand U15222 (N_15222,N_14757,N_14838);
nor U15223 (N_15223,N_14591,N_14595);
or U15224 (N_15224,N_14729,N_14604);
nor U15225 (N_15225,N_14401,N_14605);
nor U15226 (N_15226,N_14918,N_14535);
or U15227 (N_15227,N_14915,N_14974);
nand U15228 (N_15228,N_14877,N_14476);
xor U15229 (N_15229,N_14460,N_14426);
or U15230 (N_15230,N_14823,N_14447);
and U15231 (N_15231,N_14590,N_14896);
xor U15232 (N_15232,N_14663,N_14416);
nand U15233 (N_15233,N_14562,N_14457);
nor U15234 (N_15234,N_14671,N_14758);
and U15235 (N_15235,N_14466,N_14994);
and U15236 (N_15236,N_14487,N_14948);
and U15237 (N_15237,N_14405,N_14748);
nor U15238 (N_15238,N_14913,N_14800);
nand U15239 (N_15239,N_14410,N_14690);
nor U15240 (N_15240,N_14924,N_14725);
nor U15241 (N_15241,N_14734,N_14826);
xnor U15242 (N_15242,N_14646,N_14610);
or U15243 (N_15243,N_14947,N_14607);
and U15244 (N_15244,N_14988,N_14536);
or U15245 (N_15245,N_14606,N_14545);
nor U15246 (N_15246,N_14508,N_14634);
nor U15247 (N_15247,N_14640,N_14764);
nor U15248 (N_15248,N_14908,N_14813);
or U15249 (N_15249,N_14761,N_14879);
and U15250 (N_15250,N_14685,N_14481);
xor U15251 (N_15251,N_14527,N_14916);
nand U15252 (N_15252,N_14473,N_14969);
nand U15253 (N_15253,N_14961,N_14448);
or U15254 (N_15254,N_14862,N_14777);
xor U15255 (N_15255,N_14845,N_14483);
nor U15256 (N_15256,N_14411,N_14554);
nor U15257 (N_15257,N_14754,N_14522);
and U15258 (N_15258,N_14424,N_14620);
or U15259 (N_15259,N_14404,N_14477);
nor U15260 (N_15260,N_14768,N_14443);
xnor U15261 (N_15261,N_14531,N_14975);
and U15262 (N_15262,N_14669,N_14949);
or U15263 (N_15263,N_14517,N_14832);
or U15264 (N_15264,N_14886,N_14528);
xnor U15265 (N_15265,N_14901,N_14418);
and U15266 (N_15266,N_14802,N_14744);
nand U15267 (N_15267,N_14731,N_14423);
nand U15268 (N_15268,N_14926,N_14834);
xor U15269 (N_15269,N_14985,N_14857);
xnor U15270 (N_15270,N_14544,N_14485);
or U15271 (N_15271,N_14781,N_14943);
xnor U15272 (N_15272,N_14887,N_14783);
and U15273 (N_15273,N_14927,N_14960);
nor U15274 (N_15274,N_14688,N_14455);
and U15275 (N_15275,N_14541,N_14710);
nand U15276 (N_15276,N_14552,N_14612);
xnor U15277 (N_15277,N_14583,N_14726);
and U15278 (N_15278,N_14955,N_14660);
xnor U15279 (N_15279,N_14409,N_14905);
xnor U15280 (N_15280,N_14769,N_14408);
nor U15281 (N_15281,N_14611,N_14870);
xnor U15282 (N_15282,N_14867,N_14628);
nor U15283 (N_15283,N_14507,N_14650);
nand U15284 (N_15284,N_14747,N_14666);
nand U15285 (N_15285,N_14847,N_14543);
nand U15286 (N_15286,N_14939,N_14441);
and U15287 (N_15287,N_14658,N_14885);
or U15288 (N_15288,N_14933,N_14785);
nor U15289 (N_15289,N_14488,N_14743);
nand U15290 (N_15290,N_14858,N_14497);
nor U15291 (N_15291,N_14599,N_14889);
nand U15292 (N_15292,N_14997,N_14995);
and U15293 (N_15293,N_14530,N_14941);
nor U15294 (N_15294,N_14538,N_14818);
and U15295 (N_15295,N_14434,N_14479);
nor U15296 (N_15296,N_14968,N_14717);
or U15297 (N_15297,N_14588,N_14925);
nor U15298 (N_15298,N_14759,N_14875);
nand U15299 (N_15299,N_14872,N_14580);
nor U15300 (N_15300,N_14851,N_14785);
nor U15301 (N_15301,N_14665,N_14495);
nand U15302 (N_15302,N_14857,N_14752);
and U15303 (N_15303,N_14790,N_14829);
and U15304 (N_15304,N_14722,N_14775);
and U15305 (N_15305,N_14981,N_14758);
and U15306 (N_15306,N_14579,N_14914);
nand U15307 (N_15307,N_14767,N_14727);
xor U15308 (N_15308,N_14923,N_14975);
and U15309 (N_15309,N_14681,N_14535);
nor U15310 (N_15310,N_14748,N_14741);
nand U15311 (N_15311,N_14721,N_14580);
nor U15312 (N_15312,N_14800,N_14672);
or U15313 (N_15313,N_14682,N_14519);
or U15314 (N_15314,N_14857,N_14643);
and U15315 (N_15315,N_14809,N_14828);
xor U15316 (N_15316,N_14510,N_14742);
or U15317 (N_15317,N_14941,N_14505);
nor U15318 (N_15318,N_14899,N_14603);
or U15319 (N_15319,N_14599,N_14932);
or U15320 (N_15320,N_14450,N_14754);
nand U15321 (N_15321,N_14962,N_14535);
nor U15322 (N_15322,N_14620,N_14839);
and U15323 (N_15323,N_14898,N_14672);
nand U15324 (N_15324,N_14840,N_14821);
or U15325 (N_15325,N_14461,N_14781);
and U15326 (N_15326,N_14629,N_14638);
nor U15327 (N_15327,N_14477,N_14771);
xor U15328 (N_15328,N_14781,N_14476);
nor U15329 (N_15329,N_14628,N_14583);
nand U15330 (N_15330,N_14611,N_14675);
nor U15331 (N_15331,N_14819,N_14935);
and U15332 (N_15332,N_14430,N_14472);
and U15333 (N_15333,N_14965,N_14586);
xnor U15334 (N_15334,N_14908,N_14751);
nor U15335 (N_15335,N_14819,N_14553);
nor U15336 (N_15336,N_14519,N_14633);
and U15337 (N_15337,N_14796,N_14791);
nor U15338 (N_15338,N_14983,N_14897);
xnor U15339 (N_15339,N_14656,N_14769);
and U15340 (N_15340,N_14530,N_14560);
nor U15341 (N_15341,N_14573,N_14821);
and U15342 (N_15342,N_14556,N_14608);
or U15343 (N_15343,N_14576,N_14808);
nor U15344 (N_15344,N_14581,N_14887);
nand U15345 (N_15345,N_14638,N_14459);
or U15346 (N_15346,N_14873,N_14475);
or U15347 (N_15347,N_14655,N_14582);
and U15348 (N_15348,N_14430,N_14737);
or U15349 (N_15349,N_14627,N_14568);
or U15350 (N_15350,N_14468,N_14403);
nand U15351 (N_15351,N_14962,N_14636);
xor U15352 (N_15352,N_14917,N_14432);
nand U15353 (N_15353,N_14919,N_14793);
nor U15354 (N_15354,N_14952,N_14937);
or U15355 (N_15355,N_14537,N_14945);
and U15356 (N_15356,N_14525,N_14640);
or U15357 (N_15357,N_14771,N_14873);
nand U15358 (N_15358,N_14488,N_14796);
nor U15359 (N_15359,N_14881,N_14462);
xor U15360 (N_15360,N_14410,N_14964);
nor U15361 (N_15361,N_14488,N_14808);
xnor U15362 (N_15362,N_14702,N_14460);
nor U15363 (N_15363,N_14432,N_14929);
and U15364 (N_15364,N_14689,N_14820);
and U15365 (N_15365,N_14556,N_14515);
nor U15366 (N_15366,N_14641,N_14460);
and U15367 (N_15367,N_14611,N_14678);
xor U15368 (N_15368,N_14767,N_14683);
xor U15369 (N_15369,N_14707,N_14425);
and U15370 (N_15370,N_14745,N_14513);
and U15371 (N_15371,N_14743,N_14668);
nand U15372 (N_15372,N_14696,N_14629);
nor U15373 (N_15373,N_14457,N_14407);
nor U15374 (N_15374,N_14514,N_14499);
xor U15375 (N_15375,N_14742,N_14726);
nor U15376 (N_15376,N_14409,N_14990);
nand U15377 (N_15377,N_14765,N_14482);
nor U15378 (N_15378,N_14988,N_14927);
or U15379 (N_15379,N_14535,N_14759);
or U15380 (N_15380,N_14796,N_14859);
xor U15381 (N_15381,N_14629,N_14994);
nor U15382 (N_15382,N_14738,N_14684);
nor U15383 (N_15383,N_14710,N_14540);
nor U15384 (N_15384,N_14457,N_14620);
xnor U15385 (N_15385,N_14638,N_14402);
or U15386 (N_15386,N_14819,N_14618);
xnor U15387 (N_15387,N_14565,N_14813);
nand U15388 (N_15388,N_14843,N_14516);
nand U15389 (N_15389,N_14734,N_14600);
nor U15390 (N_15390,N_14476,N_14943);
xnor U15391 (N_15391,N_14770,N_14905);
and U15392 (N_15392,N_14726,N_14776);
and U15393 (N_15393,N_14841,N_14416);
and U15394 (N_15394,N_14931,N_14514);
nand U15395 (N_15395,N_14944,N_14860);
xnor U15396 (N_15396,N_14933,N_14854);
nor U15397 (N_15397,N_14836,N_14956);
and U15398 (N_15398,N_14509,N_14991);
xnor U15399 (N_15399,N_14434,N_14549);
nand U15400 (N_15400,N_14841,N_14667);
or U15401 (N_15401,N_14979,N_14851);
nand U15402 (N_15402,N_14677,N_14828);
and U15403 (N_15403,N_14843,N_14959);
xnor U15404 (N_15404,N_14404,N_14610);
or U15405 (N_15405,N_14853,N_14988);
and U15406 (N_15406,N_14445,N_14691);
xor U15407 (N_15407,N_14441,N_14449);
and U15408 (N_15408,N_14735,N_14469);
nor U15409 (N_15409,N_14859,N_14992);
nor U15410 (N_15410,N_14432,N_14706);
nor U15411 (N_15411,N_14719,N_14994);
nand U15412 (N_15412,N_14493,N_14790);
or U15413 (N_15413,N_14414,N_14522);
nand U15414 (N_15414,N_14559,N_14532);
or U15415 (N_15415,N_14559,N_14720);
or U15416 (N_15416,N_14876,N_14668);
and U15417 (N_15417,N_14856,N_14674);
and U15418 (N_15418,N_14807,N_14463);
and U15419 (N_15419,N_14435,N_14733);
xor U15420 (N_15420,N_14428,N_14703);
and U15421 (N_15421,N_14725,N_14966);
nor U15422 (N_15422,N_14484,N_14732);
and U15423 (N_15423,N_14952,N_14877);
and U15424 (N_15424,N_14832,N_14565);
nor U15425 (N_15425,N_14770,N_14853);
xor U15426 (N_15426,N_14970,N_14424);
nand U15427 (N_15427,N_14941,N_14429);
and U15428 (N_15428,N_14483,N_14695);
and U15429 (N_15429,N_14791,N_14711);
or U15430 (N_15430,N_14451,N_14457);
nor U15431 (N_15431,N_14500,N_14745);
nor U15432 (N_15432,N_14895,N_14919);
or U15433 (N_15433,N_14975,N_14886);
nand U15434 (N_15434,N_14768,N_14855);
and U15435 (N_15435,N_14606,N_14884);
or U15436 (N_15436,N_14591,N_14810);
nand U15437 (N_15437,N_14426,N_14814);
nand U15438 (N_15438,N_14464,N_14933);
nor U15439 (N_15439,N_14786,N_14941);
or U15440 (N_15440,N_14543,N_14534);
xnor U15441 (N_15441,N_14440,N_14813);
nor U15442 (N_15442,N_14790,N_14436);
or U15443 (N_15443,N_14706,N_14637);
and U15444 (N_15444,N_14724,N_14806);
or U15445 (N_15445,N_14413,N_14596);
and U15446 (N_15446,N_14682,N_14626);
nor U15447 (N_15447,N_14693,N_14428);
nor U15448 (N_15448,N_14676,N_14787);
nand U15449 (N_15449,N_14559,N_14411);
or U15450 (N_15450,N_14824,N_14667);
or U15451 (N_15451,N_14740,N_14963);
nor U15452 (N_15452,N_14976,N_14935);
and U15453 (N_15453,N_14636,N_14458);
xnor U15454 (N_15454,N_14409,N_14747);
nand U15455 (N_15455,N_14800,N_14686);
or U15456 (N_15456,N_14507,N_14669);
nand U15457 (N_15457,N_14928,N_14719);
xnor U15458 (N_15458,N_14896,N_14630);
or U15459 (N_15459,N_14584,N_14628);
and U15460 (N_15460,N_14468,N_14681);
and U15461 (N_15461,N_14802,N_14830);
nor U15462 (N_15462,N_14533,N_14807);
and U15463 (N_15463,N_14740,N_14791);
nor U15464 (N_15464,N_14827,N_14898);
xnor U15465 (N_15465,N_14664,N_14418);
xor U15466 (N_15466,N_14417,N_14791);
and U15467 (N_15467,N_14677,N_14442);
nor U15468 (N_15468,N_14625,N_14633);
xor U15469 (N_15469,N_14471,N_14911);
xnor U15470 (N_15470,N_14724,N_14704);
nor U15471 (N_15471,N_14930,N_14754);
nand U15472 (N_15472,N_14660,N_14827);
and U15473 (N_15473,N_14837,N_14797);
nor U15474 (N_15474,N_14808,N_14672);
nor U15475 (N_15475,N_14667,N_14638);
nor U15476 (N_15476,N_14824,N_14453);
and U15477 (N_15477,N_14961,N_14716);
nand U15478 (N_15478,N_14419,N_14557);
nor U15479 (N_15479,N_14923,N_14659);
or U15480 (N_15480,N_14633,N_14523);
and U15481 (N_15481,N_14730,N_14501);
nand U15482 (N_15482,N_14568,N_14680);
and U15483 (N_15483,N_14701,N_14451);
xnor U15484 (N_15484,N_14832,N_14947);
xnor U15485 (N_15485,N_14786,N_14725);
xnor U15486 (N_15486,N_14438,N_14774);
and U15487 (N_15487,N_14480,N_14773);
xnor U15488 (N_15488,N_14716,N_14925);
nand U15489 (N_15489,N_14596,N_14564);
nor U15490 (N_15490,N_14590,N_14506);
and U15491 (N_15491,N_14806,N_14833);
nand U15492 (N_15492,N_14930,N_14545);
xnor U15493 (N_15493,N_14410,N_14955);
nand U15494 (N_15494,N_14401,N_14468);
nand U15495 (N_15495,N_14570,N_14484);
xor U15496 (N_15496,N_14968,N_14934);
and U15497 (N_15497,N_14908,N_14466);
and U15498 (N_15498,N_14668,N_14594);
or U15499 (N_15499,N_14598,N_14872);
and U15500 (N_15500,N_14602,N_14744);
xor U15501 (N_15501,N_14967,N_14945);
and U15502 (N_15502,N_14440,N_14418);
or U15503 (N_15503,N_14851,N_14558);
or U15504 (N_15504,N_14647,N_14859);
or U15505 (N_15505,N_14922,N_14636);
xor U15506 (N_15506,N_14910,N_14865);
xor U15507 (N_15507,N_14615,N_14433);
and U15508 (N_15508,N_14779,N_14592);
or U15509 (N_15509,N_14408,N_14639);
and U15510 (N_15510,N_14414,N_14907);
nand U15511 (N_15511,N_14710,N_14934);
nor U15512 (N_15512,N_14774,N_14865);
nor U15513 (N_15513,N_14734,N_14409);
nor U15514 (N_15514,N_14661,N_14923);
or U15515 (N_15515,N_14489,N_14559);
nand U15516 (N_15516,N_14417,N_14686);
or U15517 (N_15517,N_14766,N_14578);
nor U15518 (N_15518,N_14734,N_14578);
nand U15519 (N_15519,N_14596,N_14785);
nor U15520 (N_15520,N_14925,N_14684);
or U15521 (N_15521,N_14998,N_14878);
nand U15522 (N_15522,N_14614,N_14706);
nor U15523 (N_15523,N_14661,N_14480);
xnor U15524 (N_15524,N_14624,N_14925);
xor U15525 (N_15525,N_14461,N_14432);
xor U15526 (N_15526,N_14428,N_14937);
nor U15527 (N_15527,N_14500,N_14822);
or U15528 (N_15528,N_14572,N_14991);
or U15529 (N_15529,N_14560,N_14619);
and U15530 (N_15530,N_14461,N_14917);
and U15531 (N_15531,N_14863,N_14574);
xnor U15532 (N_15532,N_14910,N_14961);
nor U15533 (N_15533,N_14433,N_14903);
nor U15534 (N_15534,N_14974,N_14943);
or U15535 (N_15535,N_14976,N_14534);
or U15536 (N_15536,N_14463,N_14544);
or U15537 (N_15537,N_14801,N_14430);
nor U15538 (N_15538,N_14715,N_14974);
or U15539 (N_15539,N_14868,N_14826);
nand U15540 (N_15540,N_14764,N_14952);
xnor U15541 (N_15541,N_14750,N_14657);
xor U15542 (N_15542,N_14831,N_14962);
xor U15543 (N_15543,N_14930,N_14787);
nand U15544 (N_15544,N_14993,N_14440);
xor U15545 (N_15545,N_14802,N_14908);
or U15546 (N_15546,N_14582,N_14665);
xnor U15547 (N_15547,N_14408,N_14531);
xor U15548 (N_15548,N_14466,N_14434);
or U15549 (N_15549,N_14628,N_14744);
nand U15550 (N_15550,N_14637,N_14683);
or U15551 (N_15551,N_14910,N_14790);
or U15552 (N_15552,N_14952,N_14582);
nand U15553 (N_15553,N_14406,N_14423);
and U15554 (N_15554,N_14730,N_14490);
or U15555 (N_15555,N_14507,N_14978);
or U15556 (N_15556,N_14829,N_14856);
nor U15557 (N_15557,N_14710,N_14954);
xor U15558 (N_15558,N_14770,N_14844);
xnor U15559 (N_15559,N_14542,N_14570);
nand U15560 (N_15560,N_14833,N_14651);
nand U15561 (N_15561,N_14860,N_14871);
and U15562 (N_15562,N_14489,N_14775);
or U15563 (N_15563,N_14937,N_14827);
nand U15564 (N_15564,N_14933,N_14569);
xnor U15565 (N_15565,N_14712,N_14949);
nand U15566 (N_15566,N_14984,N_14941);
or U15567 (N_15567,N_14818,N_14434);
nor U15568 (N_15568,N_14983,N_14598);
nand U15569 (N_15569,N_14935,N_14652);
and U15570 (N_15570,N_14968,N_14962);
nand U15571 (N_15571,N_14512,N_14796);
nand U15572 (N_15572,N_14409,N_14539);
xor U15573 (N_15573,N_14748,N_14910);
nor U15574 (N_15574,N_14900,N_14977);
xor U15575 (N_15575,N_14543,N_14530);
nor U15576 (N_15576,N_14463,N_14840);
and U15577 (N_15577,N_14686,N_14555);
and U15578 (N_15578,N_14551,N_14540);
nor U15579 (N_15579,N_14797,N_14890);
or U15580 (N_15580,N_14831,N_14774);
nor U15581 (N_15581,N_14904,N_14719);
nand U15582 (N_15582,N_14688,N_14510);
and U15583 (N_15583,N_14650,N_14488);
and U15584 (N_15584,N_14815,N_14711);
and U15585 (N_15585,N_14590,N_14470);
and U15586 (N_15586,N_14799,N_14635);
xor U15587 (N_15587,N_14706,N_14653);
and U15588 (N_15588,N_14800,N_14523);
or U15589 (N_15589,N_14432,N_14760);
nor U15590 (N_15590,N_14469,N_14819);
xnor U15591 (N_15591,N_14803,N_14467);
nand U15592 (N_15592,N_14984,N_14580);
nand U15593 (N_15593,N_14673,N_14767);
xor U15594 (N_15594,N_14952,N_14493);
nand U15595 (N_15595,N_14492,N_14587);
and U15596 (N_15596,N_14863,N_14569);
nand U15597 (N_15597,N_14659,N_14670);
or U15598 (N_15598,N_14829,N_14808);
xnor U15599 (N_15599,N_14831,N_14866);
and U15600 (N_15600,N_15532,N_15555);
nand U15601 (N_15601,N_15212,N_15383);
nor U15602 (N_15602,N_15045,N_15023);
nand U15603 (N_15603,N_15021,N_15449);
and U15604 (N_15604,N_15127,N_15140);
and U15605 (N_15605,N_15432,N_15492);
and U15606 (N_15606,N_15415,N_15228);
or U15607 (N_15607,N_15149,N_15113);
and U15608 (N_15608,N_15302,N_15009);
nand U15609 (N_15609,N_15597,N_15102);
and U15610 (N_15610,N_15453,N_15423);
or U15611 (N_15611,N_15067,N_15001);
nand U15612 (N_15612,N_15184,N_15134);
nor U15613 (N_15613,N_15268,N_15549);
and U15614 (N_15614,N_15471,N_15482);
xnor U15615 (N_15615,N_15494,N_15233);
nand U15616 (N_15616,N_15565,N_15361);
nor U15617 (N_15617,N_15554,N_15217);
nor U15618 (N_15618,N_15108,N_15066);
nand U15619 (N_15619,N_15396,N_15318);
nand U15620 (N_15620,N_15427,N_15089);
nor U15621 (N_15621,N_15497,N_15296);
or U15622 (N_15622,N_15278,N_15419);
or U15623 (N_15623,N_15172,N_15343);
xor U15624 (N_15624,N_15050,N_15579);
xnor U15625 (N_15625,N_15177,N_15095);
xor U15626 (N_15626,N_15496,N_15412);
xnor U15627 (N_15627,N_15411,N_15219);
or U15628 (N_15628,N_15099,N_15539);
xnor U15629 (N_15629,N_15114,N_15012);
nor U15630 (N_15630,N_15020,N_15235);
nand U15631 (N_15631,N_15145,N_15488);
or U15632 (N_15632,N_15522,N_15298);
and U15633 (N_15633,N_15578,N_15402);
xnor U15634 (N_15634,N_15315,N_15205);
xnor U15635 (N_15635,N_15098,N_15271);
or U15636 (N_15636,N_15109,N_15175);
and U15637 (N_15637,N_15382,N_15336);
xor U15638 (N_15638,N_15292,N_15046);
and U15639 (N_15639,N_15509,N_15413);
nand U15640 (N_15640,N_15061,N_15064);
nor U15641 (N_15641,N_15056,N_15245);
or U15642 (N_15642,N_15055,N_15389);
nor U15643 (N_15643,N_15426,N_15470);
nand U15644 (N_15644,N_15520,N_15585);
or U15645 (N_15645,N_15297,N_15273);
and U15646 (N_15646,N_15444,N_15331);
nor U15647 (N_15647,N_15160,N_15232);
nand U15648 (N_15648,N_15270,N_15379);
xor U15649 (N_15649,N_15475,N_15407);
nand U15650 (N_15650,N_15211,N_15590);
or U15651 (N_15651,N_15198,N_15310);
xor U15652 (N_15652,N_15247,N_15133);
nand U15653 (N_15653,N_15169,N_15309);
xor U15654 (N_15654,N_15042,N_15370);
nor U15655 (N_15655,N_15596,N_15399);
xor U15656 (N_15656,N_15562,N_15158);
and U15657 (N_15657,N_15533,N_15529);
xnor U15658 (N_15658,N_15117,N_15484);
and U15659 (N_15659,N_15252,N_15199);
nand U15660 (N_15660,N_15346,N_15026);
and U15661 (N_15661,N_15107,N_15577);
xor U15662 (N_15662,N_15034,N_15527);
xnor U15663 (N_15663,N_15375,N_15485);
nand U15664 (N_15664,N_15225,N_15438);
and U15665 (N_15665,N_15393,N_15072);
xor U15666 (N_15666,N_15563,N_15025);
or U15667 (N_15667,N_15065,N_15478);
and U15668 (N_15668,N_15123,N_15434);
and U15669 (N_15669,N_15347,N_15377);
nand U15670 (N_15670,N_15448,N_15171);
nand U15671 (N_15671,N_15291,N_15147);
or U15672 (N_15672,N_15429,N_15017);
nand U15673 (N_15673,N_15401,N_15457);
and U15674 (N_15674,N_15598,N_15337);
nand U15675 (N_15675,N_15499,N_15155);
or U15676 (N_15676,N_15060,N_15080);
nand U15677 (N_15677,N_15358,N_15242);
nand U15678 (N_15678,N_15112,N_15222);
nor U15679 (N_15679,N_15541,N_15283);
nor U15680 (N_15680,N_15131,N_15077);
nor U15681 (N_15681,N_15557,N_15576);
nor U15682 (N_15682,N_15373,N_15574);
nand U15683 (N_15683,N_15092,N_15194);
nor U15684 (N_15684,N_15435,N_15048);
or U15685 (N_15685,N_15091,N_15011);
nand U15686 (N_15686,N_15150,N_15180);
or U15687 (N_15687,N_15129,N_15463);
or U15688 (N_15688,N_15403,N_15197);
xnor U15689 (N_15689,N_15352,N_15263);
and U15690 (N_15690,N_15459,N_15581);
xnor U15691 (N_15691,N_15570,N_15404);
nand U15692 (N_15692,N_15290,N_15493);
xor U15693 (N_15693,N_15076,N_15322);
nor U15694 (N_15694,N_15575,N_15256);
nor U15695 (N_15695,N_15239,N_15257);
or U15696 (N_15696,N_15024,N_15231);
or U15697 (N_15697,N_15359,N_15474);
nor U15698 (N_15698,N_15130,N_15390);
nor U15699 (N_15699,N_15236,N_15335);
xnor U15700 (N_15700,N_15293,N_15552);
and U15701 (N_15701,N_15274,N_15540);
and U15702 (N_15702,N_15106,N_15097);
nand U15703 (N_15703,N_15450,N_15307);
or U15704 (N_15704,N_15489,N_15571);
nor U15705 (N_15705,N_15508,N_15207);
or U15706 (N_15706,N_15506,N_15261);
xnor U15707 (N_15707,N_15308,N_15081);
and U15708 (N_15708,N_15416,N_15051);
xor U15709 (N_15709,N_15036,N_15052);
and U15710 (N_15710,N_15028,N_15258);
and U15711 (N_15711,N_15039,N_15547);
or U15712 (N_15712,N_15305,N_15264);
nor U15713 (N_15713,N_15246,N_15053);
and U15714 (N_15714,N_15487,N_15241);
and U15715 (N_15715,N_15386,N_15078);
or U15716 (N_15716,N_15101,N_15376);
nor U15717 (N_15717,N_15154,N_15148);
xor U15718 (N_15718,N_15537,N_15022);
or U15719 (N_15719,N_15572,N_15558);
and U15720 (N_15720,N_15410,N_15339);
and U15721 (N_15721,N_15151,N_15189);
and U15722 (N_15722,N_15332,N_15431);
and U15723 (N_15723,N_15128,N_15144);
xnor U15724 (N_15724,N_15044,N_15163);
nand U15725 (N_15725,N_15182,N_15203);
and U15726 (N_15726,N_15200,N_15491);
and U15727 (N_15727,N_15260,N_15063);
or U15728 (N_15728,N_15455,N_15170);
xnor U15729 (N_15729,N_15213,N_15124);
or U15730 (N_15730,N_15100,N_15248);
nor U15731 (N_15731,N_15279,N_15216);
and U15732 (N_15732,N_15530,N_15010);
or U15733 (N_15733,N_15316,N_15369);
or U15734 (N_15734,N_15334,N_15311);
xor U15735 (N_15735,N_15234,N_15179);
nor U15736 (N_15736,N_15468,N_15069);
xor U15737 (N_15737,N_15142,N_15071);
nor U15738 (N_15738,N_15187,N_15513);
and U15739 (N_15739,N_15595,N_15294);
and U15740 (N_15740,N_15462,N_15467);
nor U15741 (N_15741,N_15229,N_15543);
or U15742 (N_15742,N_15357,N_15397);
xor U15743 (N_15743,N_15090,N_15275);
xnor U15744 (N_15744,N_15227,N_15237);
nand U15745 (N_15745,N_15498,N_15249);
nand U15746 (N_15746,N_15138,N_15368);
nor U15747 (N_15747,N_15116,N_15503);
or U15748 (N_15748,N_15003,N_15230);
and U15749 (N_15749,N_15136,N_15511);
and U15750 (N_15750,N_15573,N_15037);
xor U15751 (N_15751,N_15209,N_15224);
nand U15752 (N_15752,N_15152,N_15284);
and U15753 (N_15753,N_15281,N_15002);
or U15754 (N_15754,N_15104,N_15394);
or U15755 (N_15755,N_15354,N_15313);
and U15756 (N_15756,N_15398,N_15139);
nand U15757 (N_15757,N_15599,N_15319);
xor U15758 (N_15758,N_15201,N_15580);
or U15759 (N_15759,N_15526,N_15507);
nand U15760 (N_15760,N_15159,N_15168);
xnor U15761 (N_15761,N_15110,N_15259);
nor U15762 (N_15762,N_15250,N_15303);
nand U15763 (N_15763,N_15476,N_15538);
and U15764 (N_15764,N_15439,N_15049);
or U15765 (N_15765,N_15546,N_15586);
xnor U15766 (N_15766,N_15087,N_15333);
and U15767 (N_15767,N_15162,N_15559);
and U15768 (N_15768,N_15214,N_15564);
nand U15769 (N_15769,N_15244,N_15035);
or U15770 (N_15770,N_15208,N_15340);
or U15771 (N_15771,N_15122,N_15325);
nand U15772 (N_15772,N_15165,N_15464);
or U15773 (N_15773,N_15591,N_15210);
nor U15774 (N_15774,N_15502,N_15486);
or U15775 (N_15775,N_15016,N_15501);
nand U15776 (N_15776,N_15280,N_15300);
nand U15777 (N_15777,N_15447,N_15351);
nand U15778 (N_15778,N_15567,N_15344);
and U15779 (N_15779,N_15115,N_15589);
nand U15780 (N_15780,N_15038,N_15469);
and U15781 (N_15781,N_15262,N_15041);
nor U15782 (N_15782,N_15561,N_15276);
nand U15783 (N_15783,N_15111,N_15353);
nand U15784 (N_15784,N_15592,N_15356);
nand U15785 (N_15785,N_15125,N_15460);
or U15786 (N_15786,N_15518,N_15481);
or U15787 (N_15787,N_15545,N_15442);
and U15788 (N_15788,N_15480,N_15093);
or U15789 (N_15789,N_15195,N_15582);
nor U15790 (N_15790,N_15267,N_15013);
xor U15791 (N_15791,N_15031,N_15362);
and U15792 (N_15792,N_15441,N_15040);
and U15793 (N_15793,N_15391,N_15266);
or U15794 (N_15794,N_15269,N_15371);
xnor U15795 (N_15795,N_15174,N_15166);
nand U15796 (N_15796,N_15255,N_15014);
and U15797 (N_15797,N_15190,N_15387);
xor U15798 (N_15798,N_15454,N_15583);
nand U15799 (N_15799,N_15341,N_15329);
and U15800 (N_15800,N_15425,N_15153);
xor U15801 (N_15801,N_15593,N_15196);
and U15802 (N_15802,N_15544,N_15328);
nand U15803 (N_15803,N_15495,N_15215);
xnor U15804 (N_15804,N_15027,N_15551);
and U15805 (N_15805,N_15240,N_15355);
nand U15806 (N_15806,N_15068,N_15059);
nand U15807 (N_15807,N_15521,N_15146);
and U15808 (N_15808,N_15188,N_15436);
xor U15809 (N_15809,N_15243,N_15472);
nor U15810 (N_15810,N_15384,N_15176);
xnor U15811 (N_15811,N_15047,N_15553);
and U15812 (N_15812,N_15424,N_15206);
and U15813 (N_15813,N_15084,N_15514);
xnor U15814 (N_15814,N_15032,N_15519);
nor U15815 (N_15815,N_15317,N_15320);
xnor U15816 (N_15816,N_15594,N_15289);
nand U15817 (N_15817,N_15338,N_15226);
nor U15818 (N_15818,N_15500,N_15405);
nand U15819 (N_15819,N_15445,N_15515);
and U15820 (N_15820,N_15301,N_15277);
nand U15821 (N_15821,N_15568,N_15288);
nand U15822 (N_15822,N_15350,N_15364);
or U15823 (N_15823,N_15321,N_15587);
nand U15824 (N_15824,N_15286,N_15326);
nand U15825 (N_15825,N_15330,N_15536);
and U15826 (N_15826,N_15372,N_15465);
xor U15827 (N_15827,N_15192,N_15473);
and U15828 (N_15828,N_15000,N_15086);
and U15829 (N_15829,N_15422,N_15306);
or U15830 (N_15830,N_15018,N_15121);
nand U15831 (N_15831,N_15029,N_15535);
or U15832 (N_15832,N_15265,N_15452);
or U15833 (N_15833,N_15006,N_15088);
and U15834 (N_15834,N_15304,N_15420);
nand U15835 (N_15835,N_15030,N_15181);
or U15836 (N_15836,N_15220,N_15074);
nand U15837 (N_15837,N_15033,N_15366);
or U15838 (N_15838,N_15437,N_15477);
and U15839 (N_15839,N_15388,N_15161);
and U15840 (N_15840,N_15251,N_15085);
and U15841 (N_15841,N_15505,N_15548);
or U15842 (N_15842,N_15550,N_15440);
nand U15843 (N_15843,N_15517,N_15560);
or U15844 (N_15844,N_15430,N_15054);
and U15845 (N_15845,N_15523,N_15584);
and U15846 (N_15846,N_15566,N_15421);
or U15847 (N_15847,N_15221,N_15446);
and U15848 (N_15848,N_15079,N_15374);
or U15849 (N_15849,N_15004,N_15400);
xor U15850 (N_15850,N_15414,N_15395);
or U15851 (N_15851,N_15408,N_15392);
or U15852 (N_15852,N_15119,N_15254);
xnor U15853 (N_15853,N_15282,N_15015);
and U15854 (N_15854,N_15008,N_15349);
or U15855 (N_15855,N_15167,N_15141);
nand U15856 (N_15856,N_15380,N_15556);
xnor U15857 (N_15857,N_15204,N_15191);
nor U15858 (N_15858,N_15542,N_15409);
xor U15859 (N_15859,N_15272,N_15299);
or U15860 (N_15860,N_15057,N_15238);
nor U15861 (N_15861,N_15367,N_15082);
nor U15862 (N_15862,N_15156,N_15327);
xor U15863 (N_15863,N_15178,N_15483);
nand U15864 (N_15864,N_15137,N_15451);
or U15865 (N_15865,N_15524,N_15096);
nand U15866 (N_15866,N_15588,N_15019);
nor U15867 (N_15867,N_15073,N_15183);
or U15868 (N_15868,N_15118,N_15490);
and U15869 (N_15869,N_15512,N_15525);
or U15870 (N_15870,N_15378,N_15479);
and U15871 (N_15871,N_15094,N_15143);
nor U15872 (N_15872,N_15534,N_15007);
nor U15873 (N_15873,N_15043,N_15417);
xnor U15874 (N_15874,N_15126,N_15186);
nand U15875 (N_15875,N_15363,N_15193);
xnor U15876 (N_15876,N_15406,N_15323);
or U15877 (N_15877,N_15287,N_15324);
xnor U15878 (N_15878,N_15569,N_15135);
nand U15879 (N_15879,N_15202,N_15005);
and U15880 (N_15880,N_15381,N_15253);
nand U15881 (N_15881,N_15342,N_15218);
nor U15882 (N_15882,N_15223,N_15285);
nand U15883 (N_15883,N_15083,N_15164);
nor U15884 (N_15884,N_15058,N_15314);
nand U15885 (N_15885,N_15062,N_15132);
and U15886 (N_15886,N_15456,N_15365);
or U15887 (N_15887,N_15120,N_15075);
nand U15888 (N_15888,N_15443,N_15345);
and U15889 (N_15889,N_15466,N_15458);
nand U15890 (N_15890,N_15531,N_15418);
nor U15891 (N_15891,N_15510,N_15516);
or U15892 (N_15892,N_15295,N_15173);
and U15893 (N_15893,N_15103,N_15185);
or U15894 (N_15894,N_15385,N_15504);
or U15895 (N_15895,N_15312,N_15360);
or U15896 (N_15896,N_15433,N_15461);
nor U15897 (N_15897,N_15528,N_15428);
xor U15898 (N_15898,N_15070,N_15348);
xor U15899 (N_15899,N_15157,N_15105);
nand U15900 (N_15900,N_15300,N_15093);
or U15901 (N_15901,N_15249,N_15222);
xnor U15902 (N_15902,N_15403,N_15431);
nor U15903 (N_15903,N_15482,N_15271);
nor U15904 (N_15904,N_15409,N_15221);
and U15905 (N_15905,N_15131,N_15410);
and U15906 (N_15906,N_15420,N_15099);
nor U15907 (N_15907,N_15057,N_15286);
and U15908 (N_15908,N_15307,N_15447);
xor U15909 (N_15909,N_15301,N_15439);
nor U15910 (N_15910,N_15225,N_15576);
or U15911 (N_15911,N_15575,N_15147);
nand U15912 (N_15912,N_15517,N_15422);
or U15913 (N_15913,N_15297,N_15385);
nor U15914 (N_15914,N_15535,N_15456);
xor U15915 (N_15915,N_15164,N_15114);
or U15916 (N_15916,N_15168,N_15140);
nor U15917 (N_15917,N_15238,N_15155);
nor U15918 (N_15918,N_15563,N_15032);
xor U15919 (N_15919,N_15537,N_15231);
or U15920 (N_15920,N_15400,N_15370);
and U15921 (N_15921,N_15579,N_15349);
xnor U15922 (N_15922,N_15354,N_15168);
nand U15923 (N_15923,N_15597,N_15534);
nor U15924 (N_15924,N_15474,N_15424);
or U15925 (N_15925,N_15379,N_15399);
xnor U15926 (N_15926,N_15009,N_15339);
xnor U15927 (N_15927,N_15351,N_15084);
xnor U15928 (N_15928,N_15331,N_15060);
and U15929 (N_15929,N_15032,N_15344);
and U15930 (N_15930,N_15134,N_15131);
nand U15931 (N_15931,N_15557,N_15516);
or U15932 (N_15932,N_15230,N_15544);
xnor U15933 (N_15933,N_15368,N_15139);
and U15934 (N_15934,N_15335,N_15536);
and U15935 (N_15935,N_15354,N_15113);
nor U15936 (N_15936,N_15314,N_15160);
xor U15937 (N_15937,N_15207,N_15187);
or U15938 (N_15938,N_15337,N_15439);
xnor U15939 (N_15939,N_15389,N_15289);
and U15940 (N_15940,N_15564,N_15530);
nor U15941 (N_15941,N_15348,N_15569);
or U15942 (N_15942,N_15564,N_15516);
nand U15943 (N_15943,N_15373,N_15595);
nor U15944 (N_15944,N_15342,N_15015);
and U15945 (N_15945,N_15298,N_15403);
or U15946 (N_15946,N_15098,N_15368);
nand U15947 (N_15947,N_15565,N_15359);
nor U15948 (N_15948,N_15399,N_15441);
xor U15949 (N_15949,N_15219,N_15428);
and U15950 (N_15950,N_15166,N_15092);
or U15951 (N_15951,N_15166,N_15437);
or U15952 (N_15952,N_15560,N_15196);
or U15953 (N_15953,N_15333,N_15192);
or U15954 (N_15954,N_15440,N_15594);
and U15955 (N_15955,N_15549,N_15049);
or U15956 (N_15956,N_15483,N_15308);
nor U15957 (N_15957,N_15001,N_15400);
xor U15958 (N_15958,N_15066,N_15434);
and U15959 (N_15959,N_15328,N_15543);
or U15960 (N_15960,N_15331,N_15056);
or U15961 (N_15961,N_15439,N_15053);
nor U15962 (N_15962,N_15328,N_15568);
nand U15963 (N_15963,N_15508,N_15139);
nand U15964 (N_15964,N_15317,N_15426);
or U15965 (N_15965,N_15527,N_15018);
or U15966 (N_15966,N_15336,N_15401);
and U15967 (N_15967,N_15109,N_15359);
or U15968 (N_15968,N_15247,N_15026);
or U15969 (N_15969,N_15046,N_15363);
and U15970 (N_15970,N_15119,N_15483);
nand U15971 (N_15971,N_15077,N_15561);
nor U15972 (N_15972,N_15123,N_15574);
nand U15973 (N_15973,N_15182,N_15448);
nor U15974 (N_15974,N_15570,N_15483);
or U15975 (N_15975,N_15444,N_15135);
or U15976 (N_15976,N_15250,N_15305);
xor U15977 (N_15977,N_15462,N_15005);
or U15978 (N_15978,N_15288,N_15163);
or U15979 (N_15979,N_15362,N_15167);
or U15980 (N_15980,N_15230,N_15377);
and U15981 (N_15981,N_15547,N_15163);
xnor U15982 (N_15982,N_15188,N_15143);
nor U15983 (N_15983,N_15336,N_15212);
nor U15984 (N_15984,N_15272,N_15470);
nor U15985 (N_15985,N_15437,N_15407);
xor U15986 (N_15986,N_15368,N_15575);
nor U15987 (N_15987,N_15359,N_15411);
or U15988 (N_15988,N_15517,N_15452);
or U15989 (N_15989,N_15406,N_15217);
and U15990 (N_15990,N_15136,N_15354);
nand U15991 (N_15991,N_15519,N_15493);
xnor U15992 (N_15992,N_15492,N_15104);
xnor U15993 (N_15993,N_15460,N_15492);
and U15994 (N_15994,N_15194,N_15304);
nor U15995 (N_15995,N_15391,N_15236);
or U15996 (N_15996,N_15519,N_15056);
xnor U15997 (N_15997,N_15255,N_15331);
nor U15998 (N_15998,N_15027,N_15164);
or U15999 (N_15999,N_15088,N_15106);
nand U16000 (N_16000,N_15071,N_15471);
or U16001 (N_16001,N_15367,N_15502);
nand U16002 (N_16002,N_15317,N_15241);
nand U16003 (N_16003,N_15461,N_15460);
nand U16004 (N_16004,N_15003,N_15319);
nor U16005 (N_16005,N_15158,N_15388);
xnor U16006 (N_16006,N_15277,N_15311);
xnor U16007 (N_16007,N_15399,N_15052);
nand U16008 (N_16008,N_15192,N_15031);
or U16009 (N_16009,N_15071,N_15328);
or U16010 (N_16010,N_15482,N_15532);
nor U16011 (N_16011,N_15268,N_15532);
and U16012 (N_16012,N_15048,N_15075);
or U16013 (N_16013,N_15218,N_15339);
xor U16014 (N_16014,N_15126,N_15505);
and U16015 (N_16015,N_15437,N_15028);
xor U16016 (N_16016,N_15227,N_15112);
nor U16017 (N_16017,N_15126,N_15125);
and U16018 (N_16018,N_15338,N_15371);
xnor U16019 (N_16019,N_15345,N_15586);
xnor U16020 (N_16020,N_15406,N_15316);
nor U16021 (N_16021,N_15481,N_15358);
or U16022 (N_16022,N_15169,N_15187);
xnor U16023 (N_16023,N_15358,N_15372);
nor U16024 (N_16024,N_15475,N_15245);
nand U16025 (N_16025,N_15528,N_15559);
xnor U16026 (N_16026,N_15396,N_15591);
nor U16027 (N_16027,N_15138,N_15292);
and U16028 (N_16028,N_15145,N_15361);
nor U16029 (N_16029,N_15500,N_15438);
nor U16030 (N_16030,N_15162,N_15113);
nor U16031 (N_16031,N_15203,N_15126);
xor U16032 (N_16032,N_15554,N_15080);
nor U16033 (N_16033,N_15335,N_15393);
or U16034 (N_16034,N_15280,N_15015);
xor U16035 (N_16035,N_15091,N_15533);
xor U16036 (N_16036,N_15012,N_15048);
nor U16037 (N_16037,N_15280,N_15325);
or U16038 (N_16038,N_15099,N_15523);
or U16039 (N_16039,N_15234,N_15510);
xor U16040 (N_16040,N_15379,N_15373);
or U16041 (N_16041,N_15152,N_15353);
or U16042 (N_16042,N_15392,N_15300);
or U16043 (N_16043,N_15567,N_15427);
xor U16044 (N_16044,N_15170,N_15394);
xor U16045 (N_16045,N_15300,N_15429);
or U16046 (N_16046,N_15190,N_15382);
xor U16047 (N_16047,N_15307,N_15259);
nand U16048 (N_16048,N_15508,N_15114);
and U16049 (N_16049,N_15337,N_15556);
and U16050 (N_16050,N_15247,N_15236);
or U16051 (N_16051,N_15559,N_15365);
nor U16052 (N_16052,N_15122,N_15509);
nor U16053 (N_16053,N_15218,N_15340);
nor U16054 (N_16054,N_15216,N_15272);
nor U16055 (N_16055,N_15056,N_15487);
nor U16056 (N_16056,N_15579,N_15538);
and U16057 (N_16057,N_15542,N_15334);
nor U16058 (N_16058,N_15471,N_15452);
xnor U16059 (N_16059,N_15331,N_15563);
nor U16060 (N_16060,N_15063,N_15214);
nand U16061 (N_16061,N_15224,N_15311);
nand U16062 (N_16062,N_15570,N_15224);
nand U16063 (N_16063,N_15136,N_15076);
and U16064 (N_16064,N_15293,N_15445);
nand U16065 (N_16065,N_15470,N_15544);
or U16066 (N_16066,N_15397,N_15392);
and U16067 (N_16067,N_15588,N_15121);
nor U16068 (N_16068,N_15143,N_15599);
nand U16069 (N_16069,N_15570,N_15353);
xor U16070 (N_16070,N_15258,N_15474);
xnor U16071 (N_16071,N_15266,N_15243);
and U16072 (N_16072,N_15554,N_15065);
or U16073 (N_16073,N_15134,N_15418);
and U16074 (N_16074,N_15294,N_15093);
nand U16075 (N_16075,N_15122,N_15209);
and U16076 (N_16076,N_15176,N_15480);
xnor U16077 (N_16077,N_15136,N_15304);
or U16078 (N_16078,N_15408,N_15505);
nand U16079 (N_16079,N_15045,N_15596);
xnor U16080 (N_16080,N_15109,N_15086);
nor U16081 (N_16081,N_15401,N_15339);
nand U16082 (N_16082,N_15265,N_15578);
and U16083 (N_16083,N_15029,N_15425);
nor U16084 (N_16084,N_15535,N_15078);
and U16085 (N_16085,N_15397,N_15132);
xnor U16086 (N_16086,N_15582,N_15111);
xnor U16087 (N_16087,N_15000,N_15158);
xor U16088 (N_16088,N_15197,N_15173);
and U16089 (N_16089,N_15053,N_15213);
nor U16090 (N_16090,N_15149,N_15084);
nor U16091 (N_16091,N_15137,N_15478);
or U16092 (N_16092,N_15157,N_15232);
nor U16093 (N_16093,N_15178,N_15471);
nor U16094 (N_16094,N_15248,N_15214);
and U16095 (N_16095,N_15279,N_15420);
nand U16096 (N_16096,N_15442,N_15257);
and U16097 (N_16097,N_15540,N_15170);
nand U16098 (N_16098,N_15000,N_15107);
or U16099 (N_16099,N_15160,N_15504);
nor U16100 (N_16100,N_15154,N_15222);
nand U16101 (N_16101,N_15027,N_15321);
xor U16102 (N_16102,N_15508,N_15364);
xor U16103 (N_16103,N_15161,N_15439);
xor U16104 (N_16104,N_15348,N_15426);
or U16105 (N_16105,N_15169,N_15573);
or U16106 (N_16106,N_15022,N_15349);
nand U16107 (N_16107,N_15384,N_15272);
nor U16108 (N_16108,N_15071,N_15118);
nand U16109 (N_16109,N_15238,N_15375);
nor U16110 (N_16110,N_15109,N_15449);
or U16111 (N_16111,N_15105,N_15002);
nor U16112 (N_16112,N_15507,N_15320);
nand U16113 (N_16113,N_15371,N_15475);
nand U16114 (N_16114,N_15489,N_15368);
nand U16115 (N_16115,N_15203,N_15223);
or U16116 (N_16116,N_15539,N_15483);
or U16117 (N_16117,N_15196,N_15229);
nor U16118 (N_16118,N_15502,N_15352);
or U16119 (N_16119,N_15590,N_15274);
nand U16120 (N_16120,N_15493,N_15404);
xnor U16121 (N_16121,N_15513,N_15138);
nand U16122 (N_16122,N_15558,N_15186);
xnor U16123 (N_16123,N_15259,N_15199);
and U16124 (N_16124,N_15240,N_15235);
xnor U16125 (N_16125,N_15546,N_15564);
and U16126 (N_16126,N_15026,N_15386);
nor U16127 (N_16127,N_15237,N_15545);
xnor U16128 (N_16128,N_15076,N_15430);
and U16129 (N_16129,N_15500,N_15581);
nor U16130 (N_16130,N_15169,N_15007);
and U16131 (N_16131,N_15312,N_15545);
nand U16132 (N_16132,N_15220,N_15270);
and U16133 (N_16133,N_15071,N_15199);
or U16134 (N_16134,N_15514,N_15274);
nor U16135 (N_16135,N_15085,N_15537);
xnor U16136 (N_16136,N_15537,N_15155);
or U16137 (N_16137,N_15383,N_15066);
nor U16138 (N_16138,N_15408,N_15376);
and U16139 (N_16139,N_15096,N_15447);
nor U16140 (N_16140,N_15449,N_15057);
nand U16141 (N_16141,N_15195,N_15361);
nor U16142 (N_16142,N_15567,N_15142);
xnor U16143 (N_16143,N_15080,N_15239);
nor U16144 (N_16144,N_15156,N_15190);
xor U16145 (N_16145,N_15076,N_15134);
nand U16146 (N_16146,N_15142,N_15555);
nor U16147 (N_16147,N_15476,N_15266);
or U16148 (N_16148,N_15291,N_15255);
xor U16149 (N_16149,N_15293,N_15315);
xnor U16150 (N_16150,N_15125,N_15118);
xor U16151 (N_16151,N_15456,N_15102);
xnor U16152 (N_16152,N_15167,N_15180);
or U16153 (N_16153,N_15331,N_15301);
xor U16154 (N_16154,N_15428,N_15523);
or U16155 (N_16155,N_15169,N_15402);
xnor U16156 (N_16156,N_15050,N_15201);
nand U16157 (N_16157,N_15581,N_15566);
xor U16158 (N_16158,N_15052,N_15321);
or U16159 (N_16159,N_15054,N_15550);
and U16160 (N_16160,N_15282,N_15233);
xnor U16161 (N_16161,N_15457,N_15136);
and U16162 (N_16162,N_15588,N_15277);
nand U16163 (N_16163,N_15532,N_15414);
and U16164 (N_16164,N_15181,N_15504);
xor U16165 (N_16165,N_15019,N_15502);
or U16166 (N_16166,N_15462,N_15185);
nor U16167 (N_16167,N_15421,N_15365);
or U16168 (N_16168,N_15541,N_15161);
and U16169 (N_16169,N_15222,N_15575);
xnor U16170 (N_16170,N_15257,N_15405);
and U16171 (N_16171,N_15560,N_15291);
and U16172 (N_16172,N_15062,N_15047);
nor U16173 (N_16173,N_15088,N_15338);
and U16174 (N_16174,N_15460,N_15121);
nor U16175 (N_16175,N_15126,N_15052);
xor U16176 (N_16176,N_15056,N_15430);
xnor U16177 (N_16177,N_15376,N_15591);
or U16178 (N_16178,N_15381,N_15489);
or U16179 (N_16179,N_15146,N_15354);
nand U16180 (N_16180,N_15332,N_15020);
and U16181 (N_16181,N_15395,N_15599);
nor U16182 (N_16182,N_15046,N_15293);
or U16183 (N_16183,N_15559,N_15161);
xor U16184 (N_16184,N_15387,N_15209);
or U16185 (N_16185,N_15293,N_15568);
xor U16186 (N_16186,N_15487,N_15508);
xnor U16187 (N_16187,N_15004,N_15018);
or U16188 (N_16188,N_15051,N_15506);
nor U16189 (N_16189,N_15229,N_15439);
nand U16190 (N_16190,N_15428,N_15056);
or U16191 (N_16191,N_15348,N_15517);
nor U16192 (N_16192,N_15059,N_15422);
nor U16193 (N_16193,N_15485,N_15543);
nor U16194 (N_16194,N_15200,N_15057);
and U16195 (N_16195,N_15527,N_15585);
nand U16196 (N_16196,N_15374,N_15414);
nand U16197 (N_16197,N_15293,N_15345);
nand U16198 (N_16198,N_15270,N_15210);
or U16199 (N_16199,N_15289,N_15176);
and U16200 (N_16200,N_16010,N_15645);
xnor U16201 (N_16201,N_15907,N_15940);
nand U16202 (N_16202,N_16071,N_16107);
nor U16203 (N_16203,N_15727,N_15931);
nand U16204 (N_16204,N_15612,N_16026);
nand U16205 (N_16205,N_15747,N_15871);
xor U16206 (N_16206,N_16062,N_16185);
nand U16207 (N_16207,N_15888,N_16189);
nor U16208 (N_16208,N_15811,N_15839);
nand U16209 (N_16209,N_16106,N_16080);
or U16210 (N_16210,N_15772,N_15854);
xor U16211 (N_16211,N_15729,N_16162);
xor U16212 (N_16212,N_15936,N_16149);
or U16213 (N_16213,N_15987,N_15771);
nand U16214 (N_16214,N_15915,N_16158);
and U16215 (N_16215,N_15718,N_16049);
nor U16216 (N_16216,N_16160,N_16088);
xor U16217 (N_16217,N_15670,N_16115);
nor U16218 (N_16218,N_15673,N_15789);
nand U16219 (N_16219,N_15827,N_15898);
nand U16220 (N_16220,N_15949,N_16138);
or U16221 (N_16221,N_16016,N_15722);
or U16222 (N_16222,N_16086,N_16199);
xnor U16223 (N_16223,N_16155,N_15635);
nor U16224 (N_16224,N_15976,N_15684);
or U16225 (N_16225,N_15646,N_15668);
or U16226 (N_16226,N_15737,N_15958);
or U16227 (N_16227,N_15641,N_16083);
and U16228 (N_16228,N_15875,N_15858);
xnor U16229 (N_16229,N_16125,N_15923);
nor U16230 (N_16230,N_16169,N_15969);
and U16231 (N_16231,N_16003,N_15766);
or U16232 (N_16232,N_15815,N_15748);
and U16233 (N_16233,N_15638,N_16060);
nor U16234 (N_16234,N_15607,N_16157);
xor U16235 (N_16235,N_16075,N_16153);
nor U16236 (N_16236,N_15807,N_15889);
or U16237 (N_16237,N_16108,N_15647);
nor U16238 (N_16238,N_16087,N_15819);
or U16239 (N_16239,N_16116,N_15995);
nand U16240 (N_16240,N_15939,N_15672);
nor U16241 (N_16241,N_15619,N_16066);
xor U16242 (N_16242,N_16048,N_15829);
nand U16243 (N_16243,N_15719,N_15971);
nor U16244 (N_16244,N_15917,N_16102);
and U16245 (N_16245,N_16164,N_16032);
and U16246 (N_16246,N_15860,N_15950);
or U16247 (N_16247,N_15880,N_15796);
and U16248 (N_16248,N_15680,N_16178);
nor U16249 (N_16249,N_15754,N_15629);
xor U16250 (N_16250,N_16105,N_15895);
and U16251 (N_16251,N_15894,N_15806);
and U16252 (N_16252,N_15948,N_16068);
nor U16253 (N_16253,N_15890,N_15797);
xnor U16254 (N_16254,N_16166,N_15702);
nand U16255 (N_16255,N_16132,N_16047);
nand U16256 (N_16256,N_15838,N_16101);
nand U16257 (N_16257,N_16037,N_16100);
or U16258 (N_16258,N_16156,N_15669);
nor U16259 (N_16259,N_15660,N_16076);
or U16260 (N_16260,N_15699,N_15926);
nand U16261 (N_16261,N_15818,N_15897);
nor U16262 (N_16262,N_16197,N_15834);
and U16263 (N_16263,N_15959,N_15998);
xor U16264 (N_16264,N_15882,N_16079);
nand U16265 (N_16265,N_16191,N_16146);
nor U16266 (N_16266,N_16096,N_16002);
or U16267 (N_16267,N_15755,N_16018);
nor U16268 (N_16268,N_15640,N_16024);
and U16269 (N_16269,N_15903,N_15774);
nand U16270 (N_16270,N_15698,N_16030);
or U16271 (N_16271,N_15659,N_15961);
nor U16272 (N_16272,N_15753,N_15787);
or U16273 (N_16273,N_16182,N_16020);
or U16274 (N_16274,N_15964,N_16175);
nand U16275 (N_16275,N_16194,N_15937);
xor U16276 (N_16276,N_15686,N_15919);
nand U16277 (N_16277,N_15862,N_16192);
xnor U16278 (N_16278,N_15769,N_15982);
and U16279 (N_16279,N_15655,N_16184);
and U16280 (N_16280,N_16120,N_15687);
nand U16281 (N_16281,N_15928,N_15828);
xnor U16282 (N_16282,N_15975,N_15902);
and U16283 (N_16283,N_15658,N_15996);
and U16284 (N_16284,N_15761,N_16034);
nor U16285 (N_16285,N_16198,N_16055);
xnor U16286 (N_16286,N_15911,N_15821);
and U16287 (N_16287,N_16085,N_15760);
nor U16288 (N_16288,N_16104,N_16114);
xor U16289 (N_16289,N_15681,N_16078);
or U16290 (N_16290,N_15798,N_16176);
xor U16291 (N_16291,N_15929,N_16033);
and U16292 (N_16292,N_15981,N_16006);
and U16293 (N_16293,N_15892,N_16064);
and U16294 (N_16294,N_15900,N_15914);
nand U16295 (N_16295,N_15820,N_15868);
xnor U16296 (N_16296,N_16117,N_15795);
or U16297 (N_16297,N_15803,N_15785);
or U16298 (N_16298,N_16172,N_16056);
xnor U16299 (N_16299,N_15884,N_15954);
xnor U16300 (N_16300,N_15628,N_15901);
or U16301 (N_16301,N_15865,N_15666);
or U16302 (N_16302,N_16031,N_15651);
or U16303 (N_16303,N_15767,N_15616);
nor U16304 (N_16304,N_16009,N_15763);
xor U16305 (N_16305,N_15726,N_15707);
nand U16306 (N_16306,N_15625,N_15904);
nand U16307 (N_16307,N_15848,N_16111);
nor U16308 (N_16308,N_15733,N_15816);
nand U16309 (N_16309,N_16007,N_15768);
or U16310 (N_16310,N_15750,N_15891);
nand U16311 (N_16311,N_15730,N_16040);
nand U16312 (N_16312,N_16112,N_15709);
and U16313 (N_16313,N_15801,N_15824);
nor U16314 (N_16314,N_15742,N_16130);
nand U16315 (N_16315,N_15759,N_15746);
or U16316 (N_16316,N_15953,N_15777);
nand U16317 (N_16317,N_15963,N_16163);
and U16318 (N_16318,N_15986,N_15951);
nor U16319 (N_16319,N_15810,N_16095);
xnor U16320 (N_16320,N_16063,N_16196);
nand U16321 (N_16321,N_15715,N_15675);
nor U16322 (N_16322,N_15695,N_15653);
nor U16323 (N_16323,N_15861,N_16081);
nand U16324 (N_16324,N_15621,N_15690);
nor U16325 (N_16325,N_16124,N_15930);
xor U16326 (N_16326,N_16054,N_15602);
and U16327 (N_16327,N_16186,N_15974);
xor U16328 (N_16328,N_15657,N_15704);
xor U16329 (N_16329,N_15970,N_15832);
nand U16330 (N_16330,N_15855,N_15683);
xnor U16331 (N_16331,N_15739,N_15790);
and U16332 (N_16332,N_15765,N_15946);
nor U16333 (N_16333,N_16165,N_15786);
xor U16334 (N_16334,N_16039,N_15853);
xnor U16335 (N_16335,N_15648,N_15637);
xnor U16336 (N_16336,N_16011,N_16070);
nor U16337 (N_16337,N_16084,N_16097);
xnor U16338 (N_16338,N_15905,N_15724);
nand U16339 (N_16339,N_15847,N_16029);
nor U16340 (N_16340,N_16028,N_15992);
and U16341 (N_16341,N_15751,N_16061);
or U16342 (N_16342,N_15627,N_15644);
nand U16343 (N_16343,N_16058,N_15610);
nor U16344 (N_16344,N_15706,N_16093);
nand U16345 (N_16345,N_15909,N_15994);
xnor U16346 (N_16346,N_15791,N_15682);
xor U16347 (N_16347,N_15856,N_15650);
and U16348 (N_16348,N_15631,N_16126);
nand U16349 (N_16349,N_15925,N_15843);
or U16350 (N_16350,N_15944,N_15879);
or U16351 (N_16351,N_15661,N_15967);
or U16352 (N_16352,N_15764,N_16137);
xor U16353 (N_16353,N_16065,N_16167);
nand U16354 (N_16354,N_15910,N_16131);
nand U16355 (N_16355,N_16135,N_15935);
nand U16356 (N_16356,N_16035,N_15775);
xor U16357 (N_16357,N_15700,N_15703);
or U16358 (N_16358,N_15745,N_15922);
or U16359 (N_16359,N_15857,N_16143);
nor U16360 (N_16360,N_15942,N_15988);
and U16361 (N_16361,N_16050,N_15823);
nor U16362 (N_16362,N_15979,N_15850);
xor U16363 (N_16363,N_15972,N_15649);
xnor U16364 (N_16364,N_15913,N_16103);
or U16365 (N_16365,N_15933,N_15626);
nor U16366 (N_16366,N_15980,N_15614);
xor U16367 (N_16367,N_15620,N_16113);
or U16368 (N_16368,N_15756,N_15692);
or U16369 (N_16369,N_15608,N_15749);
nand U16370 (N_16370,N_16170,N_15735);
nor U16371 (N_16371,N_15691,N_15783);
nand U16372 (N_16372,N_15656,N_16168);
or U16373 (N_16373,N_15615,N_15738);
or U16374 (N_16374,N_16001,N_16119);
nand U16375 (N_16375,N_15984,N_16193);
or U16376 (N_16376,N_16013,N_15603);
nand U16377 (N_16377,N_15717,N_15770);
or U16378 (N_16378,N_16159,N_16161);
nand U16379 (N_16379,N_15881,N_15654);
xor U16380 (N_16380,N_16091,N_16023);
and U16381 (N_16381,N_15960,N_15962);
and U16382 (N_16382,N_16183,N_15991);
nand U16383 (N_16383,N_15870,N_16110);
or U16384 (N_16384,N_15725,N_15920);
xnor U16385 (N_16385,N_15973,N_16052);
xnor U16386 (N_16386,N_16098,N_15956);
and U16387 (N_16387,N_15943,N_15697);
xnor U16388 (N_16388,N_15630,N_16123);
nor U16389 (N_16389,N_15852,N_15873);
or U16390 (N_16390,N_15613,N_15934);
nor U16391 (N_16391,N_15731,N_15983);
and U16392 (N_16392,N_15957,N_15859);
or U16393 (N_16393,N_15837,N_15711);
xor U16394 (N_16394,N_15604,N_16000);
nand U16395 (N_16395,N_15993,N_16027);
nand U16396 (N_16396,N_15864,N_16118);
nor U16397 (N_16397,N_15825,N_15849);
or U16398 (N_16398,N_15622,N_15883);
and U16399 (N_16399,N_16004,N_16129);
nor U16400 (N_16400,N_15623,N_16141);
nor U16401 (N_16401,N_15714,N_15918);
or U16402 (N_16402,N_16042,N_15841);
or U16403 (N_16403,N_16036,N_15710);
nand U16404 (N_16404,N_16152,N_15835);
xor U16405 (N_16405,N_16072,N_16046);
nand U16406 (N_16406,N_15833,N_15809);
nor U16407 (N_16407,N_15851,N_15800);
nor U16408 (N_16408,N_16077,N_16179);
or U16409 (N_16409,N_16044,N_16038);
nand U16410 (N_16410,N_15965,N_15643);
nor U16411 (N_16411,N_16059,N_15633);
and U16412 (N_16412,N_15652,N_15693);
nand U16413 (N_16413,N_15664,N_16187);
xor U16414 (N_16414,N_15966,N_15867);
xor U16415 (N_16415,N_16127,N_15696);
and U16416 (N_16416,N_15744,N_16148);
xor U16417 (N_16417,N_16090,N_15813);
xnor U16418 (N_16418,N_16043,N_15708);
xnor U16419 (N_16419,N_16017,N_15788);
or U16420 (N_16420,N_15671,N_16051);
nand U16421 (N_16421,N_16019,N_15740);
nor U16422 (N_16422,N_16134,N_15845);
nand U16423 (N_16423,N_16190,N_15872);
xnor U16424 (N_16424,N_15887,N_15694);
nor U16425 (N_16425,N_16012,N_15779);
nand U16426 (N_16426,N_16171,N_15716);
and U16427 (N_16427,N_15844,N_15878);
and U16428 (N_16428,N_16144,N_15757);
nor U16429 (N_16429,N_15721,N_16180);
xnor U16430 (N_16430,N_15938,N_15977);
nand U16431 (N_16431,N_16074,N_15600);
nand U16432 (N_16432,N_15676,N_15893);
nand U16433 (N_16433,N_15876,N_15712);
or U16434 (N_16434,N_15784,N_15874);
xor U16435 (N_16435,N_16008,N_15678);
or U16436 (N_16436,N_15822,N_16128);
xor U16437 (N_16437,N_16173,N_15906);
and U16438 (N_16438,N_16121,N_15932);
nand U16439 (N_16439,N_16139,N_15952);
nand U16440 (N_16440,N_15677,N_15831);
nor U16441 (N_16441,N_16045,N_15634);
and U16442 (N_16442,N_15978,N_15743);
and U16443 (N_16443,N_16094,N_16073);
and U16444 (N_16444,N_15812,N_15877);
xor U16445 (N_16445,N_15758,N_15762);
nor U16446 (N_16446,N_15781,N_15632);
nor U16447 (N_16447,N_16021,N_15814);
nor U16448 (N_16448,N_16082,N_16109);
nand U16449 (N_16449,N_16188,N_15705);
nand U16450 (N_16450,N_15782,N_15817);
nor U16451 (N_16451,N_15802,N_15773);
nand U16452 (N_16452,N_16145,N_15732);
and U16453 (N_16453,N_15679,N_15799);
nor U16454 (N_16454,N_15941,N_15728);
nor U16455 (N_16455,N_16150,N_16136);
and U16456 (N_16456,N_15605,N_16142);
nand U16457 (N_16457,N_15805,N_15611);
nand U16458 (N_16458,N_15793,N_15924);
and U16459 (N_16459,N_15912,N_15667);
and U16460 (N_16460,N_15990,N_15618);
or U16461 (N_16461,N_15734,N_15609);
xnor U16462 (N_16462,N_15685,N_15908);
nor U16463 (N_16463,N_15896,N_16140);
nand U16464 (N_16464,N_15863,N_15955);
and U16465 (N_16465,N_16181,N_16053);
nand U16466 (N_16466,N_15778,N_16099);
xor U16467 (N_16467,N_15663,N_15866);
xnor U16468 (N_16468,N_15921,N_15968);
nor U16469 (N_16469,N_16151,N_15720);
or U16470 (N_16470,N_15804,N_15997);
xnor U16471 (N_16471,N_15639,N_16057);
xnor U16472 (N_16472,N_15662,N_16174);
xnor U16473 (N_16473,N_15840,N_16195);
nor U16474 (N_16474,N_16089,N_15665);
or U16475 (N_16475,N_15945,N_15989);
and U16476 (N_16476,N_15642,N_15688);
nand U16477 (N_16477,N_15794,N_16177);
and U16478 (N_16478,N_16005,N_15792);
nand U16479 (N_16479,N_16041,N_15601);
or U16480 (N_16480,N_16014,N_16122);
xor U16481 (N_16481,N_15885,N_15899);
and U16482 (N_16482,N_15886,N_16154);
nor U16483 (N_16483,N_16147,N_15776);
xnor U16484 (N_16484,N_15999,N_15624);
or U16485 (N_16485,N_15689,N_15836);
and U16486 (N_16486,N_15723,N_16022);
and U16487 (N_16487,N_15830,N_15947);
and U16488 (N_16488,N_15846,N_15636);
nand U16489 (N_16489,N_15674,N_15736);
xor U16490 (N_16490,N_15741,N_15826);
nor U16491 (N_16491,N_15752,N_16069);
nand U16492 (N_16492,N_15916,N_16025);
xor U16493 (N_16493,N_16133,N_15780);
and U16494 (N_16494,N_15713,N_15808);
or U16495 (N_16495,N_16067,N_15606);
or U16496 (N_16496,N_15701,N_15617);
nand U16497 (N_16497,N_15927,N_15985);
nand U16498 (N_16498,N_16092,N_16015);
nand U16499 (N_16499,N_15869,N_15842);
and U16500 (N_16500,N_16068,N_15843);
xnor U16501 (N_16501,N_15888,N_15919);
nand U16502 (N_16502,N_15714,N_15669);
nand U16503 (N_16503,N_15907,N_16192);
or U16504 (N_16504,N_16032,N_15851);
nand U16505 (N_16505,N_16067,N_15631);
or U16506 (N_16506,N_16149,N_15869);
nor U16507 (N_16507,N_16025,N_16162);
xor U16508 (N_16508,N_15790,N_15869);
and U16509 (N_16509,N_15743,N_15816);
and U16510 (N_16510,N_15781,N_15933);
or U16511 (N_16511,N_15975,N_15792);
nand U16512 (N_16512,N_16151,N_15792);
or U16513 (N_16513,N_16188,N_15630);
or U16514 (N_16514,N_15755,N_15615);
and U16515 (N_16515,N_16054,N_15659);
xor U16516 (N_16516,N_16123,N_15985);
nand U16517 (N_16517,N_16042,N_15829);
nand U16518 (N_16518,N_15789,N_15613);
or U16519 (N_16519,N_15732,N_16181);
xnor U16520 (N_16520,N_15974,N_16082);
xor U16521 (N_16521,N_16163,N_16191);
xor U16522 (N_16522,N_15889,N_15942);
nand U16523 (N_16523,N_15747,N_15819);
nand U16524 (N_16524,N_15810,N_15609);
xor U16525 (N_16525,N_15758,N_15911);
and U16526 (N_16526,N_15682,N_15860);
nand U16527 (N_16527,N_15785,N_16112);
or U16528 (N_16528,N_16124,N_16005);
or U16529 (N_16529,N_15999,N_15673);
xor U16530 (N_16530,N_15679,N_16067);
xnor U16531 (N_16531,N_16029,N_15611);
xnor U16532 (N_16532,N_16131,N_16183);
or U16533 (N_16533,N_15832,N_15943);
xor U16534 (N_16534,N_15741,N_15670);
xnor U16535 (N_16535,N_16113,N_15925);
or U16536 (N_16536,N_15796,N_15700);
and U16537 (N_16537,N_15748,N_15984);
nand U16538 (N_16538,N_15671,N_15661);
nand U16539 (N_16539,N_15882,N_15605);
xnor U16540 (N_16540,N_15686,N_15658);
and U16541 (N_16541,N_15941,N_15632);
or U16542 (N_16542,N_15993,N_15690);
xnor U16543 (N_16543,N_15756,N_15669);
nand U16544 (N_16544,N_15709,N_15638);
nand U16545 (N_16545,N_15847,N_16011);
or U16546 (N_16546,N_16121,N_16025);
or U16547 (N_16547,N_15940,N_15836);
or U16548 (N_16548,N_16055,N_15731);
nor U16549 (N_16549,N_16035,N_15859);
and U16550 (N_16550,N_16098,N_15728);
xor U16551 (N_16551,N_15621,N_16149);
xnor U16552 (N_16552,N_16109,N_15713);
and U16553 (N_16553,N_15684,N_15812);
nand U16554 (N_16554,N_15755,N_16108);
or U16555 (N_16555,N_16101,N_16028);
xnor U16556 (N_16556,N_15751,N_15934);
and U16557 (N_16557,N_15991,N_15665);
nor U16558 (N_16558,N_15794,N_15924);
nand U16559 (N_16559,N_16153,N_15810);
and U16560 (N_16560,N_16079,N_16036);
or U16561 (N_16561,N_16196,N_15891);
nor U16562 (N_16562,N_16021,N_15734);
and U16563 (N_16563,N_15926,N_16070);
and U16564 (N_16564,N_16110,N_15756);
nand U16565 (N_16565,N_15904,N_15744);
or U16566 (N_16566,N_15988,N_15912);
or U16567 (N_16567,N_15738,N_15837);
and U16568 (N_16568,N_15609,N_16141);
xor U16569 (N_16569,N_15938,N_15876);
nor U16570 (N_16570,N_15816,N_16192);
xnor U16571 (N_16571,N_15663,N_16168);
xnor U16572 (N_16572,N_15623,N_15785);
nand U16573 (N_16573,N_16041,N_16008);
xor U16574 (N_16574,N_15760,N_15638);
xor U16575 (N_16575,N_15834,N_15957);
xnor U16576 (N_16576,N_16151,N_15713);
and U16577 (N_16577,N_16015,N_15935);
and U16578 (N_16578,N_16187,N_15692);
nand U16579 (N_16579,N_16150,N_15688);
and U16580 (N_16580,N_15789,N_15632);
nor U16581 (N_16581,N_15992,N_15941);
xor U16582 (N_16582,N_15792,N_15703);
and U16583 (N_16583,N_15987,N_15942);
nand U16584 (N_16584,N_16136,N_16003);
and U16585 (N_16585,N_15895,N_15727);
nor U16586 (N_16586,N_15923,N_16121);
nor U16587 (N_16587,N_15823,N_15759);
nor U16588 (N_16588,N_16153,N_16128);
nand U16589 (N_16589,N_15775,N_15735);
or U16590 (N_16590,N_16186,N_15689);
nor U16591 (N_16591,N_15870,N_15894);
nand U16592 (N_16592,N_15652,N_16038);
xnor U16593 (N_16593,N_15953,N_15602);
xnor U16594 (N_16594,N_15869,N_15962);
nor U16595 (N_16595,N_15909,N_16146);
nand U16596 (N_16596,N_16028,N_15818);
nor U16597 (N_16597,N_15659,N_16075);
xor U16598 (N_16598,N_15893,N_15925);
nor U16599 (N_16599,N_16154,N_15954);
and U16600 (N_16600,N_15847,N_15963);
xnor U16601 (N_16601,N_15751,N_16120);
and U16602 (N_16602,N_16044,N_15651);
nor U16603 (N_16603,N_15910,N_15602);
nor U16604 (N_16604,N_15925,N_16048);
or U16605 (N_16605,N_16134,N_15879);
nor U16606 (N_16606,N_16186,N_15804);
nor U16607 (N_16607,N_15808,N_15605);
and U16608 (N_16608,N_15844,N_15626);
nor U16609 (N_16609,N_15777,N_16185);
and U16610 (N_16610,N_15898,N_15705);
nand U16611 (N_16611,N_15638,N_15896);
and U16612 (N_16612,N_15777,N_16028);
xnor U16613 (N_16613,N_16034,N_15820);
nand U16614 (N_16614,N_16033,N_15764);
nand U16615 (N_16615,N_15989,N_15784);
or U16616 (N_16616,N_15728,N_15880);
xnor U16617 (N_16617,N_15628,N_16194);
or U16618 (N_16618,N_15703,N_15709);
nor U16619 (N_16619,N_15931,N_15839);
or U16620 (N_16620,N_15867,N_16132);
and U16621 (N_16621,N_15629,N_15600);
nand U16622 (N_16622,N_15787,N_16113);
and U16623 (N_16623,N_16061,N_16069);
or U16624 (N_16624,N_16146,N_16182);
nor U16625 (N_16625,N_16116,N_15802);
or U16626 (N_16626,N_16065,N_15747);
or U16627 (N_16627,N_15793,N_15945);
or U16628 (N_16628,N_15984,N_15982);
nand U16629 (N_16629,N_16009,N_15653);
nand U16630 (N_16630,N_16172,N_15643);
nand U16631 (N_16631,N_15669,N_15862);
nand U16632 (N_16632,N_16058,N_15678);
nor U16633 (N_16633,N_15905,N_16101);
nand U16634 (N_16634,N_15659,N_15767);
nor U16635 (N_16635,N_16024,N_15928);
nand U16636 (N_16636,N_15855,N_15944);
and U16637 (N_16637,N_16089,N_15868);
nand U16638 (N_16638,N_15990,N_15689);
nor U16639 (N_16639,N_16011,N_16088);
xnor U16640 (N_16640,N_16090,N_15939);
xnor U16641 (N_16641,N_15720,N_16089);
xnor U16642 (N_16642,N_15806,N_16065);
nand U16643 (N_16643,N_16164,N_15762);
or U16644 (N_16644,N_15754,N_16189);
or U16645 (N_16645,N_15789,N_16136);
and U16646 (N_16646,N_15798,N_16057);
nand U16647 (N_16647,N_15614,N_16185);
xnor U16648 (N_16648,N_15706,N_15675);
and U16649 (N_16649,N_15832,N_15980);
and U16650 (N_16650,N_15696,N_15781);
or U16651 (N_16651,N_15798,N_16172);
or U16652 (N_16652,N_15853,N_15893);
xnor U16653 (N_16653,N_15638,N_15822);
nor U16654 (N_16654,N_16184,N_16019);
or U16655 (N_16655,N_15608,N_16198);
nand U16656 (N_16656,N_16046,N_15636);
and U16657 (N_16657,N_15967,N_16066);
or U16658 (N_16658,N_15742,N_15889);
or U16659 (N_16659,N_15794,N_15725);
and U16660 (N_16660,N_15885,N_15918);
nor U16661 (N_16661,N_15942,N_15884);
or U16662 (N_16662,N_16193,N_15924);
xor U16663 (N_16663,N_15857,N_16106);
xnor U16664 (N_16664,N_15953,N_15651);
and U16665 (N_16665,N_15874,N_15791);
xor U16666 (N_16666,N_16144,N_16136);
and U16667 (N_16667,N_15964,N_16170);
or U16668 (N_16668,N_16081,N_16030);
or U16669 (N_16669,N_15952,N_15988);
nand U16670 (N_16670,N_15797,N_15899);
xor U16671 (N_16671,N_15652,N_15836);
nor U16672 (N_16672,N_15937,N_16141);
and U16673 (N_16673,N_15819,N_16128);
nand U16674 (N_16674,N_16181,N_15999);
and U16675 (N_16675,N_15765,N_16171);
or U16676 (N_16676,N_16194,N_16078);
nand U16677 (N_16677,N_15959,N_16059);
xnor U16678 (N_16678,N_16046,N_16092);
nand U16679 (N_16679,N_15939,N_15628);
or U16680 (N_16680,N_15673,N_15698);
or U16681 (N_16681,N_16070,N_16198);
and U16682 (N_16682,N_15605,N_16102);
and U16683 (N_16683,N_15724,N_15752);
or U16684 (N_16684,N_16100,N_15830);
or U16685 (N_16685,N_16143,N_15626);
xnor U16686 (N_16686,N_16036,N_15931);
and U16687 (N_16687,N_15859,N_15714);
and U16688 (N_16688,N_15782,N_15902);
nand U16689 (N_16689,N_16067,N_16178);
nand U16690 (N_16690,N_15891,N_15800);
or U16691 (N_16691,N_15734,N_16182);
nand U16692 (N_16692,N_15881,N_15770);
nand U16693 (N_16693,N_16020,N_15984);
nor U16694 (N_16694,N_15762,N_16095);
nand U16695 (N_16695,N_15832,N_15664);
and U16696 (N_16696,N_15724,N_16106);
nand U16697 (N_16697,N_16015,N_16083);
and U16698 (N_16698,N_16073,N_16194);
nor U16699 (N_16699,N_15609,N_16025);
and U16700 (N_16700,N_15835,N_15911);
and U16701 (N_16701,N_15739,N_15915);
or U16702 (N_16702,N_15761,N_15774);
or U16703 (N_16703,N_16179,N_15940);
nor U16704 (N_16704,N_16015,N_15762);
or U16705 (N_16705,N_15794,N_15669);
or U16706 (N_16706,N_15680,N_15726);
xor U16707 (N_16707,N_16145,N_15622);
or U16708 (N_16708,N_16039,N_16028);
or U16709 (N_16709,N_15718,N_15981);
xor U16710 (N_16710,N_16019,N_16003);
or U16711 (N_16711,N_16032,N_15972);
nand U16712 (N_16712,N_16057,N_15822);
and U16713 (N_16713,N_15848,N_15786);
xnor U16714 (N_16714,N_15740,N_16068);
nand U16715 (N_16715,N_15986,N_16181);
nor U16716 (N_16716,N_16139,N_16119);
nand U16717 (N_16717,N_15660,N_15740);
or U16718 (N_16718,N_16056,N_15611);
xnor U16719 (N_16719,N_16103,N_15997);
or U16720 (N_16720,N_15874,N_15987);
xor U16721 (N_16721,N_15690,N_15961);
nor U16722 (N_16722,N_15876,N_15846);
nor U16723 (N_16723,N_15802,N_15864);
nor U16724 (N_16724,N_16033,N_16037);
xnor U16725 (N_16725,N_16050,N_16008);
or U16726 (N_16726,N_16134,N_16146);
and U16727 (N_16727,N_15775,N_16077);
and U16728 (N_16728,N_16102,N_16049);
and U16729 (N_16729,N_16038,N_16027);
or U16730 (N_16730,N_16133,N_15830);
and U16731 (N_16731,N_15971,N_15662);
or U16732 (N_16732,N_16057,N_15884);
xor U16733 (N_16733,N_15794,N_15717);
nand U16734 (N_16734,N_16042,N_16047);
nand U16735 (N_16735,N_16016,N_15760);
or U16736 (N_16736,N_15785,N_16123);
nor U16737 (N_16737,N_16012,N_15678);
and U16738 (N_16738,N_16111,N_15900);
nand U16739 (N_16739,N_16055,N_16185);
or U16740 (N_16740,N_15729,N_15944);
or U16741 (N_16741,N_15896,N_15974);
nand U16742 (N_16742,N_15630,N_15678);
nor U16743 (N_16743,N_16042,N_15931);
nor U16744 (N_16744,N_15846,N_15616);
nand U16745 (N_16745,N_15705,N_15782);
nor U16746 (N_16746,N_15602,N_15622);
and U16747 (N_16747,N_16198,N_15883);
nor U16748 (N_16748,N_15969,N_15917);
nand U16749 (N_16749,N_15865,N_15833);
nand U16750 (N_16750,N_16137,N_15732);
xor U16751 (N_16751,N_15868,N_15628);
nor U16752 (N_16752,N_16047,N_16181);
nor U16753 (N_16753,N_16031,N_15811);
xor U16754 (N_16754,N_15654,N_16044);
xor U16755 (N_16755,N_16151,N_16096);
and U16756 (N_16756,N_15736,N_15929);
and U16757 (N_16757,N_16052,N_15825);
nor U16758 (N_16758,N_15932,N_15876);
or U16759 (N_16759,N_15712,N_16091);
or U16760 (N_16760,N_15850,N_15814);
and U16761 (N_16761,N_16156,N_15679);
xor U16762 (N_16762,N_15909,N_15679);
and U16763 (N_16763,N_16182,N_15917);
and U16764 (N_16764,N_15944,N_15758);
nor U16765 (N_16765,N_16146,N_15751);
xor U16766 (N_16766,N_15909,N_16023);
nand U16767 (N_16767,N_15958,N_16193);
xor U16768 (N_16768,N_15939,N_16113);
nand U16769 (N_16769,N_15634,N_15956);
and U16770 (N_16770,N_15886,N_15733);
nand U16771 (N_16771,N_15937,N_15629);
and U16772 (N_16772,N_15712,N_16129);
nand U16773 (N_16773,N_16188,N_15995);
or U16774 (N_16774,N_15774,N_15952);
and U16775 (N_16775,N_15762,N_15827);
or U16776 (N_16776,N_16043,N_16006);
and U16777 (N_16777,N_15641,N_15755);
or U16778 (N_16778,N_16078,N_15987);
xor U16779 (N_16779,N_16087,N_16052);
nand U16780 (N_16780,N_15732,N_15645);
nor U16781 (N_16781,N_15725,N_15743);
xnor U16782 (N_16782,N_16176,N_15701);
and U16783 (N_16783,N_15674,N_15623);
or U16784 (N_16784,N_15873,N_15974);
nor U16785 (N_16785,N_15717,N_15753);
nand U16786 (N_16786,N_15807,N_16010);
or U16787 (N_16787,N_15701,N_16036);
nor U16788 (N_16788,N_15920,N_15799);
nand U16789 (N_16789,N_15634,N_16109);
nand U16790 (N_16790,N_15654,N_15665);
and U16791 (N_16791,N_16118,N_16001);
nor U16792 (N_16792,N_16021,N_16141);
or U16793 (N_16793,N_16144,N_15792);
or U16794 (N_16794,N_15656,N_15774);
nand U16795 (N_16795,N_15876,N_15899);
nand U16796 (N_16796,N_16050,N_15801);
or U16797 (N_16797,N_15804,N_16057);
or U16798 (N_16798,N_15786,N_15677);
xnor U16799 (N_16799,N_16091,N_16028);
xor U16800 (N_16800,N_16233,N_16421);
and U16801 (N_16801,N_16296,N_16633);
or U16802 (N_16802,N_16265,N_16458);
or U16803 (N_16803,N_16485,N_16643);
nand U16804 (N_16804,N_16319,N_16362);
or U16805 (N_16805,N_16570,N_16466);
nor U16806 (N_16806,N_16252,N_16731);
or U16807 (N_16807,N_16390,N_16542);
nor U16808 (N_16808,N_16635,N_16738);
and U16809 (N_16809,N_16578,N_16728);
and U16810 (N_16810,N_16492,N_16436);
xnor U16811 (N_16811,N_16529,N_16447);
xnor U16812 (N_16812,N_16584,N_16257);
xnor U16813 (N_16813,N_16488,N_16781);
xnor U16814 (N_16814,N_16748,N_16678);
nor U16815 (N_16815,N_16750,N_16461);
nor U16816 (N_16816,N_16211,N_16293);
nand U16817 (N_16817,N_16330,N_16313);
xnor U16818 (N_16818,N_16783,N_16274);
nor U16819 (N_16819,N_16668,N_16673);
xnor U16820 (N_16820,N_16221,N_16577);
nor U16821 (N_16821,N_16796,N_16216);
nand U16822 (N_16822,N_16795,N_16652);
xnor U16823 (N_16823,N_16587,N_16444);
and U16824 (N_16824,N_16707,N_16380);
nand U16825 (N_16825,N_16660,N_16269);
or U16826 (N_16826,N_16766,N_16215);
xnor U16827 (N_16827,N_16217,N_16531);
nand U16828 (N_16828,N_16579,N_16688);
and U16829 (N_16829,N_16506,N_16454);
and U16830 (N_16830,N_16200,N_16307);
xnor U16831 (N_16831,N_16371,N_16516);
nand U16832 (N_16832,N_16367,N_16443);
xor U16833 (N_16833,N_16700,N_16694);
and U16834 (N_16834,N_16586,N_16223);
nand U16835 (N_16835,N_16758,N_16423);
and U16836 (N_16836,N_16705,N_16263);
xnor U16837 (N_16837,N_16589,N_16344);
nand U16838 (N_16838,N_16416,N_16247);
nand U16839 (N_16839,N_16358,N_16596);
nand U16840 (N_16840,N_16701,N_16314);
nor U16841 (N_16841,N_16225,N_16450);
or U16842 (N_16842,N_16222,N_16242);
nand U16843 (N_16843,N_16636,N_16679);
xnor U16844 (N_16844,N_16501,N_16267);
or U16845 (N_16845,N_16722,N_16662);
nor U16846 (N_16846,N_16602,N_16256);
nor U16847 (N_16847,N_16258,N_16550);
xor U16848 (N_16848,N_16718,N_16432);
nor U16849 (N_16849,N_16219,N_16630);
nor U16850 (N_16850,N_16312,N_16469);
or U16851 (N_16851,N_16512,N_16509);
nand U16852 (N_16852,N_16281,N_16743);
nor U16853 (N_16853,N_16655,N_16654);
and U16854 (N_16854,N_16212,N_16546);
or U16855 (N_16855,N_16321,N_16426);
nand U16856 (N_16856,N_16536,N_16207);
nor U16857 (N_16857,N_16645,N_16204);
xor U16858 (N_16858,N_16565,N_16382);
nand U16859 (N_16859,N_16505,N_16295);
xnor U16860 (N_16860,N_16272,N_16389);
nand U16861 (N_16861,N_16483,N_16490);
nor U16862 (N_16862,N_16710,N_16427);
nand U16863 (N_16863,N_16299,N_16276);
nor U16864 (N_16864,N_16661,N_16398);
and U16865 (N_16865,N_16677,N_16388);
nand U16866 (N_16866,N_16594,N_16761);
nor U16867 (N_16867,N_16338,N_16599);
or U16868 (N_16868,N_16580,N_16213);
and U16869 (N_16869,N_16764,N_16317);
xor U16870 (N_16870,N_16514,N_16508);
nor U16871 (N_16871,N_16463,N_16740);
xor U16872 (N_16872,N_16208,N_16775);
or U16873 (N_16873,N_16629,N_16537);
nor U16874 (N_16874,N_16395,N_16604);
nand U16875 (N_16875,N_16657,N_16591);
or U16876 (N_16876,N_16517,N_16359);
nand U16877 (N_16877,N_16521,N_16588);
nand U16878 (N_16878,N_16571,N_16266);
or U16879 (N_16879,N_16227,N_16741);
xnor U16880 (N_16880,N_16271,N_16736);
or U16881 (N_16881,N_16410,N_16702);
or U16882 (N_16882,N_16520,N_16791);
and U16883 (N_16883,N_16238,N_16639);
nor U16884 (N_16884,N_16511,N_16397);
xnor U16885 (N_16885,N_16291,N_16658);
nand U16886 (N_16886,N_16300,N_16343);
xnor U16887 (N_16887,N_16369,N_16502);
xnor U16888 (N_16888,N_16441,N_16309);
nand U16889 (N_16889,N_16699,N_16328);
nand U16890 (N_16890,N_16220,N_16471);
or U16891 (N_16891,N_16715,N_16228);
and U16892 (N_16892,N_16491,N_16592);
nor U16893 (N_16893,N_16459,N_16603);
nor U16894 (N_16894,N_16278,N_16341);
or U16895 (N_16895,N_16544,N_16434);
xor U16896 (N_16896,N_16757,N_16429);
xnor U16897 (N_16897,N_16575,N_16590);
and U16898 (N_16898,N_16393,N_16675);
nor U16899 (N_16899,N_16752,N_16595);
nor U16900 (N_16900,N_16452,N_16301);
or U16901 (N_16901,N_16535,N_16695);
xnor U16902 (N_16902,N_16704,N_16646);
nor U16903 (N_16903,N_16563,N_16448);
and U16904 (N_16904,N_16777,N_16782);
nor U16905 (N_16905,N_16440,N_16621);
or U16906 (N_16906,N_16373,N_16745);
nor U16907 (N_16907,N_16282,N_16486);
nand U16908 (N_16908,N_16318,N_16334);
and U16909 (N_16909,N_16431,N_16672);
nor U16910 (N_16910,N_16475,N_16402);
or U16911 (N_16911,N_16481,N_16375);
or U16912 (N_16912,N_16477,N_16774);
nor U16913 (N_16913,N_16335,N_16386);
or U16914 (N_16914,N_16494,N_16527);
nor U16915 (N_16915,N_16411,N_16457);
or U16916 (N_16916,N_16545,N_16433);
and U16917 (N_16917,N_16455,N_16598);
nand U16918 (N_16918,N_16769,N_16684);
nand U16919 (N_16919,N_16691,N_16472);
nand U16920 (N_16920,N_16790,N_16482);
nand U16921 (N_16921,N_16725,N_16532);
nor U16922 (N_16922,N_16609,N_16620);
nand U16923 (N_16923,N_16391,N_16756);
nor U16924 (N_16924,N_16418,N_16797);
nor U16925 (N_16925,N_16732,N_16417);
nor U16926 (N_16926,N_16350,N_16585);
nand U16927 (N_16927,N_16779,N_16408);
or U16928 (N_16928,N_16288,N_16496);
or U16929 (N_16929,N_16292,N_16352);
and U16930 (N_16930,N_16287,N_16364);
or U16931 (N_16931,N_16638,N_16489);
and U16932 (N_16932,N_16235,N_16414);
nor U16933 (N_16933,N_16248,N_16666);
and U16934 (N_16934,N_16538,N_16387);
nand U16935 (N_16935,N_16554,N_16474);
nor U16936 (N_16936,N_16768,N_16724);
nand U16937 (N_16937,N_16306,N_16415);
or U16938 (N_16938,N_16632,N_16453);
xor U16939 (N_16939,N_16360,N_16226);
nor U16940 (N_16940,N_16348,N_16403);
nand U16941 (N_16941,N_16607,N_16622);
and U16942 (N_16942,N_16689,N_16205);
nand U16943 (N_16943,N_16619,N_16559);
xor U16944 (N_16944,N_16776,N_16345);
xor U16945 (N_16945,N_16794,N_16412);
xnor U16946 (N_16946,N_16246,N_16273);
nor U16947 (N_16947,N_16232,N_16730);
xor U16948 (N_16948,N_16260,N_16760);
xnor U16949 (N_16949,N_16337,N_16717);
or U16950 (N_16950,N_16561,N_16703);
nand U16951 (N_16951,N_16647,N_16534);
and U16952 (N_16952,N_16612,N_16357);
nor U16953 (N_16953,N_16262,N_16480);
nor U16954 (N_16954,N_16720,N_16290);
xor U16955 (N_16955,N_16302,N_16366);
nor U16956 (N_16956,N_16311,N_16582);
nor U16957 (N_16957,N_16356,N_16210);
and U16958 (N_16958,N_16283,N_16404);
nand U16959 (N_16959,N_16510,N_16464);
nand U16960 (N_16960,N_16353,N_16614);
or U16961 (N_16961,N_16692,N_16513);
or U16962 (N_16962,N_16653,N_16413);
xnor U16963 (N_16963,N_16754,N_16249);
nand U16964 (N_16964,N_16789,N_16451);
and U16965 (N_16965,N_16493,N_16326);
or U16966 (N_16966,N_16530,N_16294);
or U16967 (N_16967,N_16478,N_16385);
or U16968 (N_16968,N_16342,N_16784);
or U16969 (N_16969,N_16304,N_16785);
xnor U16970 (N_16970,N_16244,N_16522);
or U16971 (N_16971,N_16566,N_16445);
nor U16972 (N_16972,N_16548,N_16374);
nand U16973 (N_16973,N_16659,N_16470);
and U16974 (N_16974,N_16771,N_16551);
xnor U16975 (N_16975,N_16558,N_16568);
xnor U16976 (N_16976,N_16723,N_16394);
nor U16977 (N_16977,N_16325,N_16420);
nand U16978 (N_16978,N_16329,N_16682);
or U16979 (N_16979,N_16495,N_16648);
xnor U16980 (N_16980,N_16687,N_16484);
nor U16981 (N_16981,N_16255,N_16799);
nor U16982 (N_16982,N_16401,N_16770);
xnor U16983 (N_16983,N_16327,N_16460);
nand U16984 (N_16984,N_16378,N_16528);
nand U16985 (N_16985,N_16241,N_16788);
or U16986 (N_16986,N_16683,N_16355);
nor U16987 (N_16987,N_16270,N_16605);
and U16988 (N_16988,N_16547,N_16368);
nand U16989 (N_16989,N_16405,N_16279);
and U16990 (N_16990,N_16676,N_16234);
nor U16991 (N_16991,N_16322,N_16541);
and U16992 (N_16992,N_16618,N_16525);
xor U16993 (N_16993,N_16556,N_16613);
nor U16994 (N_16994,N_16515,N_16231);
nor U16995 (N_16995,N_16384,N_16600);
and U16996 (N_16996,N_16383,N_16798);
or U16997 (N_16997,N_16762,N_16737);
or U16998 (N_16998,N_16610,N_16706);
and U16999 (N_16999,N_16560,N_16634);
and U17000 (N_17000,N_16669,N_16202);
and U17001 (N_17001,N_16637,N_16372);
nor U17002 (N_17002,N_16310,N_16712);
nand U17003 (N_17003,N_16719,N_16331);
xnor U17004 (N_17004,N_16435,N_16365);
or U17005 (N_17005,N_16336,N_16749);
xor U17006 (N_17006,N_16721,N_16376);
nor U17007 (N_17007,N_16209,N_16349);
nor U17008 (N_17008,N_16778,N_16780);
or U17009 (N_17009,N_16697,N_16539);
nor U17010 (N_17010,N_16562,N_16742);
and U17011 (N_17011,N_16351,N_16713);
xor U17012 (N_17012,N_16456,N_16438);
nand U17013 (N_17013,N_16280,N_16214);
nor U17014 (N_17014,N_16277,N_16264);
nand U17015 (N_17015,N_16409,N_16773);
and U17016 (N_17016,N_16323,N_16229);
nand U17017 (N_17017,N_16564,N_16693);
nand U17018 (N_17018,N_16370,N_16739);
nor U17019 (N_17019,N_16354,N_16716);
nand U17020 (N_17020,N_16674,N_16419);
nand U17021 (N_17021,N_16465,N_16504);
nor U17022 (N_17022,N_16245,N_16623);
nor U17023 (N_17023,N_16667,N_16543);
nand U17024 (N_17024,N_16468,N_16201);
and U17025 (N_17025,N_16361,N_16206);
nor U17026 (N_17026,N_16597,N_16316);
or U17027 (N_17027,N_16787,N_16726);
nor U17028 (N_17028,N_16497,N_16526);
and U17029 (N_17029,N_16500,N_16611);
nand U17030 (N_17030,N_16347,N_16430);
nand U17031 (N_17031,N_16399,N_16698);
nand U17032 (N_17032,N_16243,N_16651);
and U17033 (N_17033,N_16519,N_16237);
and U17034 (N_17034,N_16549,N_16407);
and U17035 (N_17035,N_16583,N_16553);
and U17036 (N_17036,N_16203,N_16400);
and U17037 (N_17037,N_16381,N_16346);
or U17038 (N_17038,N_16332,N_16767);
and U17039 (N_17039,N_16751,N_16744);
nor U17040 (N_17040,N_16308,N_16625);
nand U17041 (N_17041,N_16286,N_16406);
xor U17042 (N_17042,N_16642,N_16428);
nand U17043 (N_17043,N_16572,N_16424);
and U17044 (N_17044,N_16616,N_16425);
and U17045 (N_17045,N_16576,N_16218);
xor U17046 (N_17046,N_16696,N_16251);
or U17047 (N_17047,N_16467,N_16650);
xnor U17048 (N_17048,N_16442,N_16533);
nand U17049 (N_17049,N_16268,N_16253);
or U17050 (N_17050,N_16747,N_16680);
nor U17051 (N_17051,N_16462,N_16734);
or U17052 (N_17052,N_16567,N_16649);
xor U17053 (N_17053,N_16714,N_16540);
nand U17054 (N_17054,N_16601,N_16297);
nand U17055 (N_17055,N_16446,N_16615);
and U17056 (N_17056,N_16690,N_16664);
and U17057 (N_17057,N_16727,N_16765);
xor U17058 (N_17058,N_16320,N_16628);
xnor U17059 (N_17059,N_16665,N_16275);
xor U17060 (N_17060,N_16507,N_16670);
and U17061 (N_17061,N_16340,N_16640);
nor U17062 (N_17062,N_16641,N_16606);
nor U17063 (N_17063,N_16593,N_16735);
nand U17064 (N_17064,N_16333,N_16303);
and U17065 (N_17065,N_16499,N_16631);
and U17066 (N_17066,N_16259,N_16671);
and U17067 (N_17067,N_16437,N_16644);
nor U17068 (N_17068,N_16759,N_16236);
nor U17069 (N_17069,N_16284,N_16753);
xor U17070 (N_17070,N_16254,N_16224);
and U17071 (N_17071,N_16503,N_16763);
or U17072 (N_17072,N_16557,N_16627);
nor U17073 (N_17073,N_16498,N_16379);
nand U17074 (N_17074,N_16681,N_16772);
or U17075 (N_17075,N_16523,N_16392);
and U17076 (N_17076,N_16608,N_16298);
or U17077 (N_17077,N_16240,N_16479);
xor U17078 (N_17078,N_16377,N_16487);
nand U17079 (N_17079,N_16574,N_16261);
nor U17080 (N_17080,N_16555,N_16786);
nand U17081 (N_17081,N_16573,N_16729);
or U17082 (N_17082,N_16339,N_16755);
xor U17083 (N_17083,N_16363,N_16422);
nand U17084 (N_17084,N_16746,N_16708);
or U17085 (N_17085,N_16289,N_16518);
nor U17086 (N_17086,N_16396,N_16324);
xor U17087 (N_17087,N_16285,N_16663);
nor U17088 (N_17088,N_16476,N_16230);
xnor U17089 (N_17089,N_16624,N_16569);
nor U17090 (N_17090,N_16792,N_16250);
nand U17091 (N_17091,N_16315,N_16626);
xnor U17092 (N_17092,N_16581,N_16524);
and U17093 (N_17093,N_16449,N_16656);
xor U17094 (N_17094,N_16305,N_16709);
nor U17095 (N_17095,N_16473,N_16439);
or U17096 (N_17096,N_16686,N_16711);
nor U17097 (N_17097,N_16733,N_16239);
nor U17098 (N_17098,N_16793,N_16552);
nor U17099 (N_17099,N_16617,N_16685);
xor U17100 (N_17100,N_16642,N_16462);
and U17101 (N_17101,N_16553,N_16282);
nand U17102 (N_17102,N_16505,N_16434);
and U17103 (N_17103,N_16246,N_16733);
and U17104 (N_17104,N_16755,N_16430);
or U17105 (N_17105,N_16273,N_16773);
nor U17106 (N_17106,N_16250,N_16781);
or U17107 (N_17107,N_16575,N_16371);
nand U17108 (N_17108,N_16654,N_16390);
nor U17109 (N_17109,N_16368,N_16406);
or U17110 (N_17110,N_16786,N_16683);
or U17111 (N_17111,N_16352,N_16624);
nor U17112 (N_17112,N_16201,N_16297);
or U17113 (N_17113,N_16672,N_16382);
xor U17114 (N_17114,N_16497,N_16471);
nand U17115 (N_17115,N_16684,N_16213);
xor U17116 (N_17116,N_16526,N_16368);
and U17117 (N_17117,N_16516,N_16365);
xor U17118 (N_17118,N_16203,N_16240);
and U17119 (N_17119,N_16253,N_16251);
or U17120 (N_17120,N_16322,N_16782);
nand U17121 (N_17121,N_16564,N_16647);
or U17122 (N_17122,N_16729,N_16363);
nor U17123 (N_17123,N_16391,N_16463);
and U17124 (N_17124,N_16357,N_16283);
nand U17125 (N_17125,N_16543,N_16518);
nand U17126 (N_17126,N_16319,N_16664);
and U17127 (N_17127,N_16496,N_16342);
or U17128 (N_17128,N_16227,N_16682);
and U17129 (N_17129,N_16271,N_16546);
nor U17130 (N_17130,N_16733,N_16625);
and U17131 (N_17131,N_16684,N_16427);
or U17132 (N_17132,N_16649,N_16600);
nand U17133 (N_17133,N_16609,N_16488);
and U17134 (N_17134,N_16426,N_16658);
xnor U17135 (N_17135,N_16230,N_16767);
xnor U17136 (N_17136,N_16255,N_16541);
or U17137 (N_17137,N_16439,N_16278);
or U17138 (N_17138,N_16459,N_16780);
and U17139 (N_17139,N_16451,N_16664);
nor U17140 (N_17140,N_16268,N_16488);
xnor U17141 (N_17141,N_16253,N_16346);
nand U17142 (N_17142,N_16408,N_16751);
nor U17143 (N_17143,N_16351,N_16275);
xor U17144 (N_17144,N_16614,N_16277);
nand U17145 (N_17145,N_16705,N_16405);
xor U17146 (N_17146,N_16444,N_16204);
nor U17147 (N_17147,N_16714,N_16273);
nor U17148 (N_17148,N_16510,N_16444);
or U17149 (N_17149,N_16712,N_16521);
or U17150 (N_17150,N_16690,N_16622);
nand U17151 (N_17151,N_16718,N_16736);
nand U17152 (N_17152,N_16278,N_16464);
or U17153 (N_17153,N_16791,N_16655);
and U17154 (N_17154,N_16667,N_16356);
and U17155 (N_17155,N_16787,N_16294);
and U17156 (N_17156,N_16792,N_16467);
nor U17157 (N_17157,N_16233,N_16658);
nand U17158 (N_17158,N_16585,N_16471);
nor U17159 (N_17159,N_16590,N_16344);
nor U17160 (N_17160,N_16554,N_16750);
and U17161 (N_17161,N_16695,N_16665);
xor U17162 (N_17162,N_16694,N_16240);
xnor U17163 (N_17163,N_16227,N_16214);
and U17164 (N_17164,N_16265,N_16370);
nor U17165 (N_17165,N_16239,N_16289);
or U17166 (N_17166,N_16781,N_16304);
and U17167 (N_17167,N_16636,N_16499);
nand U17168 (N_17168,N_16421,N_16417);
nand U17169 (N_17169,N_16426,N_16732);
nor U17170 (N_17170,N_16581,N_16247);
nand U17171 (N_17171,N_16345,N_16411);
and U17172 (N_17172,N_16529,N_16355);
and U17173 (N_17173,N_16328,N_16236);
nor U17174 (N_17174,N_16253,N_16273);
nor U17175 (N_17175,N_16743,N_16557);
nand U17176 (N_17176,N_16270,N_16496);
nand U17177 (N_17177,N_16229,N_16781);
or U17178 (N_17178,N_16755,N_16749);
or U17179 (N_17179,N_16612,N_16758);
xnor U17180 (N_17180,N_16420,N_16268);
nor U17181 (N_17181,N_16481,N_16518);
or U17182 (N_17182,N_16218,N_16461);
xnor U17183 (N_17183,N_16378,N_16741);
nor U17184 (N_17184,N_16254,N_16482);
xnor U17185 (N_17185,N_16784,N_16261);
or U17186 (N_17186,N_16669,N_16373);
and U17187 (N_17187,N_16269,N_16795);
nor U17188 (N_17188,N_16322,N_16256);
and U17189 (N_17189,N_16720,N_16331);
nor U17190 (N_17190,N_16684,N_16395);
and U17191 (N_17191,N_16645,N_16526);
nand U17192 (N_17192,N_16459,N_16408);
and U17193 (N_17193,N_16461,N_16795);
and U17194 (N_17194,N_16612,N_16558);
and U17195 (N_17195,N_16685,N_16208);
nor U17196 (N_17196,N_16244,N_16352);
and U17197 (N_17197,N_16486,N_16307);
and U17198 (N_17198,N_16313,N_16439);
and U17199 (N_17199,N_16261,N_16686);
nand U17200 (N_17200,N_16230,N_16602);
nand U17201 (N_17201,N_16694,N_16547);
xnor U17202 (N_17202,N_16370,N_16423);
or U17203 (N_17203,N_16373,N_16618);
nor U17204 (N_17204,N_16612,N_16506);
nand U17205 (N_17205,N_16264,N_16350);
or U17206 (N_17206,N_16316,N_16273);
nor U17207 (N_17207,N_16409,N_16366);
nand U17208 (N_17208,N_16346,N_16772);
xnor U17209 (N_17209,N_16710,N_16749);
nor U17210 (N_17210,N_16671,N_16510);
and U17211 (N_17211,N_16570,N_16419);
and U17212 (N_17212,N_16599,N_16735);
and U17213 (N_17213,N_16700,N_16360);
xor U17214 (N_17214,N_16276,N_16438);
nand U17215 (N_17215,N_16549,N_16787);
or U17216 (N_17216,N_16715,N_16632);
xor U17217 (N_17217,N_16568,N_16538);
or U17218 (N_17218,N_16237,N_16238);
or U17219 (N_17219,N_16338,N_16283);
or U17220 (N_17220,N_16319,N_16580);
xor U17221 (N_17221,N_16646,N_16490);
xnor U17222 (N_17222,N_16715,N_16592);
nor U17223 (N_17223,N_16262,N_16777);
xnor U17224 (N_17224,N_16647,N_16259);
nand U17225 (N_17225,N_16529,N_16569);
xor U17226 (N_17226,N_16752,N_16508);
xnor U17227 (N_17227,N_16759,N_16573);
nor U17228 (N_17228,N_16476,N_16604);
and U17229 (N_17229,N_16466,N_16796);
nand U17230 (N_17230,N_16456,N_16689);
or U17231 (N_17231,N_16524,N_16211);
or U17232 (N_17232,N_16503,N_16759);
xnor U17233 (N_17233,N_16544,N_16427);
nor U17234 (N_17234,N_16234,N_16765);
nand U17235 (N_17235,N_16503,N_16500);
and U17236 (N_17236,N_16485,N_16791);
xor U17237 (N_17237,N_16285,N_16464);
and U17238 (N_17238,N_16548,N_16537);
xnor U17239 (N_17239,N_16615,N_16381);
nor U17240 (N_17240,N_16687,N_16204);
nor U17241 (N_17241,N_16294,N_16409);
or U17242 (N_17242,N_16337,N_16529);
nand U17243 (N_17243,N_16738,N_16669);
xor U17244 (N_17244,N_16241,N_16756);
or U17245 (N_17245,N_16444,N_16550);
and U17246 (N_17246,N_16222,N_16203);
xor U17247 (N_17247,N_16289,N_16406);
xor U17248 (N_17248,N_16430,N_16655);
or U17249 (N_17249,N_16644,N_16399);
nor U17250 (N_17250,N_16758,N_16742);
or U17251 (N_17251,N_16690,N_16225);
and U17252 (N_17252,N_16235,N_16467);
nor U17253 (N_17253,N_16679,N_16742);
nand U17254 (N_17254,N_16229,N_16514);
xor U17255 (N_17255,N_16531,N_16246);
and U17256 (N_17256,N_16359,N_16640);
xnor U17257 (N_17257,N_16627,N_16550);
or U17258 (N_17258,N_16238,N_16755);
xor U17259 (N_17259,N_16656,N_16209);
xor U17260 (N_17260,N_16659,N_16244);
or U17261 (N_17261,N_16450,N_16496);
or U17262 (N_17262,N_16738,N_16397);
or U17263 (N_17263,N_16240,N_16211);
or U17264 (N_17264,N_16558,N_16746);
xnor U17265 (N_17265,N_16604,N_16523);
and U17266 (N_17266,N_16566,N_16499);
nor U17267 (N_17267,N_16769,N_16210);
xnor U17268 (N_17268,N_16220,N_16544);
nor U17269 (N_17269,N_16228,N_16684);
xor U17270 (N_17270,N_16759,N_16310);
or U17271 (N_17271,N_16394,N_16330);
xor U17272 (N_17272,N_16788,N_16676);
and U17273 (N_17273,N_16649,N_16469);
nand U17274 (N_17274,N_16212,N_16469);
and U17275 (N_17275,N_16469,N_16720);
nor U17276 (N_17276,N_16375,N_16716);
or U17277 (N_17277,N_16451,N_16652);
xnor U17278 (N_17278,N_16474,N_16484);
or U17279 (N_17279,N_16544,N_16678);
nor U17280 (N_17280,N_16254,N_16452);
nand U17281 (N_17281,N_16634,N_16707);
nand U17282 (N_17282,N_16297,N_16797);
nand U17283 (N_17283,N_16693,N_16660);
and U17284 (N_17284,N_16306,N_16590);
or U17285 (N_17285,N_16510,N_16602);
or U17286 (N_17286,N_16275,N_16458);
nand U17287 (N_17287,N_16258,N_16335);
xnor U17288 (N_17288,N_16463,N_16620);
or U17289 (N_17289,N_16497,N_16708);
or U17290 (N_17290,N_16710,N_16203);
nor U17291 (N_17291,N_16630,N_16740);
and U17292 (N_17292,N_16251,N_16454);
or U17293 (N_17293,N_16299,N_16494);
or U17294 (N_17294,N_16717,N_16243);
nor U17295 (N_17295,N_16523,N_16638);
and U17296 (N_17296,N_16205,N_16244);
xor U17297 (N_17297,N_16392,N_16616);
nand U17298 (N_17298,N_16558,N_16737);
nor U17299 (N_17299,N_16545,N_16445);
xnor U17300 (N_17300,N_16511,N_16316);
and U17301 (N_17301,N_16484,N_16489);
nor U17302 (N_17302,N_16654,N_16511);
nor U17303 (N_17303,N_16747,N_16429);
and U17304 (N_17304,N_16442,N_16673);
nand U17305 (N_17305,N_16638,N_16659);
nand U17306 (N_17306,N_16380,N_16433);
and U17307 (N_17307,N_16467,N_16290);
and U17308 (N_17308,N_16406,N_16283);
nor U17309 (N_17309,N_16720,N_16584);
and U17310 (N_17310,N_16350,N_16640);
nor U17311 (N_17311,N_16732,N_16610);
xnor U17312 (N_17312,N_16604,N_16769);
and U17313 (N_17313,N_16574,N_16313);
and U17314 (N_17314,N_16619,N_16319);
xor U17315 (N_17315,N_16725,N_16358);
or U17316 (N_17316,N_16422,N_16684);
and U17317 (N_17317,N_16202,N_16323);
nand U17318 (N_17318,N_16220,N_16708);
and U17319 (N_17319,N_16483,N_16656);
nand U17320 (N_17320,N_16621,N_16384);
and U17321 (N_17321,N_16412,N_16629);
nand U17322 (N_17322,N_16551,N_16689);
nor U17323 (N_17323,N_16394,N_16562);
nand U17324 (N_17324,N_16643,N_16448);
and U17325 (N_17325,N_16770,N_16684);
xnor U17326 (N_17326,N_16349,N_16656);
xnor U17327 (N_17327,N_16246,N_16419);
or U17328 (N_17328,N_16218,N_16266);
nand U17329 (N_17329,N_16734,N_16315);
and U17330 (N_17330,N_16391,N_16797);
nand U17331 (N_17331,N_16518,N_16488);
and U17332 (N_17332,N_16233,N_16454);
xor U17333 (N_17333,N_16603,N_16618);
xor U17334 (N_17334,N_16222,N_16615);
nor U17335 (N_17335,N_16281,N_16516);
and U17336 (N_17336,N_16782,N_16743);
and U17337 (N_17337,N_16256,N_16794);
nand U17338 (N_17338,N_16397,N_16657);
nand U17339 (N_17339,N_16294,N_16476);
or U17340 (N_17340,N_16532,N_16739);
and U17341 (N_17341,N_16338,N_16534);
nand U17342 (N_17342,N_16483,N_16678);
or U17343 (N_17343,N_16526,N_16253);
or U17344 (N_17344,N_16324,N_16737);
nand U17345 (N_17345,N_16751,N_16657);
nand U17346 (N_17346,N_16745,N_16551);
xnor U17347 (N_17347,N_16467,N_16316);
xnor U17348 (N_17348,N_16327,N_16749);
nand U17349 (N_17349,N_16503,N_16687);
nor U17350 (N_17350,N_16647,N_16630);
and U17351 (N_17351,N_16398,N_16633);
nand U17352 (N_17352,N_16575,N_16283);
nor U17353 (N_17353,N_16466,N_16701);
and U17354 (N_17354,N_16514,N_16577);
or U17355 (N_17355,N_16209,N_16479);
xor U17356 (N_17356,N_16457,N_16779);
and U17357 (N_17357,N_16619,N_16454);
nand U17358 (N_17358,N_16664,N_16454);
and U17359 (N_17359,N_16749,N_16709);
nor U17360 (N_17360,N_16747,N_16273);
and U17361 (N_17361,N_16367,N_16620);
xnor U17362 (N_17362,N_16305,N_16276);
nand U17363 (N_17363,N_16254,N_16551);
and U17364 (N_17364,N_16731,N_16432);
or U17365 (N_17365,N_16286,N_16649);
nor U17366 (N_17366,N_16660,N_16485);
xor U17367 (N_17367,N_16581,N_16518);
or U17368 (N_17368,N_16272,N_16766);
or U17369 (N_17369,N_16268,N_16660);
or U17370 (N_17370,N_16420,N_16650);
and U17371 (N_17371,N_16459,N_16425);
xnor U17372 (N_17372,N_16310,N_16677);
xor U17373 (N_17373,N_16442,N_16457);
and U17374 (N_17374,N_16589,N_16503);
nor U17375 (N_17375,N_16401,N_16604);
xor U17376 (N_17376,N_16544,N_16324);
xor U17377 (N_17377,N_16201,N_16544);
nor U17378 (N_17378,N_16429,N_16624);
xor U17379 (N_17379,N_16219,N_16627);
xor U17380 (N_17380,N_16325,N_16700);
or U17381 (N_17381,N_16462,N_16287);
nor U17382 (N_17382,N_16308,N_16347);
and U17383 (N_17383,N_16235,N_16413);
xnor U17384 (N_17384,N_16290,N_16629);
and U17385 (N_17385,N_16497,N_16447);
and U17386 (N_17386,N_16619,N_16754);
xor U17387 (N_17387,N_16511,N_16268);
xnor U17388 (N_17388,N_16786,N_16690);
or U17389 (N_17389,N_16658,N_16574);
nor U17390 (N_17390,N_16524,N_16543);
or U17391 (N_17391,N_16247,N_16587);
and U17392 (N_17392,N_16294,N_16773);
and U17393 (N_17393,N_16354,N_16576);
nand U17394 (N_17394,N_16400,N_16700);
xnor U17395 (N_17395,N_16459,N_16479);
nor U17396 (N_17396,N_16748,N_16469);
nand U17397 (N_17397,N_16425,N_16635);
nor U17398 (N_17398,N_16417,N_16253);
xor U17399 (N_17399,N_16502,N_16230);
xnor U17400 (N_17400,N_17029,N_17264);
or U17401 (N_17401,N_17142,N_17135);
xor U17402 (N_17402,N_16987,N_16824);
nor U17403 (N_17403,N_17148,N_16819);
xnor U17404 (N_17404,N_16812,N_17388);
nand U17405 (N_17405,N_16905,N_17201);
and U17406 (N_17406,N_17047,N_16829);
nand U17407 (N_17407,N_17321,N_17012);
nor U17408 (N_17408,N_16914,N_16831);
nand U17409 (N_17409,N_17111,N_16965);
and U17410 (N_17410,N_16944,N_17107);
or U17411 (N_17411,N_17376,N_17244);
nand U17412 (N_17412,N_16877,N_17338);
nand U17413 (N_17413,N_17102,N_17282);
or U17414 (N_17414,N_17302,N_17105);
nand U17415 (N_17415,N_17290,N_17381);
nand U17416 (N_17416,N_17075,N_17076);
or U17417 (N_17417,N_17339,N_16936);
nor U17418 (N_17418,N_17344,N_17089);
and U17419 (N_17419,N_16932,N_17232);
nand U17420 (N_17420,N_16814,N_17250);
or U17421 (N_17421,N_17136,N_17320);
and U17422 (N_17422,N_16955,N_17168);
and U17423 (N_17423,N_17228,N_16993);
xor U17424 (N_17424,N_17134,N_16890);
nor U17425 (N_17425,N_17020,N_16870);
or U17426 (N_17426,N_17078,N_16985);
nand U17427 (N_17427,N_16970,N_16866);
nand U17428 (N_17428,N_17038,N_17373);
nor U17429 (N_17429,N_16809,N_17096);
and U17430 (N_17430,N_17298,N_17055);
nand U17431 (N_17431,N_17045,N_17097);
xnor U17432 (N_17432,N_17043,N_17115);
and U17433 (N_17433,N_17188,N_16802);
and U17434 (N_17434,N_16975,N_16826);
nor U17435 (N_17435,N_16810,N_16891);
nand U17436 (N_17436,N_16920,N_16859);
nand U17437 (N_17437,N_17066,N_17145);
nand U17438 (N_17438,N_17184,N_17313);
or U17439 (N_17439,N_17162,N_17391);
and U17440 (N_17440,N_16839,N_17117);
and U17441 (N_17441,N_17347,N_16842);
xor U17442 (N_17442,N_16878,N_16899);
nor U17443 (N_17443,N_17167,N_17099);
or U17444 (N_17444,N_16855,N_17031);
nor U17445 (N_17445,N_16811,N_17340);
xnor U17446 (N_17446,N_16848,N_17174);
nand U17447 (N_17447,N_17316,N_17077);
and U17448 (N_17448,N_17377,N_17063);
xor U17449 (N_17449,N_17072,N_17243);
xor U17450 (N_17450,N_17348,N_16933);
or U17451 (N_17451,N_17143,N_17017);
xor U17452 (N_17452,N_16942,N_16908);
nor U17453 (N_17453,N_17199,N_16919);
nor U17454 (N_17454,N_16983,N_16903);
or U17455 (N_17455,N_17194,N_16994);
xor U17456 (N_17456,N_17227,N_17110);
nor U17457 (N_17457,N_17274,N_17137);
xnor U17458 (N_17458,N_17292,N_17157);
nor U17459 (N_17459,N_16925,N_17113);
xor U17460 (N_17460,N_17385,N_17094);
or U17461 (N_17461,N_17218,N_17050);
xnor U17462 (N_17462,N_17205,N_16872);
or U17463 (N_17463,N_16897,N_17006);
and U17464 (N_17464,N_17281,N_17119);
nor U17465 (N_17465,N_17091,N_17314);
nand U17466 (N_17466,N_16882,N_17396);
or U17467 (N_17467,N_17270,N_17237);
or U17468 (N_17468,N_17248,N_17288);
xor U17469 (N_17469,N_16885,N_16845);
nor U17470 (N_17470,N_17158,N_16883);
nand U17471 (N_17471,N_17088,N_17395);
nand U17472 (N_17472,N_16963,N_17343);
and U17473 (N_17473,N_16873,N_17152);
nand U17474 (N_17474,N_17127,N_17027);
or U17475 (N_17475,N_17331,N_17086);
nor U17476 (N_17476,N_16834,N_17071);
nand U17477 (N_17477,N_16896,N_17176);
and U17478 (N_17478,N_17390,N_17258);
or U17479 (N_17479,N_17289,N_17009);
or U17480 (N_17480,N_17397,N_17095);
xnor U17481 (N_17481,N_17106,N_17165);
and U17482 (N_17482,N_17333,N_16957);
and U17483 (N_17483,N_17297,N_17062);
and U17484 (N_17484,N_17216,N_17399);
nor U17485 (N_17485,N_17280,N_17122);
xnor U17486 (N_17486,N_17175,N_17190);
or U17487 (N_17487,N_16945,N_17295);
or U17488 (N_17488,N_17335,N_17353);
or U17489 (N_17489,N_16887,N_17032);
nand U17490 (N_17490,N_16913,N_16941);
xnor U17491 (N_17491,N_17285,N_17254);
and U17492 (N_17492,N_17120,N_17308);
or U17493 (N_17493,N_17370,N_17360);
nand U17494 (N_17494,N_17182,N_16871);
or U17495 (N_17495,N_17170,N_16888);
nand U17496 (N_17496,N_17155,N_17123);
nand U17497 (N_17497,N_16803,N_17271);
nand U17498 (N_17498,N_17317,N_17256);
nor U17499 (N_17499,N_17196,N_16923);
or U17500 (N_17500,N_17132,N_16968);
or U17501 (N_17501,N_17200,N_17212);
or U17502 (N_17502,N_16835,N_17178);
xor U17503 (N_17503,N_17255,N_17073);
or U17504 (N_17504,N_17061,N_17337);
xnor U17505 (N_17505,N_17366,N_17181);
or U17506 (N_17506,N_17156,N_16931);
xnor U17507 (N_17507,N_17206,N_17296);
or U17508 (N_17508,N_16951,N_17007);
or U17509 (N_17509,N_17394,N_16969);
or U17510 (N_17510,N_17124,N_16962);
nand U17511 (N_17511,N_16850,N_17275);
nand U17512 (N_17512,N_17363,N_16998);
nor U17513 (N_17513,N_16840,N_17064);
or U17514 (N_17514,N_17149,N_16833);
xor U17515 (N_17515,N_17056,N_17018);
nor U17516 (N_17516,N_17386,N_16876);
nand U17517 (N_17517,N_17269,N_17019);
or U17518 (N_17518,N_17005,N_17249);
and U17519 (N_17519,N_17309,N_17217);
and U17520 (N_17520,N_16906,N_17189);
nor U17521 (N_17521,N_16889,N_17101);
nor U17522 (N_17522,N_17334,N_16867);
nand U17523 (N_17523,N_17085,N_17058);
or U17524 (N_17524,N_16982,N_16857);
or U17525 (N_17525,N_16961,N_16822);
xor U17526 (N_17526,N_17215,N_16804);
xor U17527 (N_17527,N_17070,N_17221);
nor U17528 (N_17528,N_17352,N_17059);
xnor U17529 (N_17529,N_17235,N_16830);
or U17530 (N_17530,N_17312,N_17131);
xor U17531 (N_17531,N_17355,N_16940);
xor U17532 (N_17532,N_17367,N_17021);
or U17533 (N_17533,N_17204,N_17109);
xnor U17534 (N_17534,N_16981,N_16821);
and U17535 (N_17535,N_16817,N_17185);
and U17536 (N_17536,N_17116,N_16916);
nor U17537 (N_17537,N_17261,N_17192);
and U17538 (N_17538,N_16907,N_16984);
xnor U17539 (N_17539,N_16960,N_17171);
and U17540 (N_17540,N_16991,N_17263);
or U17541 (N_17541,N_17041,N_16861);
nand U17542 (N_17542,N_17267,N_17311);
or U17543 (N_17543,N_17371,N_16881);
nand U17544 (N_17544,N_16828,N_17051);
xor U17545 (N_17545,N_17329,N_17266);
and U17546 (N_17546,N_17209,N_17207);
nor U17547 (N_17547,N_17379,N_17246);
nor U17548 (N_17548,N_17186,N_17208);
nor U17549 (N_17549,N_16844,N_17052);
nand U17550 (N_17550,N_17144,N_17392);
nand U17551 (N_17551,N_16875,N_17037);
or U17552 (N_17552,N_17090,N_17084);
xnor U17553 (N_17553,N_16990,N_17277);
nor U17554 (N_17554,N_16823,N_17008);
nand U17555 (N_17555,N_16912,N_16851);
nor U17556 (N_17556,N_17251,N_17383);
xor U17557 (N_17557,N_16849,N_17068);
nor U17558 (N_17558,N_17387,N_17389);
xor U17559 (N_17559,N_16926,N_16928);
nor U17560 (N_17560,N_17327,N_17108);
nand U17561 (N_17561,N_17214,N_17030);
or U17562 (N_17562,N_17129,N_16939);
nor U17563 (N_17563,N_16930,N_16806);
and U17564 (N_17564,N_17042,N_17154);
or U17565 (N_17565,N_16924,N_17159);
or U17566 (N_17566,N_17028,N_17300);
nand U17567 (N_17567,N_17166,N_17160);
or U17568 (N_17568,N_17163,N_17053);
or U17569 (N_17569,N_16902,N_17346);
or U17570 (N_17570,N_17103,N_17294);
or U17571 (N_17571,N_17093,N_17252);
xor U17572 (N_17572,N_16986,N_17060);
xnor U17573 (N_17573,N_17040,N_16852);
or U17574 (N_17574,N_17336,N_16911);
nand U17575 (N_17575,N_17210,N_17358);
or U17576 (N_17576,N_17265,N_17293);
and U17577 (N_17577,N_17310,N_16800);
nor U17578 (N_17578,N_16973,N_16825);
xnor U17579 (N_17579,N_17326,N_17024);
or U17580 (N_17580,N_16838,N_17324);
nand U17581 (N_17581,N_16854,N_16900);
or U17582 (N_17582,N_17140,N_17372);
and U17583 (N_17583,N_17253,N_17225);
or U17584 (N_17584,N_17325,N_17234);
nor U17585 (N_17585,N_16915,N_16937);
nand U17586 (N_17586,N_16884,N_17150);
or U17587 (N_17587,N_17044,N_16974);
nand U17588 (N_17588,N_17035,N_16971);
nand U17589 (N_17589,N_16954,N_17211);
xor U17590 (N_17590,N_16827,N_17067);
xnor U17591 (N_17591,N_16967,N_16868);
xnor U17592 (N_17592,N_17382,N_17284);
or U17593 (N_17593,N_17164,N_17351);
xnor U17594 (N_17594,N_16862,N_17342);
and U17595 (N_17595,N_17183,N_16958);
and U17596 (N_17596,N_17146,N_17036);
nor U17597 (N_17597,N_16805,N_16879);
or U17598 (N_17598,N_17118,N_16988);
and U17599 (N_17599,N_17180,N_16894);
nor U17600 (N_17600,N_17330,N_17004);
or U17601 (N_17601,N_17014,N_16950);
or U17602 (N_17602,N_17245,N_17349);
and U17603 (N_17603,N_17328,N_17306);
nand U17604 (N_17604,N_16874,N_17128);
nor U17605 (N_17605,N_16893,N_17003);
and U17606 (N_17606,N_16832,N_17049);
nand U17607 (N_17607,N_17247,N_17262);
nand U17608 (N_17608,N_16972,N_16880);
nor U17609 (N_17609,N_16815,N_16927);
and U17610 (N_17610,N_17138,N_16801);
nand U17611 (N_17611,N_17141,N_16843);
nand U17612 (N_17612,N_17046,N_17240);
or U17613 (N_17613,N_17307,N_17375);
nand U17614 (N_17614,N_17299,N_17224);
or U17615 (N_17615,N_16929,N_17161);
nor U17616 (N_17616,N_17286,N_17112);
xor U17617 (N_17617,N_17239,N_16864);
xnor U17618 (N_17618,N_17291,N_17048);
nand U17619 (N_17619,N_17179,N_17268);
nand U17620 (N_17620,N_16995,N_17013);
nand U17621 (N_17621,N_17000,N_17104);
or U17622 (N_17622,N_16846,N_16860);
or U17623 (N_17623,N_17272,N_17304);
xnor U17624 (N_17624,N_17305,N_17364);
or U17625 (N_17625,N_16898,N_16989);
or U17626 (N_17626,N_16976,N_17350);
and U17627 (N_17627,N_17187,N_17319);
nor U17628 (N_17628,N_17301,N_17151);
nor U17629 (N_17629,N_17057,N_17229);
or U17630 (N_17630,N_17125,N_16892);
xor U17631 (N_17631,N_17241,N_16816);
and U17632 (N_17632,N_17345,N_17191);
or U17633 (N_17633,N_17287,N_16935);
or U17634 (N_17634,N_16856,N_17133);
nor U17635 (N_17635,N_17332,N_16807);
nand U17636 (N_17636,N_17082,N_17354);
nor U17637 (N_17637,N_17177,N_16934);
nor U17638 (N_17638,N_16904,N_17260);
nor U17639 (N_17639,N_16837,N_17147);
nand U17640 (N_17640,N_17380,N_16895);
or U17641 (N_17641,N_17315,N_16910);
nand U17642 (N_17642,N_16818,N_17365);
nand U17643 (N_17643,N_17100,N_16953);
or U17644 (N_17644,N_17361,N_17016);
and U17645 (N_17645,N_17083,N_16841);
or U17646 (N_17646,N_17362,N_17033);
nor U17647 (N_17647,N_17222,N_17011);
nor U17648 (N_17648,N_16946,N_17069);
nand U17649 (N_17649,N_17393,N_16992);
nor U17650 (N_17650,N_16847,N_17022);
nand U17651 (N_17651,N_16909,N_17356);
nor U17652 (N_17652,N_17359,N_17025);
and U17653 (N_17653,N_17130,N_17126);
nand U17654 (N_17654,N_16808,N_17276);
xnor U17655 (N_17655,N_17318,N_16979);
xnor U17656 (N_17656,N_17273,N_17279);
xnor U17657 (N_17657,N_16947,N_17231);
nor U17658 (N_17658,N_17197,N_16922);
nand U17659 (N_17659,N_17384,N_16956);
xor U17660 (N_17660,N_16858,N_16836);
nor U17661 (N_17661,N_17323,N_17092);
or U17662 (N_17662,N_17034,N_17259);
or U17663 (N_17663,N_16996,N_16997);
or U17664 (N_17664,N_17001,N_16886);
nand U17665 (N_17665,N_17074,N_17398);
nand U17666 (N_17666,N_17203,N_17278);
and U17667 (N_17667,N_17368,N_17213);
xor U17668 (N_17668,N_16917,N_17169);
nand U17669 (N_17669,N_17002,N_17357);
nand U17670 (N_17670,N_17173,N_17023);
nor U17671 (N_17671,N_17341,N_17322);
nor U17672 (N_17672,N_17236,N_16977);
nor U17673 (N_17673,N_17242,N_16820);
xnor U17674 (N_17674,N_16918,N_17238);
or U17675 (N_17675,N_17283,N_17369);
nor U17676 (N_17676,N_16938,N_17153);
and U17677 (N_17677,N_17010,N_17374);
or U17678 (N_17678,N_16869,N_17378);
and U17679 (N_17679,N_17303,N_17226);
xor U17680 (N_17680,N_16863,N_16952);
nand U17681 (N_17681,N_16964,N_17098);
nand U17682 (N_17682,N_17026,N_16999);
or U17683 (N_17683,N_16980,N_17193);
nand U17684 (N_17684,N_17223,N_16966);
nand U17685 (N_17685,N_16813,N_16948);
and U17686 (N_17686,N_17081,N_17121);
nor U17687 (N_17687,N_17219,N_17220);
and U17688 (N_17688,N_17198,N_17080);
and U17689 (N_17689,N_17054,N_17233);
xor U17690 (N_17690,N_16865,N_17202);
nand U17691 (N_17691,N_17139,N_17230);
xor U17692 (N_17692,N_17257,N_16921);
or U17693 (N_17693,N_17172,N_16978);
or U17694 (N_17694,N_17039,N_17015);
or U17695 (N_17695,N_17114,N_17195);
or U17696 (N_17696,N_16853,N_16901);
nor U17697 (N_17697,N_17079,N_16943);
and U17698 (N_17698,N_16959,N_17087);
xnor U17699 (N_17699,N_16949,N_17065);
xnor U17700 (N_17700,N_17236,N_17116);
and U17701 (N_17701,N_16831,N_16832);
or U17702 (N_17702,N_17382,N_16879);
or U17703 (N_17703,N_16984,N_16843);
nand U17704 (N_17704,N_17334,N_17213);
nor U17705 (N_17705,N_17317,N_17239);
xor U17706 (N_17706,N_16871,N_17385);
and U17707 (N_17707,N_17319,N_16957);
xnor U17708 (N_17708,N_17335,N_17089);
xnor U17709 (N_17709,N_17390,N_17127);
nand U17710 (N_17710,N_17232,N_17235);
and U17711 (N_17711,N_17395,N_17363);
nand U17712 (N_17712,N_17002,N_17144);
or U17713 (N_17713,N_17227,N_16918);
nor U17714 (N_17714,N_17175,N_17165);
and U17715 (N_17715,N_16822,N_17295);
nand U17716 (N_17716,N_17318,N_17005);
xnor U17717 (N_17717,N_17279,N_17315);
nand U17718 (N_17718,N_17300,N_17139);
nand U17719 (N_17719,N_17235,N_17046);
or U17720 (N_17720,N_17034,N_17126);
xnor U17721 (N_17721,N_16950,N_17312);
nand U17722 (N_17722,N_17393,N_17278);
or U17723 (N_17723,N_17214,N_17078);
nor U17724 (N_17724,N_16846,N_16875);
nand U17725 (N_17725,N_17346,N_17349);
or U17726 (N_17726,N_17249,N_17233);
and U17727 (N_17727,N_16805,N_17267);
nand U17728 (N_17728,N_16930,N_17278);
xnor U17729 (N_17729,N_16975,N_17194);
xnor U17730 (N_17730,N_17029,N_16993);
nand U17731 (N_17731,N_17264,N_16949);
nand U17732 (N_17732,N_17381,N_17366);
and U17733 (N_17733,N_16866,N_17205);
nor U17734 (N_17734,N_17006,N_17031);
nand U17735 (N_17735,N_16949,N_17302);
nor U17736 (N_17736,N_16850,N_17232);
nand U17737 (N_17737,N_16856,N_16980);
and U17738 (N_17738,N_17113,N_17088);
or U17739 (N_17739,N_16942,N_17062);
nor U17740 (N_17740,N_17069,N_17304);
nor U17741 (N_17741,N_16831,N_17251);
nor U17742 (N_17742,N_17218,N_17337);
nand U17743 (N_17743,N_16948,N_17252);
or U17744 (N_17744,N_17291,N_17155);
nor U17745 (N_17745,N_16884,N_16806);
xnor U17746 (N_17746,N_17357,N_17085);
nand U17747 (N_17747,N_16934,N_16904);
xnor U17748 (N_17748,N_17081,N_16864);
nor U17749 (N_17749,N_17086,N_17182);
nand U17750 (N_17750,N_17010,N_17082);
xnor U17751 (N_17751,N_16891,N_17258);
nand U17752 (N_17752,N_17009,N_17301);
and U17753 (N_17753,N_17018,N_16975);
nand U17754 (N_17754,N_17023,N_16932);
nand U17755 (N_17755,N_16949,N_16838);
xnor U17756 (N_17756,N_17058,N_16933);
and U17757 (N_17757,N_17171,N_17278);
nor U17758 (N_17758,N_17130,N_16936);
or U17759 (N_17759,N_17119,N_16883);
nand U17760 (N_17760,N_17090,N_16986);
or U17761 (N_17761,N_17077,N_17022);
and U17762 (N_17762,N_17003,N_17158);
xor U17763 (N_17763,N_16933,N_17063);
and U17764 (N_17764,N_16893,N_16841);
nand U17765 (N_17765,N_17395,N_17316);
nor U17766 (N_17766,N_17338,N_16978);
or U17767 (N_17767,N_17145,N_17228);
nor U17768 (N_17768,N_17216,N_16816);
and U17769 (N_17769,N_17187,N_16875);
or U17770 (N_17770,N_17232,N_17386);
nand U17771 (N_17771,N_17028,N_16924);
or U17772 (N_17772,N_17040,N_16812);
or U17773 (N_17773,N_17180,N_17215);
nand U17774 (N_17774,N_16849,N_17127);
or U17775 (N_17775,N_16951,N_16938);
and U17776 (N_17776,N_16974,N_17180);
nor U17777 (N_17777,N_17245,N_16899);
nand U17778 (N_17778,N_17015,N_17276);
nand U17779 (N_17779,N_17058,N_17141);
nand U17780 (N_17780,N_17381,N_17018);
nor U17781 (N_17781,N_16961,N_17137);
nand U17782 (N_17782,N_17101,N_17159);
xnor U17783 (N_17783,N_16828,N_17161);
nand U17784 (N_17784,N_17358,N_17388);
xnor U17785 (N_17785,N_17145,N_16977);
or U17786 (N_17786,N_16989,N_17107);
or U17787 (N_17787,N_17303,N_16989);
xor U17788 (N_17788,N_17043,N_17379);
nand U17789 (N_17789,N_16952,N_17113);
or U17790 (N_17790,N_16914,N_17394);
nor U17791 (N_17791,N_16998,N_17176);
xnor U17792 (N_17792,N_17171,N_16959);
and U17793 (N_17793,N_17152,N_17376);
nand U17794 (N_17794,N_17260,N_17373);
nand U17795 (N_17795,N_17372,N_17023);
xnor U17796 (N_17796,N_16849,N_17352);
nor U17797 (N_17797,N_17151,N_17239);
xnor U17798 (N_17798,N_17015,N_17392);
nor U17799 (N_17799,N_17240,N_16818);
or U17800 (N_17800,N_16930,N_17275);
or U17801 (N_17801,N_17372,N_16965);
and U17802 (N_17802,N_17064,N_17115);
nand U17803 (N_17803,N_17086,N_17366);
or U17804 (N_17804,N_17213,N_16964);
and U17805 (N_17805,N_17000,N_17394);
and U17806 (N_17806,N_16915,N_17192);
or U17807 (N_17807,N_17349,N_17373);
nand U17808 (N_17808,N_16954,N_16970);
xor U17809 (N_17809,N_16842,N_17374);
nor U17810 (N_17810,N_17091,N_16934);
and U17811 (N_17811,N_16925,N_16975);
and U17812 (N_17812,N_17008,N_16833);
nand U17813 (N_17813,N_17229,N_17052);
xor U17814 (N_17814,N_17112,N_17374);
nor U17815 (N_17815,N_16924,N_16986);
xnor U17816 (N_17816,N_16948,N_17064);
nor U17817 (N_17817,N_16883,N_16905);
and U17818 (N_17818,N_16982,N_17127);
nor U17819 (N_17819,N_17079,N_16887);
xnor U17820 (N_17820,N_17001,N_16933);
and U17821 (N_17821,N_16819,N_17354);
or U17822 (N_17822,N_17072,N_17046);
xnor U17823 (N_17823,N_17211,N_16850);
nand U17824 (N_17824,N_17232,N_17335);
nor U17825 (N_17825,N_16850,N_16980);
xnor U17826 (N_17826,N_17088,N_17174);
and U17827 (N_17827,N_16921,N_16876);
nor U17828 (N_17828,N_17019,N_17288);
and U17829 (N_17829,N_17074,N_17104);
nand U17830 (N_17830,N_16803,N_17094);
nor U17831 (N_17831,N_17383,N_16987);
nand U17832 (N_17832,N_16908,N_17021);
or U17833 (N_17833,N_16848,N_17051);
and U17834 (N_17834,N_17276,N_17195);
nor U17835 (N_17835,N_17173,N_16929);
and U17836 (N_17836,N_17031,N_17292);
or U17837 (N_17837,N_16805,N_17269);
and U17838 (N_17838,N_17072,N_17154);
xnor U17839 (N_17839,N_17258,N_17323);
or U17840 (N_17840,N_16867,N_17308);
or U17841 (N_17841,N_17099,N_16972);
nand U17842 (N_17842,N_16900,N_17266);
nor U17843 (N_17843,N_17345,N_17326);
nand U17844 (N_17844,N_17275,N_17192);
nand U17845 (N_17845,N_17107,N_16846);
nand U17846 (N_17846,N_16976,N_17148);
nand U17847 (N_17847,N_17245,N_17150);
nor U17848 (N_17848,N_16904,N_16855);
xnor U17849 (N_17849,N_17211,N_16923);
nor U17850 (N_17850,N_16889,N_17069);
and U17851 (N_17851,N_17031,N_17394);
nor U17852 (N_17852,N_16885,N_17176);
nand U17853 (N_17853,N_17018,N_17025);
nor U17854 (N_17854,N_17276,N_16995);
xor U17855 (N_17855,N_16892,N_17262);
or U17856 (N_17856,N_17347,N_17399);
or U17857 (N_17857,N_17070,N_16901);
and U17858 (N_17858,N_16819,N_17152);
xor U17859 (N_17859,N_17006,N_17185);
xnor U17860 (N_17860,N_17169,N_16967);
or U17861 (N_17861,N_17328,N_16895);
and U17862 (N_17862,N_17356,N_16994);
and U17863 (N_17863,N_16881,N_17169);
nand U17864 (N_17864,N_17349,N_16817);
and U17865 (N_17865,N_16929,N_16910);
and U17866 (N_17866,N_16918,N_17276);
xnor U17867 (N_17867,N_16836,N_17248);
xor U17868 (N_17868,N_17056,N_16800);
nor U17869 (N_17869,N_17299,N_16882);
or U17870 (N_17870,N_16991,N_16888);
and U17871 (N_17871,N_16818,N_17008);
nor U17872 (N_17872,N_17064,N_17310);
or U17873 (N_17873,N_17238,N_17373);
and U17874 (N_17874,N_17218,N_17026);
nor U17875 (N_17875,N_16912,N_17145);
or U17876 (N_17876,N_16819,N_17069);
nor U17877 (N_17877,N_16931,N_16979);
nand U17878 (N_17878,N_17008,N_17180);
xnor U17879 (N_17879,N_16919,N_16867);
or U17880 (N_17880,N_17066,N_16862);
nor U17881 (N_17881,N_17375,N_17155);
nor U17882 (N_17882,N_16853,N_16816);
nand U17883 (N_17883,N_17179,N_16816);
and U17884 (N_17884,N_17291,N_17006);
nand U17885 (N_17885,N_16907,N_17156);
xnor U17886 (N_17886,N_16912,N_17275);
xnor U17887 (N_17887,N_17126,N_17162);
and U17888 (N_17888,N_16858,N_17176);
or U17889 (N_17889,N_17220,N_17218);
nor U17890 (N_17890,N_17031,N_17169);
and U17891 (N_17891,N_16963,N_16950);
nand U17892 (N_17892,N_17285,N_16975);
xor U17893 (N_17893,N_16826,N_17124);
nor U17894 (N_17894,N_17139,N_17249);
xor U17895 (N_17895,N_17241,N_16916);
nand U17896 (N_17896,N_16897,N_17102);
nor U17897 (N_17897,N_16813,N_16890);
and U17898 (N_17898,N_17002,N_16870);
xnor U17899 (N_17899,N_16885,N_17196);
nand U17900 (N_17900,N_17221,N_16834);
xor U17901 (N_17901,N_17396,N_17056);
xnor U17902 (N_17902,N_17012,N_16874);
xor U17903 (N_17903,N_17149,N_16919);
nand U17904 (N_17904,N_17199,N_16819);
xor U17905 (N_17905,N_17074,N_17189);
nor U17906 (N_17906,N_17119,N_17092);
nor U17907 (N_17907,N_16834,N_17024);
xnor U17908 (N_17908,N_17327,N_17341);
or U17909 (N_17909,N_17062,N_17001);
nor U17910 (N_17910,N_16919,N_17085);
nor U17911 (N_17911,N_16991,N_16984);
and U17912 (N_17912,N_17392,N_17185);
and U17913 (N_17913,N_17178,N_17320);
nand U17914 (N_17914,N_17207,N_16998);
and U17915 (N_17915,N_17263,N_17340);
or U17916 (N_17916,N_16992,N_17236);
or U17917 (N_17917,N_17087,N_16844);
nand U17918 (N_17918,N_17079,N_16961);
and U17919 (N_17919,N_17041,N_16855);
or U17920 (N_17920,N_16834,N_17288);
nor U17921 (N_17921,N_16868,N_17353);
xor U17922 (N_17922,N_17147,N_17263);
nor U17923 (N_17923,N_17144,N_16801);
and U17924 (N_17924,N_17324,N_16913);
nand U17925 (N_17925,N_17098,N_16872);
xor U17926 (N_17926,N_17188,N_17386);
and U17927 (N_17927,N_17164,N_17107);
and U17928 (N_17928,N_16900,N_17396);
xnor U17929 (N_17929,N_16848,N_16910);
or U17930 (N_17930,N_17281,N_16915);
nand U17931 (N_17931,N_17273,N_17342);
xor U17932 (N_17932,N_17120,N_17347);
or U17933 (N_17933,N_17004,N_17242);
nor U17934 (N_17934,N_16983,N_17288);
xnor U17935 (N_17935,N_17035,N_17362);
xor U17936 (N_17936,N_17364,N_17288);
nand U17937 (N_17937,N_17120,N_17047);
nand U17938 (N_17938,N_16812,N_17331);
xnor U17939 (N_17939,N_17194,N_17283);
and U17940 (N_17940,N_17166,N_16880);
xnor U17941 (N_17941,N_17231,N_17079);
nor U17942 (N_17942,N_17352,N_16978);
and U17943 (N_17943,N_17172,N_17036);
or U17944 (N_17944,N_17395,N_17319);
and U17945 (N_17945,N_17036,N_17035);
nor U17946 (N_17946,N_17238,N_17343);
nand U17947 (N_17947,N_16851,N_17154);
nand U17948 (N_17948,N_16906,N_17040);
and U17949 (N_17949,N_17239,N_17302);
and U17950 (N_17950,N_17293,N_17302);
xor U17951 (N_17951,N_17070,N_17013);
and U17952 (N_17952,N_17214,N_16985);
xnor U17953 (N_17953,N_16880,N_17204);
nand U17954 (N_17954,N_17141,N_17134);
and U17955 (N_17955,N_17388,N_17071);
xnor U17956 (N_17956,N_16802,N_17141);
and U17957 (N_17957,N_17367,N_17390);
and U17958 (N_17958,N_16830,N_17179);
xor U17959 (N_17959,N_17142,N_17292);
and U17960 (N_17960,N_16892,N_17301);
or U17961 (N_17961,N_17211,N_16883);
xnor U17962 (N_17962,N_17381,N_17289);
or U17963 (N_17963,N_16866,N_16812);
nand U17964 (N_17964,N_17348,N_17077);
or U17965 (N_17965,N_17130,N_17015);
and U17966 (N_17966,N_17139,N_16996);
nand U17967 (N_17967,N_16889,N_16924);
nor U17968 (N_17968,N_17369,N_16801);
nand U17969 (N_17969,N_16978,N_17144);
nor U17970 (N_17970,N_16956,N_17211);
and U17971 (N_17971,N_17039,N_17346);
nor U17972 (N_17972,N_17040,N_17024);
nor U17973 (N_17973,N_17274,N_16950);
nor U17974 (N_17974,N_17074,N_17020);
and U17975 (N_17975,N_17004,N_17290);
nand U17976 (N_17976,N_17202,N_16955);
nand U17977 (N_17977,N_17074,N_17363);
nor U17978 (N_17978,N_17212,N_17220);
or U17979 (N_17979,N_17069,N_17265);
nor U17980 (N_17980,N_17163,N_17074);
nor U17981 (N_17981,N_16865,N_16943);
xor U17982 (N_17982,N_16842,N_16918);
nor U17983 (N_17983,N_16921,N_17249);
nor U17984 (N_17984,N_17349,N_16920);
and U17985 (N_17985,N_16856,N_16992);
nor U17986 (N_17986,N_17102,N_16829);
xnor U17987 (N_17987,N_17026,N_16979);
and U17988 (N_17988,N_16974,N_16920);
and U17989 (N_17989,N_17320,N_17283);
or U17990 (N_17990,N_17198,N_17057);
nand U17991 (N_17991,N_17014,N_17284);
or U17992 (N_17992,N_17138,N_16925);
nor U17993 (N_17993,N_17255,N_16821);
xnor U17994 (N_17994,N_17116,N_16852);
nor U17995 (N_17995,N_17277,N_17320);
and U17996 (N_17996,N_17188,N_17358);
nand U17997 (N_17997,N_17163,N_17271);
or U17998 (N_17998,N_16925,N_17009);
nor U17999 (N_17999,N_17180,N_17384);
nor U18000 (N_18000,N_17582,N_17444);
nor U18001 (N_18001,N_17401,N_17613);
nor U18002 (N_18002,N_17979,N_17866);
or U18003 (N_18003,N_17445,N_17563);
or U18004 (N_18004,N_17455,N_17650);
or U18005 (N_18005,N_17480,N_17681);
or U18006 (N_18006,N_17605,N_17589);
and U18007 (N_18007,N_17701,N_17406);
nand U18008 (N_18008,N_17891,N_17544);
nor U18009 (N_18009,N_17792,N_17910);
nand U18010 (N_18010,N_17721,N_17590);
xnor U18011 (N_18011,N_17657,N_17500);
and U18012 (N_18012,N_17606,N_17976);
nor U18013 (N_18013,N_17646,N_17689);
nor U18014 (N_18014,N_17411,N_17895);
nand U18015 (N_18015,N_17964,N_17461);
and U18016 (N_18016,N_17817,N_17495);
nor U18017 (N_18017,N_17628,N_17512);
nor U18018 (N_18018,N_17803,N_17953);
nor U18019 (N_18019,N_17728,N_17928);
xor U18020 (N_18020,N_17741,N_17614);
xor U18021 (N_18021,N_17631,N_17536);
or U18022 (N_18022,N_17975,N_17905);
or U18023 (N_18023,N_17715,N_17846);
nand U18024 (N_18024,N_17777,N_17610);
nor U18025 (N_18025,N_17601,N_17796);
nand U18026 (N_18026,N_17597,N_17934);
or U18027 (N_18027,N_17694,N_17938);
nand U18028 (N_18028,N_17894,N_17767);
xor U18029 (N_18029,N_17424,N_17824);
and U18030 (N_18030,N_17965,N_17983);
nor U18031 (N_18031,N_17408,N_17751);
nor U18032 (N_18032,N_17914,N_17477);
or U18033 (N_18033,N_17652,N_17471);
xor U18034 (N_18034,N_17580,N_17572);
xnor U18035 (N_18035,N_17729,N_17991);
or U18036 (N_18036,N_17760,N_17437);
or U18037 (N_18037,N_17873,N_17821);
nand U18038 (N_18038,N_17837,N_17643);
or U18039 (N_18039,N_17476,N_17510);
and U18040 (N_18040,N_17430,N_17562);
or U18041 (N_18041,N_17850,N_17519);
xor U18042 (N_18042,N_17774,N_17770);
or U18043 (N_18043,N_17505,N_17603);
nor U18044 (N_18044,N_17484,N_17506);
or U18045 (N_18045,N_17448,N_17849);
nor U18046 (N_18046,N_17787,N_17638);
nor U18047 (N_18047,N_17750,N_17680);
nand U18048 (N_18048,N_17452,N_17920);
nor U18049 (N_18049,N_17665,N_17911);
xor U18050 (N_18050,N_17804,N_17919);
or U18051 (N_18051,N_17888,N_17443);
and U18052 (N_18052,N_17441,N_17418);
nor U18053 (N_18053,N_17555,N_17768);
or U18054 (N_18054,N_17784,N_17875);
nand U18055 (N_18055,N_17440,N_17602);
nor U18056 (N_18056,N_17838,N_17662);
and U18057 (N_18057,N_17859,N_17799);
nor U18058 (N_18058,N_17529,N_17465);
or U18059 (N_18059,N_17672,N_17966);
or U18060 (N_18060,N_17608,N_17731);
nor U18061 (N_18061,N_17781,N_17982);
nand U18062 (N_18062,N_17592,N_17463);
and U18063 (N_18063,N_17835,N_17503);
nor U18064 (N_18064,N_17901,N_17973);
xnor U18065 (N_18065,N_17707,N_17704);
xnor U18066 (N_18066,N_17676,N_17648);
and U18067 (N_18067,N_17742,N_17712);
and U18068 (N_18068,N_17773,N_17611);
xor U18069 (N_18069,N_17706,N_17940);
and U18070 (N_18070,N_17852,N_17933);
and U18071 (N_18071,N_17696,N_17421);
nor U18072 (N_18072,N_17764,N_17997);
or U18073 (N_18073,N_17730,N_17615);
nand U18074 (N_18074,N_17474,N_17422);
or U18075 (N_18075,N_17412,N_17833);
nand U18076 (N_18076,N_17913,N_17753);
and U18077 (N_18077,N_17591,N_17878);
xor U18078 (N_18078,N_17483,N_17625);
or U18079 (N_18079,N_17703,N_17797);
nand U18080 (N_18080,N_17860,N_17549);
xnor U18081 (N_18081,N_17488,N_17486);
nand U18082 (N_18082,N_17619,N_17624);
and U18083 (N_18083,N_17433,N_17658);
nand U18084 (N_18084,N_17863,N_17726);
nand U18085 (N_18085,N_17647,N_17818);
or U18086 (N_18086,N_17559,N_17840);
xnor U18087 (N_18087,N_17565,N_17598);
nor U18088 (N_18088,N_17702,N_17989);
nand U18089 (N_18089,N_17524,N_17851);
nand U18090 (N_18090,N_17434,N_17865);
nor U18091 (N_18091,N_17766,N_17889);
nor U18092 (N_18092,N_17716,N_17780);
nor U18093 (N_18093,N_17747,N_17718);
xnor U18094 (N_18094,N_17684,N_17816);
and U18095 (N_18095,N_17834,N_17502);
xnor U18096 (N_18096,N_17537,N_17775);
nor U18097 (N_18097,N_17692,N_17479);
and U18098 (N_18098,N_17705,N_17746);
nand U18099 (N_18099,N_17884,N_17595);
nor U18100 (N_18100,N_17732,N_17688);
xnor U18101 (N_18101,N_17987,N_17902);
nand U18102 (N_18102,N_17986,N_17513);
nand U18103 (N_18103,N_17890,N_17578);
or U18104 (N_18104,N_17808,N_17990);
nor U18105 (N_18105,N_17467,N_17785);
nor U18106 (N_18106,N_17558,N_17687);
and U18107 (N_18107,N_17829,N_17581);
nor U18108 (N_18108,N_17737,N_17954);
nand U18109 (N_18109,N_17814,N_17641);
nand U18110 (N_18110,N_17548,N_17872);
nor U18111 (N_18111,N_17475,N_17653);
xor U18112 (N_18112,N_17621,N_17815);
nor U18113 (N_18113,N_17809,N_17725);
or U18114 (N_18114,N_17822,N_17534);
or U18115 (N_18115,N_17869,N_17607);
and U18116 (N_18116,N_17828,N_17700);
and U18117 (N_18117,N_17404,N_17617);
nand U18118 (N_18118,N_17930,N_17917);
or U18119 (N_18119,N_17636,N_17627);
xnor U18120 (N_18120,N_17675,N_17862);
or U18121 (N_18121,N_17584,N_17664);
or U18122 (N_18122,N_17487,N_17970);
and U18123 (N_18123,N_17683,N_17922);
and U18124 (N_18124,N_17633,N_17736);
or U18125 (N_18125,N_17561,N_17845);
xnor U18126 (N_18126,N_17795,N_17629);
nand U18127 (N_18127,N_17868,N_17654);
and U18128 (N_18128,N_17575,N_17670);
and U18129 (N_18129,N_17454,N_17724);
xor U18130 (N_18130,N_17793,N_17660);
xor U18131 (N_18131,N_17844,N_17535);
and U18132 (N_18132,N_17936,N_17813);
and U18133 (N_18133,N_17539,N_17402);
nand U18134 (N_18134,N_17727,N_17880);
or U18135 (N_18135,N_17493,N_17415);
or U18136 (N_18136,N_17466,N_17831);
nand U18137 (N_18137,N_17820,N_17546);
and U18138 (N_18138,N_17843,N_17508);
nand U18139 (N_18139,N_17618,N_17887);
nor U18140 (N_18140,N_17413,N_17588);
nor U18141 (N_18141,N_17935,N_17527);
nand U18142 (N_18142,N_17511,N_17407);
xnor U18143 (N_18143,N_17516,N_17651);
nand U18144 (N_18144,N_17722,N_17576);
xor U18145 (N_18145,N_17848,N_17962);
xor U18146 (N_18146,N_17553,N_17945);
or U18147 (N_18147,N_17984,N_17832);
nor U18148 (N_18148,N_17789,N_17950);
nand U18149 (N_18149,N_17557,N_17570);
nor U18150 (N_18150,N_17957,N_17420);
nor U18151 (N_18151,N_17881,N_17893);
nand U18152 (N_18152,N_17645,N_17594);
and U18153 (N_18153,N_17963,N_17802);
and U18154 (N_18154,N_17711,N_17874);
xor U18155 (N_18155,N_17447,N_17717);
nor U18156 (N_18156,N_17697,N_17709);
and U18157 (N_18157,N_17959,N_17659);
and U18158 (N_18158,N_17757,N_17755);
xnor U18159 (N_18159,N_17504,N_17490);
nor U18160 (N_18160,N_17497,N_17426);
xor U18161 (N_18161,N_17518,N_17918);
nand U18162 (N_18162,N_17871,N_17879);
xnor U18163 (N_18163,N_17446,N_17853);
or U18164 (N_18164,N_17533,N_17442);
nor U18165 (N_18165,N_17765,N_17509);
and U18166 (N_18166,N_17735,N_17972);
nor U18167 (N_18167,N_17669,N_17656);
nor U18168 (N_18168,N_17417,N_17839);
xnor U18169 (N_18169,N_17435,N_17942);
xnor U18170 (N_18170,N_17679,N_17977);
and U18171 (N_18171,N_17685,N_17531);
nand U18172 (N_18172,N_17739,N_17995);
nand U18173 (N_18173,N_17886,N_17836);
nor U18174 (N_18174,N_17550,N_17958);
or U18175 (N_18175,N_17826,N_17642);
nand U18176 (N_18176,N_17449,N_17806);
and U18177 (N_18177,N_17961,N_17939);
or U18178 (N_18178,N_17457,N_17779);
xor U18179 (N_18179,N_17423,N_17955);
nor U18180 (N_18180,N_17492,N_17460);
nand U18181 (N_18181,N_17690,N_17823);
xnor U18182 (N_18182,N_17778,N_17714);
or U18183 (N_18183,N_17514,N_17996);
nand U18184 (N_18184,N_17593,N_17432);
or U18185 (N_18185,N_17405,N_17926);
or U18186 (N_18186,N_17967,N_17456);
xor U18187 (N_18187,N_17956,N_17897);
xnor U18188 (N_18188,N_17678,N_17551);
and U18189 (N_18189,N_17708,N_17587);
and U18190 (N_18190,N_17462,N_17499);
or U18191 (N_18191,N_17798,N_17772);
nor U18192 (N_18192,N_17812,N_17943);
or U18193 (N_18193,N_17567,N_17927);
xor U18194 (N_18194,N_17969,N_17612);
or U18195 (N_18195,N_17428,N_17691);
or U18196 (N_18196,N_17521,N_17855);
and U18197 (N_18197,N_17949,N_17783);
or U18198 (N_18198,N_17482,N_17762);
and U18199 (N_18199,N_17929,N_17841);
nand U18200 (N_18200,N_17907,N_17695);
or U18201 (N_18201,N_17574,N_17450);
and U18202 (N_18202,N_17556,N_17632);
xor U18203 (N_18203,N_17596,N_17526);
or U18204 (N_18204,N_17925,N_17425);
nor U18205 (N_18205,N_17857,N_17947);
and U18206 (N_18206,N_17517,N_17501);
nand U18207 (N_18207,N_17698,N_17637);
xnor U18208 (N_18208,N_17666,N_17566);
or U18209 (N_18209,N_17552,N_17674);
or U18210 (N_18210,N_17403,N_17661);
xnor U18211 (N_18211,N_17523,N_17748);
nor U18212 (N_18212,N_17682,N_17667);
and U18213 (N_18213,N_17481,N_17885);
or U18214 (N_18214,N_17807,N_17616);
and U18215 (N_18215,N_17410,N_17906);
nand U18216 (N_18216,N_17994,N_17931);
nor U18217 (N_18217,N_17790,N_17464);
nor U18218 (N_18218,N_17507,N_17620);
xnor U18219 (N_18219,N_17960,N_17622);
xnor U18220 (N_18220,N_17937,N_17568);
or U18221 (N_18221,N_17469,N_17644);
nand U18222 (N_18222,N_17649,N_17740);
xnor U18223 (N_18223,N_17743,N_17585);
and U18224 (N_18224,N_17541,N_17543);
nand U18225 (N_18225,N_17791,N_17909);
or U18226 (N_18226,N_17400,N_17655);
and U18227 (N_18227,N_17470,N_17974);
nand U18228 (N_18228,N_17761,N_17861);
nor U18229 (N_18229,N_17981,N_17416);
nand U18230 (N_18230,N_17763,N_17998);
nor U18231 (N_18231,N_17842,N_17946);
or U18232 (N_18232,N_17528,N_17604);
nand U18233 (N_18233,N_17899,N_17577);
and U18234 (N_18234,N_17564,N_17573);
nor U18235 (N_18235,N_17525,N_17453);
nand U18236 (N_18236,N_17819,N_17924);
nand U18237 (N_18237,N_17600,N_17847);
xor U18238 (N_18238,N_17794,N_17800);
or U18239 (N_18239,N_17498,N_17985);
nor U18240 (N_18240,N_17999,N_17473);
nand U18241 (N_18241,N_17673,N_17903);
nand U18242 (N_18242,N_17892,N_17870);
or U18243 (N_18243,N_17569,N_17414);
or U18244 (N_18244,N_17538,N_17825);
and U18245 (N_18245,N_17734,N_17677);
and U18246 (N_18246,N_17560,N_17439);
or U18247 (N_18247,N_17867,N_17671);
xnor U18248 (N_18248,N_17908,N_17427);
nor U18249 (N_18249,N_17951,N_17978);
and U18250 (N_18250,N_17542,N_17745);
nand U18251 (N_18251,N_17915,N_17776);
and U18252 (N_18252,N_17749,N_17921);
nand U18253 (N_18253,N_17723,N_17810);
nor U18254 (N_18254,N_17713,N_17882);
nor U18255 (N_18255,N_17520,N_17858);
nor U18256 (N_18256,N_17699,N_17491);
or U18257 (N_18257,N_17744,N_17932);
nor U18258 (N_18258,N_17686,N_17409);
and U18259 (N_18259,N_17663,N_17496);
and U18260 (N_18260,N_17759,N_17668);
nor U18261 (N_18261,N_17472,N_17583);
and U18262 (N_18262,N_17898,N_17877);
and U18263 (N_18263,N_17554,N_17710);
xnor U18264 (N_18264,N_17640,N_17522);
nor U18265 (N_18265,N_17733,N_17752);
or U18266 (N_18266,N_17579,N_17923);
and U18267 (N_18267,N_17436,N_17494);
and U18268 (N_18268,N_17782,N_17693);
or U18269 (N_18269,N_17988,N_17896);
xnor U18270 (N_18270,N_17419,N_17438);
or U18271 (N_18271,N_17771,N_17827);
nand U18272 (N_18272,N_17431,N_17941);
nand U18273 (N_18273,N_17738,N_17515);
nor U18274 (N_18274,N_17720,N_17635);
and U18275 (N_18275,N_17599,N_17489);
and U18276 (N_18276,N_17468,N_17532);
nor U18277 (N_18277,N_17626,N_17864);
or U18278 (N_18278,N_17609,N_17992);
nor U18279 (N_18279,N_17971,N_17948);
or U18280 (N_18280,N_17540,N_17788);
and U18281 (N_18281,N_17805,N_17952);
xor U18282 (N_18282,N_17916,N_17944);
and U18283 (N_18283,N_17571,N_17900);
and U18284 (N_18284,N_17856,N_17811);
nand U18285 (N_18285,N_17912,N_17545);
nand U18286 (N_18286,N_17623,N_17876);
nor U18287 (N_18287,N_17547,N_17485);
xnor U18288 (N_18288,N_17769,N_17980);
nor U18289 (N_18289,N_17630,N_17586);
xnor U18290 (N_18290,N_17854,N_17639);
xnor U18291 (N_18291,N_17883,N_17478);
and U18292 (N_18292,N_17459,N_17758);
nor U18293 (N_18293,N_17993,N_17968);
and U18294 (N_18294,N_17801,N_17634);
nand U18295 (N_18295,N_17458,N_17451);
and U18296 (N_18296,N_17719,N_17904);
xnor U18297 (N_18297,N_17429,N_17530);
nand U18298 (N_18298,N_17786,N_17830);
nand U18299 (N_18299,N_17754,N_17756);
xnor U18300 (N_18300,N_17846,N_17425);
or U18301 (N_18301,N_17527,N_17622);
nand U18302 (N_18302,N_17621,N_17689);
nor U18303 (N_18303,N_17429,N_17970);
nor U18304 (N_18304,N_17751,N_17573);
nor U18305 (N_18305,N_17877,N_17661);
or U18306 (N_18306,N_17703,N_17518);
nand U18307 (N_18307,N_17702,N_17607);
xnor U18308 (N_18308,N_17862,N_17569);
and U18309 (N_18309,N_17787,N_17818);
or U18310 (N_18310,N_17524,N_17835);
xor U18311 (N_18311,N_17724,N_17765);
nor U18312 (N_18312,N_17925,N_17885);
or U18313 (N_18313,N_17587,N_17894);
and U18314 (N_18314,N_17751,N_17419);
or U18315 (N_18315,N_17685,N_17976);
or U18316 (N_18316,N_17680,N_17405);
xor U18317 (N_18317,N_17832,N_17668);
or U18318 (N_18318,N_17922,N_17523);
xor U18319 (N_18319,N_17842,N_17980);
and U18320 (N_18320,N_17765,N_17828);
nand U18321 (N_18321,N_17754,N_17807);
nor U18322 (N_18322,N_17605,N_17865);
nor U18323 (N_18323,N_17572,N_17521);
and U18324 (N_18324,N_17678,N_17812);
nor U18325 (N_18325,N_17919,N_17829);
and U18326 (N_18326,N_17788,N_17777);
and U18327 (N_18327,N_17729,N_17795);
nand U18328 (N_18328,N_17521,N_17682);
nand U18329 (N_18329,N_17610,N_17509);
xor U18330 (N_18330,N_17933,N_17450);
xor U18331 (N_18331,N_17995,N_17713);
xnor U18332 (N_18332,N_17690,N_17912);
xnor U18333 (N_18333,N_17561,N_17519);
nor U18334 (N_18334,N_17920,N_17709);
or U18335 (N_18335,N_17804,N_17558);
or U18336 (N_18336,N_17508,N_17437);
nand U18337 (N_18337,N_17935,N_17916);
and U18338 (N_18338,N_17541,N_17930);
or U18339 (N_18339,N_17631,N_17456);
nor U18340 (N_18340,N_17500,N_17619);
and U18341 (N_18341,N_17506,N_17893);
nand U18342 (N_18342,N_17478,N_17712);
nand U18343 (N_18343,N_17595,N_17857);
nand U18344 (N_18344,N_17782,N_17871);
xnor U18345 (N_18345,N_17493,N_17955);
or U18346 (N_18346,N_17565,N_17689);
nand U18347 (N_18347,N_17960,N_17422);
nor U18348 (N_18348,N_17748,N_17404);
nor U18349 (N_18349,N_17945,N_17784);
nand U18350 (N_18350,N_17973,N_17643);
xnor U18351 (N_18351,N_17864,N_17557);
nand U18352 (N_18352,N_17762,N_17985);
nor U18353 (N_18353,N_17462,N_17703);
and U18354 (N_18354,N_17709,N_17934);
nand U18355 (N_18355,N_17539,N_17695);
or U18356 (N_18356,N_17560,N_17886);
or U18357 (N_18357,N_17931,N_17712);
xor U18358 (N_18358,N_17423,N_17687);
xor U18359 (N_18359,N_17942,N_17623);
nor U18360 (N_18360,N_17904,N_17899);
and U18361 (N_18361,N_17834,N_17641);
xor U18362 (N_18362,N_17493,N_17805);
nor U18363 (N_18363,N_17808,N_17953);
or U18364 (N_18364,N_17420,N_17728);
nor U18365 (N_18365,N_17421,N_17541);
and U18366 (N_18366,N_17693,N_17454);
nor U18367 (N_18367,N_17649,N_17596);
nor U18368 (N_18368,N_17938,N_17706);
nand U18369 (N_18369,N_17953,N_17610);
xor U18370 (N_18370,N_17871,N_17513);
and U18371 (N_18371,N_17574,N_17939);
nor U18372 (N_18372,N_17744,N_17458);
nand U18373 (N_18373,N_17478,N_17852);
xnor U18374 (N_18374,N_17813,N_17905);
xor U18375 (N_18375,N_17748,N_17847);
nor U18376 (N_18376,N_17862,N_17984);
nand U18377 (N_18377,N_17624,N_17972);
nor U18378 (N_18378,N_17504,N_17803);
nand U18379 (N_18379,N_17866,N_17604);
xor U18380 (N_18380,N_17641,N_17403);
or U18381 (N_18381,N_17955,N_17400);
nor U18382 (N_18382,N_17756,N_17701);
and U18383 (N_18383,N_17656,N_17466);
nor U18384 (N_18384,N_17491,N_17589);
nand U18385 (N_18385,N_17789,N_17446);
or U18386 (N_18386,N_17489,N_17527);
and U18387 (N_18387,N_17428,N_17920);
and U18388 (N_18388,N_17916,N_17608);
and U18389 (N_18389,N_17514,N_17724);
nor U18390 (N_18390,N_17678,N_17513);
nor U18391 (N_18391,N_17939,N_17833);
and U18392 (N_18392,N_17702,N_17871);
nand U18393 (N_18393,N_17780,N_17845);
nor U18394 (N_18394,N_17424,N_17870);
nor U18395 (N_18395,N_17484,N_17693);
and U18396 (N_18396,N_17810,N_17738);
or U18397 (N_18397,N_17568,N_17482);
and U18398 (N_18398,N_17452,N_17404);
nand U18399 (N_18399,N_17866,N_17567);
xor U18400 (N_18400,N_17620,N_17822);
xor U18401 (N_18401,N_17978,N_17448);
or U18402 (N_18402,N_17858,N_17560);
xor U18403 (N_18403,N_17892,N_17898);
nor U18404 (N_18404,N_17761,N_17693);
nor U18405 (N_18405,N_17467,N_17787);
xnor U18406 (N_18406,N_17423,N_17548);
xor U18407 (N_18407,N_17439,N_17406);
nand U18408 (N_18408,N_17534,N_17607);
or U18409 (N_18409,N_17753,N_17825);
nor U18410 (N_18410,N_17511,N_17725);
nor U18411 (N_18411,N_17436,N_17943);
nor U18412 (N_18412,N_17496,N_17920);
xor U18413 (N_18413,N_17474,N_17917);
xnor U18414 (N_18414,N_17716,N_17991);
and U18415 (N_18415,N_17621,N_17532);
nor U18416 (N_18416,N_17434,N_17626);
xor U18417 (N_18417,N_17855,N_17617);
nand U18418 (N_18418,N_17960,N_17811);
and U18419 (N_18419,N_17943,N_17734);
xnor U18420 (N_18420,N_17812,N_17632);
nand U18421 (N_18421,N_17604,N_17862);
nor U18422 (N_18422,N_17529,N_17913);
nor U18423 (N_18423,N_17673,N_17824);
nand U18424 (N_18424,N_17876,N_17633);
xor U18425 (N_18425,N_17538,N_17915);
and U18426 (N_18426,N_17653,N_17638);
nor U18427 (N_18427,N_17683,N_17814);
xnor U18428 (N_18428,N_17640,N_17998);
nor U18429 (N_18429,N_17540,N_17908);
xnor U18430 (N_18430,N_17670,N_17726);
xor U18431 (N_18431,N_17834,N_17488);
and U18432 (N_18432,N_17761,N_17835);
nand U18433 (N_18433,N_17615,N_17593);
nor U18434 (N_18434,N_17950,N_17808);
and U18435 (N_18435,N_17803,N_17874);
and U18436 (N_18436,N_17743,N_17944);
xnor U18437 (N_18437,N_17856,N_17572);
and U18438 (N_18438,N_17550,N_17982);
nor U18439 (N_18439,N_17402,N_17711);
or U18440 (N_18440,N_17951,N_17405);
xor U18441 (N_18441,N_17590,N_17748);
or U18442 (N_18442,N_17865,N_17670);
nand U18443 (N_18443,N_17440,N_17541);
nor U18444 (N_18444,N_17414,N_17872);
or U18445 (N_18445,N_17659,N_17902);
and U18446 (N_18446,N_17804,N_17923);
and U18447 (N_18447,N_17756,N_17707);
and U18448 (N_18448,N_17464,N_17911);
nor U18449 (N_18449,N_17502,N_17712);
xor U18450 (N_18450,N_17562,N_17668);
and U18451 (N_18451,N_17408,N_17734);
nor U18452 (N_18452,N_17440,N_17598);
nor U18453 (N_18453,N_17755,N_17479);
nor U18454 (N_18454,N_17713,N_17754);
or U18455 (N_18455,N_17577,N_17824);
nand U18456 (N_18456,N_17790,N_17443);
or U18457 (N_18457,N_17441,N_17943);
and U18458 (N_18458,N_17812,N_17860);
xor U18459 (N_18459,N_17419,N_17989);
and U18460 (N_18460,N_17539,N_17407);
nor U18461 (N_18461,N_17954,N_17557);
and U18462 (N_18462,N_17874,N_17652);
nand U18463 (N_18463,N_17540,N_17671);
xor U18464 (N_18464,N_17711,N_17808);
or U18465 (N_18465,N_17819,N_17526);
nand U18466 (N_18466,N_17906,N_17723);
xor U18467 (N_18467,N_17820,N_17748);
nor U18468 (N_18468,N_17631,N_17857);
nor U18469 (N_18469,N_17820,N_17735);
xor U18470 (N_18470,N_17579,N_17892);
nand U18471 (N_18471,N_17896,N_17515);
nor U18472 (N_18472,N_17725,N_17739);
or U18473 (N_18473,N_17556,N_17642);
or U18474 (N_18474,N_17893,N_17447);
xnor U18475 (N_18475,N_17967,N_17502);
nand U18476 (N_18476,N_17567,N_17718);
nand U18477 (N_18477,N_17656,N_17560);
nor U18478 (N_18478,N_17808,N_17666);
xnor U18479 (N_18479,N_17940,N_17604);
and U18480 (N_18480,N_17725,N_17720);
or U18481 (N_18481,N_17753,N_17427);
nand U18482 (N_18482,N_17999,N_17729);
or U18483 (N_18483,N_17582,N_17446);
and U18484 (N_18484,N_17613,N_17855);
xor U18485 (N_18485,N_17674,N_17691);
xor U18486 (N_18486,N_17966,N_17736);
or U18487 (N_18487,N_17478,N_17844);
nor U18488 (N_18488,N_17469,N_17696);
nor U18489 (N_18489,N_17866,N_17637);
or U18490 (N_18490,N_17687,N_17912);
nor U18491 (N_18491,N_17515,N_17674);
and U18492 (N_18492,N_17798,N_17776);
xor U18493 (N_18493,N_17766,N_17615);
xnor U18494 (N_18494,N_17605,N_17533);
nor U18495 (N_18495,N_17695,N_17879);
nor U18496 (N_18496,N_17503,N_17955);
or U18497 (N_18497,N_17733,N_17964);
nand U18498 (N_18498,N_17763,N_17823);
xor U18499 (N_18499,N_17755,N_17743);
nand U18500 (N_18500,N_17899,N_17642);
nand U18501 (N_18501,N_17568,N_17653);
nor U18502 (N_18502,N_17666,N_17565);
or U18503 (N_18503,N_17497,N_17428);
and U18504 (N_18504,N_17657,N_17454);
and U18505 (N_18505,N_17466,N_17419);
and U18506 (N_18506,N_17808,N_17463);
xor U18507 (N_18507,N_17839,N_17668);
nor U18508 (N_18508,N_17456,N_17534);
and U18509 (N_18509,N_17740,N_17723);
xor U18510 (N_18510,N_17760,N_17855);
or U18511 (N_18511,N_17942,N_17484);
or U18512 (N_18512,N_17412,N_17830);
nand U18513 (N_18513,N_17587,N_17983);
xor U18514 (N_18514,N_17492,N_17877);
and U18515 (N_18515,N_17646,N_17901);
or U18516 (N_18516,N_17484,N_17432);
and U18517 (N_18517,N_17903,N_17415);
or U18518 (N_18518,N_17673,N_17669);
and U18519 (N_18519,N_17857,N_17627);
and U18520 (N_18520,N_17923,N_17845);
or U18521 (N_18521,N_17411,N_17857);
xor U18522 (N_18522,N_17587,N_17917);
and U18523 (N_18523,N_17846,N_17489);
or U18524 (N_18524,N_17583,N_17507);
and U18525 (N_18525,N_17728,N_17931);
nor U18526 (N_18526,N_17609,N_17678);
xor U18527 (N_18527,N_17470,N_17489);
nand U18528 (N_18528,N_17773,N_17642);
xor U18529 (N_18529,N_17567,N_17665);
or U18530 (N_18530,N_17695,N_17498);
or U18531 (N_18531,N_17827,N_17519);
nand U18532 (N_18532,N_17711,N_17549);
and U18533 (N_18533,N_17750,N_17853);
xnor U18534 (N_18534,N_17788,N_17719);
or U18535 (N_18535,N_17708,N_17616);
xor U18536 (N_18536,N_17896,N_17639);
or U18537 (N_18537,N_17906,N_17888);
or U18538 (N_18538,N_17536,N_17595);
xor U18539 (N_18539,N_17715,N_17515);
or U18540 (N_18540,N_17406,N_17934);
or U18541 (N_18541,N_17915,N_17445);
or U18542 (N_18542,N_17992,N_17511);
nand U18543 (N_18543,N_17906,N_17964);
nor U18544 (N_18544,N_17719,N_17874);
or U18545 (N_18545,N_17795,N_17608);
nor U18546 (N_18546,N_17563,N_17506);
xnor U18547 (N_18547,N_17881,N_17430);
and U18548 (N_18548,N_17852,N_17521);
nand U18549 (N_18549,N_17642,N_17531);
nand U18550 (N_18550,N_17547,N_17671);
and U18551 (N_18551,N_17487,N_17877);
nor U18552 (N_18552,N_17892,N_17692);
or U18553 (N_18553,N_17690,N_17678);
nor U18554 (N_18554,N_17977,N_17781);
and U18555 (N_18555,N_17567,N_17732);
nor U18556 (N_18556,N_17802,N_17993);
and U18557 (N_18557,N_17843,N_17400);
xnor U18558 (N_18558,N_17468,N_17812);
nand U18559 (N_18559,N_17548,N_17472);
nor U18560 (N_18560,N_17569,N_17780);
nor U18561 (N_18561,N_17968,N_17892);
nor U18562 (N_18562,N_17677,N_17724);
or U18563 (N_18563,N_17815,N_17598);
xor U18564 (N_18564,N_17958,N_17835);
xnor U18565 (N_18565,N_17440,N_17892);
nand U18566 (N_18566,N_17910,N_17542);
xor U18567 (N_18567,N_17555,N_17926);
or U18568 (N_18568,N_17880,N_17438);
xnor U18569 (N_18569,N_17483,N_17459);
or U18570 (N_18570,N_17615,N_17524);
nor U18571 (N_18571,N_17861,N_17953);
nor U18572 (N_18572,N_17974,N_17954);
nand U18573 (N_18573,N_17956,N_17873);
xnor U18574 (N_18574,N_17410,N_17993);
nor U18575 (N_18575,N_17980,N_17612);
nor U18576 (N_18576,N_17653,N_17745);
xnor U18577 (N_18577,N_17636,N_17888);
xnor U18578 (N_18578,N_17931,N_17442);
or U18579 (N_18579,N_17421,N_17794);
and U18580 (N_18580,N_17999,N_17606);
nand U18581 (N_18581,N_17957,N_17999);
nand U18582 (N_18582,N_17553,N_17966);
nand U18583 (N_18583,N_17552,N_17994);
nand U18584 (N_18584,N_17475,N_17899);
or U18585 (N_18585,N_17500,N_17803);
nand U18586 (N_18586,N_17683,N_17690);
and U18587 (N_18587,N_17756,N_17827);
or U18588 (N_18588,N_17717,N_17616);
nand U18589 (N_18589,N_17640,N_17536);
nand U18590 (N_18590,N_17631,N_17489);
or U18591 (N_18591,N_17874,N_17751);
nor U18592 (N_18592,N_17557,N_17648);
nor U18593 (N_18593,N_17441,N_17861);
or U18594 (N_18594,N_17496,N_17991);
nand U18595 (N_18595,N_17701,N_17902);
xor U18596 (N_18596,N_17505,N_17587);
xor U18597 (N_18597,N_17928,N_17980);
nor U18598 (N_18598,N_17690,N_17609);
nor U18599 (N_18599,N_17725,N_17963);
or U18600 (N_18600,N_18142,N_18044);
xor U18601 (N_18601,N_18259,N_18129);
nor U18602 (N_18602,N_18458,N_18228);
nor U18603 (N_18603,N_18521,N_18094);
nor U18604 (N_18604,N_18515,N_18013);
nand U18605 (N_18605,N_18527,N_18053);
nor U18606 (N_18606,N_18092,N_18093);
or U18607 (N_18607,N_18191,N_18154);
nor U18608 (N_18608,N_18186,N_18100);
or U18609 (N_18609,N_18345,N_18274);
or U18610 (N_18610,N_18349,N_18353);
and U18611 (N_18611,N_18409,N_18153);
nand U18612 (N_18612,N_18238,N_18447);
xnor U18613 (N_18613,N_18315,N_18473);
or U18614 (N_18614,N_18309,N_18247);
xor U18615 (N_18615,N_18034,N_18120);
and U18616 (N_18616,N_18086,N_18384);
and U18617 (N_18617,N_18234,N_18256);
or U18618 (N_18618,N_18155,N_18331);
nor U18619 (N_18619,N_18198,N_18321);
nand U18620 (N_18620,N_18569,N_18314);
nand U18621 (N_18621,N_18004,N_18365);
or U18622 (N_18622,N_18324,N_18303);
xor U18623 (N_18623,N_18300,N_18399);
and U18624 (N_18624,N_18596,N_18209);
nand U18625 (N_18625,N_18114,N_18297);
nor U18626 (N_18626,N_18235,N_18284);
xor U18627 (N_18627,N_18449,N_18492);
nand U18628 (N_18628,N_18137,N_18403);
nand U18629 (N_18629,N_18337,N_18535);
or U18630 (N_18630,N_18549,N_18060);
or U18631 (N_18631,N_18022,N_18390);
and U18632 (N_18632,N_18266,N_18176);
nor U18633 (N_18633,N_18233,N_18488);
xor U18634 (N_18634,N_18199,N_18109);
nor U18635 (N_18635,N_18587,N_18222);
nor U18636 (N_18636,N_18215,N_18461);
nor U18637 (N_18637,N_18340,N_18428);
nand U18638 (N_18638,N_18431,N_18252);
xnor U18639 (N_18639,N_18419,N_18372);
or U18640 (N_18640,N_18224,N_18019);
nand U18641 (N_18641,N_18205,N_18217);
xor U18642 (N_18642,N_18071,N_18378);
and U18643 (N_18643,N_18302,N_18000);
and U18644 (N_18644,N_18460,N_18091);
nor U18645 (N_18645,N_18166,N_18508);
or U18646 (N_18646,N_18267,N_18575);
nand U18647 (N_18647,N_18469,N_18318);
nand U18648 (N_18648,N_18089,N_18420);
nand U18649 (N_18649,N_18594,N_18240);
or U18650 (N_18650,N_18454,N_18127);
and U18651 (N_18651,N_18167,N_18369);
nor U18652 (N_18652,N_18021,N_18572);
and U18653 (N_18653,N_18212,N_18566);
xor U18654 (N_18654,N_18286,N_18326);
and U18655 (N_18655,N_18255,N_18463);
and U18656 (N_18656,N_18119,N_18292);
nand U18657 (N_18657,N_18573,N_18253);
nand U18658 (N_18658,N_18505,N_18531);
or U18659 (N_18659,N_18568,N_18437);
and U18660 (N_18660,N_18328,N_18008);
or U18661 (N_18661,N_18017,N_18588);
nand U18662 (N_18662,N_18544,N_18424);
nand U18663 (N_18663,N_18481,N_18136);
and U18664 (N_18664,N_18181,N_18035);
xor U18665 (N_18665,N_18502,N_18095);
or U18666 (N_18666,N_18452,N_18069);
nand U18667 (N_18667,N_18557,N_18225);
xnor U18668 (N_18668,N_18160,N_18223);
or U18669 (N_18669,N_18582,N_18564);
and U18670 (N_18670,N_18581,N_18497);
xnor U18671 (N_18671,N_18580,N_18418);
nor U18672 (N_18672,N_18417,N_18386);
and U18673 (N_18673,N_18362,N_18107);
and U18674 (N_18674,N_18106,N_18422);
nor U18675 (N_18675,N_18056,N_18509);
nand U18676 (N_18676,N_18304,N_18049);
and U18677 (N_18677,N_18382,N_18257);
nand U18678 (N_18678,N_18131,N_18501);
or U18679 (N_18679,N_18174,N_18472);
and U18680 (N_18680,N_18516,N_18457);
or U18681 (N_18681,N_18207,N_18595);
or U18682 (N_18682,N_18051,N_18026);
or U18683 (N_18683,N_18015,N_18058);
or U18684 (N_18684,N_18159,N_18426);
or U18685 (N_18685,N_18081,N_18172);
or U18686 (N_18686,N_18411,N_18339);
xor U18687 (N_18687,N_18263,N_18366);
nand U18688 (N_18688,N_18230,N_18029);
or U18689 (N_18689,N_18294,N_18565);
nand U18690 (N_18690,N_18202,N_18306);
or U18691 (N_18691,N_18296,N_18393);
or U18692 (N_18692,N_18003,N_18299);
and U18693 (N_18693,N_18206,N_18322);
nand U18694 (N_18694,N_18520,N_18559);
or U18695 (N_18695,N_18162,N_18031);
or U18696 (N_18696,N_18561,N_18512);
nor U18697 (N_18697,N_18313,N_18542);
xnor U18698 (N_18698,N_18168,N_18145);
nor U18699 (N_18699,N_18088,N_18057);
or U18700 (N_18700,N_18291,N_18141);
or U18701 (N_18701,N_18389,N_18175);
nor U18702 (N_18702,N_18478,N_18597);
or U18703 (N_18703,N_18523,N_18405);
nand U18704 (N_18704,N_18138,N_18090);
nor U18705 (N_18705,N_18487,N_18196);
or U18706 (N_18706,N_18351,N_18537);
or U18707 (N_18707,N_18485,N_18524);
nor U18708 (N_18708,N_18045,N_18179);
xnor U18709 (N_18709,N_18165,N_18396);
and U18710 (N_18710,N_18506,N_18379);
xor U18711 (N_18711,N_18112,N_18260);
or U18712 (N_18712,N_18002,N_18585);
or U18713 (N_18713,N_18357,N_18128);
or U18714 (N_18714,N_18268,N_18493);
or U18715 (N_18715,N_18038,N_18083);
nand U18716 (N_18716,N_18342,N_18538);
and U18717 (N_18717,N_18183,N_18539);
or U18718 (N_18718,N_18133,N_18147);
xnor U18719 (N_18719,N_18262,N_18555);
nor U18720 (N_18720,N_18105,N_18586);
or U18721 (N_18721,N_18061,N_18012);
and U18722 (N_18722,N_18011,N_18320);
nand U18723 (N_18723,N_18062,N_18099);
nand U18724 (N_18724,N_18475,N_18344);
and U18725 (N_18725,N_18020,N_18468);
xor U18726 (N_18726,N_18173,N_18408);
xor U18727 (N_18727,N_18059,N_18474);
xor U18728 (N_18728,N_18376,N_18360);
nor U18729 (N_18729,N_18041,N_18148);
xor U18730 (N_18730,N_18006,N_18213);
nor U18731 (N_18731,N_18080,N_18562);
and U18732 (N_18732,N_18067,N_18157);
and U18733 (N_18733,N_18325,N_18514);
or U18734 (N_18734,N_18152,N_18383);
nand U18735 (N_18735,N_18395,N_18385);
nand U18736 (N_18736,N_18423,N_18227);
and U18737 (N_18737,N_18115,N_18295);
nand U18738 (N_18738,N_18150,N_18079);
nand U18739 (N_18739,N_18364,N_18536);
or U18740 (N_18740,N_18510,N_18436);
and U18741 (N_18741,N_18250,N_18278);
or U18742 (N_18742,N_18484,N_18214);
or U18743 (N_18743,N_18400,N_18289);
nor U18744 (N_18744,N_18526,N_18052);
and U18745 (N_18745,N_18550,N_18308);
nor U18746 (N_18746,N_18576,N_18182);
nor U18747 (N_18747,N_18108,N_18343);
nor U18748 (N_18748,N_18415,N_18073);
and U18749 (N_18749,N_18498,N_18158);
xnor U18750 (N_18750,N_18459,N_18525);
nor U18751 (N_18751,N_18243,N_18195);
and U18752 (N_18752,N_18221,N_18504);
and U18753 (N_18753,N_18097,N_18528);
xor U18754 (N_18754,N_18476,N_18254);
nor U18755 (N_18755,N_18290,N_18305);
or U18756 (N_18756,N_18054,N_18047);
nor U18757 (N_18757,N_18394,N_18567);
xor U18758 (N_18758,N_18219,N_18477);
xnor U18759 (N_18759,N_18470,N_18401);
and U18760 (N_18760,N_18113,N_18123);
xnor U18761 (N_18761,N_18229,N_18551);
nand U18762 (N_18762,N_18126,N_18189);
or U18763 (N_18763,N_18014,N_18251);
nand U18764 (N_18764,N_18592,N_18453);
nand U18765 (N_18765,N_18332,N_18194);
xnor U18766 (N_18766,N_18450,N_18354);
nor U18767 (N_18767,N_18370,N_18282);
xnor U18768 (N_18768,N_18293,N_18007);
or U18769 (N_18769,N_18517,N_18201);
xnor U18770 (N_18770,N_18009,N_18547);
xnor U18771 (N_18771,N_18216,N_18132);
and U18772 (N_18772,N_18023,N_18483);
nor U18773 (N_18773,N_18244,N_18499);
or U18774 (N_18774,N_18388,N_18495);
xnor U18775 (N_18775,N_18018,N_18334);
nor U18776 (N_18776,N_18048,N_18046);
nor U18777 (N_18777,N_18279,N_18430);
or U18778 (N_18778,N_18203,N_18287);
and U18779 (N_18779,N_18432,N_18110);
or U18780 (N_18780,N_18211,N_18248);
and U18781 (N_18781,N_18451,N_18116);
nand U18782 (N_18782,N_18170,N_18435);
or U18783 (N_18783,N_18464,N_18117);
nor U18784 (N_18784,N_18348,N_18479);
and U18785 (N_18785,N_18103,N_18532);
nand U18786 (N_18786,N_18563,N_18489);
nand U18787 (N_18787,N_18271,N_18433);
and U18788 (N_18788,N_18371,N_18169);
nand U18789 (N_18789,N_18496,N_18231);
and U18790 (N_18790,N_18118,N_18121);
nor U18791 (N_18791,N_18513,N_18429);
nand U18792 (N_18792,N_18494,N_18491);
or U18793 (N_18793,N_18301,N_18135);
xor U18794 (N_18794,N_18024,N_18414);
nand U18795 (N_18795,N_18346,N_18226);
xnor U18796 (N_18796,N_18070,N_18543);
and U18797 (N_18797,N_18560,N_18218);
or U18798 (N_18798,N_18055,N_18361);
or U18799 (N_18799,N_18327,N_18553);
xor U18800 (N_18800,N_18462,N_18124);
nand U18801 (N_18801,N_18406,N_18591);
xnor U18802 (N_18802,N_18578,N_18574);
and U18803 (N_18803,N_18448,N_18085);
and U18804 (N_18804,N_18028,N_18471);
nand U18805 (N_18805,N_18347,N_18465);
nand U18806 (N_18806,N_18040,N_18518);
xor U18807 (N_18807,N_18249,N_18590);
nand U18808 (N_18808,N_18375,N_18579);
and U18809 (N_18809,N_18446,N_18584);
nand U18810 (N_18810,N_18261,N_18554);
and U18811 (N_18811,N_18074,N_18455);
or U18812 (N_18812,N_18140,N_18534);
and U18813 (N_18813,N_18507,N_18210);
nand U18814 (N_18814,N_18500,N_18016);
or U18815 (N_18815,N_18335,N_18010);
or U18816 (N_18816,N_18397,N_18533);
nand U18817 (N_18817,N_18025,N_18078);
nand U18818 (N_18818,N_18355,N_18096);
nor U18819 (N_18819,N_18404,N_18410);
xor U18820 (N_18820,N_18341,N_18593);
xnor U18821 (N_18821,N_18063,N_18380);
nor U18822 (N_18822,N_18374,N_18519);
and U18823 (N_18823,N_18391,N_18077);
nor U18824 (N_18824,N_18276,N_18529);
nand U18825 (N_18825,N_18005,N_18076);
nand U18826 (N_18826,N_18033,N_18050);
and U18827 (N_18827,N_18545,N_18144);
xnor U18828 (N_18828,N_18264,N_18193);
xnor U18829 (N_18829,N_18336,N_18358);
or U18830 (N_18830,N_18456,N_18571);
nor U18831 (N_18831,N_18001,N_18204);
or U18832 (N_18832,N_18356,N_18317);
nor U18833 (N_18833,N_18098,N_18281);
nor U18834 (N_18834,N_18541,N_18438);
nand U18835 (N_18835,N_18270,N_18556);
nand U18836 (N_18836,N_18552,N_18042);
nor U18837 (N_18837,N_18398,N_18246);
and U18838 (N_18838,N_18241,N_18307);
nor U18839 (N_18839,N_18323,N_18272);
and U18840 (N_18840,N_18285,N_18589);
nand U18841 (N_18841,N_18283,N_18540);
xnor U18842 (N_18842,N_18333,N_18583);
nand U18843 (N_18843,N_18548,N_18220);
xnor U18844 (N_18844,N_18407,N_18066);
and U18845 (N_18845,N_18237,N_18275);
and U18846 (N_18846,N_18139,N_18269);
nor U18847 (N_18847,N_18319,N_18032);
or U18848 (N_18848,N_18197,N_18503);
xor U18849 (N_18849,N_18443,N_18363);
and U18850 (N_18850,N_18442,N_18082);
and U18851 (N_18851,N_18122,N_18072);
and U18852 (N_18852,N_18316,N_18480);
nor U18853 (N_18853,N_18352,N_18163);
or U18854 (N_18854,N_18558,N_18427);
and U18855 (N_18855,N_18570,N_18373);
and U18856 (N_18856,N_18413,N_18037);
nor U18857 (N_18857,N_18402,N_18392);
xor U18858 (N_18858,N_18288,N_18530);
or U18859 (N_18859,N_18482,N_18329);
xnor U18860 (N_18860,N_18187,N_18101);
nor U18861 (N_18861,N_18265,N_18421);
nor U18862 (N_18862,N_18164,N_18068);
nand U18863 (N_18863,N_18143,N_18125);
and U18864 (N_18864,N_18273,N_18312);
nor U18865 (N_18865,N_18208,N_18546);
xnor U18866 (N_18866,N_18030,N_18185);
and U18867 (N_18867,N_18036,N_18084);
nand U18868 (N_18868,N_18245,N_18440);
and U18869 (N_18869,N_18258,N_18280);
nor U18870 (N_18870,N_18330,N_18134);
nor U18871 (N_18871,N_18367,N_18146);
xor U18872 (N_18872,N_18177,N_18425);
nand U18873 (N_18873,N_18445,N_18599);
and U18874 (N_18874,N_18242,N_18466);
or U18875 (N_18875,N_18161,N_18467);
xor U18876 (N_18876,N_18239,N_18277);
xnor U18877 (N_18877,N_18387,N_18104);
nand U18878 (N_18878,N_18439,N_18178);
and U18879 (N_18879,N_18111,N_18156);
xor U18880 (N_18880,N_18412,N_18490);
or U18881 (N_18881,N_18102,N_18190);
or U18882 (N_18882,N_18377,N_18311);
and U18883 (N_18883,N_18368,N_18180);
and U18884 (N_18884,N_18151,N_18192);
nand U18885 (N_18885,N_18200,N_18027);
xor U18886 (N_18886,N_18065,N_18171);
or U18887 (N_18887,N_18039,N_18064);
and U18888 (N_18888,N_18522,N_18381);
xnor U18889 (N_18889,N_18298,N_18184);
nor U18890 (N_18890,N_18130,N_18087);
nand U18891 (N_18891,N_18338,N_18511);
nand U18892 (N_18892,N_18577,N_18359);
nand U18893 (N_18893,N_18486,N_18075);
xor U18894 (N_18894,N_18441,N_18416);
or U18895 (N_18895,N_18350,N_18043);
nor U18896 (N_18896,N_18310,N_18236);
nor U18897 (N_18897,N_18232,N_18188);
xnor U18898 (N_18898,N_18434,N_18444);
xnor U18899 (N_18899,N_18598,N_18149);
and U18900 (N_18900,N_18280,N_18297);
and U18901 (N_18901,N_18151,N_18120);
nand U18902 (N_18902,N_18411,N_18365);
nor U18903 (N_18903,N_18227,N_18082);
xnor U18904 (N_18904,N_18077,N_18245);
and U18905 (N_18905,N_18158,N_18115);
xnor U18906 (N_18906,N_18061,N_18178);
nor U18907 (N_18907,N_18052,N_18304);
or U18908 (N_18908,N_18375,N_18396);
or U18909 (N_18909,N_18350,N_18303);
or U18910 (N_18910,N_18002,N_18077);
nand U18911 (N_18911,N_18372,N_18026);
nand U18912 (N_18912,N_18404,N_18369);
xor U18913 (N_18913,N_18038,N_18265);
and U18914 (N_18914,N_18217,N_18498);
nand U18915 (N_18915,N_18101,N_18033);
nor U18916 (N_18916,N_18376,N_18587);
xor U18917 (N_18917,N_18344,N_18034);
nand U18918 (N_18918,N_18442,N_18583);
or U18919 (N_18919,N_18327,N_18068);
nand U18920 (N_18920,N_18095,N_18008);
nand U18921 (N_18921,N_18315,N_18094);
nor U18922 (N_18922,N_18520,N_18385);
or U18923 (N_18923,N_18149,N_18410);
or U18924 (N_18924,N_18500,N_18110);
nor U18925 (N_18925,N_18361,N_18075);
or U18926 (N_18926,N_18369,N_18597);
xor U18927 (N_18927,N_18085,N_18501);
or U18928 (N_18928,N_18497,N_18567);
xnor U18929 (N_18929,N_18354,N_18493);
nand U18930 (N_18930,N_18011,N_18518);
and U18931 (N_18931,N_18354,N_18242);
or U18932 (N_18932,N_18343,N_18302);
and U18933 (N_18933,N_18209,N_18415);
or U18934 (N_18934,N_18341,N_18424);
xnor U18935 (N_18935,N_18127,N_18285);
and U18936 (N_18936,N_18214,N_18530);
and U18937 (N_18937,N_18230,N_18473);
xnor U18938 (N_18938,N_18097,N_18347);
xor U18939 (N_18939,N_18387,N_18468);
xnor U18940 (N_18940,N_18227,N_18375);
or U18941 (N_18941,N_18408,N_18295);
or U18942 (N_18942,N_18313,N_18409);
and U18943 (N_18943,N_18575,N_18541);
and U18944 (N_18944,N_18456,N_18343);
xnor U18945 (N_18945,N_18325,N_18075);
or U18946 (N_18946,N_18056,N_18278);
and U18947 (N_18947,N_18138,N_18401);
or U18948 (N_18948,N_18079,N_18218);
or U18949 (N_18949,N_18352,N_18235);
or U18950 (N_18950,N_18087,N_18093);
and U18951 (N_18951,N_18256,N_18403);
nand U18952 (N_18952,N_18329,N_18415);
and U18953 (N_18953,N_18465,N_18390);
nand U18954 (N_18954,N_18170,N_18427);
nand U18955 (N_18955,N_18016,N_18134);
nor U18956 (N_18956,N_18299,N_18422);
nand U18957 (N_18957,N_18563,N_18338);
nand U18958 (N_18958,N_18403,N_18217);
and U18959 (N_18959,N_18551,N_18330);
or U18960 (N_18960,N_18089,N_18072);
or U18961 (N_18961,N_18391,N_18117);
nand U18962 (N_18962,N_18268,N_18481);
xor U18963 (N_18963,N_18035,N_18534);
nor U18964 (N_18964,N_18057,N_18045);
or U18965 (N_18965,N_18405,N_18505);
nor U18966 (N_18966,N_18447,N_18502);
nor U18967 (N_18967,N_18594,N_18444);
nand U18968 (N_18968,N_18073,N_18027);
or U18969 (N_18969,N_18121,N_18427);
xor U18970 (N_18970,N_18169,N_18440);
and U18971 (N_18971,N_18495,N_18305);
nand U18972 (N_18972,N_18388,N_18586);
and U18973 (N_18973,N_18598,N_18044);
nor U18974 (N_18974,N_18174,N_18461);
nor U18975 (N_18975,N_18561,N_18533);
or U18976 (N_18976,N_18556,N_18149);
or U18977 (N_18977,N_18556,N_18565);
or U18978 (N_18978,N_18531,N_18090);
nor U18979 (N_18979,N_18071,N_18280);
nor U18980 (N_18980,N_18551,N_18461);
nor U18981 (N_18981,N_18363,N_18084);
nor U18982 (N_18982,N_18080,N_18598);
or U18983 (N_18983,N_18325,N_18311);
or U18984 (N_18984,N_18237,N_18143);
or U18985 (N_18985,N_18541,N_18027);
or U18986 (N_18986,N_18597,N_18588);
nor U18987 (N_18987,N_18262,N_18389);
or U18988 (N_18988,N_18182,N_18180);
or U18989 (N_18989,N_18004,N_18257);
and U18990 (N_18990,N_18235,N_18477);
xnor U18991 (N_18991,N_18201,N_18411);
nor U18992 (N_18992,N_18329,N_18131);
and U18993 (N_18993,N_18016,N_18333);
xnor U18994 (N_18994,N_18096,N_18568);
nand U18995 (N_18995,N_18458,N_18451);
xor U18996 (N_18996,N_18581,N_18571);
nor U18997 (N_18997,N_18530,N_18291);
xnor U18998 (N_18998,N_18198,N_18016);
xor U18999 (N_18999,N_18263,N_18347);
and U19000 (N_19000,N_18374,N_18024);
nor U19001 (N_19001,N_18340,N_18532);
and U19002 (N_19002,N_18572,N_18372);
xor U19003 (N_19003,N_18317,N_18119);
nor U19004 (N_19004,N_18217,N_18225);
nor U19005 (N_19005,N_18429,N_18258);
nor U19006 (N_19006,N_18510,N_18435);
nand U19007 (N_19007,N_18054,N_18102);
nand U19008 (N_19008,N_18425,N_18125);
or U19009 (N_19009,N_18105,N_18481);
or U19010 (N_19010,N_18516,N_18430);
nand U19011 (N_19011,N_18341,N_18458);
or U19012 (N_19012,N_18172,N_18470);
xor U19013 (N_19013,N_18016,N_18306);
and U19014 (N_19014,N_18568,N_18294);
or U19015 (N_19015,N_18492,N_18561);
xor U19016 (N_19016,N_18546,N_18575);
and U19017 (N_19017,N_18311,N_18051);
and U19018 (N_19018,N_18194,N_18285);
or U19019 (N_19019,N_18223,N_18342);
or U19020 (N_19020,N_18073,N_18245);
nor U19021 (N_19021,N_18199,N_18553);
nor U19022 (N_19022,N_18318,N_18073);
nor U19023 (N_19023,N_18097,N_18145);
nor U19024 (N_19024,N_18059,N_18121);
nand U19025 (N_19025,N_18262,N_18585);
xor U19026 (N_19026,N_18276,N_18178);
and U19027 (N_19027,N_18234,N_18426);
nor U19028 (N_19028,N_18137,N_18474);
nor U19029 (N_19029,N_18566,N_18051);
and U19030 (N_19030,N_18299,N_18412);
or U19031 (N_19031,N_18191,N_18160);
and U19032 (N_19032,N_18590,N_18079);
nor U19033 (N_19033,N_18182,N_18446);
nor U19034 (N_19034,N_18019,N_18511);
nor U19035 (N_19035,N_18076,N_18178);
nand U19036 (N_19036,N_18154,N_18179);
nand U19037 (N_19037,N_18031,N_18511);
and U19038 (N_19038,N_18320,N_18415);
xor U19039 (N_19039,N_18285,N_18153);
xor U19040 (N_19040,N_18305,N_18516);
nand U19041 (N_19041,N_18559,N_18460);
nand U19042 (N_19042,N_18142,N_18120);
xor U19043 (N_19043,N_18134,N_18037);
nand U19044 (N_19044,N_18160,N_18384);
nand U19045 (N_19045,N_18548,N_18285);
xor U19046 (N_19046,N_18197,N_18026);
and U19047 (N_19047,N_18336,N_18126);
and U19048 (N_19048,N_18311,N_18599);
nand U19049 (N_19049,N_18266,N_18504);
xor U19050 (N_19050,N_18090,N_18196);
xnor U19051 (N_19051,N_18530,N_18140);
or U19052 (N_19052,N_18092,N_18294);
or U19053 (N_19053,N_18315,N_18596);
and U19054 (N_19054,N_18342,N_18097);
nand U19055 (N_19055,N_18500,N_18561);
nor U19056 (N_19056,N_18565,N_18472);
nor U19057 (N_19057,N_18341,N_18573);
xor U19058 (N_19058,N_18208,N_18411);
nand U19059 (N_19059,N_18547,N_18239);
and U19060 (N_19060,N_18531,N_18229);
nand U19061 (N_19061,N_18585,N_18432);
nand U19062 (N_19062,N_18197,N_18105);
or U19063 (N_19063,N_18369,N_18478);
xor U19064 (N_19064,N_18594,N_18171);
nor U19065 (N_19065,N_18070,N_18038);
nor U19066 (N_19066,N_18155,N_18391);
xnor U19067 (N_19067,N_18599,N_18233);
and U19068 (N_19068,N_18455,N_18356);
nand U19069 (N_19069,N_18121,N_18143);
and U19070 (N_19070,N_18338,N_18225);
or U19071 (N_19071,N_18363,N_18319);
nand U19072 (N_19072,N_18217,N_18507);
or U19073 (N_19073,N_18216,N_18195);
nor U19074 (N_19074,N_18156,N_18110);
nand U19075 (N_19075,N_18014,N_18156);
and U19076 (N_19076,N_18099,N_18092);
nand U19077 (N_19077,N_18100,N_18064);
xnor U19078 (N_19078,N_18165,N_18027);
or U19079 (N_19079,N_18499,N_18305);
or U19080 (N_19080,N_18454,N_18389);
nor U19081 (N_19081,N_18070,N_18238);
nor U19082 (N_19082,N_18181,N_18536);
nand U19083 (N_19083,N_18238,N_18246);
xor U19084 (N_19084,N_18517,N_18485);
and U19085 (N_19085,N_18240,N_18203);
or U19086 (N_19086,N_18027,N_18161);
xnor U19087 (N_19087,N_18501,N_18075);
and U19088 (N_19088,N_18520,N_18222);
or U19089 (N_19089,N_18365,N_18091);
nor U19090 (N_19090,N_18583,N_18210);
nor U19091 (N_19091,N_18276,N_18342);
nand U19092 (N_19092,N_18590,N_18411);
or U19093 (N_19093,N_18294,N_18150);
and U19094 (N_19094,N_18036,N_18394);
and U19095 (N_19095,N_18019,N_18201);
and U19096 (N_19096,N_18217,N_18576);
nand U19097 (N_19097,N_18314,N_18182);
xor U19098 (N_19098,N_18566,N_18105);
nand U19099 (N_19099,N_18117,N_18349);
and U19100 (N_19100,N_18462,N_18260);
nand U19101 (N_19101,N_18372,N_18364);
nand U19102 (N_19102,N_18288,N_18008);
or U19103 (N_19103,N_18392,N_18422);
xor U19104 (N_19104,N_18421,N_18097);
and U19105 (N_19105,N_18495,N_18216);
and U19106 (N_19106,N_18049,N_18580);
nor U19107 (N_19107,N_18278,N_18120);
nor U19108 (N_19108,N_18171,N_18148);
nor U19109 (N_19109,N_18540,N_18418);
or U19110 (N_19110,N_18001,N_18561);
xor U19111 (N_19111,N_18053,N_18378);
or U19112 (N_19112,N_18415,N_18064);
or U19113 (N_19113,N_18459,N_18512);
xor U19114 (N_19114,N_18180,N_18283);
and U19115 (N_19115,N_18496,N_18555);
nor U19116 (N_19116,N_18162,N_18033);
and U19117 (N_19117,N_18136,N_18578);
or U19118 (N_19118,N_18063,N_18141);
nor U19119 (N_19119,N_18093,N_18342);
and U19120 (N_19120,N_18327,N_18514);
or U19121 (N_19121,N_18179,N_18364);
xnor U19122 (N_19122,N_18279,N_18116);
or U19123 (N_19123,N_18240,N_18056);
nand U19124 (N_19124,N_18081,N_18307);
nor U19125 (N_19125,N_18501,N_18496);
nand U19126 (N_19126,N_18078,N_18492);
or U19127 (N_19127,N_18544,N_18481);
xor U19128 (N_19128,N_18504,N_18223);
or U19129 (N_19129,N_18231,N_18099);
nor U19130 (N_19130,N_18524,N_18380);
xor U19131 (N_19131,N_18537,N_18013);
nor U19132 (N_19132,N_18324,N_18086);
xor U19133 (N_19133,N_18107,N_18522);
xor U19134 (N_19134,N_18005,N_18388);
xor U19135 (N_19135,N_18286,N_18263);
or U19136 (N_19136,N_18317,N_18086);
nand U19137 (N_19137,N_18152,N_18513);
and U19138 (N_19138,N_18576,N_18528);
nand U19139 (N_19139,N_18511,N_18092);
and U19140 (N_19140,N_18236,N_18487);
nor U19141 (N_19141,N_18137,N_18029);
nand U19142 (N_19142,N_18511,N_18155);
nor U19143 (N_19143,N_18277,N_18078);
nor U19144 (N_19144,N_18316,N_18044);
xor U19145 (N_19145,N_18521,N_18539);
and U19146 (N_19146,N_18283,N_18550);
and U19147 (N_19147,N_18302,N_18341);
and U19148 (N_19148,N_18127,N_18070);
nand U19149 (N_19149,N_18059,N_18397);
and U19150 (N_19150,N_18201,N_18135);
xor U19151 (N_19151,N_18444,N_18483);
and U19152 (N_19152,N_18175,N_18145);
xnor U19153 (N_19153,N_18152,N_18084);
xnor U19154 (N_19154,N_18334,N_18214);
nor U19155 (N_19155,N_18590,N_18225);
nor U19156 (N_19156,N_18455,N_18425);
xor U19157 (N_19157,N_18202,N_18116);
xnor U19158 (N_19158,N_18559,N_18534);
nand U19159 (N_19159,N_18295,N_18149);
or U19160 (N_19160,N_18366,N_18147);
and U19161 (N_19161,N_18065,N_18244);
nand U19162 (N_19162,N_18108,N_18149);
nor U19163 (N_19163,N_18032,N_18078);
or U19164 (N_19164,N_18081,N_18454);
or U19165 (N_19165,N_18337,N_18409);
xor U19166 (N_19166,N_18470,N_18321);
xnor U19167 (N_19167,N_18351,N_18278);
and U19168 (N_19168,N_18554,N_18106);
nor U19169 (N_19169,N_18539,N_18347);
nor U19170 (N_19170,N_18461,N_18434);
nand U19171 (N_19171,N_18544,N_18588);
nor U19172 (N_19172,N_18331,N_18191);
nor U19173 (N_19173,N_18069,N_18599);
or U19174 (N_19174,N_18250,N_18507);
xor U19175 (N_19175,N_18152,N_18246);
and U19176 (N_19176,N_18054,N_18218);
and U19177 (N_19177,N_18363,N_18020);
and U19178 (N_19178,N_18265,N_18223);
or U19179 (N_19179,N_18496,N_18099);
and U19180 (N_19180,N_18267,N_18492);
or U19181 (N_19181,N_18338,N_18548);
nor U19182 (N_19182,N_18126,N_18182);
nand U19183 (N_19183,N_18472,N_18422);
xnor U19184 (N_19184,N_18448,N_18142);
and U19185 (N_19185,N_18521,N_18380);
and U19186 (N_19186,N_18395,N_18147);
or U19187 (N_19187,N_18021,N_18576);
nand U19188 (N_19188,N_18487,N_18315);
and U19189 (N_19189,N_18054,N_18093);
xnor U19190 (N_19190,N_18225,N_18332);
or U19191 (N_19191,N_18276,N_18066);
nor U19192 (N_19192,N_18259,N_18441);
nand U19193 (N_19193,N_18321,N_18073);
xor U19194 (N_19194,N_18025,N_18067);
nand U19195 (N_19195,N_18236,N_18220);
nand U19196 (N_19196,N_18507,N_18405);
or U19197 (N_19197,N_18463,N_18115);
or U19198 (N_19198,N_18401,N_18574);
or U19199 (N_19199,N_18048,N_18467);
nand U19200 (N_19200,N_18712,N_18985);
nor U19201 (N_19201,N_19178,N_18650);
nor U19202 (N_19202,N_19199,N_18927);
xor U19203 (N_19203,N_19173,N_18735);
nor U19204 (N_19204,N_18673,N_19097);
nor U19205 (N_19205,N_18924,N_18696);
or U19206 (N_19206,N_18617,N_18666);
and U19207 (N_19207,N_18640,N_18866);
nor U19208 (N_19208,N_18728,N_18815);
or U19209 (N_19209,N_18723,N_19043);
and U19210 (N_19210,N_18615,N_19102);
nor U19211 (N_19211,N_18945,N_18779);
nor U19212 (N_19212,N_19040,N_18767);
or U19213 (N_19213,N_18995,N_18901);
nor U19214 (N_19214,N_19164,N_19091);
nor U19215 (N_19215,N_18755,N_18722);
nand U19216 (N_19216,N_18870,N_19026);
nor U19217 (N_19217,N_18873,N_18987);
nor U19218 (N_19218,N_18678,N_18794);
or U19219 (N_19219,N_18654,N_18918);
nand U19220 (N_19220,N_18928,N_18768);
and U19221 (N_19221,N_19099,N_18684);
and U19222 (N_19222,N_19068,N_18796);
nor U19223 (N_19223,N_19060,N_19001);
xnor U19224 (N_19224,N_18705,N_18810);
xnor U19225 (N_19225,N_18703,N_18816);
or U19226 (N_19226,N_18833,N_18829);
nor U19227 (N_19227,N_19193,N_18659);
or U19228 (N_19228,N_18981,N_19019);
or U19229 (N_19229,N_18975,N_18885);
xnor U19230 (N_19230,N_18902,N_18900);
xor U19231 (N_19231,N_18633,N_18936);
or U19232 (N_19232,N_18840,N_19184);
and U19233 (N_19233,N_19035,N_18955);
and U19234 (N_19234,N_19034,N_19196);
nor U19235 (N_19235,N_18940,N_18921);
nor U19236 (N_19236,N_18807,N_18871);
nor U19237 (N_19237,N_18908,N_19195);
or U19238 (N_19238,N_18999,N_18627);
or U19239 (N_19239,N_18716,N_19123);
or U19240 (N_19240,N_19122,N_18973);
and U19241 (N_19241,N_18930,N_18874);
nand U19242 (N_19242,N_18729,N_18911);
xor U19243 (N_19243,N_18806,N_19053);
nand U19244 (N_19244,N_18850,N_18687);
nand U19245 (N_19245,N_19139,N_18667);
and U19246 (N_19246,N_18878,N_18753);
nand U19247 (N_19247,N_18883,N_18663);
xnor U19248 (N_19248,N_19025,N_19046);
or U19249 (N_19249,N_18621,N_19065);
xor U19250 (N_19250,N_18637,N_18763);
nand U19251 (N_19251,N_19084,N_18731);
and U19252 (N_19252,N_18819,N_19114);
or U19253 (N_19253,N_19179,N_19156);
nand U19254 (N_19254,N_19175,N_19130);
nand U19255 (N_19255,N_18744,N_18649);
and U19256 (N_19256,N_18718,N_19031);
and U19257 (N_19257,N_19090,N_18826);
nor U19258 (N_19258,N_18830,N_18896);
and U19259 (N_19259,N_18891,N_18745);
nor U19260 (N_19260,N_18675,N_18674);
xor U19261 (N_19261,N_18959,N_18837);
nand U19262 (N_19262,N_18604,N_18888);
and U19263 (N_19263,N_19141,N_18876);
nor U19264 (N_19264,N_18892,N_18784);
nor U19265 (N_19265,N_19182,N_18620);
nand U19266 (N_19266,N_19100,N_19168);
nor U19267 (N_19267,N_18761,N_18766);
xor U19268 (N_19268,N_18726,N_19048);
xor U19269 (N_19269,N_18855,N_19128);
and U19270 (N_19270,N_18827,N_19144);
or U19271 (N_19271,N_18715,N_18904);
and U19272 (N_19272,N_18694,N_19057);
or U19273 (N_19273,N_18710,N_18968);
or U19274 (N_19274,N_18798,N_19028);
xor U19275 (N_19275,N_19021,N_19143);
nand U19276 (N_19276,N_19094,N_18656);
nand U19277 (N_19277,N_18626,N_19154);
or U19278 (N_19278,N_18944,N_18998);
or U19279 (N_19279,N_18939,N_18732);
nor U19280 (N_19280,N_18747,N_19160);
or U19281 (N_19281,N_18811,N_19105);
nand U19282 (N_19282,N_18630,N_19085);
nand U19283 (N_19283,N_18812,N_18702);
xnor U19284 (N_19284,N_19096,N_18856);
or U19285 (N_19285,N_19089,N_18844);
or U19286 (N_19286,N_18781,N_19172);
nand U19287 (N_19287,N_18823,N_18967);
nor U19288 (N_19288,N_19003,N_18990);
xnor U19289 (N_19289,N_18882,N_18771);
xor U19290 (N_19290,N_18601,N_19066);
xnor U19291 (N_19291,N_18865,N_19133);
xor U19292 (N_19292,N_19024,N_19063);
and U19293 (N_19293,N_18841,N_19146);
nor U19294 (N_19294,N_19008,N_19189);
nor U19295 (N_19295,N_18954,N_19135);
or U19296 (N_19296,N_18943,N_18651);
xnor U19297 (N_19297,N_18616,N_18776);
or U19298 (N_19298,N_19118,N_18629);
nand U19299 (N_19299,N_19159,N_19157);
nor U19300 (N_19300,N_18748,N_18724);
nor U19301 (N_19301,N_19076,N_18734);
xnor U19302 (N_19302,N_19132,N_18680);
nor U19303 (N_19303,N_18926,N_19072);
or U19304 (N_19304,N_18802,N_19032);
and U19305 (N_19305,N_18752,N_18609);
and U19306 (N_19306,N_18847,N_18772);
nor U19307 (N_19307,N_18644,N_18671);
nor U19308 (N_19308,N_18831,N_19155);
nand U19309 (N_19309,N_18966,N_18915);
xnor U19310 (N_19310,N_18669,N_19078);
xor U19311 (N_19311,N_18804,N_18933);
nor U19312 (N_19312,N_18895,N_19059);
xor U19313 (N_19313,N_18725,N_19054);
and U19314 (N_19314,N_18905,N_19148);
or U19315 (N_19315,N_18643,N_18742);
or U19316 (N_19316,N_18720,N_18913);
or U19317 (N_19317,N_18979,N_18783);
xnor U19318 (N_19318,N_19181,N_18792);
or U19319 (N_19319,N_19151,N_19165);
xnor U19320 (N_19320,N_18786,N_19012);
or U19321 (N_19321,N_18805,N_18670);
xnor U19322 (N_19322,N_19120,N_18938);
and U19323 (N_19323,N_18603,N_18765);
and U19324 (N_19324,N_19169,N_19117);
or U19325 (N_19325,N_18733,N_18877);
or U19326 (N_19326,N_18853,N_19002);
nand U19327 (N_19327,N_19045,N_19007);
xor U19328 (N_19328,N_19013,N_18791);
nor U19329 (N_19329,N_19070,N_19055);
and U19330 (N_19330,N_18897,N_19038);
or U19331 (N_19331,N_19145,N_18634);
or U19332 (N_19332,N_18828,N_18689);
xor U19333 (N_19333,N_19150,N_18717);
nand U19334 (N_19334,N_18958,N_18989);
nand U19335 (N_19335,N_19023,N_19039);
xor U19336 (N_19336,N_19110,N_18956);
xor U19337 (N_19337,N_18727,N_18884);
xnor U19338 (N_19338,N_18960,N_18612);
nand U19339 (N_19339,N_18868,N_18906);
nor U19340 (N_19340,N_18665,N_18909);
xor U19341 (N_19341,N_18842,N_18711);
nand U19342 (N_19342,N_19049,N_18739);
xnor U19343 (N_19343,N_18760,N_18706);
nand U19344 (N_19344,N_18655,N_18764);
xnor U19345 (N_19345,N_18770,N_18622);
and U19346 (N_19346,N_18787,N_18757);
and U19347 (N_19347,N_18984,N_19061);
and U19348 (N_19348,N_18978,N_18635);
nand U19349 (N_19349,N_18809,N_18625);
nand U19350 (N_19350,N_18992,N_19192);
nor U19351 (N_19351,N_19171,N_18708);
xor U19352 (N_19352,N_18730,N_19075);
nand U19353 (N_19353,N_19015,N_18657);
xnor U19354 (N_19354,N_19149,N_18690);
nand U19355 (N_19355,N_18875,N_19069);
and U19356 (N_19356,N_18756,N_19194);
xor U19357 (N_19357,N_19027,N_19077);
or U19358 (N_19358,N_19174,N_18777);
or U19359 (N_19359,N_18951,N_18797);
xnor U19360 (N_19360,N_18789,N_18701);
and U19361 (N_19361,N_18688,N_19103);
and U19362 (N_19362,N_19163,N_19000);
or U19363 (N_19363,N_19093,N_18822);
and U19364 (N_19364,N_18824,N_18843);
and U19365 (N_19365,N_19176,N_18825);
and U19366 (N_19366,N_18962,N_19020);
and U19367 (N_19367,N_19188,N_18969);
or U19368 (N_19368,N_19016,N_18957);
nand U19369 (N_19369,N_18778,N_18965);
nor U19370 (N_19370,N_18638,N_18851);
or U19371 (N_19371,N_19017,N_18949);
nand U19372 (N_19372,N_18737,N_18808);
nand U19373 (N_19373,N_19011,N_19033);
and U19374 (N_19374,N_18681,N_18852);
xor U19375 (N_19375,N_18894,N_19108);
xor U19376 (N_19376,N_18934,N_18886);
and U19377 (N_19377,N_18646,N_19067);
nand U19378 (N_19378,N_18700,N_18709);
nor U19379 (N_19379,N_19121,N_18664);
nor U19380 (N_19380,N_18907,N_18658);
or U19381 (N_19381,N_18914,N_18614);
xor U19382 (N_19382,N_18997,N_19177);
or U19383 (N_19383,N_18813,N_19198);
and U19384 (N_19384,N_19136,N_18925);
or U19385 (N_19385,N_18721,N_18867);
or U19386 (N_19386,N_18672,N_18845);
nand U19387 (N_19387,N_18916,N_18980);
or U19388 (N_19388,N_18893,N_19126);
nor U19389 (N_19389,N_19092,N_18759);
xor U19390 (N_19390,N_19073,N_18838);
and U19391 (N_19391,N_18977,N_19006);
nand U19392 (N_19392,N_18740,N_18704);
nor U19393 (N_19393,N_18858,N_18988);
or U19394 (N_19394,N_18935,N_18950);
xor U19395 (N_19395,N_18762,N_19197);
xnor U19396 (N_19396,N_19129,N_18832);
nand U19397 (N_19397,N_18628,N_18692);
nand U19398 (N_19398,N_18801,N_19064);
nor U19399 (N_19399,N_18631,N_18835);
xnor U19400 (N_19400,N_18952,N_18814);
or U19401 (N_19401,N_18863,N_19074);
nand U19402 (N_19402,N_18713,N_19087);
xor U19403 (N_19403,N_19018,N_18623);
xor U19404 (N_19404,N_18846,N_18610);
xor U19405 (N_19405,N_18864,N_18754);
nand U19406 (N_19406,N_19004,N_18946);
nor U19407 (N_19407,N_18889,N_19170);
or U19408 (N_19408,N_18639,N_18602);
xor U19409 (N_19409,N_18683,N_19058);
or U19410 (N_19410,N_18994,N_19082);
xor U19411 (N_19411,N_18922,N_18993);
or U19412 (N_19412,N_19166,N_18647);
nor U19413 (N_19413,N_19014,N_18738);
xor U19414 (N_19414,N_18736,N_18929);
or U19415 (N_19415,N_19037,N_19080);
and U19416 (N_19416,N_19138,N_18699);
nor U19417 (N_19417,N_18758,N_18974);
and U19418 (N_19418,N_18803,N_19010);
and U19419 (N_19419,N_19186,N_18971);
xor U19420 (N_19420,N_18662,N_18653);
nand U19421 (N_19421,N_18645,N_18947);
xor U19422 (N_19422,N_19109,N_19147);
nand U19423 (N_19423,N_19005,N_18749);
and U19424 (N_19424,N_18821,N_19167);
or U19425 (N_19425,N_19119,N_19112);
nor U19426 (N_19426,N_18917,N_18775);
and U19427 (N_19427,N_19056,N_18849);
or U19428 (N_19428,N_18800,N_18881);
nor U19429 (N_19429,N_19185,N_18931);
xnor U19430 (N_19430,N_18890,N_18697);
nor U19431 (N_19431,N_18942,N_18660);
or U19432 (N_19432,N_18773,N_19044);
xnor U19433 (N_19433,N_18983,N_18636);
nand U19434 (N_19434,N_18795,N_18632);
and U19435 (N_19435,N_18880,N_19071);
nor U19436 (N_19436,N_19095,N_18613);
nor U19437 (N_19437,N_18976,N_18919);
nand U19438 (N_19438,N_18750,N_19116);
and U19439 (N_19439,N_18668,N_19124);
or U19440 (N_19440,N_19115,N_18920);
nor U19441 (N_19441,N_18862,N_18991);
xor U19442 (N_19442,N_19101,N_19158);
and U19443 (N_19443,N_18741,N_18641);
nor U19444 (N_19444,N_19127,N_18961);
xor U19445 (N_19445,N_18600,N_18857);
xor U19446 (N_19446,N_19152,N_18624);
or U19447 (N_19447,N_19131,N_18780);
xor U19448 (N_19448,N_18948,N_18859);
and U19449 (N_19449,N_18963,N_19030);
nand U19450 (N_19450,N_18611,N_19050);
and U19451 (N_19451,N_18869,N_18642);
nand U19452 (N_19452,N_19111,N_18910);
or U19453 (N_19453,N_18899,N_18903);
or U19454 (N_19454,N_18854,N_18774);
and U19455 (N_19455,N_18836,N_18817);
nor U19456 (N_19456,N_18652,N_18972);
nand U19457 (N_19457,N_18691,N_19191);
nor U19458 (N_19458,N_19079,N_19098);
or U19459 (N_19459,N_18932,N_18860);
xnor U19460 (N_19460,N_18605,N_18887);
xnor U19461 (N_19461,N_18676,N_18607);
or U19462 (N_19462,N_19086,N_19009);
or U19463 (N_19463,N_18661,N_19153);
and U19464 (N_19464,N_19041,N_19107);
nor U19465 (N_19465,N_19104,N_18648);
nor U19466 (N_19466,N_18608,N_18937);
nand U19467 (N_19467,N_18769,N_18839);
xor U19468 (N_19468,N_19134,N_18799);
nor U19469 (N_19469,N_19036,N_18618);
nand U19470 (N_19470,N_18685,N_19113);
nor U19471 (N_19471,N_19161,N_18782);
nand U19472 (N_19472,N_19190,N_19047);
xor U19473 (N_19473,N_18619,N_18785);
nand U19474 (N_19474,N_19088,N_18898);
nor U19475 (N_19475,N_18818,N_18788);
xnor U19476 (N_19476,N_19187,N_18677);
xnor U19477 (N_19477,N_18746,N_18912);
nor U19478 (N_19478,N_18751,N_18986);
xor U19479 (N_19479,N_18714,N_19052);
nand U19480 (N_19480,N_18879,N_18793);
nand U19481 (N_19481,N_18923,N_18682);
and U19482 (N_19482,N_19183,N_19137);
and U19483 (N_19483,N_18719,N_18695);
nand U19484 (N_19484,N_19062,N_18941);
xor U19485 (N_19485,N_18982,N_18790);
or U19486 (N_19486,N_18970,N_18964);
nor U19487 (N_19487,N_19051,N_19142);
and U19488 (N_19488,N_19022,N_19162);
and U19489 (N_19489,N_18820,N_19081);
nand U19490 (N_19490,N_18834,N_18679);
or U19491 (N_19491,N_19140,N_19125);
nor U19492 (N_19492,N_18861,N_18872);
xnor U19493 (N_19493,N_18606,N_18686);
and U19494 (N_19494,N_18743,N_18996);
nor U19495 (N_19495,N_18707,N_18693);
or U19496 (N_19496,N_18953,N_19106);
nand U19497 (N_19497,N_19042,N_19083);
and U19498 (N_19498,N_19180,N_18698);
and U19499 (N_19499,N_18848,N_19029);
nor U19500 (N_19500,N_19057,N_18717);
xnor U19501 (N_19501,N_18987,N_18619);
nor U19502 (N_19502,N_18864,N_19060);
and U19503 (N_19503,N_18924,N_18651);
xor U19504 (N_19504,N_18871,N_19161);
or U19505 (N_19505,N_18732,N_18673);
nand U19506 (N_19506,N_18701,N_19029);
xor U19507 (N_19507,N_18667,N_18813);
and U19508 (N_19508,N_18770,N_18955);
or U19509 (N_19509,N_18763,N_19153);
and U19510 (N_19510,N_18964,N_18805);
nand U19511 (N_19511,N_19100,N_18696);
and U19512 (N_19512,N_19097,N_19058);
nand U19513 (N_19513,N_19114,N_18822);
xnor U19514 (N_19514,N_19005,N_18844);
nand U19515 (N_19515,N_18743,N_19157);
nor U19516 (N_19516,N_19146,N_18622);
and U19517 (N_19517,N_18926,N_18707);
or U19518 (N_19518,N_18617,N_19151);
and U19519 (N_19519,N_19183,N_18957);
nand U19520 (N_19520,N_18886,N_18708);
nor U19521 (N_19521,N_18856,N_18893);
xor U19522 (N_19522,N_19116,N_18663);
and U19523 (N_19523,N_18983,N_19186);
and U19524 (N_19524,N_18740,N_19117);
or U19525 (N_19525,N_18766,N_18629);
nor U19526 (N_19526,N_18658,N_18613);
nand U19527 (N_19527,N_18635,N_18910);
nand U19528 (N_19528,N_18830,N_19042);
and U19529 (N_19529,N_18739,N_18712);
xnor U19530 (N_19530,N_18744,N_19191);
or U19531 (N_19531,N_18785,N_18969);
nand U19532 (N_19532,N_19040,N_19037);
or U19533 (N_19533,N_18791,N_18806);
xnor U19534 (N_19534,N_18684,N_19105);
xnor U19535 (N_19535,N_18774,N_19171);
xnor U19536 (N_19536,N_18876,N_19092);
nor U19537 (N_19537,N_18736,N_19116);
and U19538 (N_19538,N_18933,N_18825);
nor U19539 (N_19539,N_18787,N_19076);
nor U19540 (N_19540,N_19032,N_18735);
and U19541 (N_19541,N_18704,N_19005);
nor U19542 (N_19542,N_18821,N_18912);
or U19543 (N_19543,N_18727,N_18828);
or U19544 (N_19544,N_18702,N_19191);
xnor U19545 (N_19545,N_19060,N_19102);
nor U19546 (N_19546,N_18877,N_18893);
xor U19547 (N_19547,N_18780,N_19195);
or U19548 (N_19548,N_18822,N_18670);
and U19549 (N_19549,N_18742,N_19072);
and U19550 (N_19550,N_18762,N_19116);
and U19551 (N_19551,N_18603,N_18655);
nand U19552 (N_19552,N_18632,N_18944);
or U19553 (N_19553,N_18984,N_19069);
or U19554 (N_19554,N_18614,N_19110);
nand U19555 (N_19555,N_18614,N_18849);
xor U19556 (N_19556,N_18617,N_18779);
and U19557 (N_19557,N_19199,N_19187);
xnor U19558 (N_19558,N_18713,N_18948);
nand U19559 (N_19559,N_18837,N_18737);
nand U19560 (N_19560,N_18866,N_18628);
or U19561 (N_19561,N_18694,N_18816);
or U19562 (N_19562,N_19046,N_18812);
nand U19563 (N_19563,N_19194,N_18759);
nand U19564 (N_19564,N_18832,N_19144);
nand U19565 (N_19565,N_18724,N_18995);
xnor U19566 (N_19566,N_19173,N_18762);
or U19567 (N_19567,N_18637,N_19193);
and U19568 (N_19568,N_19013,N_18786);
xor U19569 (N_19569,N_18890,N_18629);
xor U19570 (N_19570,N_19049,N_18623);
nand U19571 (N_19571,N_19052,N_18662);
xnor U19572 (N_19572,N_19076,N_18829);
nand U19573 (N_19573,N_18929,N_18621);
and U19574 (N_19574,N_19171,N_18677);
and U19575 (N_19575,N_18917,N_18808);
nand U19576 (N_19576,N_18774,N_18813);
xor U19577 (N_19577,N_18947,N_18881);
and U19578 (N_19578,N_18614,N_19120);
nor U19579 (N_19579,N_18809,N_19049);
nor U19580 (N_19580,N_19137,N_18709);
nor U19581 (N_19581,N_19145,N_18814);
xor U19582 (N_19582,N_18910,N_18712);
or U19583 (N_19583,N_18645,N_18888);
nand U19584 (N_19584,N_18743,N_18749);
or U19585 (N_19585,N_18857,N_18604);
and U19586 (N_19586,N_19110,N_19168);
nor U19587 (N_19587,N_18890,N_18901);
nand U19588 (N_19588,N_18855,N_18898);
nand U19589 (N_19589,N_18659,N_18691);
nand U19590 (N_19590,N_18655,N_18633);
or U19591 (N_19591,N_18814,N_18883);
nand U19592 (N_19592,N_18795,N_18851);
nor U19593 (N_19593,N_19191,N_19141);
or U19594 (N_19594,N_19173,N_18776);
nand U19595 (N_19595,N_19195,N_18603);
xor U19596 (N_19596,N_19114,N_19060);
xor U19597 (N_19597,N_18665,N_18804);
or U19598 (N_19598,N_19064,N_18726);
or U19599 (N_19599,N_19095,N_19035);
and U19600 (N_19600,N_18922,N_18775);
xnor U19601 (N_19601,N_19144,N_18924);
or U19602 (N_19602,N_19068,N_18907);
nor U19603 (N_19603,N_18606,N_18829);
and U19604 (N_19604,N_18628,N_19010);
or U19605 (N_19605,N_19004,N_18639);
nor U19606 (N_19606,N_18994,N_18795);
nor U19607 (N_19607,N_18824,N_18642);
and U19608 (N_19608,N_18987,N_18676);
xor U19609 (N_19609,N_18961,N_18764);
nand U19610 (N_19610,N_19003,N_18969);
nand U19611 (N_19611,N_18774,N_18684);
or U19612 (N_19612,N_18876,N_18783);
xor U19613 (N_19613,N_18834,N_19095);
nor U19614 (N_19614,N_18824,N_18809);
nand U19615 (N_19615,N_19084,N_18902);
nor U19616 (N_19616,N_18761,N_18949);
nand U19617 (N_19617,N_19111,N_19018);
and U19618 (N_19618,N_18962,N_19057);
and U19619 (N_19619,N_18927,N_18779);
nor U19620 (N_19620,N_18663,N_18677);
and U19621 (N_19621,N_19042,N_18793);
nand U19622 (N_19622,N_18871,N_19032);
nand U19623 (N_19623,N_19117,N_18927);
and U19624 (N_19624,N_19107,N_18847);
or U19625 (N_19625,N_18652,N_18844);
or U19626 (N_19626,N_19089,N_19068);
xor U19627 (N_19627,N_18888,N_18756);
nand U19628 (N_19628,N_18607,N_19017);
and U19629 (N_19629,N_18935,N_18692);
nor U19630 (N_19630,N_18634,N_18903);
nor U19631 (N_19631,N_18952,N_18821);
or U19632 (N_19632,N_18658,N_18727);
and U19633 (N_19633,N_18721,N_18763);
nand U19634 (N_19634,N_19126,N_19064);
and U19635 (N_19635,N_18743,N_18938);
or U19636 (N_19636,N_18782,N_18868);
or U19637 (N_19637,N_18735,N_19099);
nand U19638 (N_19638,N_18685,N_19080);
and U19639 (N_19639,N_18812,N_18796);
and U19640 (N_19640,N_18792,N_18742);
xnor U19641 (N_19641,N_19118,N_18958);
xnor U19642 (N_19642,N_18832,N_18688);
or U19643 (N_19643,N_19071,N_18708);
or U19644 (N_19644,N_19186,N_18780);
xor U19645 (N_19645,N_19119,N_18943);
and U19646 (N_19646,N_19107,N_18907);
nand U19647 (N_19647,N_18822,N_18707);
or U19648 (N_19648,N_18800,N_18921);
nor U19649 (N_19649,N_18903,N_18883);
xnor U19650 (N_19650,N_19034,N_18622);
xnor U19651 (N_19651,N_18903,N_18887);
nor U19652 (N_19652,N_18663,N_18820);
and U19653 (N_19653,N_18930,N_18770);
nor U19654 (N_19654,N_18889,N_19006);
nor U19655 (N_19655,N_19188,N_19050);
nor U19656 (N_19656,N_18852,N_19029);
or U19657 (N_19657,N_19142,N_18811);
nand U19658 (N_19658,N_18832,N_18920);
xnor U19659 (N_19659,N_18896,N_18978);
nor U19660 (N_19660,N_18917,N_18902);
or U19661 (N_19661,N_18672,N_18982);
nor U19662 (N_19662,N_18879,N_18893);
or U19663 (N_19663,N_18826,N_18660);
xnor U19664 (N_19664,N_18604,N_18897);
nand U19665 (N_19665,N_18658,N_18947);
xor U19666 (N_19666,N_19147,N_18958);
xor U19667 (N_19667,N_19066,N_18870);
nor U19668 (N_19668,N_18893,N_19006);
or U19669 (N_19669,N_18781,N_19081);
nand U19670 (N_19670,N_19020,N_19048);
and U19671 (N_19671,N_19095,N_18841);
or U19672 (N_19672,N_18672,N_18963);
nand U19673 (N_19673,N_19148,N_19010);
nand U19674 (N_19674,N_19123,N_18825);
or U19675 (N_19675,N_18974,N_18769);
xor U19676 (N_19676,N_18954,N_19165);
nor U19677 (N_19677,N_18976,N_18729);
xor U19678 (N_19678,N_18822,N_18923);
nand U19679 (N_19679,N_18897,N_19119);
and U19680 (N_19680,N_18826,N_19158);
nor U19681 (N_19681,N_19063,N_18652);
xor U19682 (N_19682,N_18770,N_19197);
xnor U19683 (N_19683,N_18915,N_18611);
nor U19684 (N_19684,N_18845,N_18976);
nand U19685 (N_19685,N_19143,N_19036);
or U19686 (N_19686,N_19051,N_18680);
and U19687 (N_19687,N_18822,N_18603);
nand U19688 (N_19688,N_18859,N_18937);
and U19689 (N_19689,N_19008,N_18708);
nor U19690 (N_19690,N_18909,N_18671);
or U19691 (N_19691,N_19187,N_19072);
and U19692 (N_19692,N_18822,N_18998);
or U19693 (N_19693,N_18675,N_18758);
nand U19694 (N_19694,N_18778,N_18737);
and U19695 (N_19695,N_19076,N_19171);
or U19696 (N_19696,N_18855,N_18610);
nand U19697 (N_19697,N_18679,N_19188);
nand U19698 (N_19698,N_19142,N_19064);
or U19699 (N_19699,N_18706,N_18680);
nor U19700 (N_19700,N_19032,N_18745);
nand U19701 (N_19701,N_18622,N_18965);
and U19702 (N_19702,N_18843,N_18771);
xnor U19703 (N_19703,N_18758,N_18822);
and U19704 (N_19704,N_19070,N_18633);
nor U19705 (N_19705,N_18724,N_18636);
or U19706 (N_19706,N_18910,N_18678);
or U19707 (N_19707,N_18988,N_19059);
xor U19708 (N_19708,N_18695,N_18782);
nor U19709 (N_19709,N_19038,N_19165);
nand U19710 (N_19710,N_19175,N_18931);
and U19711 (N_19711,N_18790,N_18903);
xnor U19712 (N_19712,N_18667,N_19175);
nor U19713 (N_19713,N_18696,N_18653);
and U19714 (N_19714,N_19090,N_18747);
nor U19715 (N_19715,N_18936,N_18825);
or U19716 (N_19716,N_18768,N_19038);
xor U19717 (N_19717,N_18856,N_18630);
nand U19718 (N_19718,N_19047,N_19169);
nor U19719 (N_19719,N_18965,N_18937);
nand U19720 (N_19720,N_18821,N_18625);
or U19721 (N_19721,N_18958,N_18614);
nor U19722 (N_19722,N_18700,N_19107);
nor U19723 (N_19723,N_19035,N_19041);
and U19724 (N_19724,N_18762,N_18926);
or U19725 (N_19725,N_18854,N_18984);
xnor U19726 (N_19726,N_18861,N_19051);
nor U19727 (N_19727,N_19140,N_18744);
or U19728 (N_19728,N_19018,N_18984);
nand U19729 (N_19729,N_18854,N_18970);
nand U19730 (N_19730,N_18829,N_18643);
nand U19731 (N_19731,N_18762,N_18664);
or U19732 (N_19732,N_18812,N_19083);
nand U19733 (N_19733,N_18957,N_19087);
nor U19734 (N_19734,N_18665,N_19073);
xnor U19735 (N_19735,N_19177,N_18703);
nor U19736 (N_19736,N_18744,N_18608);
xnor U19737 (N_19737,N_18991,N_18699);
nand U19738 (N_19738,N_19020,N_18891);
and U19739 (N_19739,N_18767,N_18836);
xnor U19740 (N_19740,N_18968,N_19160);
nand U19741 (N_19741,N_18831,N_19126);
and U19742 (N_19742,N_19107,N_18934);
nor U19743 (N_19743,N_18681,N_19129);
and U19744 (N_19744,N_18881,N_18811);
nand U19745 (N_19745,N_18683,N_19013);
and U19746 (N_19746,N_18756,N_19037);
xor U19747 (N_19747,N_19047,N_18954);
nand U19748 (N_19748,N_18616,N_18752);
nor U19749 (N_19749,N_19036,N_18692);
nor U19750 (N_19750,N_19128,N_18886);
or U19751 (N_19751,N_18909,N_19164);
and U19752 (N_19752,N_19111,N_18987);
xnor U19753 (N_19753,N_18812,N_19143);
nand U19754 (N_19754,N_18643,N_18686);
and U19755 (N_19755,N_19069,N_18753);
and U19756 (N_19756,N_18897,N_18912);
nor U19757 (N_19757,N_18833,N_18819);
or U19758 (N_19758,N_18900,N_18880);
nor U19759 (N_19759,N_18877,N_19116);
and U19760 (N_19760,N_19051,N_19062);
nor U19761 (N_19761,N_18851,N_18668);
nand U19762 (N_19762,N_18673,N_18639);
xor U19763 (N_19763,N_19124,N_18727);
and U19764 (N_19764,N_18695,N_18898);
nand U19765 (N_19765,N_19162,N_18831);
xnor U19766 (N_19766,N_18783,N_19177);
and U19767 (N_19767,N_18786,N_18752);
and U19768 (N_19768,N_18664,N_19186);
and U19769 (N_19769,N_18954,N_18651);
or U19770 (N_19770,N_18761,N_19093);
xnor U19771 (N_19771,N_18709,N_18795);
and U19772 (N_19772,N_18816,N_19156);
nand U19773 (N_19773,N_18924,N_18831);
and U19774 (N_19774,N_18828,N_18807);
xor U19775 (N_19775,N_18793,N_19068);
or U19776 (N_19776,N_18877,N_18847);
nor U19777 (N_19777,N_18902,N_18903);
or U19778 (N_19778,N_18660,N_19022);
or U19779 (N_19779,N_18771,N_18793);
and U19780 (N_19780,N_18761,N_18960);
nand U19781 (N_19781,N_18991,N_18743);
xnor U19782 (N_19782,N_18926,N_19052);
and U19783 (N_19783,N_18666,N_19054);
or U19784 (N_19784,N_19096,N_18885);
xor U19785 (N_19785,N_18607,N_18923);
nor U19786 (N_19786,N_19004,N_18625);
nor U19787 (N_19787,N_18740,N_18936);
xor U19788 (N_19788,N_19055,N_18832);
nand U19789 (N_19789,N_19158,N_19083);
and U19790 (N_19790,N_18672,N_18833);
or U19791 (N_19791,N_19145,N_19149);
or U19792 (N_19792,N_18913,N_19195);
nand U19793 (N_19793,N_18710,N_18999);
or U19794 (N_19794,N_19080,N_19164);
and U19795 (N_19795,N_18711,N_18819);
xnor U19796 (N_19796,N_19109,N_19080);
xnor U19797 (N_19797,N_19117,N_19097);
nand U19798 (N_19798,N_18660,N_18945);
nor U19799 (N_19799,N_18766,N_18676);
nor U19800 (N_19800,N_19440,N_19705);
or U19801 (N_19801,N_19637,N_19731);
nand U19802 (N_19802,N_19538,N_19508);
nor U19803 (N_19803,N_19535,N_19729);
or U19804 (N_19804,N_19706,N_19693);
or U19805 (N_19805,N_19794,N_19524);
nor U19806 (N_19806,N_19733,N_19695);
or U19807 (N_19807,N_19320,N_19501);
xor U19808 (N_19808,N_19607,N_19278);
and U19809 (N_19809,N_19398,N_19448);
nor U19810 (N_19810,N_19276,N_19312);
nor U19811 (N_19811,N_19658,N_19240);
xor U19812 (N_19812,N_19670,N_19404);
xnor U19813 (N_19813,N_19460,N_19313);
xnor U19814 (N_19814,N_19761,N_19392);
nor U19815 (N_19815,N_19441,N_19283);
nor U19816 (N_19816,N_19744,N_19742);
nand U19817 (N_19817,N_19598,N_19597);
nand U19818 (N_19818,N_19580,N_19261);
xor U19819 (N_19819,N_19436,N_19287);
and U19820 (N_19820,N_19771,N_19371);
nor U19821 (N_19821,N_19447,N_19410);
nand U19822 (N_19822,N_19792,N_19745);
nor U19823 (N_19823,N_19568,N_19424);
nand U19824 (N_19824,N_19730,N_19358);
and U19825 (N_19825,N_19395,N_19725);
nand U19826 (N_19826,N_19323,N_19207);
and U19827 (N_19827,N_19361,N_19333);
or U19828 (N_19828,N_19582,N_19243);
xnor U19829 (N_19829,N_19482,N_19717);
and U19830 (N_19830,N_19306,N_19563);
nand U19831 (N_19831,N_19595,N_19336);
nand U19832 (N_19832,N_19768,N_19633);
nand U19833 (N_19833,N_19709,N_19663);
xor U19834 (N_19834,N_19669,N_19684);
or U19835 (N_19835,N_19774,N_19626);
nor U19836 (N_19836,N_19406,N_19746);
xor U19837 (N_19837,N_19701,N_19710);
and U19838 (N_19838,N_19239,N_19542);
and U19839 (N_19839,N_19412,N_19530);
or U19840 (N_19840,N_19788,N_19541);
and U19841 (N_19841,N_19326,N_19564);
xor U19842 (N_19842,N_19376,N_19439);
and U19843 (N_19843,N_19485,N_19660);
or U19844 (N_19844,N_19233,N_19795);
nand U19845 (N_19845,N_19522,N_19429);
or U19846 (N_19846,N_19609,N_19783);
or U19847 (N_19847,N_19519,N_19483);
and U19848 (N_19848,N_19380,N_19790);
nand U19849 (N_19849,N_19355,N_19246);
or U19850 (N_19850,N_19791,N_19735);
nand U19851 (N_19851,N_19211,N_19578);
and U19852 (N_19852,N_19282,N_19570);
nor U19853 (N_19853,N_19286,N_19652);
nand U19854 (N_19854,N_19421,N_19699);
nor U19855 (N_19855,N_19712,N_19471);
or U19856 (N_19856,N_19533,N_19462);
nand U19857 (N_19857,N_19648,N_19591);
xor U19858 (N_19858,N_19388,N_19691);
or U19859 (N_19859,N_19290,N_19571);
or U19860 (N_19860,N_19399,N_19437);
or U19861 (N_19861,N_19645,N_19346);
and U19862 (N_19862,N_19719,N_19270);
xor U19863 (N_19863,N_19650,N_19269);
or U19864 (N_19864,N_19664,N_19377);
and U19865 (N_19865,N_19277,N_19428);
nand U19866 (N_19866,N_19451,N_19770);
xnor U19867 (N_19867,N_19704,N_19433);
xnor U19868 (N_19868,N_19367,N_19305);
nor U19869 (N_19869,N_19734,N_19552);
nor U19870 (N_19870,N_19469,N_19720);
xnor U19871 (N_19871,N_19726,N_19521);
nand U19872 (N_19872,N_19452,N_19702);
or U19873 (N_19873,N_19752,N_19241);
or U19874 (N_19874,N_19213,N_19772);
nand U19875 (N_19875,N_19206,N_19222);
and U19876 (N_19876,N_19723,N_19671);
or U19877 (N_19877,N_19784,N_19294);
nor U19878 (N_19878,N_19724,N_19321);
nand U19879 (N_19879,N_19610,N_19453);
or U19880 (N_19880,N_19430,N_19472);
or U19881 (N_19881,N_19438,N_19748);
or U19882 (N_19882,N_19778,N_19318);
nor U19883 (N_19883,N_19267,N_19235);
and U19884 (N_19884,N_19255,N_19740);
nor U19885 (N_19885,N_19590,N_19688);
nand U19886 (N_19886,N_19348,N_19750);
and U19887 (N_19887,N_19621,N_19511);
or U19888 (N_19888,N_19515,N_19225);
or U19889 (N_19889,N_19315,N_19692);
nand U19890 (N_19890,N_19549,N_19588);
nor U19891 (N_19891,N_19343,N_19491);
nor U19892 (N_19892,N_19666,N_19608);
or U19893 (N_19893,N_19427,N_19565);
or U19894 (N_19894,N_19350,N_19529);
and U19895 (N_19895,N_19423,N_19727);
xor U19896 (N_19896,N_19411,N_19434);
nand U19897 (N_19897,N_19481,N_19581);
and U19898 (N_19898,N_19754,N_19363);
nand U19899 (N_19899,N_19518,N_19760);
nor U19900 (N_19900,N_19218,N_19732);
nand U19901 (N_19901,N_19219,N_19583);
nor U19902 (N_19902,N_19273,N_19776);
and U19903 (N_19903,N_19209,N_19554);
nand U19904 (N_19904,N_19536,N_19227);
xnor U19905 (N_19905,N_19299,N_19340);
or U19906 (N_19906,N_19574,N_19560);
nor U19907 (N_19907,N_19217,N_19496);
nor U19908 (N_19908,N_19722,N_19514);
and U19909 (N_19909,N_19532,N_19446);
nand U19910 (N_19910,N_19493,N_19548);
nand U19911 (N_19911,N_19203,N_19600);
nor U19912 (N_19912,N_19618,N_19668);
and U19913 (N_19913,N_19716,N_19512);
or U19914 (N_19914,N_19301,N_19259);
nor U19915 (N_19915,N_19527,N_19573);
nand U19916 (N_19916,N_19466,N_19444);
nor U19917 (N_19917,N_19615,N_19516);
and U19918 (N_19918,N_19293,N_19289);
nor U19919 (N_19919,N_19201,N_19576);
xor U19920 (N_19920,N_19679,N_19526);
xnor U19921 (N_19921,N_19338,N_19486);
xor U19922 (N_19922,N_19628,N_19537);
and U19923 (N_19923,N_19539,N_19417);
or U19924 (N_19924,N_19409,N_19463);
xor U19925 (N_19925,N_19480,N_19585);
xor U19926 (N_19926,N_19556,N_19540);
xnor U19927 (N_19927,N_19632,N_19718);
xor U19928 (N_19928,N_19685,N_19374);
and U19929 (N_19929,N_19640,N_19579);
nand U19930 (N_19930,N_19762,N_19384);
nand U19931 (N_19931,N_19620,N_19780);
nor U19932 (N_19932,N_19674,N_19407);
xor U19933 (N_19933,N_19260,N_19566);
xor U19934 (N_19934,N_19677,N_19789);
nor U19935 (N_19935,N_19248,N_19756);
nand U19936 (N_19936,N_19779,N_19476);
and U19937 (N_19937,N_19464,N_19465);
or U19938 (N_19938,N_19329,N_19455);
nor U19939 (N_19939,N_19349,N_19602);
or U19940 (N_19940,N_19767,N_19475);
xor U19941 (N_19941,N_19275,N_19359);
nor U19942 (N_19942,N_19711,N_19559);
or U19943 (N_19943,N_19528,N_19322);
nor U19944 (N_19944,N_19657,N_19319);
nor U19945 (N_19945,N_19506,N_19468);
nor U19946 (N_19946,N_19781,N_19456);
nand U19947 (N_19947,N_19467,N_19347);
nor U19948 (N_19948,N_19403,N_19584);
or U19949 (N_19949,N_19229,N_19419);
or U19950 (N_19950,N_19749,N_19297);
or U19951 (N_19951,N_19596,N_19341);
or U19952 (N_19952,N_19344,N_19517);
or U19953 (N_19953,N_19252,N_19787);
nor U19954 (N_19954,N_19694,N_19425);
nand U19955 (N_19955,N_19775,N_19263);
nand U19956 (N_19956,N_19234,N_19547);
or U19957 (N_19957,N_19703,N_19400);
or U19958 (N_19958,N_19531,N_19586);
or U19959 (N_19959,N_19414,N_19231);
nor U19960 (N_19960,N_19272,N_19649);
or U19961 (N_19961,N_19274,N_19328);
and U19962 (N_19962,N_19354,N_19310);
nor U19963 (N_19963,N_19226,N_19311);
nand U19964 (N_19964,N_19208,N_19629);
nand U19965 (N_19965,N_19280,N_19309);
xnor U19966 (N_19966,N_19708,N_19281);
or U19967 (N_19967,N_19592,N_19431);
and U19968 (N_19968,N_19606,N_19696);
nand U19969 (N_19969,N_19777,N_19636);
or U19970 (N_19970,N_19382,N_19545);
nand U19971 (N_19971,N_19498,N_19715);
and U19972 (N_19972,N_19351,N_19550);
and U19973 (N_19973,N_19655,N_19569);
nor U19974 (N_19974,N_19553,N_19622);
nor U19975 (N_19975,N_19449,N_19689);
and U19976 (N_19976,N_19534,N_19613);
or U19977 (N_19977,N_19551,N_19786);
and U19978 (N_19978,N_19461,N_19638);
nor U19979 (N_19979,N_19601,N_19249);
or U19980 (N_19980,N_19215,N_19646);
nand U19981 (N_19981,N_19676,N_19525);
or U19982 (N_19982,N_19793,N_19488);
xor U19983 (N_19983,N_19785,N_19639);
nor U19984 (N_19984,N_19230,N_19562);
nand U19985 (N_19985,N_19490,N_19221);
xnor U19986 (N_19986,N_19544,N_19303);
nor U19987 (N_19987,N_19594,N_19258);
or U19988 (N_19988,N_19375,N_19470);
nor U19989 (N_19989,N_19223,N_19237);
nor U19990 (N_19990,N_19751,N_19205);
and U19991 (N_19991,N_19330,N_19766);
and U19992 (N_19992,N_19391,N_19651);
nand U19993 (N_19993,N_19288,N_19339);
xor U19994 (N_19994,N_19625,N_19782);
nor U19995 (N_19995,N_19291,N_19279);
nor U19996 (N_19996,N_19271,N_19457);
and U19997 (N_19997,N_19383,N_19543);
xnor U19998 (N_19998,N_19707,N_19216);
nand U19999 (N_19999,N_19567,N_19523);
nor U20000 (N_20000,N_19678,N_19497);
xnor U20001 (N_20001,N_19763,N_19251);
nand U20002 (N_20002,N_19385,N_19690);
nand U20003 (N_20003,N_19499,N_19373);
or U20004 (N_20004,N_19416,N_19617);
nor U20005 (N_20005,N_19331,N_19262);
or U20006 (N_20006,N_19302,N_19370);
nor U20007 (N_20007,N_19558,N_19661);
nand U20008 (N_20008,N_19687,N_19682);
nand U20009 (N_20009,N_19324,N_19426);
and U20010 (N_20010,N_19212,N_19316);
xor U20011 (N_20011,N_19342,N_19555);
xor U20012 (N_20012,N_19224,N_19300);
nand U20013 (N_20013,N_19603,N_19799);
xor U20014 (N_20014,N_19624,N_19623);
and U20015 (N_20015,N_19713,N_19673);
and U20016 (N_20016,N_19334,N_19378);
nand U20017 (N_20017,N_19292,N_19256);
or U20018 (N_20018,N_19681,N_19757);
nand U20019 (N_20019,N_19504,N_19200);
or U20020 (N_20020,N_19204,N_19728);
nor U20021 (N_20021,N_19502,N_19654);
nand U20022 (N_20022,N_19647,N_19477);
nand U20023 (N_20023,N_19394,N_19614);
nand U20024 (N_20024,N_19686,N_19220);
nor U20025 (N_20025,N_19397,N_19641);
xor U20026 (N_20026,N_19325,N_19415);
xor U20027 (N_20027,N_19500,N_19432);
xnor U20028 (N_20028,N_19459,N_19314);
nand U20029 (N_20029,N_19572,N_19360);
xnor U20030 (N_20030,N_19236,N_19662);
and U20031 (N_20031,N_19589,N_19435);
xnor U20032 (N_20032,N_19317,N_19492);
nor U20033 (N_20033,N_19386,N_19659);
or U20034 (N_20034,N_19736,N_19509);
nand U20035 (N_20035,N_19796,N_19285);
nor U20036 (N_20036,N_19495,N_19232);
nor U20037 (N_20037,N_19362,N_19422);
xnor U20038 (N_20038,N_19401,N_19345);
nor U20039 (N_20039,N_19253,N_19210);
nand U20040 (N_20040,N_19630,N_19616);
nand U20041 (N_20041,N_19266,N_19714);
xor U20042 (N_20042,N_19634,N_19372);
xor U20043 (N_20043,N_19764,N_19605);
and U20044 (N_20044,N_19721,N_19520);
and U20045 (N_20045,N_19228,N_19364);
nand U20046 (N_20046,N_19365,N_19238);
xor U20047 (N_20047,N_19379,N_19513);
nand U20048 (N_20048,N_19387,N_19769);
or U20049 (N_20049,N_19737,N_19214);
nor U20050 (N_20050,N_19631,N_19643);
and U20051 (N_20051,N_19680,N_19593);
and U20052 (N_20052,N_19254,N_19798);
nor U20053 (N_20053,N_19250,N_19575);
xnor U20054 (N_20054,N_19478,N_19561);
nand U20055 (N_20055,N_19454,N_19773);
or U20056 (N_20056,N_19408,N_19604);
or U20057 (N_20057,N_19507,N_19479);
and U20058 (N_20058,N_19741,N_19420);
or U20059 (N_20059,N_19443,N_19667);
and U20060 (N_20060,N_19368,N_19257);
xnor U20061 (N_20061,N_19284,N_19245);
xor U20062 (N_20062,N_19642,N_19332);
xnor U20063 (N_20063,N_19738,N_19473);
nand U20064 (N_20064,N_19577,N_19489);
nand U20065 (N_20065,N_19242,N_19697);
or U20066 (N_20066,N_19244,N_19653);
nand U20067 (N_20067,N_19335,N_19357);
or U20068 (N_20068,N_19510,N_19337);
xor U20069 (N_20069,N_19675,N_19619);
nor U20070 (N_20070,N_19202,N_19381);
or U20071 (N_20071,N_19612,N_19611);
xor U20072 (N_20072,N_19308,N_19296);
or U20073 (N_20073,N_19503,N_19672);
xnor U20074 (N_20074,N_19352,N_19418);
or U20075 (N_20075,N_19369,N_19494);
nand U20076 (N_20076,N_19758,N_19557);
nor U20077 (N_20077,N_19587,N_19304);
or U20078 (N_20078,N_19445,N_19759);
nand U20079 (N_20079,N_19405,N_19743);
nor U20080 (N_20080,N_19797,N_19644);
nor U20081 (N_20081,N_19264,N_19665);
and U20082 (N_20082,N_19487,N_19755);
nand U20083 (N_20083,N_19656,N_19484);
nand U20084 (N_20084,N_19295,N_19546);
and U20085 (N_20085,N_19627,N_19393);
nor U20086 (N_20086,N_19474,N_19683);
xor U20087 (N_20087,N_19635,N_19753);
xor U20088 (N_20088,N_19765,N_19700);
and U20089 (N_20089,N_19747,N_19413);
and U20090 (N_20090,N_19265,N_19327);
xor U20091 (N_20091,N_19458,N_19366);
nand U20092 (N_20092,N_19353,N_19390);
and U20093 (N_20093,N_19247,N_19505);
or U20094 (N_20094,N_19268,N_19698);
nand U20095 (N_20095,N_19739,N_19389);
and U20096 (N_20096,N_19298,N_19450);
or U20097 (N_20097,N_19402,N_19442);
and U20098 (N_20098,N_19396,N_19356);
and U20099 (N_20099,N_19307,N_19599);
or U20100 (N_20100,N_19387,N_19516);
nor U20101 (N_20101,N_19641,N_19745);
or U20102 (N_20102,N_19225,N_19675);
nand U20103 (N_20103,N_19560,N_19248);
nor U20104 (N_20104,N_19244,N_19607);
nor U20105 (N_20105,N_19702,N_19666);
or U20106 (N_20106,N_19210,N_19444);
and U20107 (N_20107,N_19391,N_19316);
xor U20108 (N_20108,N_19499,N_19522);
nand U20109 (N_20109,N_19635,N_19456);
and U20110 (N_20110,N_19655,N_19547);
nor U20111 (N_20111,N_19609,N_19219);
or U20112 (N_20112,N_19780,N_19200);
xnor U20113 (N_20113,N_19295,N_19501);
nand U20114 (N_20114,N_19505,N_19463);
nor U20115 (N_20115,N_19445,N_19341);
xnor U20116 (N_20116,N_19548,N_19610);
and U20117 (N_20117,N_19727,N_19674);
or U20118 (N_20118,N_19374,N_19796);
nor U20119 (N_20119,N_19212,N_19684);
and U20120 (N_20120,N_19745,N_19418);
and U20121 (N_20121,N_19226,N_19754);
xor U20122 (N_20122,N_19547,N_19636);
nor U20123 (N_20123,N_19369,N_19718);
nand U20124 (N_20124,N_19418,N_19559);
xor U20125 (N_20125,N_19644,N_19406);
or U20126 (N_20126,N_19640,N_19488);
xnor U20127 (N_20127,N_19377,N_19415);
xnor U20128 (N_20128,N_19564,N_19393);
or U20129 (N_20129,N_19585,N_19372);
xor U20130 (N_20130,N_19563,N_19750);
xor U20131 (N_20131,N_19436,N_19718);
nor U20132 (N_20132,N_19471,N_19524);
xor U20133 (N_20133,N_19707,N_19373);
or U20134 (N_20134,N_19316,N_19792);
xor U20135 (N_20135,N_19336,N_19276);
and U20136 (N_20136,N_19200,N_19628);
nor U20137 (N_20137,N_19243,N_19772);
nor U20138 (N_20138,N_19306,N_19429);
nand U20139 (N_20139,N_19297,N_19725);
xor U20140 (N_20140,N_19573,N_19656);
xnor U20141 (N_20141,N_19674,N_19369);
and U20142 (N_20142,N_19258,N_19310);
xor U20143 (N_20143,N_19212,N_19401);
xnor U20144 (N_20144,N_19694,N_19762);
and U20145 (N_20145,N_19769,N_19504);
nand U20146 (N_20146,N_19485,N_19478);
and U20147 (N_20147,N_19612,N_19691);
nor U20148 (N_20148,N_19279,N_19207);
nor U20149 (N_20149,N_19449,N_19242);
xor U20150 (N_20150,N_19281,N_19755);
or U20151 (N_20151,N_19342,N_19365);
xor U20152 (N_20152,N_19734,N_19601);
or U20153 (N_20153,N_19521,N_19506);
and U20154 (N_20154,N_19581,N_19680);
nor U20155 (N_20155,N_19210,N_19385);
nand U20156 (N_20156,N_19234,N_19339);
or U20157 (N_20157,N_19668,N_19705);
nor U20158 (N_20158,N_19680,N_19223);
xor U20159 (N_20159,N_19258,N_19251);
nor U20160 (N_20160,N_19306,N_19419);
nand U20161 (N_20161,N_19268,N_19637);
and U20162 (N_20162,N_19641,N_19455);
nor U20163 (N_20163,N_19763,N_19281);
xor U20164 (N_20164,N_19610,N_19351);
or U20165 (N_20165,N_19234,N_19657);
or U20166 (N_20166,N_19583,N_19653);
nand U20167 (N_20167,N_19663,N_19229);
and U20168 (N_20168,N_19466,N_19257);
and U20169 (N_20169,N_19305,N_19418);
xnor U20170 (N_20170,N_19461,N_19355);
nor U20171 (N_20171,N_19206,N_19646);
nand U20172 (N_20172,N_19587,N_19717);
nand U20173 (N_20173,N_19636,N_19651);
nor U20174 (N_20174,N_19423,N_19501);
nand U20175 (N_20175,N_19200,N_19321);
nor U20176 (N_20176,N_19786,N_19387);
xnor U20177 (N_20177,N_19767,N_19765);
or U20178 (N_20178,N_19251,N_19646);
nand U20179 (N_20179,N_19627,N_19341);
nand U20180 (N_20180,N_19325,N_19329);
nor U20181 (N_20181,N_19348,N_19284);
or U20182 (N_20182,N_19767,N_19580);
xnor U20183 (N_20183,N_19507,N_19367);
xor U20184 (N_20184,N_19586,N_19466);
nor U20185 (N_20185,N_19616,N_19538);
xnor U20186 (N_20186,N_19359,N_19646);
xnor U20187 (N_20187,N_19285,N_19367);
nor U20188 (N_20188,N_19374,N_19492);
or U20189 (N_20189,N_19253,N_19291);
nor U20190 (N_20190,N_19411,N_19681);
nand U20191 (N_20191,N_19776,N_19265);
nor U20192 (N_20192,N_19352,N_19760);
or U20193 (N_20193,N_19743,N_19616);
or U20194 (N_20194,N_19575,N_19702);
nand U20195 (N_20195,N_19563,N_19537);
or U20196 (N_20196,N_19250,N_19281);
or U20197 (N_20197,N_19546,N_19794);
xnor U20198 (N_20198,N_19374,N_19206);
nor U20199 (N_20199,N_19405,N_19625);
or U20200 (N_20200,N_19538,N_19230);
nand U20201 (N_20201,N_19317,N_19200);
xnor U20202 (N_20202,N_19233,N_19409);
nand U20203 (N_20203,N_19353,N_19424);
or U20204 (N_20204,N_19644,N_19688);
or U20205 (N_20205,N_19798,N_19580);
nand U20206 (N_20206,N_19432,N_19762);
xor U20207 (N_20207,N_19407,N_19505);
or U20208 (N_20208,N_19559,N_19596);
xnor U20209 (N_20209,N_19491,N_19340);
and U20210 (N_20210,N_19422,N_19654);
nand U20211 (N_20211,N_19308,N_19695);
nor U20212 (N_20212,N_19522,N_19479);
nand U20213 (N_20213,N_19526,N_19245);
and U20214 (N_20214,N_19756,N_19208);
or U20215 (N_20215,N_19399,N_19273);
or U20216 (N_20216,N_19643,N_19429);
or U20217 (N_20217,N_19320,N_19728);
and U20218 (N_20218,N_19504,N_19282);
and U20219 (N_20219,N_19263,N_19272);
nor U20220 (N_20220,N_19705,N_19670);
or U20221 (N_20221,N_19404,N_19504);
nor U20222 (N_20222,N_19614,N_19281);
nor U20223 (N_20223,N_19404,N_19436);
and U20224 (N_20224,N_19655,N_19402);
nand U20225 (N_20225,N_19692,N_19269);
xnor U20226 (N_20226,N_19441,N_19344);
nor U20227 (N_20227,N_19319,N_19602);
nand U20228 (N_20228,N_19437,N_19253);
or U20229 (N_20229,N_19690,N_19266);
and U20230 (N_20230,N_19322,N_19329);
or U20231 (N_20231,N_19752,N_19772);
or U20232 (N_20232,N_19580,N_19554);
nor U20233 (N_20233,N_19432,N_19522);
and U20234 (N_20234,N_19749,N_19656);
xnor U20235 (N_20235,N_19664,N_19321);
or U20236 (N_20236,N_19550,N_19670);
xor U20237 (N_20237,N_19277,N_19580);
nor U20238 (N_20238,N_19229,N_19642);
nor U20239 (N_20239,N_19333,N_19513);
and U20240 (N_20240,N_19738,N_19596);
and U20241 (N_20241,N_19296,N_19233);
nand U20242 (N_20242,N_19507,N_19506);
nand U20243 (N_20243,N_19653,N_19725);
or U20244 (N_20244,N_19443,N_19307);
xor U20245 (N_20245,N_19436,N_19426);
and U20246 (N_20246,N_19241,N_19343);
nor U20247 (N_20247,N_19329,N_19723);
xor U20248 (N_20248,N_19253,N_19652);
nor U20249 (N_20249,N_19414,N_19406);
xor U20250 (N_20250,N_19294,N_19551);
or U20251 (N_20251,N_19204,N_19300);
xnor U20252 (N_20252,N_19340,N_19592);
nor U20253 (N_20253,N_19608,N_19442);
nor U20254 (N_20254,N_19590,N_19684);
or U20255 (N_20255,N_19668,N_19600);
nand U20256 (N_20256,N_19544,N_19416);
or U20257 (N_20257,N_19765,N_19712);
or U20258 (N_20258,N_19279,N_19226);
and U20259 (N_20259,N_19691,N_19767);
nand U20260 (N_20260,N_19753,N_19639);
or U20261 (N_20261,N_19617,N_19507);
nand U20262 (N_20262,N_19694,N_19621);
and U20263 (N_20263,N_19423,N_19679);
xor U20264 (N_20264,N_19662,N_19717);
or U20265 (N_20265,N_19697,N_19526);
nor U20266 (N_20266,N_19624,N_19229);
nand U20267 (N_20267,N_19344,N_19618);
nor U20268 (N_20268,N_19201,N_19323);
nor U20269 (N_20269,N_19657,N_19765);
xor U20270 (N_20270,N_19401,N_19787);
or U20271 (N_20271,N_19347,N_19497);
xor U20272 (N_20272,N_19493,N_19305);
and U20273 (N_20273,N_19584,N_19684);
nand U20274 (N_20274,N_19450,N_19697);
or U20275 (N_20275,N_19468,N_19671);
xor U20276 (N_20276,N_19274,N_19309);
nor U20277 (N_20277,N_19428,N_19249);
and U20278 (N_20278,N_19518,N_19235);
nand U20279 (N_20279,N_19656,N_19718);
xnor U20280 (N_20280,N_19637,N_19422);
nor U20281 (N_20281,N_19773,N_19287);
xor U20282 (N_20282,N_19358,N_19673);
nand U20283 (N_20283,N_19597,N_19311);
nand U20284 (N_20284,N_19455,N_19611);
or U20285 (N_20285,N_19373,N_19410);
nor U20286 (N_20286,N_19205,N_19465);
or U20287 (N_20287,N_19477,N_19451);
xnor U20288 (N_20288,N_19308,N_19717);
xor U20289 (N_20289,N_19381,N_19703);
nor U20290 (N_20290,N_19331,N_19712);
and U20291 (N_20291,N_19275,N_19767);
or U20292 (N_20292,N_19740,N_19309);
nor U20293 (N_20293,N_19408,N_19555);
or U20294 (N_20294,N_19603,N_19417);
xor U20295 (N_20295,N_19633,N_19278);
nor U20296 (N_20296,N_19440,N_19265);
nand U20297 (N_20297,N_19664,N_19537);
and U20298 (N_20298,N_19764,N_19693);
nor U20299 (N_20299,N_19563,N_19746);
nor U20300 (N_20300,N_19728,N_19561);
and U20301 (N_20301,N_19556,N_19594);
xor U20302 (N_20302,N_19370,N_19402);
or U20303 (N_20303,N_19493,N_19683);
nand U20304 (N_20304,N_19237,N_19315);
xor U20305 (N_20305,N_19713,N_19662);
nor U20306 (N_20306,N_19523,N_19218);
and U20307 (N_20307,N_19443,N_19584);
or U20308 (N_20308,N_19517,N_19590);
or U20309 (N_20309,N_19411,N_19378);
or U20310 (N_20310,N_19496,N_19291);
nor U20311 (N_20311,N_19725,N_19254);
xnor U20312 (N_20312,N_19270,N_19668);
nand U20313 (N_20313,N_19436,N_19574);
and U20314 (N_20314,N_19780,N_19245);
or U20315 (N_20315,N_19393,N_19637);
nor U20316 (N_20316,N_19383,N_19421);
and U20317 (N_20317,N_19341,N_19427);
xor U20318 (N_20318,N_19742,N_19523);
nor U20319 (N_20319,N_19620,N_19506);
or U20320 (N_20320,N_19306,N_19534);
nand U20321 (N_20321,N_19490,N_19342);
or U20322 (N_20322,N_19689,N_19480);
nor U20323 (N_20323,N_19294,N_19799);
xnor U20324 (N_20324,N_19263,N_19258);
or U20325 (N_20325,N_19662,N_19711);
nand U20326 (N_20326,N_19247,N_19290);
and U20327 (N_20327,N_19774,N_19639);
or U20328 (N_20328,N_19730,N_19443);
nand U20329 (N_20329,N_19622,N_19430);
nor U20330 (N_20330,N_19584,N_19305);
xor U20331 (N_20331,N_19498,N_19215);
nand U20332 (N_20332,N_19329,N_19526);
nor U20333 (N_20333,N_19495,N_19478);
xnor U20334 (N_20334,N_19641,N_19212);
nor U20335 (N_20335,N_19603,N_19392);
nor U20336 (N_20336,N_19577,N_19749);
nand U20337 (N_20337,N_19229,N_19307);
xor U20338 (N_20338,N_19781,N_19425);
or U20339 (N_20339,N_19746,N_19653);
nor U20340 (N_20340,N_19596,N_19501);
nand U20341 (N_20341,N_19501,N_19492);
nand U20342 (N_20342,N_19215,N_19741);
nand U20343 (N_20343,N_19309,N_19458);
xor U20344 (N_20344,N_19357,N_19496);
and U20345 (N_20345,N_19594,N_19307);
or U20346 (N_20346,N_19653,N_19513);
and U20347 (N_20347,N_19752,N_19202);
xor U20348 (N_20348,N_19789,N_19563);
or U20349 (N_20349,N_19794,N_19221);
xor U20350 (N_20350,N_19643,N_19431);
and U20351 (N_20351,N_19396,N_19654);
and U20352 (N_20352,N_19449,N_19340);
nand U20353 (N_20353,N_19792,N_19532);
nand U20354 (N_20354,N_19573,N_19564);
nor U20355 (N_20355,N_19725,N_19256);
or U20356 (N_20356,N_19688,N_19559);
and U20357 (N_20357,N_19689,N_19355);
xnor U20358 (N_20358,N_19787,N_19243);
nor U20359 (N_20359,N_19440,N_19368);
xnor U20360 (N_20360,N_19732,N_19345);
or U20361 (N_20361,N_19795,N_19397);
nand U20362 (N_20362,N_19243,N_19321);
xnor U20363 (N_20363,N_19278,N_19417);
nand U20364 (N_20364,N_19712,N_19683);
and U20365 (N_20365,N_19664,N_19226);
nand U20366 (N_20366,N_19201,N_19406);
and U20367 (N_20367,N_19368,N_19263);
and U20368 (N_20368,N_19778,N_19289);
or U20369 (N_20369,N_19543,N_19261);
or U20370 (N_20370,N_19695,N_19484);
nor U20371 (N_20371,N_19377,N_19697);
and U20372 (N_20372,N_19396,N_19642);
xor U20373 (N_20373,N_19741,N_19452);
xnor U20374 (N_20374,N_19550,N_19349);
nand U20375 (N_20375,N_19712,N_19490);
xnor U20376 (N_20376,N_19492,N_19349);
and U20377 (N_20377,N_19299,N_19219);
and U20378 (N_20378,N_19588,N_19674);
xor U20379 (N_20379,N_19674,N_19281);
nor U20380 (N_20380,N_19266,N_19327);
nor U20381 (N_20381,N_19601,N_19248);
or U20382 (N_20382,N_19209,N_19777);
and U20383 (N_20383,N_19299,N_19327);
nand U20384 (N_20384,N_19211,N_19596);
xnor U20385 (N_20385,N_19241,N_19302);
xnor U20386 (N_20386,N_19307,N_19777);
nand U20387 (N_20387,N_19277,N_19367);
nand U20388 (N_20388,N_19392,N_19738);
or U20389 (N_20389,N_19232,N_19794);
nand U20390 (N_20390,N_19790,N_19507);
and U20391 (N_20391,N_19786,N_19542);
and U20392 (N_20392,N_19558,N_19240);
xnor U20393 (N_20393,N_19455,N_19499);
nand U20394 (N_20394,N_19756,N_19284);
nand U20395 (N_20395,N_19670,N_19406);
nand U20396 (N_20396,N_19351,N_19436);
nor U20397 (N_20397,N_19666,N_19244);
nand U20398 (N_20398,N_19529,N_19791);
nor U20399 (N_20399,N_19405,N_19747);
or U20400 (N_20400,N_19849,N_20384);
nand U20401 (N_20401,N_20060,N_20132);
nor U20402 (N_20402,N_20079,N_20390);
xnor U20403 (N_20403,N_20064,N_20108);
or U20404 (N_20404,N_20349,N_19815);
nand U20405 (N_20405,N_20118,N_20270);
xnor U20406 (N_20406,N_20388,N_20025);
nor U20407 (N_20407,N_20254,N_20179);
nor U20408 (N_20408,N_20346,N_20047);
nor U20409 (N_20409,N_20114,N_19968);
nand U20410 (N_20410,N_19884,N_19911);
or U20411 (N_20411,N_19882,N_20219);
nor U20412 (N_20412,N_20323,N_20351);
xnor U20413 (N_20413,N_19905,N_19890);
or U20414 (N_20414,N_19820,N_20268);
nor U20415 (N_20415,N_19975,N_20028);
or U20416 (N_20416,N_19871,N_20297);
or U20417 (N_20417,N_19955,N_19864);
nand U20418 (N_20418,N_20001,N_20377);
or U20419 (N_20419,N_19943,N_20216);
xor U20420 (N_20420,N_20020,N_19959);
or U20421 (N_20421,N_20033,N_20081);
xnor U20422 (N_20422,N_20151,N_20241);
nor U20423 (N_20423,N_20021,N_19875);
xor U20424 (N_20424,N_20106,N_20343);
nand U20425 (N_20425,N_19831,N_20141);
xnor U20426 (N_20426,N_19936,N_20085);
and U20427 (N_20427,N_20080,N_20253);
or U20428 (N_20428,N_20215,N_20282);
nor U20429 (N_20429,N_19851,N_19869);
or U20430 (N_20430,N_19992,N_19948);
and U20431 (N_20431,N_20133,N_20029);
or U20432 (N_20432,N_20093,N_19967);
xnor U20433 (N_20433,N_19862,N_20199);
nor U20434 (N_20434,N_20014,N_20249);
nor U20435 (N_20435,N_20231,N_20267);
nand U20436 (N_20436,N_20065,N_20069);
or U20437 (N_20437,N_20149,N_19824);
nor U20438 (N_20438,N_20105,N_19819);
nor U20439 (N_20439,N_20389,N_20163);
xnor U20440 (N_20440,N_20359,N_20110);
nand U20441 (N_20441,N_19900,N_20126);
xnor U20442 (N_20442,N_20112,N_20116);
nor U20443 (N_20443,N_20287,N_20053);
nor U20444 (N_20444,N_20102,N_19902);
and U20445 (N_20445,N_20256,N_19913);
nor U20446 (N_20446,N_19969,N_20067);
or U20447 (N_20447,N_20258,N_20094);
xor U20448 (N_20448,N_19855,N_20202);
nor U20449 (N_20449,N_19832,N_20210);
nand U20450 (N_20450,N_20096,N_20058);
nor U20451 (N_20451,N_20399,N_19939);
nor U20452 (N_20452,N_20154,N_20304);
and U20453 (N_20453,N_20095,N_19972);
and U20454 (N_20454,N_20023,N_20172);
xnor U20455 (N_20455,N_20288,N_20034);
xnor U20456 (N_20456,N_20211,N_20123);
xor U20457 (N_20457,N_20305,N_20223);
nand U20458 (N_20458,N_20235,N_20084);
nor U20459 (N_20459,N_20348,N_19870);
nor U20460 (N_20460,N_19945,N_20073);
and U20461 (N_20461,N_19904,N_20015);
xor U20462 (N_20462,N_20307,N_19912);
nand U20463 (N_20463,N_20275,N_20055);
xnor U20464 (N_20464,N_19839,N_20119);
nor U20465 (N_20465,N_19907,N_20208);
nor U20466 (N_20466,N_20378,N_19830);
xor U20467 (N_20467,N_20212,N_19833);
nor U20468 (N_20468,N_20295,N_20313);
nand U20469 (N_20469,N_20056,N_19963);
nand U20470 (N_20470,N_19837,N_20382);
nand U20471 (N_20471,N_19937,N_20276);
nand U20472 (N_20472,N_19922,N_19990);
and U20473 (N_20473,N_19933,N_19858);
nor U20474 (N_20474,N_20257,N_19910);
nand U20475 (N_20475,N_19927,N_20315);
nand U20476 (N_20476,N_20204,N_20309);
nor U20477 (N_20477,N_20319,N_19845);
xor U20478 (N_20478,N_20049,N_20003);
nor U20479 (N_20479,N_20146,N_20035);
nand U20480 (N_20480,N_20284,N_20018);
nor U20481 (N_20481,N_20252,N_20063);
nand U20482 (N_20482,N_20243,N_19853);
xnor U20483 (N_20483,N_19818,N_20166);
xor U20484 (N_20484,N_19800,N_20225);
xor U20485 (N_20485,N_20331,N_19957);
nor U20486 (N_20486,N_19810,N_20074);
nand U20487 (N_20487,N_20228,N_19899);
or U20488 (N_20488,N_20037,N_20168);
nand U20489 (N_20489,N_19821,N_20277);
xnor U20490 (N_20490,N_20261,N_20247);
xor U20491 (N_20491,N_19987,N_19892);
nor U20492 (N_20492,N_19895,N_20008);
nand U20493 (N_20493,N_20042,N_19893);
or U20494 (N_20494,N_20338,N_19982);
and U20495 (N_20495,N_20143,N_20005);
and U20496 (N_20496,N_19838,N_19852);
xor U20497 (N_20497,N_19984,N_19879);
and U20498 (N_20498,N_19932,N_20145);
or U20499 (N_20499,N_19919,N_20156);
or U20500 (N_20500,N_19897,N_20299);
and U20501 (N_20501,N_20242,N_19876);
or U20502 (N_20502,N_20398,N_19966);
or U20503 (N_20503,N_19944,N_20387);
and U20504 (N_20504,N_20396,N_20341);
nor U20505 (N_20505,N_19938,N_20158);
nand U20506 (N_20506,N_20367,N_19965);
and U20507 (N_20507,N_20054,N_19964);
or U20508 (N_20508,N_20109,N_19806);
or U20509 (N_20509,N_20027,N_19998);
and U20510 (N_20510,N_20385,N_20153);
nand U20511 (N_20511,N_19813,N_19925);
nor U20512 (N_20512,N_19835,N_19951);
xnor U20513 (N_20513,N_19881,N_20302);
nand U20514 (N_20514,N_20129,N_19947);
nand U20515 (N_20515,N_20329,N_19986);
nand U20516 (N_20516,N_20115,N_19974);
nand U20517 (N_20517,N_20052,N_20381);
xnor U20518 (N_20518,N_20190,N_20019);
and U20519 (N_20519,N_20180,N_20236);
nor U20520 (N_20520,N_20357,N_19809);
and U20521 (N_20521,N_19954,N_20328);
or U20522 (N_20522,N_20188,N_20321);
and U20523 (N_20523,N_19917,N_19956);
or U20524 (N_20524,N_20195,N_20246);
nor U20525 (N_20525,N_20237,N_20292);
xnor U20526 (N_20526,N_20167,N_20009);
or U20527 (N_20527,N_20193,N_19916);
and U20528 (N_20528,N_20317,N_20135);
or U20529 (N_20529,N_20233,N_20379);
or U20530 (N_20530,N_20181,N_19977);
xor U20531 (N_20531,N_19908,N_19867);
xnor U20532 (N_20532,N_20333,N_20250);
nand U20533 (N_20533,N_19903,N_20248);
xor U20534 (N_20534,N_19920,N_20010);
nor U20535 (N_20535,N_20362,N_20170);
or U20536 (N_20536,N_20368,N_20306);
nor U20537 (N_20537,N_20087,N_20113);
or U20538 (N_20538,N_19921,N_20344);
nand U20539 (N_20539,N_20002,N_19880);
and U20540 (N_20540,N_19953,N_20314);
and U20541 (N_20541,N_19988,N_19811);
nand U20542 (N_20542,N_20312,N_20334);
nor U20543 (N_20543,N_19914,N_20030);
nand U20544 (N_20544,N_20175,N_20298);
or U20545 (N_20545,N_20140,N_20206);
nor U20546 (N_20546,N_20209,N_20361);
nand U20547 (N_20547,N_19841,N_19950);
nor U20548 (N_20548,N_20251,N_20061);
nand U20549 (N_20549,N_19889,N_19850);
or U20550 (N_20550,N_20092,N_19981);
nand U20551 (N_20551,N_20189,N_20320);
nand U20552 (N_20552,N_20201,N_19842);
nand U20553 (N_20553,N_20230,N_20150);
or U20554 (N_20554,N_19995,N_20066);
xnor U20555 (N_20555,N_20335,N_20264);
and U20556 (N_20556,N_20383,N_20301);
or U20557 (N_20557,N_20183,N_20192);
xnor U20558 (N_20558,N_20038,N_20281);
and U20559 (N_20559,N_19847,N_20148);
and U20560 (N_20560,N_19989,N_20220);
and U20561 (N_20561,N_19859,N_19861);
or U20562 (N_20562,N_19874,N_20017);
xnor U20563 (N_20563,N_20043,N_20280);
xor U20564 (N_20564,N_20016,N_19926);
nand U20565 (N_20565,N_20300,N_19823);
and U20566 (N_20566,N_20200,N_20380);
xor U20567 (N_20567,N_19808,N_20031);
and U20568 (N_20568,N_20296,N_20391);
nand U20569 (N_20569,N_20138,N_20173);
xor U20570 (N_20570,N_20157,N_20244);
xnor U20571 (N_20571,N_20229,N_20086);
nor U20572 (N_20572,N_20185,N_20291);
and U20573 (N_20573,N_20271,N_20041);
nand U20574 (N_20574,N_20234,N_19886);
nor U20575 (N_20575,N_20187,N_20012);
or U20576 (N_20576,N_20191,N_20286);
and U20577 (N_20577,N_20059,N_19976);
nand U20578 (N_20578,N_20144,N_19878);
and U20579 (N_20579,N_20360,N_20325);
and U20580 (N_20580,N_20217,N_19906);
and U20581 (N_20581,N_20111,N_19931);
or U20582 (N_20582,N_20356,N_19877);
nor U20583 (N_20583,N_20071,N_19901);
xor U20584 (N_20584,N_19940,N_20162);
xor U20585 (N_20585,N_19962,N_19865);
and U20586 (N_20586,N_20178,N_19896);
xor U20587 (N_20587,N_20026,N_19996);
or U20588 (N_20588,N_19848,N_20006);
or U20589 (N_20589,N_20121,N_19985);
or U20590 (N_20590,N_19812,N_20363);
and U20591 (N_20591,N_19804,N_20130);
nand U20592 (N_20592,N_20330,N_19816);
and U20593 (N_20593,N_20366,N_19873);
and U20594 (N_20594,N_20186,N_20039);
or U20595 (N_20595,N_20197,N_20050);
nand U20596 (N_20596,N_20177,N_19872);
and U20597 (N_20597,N_20290,N_20207);
or U20598 (N_20598,N_19843,N_20278);
xor U20599 (N_20599,N_20160,N_20048);
nor U20600 (N_20600,N_20159,N_20373);
xnor U20601 (N_20601,N_19826,N_20164);
and U20602 (N_20602,N_20392,N_20337);
nor U20603 (N_20603,N_20024,N_20322);
nand U20604 (N_20604,N_20386,N_19817);
and U20605 (N_20605,N_19979,N_20355);
xor U20606 (N_20606,N_20353,N_19929);
or U20607 (N_20607,N_20262,N_20013);
nand U20608 (N_20608,N_20098,N_20097);
nor U20609 (N_20609,N_19840,N_20255);
and U20610 (N_20610,N_19803,N_20032);
xnor U20611 (N_20611,N_20125,N_19997);
nand U20612 (N_20612,N_20263,N_20342);
or U20613 (N_20613,N_20269,N_19814);
nor U20614 (N_20614,N_19888,N_19822);
or U20615 (N_20615,N_19894,N_20137);
nand U20616 (N_20616,N_20226,N_19999);
or U20617 (N_20617,N_20293,N_19891);
nor U20618 (N_20618,N_20265,N_20283);
or U20619 (N_20619,N_19883,N_20107);
or U20620 (N_20620,N_20345,N_20104);
and U20621 (N_20621,N_20311,N_20174);
xnor U20622 (N_20622,N_20161,N_19856);
xnor U20623 (N_20623,N_19898,N_20101);
xnor U20624 (N_20624,N_20395,N_19994);
or U20625 (N_20625,N_20303,N_19935);
xor U20626 (N_20626,N_20134,N_19961);
nor U20627 (N_20627,N_20279,N_20176);
and U20628 (N_20628,N_20272,N_20376);
or U20629 (N_20629,N_20289,N_19960);
or U20630 (N_20630,N_19983,N_19829);
nor U20631 (N_20631,N_20222,N_20308);
and U20632 (N_20632,N_20182,N_20318);
xor U20633 (N_20633,N_20044,N_19846);
and U20634 (N_20634,N_20294,N_20128);
xnor U20635 (N_20635,N_20324,N_20165);
or U20636 (N_20636,N_20310,N_20045);
xnor U20637 (N_20637,N_20122,N_20062);
nand U20638 (N_20638,N_19993,N_20022);
and U20639 (N_20639,N_20224,N_20078);
nor U20640 (N_20640,N_20273,N_20046);
nand U20641 (N_20641,N_20371,N_19978);
or U20642 (N_20642,N_19958,N_20394);
xor U20643 (N_20643,N_20011,N_20198);
nor U20644 (N_20644,N_20365,N_20089);
and U20645 (N_20645,N_20239,N_19923);
xnor U20646 (N_20646,N_20051,N_19930);
or U20647 (N_20647,N_20375,N_19827);
or U20648 (N_20648,N_20099,N_19909);
xnor U20649 (N_20649,N_20169,N_20120);
xor U20650 (N_20650,N_19834,N_19941);
nand U20651 (N_20651,N_19866,N_20124);
and U20652 (N_20652,N_20326,N_19825);
or U20653 (N_20653,N_20088,N_20076);
nand U20654 (N_20654,N_19952,N_20354);
or U20655 (N_20655,N_20332,N_20370);
xnor U20656 (N_20656,N_20036,N_19802);
and U20657 (N_20657,N_20007,N_20194);
nor U20658 (N_20658,N_19973,N_20091);
nand U20659 (N_20659,N_19946,N_20260);
xnor U20660 (N_20660,N_19805,N_19857);
and U20661 (N_20661,N_19887,N_19915);
nor U20662 (N_20662,N_20218,N_20117);
nor U20663 (N_20663,N_20147,N_19836);
xor U20664 (N_20664,N_20374,N_19801);
or U20665 (N_20665,N_20327,N_20372);
or U20666 (N_20666,N_20227,N_20100);
or U20667 (N_20667,N_20340,N_20203);
or U20668 (N_20668,N_20364,N_20238);
nor U20669 (N_20669,N_20393,N_20127);
or U20670 (N_20670,N_20214,N_20083);
nor U20671 (N_20671,N_20090,N_20232);
and U20672 (N_20672,N_20245,N_20339);
nand U20673 (N_20673,N_20316,N_20136);
or U20674 (N_20674,N_20139,N_19980);
nand U20675 (N_20675,N_19970,N_20077);
nor U20676 (N_20676,N_19868,N_20142);
nor U20677 (N_20677,N_19860,N_20266);
or U20678 (N_20678,N_19934,N_20075);
or U20679 (N_20679,N_20131,N_19863);
nor U20680 (N_20680,N_20205,N_19844);
nor U20681 (N_20681,N_20155,N_20082);
and U20682 (N_20682,N_20171,N_19949);
xor U20683 (N_20683,N_20196,N_20350);
or U20684 (N_20684,N_20068,N_20184);
nor U20685 (N_20685,N_20336,N_20274);
nor U20686 (N_20686,N_19928,N_20369);
xor U20687 (N_20687,N_19971,N_20259);
or U20688 (N_20688,N_20072,N_20358);
or U20689 (N_20689,N_20347,N_20285);
nor U20690 (N_20690,N_20240,N_20397);
and U20691 (N_20691,N_20000,N_19828);
xnor U20692 (N_20692,N_19924,N_19807);
and U20693 (N_20693,N_19991,N_20152);
nand U20694 (N_20694,N_20221,N_19885);
or U20695 (N_20695,N_20057,N_20004);
or U20696 (N_20696,N_19918,N_20040);
nor U20697 (N_20697,N_20213,N_19942);
or U20698 (N_20698,N_20070,N_19854);
and U20699 (N_20699,N_20103,N_20352);
or U20700 (N_20700,N_20129,N_20231);
xnor U20701 (N_20701,N_20224,N_20352);
and U20702 (N_20702,N_19881,N_20139);
nand U20703 (N_20703,N_20197,N_20342);
and U20704 (N_20704,N_19924,N_20173);
nor U20705 (N_20705,N_20300,N_19992);
nand U20706 (N_20706,N_19974,N_20199);
nand U20707 (N_20707,N_20240,N_20144);
or U20708 (N_20708,N_19958,N_19843);
or U20709 (N_20709,N_20129,N_20056);
or U20710 (N_20710,N_20319,N_20180);
xor U20711 (N_20711,N_19836,N_20327);
or U20712 (N_20712,N_20102,N_19831);
and U20713 (N_20713,N_20394,N_20030);
or U20714 (N_20714,N_20379,N_20380);
nand U20715 (N_20715,N_20303,N_20252);
xnor U20716 (N_20716,N_19931,N_19942);
nand U20717 (N_20717,N_20307,N_20066);
xnor U20718 (N_20718,N_20075,N_19854);
or U20719 (N_20719,N_20316,N_19866);
and U20720 (N_20720,N_20169,N_19974);
xnor U20721 (N_20721,N_19888,N_20252);
or U20722 (N_20722,N_20019,N_20336);
nand U20723 (N_20723,N_20139,N_20130);
nor U20724 (N_20724,N_20318,N_20121);
nand U20725 (N_20725,N_20266,N_20025);
or U20726 (N_20726,N_19979,N_20153);
or U20727 (N_20727,N_20087,N_19813);
nor U20728 (N_20728,N_19900,N_20095);
and U20729 (N_20729,N_19979,N_20042);
nor U20730 (N_20730,N_19965,N_20356);
and U20731 (N_20731,N_20076,N_19845);
xor U20732 (N_20732,N_20368,N_19892);
nand U20733 (N_20733,N_20279,N_19946);
or U20734 (N_20734,N_20032,N_20365);
nand U20735 (N_20735,N_20028,N_20236);
or U20736 (N_20736,N_20130,N_19815);
nand U20737 (N_20737,N_20058,N_19975);
xor U20738 (N_20738,N_20188,N_20327);
or U20739 (N_20739,N_19951,N_19856);
xnor U20740 (N_20740,N_19840,N_20091);
nor U20741 (N_20741,N_20391,N_19901);
and U20742 (N_20742,N_20393,N_20192);
or U20743 (N_20743,N_20281,N_20241);
or U20744 (N_20744,N_20294,N_19810);
xor U20745 (N_20745,N_19827,N_20257);
or U20746 (N_20746,N_19855,N_19931);
nor U20747 (N_20747,N_19990,N_19974);
or U20748 (N_20748,N_20336,N_20102);
xor U20749 (N_20749,N_20273,N_20365);
nand U20750 (N_20750,N_20076,N_20025);
or U20751 (N_20751,N_19920,N_19851);
and U20752 (N_20752,N_19946,N_20320);
nor U20753 (N_20753,N_20236,N_20192);
or U20754 (N_20754,N_20245,N_20325);
and U20755 (N_20755,N_20152,N_19937);
or U20756 (N_20756,N_20364,N_20147);
nand U20757 (N_20757,N_20290,N_20279);
nor U20758 (N_20758,N_20004,N_20082);
or U20759 (N_20759,N_20220,N_20244);
nand U20760 (N_20760,N_20398,N_20241);
nand U20761 (N_20761,N_20176,N_20239);
xor U20762 (N_20762,N_20021,N_20209);
or U20763 (N_20763,N_20080,N_19820);
or U20764 (N_20764,N_20113,N_19851);
nor U20765 (N_20765,N_20128,N_20194);
or U20766 (N_20766,N_20223,N_20216);
nor U20767 (N_20767,N_20282,N_20230);
and U20768 (N_20768,N_20002,N_20365);
and U20769 (N_20769,N_20374,N_20105);
and U20770 (N_20770,N_20084,N_20265);
xor U20771 (N_20771,N_20067,N_20198);
or U20772 (N_20772,N_19964,N_20322);
nor U20773 (N_20773,N_19801,N_20081);
and U20774 (N_20774,N_19923,N_20257);
and U20775 (N_20775,N_20094,N_20237);
nand U20776 (N_20776,N_19919,N_20136);
nand U20777 (N_20777,N_20158,N_20012);
nand U20778 (N_20778,N_19929,N_19883);
nor U20779 (N_20779,N_20353,N_19803);
nand U20780 (N_20780,N_20166,N_19864);
nor U20781 (N_20781,N_20030,N_20029);
or U20782 (N_20782,N_20225,N_20129);
and U20783 (N_20783,N_20363,N_19978);
nand U20784 (N_20784,N_20155,N_20215);
xor U20785 (N_20785,N_20248,N_20116);
nor U20786 (N_20786,N_20186,N_20270);
or U20787 (N_20787,N_19863,N_20104);
xor U20788 (N_20788,N_20234,N_20151);
and U20789 (N_20789,N_20385,N_20374);
or U20790 (N_20790,N_20183,N_20097);
and U20791 (N_20791,N_20091,N_20389);
or U20792 (N_20792,N_19809,N_20134);
nand U20793 (N_20793,N_20248,N_20012);
or U20794 (N_20794,N_19901,N_20155);
or U20795 (N_20795,N_20233,N_20365);
nor U20796 (N_20796,N_20156,N_20175);
or U20797 (N_20797,N_20352,N_20136);
nand U20798 (N_20798,N_20312,N_19940);
xnor U20799 (N_20799,N_20218,N_20009);
nand U20800 (N_20800,N_20085,N_20136);
nand U20801 (N_20801,N_20018,N_19908);
nor U20802 (N_20802,N_20282,N_19983);
nor U20803 (N_20803,N_20059,N_20101);
nor U20804 (N_20804,N_20006,N_20093);
xnor U20805 (N_20805,N_19977,N_19984);
or U20806 (N_20806,N_20050,N_20062);
and U20807 (N_20807,N_19985,N_20380);
and U20808 (N_20808,N_20286,N_20066);
and U20809 (N_20809,N_20215,N_20032);
nand U20810 (N_20810,N_19848,N_20201);
nand U20811 (N_20811,N_20351,N_20008);
nor U20812 (N_20812,N_19983,N_20360);
and U20813 (N_20813,N_19869,N_19980);
or U20814 (N_20814,N_20027,N_20392);
and U20815 (N_20815,N_20301,N_20156);
xor U20816 (N_20816,N_20262,N_20329);
or U20817 (N_20817,N_20042,N_19858);
nand U20818 (N_20818,N_20392,N_20048);
xor U20819 (N_20819,N_20351,N_19811);
nor U20820 (N_20820,N_20194,N_20058);
nor U20821 (N_20821,N_20008,N_19910);
xnor U20822 (N_20822,N_20147,N_19865);
or U20823 (N_20823,N_20338,N_20173);
or U20824 (N_20824,N_20259,N_20117);
and U20825 (N_20825,N_20027,N_20044);
and U20826 (N_20826,N_20363,N_20287);
nor U20827 (N_20827,N_19982,N_20014);
xnor U20828 (N_20828,N_19841,N_20109);
and U20829 (N_20829,N_19823,N_20198);
nand U20830 (N_20830,N_19805,N_20258);
or U20831 (N_20831,N_20204,N_20125);
or U20832 (N_20832,N_20122,N_19972);
and U20833 (N_20833,N_20063,N_20117);
nor U20834 (N_20834,N_20355,N_20054);
or U20835 (N_20835,N_20384,N_19976);
xor U20836 (N_20836,N_20338,N_19961);
nor U20837 (N_20837,N_20328,N_19909);
or U20838 (N_20838,N_19948,N_20322);
xor U20839 (N_20839,N_19987,N_20135);
nor U20840 (N_20840,N_20321,N_19842);
xor U20841 (N_20841,N_20275,N_20067);
or U20842 (N_20842,N_20300,N_20395);
nand U20843 (N_20843,N_20224,N_20127);
nor U20844 (N_20844,N_19893,N_19854);
nand U20845 (N_20845,N_20004,N_20025);
and U20846 (N_20846,N_20097,N_19853);
and U20847 (N_20847,N_19902,N_20377);
xor U20848 (N_20848,N_19977,N_20351);
nand U20849 (N_20849,N_19839,N_20082);
nand U20850 (N_20850,N_20168,N_20102);
nand U20851 (N_20851,N_20162,N_20067);
nand U20852 (N_20852,N_20286,N_20169);
nand U20853 (N_20853,N_20126,N_19873);
nor U20854 (N_20854,N_20076,N_20082);
xor U20855 (N_20855,N_19931,N_20317);
and U20856 (N_20856,N_19839,N_19928);
nand U20857 (N_20857,N_20216,N_20188);
nor U20858 (N_20858,N_20198,N_20389);
and U20859 (N_20859,N_20300,N_19929);
nor U20860 (N_20860,N_20015,N_19921);
and U20861 (N_20861,N_20065,N_19951);
nor U20862 (N_20862,N_19957,N_20399);
and U20863 (N_20863,N_19860,N_20062);
xor U20864 (N_20864,N_20007,N_20150);
nor U20865 (N_20865,N_20056,N_20097);
or U20866 (N_20866,N_20397,N_20378);
or U20867 (N_20867,N_20341,N_20275);
or U20868 (N_20868,N_20189,N_20119);
nor U20869 (N_20869,N_20308,N_20185);
nand U20870 (N_20870,N_20388,N_19842);
or U20871 (N_20871,N_20261,N_19828);
nor U20872 (N_20872,N_19931,N_20139);
xnor U20873 (N_20873,N_19875,N_20160);
xnor U20874 (N_20874,N_20077,N_20047);
or U20875 (N_20875,N_20088,N_20062);
or U20876 (N_20876,N_19865,N_20307);
and U20877 (N_20877,N_20023,N_20357);
and U20878 (N_20878,N_20095,N_19998);
xor U20879 (N_20879,N_20229,N_20234);
or U20880 (N_20880,N_20078,N_20302);
and U20881 (N_20881,N_20334,N_19903);
nor U20882 (N_20882,N_19878,N_20182);
or U20883 (N_20883,N_20333,N_20156);
nand U20884 (N_20884,N_19879,N_20248);
or U20885 (N_20885,N_19814,N_20134);
xor U20886 (N_20886,N_19986,N_20315);
or U20887 (N_20887,N_20200,N_20005);
or U20888 (N_20888,N_20179,N_20242);
nand U20889 (N_20889,N_20283,N_19851);
nand U20890 (N_20890,N_19933,N_19961);
nor U20891 (N_20891,N_19835,N_20035);
nand U20892 (N_20892,N_20240,N_19819);
nand U20893 (N_20893,N_20059,N_19839);
nor U20894 (N_20894,N_20137,N_19825);
or U20895 (N_20895,N_19926,N_19879);
or U20896 (N_20896,N_20058,N_20209);
and U20897 (N_20897,N_20222,N_20383);
nand U20898 (N_20898,N_19801,N_19849);
and U20899 (N_20899,N_20034,N_20170);
nor U20900 (N_20900,N_20143,N_20166);
and U20901 (N_20901,N_20140,N_19869);
and U20902 (N_20902,N_20155,N_20216);
nand U20903 (N_20903,N_19852,N_20203);
or U20904 (N_20904,N_19813,N_20284);
xnor U20905 (N_20905,N_20304,N_20252);
nor U20906 (N_20906,N_20137,N_20118);
nand U20907 (N_20907,N_20273,N_20325);
nor U20908 (N_20908,N_19966,N_20136);
and U20909 (N_20909,N_20235,N_20355);
or U20910 (N_20910,N_20024,N_20013);
and U20911 (N_20911,N_19855,N_20316);
nor U20912 (N_20912,N_20169,N_19925);
and U20913 (N_20913,N_19979,N_20323);
xor U20914 (N_20914,N_20293,N_20284);
and U20915 (N_20915,N_20077,N_20054);
and U20916 (N_20916,N_19807,N_20160);
or U20917 (N_20917,N_19892,N_20285);
or U20918 (N_20918,N_20226,N_19904);
and U20919 (N_20919,N_20365,N_20012);
xnor U20920 (N_20920,N_20186,N_20041);
and U20921 (N_20921,N_20342,N_20268);
and U20922 (N_20922,N_19943,N_19818);
nor U20923 (N_20923,N_20223,N_20337);
nor U20924 (N_20924,N_20170,N_20108);
nor U20925 (N_20925,N_19877,N_20045);
nor U20926 (N_20926,N_19819,N_19868);
and U20927 (N_20927,N_20110,N_19975);
nand U20928 (N_20928,N_19963,N_20238);
or U20929 (N_20929,N_20398,N_19967);
nand U20930 (N_20930,N_19903,N_19838);
and U20931 (N_20931,N_20160,N_19842);
xor U20932 (N_20932,N_20116,N_20383);
xor U20933 (N_20933,N_19818,N_20194);
nand U20934 (N_20934,N_19971,N_20347);
or U20935 (N_20935,N_20342,N_20304);
nor U20936 (N_20936,N_20285,N_19850);
nand U20937 (N_20937,N_20135,N_20222);
xnor U20938 (N_20938,N_20120,N_19901);
nor U20939 (N_20939,N_20193,N_20212);
and U20940 (N_20940,N_20215,N_19920);
xor U20941 (N_20941,N_20335,N_19913);
nor U20942 (N_20942,N_19833,N_20068);
nor U20943 (N_20943,N_20285,N_20245);
nor U20944 (N_20944,N_20124,N_19854);
nor U20945 (N_20945,N_20248,N_20258);
and U20946 (N_20946,N_20115,N_20296);
and U20947 (N_20947,N_20105,N_20278);
and U20948 (N_20948,N_20078,N_19855);
or U20949 (N_20949,N_19865,N_19824);
nand U20950 (N_20950,N_20233,N_20164);
and U20951 (N_20951,N_20383,N_19807);
nor U20952 (N_20952,N_20302,N_20355);
xnor U20953 (N_20953,N_20012,N_20131);
nor U20954 (N_20954,N_20376,N_19959);
nand U20955 (N_20955,N_20095,N_20051);
or U20956 (N_20956,N_20063,N_20050);
or U20957 (N_20957,N_19936,N_19876);
and U20958 (N_20958,N_20001,N_20163);
xnor U20959 (N_20959,N_19824,N_20107);
or U20960 (N_20960,N_19967,N_19827);
nor U20961 (N_20961,N_19881,N_20366);
and U20962 (N_20962,N_20319,N_20141);
xor U20963 (N_20963,N_20121,N_20326);
nand U20964 (N_20964,N_20121,N_19940);
nand U20965 (N_20965,N_20156,N_19952);
or U20966 (N_20966,N_20115,N_20317);
and U20967 (N_20967,N_20113,N_20329);
or U20968 (N_20968,N_20029,N_20250);
and U20969 (N_20969,N_20097,N_19993);
xor U20970 (N_20970,N_19877,N_20185);
nand U20971 (N_20971,N_20119,N_20019);
and U20972 (N_20972,N_19827,N_19839);
nand U20973 (N_20973,N_20202,N_19831);
nor U20974 (N_20974,N_19923,N_19999);
xor U20975 (N_20975,N_20221,N_19936);
nor U20976 (N_20976,N_20056,N_20006);
nand U20977 (N_20977,N_20196,N_19846);
xnor U20978 (N_20978,N_20399,N_20082);
xor U20979 (N_20979,N_20301,N_20118);
xor U20980 (N_20980,N_19828,N_20002);
and U20981 (N_20981,N_19846,N_20349);
and U20982 (N_20982,N_20080,N_20384);
or U20983 (N_20983,N_20212,N_19886);
nand U20984 (N_20984,N_19865,N_19985);
nand U20985 (N_20985,N_20049,N_19823);
xor U20986 (N_20986,N_20042,N_20213);
nor U20987 (N_20987,N_19980,N_19859);
or U20988 (N_20988,N_19886,N_20268);
or U20989 (N_20989,N_20097,N_20086);
nand U20990 (N_20990,N_20137,N_20152);
or U20991 (N_20991,N_19967,N_20313);
xor U20992 (N_20992,N_20217,N_20095);
or U20993 (N_20993,N_19827,N_19945);
nor U20994 (N_20994,N_20294,N_19816);
nor U20995 (N_20995,N_20327,N_19808);
xnor U20996 (N_20996,N_20297,N_20155);
nor U20997 (N_20997,N_20057,N_20107);
nand U20998 (N_20998,N_20030,N_19801);
nor U20999 (N_20999,N_19817,N_20252);
nor U21000 (N_21000,N_20443,N_20942);
nor U21001 (N_21001,N_20422,N_20845);
xor U21002 (N_21002,N_20566,N_20658);
nand U21003 (N_21003,N_20441,N_20812);
xnor U21004 (N_21004,N_20770,N_20484);
xor U21005 (N_21005,N_20819,N_20557);
or U21006 (N_21006,N_20787,N_20535);
nand U21007 (N_21007,N_20984,N_20705);
nand U21008 (N_21008,N_20788,N_20592);
xnor U21009 (N_21009,N_20807,N_20944);
nor U21010 (N_21010,N_20527,N_20813);
or U21011 (N_21011,N_20828,N_20683);
nand U21012 (N_21012,N_20682,N_20684);
and U21013 (N_21013,N_20790,N_20718);
xor U21014 (N_21014,N_20757,N_20693);
and U21015 (N_21015,N_20425,N_20629);
nor U21016 (N_21016,N_20521,N_20438);
and U21017 (N_21017,N_20724,N_20404);
nand U21018 (N_21018,N_20667,N_20554);
and U21019 (N_21019,N_20433,N_20940);
or U21020 (N_21020,N_20478,N_20897);
and U21021 (N_21021,N_20495,N_20687);
and U21022 (N_21022,N_20526,N_20427);
xor U21023 (N_21023,N_20926,N_20910);
and U21024 (N_21024,N_20922,N_20925);
and U21025 (N_21025,N_20990,N_20852);
and U21026 (N_21026,N_20830,N_20958);
and U21027 (N_21027,N_20768,N_20500);
nor U21028 (N_21028,N_20496,N_20955);
nor U21029 (N_21029,N_20678,N_20749);
nand U21030 (N_21030,N_20440,N_20502);
nand U21031 (N_21031,N_20746,N_20837);
nand U21032 (N_21032,N_20929,N_20689);
xor U21033 (N_21033,N_20414,N_20664);
nor U21034 (N_21034,N_20821,N_20780);
nor U21035 (N_21035,N_20656,N_20628);
or U21036 (N_21036,N_20459,N_20784);
or U21037 (N_21037,N_20820,N_20983);
xnor U21038 (N_21038,N_20765,N_20904);
and U21039 (N_21039,N_20987,N_20977);
and U21040 (N_21040,N_20593,N_20434);
or U21041 (N_21041,N_20574,N_20832);
nor U21042 (N_21042,N_20776,N_20988);
xnor U21043 (N_21043,N_20709,N_20510);
xnor U21044 (N_21044,N_20612,N_20560);
or U21045 (N_21045,N_20411,N_20453);
nor U21046 (N_21046,N_20786,N_20985);
xnor U21047 (N_21047,N_20512,N_20551);
and U21048 (N_21048,N_20912,N_20748);
nor U21049 (N_21049,N_20546,N_20677);
or U21050 (N_21050,N_20556,N_20669);
or U21051 (N_21051,N_20783,N_20796);
nor U21052 (N_21052,N_20891,N_20811);
or U21053 (N_21053,N_20504,N_20491);
xor U21054 (N_21054,N_20951,N_20753);
and U21055 (N_21055,N_20623,N_20595);
or U21056 (N_21056,N_20727,N_20824);
and U21057 (N_21057,N_20671,N_20485);
and U21058 (N_21058,N_20716,N_20871);
xor U21059 (N_21059,N_20847,N_20465);
and U21060 (N_21060,N_20860,N_20649);
nor U21061 (N_21061,N_20769,N_20948);
or U21062 (N_21062,N_20722,N_20407);
and U21063 (N_21063,N_20594,N_20552);
xnor U21064 (N_21064,N_20581,N_20639);
and U21065 (N_21065,N_20997,N_20607);
nor U21066 (N_21066,N_20516,N_20509);
and U21067 (N_21067,N_20596,N_20720);
or U21068 (N_21068,N_20403,N_20419);
nand U21069 (N_21069,N_20936,N_20890);
nand U21070 (N_21070,N_20576,N_20865);
nand U21071 (N_21071,N_20763,N_20573);
xnor U21072 (N_21072,N_20466,N_20999);
xnor U21073 (N_21073,N_20982,N_20778);
and U21074 (N_21074,N_20801,N_20692);
and U21075 (N_21075,N_20804,N_20672);
xor U21076 (N_21076,N_20809,N_20643);
or U21077 (N_21077,N_20499,N_20698);
nand U21078 (N_21078,N_20651,N_20542);
or U21079 (N_21079,N_20539,N_20442);
and U21080 (N_21080,N_20793,N_20599);
and U21081 (N_21081,N_20645,N_20848);
and U21082 (N_21082,N_20802,N_20879);
or U21083 (N_21083,N_20586,N_20446);
xnor U21084 (N_21084,N_20759,N_20690);
nor U21085 (N_21085,N_20642,N_20590);
and U21086 (N_21086,N_20454,N_20408);
and U21087 (N_21087,N_20471,N_20732);
nand U21088 (N_21088,N_20544,N_20971);
or U21089 (N_21089,N_20436,N_20475);
or U21090 (N_21090,N_20638,N_20700);
nand U21091 (N_21091,N_20470,N_20674);
xnor U21092 (N_21092,N_20726,N_20933);
and U21093 (N_21093,N_20892,N_20834);
xor U21094 (N_21094,N_20872,N_20703);
xnor U21095 (N_21095,N_20901,N_20697);
nor U21096 (N_21096,N_20634,N_20636);
nor U21097 (N_21097,N_20562,N_20616);
xnor U21098 (N_21098,N_20911,N_20917);
and U21099 (N_21099,N_20532,N_20941);
nand U21100 (N_21100,N_20719,N_20928);
or U21101 (N_21101,N_20695,N_20622);
xor U21102 (N_21102,N_20932,N_20754);
or U21103 (N_21103,N_20743,N_20624);
or U21104 (N_21104,N_20898,N_20522);
nand U21105 (N_21105,N_20795,N_20902);
nand U21106 (N_21106,N_20563,N_20827);
and U21107 (N_21107,N_20600,N_20934);
xnor U21108 (N_21108,N_20842,N_20953);
nand U21109 (N_21109,N_20741,N_20733);
or U21110 (N_21110,N_20657,N_20514);
or U21111 (N_21111,N_20416,N_20598);
and U21112 (N_21112,N_20905,N_20742);
or U21113 (N_21113,N_20838,N_20640);
and U21114 (N_21114,N_20931,N_20939);
xnor U21115 (N_21115,N_20791,N_20736);
and U21116 (N_21116,N_20751,N_20921);
nand U21117 (N_21117,N_20670,N_20959);
nand U21118 (N_21118,N_20477,N_20919);
nand U21119 (N_21119,N_20721,N_20655);
nor U21120 (N_21120,N_20960,N_20935);
and U21121 (N_21121,N_20665,N_20775);
and U21122 (N_21122,N_20474,N_20569);
and U21123 (N_21123,N_20806,N_20659);
and U21124 (N_21124,N_20923,N_20980);
and U21125 (N_21125,N_20447,N_20473);
nor U21126 (N_21126,N_20981,N_20601);
nor U21127 (N_21127,N_20895,N_20975);
xnor U21128 (N_21128,N_20798,N_20481);
and U21129 (N_21129,N_20704,N_20409);
xnor U21130 (N_21130,N_20849,N_20861);
and U21131 (N_21131,N_20918,N_20758);
nand U21132 (N_21132,N_20764,N_20702);
nor U21133 (N_21133,N_20762,N_20603);
and U21134 (N_21134,N_20415,N_20448);
xnor U21135 (N_21135,N_20506,N_20854);
nor U21136 (N_21136,N_20886,N_20893);
xor U21137 (N_21137,N_20531,N_20618);
or U21138 (N_21138,N_20549,N_20402);
or U21139 (N_21139,N_20996,N_20688);
or U21140 (N_21140,N_20840,N_20580);
and U21141 (N_21141,N_20881,N_20617);
nand U21142 (N_21142,N_20712,N_20777);
and U21143 (N_21143,N_20497,N_20822);
xnor U21144 (N_21144,N_20545,N_20808);
nand U21145 (N_21145,N_20501,N_20841);
nor U21146 (N_21146,N_20870,N_20486);
and U21147 (N_21147,N_20961,N_20587);
nor U21148 (N_21148,N_20691,N_20851);
xor U21149 (N_21149,N_20467,N_20663);
nor U21150 (N_21150,N_20468,N_20493);
nor U21151 (N_21151,N_20823,N_20550);
nand U21152 (N_21152,N_20469,N_20740);
and U21153 (N_21153,N_20880,N_20737);
xnor U21154 (N_21154,N_20513,N_20745);
xor U21155 (N_21155,N_20952,N_20992);
nor U21156 (N_21156,N_20710,N_20773);
xnor U21157 (N_21157,N_20766,N_20831);
nor U21158 (N_21158,N_20818,N_20458);
nor U21159 (N_21159,N_20701,N_20589);
or U21160 (N_21160,N_20694,N_20767);
xor U21161 (N_21161,N_20924,N_20602);
nor U21162 (N_21162,N_20676,N_20613);
or U21163 (N_21163,N_20815,N_20424);
xor U21164 (N_21164,N_20972,N_20578);
xnor U21165 (N_21165,N_20888,N_20876);
nand U21166 (N_21166,N_20875,N_20826);
nor U21167 (N_21167,N_20614,N_20857);
or U21168 (N_21168,N_20555,N_20947);
and U21169 (N_21169,N_20973,N_20583);
xnor U21170 (N_21170,N_20604,N_20547);
xnor U21171 (N_21171,N_20487,N_20906);
nor U21172 (N_21172,N_20401,N_20445);
and U21173 (N_21173,N_20882,N_20889);
and U21174 (N_21174,N_20456,N_20619);
and U21175 (N_21175,N_20633,N_20885);
nor U21176 (N_21176,N_20797,N_20913);
nand U21177 (N_21177,N_20850,N_20452);
and U21178 (N_21178,N_20418,N_20530);
xnor U21179 (N_21179,N_20630,N_20782);
nand U21180 (N_21180,N_20867,N_20426);
nor U21181 (N_21181,N_20582,N_20538);
nand U21182 (N_21182,N_20877,N_20781);
nor U21183 (N_21183,N_20611,N_20428);
and U21184 (N_21184,N_20711,N_20728);
nor U21185 (N_21185,N_20699,N_20779);
or U21186 (N_21186,N_20579,N_20998);
nor U21187 (N_21187,N_20641,N_20839);
and U21188 (N_21188,N_20654,N_20956);
xor U21189 (N_21189,N_20540,N_20750);
xnor U21190 (N_21190,N_20537,N_20627);
xor U21191 (N_21191,N_20489,N_20863);
and U21192 (N_21192,N_20462,N_20508);
xor U21193 (N_21193,N_20943,N_20853);
and U21194 (N_21194,N_20715,N_20479);
xor U21195 (N_21195,N_20644,N_20605);
and U21196 (N_21196,N_20785,N_20457);
nor U21197 (N_21197,N_20417,N_20978);
nand U21198 (N_21198,N_20472,N_20957);
nor U21199 (N_21199,N_20883,N_20950);
xor U21200 (N_21200,N_20967,N_20615);
nor U21201 (N_21201,N_20874,N_20761);
xor U21202 (N_21202,N_20518,N_20482);
and U21203 (N_21203,N_20606,N_20423);
and U21204 (N_21204,N_20548,N_20543);
nand U21205 (N_21205,N_20650,N_20480);
nand U21206 (N_21206,N_20899,N_20962);
nor U21207 (N_21207,N_20681,N_20439);
and U21208 (N_21208,N_20435,N_20505);
nor U21209 (N_21209,N_20735,N_20631);
and U21210 (N_21210,N_20731,N_20449);
and U21211 (N_21211,N_20564,N_20836);
and U21212 (N_21212,N_20541,N_20561);
nand U21213 (N_21213,N_20954,N_20679);
xnor U21214 (N_21214,N_20507,N_20729);
xnor U21215 (N_21215,N_20575,N_20515);
nand U21216 (N_21216,N_20450,N_20400);
and U21217 (N_21217,N_20844,N_20652);
nor U21218 (N_21218,N_20946,N_20570);
nand U21219 (N_21219,N_20647,N_20829);
and U21220 (N_21220,N_20536,N_20771);
nand U21221 (N_21221,N_20517,N_20523);
nand U21222 (N_21222,N_20963,N_20432);
and U21223 (N_21223,N_20451,N_20637);
and U21224 (N_21224,N_20406,N_20835);
xnor U21225 (N_21225,N_20995,N_20565);
or U21226 (N_21226,N_20744,N_20991);
nor U21227 (N_21227,N_20817,N_20696);
or U21228 (N_21228,N_20410,N_20597);
nand U21229 (N_21229,N_20464,N_20577);
xnor U21230 (N_21230,N_20755,N_20965);
nand U21231 (N_21231,N_20685,N_20666);
xor U21232 (N_21232,N_20794,N_20528);
nand U21233 (N_21233,N_20492,N_20660);
and U21234 (N_21234,N_20520,N_20723);
and U21235 (N_21235,N_20799,N_20585);
nand U21236 (N_21236,N_20909,N_20949);
and U21237 (N_21237,N_20964,N_20412);
or U21238 (N_21238,N_20567,N_20816);
and U21239 (N_21239,N_20534,N_20430);
nand U21240 (N_21240,N_20994,N_20463);
or U21241 (N_21241,N_20490,N_20455);
xnor U21242 (N_21242,N_20814,N_20833);
nand U21243 (N_21243,N_20803,N_20878);
xor U21244 (N_21244,N_20498,N_20646);
nand U21245 (N_21245,N_20460,N_20461);
or U21246 (N_21246,N_20444,N_20713);
nand U21247 (N_21247,N_20900,N_20864);
nand U21248 (N_21248,N_20914,N_20789);
nor U21249 (N_21249,N_20608,N_20553);
nor U21250 (N_21250,N_20869,N_20970);
and U21251 (N_21251,N_20756,N_20989);
nand U21252 (N_21252,N_20525,N_20966);
and U21253 (N_21253,N_20437,N_20862);
nor U21254 (N_21254,N_20421,N_20431);
xor U21255 (N_21255,N_20887,N_20739);
nor U21256 (N_21256,N_20568,N_20420);
or U21257 (N_21257,N_20503,N_20675);
or U21258 (N_21258,N_20571,N_20974);
nand U21259 (N_21259,N_20706,N_20937);
nand U21260 (N_21260,N_20494,N_20686);
xor U21261 (N_21261,N_20609,N_20524);
nand U21262 (N_21262,N_20896,N_20483);
nand U21263 (N_21263,N_20855,N_20846);
or U21264 (N_21264,N_20734,N_20907);
and U21265 (N_21265,N_20635,N_20529);
xnor U21266 (N_21266,N_20976,N_20632);
and U21267 (N_21267,N_20714,N_20730);
or U21268 (N_21268,N_20969,N_20774);
and U21269 (N_21269,N_20866,N_20584);
nand U21270 (N_21270,N_20653,N_20488);
nor U21271 (N_21271,N_20908,N_20738);
and U21272 (N_21272,N_20856,N_20938);
or U21273 (N_21273,N_20413,N_20558);
xor U21274 (N_21274,N_20591,N_20800);
and U21275 (N_21275,N_20626,N_20986);
xnor U21276 (N_21276,N_20873,N_20772);
nand U21277 (N_21277,N_20725,N_20747);
xor U21278 (N_21278,N_20810,N_20621);
nand U21279 (N_21279,N_20519,N_20661);
or U21280 (N_21280,N_20927,N_20945);
nor U21281 (N_21281,N_20668,N_20405);
nor U21282 (N_21282,N_20843,N_20717);
nand U21283 (N_21283,N_20648,N_20792);
xnor U21284 (N_21284,N_20858,N_20708);
nand U21285 (N_21285,N_20884,N_20805);
xor U21286 (N_21286,N_20930,N_20894);
and U21287 (N_21287,N_20915,N_20979);
or U21288 (N_21288,N_20868,N_20859);
and U21289 (N_21289,N_20610,N_20620);
xor U21290 (N_21290,N_20662,N_20760);
or U21291 (N_21291,N_20680,N_20429);
nor U21292 (N_21292,N_20572,N_20993);
xnor U21293 (N_21293,N_20476,N_20920);
and U21294 (N_21294,N_20673,N_20916);
and U21295 (N_21295,N_20559,N_20968);
xor U21296 (N_21296,N_20752,N_20533);
nor U21297 (N_21297,N_20903,N_20625);
or U21298 (N_21298,N_20588,N_20825);
nor U21299 (N_21299,N_20511,N_20707);
nor U21300 (N_21300,N_20993,N_20428);
or U21301 (N_21301,N_20443,N_20612);
and U21302 (N_21302,N_20521,N_20739);
nor U21303 (N_21303,N_20493,N_20439);
xor U21304 (N_21304,N_20759,N_20635);
nand U21305 (N_21305,N_20472,N_20728);
or U21306 (N_21306,N_20441,N_20492);
and U21307 (N_21307,N_20418,N_20861);
or U21308 (N_21308,N_20524,N_20848);
and U21309 (N_21309,N_20519,N_20892);
nor U21310 (N_21310,N_20408,N_20566);
nand U21311 (N_21311,N_20558,N_20688);
or U21312 (N_21312,N_20929,N_20955);
nand U21313 (N_21313,N_20507,N_20525);
and U21314 (N_21314,N_20642,N_20687);
nand U21315 (N_21315,N_20521,N_20792);
nor U21316 (N_21316,N_20752,N_20724);
nand U21317 (N_21317,N_20763,N_20578);
or U21318 (N_21318,N_20630,N_20556);
or U21319 (N_21319,N_20469,N_20819);
or U21320 (N_21320,N_20887,N_20729);
xnor U21321 (N_21321,N_20480,N_20764);
nor U21322 (N_21322,N_20611,N_20435);
xnor U21323 (N_21323,N_20606,N_20693);
and U21324 (N_21324,N_20842,N_20824);
xnor U21325 (N_21325,N_20849,N_20919);
nor U21326 (N_21326,N_20864,N_20653);
nand U21327 (N_21327,N_20519,N_20455);
nand U21328 (N_21328,N_20793,N_20651);
or U21329 (N_21329,N_20419,N_20678);
or U21330 (N_21330,N_20694,N_20729);
xor U21331 (N_21331,N_20635,N_20998);
or U21332 (N_21332,N_20707,N_20549);
nor U21333 (N_21333,N_20949,N_20684);
nand U21334 (N_21334,N_20552,N_20691);
or U21335 (N_21335,N_20793,N_20440);
nor U21336 (N_21336,N_20807,N_20665);
nor U21337 (N_21337,N_20764,N_20437);
nand U21338 (N_21338,N_20888,N_20714);
and U21339 (N_21339,N_20849,N_20988);
nor U21340 (N_21340,N_20730,N_20457);
xnor U21341 (N_21341,N_20758,N_20987);
or U21342 (N_21342,N_20804,N_20898);
xor U21343 (N_21343,N_20757,N_20426);
or U21344 (N_21344,N_20957,N_20809);
and U21345 (N_21345,N_20644,N_20872);
or U21346 (N_21346,N_20580,N_20691);
nand U21347 (N_21347,N_20704,N_20666);
and U21348 (N_21348,N_20755,N_20869);
nor U21349 (N_21349,N_20905,N_20833);
and U21350 (N_21350,N_20697,N_20835);
nand U21351 (N_21351,N_20460,N_20566);
nor U21352 (N_21352,N_20676,N_20678);
xor U21353 (N_21353,N_20459,N_20894);
nor U21354 (N_21354,N_20684,N_20628);
nor U21355 (N_21355,N_20574,N_20732);
nor U21356 (N_21356,N_20489,N_20556);
nor U21357 (N_21357,N_20854,N_20586);
and U21358 (N_21358,N_20815,N_20600);
nand U21359 (N_21359,N_20641,N_20852);
xor U21360 (N_21360,N_20763,N_20494);
nor U21361 (N_21361,N_20898,N_20507);
nor U21362 (N_21362,N_20583,N_20476);
nand U21363 (N_21363,N_20465,N_20568);
or U21364 (N_21364,N_20765,N_20671);
nor U21365 (N_21365,N_20838,N_20867);
or U21366 (N_21366,N_20470,N_20997);
or U21367 (N_21367,N_20709,N_20852);
and U21368 (N_21368,N_20406,N_20652);
or U21369 (N_21369,N_20816,N_20415);
and U21370 (N_21370,N_20844,N_20528);
and U21371 (N_21371,N_20751,N_20980);
or U21372 (N_21372,N_20928,N_20823);
and U21373 (N_21373,N_20835,N_20563);
nand U21374 (N_21374,N_20576,N_20926);
nor U21375 (N_21375,N_20951,N_20601);
and U21376 (N_21376,N_20884,N_20417);
or U21377 (N_21377,N_20408,N_20757);
xor U21378 (N_21378,N_20771,N_20517);
nand U21379 (N_21379,N_20424,N_20843);
or U21380 (N_21380,N_20717,N_20426);
xnor U21381 (N_21381,N_20770,N_20660);
and U21382 (N_21382,N_20575,N_20588);
xor U21383 (N_21383,N_20841,N_20723);
nand U21384 (N_21384,N_20977,N_20787);
or U21385 (N_21385,N_20863,N_20730);
and U21386 (N_21386,N_20422,N_20557);
nor U21387 (N_21387,N_20725,N_20882);
nand U21388 (N_21388,N_20616,N_20544);
nand U21389 (N_21389,N_20693,N_20521);
nor U21390 (N_21390,N_20503,N_20791);
and U21391 (N_21391,N_20758,N_20746);
and U21392 (N_21392,N_20405,N_20606);
and U21393 (N_21393,N_20617,N_20810);
xnor U21394 (N_21394,N_20713,N_20904);
xnor U21395 (N_21395,N_20909,N_20747);
xnor U21396 (N_21396,N_20414,N_20742);
or U21397 (N_21397,N_20422,N_20634);
or U21398 (N_21398,N_20789,N_20888);
xor U21399 (N_21399,N_20442,N_20931);
and U21400 (N_21400,N_20801,N_20826);
or U21401 (N_21401,N_20934,N_20719);
and U21402 (N_21402,N_20421,N_20650);
nand U21403 (N_21403,N_20714,N_20845);
and U21404 (N_21404,N_20864,N_20629);
xnor U21405 (N_21405,N_20760,N_20686);
nand U21406 (N_21406,N_20484,N_20551);
nor U21407 (N_21407,N_20654,N_20539);
xnor U21408 (N_21408,N_20831,N_20877);
and U21409 (N_21409,N_20551,N_20940);
xor U21410 (N_21410,N_20873,N_20928);
and U21411 (N_21411,N_20605,N_20773);
or U21412 (N_21412,N_20572,N_20888);
or U21413 (N_21413,N_20786,N_20722);
and U21414 (N_21414,N_20952,N_20887);
nand U21415 (N_21415,N_20905,N_20444);
and U21416 (N_21416,N_20847,N_20539);
or U21417 (N_21417,N_20961,N_20571);
nor U21418 (N_21418,N_20829,N_20621);
or U21419 (N_21419,N_20539,N_20586);
nor U21420 (N_21420,N_20685,N_20490);
nor U21421 (N_21421,N_20988,N_20590);
xor U21422 (N_21422,N_20427,N_20764);
and U21423 (N_21423,N_20639,N_20793);
and U21424 (N_21424,N_20882,N_20536);
nor U21425 (N_21425,N_20694,N_20830);
nor U21426 (N_21426,N_20527,N_20428);
and U21427 (N_21427,N_20411,N_20518);
xor U21428 (N_21428,N_20606,N_20535);
or U21429 (N_21429,N_20724,N_20959);
nand U21430 (N_21430,N_20538,N_20752);
nand U21431 (N_21431,N_20413,N_20577);
nand U21432 (N_21432,N_20857,N_20733);
nand U21433 (N_21433,N_20780,N_20743);
and U21434 (N_21434,N_20890,N_20749);
nand U21435 (N_21435,N_20961,N_20599);
xnor U21436 (N_21436,N_20966,N_20936);
nor U21437 (N_21437,N_20823,N_20954);
nor U21438 (N_21438,N_20695,N_20943);
and U21439 (N_21439,N_20720,N_20406);
and U21440 (N_21440,N_20900,N_20678);
nor U21441 (N_21441,N_20625,N_20601);
xnor U21442 (N_21442,N_20661,N_20772);
or U21443 (N_21443,N_20875,N_20818);
and U21444 (N_21444,N_20480,N_20599);
xor U21445 (N_21445,N_20571,N_20727);
or U21446 (N_21446,N_20796,N_20926);
xor U21447 (N_21447,N_20461,N_20662);
nand U21448 (N_21448,N_20471,N_20453);
xnor U21449 (N_21449,N_20965,N_20879);
or U21450 (N_21450,N_20938,N_20840);
xnor U21451 (N_21451,N_20856,N_20973);
and U21452 (N_21452,N_20571,N_20964);
nor U21453 (N_21453,N_20590,N_20899);
nand U21454 (N_21454,N_20538,N_20484);
nand U21455 (N_21455,N_20892,N_20929);
xor U21456 (N_21456,N_20477,N_20980);
and U21457 (N_21457,N_20655,N_20431);
or U21458 (N_21458,N_20943,N_20890);
and U21459 (N_21459,N_20913,N_20586);
nand U21460 (N_21460,N_20569,N_20793);
or U21461 (N_21461,N_20894,N_20503);
and U21462 (N_21462,N_20621,N_20530);
xnor U21463 (N_21463,N_20503,N_20400);
and U21464 (N_21464,N_20617,N_20468);
and U21465 (N_21465,N_20590,N_20409);
nor U21466 (N_21466,N_20602,N_20940);
and U21467 (N_21467,N_20802,N_20853);
nor U21468 (N_21468,N_20587,N_20511);
xor U21469 (N_21469,N_20688,N_20796);
xor U21470 (N_21470,N_20998,N_20421);
nand U21471 (N_21471,N_20956,N_20553);
or U21472 (N_21472,N_20437,N_20996);
nand U21473 (N_21473,N_20602,N_20747);
nor U21474 (N_21474,N_20834,N_20403);
or U21475 (N_21475,N_20859,N_20838);
and U21476 (N_21476,N_20699,N_20609);
or U21477 (N_21477,N_20626,N_20628);
or U21478 (N_21478,N_20722,N_20628);
and U21479 (N_21479,N_20547,N_20823);
nand U21480 (N_21480,N_20769,N_20929);
xnor U21481 (N_21481,N_20866,N_20832);
xor U21482 (N_21482,N_20512,N_20645);
or U21483 (N_21483,N_20421,N_20779);
or U21484 (N_21484,N_20570,N_20974);
and U21485 (N_21485,N_20679,N_20639);
or U21486 (N_21486,N_20922,N_20480);
or U21487 (N_21487,N_20889,N_20621);
nor U21488 (N_21488,N_20965,N_20528);
nor U21489 (N_21489,N_20919,N_20690);
nand U21490 (N_21490,N_20732,N_20797);
and U21491 (N_21491,N_20457,N_20810);
and U21492 (N_21492,N_20913,N_20491);
xor U21493 (N_21493,N_20526,N_20843);
or U21494 (N_21494,N_20740,N_20644);
xor U21495 (N_21495,N_20801,N_20542);
nor U21496 (N_21496,N_20786,N_20700);
xor U21497 (N_21497,N_20564,N_20852);
nand U21498 (N_21498,N_20642,N_20546);
or U21499 (N_21499,N_20812,N_20728);
xnor U21500 (N_21500,N_20560,N_20628);
nor U21501 (N_21501,N_20989,N_20470);
or U21502 (N_21502,N_20928,N_20761);
and U21503 (N_21503,N_20627,N_20415);
nand U21504 (N_21504,N_20676,N_20686);
xnor U21505 (N_21505,N_20656,N_20835);
nor U21506 (N_21506,N_20905,N_20951);
xor U21507 (N_21507,N_20524,N_20680);
and U21508 (N_21508,N_20415,N_20432);
nand U21509 (N_21509,N_20590,N_20982);
or U21510 (N_21510,N_20692,N_20776);
nor U21511 (N_21511,N_20916,N_20905);
or U21512 (N_21512,N_20699,N_20892);
nor U21513 (N_21513,N_20938,N_20416);
or U21514 (N_21514,N_20508,N_20577);
or U21515 (N_21515,N_20881,N_20544);
xor U21516 (N_21516,N_20514,N_20438);
and U21517 (N_21517,N_20458,N_20616);
xor U21518 (N_21518,N_20564,N_20952);
xnor U21519 (N_21519,N_20457,N_20837);
and U21520 (N_21520,N_20547,N_20754);
and U21521 (N_21521,N_20423,N_20627);
nand U21522 (N_21522,N_20524,N_20826);
nand U21523 (N_21523,N_20700,N_20403);
nand U21524 (N_21524,N_20539,N_20900);
nand U21525 (N_21525,N_20606,N_20471);
or U21526 (N_21526,N_20543,N_20933);
nand U21527 (N_21527,N_20638,N_20923);
and U21528 (N_21528,N_20884,N_20507);
nor U21529 (N_21529,N_20636,N_20760);
and U21530 (N_21530,N_20626,N_20551);
nand U21531 (N_21531,N_20888,N_20555);
or U21532 (N_21532,N_20757,N_20799);
nor U21533 (N_21533,N_20994,N_20497);
or U21534 (N_21534,N_20575,N_20694);
and U21535 (N_21535,N_20871,N_20990);
and U21536 (N_21536,N_20639,N_20435);
nand U21537 (N_21537,N_20697,N_20879);
and U21538 (N_21538,N_20588,N_20754);
nor U21539 (N_21539,N_20955,N_20819);
or U21540 (N_21540,N_20673,N_20863);
and U21541 (N_21541,N_20737,N_20936);
nor U21542 (N_21542,N_20907,N_20848);
or U21543 (N_21543,N_20920,N_20996);
and U21544 (N_21544,N_20553,N_20466);
and U21545 (N_21545,N_20944,N_20556);
or U21546 (N_21546,N_20791,N_20952);
or U21547 (N_21547,N_20420,N_20940);
xnor U21548 (N_21548,N_20696,N_20601);
xnor U21549 (N_21549,N_20962,N_20890);
nand U21550 (N_21550,N_20835,N_20921);
nor U21551 (N_21551,N_20510,N_20875);
nand U21552 (N_21552,N_20456,N_20802);
nand U21553 (N_21553,N_20822,N_20832);
and U21554 (N_21554,N_20554,N_20866);
xor U21555 (N_21555,N_20599,N_20993);
and U21556 (N_21556,N_20633,N_20940);
and U21557 (N_21557,N_20933,N_20785);
nand U21558 (N_21558,N_20914,N_20706);
nand U21559 (N_21559,N_20975,N_20773);
and U21560 (N_21560,N_20480,N_20533);
or U21561 (N_21561,N_20545,N_20910);
and U21562 (N_21562,N_20847,N_20414);
xnor U21563 (N_21563,N_20557,N_20615);
nor U21564 (N_21564,N_20443,N_20737);
or U21565 (N_21565,N_20802,N_20695);
nor U21566 (N_21566,N_20448,N_20781);
and U21567 (N_21567,N_20433,N_20591);
and U21568 (N_21568,N_20750,N_20800);
nand U21569 (N_21569,N_20751,N_20720);
xnor U21570 (N_21570,N_20692,N_20672);
and U21571 (N_21571,N_20923,N_20518);
or U21572 (N_21572,N_20702,N_20408);
nand U21573 (N_21573,N_20707,N_20820);
nor U21574 (N_21574,N_20754,N_20845);
nand U21575 (N_21575,N_20604,N_20811);
nor U21576 (N_21576,N_20785,N_20909);
or U21577 (N_21577,N_20446,N_20459);
or U21578 (N_21578,N_20706,N_20970);
xor U21579 (N_21579,N_20685,N_20970);
or U21580 (N_21580,N_20562,N_20789);
nor U21581 (N_21581,N_20775,N_20863);
or U21582 (N_21582,N_20574,N_20523);
and U21583 (N_21583,N_20785,N_20665);
nor U21584 (N_21584,N_20492,N_20995);
xor U21585 (N_21585,N_20833,N_20942);
and U21586 (N_21586,N_20552,N_20824);
nor U21587 (N_21587,N_20537,N_20540);
and U21588 (N_21588,N_20783,N_20748);
nor U21589 (N_21589,N_20576,N_20773);
nor U21590 (N_21590,N_20929,N_20480);
xnor U21591 (N_21591,N_20942,N_20861);
and U21592 (N_21592,N_20879,N_20767);
or U21593 (N_21593,N_20494,N_20828);
xor U21594 (N_21594,N_20838,N_20711);
nor U21595 (N_21595,N_20467,N_20825);
or U21596 (N_21596,N_20867,N_20760);
xor U21597 (N_21597,N_20816,N_20578);
nand U21598 (N_21598,N_20869,N_20863);
or U21599 (N_21599,N_20474,N_20967);
xnor U21600 (N_21600,N_21515,N_21217);
and U21601 (N_21601,N_21205,N_21302);
and U21602 (N_21602,N_21142,N_21184);
nand U21603 (N_21603,N_21343,N_21255);
or U21604 (N_21604,N_21113,N_21376);
nor U21605 (N_21605,N_21517,N_21228);
nand U21606 (N_21606,N_21103,N_21300);
and U21607 (N_21607,N_21193,N_21249);
and U21608 (N_21608,N_21396,N_21124);
and U21609 (N_21609,N_21083,N_21108);
nand U21610 (N_21610,N_21241,N_21002);
or U21611 (N_21611,N_21243,N_21106);
nand U21612 (N_21612,N_21085,N_21324);
and U21613 (N_21613,N_21474,N_21318);
and U21614 (N_21614,N_21424,N_21366);
xnor U21615 (N_21615,N_21275,N_21251);
nand U21616 (N_21616,N_21309,N_21279);
nand U21617 (N_21617,N_21528,N_21039);
nand U21618 (N_21618,N_21263,N_21478);
nor U21619 (N_21619,N_21487,N_21281);
nor U21620 (N_21620,N_21258,N_21354);
xnor U21621 (N_21621,N_21477,N_21564);
nor U21622 (N_21622,N_21295,N_21118);
nand U21623 (N_21623,N_21047,N_21014);
xnor U21624 (N_21624,N_21015,N_21472);
nand U21625 (N_21625,N_21434,N_21535);
or U21626 (N_21626,N_21270,N_21316);
xnor U21627 (N_21627,N_21598,N_21395);
nor U21628 (N_21628,N_21529,N_21551);
nand U21629 (N_21629,N_21264,N_21596);
or U21630 (N_21630,N_21061,N_21508);
or U21631 (N_21631,N_21076,N_21063);
and U21632 (N_21632,N_21565,N_21233);
nor U21633 (N_21633,N_21473,N_21332);
nand U21634 (N_21634,N_21416,N_21071);
or U21635 (N_21635,N_21078,N_21104);
nor U21636 (N_21636,N_21240,N_21189);
and U21637 (N_21637,N_21326,N_21520);
xor U21638 (N_21638,N_21011,N_21456);
xor U21639 (N_21639,N_21364,N_21589);
and U21640 (N_21640,N_21070,N_21420);
nand U21641 (N_21641,N_21433,N_21499);
nor U21642 (N_21642,N_21563,N_21492);
nor U21643 (N_21643,N_21439,N_21356);
nor U21644 (N_21644,N_21329,N_21448);
and U21645 (N_21645,N_21278,N_21536);
or U21646 (N_21646,N_21408,N_21504);
nor U21647 (N_21647,N_21152,N_21491);
and U21648 (N_21648,N_21144,N_21432);
nand U21649 (N_21649,N_21502,N_21026);
xor U21650 (N_21650,N_21028,N_21007);
or U21651 (N_21651,N_21261,N_21531);
xnor U21652 (N_21652,N_21033,N_21050);
xnor U21653 (N_21653,N_21000,N_21308);
or U21654 (N_21654,N_21120,N_21091);
and U21655 (N_21655,N_21347,N_21181);
or U21656 (N_21656,N_21540,N_21182);
nor U21657 (N_21657,N_21562,N_21032);
nor U21658 (N_21658,N_21558,N_21016);
xnor U21659 (N_21659,N_21280,N_21130);
xor U21660 (N_21660,N_21247,N_21582);
xor U21661 (N_21661,N_21148,N_21094);
and U21662 (N_21662,N_21183,N_21344);
nor U21663 (N_21663,N_21510,N_21315);
xnor U21664 (N_21664,N_21192,N_21284);
nand U21665 (N_21665,N_21579,N_21199);
xnor U21666 (N_21666,N_21285,N_21216);
nand U21667 (N_21667,N_21186,N_21226);
nand U21668 (N_21668,N_21077,N_21069);
nor U21669 (N_21669,N_21330,N_21505);
nand U21670 (N_21670,N_21546,N_21082);
nand U21671 (N_21671,N_21549,N_21494);
nand U21672 (N_21672,N_21321,N_21001);
and U21673 (N_21673,N_21191,N_21572);
nand U21674 (N_21674,N_21341,N_21336);
or U21675 (N_21675,N_21107,N_21252);
nand U21676 (N_21676,N_21170,N_21210);
and U21677 (N_21677,N_21273,N_21570);
nor U21678 (N_21678,N_21381,N_21405);
nand U21679 (N_21679,N_21030,N_21484);
nor U21680 (N_21680,N_21465,N_21274);
nor U21681 (N_21681,N_21559,N_21401);
xor U21682 (N_21682,N_21175,N_21475);
nand U21683 (N_21683,N_21065,N_21455);
or U21684 (N_21684,N_21544,N_21503);
or U21685 (N_21685,N_21486,N_21340);
xor U21686 (N_21686,N_21294,N_21242);
nor U21687 (N_21687,N_21208,N_21173);
xor U21688 (N_21688,N_21483,N_21567);
and U21689 (N_21689,N_21292,N_21522);
nand U21690 (N_21690,N_21176,N_21129);
or U21691 (N_21691,N_21167,N_21542);
xnor U21692 (N_21692,N_21357,N_21196);
xor U21693 (N_21693,N_21037,N_21585);
or U21694 (N_21694,N_21056,N_21360);
and U21695 (N_21695,N_21171,N_21134);
or U21696 (N_21696,N_21438,N_21453);
xnor U21697 (N_21697,N_21010,N_21352);
and U21698 (N_21698,N_21248,N_21121);
xor U21699 (N_21699,N_21501,N_21586);
nand U21700 (N_21700,N_21232,N_21036);
and U21701 (N_21701,N_21337,N_21161);
nor U21702 (N_21702,N_21372,N_21584);
or U21703 (N_21703,N_21268,N_21373);
nand U21704 (N_21704,N_21489,N_21207);
nand U21705 (N_21705,N_21064,N_21402);
or U21706 (N_21706,N_21225,N_21523);
xor U21707 (N_21707,N_21496,N_21224);
xnor U21708 (N_21708,N_21479,N_21490);
nor U21709 (N_21709,N_21098,N_21271);
nor U21710 (N_21710,N_21413,N_21342);
and U21711 (N_21711,N_21172,N_21277);
xor U21712 (N_21712,N_21136,N_21053);
nor U21713 (N_21713,N_21594,N_21051);
or U21714 (N_21714,N_21431,N_21442);
and U21715 (N_21715,N_21404,N_21146);
or U21716 (N_21716,N_21362,N_21027);
nor U21717 (N_21717,N_21304,N_21230);
nand U21718 (N_21718,N_21481,N_21447);
xor U21719 (N_21719,N_21452,N_21338);
or U21720 (N_21720,N_21525,N_21128);
nand U21721 (N_21721,N_21296,N_21310);
nand U21722 (N_21722,N_21539,N_21163);
nor U21723 (N_21723,N_21072,N_21153);
nand U21724 (N_21724,N_21383,N_21157);
xnor U21725 (N_21725,N_21548,N_21417);
xor U21726 (N_21726,N_21080,N_21282);
or U21727 (N_21727,N_21466,N_21099);
or U21728 (N_21728,N_21025,N_21114);
or U21729 (N_21729,N_21235,N_21460);
nand U21730 (N_21730,N_21314,N_21206);
and U21731 (N_21731,N_21555,N_21561);
and U21732 (N_21732,N_21234,N_21526);
nor U21733 (N_21733,N_21110,N_21375);
and U21734 (N_21734,N_21013,N_21493);
nor U21735 (N_21735,N_21265,N_21306);
nor U21736 (N_21736,N_21102,N_21218);
and U21737 (N_21737,N_21412,N_21449);
or U21738 (N_21738,N_21127,N_21334);
and U21739 (N_21739,N_21350,N_21587);
or U21740 (N_21740,N_21188,N_21074);
and U21741 (N_21741,N_21054,N_21131);
nor U21742 (N_21742,N_21327,N_21514);
and U21743 (N_21743,N_21038,N_21174);
nor U21744 (N_21744,N_21155,N_21422);
xnor U21745 (N_21745,N_21221,N_21597);
or U21746 (N_21746,N_21005,N_21214);
nand U21747 (N_21747,N_21397,N_21213);
nor U21748 (N_21748,N_21133,N_21084);
nor U21749 (N_21749,N_21411,N_21035);
nor U21750 (N_21750,N_21569,N_21361);
or U21751 (N_21751,N_21445,N_21331);
and U21752 (N_21752,N_21457,N_21105);
and U21753 (N_21753,N_21394,N_21349);
nand U21754 (N_21754,N_21022,N_21018);
and U21755 (N_21755,N_21003,N_21117);
and U21756 (N_21756,N_21406,N_21165);
or U21757 (N_21757,N_21575,N_21178);
xnor U21758 (N_21758,N_21581,N_21052);
or U21759 (N_21759,N_21593,N_21382);
nor U21760 (N_21760,N_21320,N_21075);
nand U21761 (N_21761,N_21020,N_21081);
and U21762 (N_21762,N_21440,N_21384);
xnor U21763 (N_21763,N_21021,N_21160);
or U21764 (N_21764,N_21513,N_21126);
nor U21765 (N_21765,N_21211,N_21250);
xnor U21766 (N_21766,N_21132,N_21288);
nand U21767 (N_21767,N_21154,N_21556);
nor U21768 (N_21768,N_21290,N_21371);
or U21769 (N_21769,N_21532,N_21599);
or U21770 (N_21770,N_21185,N_21369);
or U21771 (N_21771,N_21591,N_21112);
nor U21772 (N_21772,N_21451,N_21187);
xor U21773 (N_21773,N_21111,N_21253);
or U21774 (N_21774,N_21150,N_21223);
or U21775 (N_21775,N_21500,N_21497);
xnor U21776 (N_21776,N_21339,N_21055);
nor U21777 (N_21777,N_21066,N_21286);
nor U21778 (N_21778,N_21400,N_21348);
and U21779 (N_21779,N_21553,N_21291);
nor U21780 (N_21780,N_21576,N_21059);
or U21781 (N_21781,N_21109,N_21511);
xnor U21782 (N_21782,N_21227,N_21093);
nor U21783 (N_21783,N_21198,N_21518);
nand U21784 (N_21784,N_21380,N_21498);
xnor U21785 (N_21785,N_21436,N_21209);
and U21786 (N_21786,N_21415,N_21495);
nand U21787 (N_21787,N_21123,N_21023);
nand U21788 (N_21788,N_21293,N_21312);
or U21789 (N_21789,N_21289,N_21203);
xor U21790 (N_21790,N_21044,N_21595);
xnor U21791 (N_21791,N_21398,N_21239);
nor U21792 (N_21792,N_21426,N_21096);
or U21793 (N_21793,N_21087,N_21437);
nor U21794 (N_21794,N_21204,N_21097);
and U21795 (N_21795,N_21463,N_21554);
nor U21796 (N_21796,N_21461,N_21159);
or U21797 (N_21797,N_21480,N_21222);
and U21798 (N_21798,N_21201,N_21031);
or U21799 (N_21799,N_21058,N_21399);
nand U21800 (N_21800,N_21244,N_21470);
xor U21801 (N_21801,N_21215,N_21237);
and U21802 (N_21802,N_21212,N_21138);
or U21803 (N_21803,N_21578,N_21393);
nand U21804 (N_21804,N_21158,N_21229);
or U21805 (N_21805,N_21527,N_21267);
nand U21806 (N_21806,N_21335,N_21390);
nor U21807 (N_21807,N_21303,N_21004);
xnor U21808 (N_21808,N_21116,N_21313);
nor U21809 (N_21809,N_21040,N_21177);
and U21810 (N_21810,N_21180,N_21409);
xnor U21811 (N_21811,N_21557,N_21092);
xnor U21812 (N_21812,N_21387,N_21143);
and U21813 (N_21813,N_21179,N_21482);
or U21814 (N_21814,N_21485,N_21122);
nor U21815 (N_21815,N_21137,N_21245);
or U21816 (N_21816,N_21538,N_21574);
xor U21817 (N_21817,N_21086,N_21365);
and U21818 (N_21818,N_21311,N_21141);
nor U21819 (N_21819,N_21101,N_21095);
nand U21820 (N_21820,N_21552,N_21236);
nor U21821 (N_21821,N_21471,N_21287);
or U21822 (N_21822,N_21543,N_21301);
and U21823 (N_21823,N_21467,N_21443);
nand U21824 (N_21824,N_21149,N_21317);
xor U21825 (N_21825,N_21363,N_21430);
nor U21826 (N_21826,N_21389,N_21385);
or U21827 (N_21827,N_21017,N_21043);
or U21828 (N_21828,N_21088,N_21298);
nor U21829 (N_21829,N_21333,N_21029);
and U21830 (N_21830,N_21592,N_21168);
nand U21831 (N_21831,N_21115,N_21519);
nor U21832 (N_21832,N_21260,N_21462);
nand U21833 (N_21833,N_21266,N_21435);
and U21834 (N_21834,N_21571,N_21200);
nor U21835 (N_21835,N_21269,N_21524);
and U21836 (N_21836,N_21568,N_21469);
xnor U21837 (N_21837,N_21046,N_21425);
or U21838 (N_21838,N_21533,N_21060);
and U21839 (N_21839,N_21006,N_21057);
and U21840 (N_21840,N_21194,N_21351);
xor U21841 (N_21841,N_21162,N_21276);
and U21842 (N_21842,N_21307,N_21012);
or U21843 (N_21843,N_21444,N_21164);
nor U21844 (N_21844,N_21345,N_21534);
xnor U21845 (N_21845,N_21246,N_21089);
nor U21846 (N_21846,N_21305,N_21590);
nor U21847 (N_21847,N_21421,N_21140);
or U21848 (N_21848,N_21195,N_21407);
and U21849 (N_21849,N_21045,N_21262);
nand U21850 (N_21850,N_21139,N_21151);
and U21851 (N_21851,N_21545,N_21283);
xnor U21852 (N_21852,N_21377,N_21272);
nand U21853 (N_21853,N_21580,N_21392);
nor U21854 (N_21854,N_21464,N_21516);
xor U21855 (N_21855,N_21560,N_21506);
or U21856 (N_21856,N_21049,N_21458);
or U21857 (N_21857,N_21202,N_21062);
nand U21858 (N_21858,N_21521,N_21573);
or U21859 (N_21859,N_21370,N_21374);
nand U21860 (N_21860,N_21299,N_21429);
and U21861 (N_21861,N_21319,N_21019);
nand U21862 (N_21862,N_21125,N_21135);
nor U21863 (N_21863,N_21537,N_21358);
or U21864 (N_21864,N_21588,N_21197);
nor U21865 (N_21865,N_21378,N_21067);
xnor U21866 (N_21866,N_21119,N_21427);
or U21867 (N_21867,N_21238,N_21169);
and U21868 (N_21868,N_21386,N_21550);
nor U21869 (N_21869,N_21403,N_21068);
xnor U21870 (N_21870,N_21476,N_21512);
xnor U21871 (N_21871,N_21034,N_21450);
nor U21872 (N_21872,N_21322,N_21048);
nor U21873 (N_21873,N_21024,N_21256);
nor U21874 (N_21874,N_21414,N_21418);
and U21875 (N_21875,N_21419,N_21073);
nor U21876 (N_21876,N_21379,N_21325);
and U21877 (N_21877,N_21359,N_21423);
and U21878 (N_21878,N_21488,N_21388);
and U21879 (N_21879,N_21090,N_21259);
xor U21880 (N_21880,N_21367,N_21509);
and U21881 (N_21881,N_21219,N_21041);
or U21882 (N_21882,N_21190,N_21008);
or U21883 (N_21883,N_21297,N_21577);
nand U21884 (N_21884,N_21353,N_21391);
or U21885 (N_21885,N_21147,N_21042);
and U21886 (N_21886,N_21428,N_21441);
nor U21887 (N_21887,N_21541,N_21323);
and U21888 (N_21888,N_21079,N_21547);
or U21889 (N_21889,N_21368,N_21166);
or U21890 (N_21890,N_21454,N_21009);
nor U21891 (N_21891,N_21530,N_21156);
or U21892 (N_21892,N_21145,N_21507);
nor U21893 (N_21893,N_21583,N_21410);
and U21894 (N_21894,N_21566,N_21100);
nor U21895 (N_21895,N_21220,N_21346);
xor U21896 (N_21896,N_21459,N_21257);
nor U21897 (N_21897,N_21254,N_21446);
or U21898 (N_21898,N_21468,N_21355);
or U21899 (N_21899,N_21328,N_21231);
or U21900 (N_21900,N_21534,N_21375);
or U21901 (N_21901,N_21247,N_21504);
xnor U21902 (N_21902,N_21332,N_21199);
nor U21903 (N_21903,N_21070,N_21503);
xor U21904 (N_21904,N_21222,N_21047);
nand U21905 (N_21905,N_21103,N_21043);
and U21906 (N_21906,N_21140,N_21289);
nand U21907 (N_21907,N_21495,N_21566);
nor U21908 (N_21908,N_21533,N_21439);
nand U21909 (N_21909,N_21253,N_21526);
and U21910 (N_21910,N_21566,N_21460);
nor U21911 (N_21911,N_21515,N_21578);
xor U21912 (N_21912,N_21542,N_21467);
and U21913 (N_21913,N_21315,N_21070);
nor U21914 (N_21914,N_21052,N_21236);
or U21915 (N_21915,N_21366,N_21432);
or U21916 (N_21916,N_21320,N_21232);
or U21917 (N_21917,N_21350,N_21422);
or U21918 (N_21918,N_21207,N_21585);
xnor U21919 (N_21919,N_21138,N_21281);
xnor U21920 (N_21920,N_21470,N_21268);
nor U21921 (N_21921,N_21382,N_21040);
and U21922 (N_21922,N_21245,N_21263);
xor U21923 (N_21923,N_21315,N_21582);
nor U21924 (N_21924,N_21116,N_21052);
nor U21925 (N_21925,N_21482,N_21195);
nand U21926 (N_21926,N_21058,N_21329);
and U21927 (N_21927,N_21469,N_21517);
or U21928 (N_21928,N_21081,N_21052);
nand U21929 (N_21929,N_21174,N_21426);
or U21930 (N_21930,N_21512,N_21184);
or U21931 (N_21931,N_21308,N_21489);
nand U21932 (N_21932,N_21365,N_21306);
and U21933 (N_21933,N_21405,N_21306);
xor U21934 (N_21934,N_21398,N_21167);
xnor U21935 (N_21935,N_21096,N_21055);
and U21936 (N_21936,N_21121,N_21009);
and U21937 (N_21937,N_21065,N_21211);
nor U21938 (N_21938,N_21549,N_21197);
or U21939 (N_21939,N_21002,N_21212);
xor U21940 (N_21940,N_21402,N_21249);
nand U21941 (N_21941,N_21089,N_21327);
and U21942 (N_21942,N_21570,N_21313);
and U21943 (N_21943,N_21491,N_21162);
nor U21944 (N_21944,N_21310,N_21145);
nor U21945 (N_21945,N_21276,N_21272);
or U21946 (N_21946,N_21336,N_21163);
nand U21947 (N_21947,N_21298,N_21212);
nor U21948 (N_21948,N_21480,N_21407);
and U21949 (N_21949,N_21378,N_21107);
nor U21950 (N_21950,N_21235,N_21516);
nand U21951 (N_21951,N_21489,N_21194);
nand U21952 (N_21952,N_21222,N_21456);
nand U21953 (N_21953,N_21337,N_21062);
and U21954 (N_21954,N_21378,N_21227);
and U21955 (N_21955,N_21046,N_21138);
and U21956 (N_21956,N_21031,N_21571);
nor U21957 (N_21957,N_21202,N_21178);
nand U21958 (N_21958,N_21511,N_21475);
nand U21959 (N_21959,N_21085,N_21072);
xnor U21960 (N_21960,N_21244,N_21395);
nand U21961 (N_21961,N_21254,N_21142);
or U21962 (N_21962,N_21530,N_21228);
and U21963 (N_21963,N_21435,N_21584);
xor U21964 (N_21964,N_21000,N_21428);
and U21965 (N_21965,N_21460,N_21130);
nand U21966 (N_21966,N_21301,N_21430);
xor U21967 (N_21967,N_21501,N_21094);
or U21968 (N_21968,N_21217,N_21138);
nand U21969 (N_21969,N_21047,N_21294);
xnor U21970 (N_21970,N_21530,N_21342);
and U21971 (N_21971,N_21044,N_21292);
nand U21972 (N_21972,N_21096,N_21399);
xor U21973 (N_21973,N_21288,N_21252);
or U21974 (N_21974,N_21154,N_21198);
or U21975 (N_21975,N_21084,N_21577);
or U21976 (N_21976,N_21199,N_21274);
nand U21977 (N_21977,N_21198,N_21139);
nor U21978 (N_21978,N_21356,N_21205);
nor U21979 (N_21979,N_21520,N_21564);
or U21980 (N_21980,N_21115,N_21002);
or U21981 (N_21981,N_21002,N_21008);
or U21982 (N_21982,N_21086,N_21080);
xor U21983 (N_21983,N_21542,N_21594);
xor U21984 (N_21984,N_21236,N_21032);
xnor U21985 (N_21985,N_21397,N_21282);
or U21986 (N_21986,N_21184,N_21524);
xor U21987 (N_21987,N_21161,N_21513);
xnor U21988 (N_21988,N_21363,N_21054);
xor U21989 (N_21989,N_21161,N_21470);
xnor U21990 (N_21990,N_21298,N_21418);
xnor U21991 (N_21991,N_21007,N_21344);
or U21992 (N_21992,N_21481,N_21333);
and U21993 (N_21993,N_21343,N_21350);
and U21994 (N_21994,N_21481,N_21518);
xnor U21995 (N_21995,N_21485,N_21168);
nand U21996 (N_21996,N_21478,N_21368);
nor U21997 (N_21997,N_21156,N_21377);
or U21998 (N_21998,N_21472,N_21239);
and U21999 (N_21999,N_21395,N_21454);
and U22000 (N_22000,N_21061,N_21538);
xnor U22001 (N_22001,N_21118,N_21177);
nand U22002 (N_22002,N_21137,N_21494);
and U22003 (N_22003,N_21543,N_21533);
nand U22004 (N_22004,N_21354,N_21417);
and U22005 (N_22005,N_21427,N_21272);
xnor U22006 (N_22006,N_21460,N_21100);
nand U22007 (N_22007,N_21138,N_21490);
or U22008 (N_22008,N_21490,N_21528);
xnor U22009 (N_22009,N_21290,N_21376);
xnor U22010 (N_22010,N_21296,N_21265);
and U22011 (N_22011,N_21348,N_21064);
nand U22012 (N_22012,N_21434,N_21006);
and U22013 (N_22013,N_21544,N_21498);
xnor U22014 (N_22014,N_21508,N_21276);
nor U22015 (N_22015,N_21133,N_21593);
or U22016 (N_22016,N_21302,N_21457);
xor U22017 (N_22017,N_21439,N_21105);
xor U22018 (N_22018,N_21265,N_21056);
or U22019 (N_22019,N_21234,N_21099);
nand U22020 (N_22020,N_21068,N_21168);
nand U22021 (N_22021,N_21336,N_21081);
or U22022 (N_22022,N_21012,N_21086);
or U22023 (N_22023,N_21365,N_21305);
or U22024 (N_22024,N_21246,N_21278);
and U22025 (N_22025,N_21457,N_21551);
xor U22026 (N_22026,N_21219,N_21180);
and U22027 (N_22027,N_21464,N_21195);
or U22028 (N_22028,N_21297,N_21517);
or U22029 (N_22029,N_21596,N_21191);
or U22030 (N_22030,N_21094,N_21288);
and U22031 (N_22031,N_21498,N_21300);
xnor U22032 (N_22032,N_21358,N_21192);
or U22033 (N_22033,N_21108,N_21384);
nand U22034 (N_22034,N_21455,N_21112);
nor U22035 (N_22035,N_21404,N_21092);
nand U22036 (N_22036,N_21054,N_21020);
or U22037 (N_22037,N_21528,N_21111);
or U22038 (N_22038,N_21432,N_21126);
xnor U22039 (N_22039,N_21205,N_21026);
or U22040 (N_22040,N_21454,N_21264);
nand U22041 (N_22041,N_21329,N_21520);
nor U22042 (N_22042,N_21469,N_21588);
nand U22043 (N_22043,N_21354,N_21368);
xor U22044 (N_22044,N_21590,N_21326);
xnor U22045 (N_22045,N_21554,N_21577);
nor U22046 (N_22046,N_21467,N_21587);
nor U22047 (N_22047,N_21168,N_21293);
and U22048 (N_22048,N_21517,N_21565);
nor U22049 (N_22049,N_21397,N_21310);
xnor U22050 (N_22050,N_21243,N_21591);
and U22051 (N_22051,N_21011,N_21558);
and U22052 (N_22052,N_21028,N_21552);
or U22053 (N_22053,N_21117,N_21507);
or U22054 (N_22054,N_21301,N_21598);
xnor U22055 (N_22055,N_21132,N_21559);
xnor U22056 (N_22056,N_21100,N_21445);
nor U22057 (N_22057,N_21052,N_21144);
nand U22058 (N_22058,N_21352,N_21524);
nand U22059 (N_22059,N_21201,N_21384);
and U22060 (N_22060,N_21594,N_21230);
nor U22061 (N_22061,N_21110,N_21472);
and U22062 (N_22062,N_21358,N_21404);
nor U22063 (N_22063,N_21098,N_21094);
or U22064 (N_22064,N_21010,N_21443);
or U22065 (N_22065,N_21474,N_21423);
xnor U22066 (N_22066,N_21246,N_21160);
nand U22067 (N_22067,N_21077,N_21342);
nand U22068 (N_22068,N_21245,N_21495);
nor U22069 (N_22069,N_21168,N_21142);
xnor U22070 (N_22070,N_21101,N_21425);
nor U22071 (N_22071,N_21046,N_21126);
xor U22072 (N_22072,N_21146,N_21428);
nand U22073 (N_22073,N_21253,N_21307);
or U22074 (N_22074,N_21099,N_21476);
nor U22075 (N_22075,N_21269,N_21002);
nor U22076 (N_22076,N_21349,N_21583);
nor U22077 (N_22077,N_21013,N_21388);
and U22078 (N_22078,N_21202,N_21444);
xor U22079 (N_22079,N_21242,N_21259);
nor U22080 (N_22080,N_21267,N_21446);
nor U22081 (N_22081,N_21499,N_21379);
or U22082 (N_22082,N_21520,N_21526);
xor U22083 (N_22083,N_21031,N_21392);
and U22084 (N_22084,N_21567,N_21331);
nor U22085 (N_22085,N_21505,N_21314);
or U22086 (N_22086,N_21165,N_21025);
xnor U22087 (N_22087,N_21131,N_21543);
or U22088 (N_22088,N_21274,N_21186);
nand U22089 (N_22089,N_21283,N_21179);
nor U22090 (N_22090,N_21221,N_21401);
and U22091 (N_22091,N_21380,N_21503);
xnor U22092 (N_22092,N_21055,N_21418);
or U22093 (N_22093,N_21238,N_21162);
nand U22094 (N_22094,N_21483,N_21161);
nand U22095 (N_22095,N_21104,N_21226);
and U22096 (N_22096,N_21229,N_21457);
nand U22097 (N_22097,N_21244,N_21496);
nand U22098 (N_22098,N_21337,N_21048);
nand U22099 (N_22099,N_21540,N_21395);
nand U22100 (N_22100,N_21043,N_21406);
or U22101 (N_22101,N_21192,N_21446);
xnor U22102 (N_22102,N_21147,N_21522);
xnor U22103 (N_22103,N_21582,N_21291);
nor U22104 (N_22104,N_21023,N_21330);
and U22105 (N_22105,N_21022,N_21176);
nand U22106 (N_22106,N_21198,N_21034);
nor U22107 (N_22107,N_21558,N_21083);
nor U22108 (N_22108,N_21211,N_21506);
or U22109 (N_22109,N_21152,N_21108);
or U22110 (N_22110,N_21062,N_21327);
and U22111 (N_22111,N_21433,N_21109);
nor U22112 (N_22112,N_21429,N_21509);
or U22113 (N_22113,N_21105,N_21417);
nand U22114 (N_22114,N_21379,N_21392);
nor U22115 (N_22115,N_21279,N_21303);
nor U22116 (N_22116,N_21439,N_21307);
nor U22117 (N_22117,N_21227,N_21107);
or U22118 (N_22118,N_21019,N_21277);
xnor U22119 (N_22119,N_21334,N_21188);
and U22120 (N_22120,N_21256,N_21569);
nand U22121 (N_22121,N_21276,N_21288);
nor U22122 (N_22122,N_21102,N_21512);
nand U22123 (N_22123,N_21481,N_21455);
nor U22124 (N_22124,N_21117,N_21119);
nor U22125 (N_22125,N_21223,N_21154);
nor U22126 (N_22126,N_21039,N_21090);
nor U22127 (N_22127,N_21357,N_21205);
nand U22128 (N_22128,N_21518,N_21106);
nand U22129 (N_22129,N_21120,N_21090);
nor U22130 (N_22130,N_21122,N_21001);
nand U22131 (N_22131,N_21292,N_21110);
xor U22132 (N_22132,N_21462,N_21092);
and U22133 (N_22133,N_21045,N_21322);
xnor U22134 (N_22134,N_21148,N_21496);
or U22135 (N_22135,N_21455,N_21090);
and U22136 (N_22136,N_21422,N_21202);
xnor U22137 (N_22137,N_21460,N_21590);
xnor U22138 (N_22138,N_21370,N_21016);
nand U22139 (N_22139,N_21411,N_21567);
nand U22140 (N_22140,N_21099,N_21574);
and U22141 (N_22141,N_21591,N_21524);
nand U22142 (N_22142,N_21231,N_21397);
or U22143 (N_22143,N_21227,N_21404);
nand U22144 (N_22144,N_21061,N_21188);
nor U22145 (N_22145,N_21330,N_21222);
or U22146 (N_22146,N_21417,N_21299);
or U22147 (N_22147,N_21260,N_21500);
xnor U22148 (N_22148,N_21547,N_21290);
nand U22149 (N_22149,N_21381,N_21480);
xor U22150 (N_22150,N_21400,N_21524);
and U22151 (N_22151,N_21515,N_21343);
nor U22152 (N_22152,N_21045,N_21237);
and U22153 (N_22153,N_21034,N_21325);
or U22154 (N_22154,N_21297,N_21199);
xnor U22155 (N_22155,N_21045,N_21483);
nand U22156 (N_22156,N_21170,N_21328);
or U22157 (N_22157,N_21315,N_21000);
or U22158 (N_22158,N_21096,N_21003);
nor U22159 (N_22159,N_21498,N_21143);
or U22160 (N_22160,N_21552,N_21339);
or U22161 (N_22161,N_21154,N_21454);
and U22162 (N_22162,N_21027,N_21033);
or U22163 (N_22163,N_21164,N_21513);
xor U22164 (N_22164,N_21031,N_21160);
or U22165 (N_22165,N_21163,N_21246);
or U22166 (N_22166,N_21329,N_21304);
and U22167 (N_22167,N_21367,N_21404);
xnor U22168 (N_22168,N_21280,N_21241);
xor U22169 (N_22169,N_21495,N_21036);
and U22170 (N_22170,N_21256,N_21315);
nand U22171 (N_22171,N_21497,N_21267);
nand U22172 (N_22172,N_21115,N_21263);
or U22173 (N_22173,N_21380,N_21049);
or U22174 (N_22174,N_21513,N_21549);
and U22175 (N_22175,N_21039,N_21323);
nor U22176 (N_22176,N_21069,N_21454);
or U22177 (N_22177,N_21559,N_21042);
nand U22178 (N_22178,N_21106,N_21240);
nand U22179 (N_22179,N_21136,N_21155);
xor U22180 (N_22180,N_21529,N_21138);
or U22181 (N_22181,N_21236,N_21046);
xnor U22182 (N_22182,N_21194,N_21547);
and U22183 (N_22183,N_21228,N_21266);
and U22184 (N_22184,N_21462,N_21406);
nor U22185 (N_22185,N_21127,N_21355);
or U22186 (N_22186,N_21594,N_21251);
xor U22187 (N_22187,N_21470,N_21505);
nand U22188 (N_22188,N_21142,N_21037);
and U22189 (N_22189,N_21015,N_21026);
and U22190 (N_22190,N_21366,N_21474);
xor U22191 (N_22191,N_21131,N_21426);
and U22192 (N_22192,N_21260,N_21186);
nand U22193 (N_22193,N_21326,N_21322);
and U22194 (N_22194,N_21522,N_21123);
nand U22195 (N_22195,N_21040,N_21314);
or U22196 (N_22196,N_21555,N_21208);
and U22197 (N_22197,N_21383,N_21336);
nor U22198 (N_22198,N_21441,N_21580);
xor U22199 (N_22199,N_21460,N_21357);
nor U22200 (N_22200,N_21926,N_21614);
or U22201 (N_22201,N_21935,N_21988);
nor U22202 (N_22202,N_21895,N_21715);
or U22203 (N_22203,N_22003,N_22129);
nand U22204 (N_22204,N_22033,N_21906);
nand U22205 (N_22205,N_21777,N_21620);
or U22206 (N_22206,N_21981,N_21821);
and U22207 (N_22207,N_21698,N_22061);
nand U22208 (N_22208,N_21722,N_21862);
or U22209 (N_22209,N_22029,N_21707);
or U22210 (N_22210,N_22149,N_21986);
nor U22211 (N_22211,N_21946,N_22187);
and U22212 (N_22212,N_21762,N_21867);
xor U22213 (N_22213,N_22116,N_21728);
or U22214 (N_22214,N_21699,N_21887);
xnor U22215 (N_22215,N_21782,N_21880);
xnor U22216 (N_22216,N_21677,N_21802);
nor U22217 (N_22217,N_22125,N_22131);
nand U22218 (N_22218,N_21754,N_22066);
nand U22219 (N_22219,N_21953,N_22106);
and U22220 (N_22220,N_21847,N_21965);
and U22221 (N_22221,N_21818,N_22041);
nor U22222 (N_22222,N_22028,N_21668);
nand U22223 (N_22223,N_21779,N_21774);
xor U22224 (N_22224,N_22088,N_22005);
and U22225 (N_22225,N_21697,N_22161);
or U22226 (N_22226,N_21748,N_22082);
nand U22227 (N_22227,N_21873,N_22002);
nand U22228 (N_22228,N_21914,N_21733);
nor U22229 (N_22229,N_21747,N_22091);
and U22230 (N_22230,N_21934,N_21630);
and U22231 (N_22231,N_21768,N_22193);
or U22232 (N_22232,N_21928,N_21643);
xnor U22233 (N_22233,N_22175,N_21925);
nor U22234 (N_22234,N_21898,N_22067);
xnor U22235 (N_22235,N_22037,N_21827);
and U22236 (N_22236,N_22188,N_21797);
xnor U22237 (N_22237,N_21691,N_22089);
xor U22238 (N_22238,N_21674,N_22045);
nand U22239 (N_22239,N_22031,N_21730);
nand U22240 (N_22240,N_22098,N_22060);
nand U22241 (N_22241,N_21853,N_21949);
and U22242 (N_22242,N_21772,N_21921);
and U22243 (N_22243,N_21684,N_21805);
or U22244 (N_22244,N_21646,N_21750);
xor U22245 (N_22245,N_22073,N_21605);
and U22246 (N_22246,N_22139,N_22077);
or U22247 (N_22247,N_21979,N_21855);
nor U22248 (N_22248,N_21687,N_21900);
or U22249 (N_22249,N_21839,N_21841);
nor U22250 (N_22250,N_22011,N_21823);
xor U22251 (N_22251,N_21929,N_22000);
xor U22252 (N_22252,N_21840,N_21967);
nand U22253 (N_22253,N_21666,N_21692);
and U22254 (N_22254,N_22142,N_21603);
and U22255 (N_22255,N_21924,N_21601);
or U22256 (N_22256,N_22009,N_21792);
and U22257 (N_22257,N_21660,N_21972);
or U22258 (N_22258,N_21901,N_21982);
or U22259 (N_22259,N_21834,N_21765);
xnor U22260 (N_22260,N_21820,N_21703);
xnor U22261 (N_22261,N_21952,N_22013);
or U22262 (N_22262,N_22172,N_22035);
nand U22263 (N_22263,N_22124,N_22148);
nor U22264 (N_22264,N_22113,N_21667);
nor U22265 (N_22265,N_21975,N_21997);
nor U22266 (N_22266,N_21908,N_22117);
xnor U22267 (N_22267,N_22140,N_21623);
xor U22268 (N_22268,N_21916,N_21864);
nor U22269 (N_22269,N_21803,N_21763);
nand U22270 (N_22270,N_22178,N_22155);
or U22271 (N_22271,N_21993,N_22008);
nor U22272 (N_22272,N_21683,N_22166);
nor U22273 (N_22273,N_22136,N_22078);
xor U22274 (N_22274,N_21721,N_22055);
nor U22275 (N_22275,N_21608,N_21959);
or U22276 (N_22276,N_21662,N_21784);
or U22277 (N_22277,N_21848,N_21672);
nor U22278 (N_22278,N_21842,N_21678);
or U22279 (N_22279,N_22093,N_21776);
nand U22280 (N_22280,N_21844,N_21717);
and U22281 (N_22281,N_21770,N_21962);
and U22282 (N_22282,N_21868,N_21710);
xor U22283 (N_22283,N_21689,N_21602);
xor U22284 (N_22284,N_21787,N_21759);
xnor U22285 (N_22285,N_21663,N_22081);
nand U22286 (N_22286,N_21892,N_22165);
nand U22287 (N_22287,N_22063,N_22048);
nor U22288 (N_22288,N_21974,N_21889);
nor U22289 (N_22289,N_22047,N_22177);
xnor U22290 (N_22290,N_21628,N_21830);
xor U22291 (N_22291,N_22100,N_21751);
xnor U22292 (N_22292,N_21738,N_21612);
and U22293 (N_22293,N_21635,N_21884);
nand U22294 (N_22294,N_21822,N_22058);
and U22295 (N_22295,N_21833,N_22097);
or U22296 (N_22296,N_21609,N_21800);
nor U22297 (N_22297,N_21854,N_22176);
or U22298 (N_22298,N_21915,N_21815);
and U22299 (N_22299,N_21980,N_21958);
nand U22300 (N_22300,N_22181,N_21992);
nor U22301 (N_22301,N_21918,N_22171);
xor U22302 (N_22302,N_21955,N_22085);
nand U22303 (N_22303,N_22153,N_21956);
and U22304 (N_22304,N_22065,N_21983);
xnor U22305 (N_22305,N_21969,N_21945);
and U22306 (N_22306,N_21753,N_21865);
and U22307 (N_22307,N_22025,N_21785);
nand U22308 (N_22308,N_21960,N_22105);
or U22309 (N_22309,N_22173,N_22137);
or U22310 (N_22310,N_21659,N_21723);
and U22311 (N_22311,N_21871,N_22084);
or U22312 (N_22312,N_21919,N_22130);
nand U22313 (N_22313,N_21922,N_21883);
or U22314 (N_22314,N_21607,N_21786);
or U22315 (N_22315,N_22074,N_22199);
nor U22316 (N_22316,N_22151,N_21904);
nand U22317 (N_22317,N_21963,N_21936);
and U22318 (N_22318,N_22034,N_21706);
nand U22319 (N_22319,N_21679,N_21651);
xor U22320 (N_22320,N_22032,N_21794);
and U22321 (N_22321,N_21718,N_22007);
xor U22322 (N_22322,N_21888,N_21954);
and U22323 (N_22323,N_22180,N_22051);
and U22324 (N_22324,N_21700,N_21902);
and U22325 (N_22325,N_21645,N_21775);
nand U22326 (N_22326,N_21801,N_21825);
xnor U22327 (N_22327,N_21941,N_21604);
xnor U22328 (N_22328,N_21940,N_21923);
and U22329 (N_22329,N_21727,N_22050);
xnor U22330 (N_22330,N_21615,N_21807);
xnor U22331 (N_22331,N_21633,N_21957);
nand U22332 (N_22332,N_22112,N_21920);
nor U22333 (N_22333,N_21616,N_21882);
or U22334 (N_22334,N_21647,N_22186);
nor U22335 (N_22335,N_21675,N_22184);
xnor U22336 (N_22336,N_22010,N_22030);
nor U22337 (N_22337,N_22160,N_22023);
and U22338 (N_22338,N_21613,N_21907);
nor U22339 (N_22339,N_22185,N_21654);
nand U22340 (N_22340,N_21857,N_22135);
and U22341 (N_22341,N_21746,N_22169);
nor U22342 (N_22342,N_22057,N_21642);
nand U22343 (N_22343,N_22197,N_22121);
xor U22344 (N_22344,N_22126,N_21644);
nand U22345 (N_22345,N_21756,N_22162);
and U22346 (N_22346,N_22134,N_21879);
or U22347 (N_22347,N_22190,N_21944);
or U22348 (N_22348,N_22038,N_21795);
nor U22349 (N_22349,N_21810,N_21851);
or U22350 (N_22350,N_21829,N_21670);
xnor U22351 (N_22351,N_21832,N_22192);
nor U22352 (N_22352,N_21813,N_21849);
nand U22353 (N_22353,N_22120,N_22069);
or U22354 (N_22354,N_21744,N_21896);
and U22355 (N_22355,N_22090,N_21806);
and U22356 (N_22356,N_21716,N_22059);
nand U22357 (N_22357,N_21638,N_21826);
or U22358 (N_22358,N_21653,N_21652);
nand U22359 (N_22359,N_22016,N_21790);
xnor U22360 (N_22360,N_21942,N_21690);
nor U22361 (N_22361,N_21617,N_22092);
nand U22362 (N_22362,N_22159,N_21863);
and U22363 (N_22363,N_22118,N_21874);
xnor U22364 (N_22364,N_22094,N_21640);
nor U22365 (N_22365,N_22146,N_21637);
nand U22366 (N_22366,N_21655,N_22123);
or U22367 (N_22367,N_21626,N_21927);
nor U22368 (N_22368,N_21636,N_21869);
and U22369 (N_22369,N_21724,N_21816);
nand U22370 (N_22370,N_22052,N_21973);
xor U22371 (N_22371,N_21950,N_21791);
and U22372 (N_22372,N_21618,N_21930);
or U22373 (N_22373,N_22167,N_21860);
nand U22374 (N_22374,N_22145,N_22099);
and U22375 (N_22375,N_21976,N_21769);
and U22376 (N_22376,N_21758,N_21704);
nor U22377 (N_22377,N_21948,N_21725);
nor U22378 (N_22378,N_21872,N_22143);
xor U22379 (N_22379,N_21611,N_21814);
nand U22380 (N_22380,N_21743,N_22019);
and U22381 (N_22381,N_21767,N_21843);
or U22382 (N_22382,N_21964,N_22021);
or U22383 (N_22383,N_21755,N_21891);
nand U22384 (N_22384,N_21624,N_21682);
xor U22385 (N_22385,N_21729,N_22179);
nor U22386 (N_22386,N_21994,N_21987);
xor U22387 (N_22387,N_21828,N_21903);
xor U22388 (N_22388,N_22068,N_21951);
or U22389 (N_22389,N_21665,N_21621);
nor U22390 (N_22390,N_22182,N_22012);
nor U22391 (N_22391,N_22056,N_21991);
or U22392 (N_22392,N_22147,N_22018);
and U22393 (N_22393,N_21913,N_22087);
nand U22394 (N_22394,N_21966,N_22006);
or U22395 (N_22395,N_21600,N_21701);
or U22396 (N_22396,N_22141,N_22070);
nand U22397 (N_22397,N_22086,N_21773);
nand U22398 (N_22398,N_22158,N_21749);
and U22399 (N_22399,N_21796,N_21938);
or U22400 (N_22400,N_21629,N_21737);
and U22401 (N_22401,N_21745,N_22128);
or U22402 (N_22402,N_21676,N_21757);
nand U22403 (N_22403,N_21837,N_21661);
nor U22404 (N_22404,N_21793,N_21998);
and U22405 (N_22405,N_21671,N_21894);
nand U22406 (N_22406,N_21720,N_21876);
or U22407 (N_22407,N_21788,N_22163);
or U22408 (N_22408,N_22022,N_21978);
xnor U22409 (N_22409,N_21760,N_21911);
nor U22410 (N_22410,N_22049,N_22154);
xnor U22411 (N_22411,N_21870,N_21852);
nor U22412 (N_22412,N_21824,N_22191);
or U22413 (N_22413,N_22119,N_21783);
nor U22414 (N_22414,N_21649,N_22075);
nand U22415 (N_22415,N_21685,N_21752);
and U22416 (N_22416,N_21968,N_21713);
nand U22417 (N_22417,N_22001,N_21632);
nor U22418 (N_22418,N_21910,N_21702);
xnor U22419 (N_22419,N_22042,N_21719);
nand U22420 (N_22420,N_21648,N_21836);
and U22421 (N_22421,N_21917,N_21688);
or U22422 (N_22422,N_21859,N_21669);
xnor U22423 (N_22423,N_22024,N_22101);
and U22424 (N_22424,N_21939,N_21912);
nand U22425 (N_22425,N_21711,N_21861);
nor U22426 (N_22426,N_21850,N_22095);
xor U22427 (N_22427,N_21695,N_21778);
nand U22428 (N_22428,N_22168,N_21804);
nor U22429 (N_22429,N_22072,N_21947);
nand U22430 (N_22430,N_21789,N_21764);
nor U22431 (N_22431,N_22027,N_21932);
or U22432 (N_22432,N_21606,N_21634);
xnor U22433 (N_22433,N_22015,N_22144);
nand U22434 (N_22434,N_22053,N_22039);
or U22435 (N_22435,N_22109,N_22046);
xnor U22436 (N_22436,N_21893,N_21627);
or U22437 (N_22437,N_22189,N_22103);
xor U22438 (N_22438,N_22036,N_21735);
or U22439 (N_22439,N_21809,N_21656);
xnor U22440 (N_22440,N_22110,N_21819);
or U22441 (N_22441,N_22071,N_22083);
nor U22442 (N_22442,N_21781,N_22026);
xnor U22443 (N_22443,N_21989,N_21657);
nand U22444 (N_22444,N_21708,N_21937);
or U22445 (N_22445,N_21881,N_22014);
and U22446 (N_22446,N_21984,N_21712);
and U22447 (N_22447,N_22064,N_21905);
or U22448 (N_22448,N_22198,N_22107);
or U22449 (N_22449,N_22127,N_21875);
or U22450 (N_22450,N_21846,N_21961);
nor U22451 (N_22451,N_21639,N_21996);
nor U22452 (N_22452,N_21845,N_21766);
or U22453 (N_22453,N_21714,N_21886);
nand U22454 (N_22454,N_21705,N_21890);
xor U22455 (N_22455,N_22108,N_22133);
nand U22456 (N_22456,N_21970,N_22156);
or U22457 (N_22457,N_21625,N_22196);
or U22458 (N_22458,N_22132,N_21971);
xnor U22459 (N_22459,N_21641,N_21771);
xnor U22460 (N_22460,N_22080,N_21866);
xor U22461 (N_22461,N_22020,N_22122);
nand U22462 (N_22462,N_21878,N_21736);
or U22463 (N_22463,N_21985,N_21739);
nand U22464 (N_22464,N_21799,N_22170);
nor U22465 (N_22465,N_21798,N_21856);
xnor U22466 (N_22466,N_21693,N_22104);
and U22467 (N_22467,N_21619,N_21694);
and U22468 (N_22468,N_22138,N_21817);
and U22469 (N_22469,N_21990,N_22079);
nand U22470 (N_22470,N_21999,N_21977);
xnor U22471 (N_22471,N_21831,N_21780);
xor U22472 (N_22472,N_22157,N_21885);
nor U22473 (N_22473,N_21933,N_21658);
xnor U22474 (N_22474,N_21811,N_21622);
xor U22475 (N_22475,N_22174,N_22043);
nand U22476 (N_22476,N_22062,N_21899);
or U22477 (N_22477,N_21631,N_21858);
or U22478 (N_22478,N_22017,N_21995);
xor U22479 (N_22479,N_21610,N_21732);
xor U22480 (N_22480,N_21812,N_21835);
and U22481 (N_22481,N_21709,N_21696);
nand U22482 (N_22482,N_21931,N_22114);
nand U22483 (N_22483,N_22195,N_22040);
and U22484 (N_22484,N_21838,N_21731);
nor U22485 (N_22485,N_21808,N_21943);
nor U22486 (N_22486,N_22115,N_21761);
nand U22487 (N_22487,N_21897,N_22102);
nand U22488 (N_22488,N_22096,N_21877);
nand U22489 (N_22489,N_21681,N_21726);
nand U22490 (N_22490,N_22164,N_21673);
xor U22491 (N_22491,N_22111,N_21686);
nor U22492 (N_22492,N_21650,N_22150);
or U22493 (N_22493,N_21734,N_21664);
or U22494 (N_22494,N_22194,N_22183);
or U22495 (N_22495,N_22076,N_21680);
nor U22496 (N_22496,N_21740,N_22152);
nand U22497 (N_22497,N_22044,N_22054);
nand U22498 (N_22498,N_21741,N_21909);
nor U22499 (N_22499,N_21742,N_22004);
and U22500 (N_22500,N_21828,N_21627);
and U22501 (N_22501,N_22074,N_21671);
and U22502 (N_22502,N_22152,N_21680);
nor U22503 (N_22503,N_21913,N_22089);
or U22504 (N_22504,N_21699,N_22014);
xnor U22505 (N_22505,N_21609,N_22112);
xor U22506 (N_22506,N_22132,N_21876);
xor U22507 (N_22507,N_21975,N_21907);
or U22508 (N_22508,N_21611,N_21612);
nor U22509 (N_22509,N_22139,N_22081);
and U22510 (N_22510,N_21951,N_22018);
or U22511 (N_22511,N_22091,N_21685);
nand U22512 (N_22512,N_21880,N_21930);
or U22513 (N_22513,N_21677,N_21682);
xor U22514 (N_22514,N_21943,N_22193);
xnor U22515 (N_22515,N_21726,N_21898);
or U22516 (N_22516,N_21616,N_21636);
xor U22517 (N_22517,N_21935,N_21861);
or U22518 (N_22518,N_22084,N_21602);
and U22519 (N_22519,N_22039,N_21928);
xor U22520 (N_22520,N_21604,N_21798);
nor U22521 (N_22521,N_21957,N_21832);
xor U22522 (N_22522,N_21855,N_22031);
nor U22523 (N_22523,N_21650,N_21749);
nand U22524 (N_22524,N_21960,N_22143);
nand U22525 (N_22525,N_21688,N_21641);
or U22526 (N_22526,N_21664,N_22149);
xor U22527 (N_22527,N_22087,N_21801);
and U22528 (N_22528,N_21959,N_22116);
or U22529 (N_22529,N_22061,N_21894);
nand U22530 (N_22530,N_22009,N_21797);
xor U22531 (N_22531,N_21891,N_21761);
nand U22532 (N_22532,N_21770,N_22125);
nor U22533 (N_22533,N_21701,N_21634);
nor U22534 (N_22534,N_21751,N_21691);
nand U22535 (N_22535,N_21662,N_22044);
xor U22536 (N_22536,N_21659,N_21995);
xnor U22537 (N_22537,N_21698,N_21616);
xnor U22538 (N_22538,N_22035,N_22100);
xnor U22539 (N_22539,N_21639,N_22102);
or U22540 (N_22540,N_22086,N_21792);
nand U22541 (N_22541,N_21704,N_21970);
nand U22542 (N_22542,N_21929,N_22176);
nand U22543 (N_22543,N_22070,N_21739);
nand U22544 (N_22544,N_21717,N_21835);
and U22545 (N_22545,N_21997,N_22161);
xnor U22546 (N_22546,N_21952,N_21651);
and U22547 (N_22547,N_21721,N_21846);
and U22548 (N_22548,N_22007,N_21617);
xor U22549 (N_22549,N_22154,N_21828);
or U22550 (N_22550,N_22053,N_21665);
xor U22551 (N_22551,N_22159,N_22024);
and U22552 (N_22552,N_21849,N_21647);
nand U22553 (N_22553,N_22009,N_21677);
xor U22554 (N_22554,N_22029,N_21633);
nand U22555 (N_22555,N_22141,N_21693);
xor U22556 (N_22556,N_22125,N_22157);
or U22557 (N_22557,N_21972,N_22078);
xor U22558 (N_22558,N_22148,N_21615);
nor U22559 (N_22559,N_21659,N_22184);
nor U22560 (N_22560,N_22096,N_21977);
or U22561 (N_22561,N_22039,N_21850);
xor U22562 (N_22562,N_22196,N_21985);
and U22563 (N_22563,N_22045,N_22035);
nor U22564 (N_22564,N_21955,N_21725);
nor U22565 (N_22565,N_21737,N_22196);
and U22566 (N_22566,N_22072,N_21762);
nor U22567 (N_22567,N_21859,N_22046);
or U22568 (N_22568,N_21944,N_21733);
nor U22569 (N_22569,N_21820,N_21866);
or U22570 (N_22570,N_21983,N_22110);
xor U22571 (N_22571,N_22199,N_22172);
and U22572 (N_22572,N_21753,N_21905);
or U22573 (N_22573,N_21983,N_21938);
or U22574 (N_22574,N_21648,N_21976);
or U22575 (N_22575,N_21731,N_22090);
xnor U22576 (N_22576,N_22158,N_22077);
or U22577 (N_22577,N_22072,N_21911);
or U22578 (N_22578,N_21943,N_22086);
nor U22579 (N_22579,N_22049,N_21913);
nor U22580 (N_22580,N_22182,N_21867);
nand U22581 (N_22581,N_22192,N_22076);
or U22582 (N_22582,N_21808,N_22063);
and U22583 (N_22583,N_21941,N_21961);
nor U22584 (N_22584,N_22019,N_22064);
or U22585 (N_22585,N_21618,N_21633);
or U22586 (N_22586,N_22080,N_22016);
and U22587 (N_22587,N_21947,N_21812);
nand U22588 (N_22588,N_21958,N_21867);
or U22589 (N_22589,N_21934,N_21892);
xor U22590 (N_22590,N_21869,N_22137);
and U22591 (N_22591,N_22068,N_21945);
and U22592 (N_22592,N_21785,N_21628);
xor U22593 (N_22593,N_21996,N_21871);
nor U22594 (N_22594,N_21848,N_21746);
and U22595 (N_22595,N_22038,N_22177);
nand U22596 (N_22596,N_21610,N_21660);
and U22597 (N_22597,N_21629,N_21703);
nand U22598 (N_22598,N_22152,N_22009);
or U22599 (N_22599,N_21878,N_21620);
or U22600 (N_22600,N_21837,N_21992);
and U22601 (N_22601,N_21600,N_22180);
xor U22602 (N_22602,N_21912,N_21955);
xor U22603 (N_22603,N_21608,N_22129);
xnor U22604 (N_22604,N_22052,N_22012);
nor U22605 (N_22605,N_21969,N_21979);
nand U22606 (N_22606,N_22059,N_21974);
and U22607 (N_22607,N_21959,N_22174);
nor U22608 (N_22608,N_21641,N_21887);
nand U22609 (N_22609,N_21819,N_21687);
nor U22610 (N_22610,N_22043,N_21923);
xor U22611 (N_22611,N_22067,N_21862);
and U22612 (N_22612,N_21869,N_22174);
or U22613 (N_22613,N_21673,N_21933);
nand U22614 (N_22614,N_21942,N_21892);
xor U22615 (N_22615,N_22009,N_21943);
and U22616 (N_22616,N_22087,N_21709);
and U22617 (N_22617,N_21748,N_21610);
xnor U22618 (N_22618,N_21608,N_21943);
and U22619 (N_22619,N_22186,N_22055);
nand U22620 (N_22620,N_21644,N_22087);
or U22621 (N_22621,N_22152,N_22085);
nand U22622 (N_22622,N_21643,N_21934);
or U22623 (N_22623,N_21663,N_22169);
xor U22624 (N_22624,N_21818,N_21738);
and U22625 (N_22625,N_21674,N_22071);
nand U22626 (N_22626,N_22159,N_21679);
or U22627 (N_22627,N_22052,N_21786);
or U22628 (N_22628,N_21699,N_21769);
xnor U22629 (N_22629,N_21830,N_21707);
nor U22630 (N_22630,N_22146,N_21654);
and U22631 (N_22631,N_21743,N_21765);
xnor U22632 (N_22632,N_21666,N_21935);
nor U22633 (N_22633,N_22011,N_21730);
xor U22634 (N_22634,N_22139,N_21893);
and U22635 (N_22635,N_22047,N_21662);
nand U22636 (N_22636,N_21975,N_21845);
or U22637 (N_22637,N_22095,N_22006);
xnor U22638 (N_22638,N_22186,N_21794);
or U22639 (N_22639,N_22059,N_22162);
nor U22640 (N_22640,N_21849,N_21841);
xor U22641 (N_22641,N_21643,N_22144);
nor U22642 (N_22642,N_21600,N_21843);
nand U22643 (N_22643,N_22010,N_21864);
nand U22644 (N_22644,N_22095,N_21838);
and U22645 (N_22645,N_21996,N_21817);
nor U22646 (N_22646,N_21737,N_21846);
xnor U22647 (N_22647,N_21890,N_22123);
nor U22648 (N_22648,N_21670,N_21873);
xnor U22649 (N_22649,N_21762,N_22162);
or U22650 (N_22650,N_22028,N_22007);
and U22651 (N_22651,N_21903,N_22015);
xnor U22652 (N_22652,N_22090,N_22147);
nor U22653 (N_22653,N_21951,N_22110);
and U22654 (N_22654,N_21766,N_21811);
and U22655 (N_22655,N_21697,N_21768);
xor U22656 (N_22656,N_21743,N_21963);
nand U22657 (N_22657,N_22121,N_21928);
or U22658 (N_22658,N_22160,N_21701);
nand U22659 (N_22659,N_22049,N_22115);
xor U22660 (N_22660,N_21659,N_22113);
nand U22661 (N_22661,N_22173,N_22181);
nand U22662 (N_22662,N_21616,N_21905);
and U22663 (N_22663,N_21863,N_21704);
and U22664 (N_22664,N_21979,N_21835);
or U22665 (N_22665,N_22187,N_22076);
xor U22666 (N_22666,N_21750,N_21888);
nor U22667 (N_22667,N_21869,N_21799);
xor U22668 (N_22668,N_21763,N_21950);
or U22669 (N_22669,N_22055,N_21874);
nor U22670 (N_22670,N_21740,N_21921);
xor U22671 (N_22671,N_21669,N_21992);
and U22672 (N_22672,N_22106,N_21976);
and U22673 (N_22673,N_21702,N_21988);
or U22674 (N_22674,N_21646,N_21979);
xnor U22675 (N_22675,N_22149,N_21660);
and U22676 (N_22676,N_22121,N_22183);
xnor U22677 (N_22677,N_21662,N_21682);
and U22678 (N_22678,N_21892,N_21742);
xnor U22679 (N_22679,N_22089,N_21981);
and U22680 (N_22680,N_21925,N_21711);
and U22681 (N_22681,N_22100,N_22070);
nor U22682 (N_22682,N_21885,N_22068);
nand U22683 (N_22683,N_22031,N_21668);
or U22684 (N_22684,N_21857,N_21716);
nand U22685 (N_22685,N_21716,N_21751);
or U22686 (N_22686,N_22017,N_21960);
and U22687 (N_22687,N_21758,N_22031);
or U22688 (N_22688,N_21745,N_22139);
and U22689 (N_22689,N_21846,N_21735);
and U22690 (N_22690,N_21703,N_21638);
xnor U22691 (N_22691,N_21815,N_21606);
nor U22692 (N_22692,N_21885,N_21839);
xor U22693 (N_22693,N_22161,N_21970);
nor U22694 (N_22694,N_21735,N_22148);
xor U22695 (N_22695,N_21668,N_21708);
nand U22696 (N_22696,N_22163,N_21985);
and U22697 (N_22697,N_21780,N_21980);
nor U22698 (N_22698,N_21674,N_21730);
nor U22699 (N_22699,N_21847,N_22041);
nand U22700 (N_22700,N_21826,N_21847);
and U22701 (N_22701,N_21746,N_21654);
nor U22702 (N_22702,N_21660,N_22162);
and U22703 (N_22703,N_21732,N_21658);
and U22704 (N_22704,N_21862,N_21741);
and U22705 (N_22705,N_22088,N_21893);
and U22706 (N_22706,N_21686,N_22030);
xnor U22707 (N_22707,N_21648,N_21801);
nand U22708 (N_22708,N_22161,N_22022);
and U22709 (N_22709,N_22056,N_21633);
xor U22710 (N_22710,N_21782,N_21739);
xnor U22711 (N_22711,N_21910,N_21949);
nor U22712 (N_22712,N_22047,N_22075);
xor U22713 (N_22713,N_22097,N_21988);
and U22714 (N_22714,N_21695,N_21961);
nor U22715 (N_22715,N_21816,N_22136);
nand U22716 (N_22716,N_21742,N_21800);
or U22717 (N_22717,N_21867,N_21712);
xnor U22718 (N_22718,N_21929,N_21688);
nand U22719 (N_22719,N_21996,N_21902);
nand U22720 (N_22720,N_21849,N_21672);
or U22721 (N_22721,N_21854,N_22115);
xor U22722 (N_22722,N_21766,N_21853);
or U22723 (N_22723,N_22039,N_22153);
or U22724 (N_22724,N_21779,N_21998);
nand U22725 (N_22725,N_21989,N_21739);
and U22726 (N_22726,N_21811,N_21853);
nand U22727 (N_22727,N_21625,N_21828);
nor U22728 (N_22728,N_21721,N_22091);
xor U22729 (N_22729,N_21719,N_21912);
nor U22730 (N_22730,N_22012,N_21905);
nor U22731 (N_22731,N_21851,N_21994);
or U22732 (N_22732,N_21875,N_21637);
or U22733 (N_22733,N_21617,N_21686);
or U22734 (N_22734,N_22028,N_21955);
xnor U22735 (N_22735,N_21833,N_22100);
nand U22736 (N_22736,N_22027,N_22160);
nand U22737 (N_22737,N_21945,N_21637);
xnor U22738 (N_22738,N_21696,N_21909);
xnor U22739 (N_22739,N_21952,N_21763);
nand U22740 (N_22740,N_22081,N_22158);
xnor U22741 (N_22741,N_21946,N_21984);
and U22742 (N_22742,N_21732,N_21628);
xnor U22743 (N_22743,N_21850,N_22143);
and U22744 (N_22744,N_21755,N_22029);
nor U22745 (N_22745,N_22068,N_22144);
xor U22746 (N_22746,N_22147,N_22057);
xor U22747 (N_22747,N_21873,N_22177);
or U22748 (N_22748,N_22111,N_22094);
and U22749 (N_22749,N_22165,N_22029);
xnor U22750 (N_22750,N_21766,N_21836);
xnor U22751 (N_22751,N_21735,N_21766);
nor U22752 (N_22752,N_22094,N_21646);
or U22753 (N_22753,N_21686,N_21833);
nor U22754 (N_22754,N_21985,N_22164);
or U22755 (N_22755,N_22183,N_21846);
nand U22756 (N_22756,N_21711,N_22125);
or U22757 (N_22757,N_22148,N_22066);
nor U22758 (N_22758,N_21887,N_21974);
or U22759 (N_22759,N_22054,N_21744);
and U22760 (N_22760,N_21634,N_22174);
nor U22761 (N_22761,N_21936,N_21851);
nor U22762 (N_22762,N_21957,N_22027);
nor U22763 (N_22763,N_22179,N_21847);
xnor U22764 (N_22764,N_21633,N_21958);
xor U22765 (N_22765,N_22073,N_21736);
nand U22766 (N_22766,N_21868,N_22032);
or U22767 (N_22767,N_22046,N_21643);
or U22768 (N_22768,N_21784,N_22073);
xor U22769 (N_22769,N_22121,N_21987);
nand U22770 (N_22770,N_21737,N_21714);
nand U22771 (N_22771,N_22146,N_21839);
xor U22772 (N_22772,N_21948,N_22036);
and U22773 (N_22773,N_22031,N_21983);
or U22774 (N_22774,N_22104,N_21717);
or U22775 (N_22775,N_21664,N_22044);
nand U22776 (N_22776,N_21758,N_21832);
xnor U22777 (N_22777,N_22013,N_22111);
xor U22778 (N_22778,N_21786,N_21835);
nand U22779 (N_22779,N_22031,N_21728);
nand U22780 (N_22780,N_22181,N_21712);
nand U22781 (N_22781,N_21776,N_22135);
nor U22782 (N_22782,N_21983,N_21849);
and U22783 (N_22783,N_21987,N_21997);
or U22784 (N_22784,N_21709,N_22188);
xnor U22785 (N_22785,N_21622,N_21824);
nand U22786 (N_22786,N_22131,N_22087);
and U22787 (N_22787,N_21648,N_21652);
nand U22788 (N_22788,N_21784,N_21777);
nand U22789 (N_22789,N_22124,N_21788);
and U22790 (N_22790,N_22091,N_21945);
and U22791 (N_22791,N_21971,N_21665);
nor U22792 (N_22792,N_22017,N_21752);
and U22793 (N_22793,N_21957,N_21635);
xor U22794 (N_22794,N_21965,N_21827);
nor U22795 (N_22795,N_22157,N_22104);
xnor U22796 (N_22796,N_21993,N_21928);
xnor U22797 (N_22797,N_21636,N_21879);
xor U22798 (N_22798,N_22147,N_21636);
or U22799 (N_22799,N_21950,N_21896);
and U22800 (N_22800,N_22558,N_22651);
or U22801 (N_22801,N_22754,N_22676);
or U22802 (N_22802,N_22387,N_22697);
xnor U22803 (N_22803,N_22493,N_22263);
or U22804 (N_22804,N_22535,N_22637);
nor U22805 (N_22805,N_22518,N_22729);
or U22806 (N_22806,N_22526,N_22704);
and U22807 (N_22807,N_22600,N_22582);
xor U22808 (N_22808,N_22415,N_22723);
nand U22809 (N_22809,N_22601,N_22540);
or U22810 (N_22810,N_22780,N_22332);
or U22811 (N_22811,N_22334,N_22798);
nand U22812 (N_22812,N_22236,N_22421);
xnor U22813 (N_22813,N_22519,N_22251);
nand U22814 (N_22814,N_22219,N_22490);
nor U22815 (N_22815,N_22442,N_22777);
or U22816 (N_22816,N_22364,N_22668);
nor U22817 (N_22817,N_22650,N_22209);
xor U22818 (N_22818,N_22370,N_22583);
xnor U22819 (N_22819,N_22311,N_22769);
or U22820 (N_22820,N_22397,N_22683);
or U22821 (N_22821,N_22680,N_22521);
xnor U22822 (N_22822,N_22720,N_22572);
nor U22823 (N_22823,N_22256,N_22294);
nor U22824 (N_22824,N_22630,N_22214);
or U22825 (N_22825,N_22770,N_22455);
nand U22826 (N_22826,N_22302,N_22606);
and U22827 (N_22827,N_22344,N_22288);
xor U22828 (N_22828,N_22785,N_22789);
nand U22829 (N_22829,N_22226,N_22329);
xnor U22830 (N_22830,N_22552,N_22274);
xor U22831 (N_22831,N_22466,N_22475);
nand U22832 (N_22832,N_22750,N_22459);
nand U22833 (N_22833,N_22452,N_22632);
nand U22834 (N_22834,N_22391,N_22618);
and U22835 (N_22835,N_22756,N_22372);
and U22836 (N_22836,N_22774,N_22746);
or U22837 (N_22837,N_22677,N_22402);
or U22838 (N_22838,N_22545,N_22661);
and U22839 (N_22839,N_22347,N_22762);
nand U22840 (N_22840,N_22793,N_22299);
nand U22841 (N_22841,N_22380,N_22222);
and U22842 (N_22842,N_22679,N_22759);
and U22843 (N_22843,N_22427,N_22355);
xor U22844 (N_22844,N_22666,N_22373);
or U22845 (N_22845,N_22237,N_22597);
and U22846 (N_22846,N_22654,N_22547);
nor U22847 (N_22847,N_22553,N_22571);
or U22848 (N_22848,N_22505,N_22625);
nand U22849 (N_22849,N_22724,N_22691);
xnor U22850 (N_22850,N_22439,N_22333);
or U22851 (N_22851,N_22736,N_22586);
nand U22852 (N_22852,N_22574,N_22531);
and U22853 (N_22853,N_22737,N_22282);
xnor U22854 (N_22854,N_22779,N_22730);
and U22855 (N_22855,N_22690,N_22412);
nor U22856 (N_22856,N_22658,N_22563);
nor U22857 (N_22857,N_22783,N_22242);
xnor U22858 (N_22858,N_22568,N_22522);
or U22859 (N_22859,N_22223,N_22634);
nand U22860 (N_22860,N_22417,N_22491);
xor U22861 (N_22861,N_22575,N_22570);
xor U22862 (N_22862,N_22515,N_22554);
nor U22863 (N_22863,N_22749,N_22233);
or U22864 (N_22864,N_22734,N_22566);
xor U22865 (N_22865,N_22394,N_22318);
nor U22866 (N_22866,N_22351,N_22349);
nand U22867 (N_22867,N_22411,N_22556);
nand U22868 (N_22868,N_22482,N_22492);
nor U22869 (N_22869,N_22249,N_22213);
nor U22870 (N_22870,N_22216,N_22671);
xor U22871 (N_22871,N_22315,N_22792);
or U22872 (N_22872,N_22448,N_22511);
nand U22873 (N_22873,N_22660,N_22706);
and U22874 (N_22874,N_22748,N_22420);
nand U22875 (N_22875,N_22592,N_22794);
nor U22876 (N_22876,N_22323,N_22278);
xnor U22877 (N_22877,N_22498,N_22569);
nor U22878 (N_22878,N_22424,N_22524);
xor U22879 (N_22879,N_22395,N_22584);
nor U22880 (N_22880,N_22356,N_22434);
nand U22881 (N_22881,N_22445,N_22509);
nor U22882 (N_22882,N_22639,N_22207);
or U22883 (N_22883,N_22670,N_22437);
and U22884 (N_22884,N_22663,N_22450);
and U22885 (N_22885,N_22306,N_22483);
and U22886 (N_22886,N_22408,N_22230);
nor U22887 (N_22887,N_22290,N_22324);
nand U22888 (N_22888,N_22773,N_22285);
xor U22889 (N_22889,N_22376,N_22458);
nor U22890 (N_22890,N_22354,N_22353);
and U22891 (N_22891,N_22687,N_22407);
nand U22892 (N_22892,N_22782,N_22738);
nand U22893 (N_22893,N_22365,N_22751);
and U22894 (N_22894,N_22537,N_22453);
nor U22895 (N_22895,N_22539,N_22550);
nand U22896 (N_22896,N_22447,N_22357);
or U22897 (N_22897,N_22238,N_22594);
nor U22898 (N_22898,N_22390,N_22465);
xnor U22899 (N_22899,N_22396,N_22562);
nor U22900 (N_22900,N_22722,N_22284);
nand U22901 (N_22901,N_22352,N_22588);
and U22902 (N_22902,N_22747,N_22406);
nand U22903 (N_22903,N_22293,N_22405);
and U22904 (N_22904,N_22457,N_22462);
nand U22905 (N_22905,N_22438,N_22719);
or U22906 (N_22906,N_22673,N_22638);
or U22907 (N_22907,N_22693,N_22217);
and U22908 (N_22908,N_22441,N_22507);
or U22909 (N_22909,N_22319,N_22525);
nand U22910 (N_22910,N_22786,N_22460);
and U22911 (N_22911,N_22346,N_22327);
nand U22912 (N_22912,N_22231,N_22205);
nand U22913 (N_22913,N_22435,N_22454);
xnor U22914 (N_22914,N_22361,N_22321);
xor U22915 (N_22915,N_22212,N_22326);
xor U22916 (N_22916,N_22300,N_22422);
nor U22917 (N_22917,N_22423,N_22227);
xor U22918 (N_22918,N_22520,N_22768);
nand U22919 (N_22919,N_22610,N_22655);
xor U22920 (N_22920,N_22781,N_22613);
nand U22921 (N_22921,N_22757,N_22771);
nand U22922 (N_22922,N_22481,N_22579);
or U22923 (N_22923,N_22631,N_22725);
nand U22924 (N_22924,N_22739,N_22265);
xnor U22925 (N_22925,N_22331,N_22640);
nor U22926 (N_22926,N_22210,N_22425);
or U22927 (N_22927,N_22716,N_22418);
nand U22928 (N_22928,N_22612,N_22262);
and U22929 (N_22929,N_22476,N_22644);
nor U22930 (N_22930,N_22449,N_22692);
and U22931 (N_22931,N_22292,N_22268);
or U22932 (N_22932,N_22267,N_22731);
or U22933 (N_22933,N_22776,N_22752);
or U22934 (N_22934,N_22338,N_22627);
or U22935 (N_22935,N_22527,N_22500);
nor U22936 (N_22936,N_22487,N_22416);
nand U22937 (N_22937,N_22528,N_22443);
or U22938 (N_22938,N_22617,N_22385);
nor U22939 (N_22939,N_22204,N_22201);
and U22940 (N_22940,N_22772,N_22686);
xnor U22941 (N_22941,N_22494,N_22790);
nand U22942 (N_22942,N_22477,N_22514);
xnor U22943 (N_22943,N_22733,N_22712);
xor U22944 (N_22944,N_22430,N_22513);
nand U22945 (N_22945,N_22480,N_22283);
nor U22946 (N_22946,N_22542,N_22348);
nand U22947 (N_22947,N_22279,N_22208);
or U22948 (N_22948,N_22440,N_22598);
nor U22949 (N_22949,N_22456,N_22512);
nand U22950 (N_22950,N_22665,N_22382);
nand U22951 (N_22951,N_22523,N_22314);
or U22952 (N_22952,N_22399,N_22471);
xnor U22953 (N_22953,N_22544,N_22576);
nand U22954 (N_22954,N_22694,N_22765);
and U22955 (N_22955,N_22255,N_22428);
nor U22956 (N_22956,N_22474,N_22605);
or U22957 (N_22957,N_22797,N_22296);
and U22958 (N_22958,N_22591,N_22247);
nand U22959 (N_22959,N_22698,N_22799);
nor U22960 (N_22960,N_22564,N_22715);
xnor U22961 (N_22961,N_22745,N_22495);
nor U22962 (N_22962,N_22224,N_22383);
xor U22963 (N_22963,N_22473,N_22414);
xor U22964 (N_22964,N_22656,N_22662);
nand U22965 (N_22965,N_22360,N_22497);
and U22966 (N_22966,N_22620,N_22534);
nand U22967 (N_22967,N_22758,N_22270);
nand U22968 (N_22968,N_22567,N_22275);
xor U22969 (N_22969,N_22499,N_22375);
xnor U22970 (N_22970,N_22257,N_22635);
xnor U22971 (N_22971,N_22404,N_22225);
nand U22972 (N_22972,N_22289,N_22379);
xnor U22973 (N_22973,N_22695,N_22280);
xor U22974 (N_22974,N_22510,N_22621);
and U22975 (N_22975,N_22727,N_22767);
xnor U22976 (N_22976,N_22429,N_22221);
nand U22977 (N_22977,N_22489,N_22235);
and U22978 (N_22978,N_22766,N_22358);
or U22979 (N_22979,N_22641,N_22599);
nor U22980 (N_22980,N_22726,N_22272);
or U22981 (N_22981,N_22503,N_22464);
nand U22982 (N_22982,N_22202,N_22517);
xnor U22983 (N_22983,N_22787,N_22316);
xnor U22984 (N_22984,N_22363,N_22269);
nor U22985 (N_22985,N_22342,N_22744);
xor U22986 (N_22986,N_22384,N_22260);
nand U22987 (N_22987,N_22502,N_22273);
or U22988 (N_22988,N_22451,N_22614);
nor U22989 (N_22989,N_22532,N_22378);
nand U22990 (N_22990,N_22763,N_22669);
or U22991 (N_22991,N_22245,N_22444);
xnor U22992 (N_22992,N_22672,N_22461);
and U22993 (N_22993,N_22261,N_22307);
nor U22994 (N_22994,N_22381,N_22795);
nor U22995 (N_22995,N_22699,N_22496);
xor U22996 (N_22996,N_22796,N_22345);
nor U22997 (N_22997,N_22616,N_22647);
nand U22998 (N_22998,N_22336,N_22743);
xor U22999 (N_22999,N_22310,N_22714);
or U23000 (N_23000,N_22652,N_22228);
xnor U23001 (N_23001,N_22367,N_22742);
xnor U23002 (N_23002,N_22463,N_22371);
and U23003 (N_23003,N_22760,N_22258);
nor U23004 (N_23004,N_22682,N_22304);
and U23005 (N_23005,N_22607,N_22340);
or U23006 (N_23006,N_22468,N_22350);
nor U23007 (N_23007,N_22565,N_22589);
nand U23008 (N_23008,N_22388,N_22401);
nand U23009 (N_23009,N_22234,N_22681);
and U23010 (N_23010,N_22657,N_22784);
nand U23011 (N_23011,N_22700,N_22506);
nor U23012 (N_23012,N_22446,N_22281);
nand U23013 (N_23013,N_22626,N_22708);
or U23014 (N_23014,N_22529,N_22276);
or U23015 (N_23015,N_22295,N_22312);
or U23016 (N_23016,N_22309,N_22633);
or U23017 (N_23017,N_22603,N_22211);
and U23018 (N_23018,N_22791,N_22271);
or U23019 (N_23019,N_22266,N_22710);
nand U23020 (N_23020,N_22548,N_22578);
nor U23021 (N_23021,N_22688,N_22619);
xor U23022 (N_23022,N_22246,N_22555);
or U23023 (N_23023,N_22206,N_22244);
nor U23024 (N_23024,N_22488,N_22713);
nand U23025 (N_23025,N_22239,N_22479);
and U23026 (N_23026,N_22386,N_22264);
xnor U23027 (N_23027,N_22484,N_22705);
nor U23028 (N_23028,N_22559,N_22504);
xor U23029 (N_23029,N_22410,N_22392);
nand U23030 (N_23030,N_22764,N_22341);
xnor U23031 (N_23031,N_22653,N_22624);
or U23032 (N_23032,N_22508,N_22778);
nor U23033 (N_23033,N_22549,N_22611);
and U23034 (N_23034,N_22608,N_22561);
or U23035 (N_23035,N_22703,N_22203);
or U23036 (N_23036,N_22248,N_22643);
and U23037 (N_23037,N_22557,N_22337);
or U23038 (N_23038,N_22325,N_22689);
or U23039 (N_23039,N_22702,N_22740);
xnor U23040 (N_23040,N_22646,N_22339);
and U23041 (N_23041,N_22536,N_22250);
xnor U23042 (N_23042,N_22685,N_22335);
nor U23043 (N_23043,N_22374,N_22220);
nand U23044 (N_23044,N_22775,N_22560);
or U23045 (N_23045,N_22587,N_22501);
nand U23046 (N_23046,N_22615,N_22628);
xnor U23047 (N_23047,N_22426,N_22433);
nor U23048 (N_23048,N_22642,N_22252);
or U23049 (N_23049,N_22788,N_22436);
nand U23050 (N_23050,N_22648,N_22467);
nor U23051 (N_23051,N_22298,N_22585);
xor U23052 (N_23052,N_22577,N_22667);
and U23053 (N_23053,N_22362,N_22684);
xor U23054 (N_23054,N_22377,N_22664);
or U23055 (N_23055,N_22675,N_22431);
xnor U23056 (N_23056,N_22530,N_22286);
nor U23057 (N_23057,N_22623,N_22541);
or U23058 (N_23058,N_22543,N_22538);
and U23059 (N_23059,N_22636,N_22287);
nand U23060 (N_23060,N_22328,N_22419);
xnor U23061 (N_23061,N_22400,N_22546);
xor U23062 (N_23062,N_22581,N_22593);
nand U23063 (N_23063,N_22409,N_22253);
nand U23064 (N_23064,N_22301,N_22413);
nor U23065 (N_23065,N_22359,N_22604);
and U23066 (N_23066,N_22696,N_22709);
nand U23067 (N_23067,N_22229,N_22291);
and U23068 (N_23068,N_22755,N_22645);
or U23069 (N_23069,N_22735,N_22308);
and U23070 (N_23070,N_22469,N_22403);
and U23071 (N_23071,N_22200,N_22602);
nor U23072 (N_23072,N_22303,N_22721);
xnor U23073 (N_23073,N_22718,N_22393);
and U23074 (N_23074,N_22215,N_22732);
and U23075 (N_23075,N_22741,N_22313);
and U23076 (N_23076,N_22551,N_22320);
nand U23077 (N_23077,N_22622,N_22649);
nor U23078 (N_23078,N_22240,N_22533);
or U23079 (N_23079,N_22717,N_22516);
nor U23080 (N_23080,N_22322,N_22297);
or U23081 (N_23081,N_22305,N_22486);
nand U23082 (N_23082,N_22218,N_22277);
nor U23083 (N_23083,N_22389,N_22472);
and U23084 (N_23084,N_22470,N_22432);
or U23085 (N_23085,N_22580,N_22366);
or U23086 (N_23086,N_22254,N_22485);
nor U23087 (N_23087,N_22573,N_22728);
nor U23088 (N_23088,N_22674,N_22590);
xnor U23089 (N_23089,N_22609,N_22243);
nand U23090 (N_23090,N_22659,N_22596);
and U23091 (N_23091,N_22398,N_22478);
nor U23092 (N_23092,N_22711,N_22317);
nand U23093 (N_23093,N_22678,N_22753);
nand U23094 (N_23094,N_22595,N_22707);
or U23095 (N_23095,N_22368,N_22330);
xor U23096 (N_23096,N_22241,N_22369);
and U23097 (N_23097,N_22343,N_22761);
xnor U23098 (N_23098,N_22259,N_22629);
and U23099 (N_23099,N_22232,N_22701);
nand U23100 (N_23100,N_22277,N_22317);
or U23101 (N_23101,N_22624,N_22310);
and U23102 (N_23102,N_22211,N_22498);
nor U23103 (N_23103,N_22656,N_22459);
nand U23104 (N_23104,N_22254,N_22550);
xor U23105 (N_23105,N_22651,N_22614);
and U23106 (N_23106,N_22230,N_22274);
xnor U23107 (N_23107,N_22339,N_22394);
or U23108 (N_23108,N_22288,N_22340);
nand U23109 (N_23109,N_22660,N_22611);
nor U23110 (N_23110,N_22377,N_22718);
nand U23111 (N_23111,N_22648,N_22561);
nor U23112 (N_23112,N_22490,N_22700);
or U23113 (N_23113,N_22765,N_22662);
nor U23114 (N_23114,N_22301,N_22480);
or U23115 (N_23115,N_22779,N_22650);
or U23116 (N_23116,N_22484,N_22358);
xnor U23117 (N_23117,N_22296,N_22259);
nand U23118 (N_23118,N_22215,N_22337);
or U23119 (N_23119,N_22521,N_22228);
nand U23120 (N_23120,N_22283,N_22693);
xor U23121 (N_23121,N_22234,N_22265);
nor U23122 (N_23122,N_22562,N_22264);
or U23123 (N_23123,N_22762,N_22735);
nor U23124 (N_23124,N_22501,N_22693);
nor U23125 (N_23125,N_22492,N_22301);
and U23126 (N_23126,N_22347,N_22380);
nand U23127 (N_23127,N_22660,N_22635);
or U23128 (N_23128,N_22205,N_22637);
and U23129 (N_23129,N_22381,N_22225);
xor U23130 (N_23130,N_22701,N_22686);
xnor U23131 (N_23131,N_22372,N_22783);
or U23132 (N_23132,N_22275,N_22721);
xor U23133 (N_23133,N_22261,N_22660);
and U23134 (N_23134,N_22226,N_22557);
nor U23135 (N_23135,N_22293,N_22341);
nor U23136 (N_23136,N_22736,N_22672);
nor U23137 (N_23137,N_22769,N_22422);
xor U23138 (N_23138,N_22541,N_22569);
nand U23139 (N_23139,N_22226,N_22603);
xor U23140 (N_23140,N_22590,N_22390);
nor U23141 (N_23141,N_22282,N_22461);
nand U23142 (N_23142,N_22740,N_22321);
nor U23143 (N_23143,N_22208,N_22207);
nand U23144 (N_23144,N_22550,N_22276);
and U23145 (N_23145,N_22578,N_22264);
nor U23146 (N_23146,N_22371,N_22745);
xnor U23147 (N_23147,N_22615,N_22392);
nand U23148 (N_23148,N_22486,N_22337);
and U23149 (N_23149,N_22675,N_22212);
and U23150 (N_23150,N_22499,N_22515);
xnor U23151 (N_23151,N_22341,N_22486);
xnor U23152 (N_23152,N_22730,N_22473);
xnor U23153 (N_23153,N_22787,N_22735);
or U23154 (N_23154,N_22450,N_22688);
nor U23155 (N_23155,N_22302,N_22314);
or U23156 (N_23156,N_22790,N_22792);
nor U23157 (N_23157,N_22684,N_22590);
xnor U23158 (N_23158,N_22615,N_22432);
nor U23159 (N_23159,N_22248,N_22294);
nor U23160 (N_23160,N_22778,N_22642);
xor U23161 (N_23161,N_22692,N_22586);
and U23162 (N_23162,N_22762,N_22758);
nor U23163 (N_23163,N_22264,N_22783);
nor U23164 (N_23164,N_22645,N_22426);
nand U23165 (N_23165,N_22233,N_22238);
nor U23166 (N_23166,N_22541,N_22256);
and U23167 (N_23167,N_22337,N_22307);
or U23168 (N_23168,N_22414,N_22490);
nand U23169 (N_23169,N_22351,N_22560);
xor U23170 (N_23170,N_22356,N_22468);
nor U23171 (N_23171,N_22548,N_22793);
nor U23172 (N_23172,N_22202,N_22378);
and U23173 (N_23173,N_22705,N_22613);
and U23174 (N_23174,N_22750,N_22274);
and U23175 (N_23175,N_22258,N_22558);
nand U23176 (N_23176,N_22645,N_22627);
nand U23177 (N_23177,N_22678,N_22260);
and U23178 (N_23178,N_22353,N_22441);
nand U23179 (N_23179,N_22716,N_22622);
nand U23180 (N_23180,N_22399,N_22635);
and U23181 (N_23181,N_22232,N_22491);
xnor U23182 (N_23182,N_22721,N_22255);
or U23183 (N_23183,N_22546,N_22321);
xnor U23184 (N_23184,N_22780,N_22275);
nand U23185 (N_23185,N_22638,N_22664);
or U23186 (N_23186,N_22443,N_22295);
and U23187 (N_23187,N_22787,N_22726);
nand U23188 (N_23188,N_22217,N_22255);
nor U23189 (N_23189,N_22548,N_22372);
xnor U23190 (N_23190,N_22605,N_22628);
and U23191 (N_23191,N_22775,N_22244);
nor U23192 (N_23192,N_22245,N_22657);
or U23193 (N_23193,N_22734,N_22533);
or U23194 (N_23194,N_22399,N_22631);
and U23195 (N_23195,N_22204,N_22785);
and U23196 (N_23196,N_22697,N_22337);
or U23197 (N_23197,N_22478,N_22762);
or U23198 (N_23198,N_22527,N_22203);
and U23199 (N_23199,N_22397,N_22314);
and U23200 (N_23200,N_22716,N_22338);
and U23201 (N_23201,N_22437,N_22416);
xnor U23202 (N_23202,N_22572,N_22389);
nand U23203 (N_23203,N_22205,N_22338);
and U23204 (N_23204,N_22301,N_22263);
or U23205 (N_23205,N_22759,N_22560);
or U23206 (N_23206,N_22440,N_22769);
nor U23207 (N_23207,N_22329,N_22530);
nand U23208 (N_23208,N_22450,N_22626);
or U23209 (N_23209,N_22466,N_22301);
xnor U23210 (N_23210,N_22663,N_22690);
xnor U23211 (N_23211,N_22429,N_22503);
nand U23212 (N_23212,N_22589,N_22509);
xnor U23213 (N_23213,N_22235,N_22704);
or U23214 (N_23214,N_22569,N_22690);
nand U23215 (N_23215,N_22598,N_22442);
xnor U23216 (N_23216,N_22579,N_22435);
nand U23217 (N_23217,N_22222,N_22792);
xor U23218 (N_23218,N_22536,N_22799);
or U23219 (N_23219,N_22256,N_22205);
or U23220 (N_23220,N_22485,N_22238);
nor U23221 (N_23221,N_22698,N_22390);
nand U23222 (N_23222,N_22228,N_22338);
nand U23223 (N_23223,N_22549,N_22463);
nor U23224 (N_23224,N_22301,N_22399);
nor U23225 (N_23225,N_22697,N_22571);
nand U23226 (N_23226,N_22559,N_22459);
and U23227 (N_23227,N_22323,N_22617);
and U23228 (N_23228,N_22538,N_22768);
and U23229 (N_23229,N_22646,N_22395);
xor U23230 (N_23230,N_22332,N_22484);
or U23231 (N_23231,N_22400,N_22758);
xnor U23232 (N_23232,N_22702,N_22229);
nand U23233 (N_23233,N_22399,N_22249);
and U23234 (N_23234,N_22453,N_22672);
nand U23235 (N_23235,N_22602,N_22354);
nor U23236 (N_23236,N_22329,N_22501);
xnor U23237 (N_23237,N_22567,N_22551);
xor U23238 (N_23238,N_22712,N_22243);
nand U23239 (N_23239,N_22430,N_22675);
nor U23240 (N_23240,N_22598,N_22234);
or U23241 (N_23241,N_22472,N_22455);
nor U23242 (N_23242,N_22473,N_22491);
xor U23243 (N_23243,N_22673,N_22451);
and U23244 (N_23244,N_22304,N_22691);
or U23245 (N_23245,N_22391,N_22244);
nand U23246 (N_23246,N_22218,N_22574);
xnor U23247 (N_23247,N_22285,N_22313);
xnor U23248 (N_23248,N_22371,N_22309);
xor U23249 (N_23249,N_22510,N_22201);
or U23250 (N_23250,N_22383,N_22619);
nand U23251 (N_23251,N_22465,N_22315);
xnor U23252 (N_23252,N_22574,N_22681);
xor U23253 (N_23253,N_22571,N_22325);
and U23254 (N_23254,N_22596,N_22584);
or U23255 (N_23255,N_22303,N_22362);
nor U23256 (N_23256,N_22489,N_22454);
xnor U23257 (N_23257,N_22449,N_22601);
and U23258 (N_23258,N_22671,N_22260);
or U23259 (N_23259,N_22788,N_22461);
nand U23260 (N_23260,N_22519,N_22661);
and U23261 (N_23261,N_22259,N_22512);
xnor U23262 (N_23262,N_22317,N_22572);
and U23263 (N_23263,N_22775,N_22464);
nor U23264 (N_23264,N_22794,N_22201);
and U23265 (N_23265,N_22729,N_22629);
or U23266 (N_23266,N_22641,N_22592);
nor U23267 (N_23267,N_22225,N_22419);
and U23268 (N_23268,N_22487,N_22532);
or U23269 (N_23269,N_22434,N_22352);
nand U23270 (N_23270,N_22648,N_22721);
nand U23271 (N_23271,N_22207,N_22298);
nor U23272 (N_23272,N_22625,N_22610);
nand U23273 (N_23273,N_22268,N_22513);
or U23274 (N_23274,N_22234,N_22428);
nand U23275 (N_23275,N_22752,N_22450);
xor U23276 (N_23276,N_22466,N_22394);
nand U23277 (N_23277,N_22795,N_22742);
nor U23278 (N_23278,N_22245,N_22537);
nand U23279 (N_23279,N_22657,N_22396);
xnor U23280 (N_23280,N_22724,N_22376);
nor U23281 (N_23281,N_22454,N_22481);
xnor U23282 (N_23282,N_22233,N_22535);
and U23283 (N_23283,N_22342,N_22701);
nand U23284 (N_23284,N_22230,N_22761);
nor U23285 (N_23285,N_22435,N_22554);
xor U23286 (N_23286,N_22363,N_22259);
and U23287 (N_23287,N_22633,N_22798);
nand U23288 (N_23288,N_22685,N_22438);
nor U23289 (N_23289,N_22253,N_22433);
nor U23290 (N_23290,N_22442,N_22508);
or U23291 (N_23291,N_22732,N_22222);
nor U23292 (N_23292,N_22759,N_22652);
and U23293 (N_23293,N_22662,N_22352);
nand U23294 (N_23294,N_22798,N_22327);
or U23295 (N_23295,N_22468,N_22783);
nor U23296 (N_23296,N_22224,N_22711);
and U23297 (N_23297,N_22452,N_22648);
and U23298 (N_23298,N_22769,N_22367);
and U23299 (N_23299,N_22284,N_22469);
xor U23300 (N_23300,N_22628,N_22258);
and U23301 (N_23301,N_22531,N_22669);
xnor U23302 (N_23302,N_22216,N_22556);
xnor U23303 (N_23303,N_22662,N_22474);
nand U23304 (N_23304,N_22755,N_22696);
nand U23305 (N_23305,N_22661,N_22739);
nor U23306 (N_23306,N_22290,N_22397);
nand U23307 (N_23307,N_22483,N_22367);
and U23308 (N_23308,N_22237,N_22619);
or U23309 (N_23309,N_22379,N_22543);
and U23310 (N_23310,N_22560,N_22694);
nand U23311 (N_23311,N_22527,N_22329);
and U23312 (N_23312,N_22388,N_22462);
or U23313 (N_23313,N_22799,N_22274);
nand U23314 (N_23314,N_22468,N_22741);
xor U23315 (N_23315,N_22393,N_22249);
xor U23316 (N_23316,N_22280,N_22286);
or U23317 (N_23317,N_22503,N_22683);
xor U23318 (N_23318,N_22697,N_22323);
nor U23319 (N_23319,N_22443,N_22698);
or U23320 (N_23320,N_22471,N_22709);
nor U23321 (N_23321,N_22618,N_22404);
nor U23322 (N_23322,N_22259,N_22216);
and U23323 (N_23323,N_22273,N_22430);
or U23324 (N_23324,N_22536,N_22590);
xnor U23325 (N_23325,N_22450,N_22783);
or U23326 (N_23326,N_22528,N_22383);
nand U23327 (N_23327,N_22697,N_22225);
and U23328 (N_23328,N_22507,N_22766);
nand U23329 (N_23329,N_22758,N_22219);
or U23330 (N_23330,N_22437,N_22362);
nand U23331 (N_23331,N_22642,N_22229);
nand U23332 (N_23332,N_22321,N_22396);
nand U23333 (N_23333,N_22632,N_22540);
nor U23334 (N_23334,N_22589,N_22414);
xor U23335 (N_23335,N_22750,N_22353);
or U23336 (N_23336,N_22266,N_22638);
or U23337 (N_23337,N_22743,N_22263);
nand U23338 (N_23338,N_22364,N_22779);
nand U23339 (N_23339,N_22549,N_22645);
nand U23340 (N_23340,N_22396,N_22689);
nand U23341 (N_23341,N_22460,N_22203);
and U23342 (N_23342,N_22332,N_22500);
and U23343 (N_23343,N_22466,N_22411);
xnor U23344 (N_23344,N_22303,N_22723);
or U23345 (N_23345,N_22458,N_22798);
and U23346 (N_23346,N_22636,N_22472);
nor U23347 (N_23347,N_22566,N_22676);
nor U23348 (N_23348,N_22684,N_22568);
nor U23349 (N_23349,N_22693,N_22312);
nor U23350 (N_23350,N_22617,N_22471);
nand U23351 (N_23351,N_22630,N_22223);
xor U23352 (N_23352,N_22621,N_22253);
nor U23353 (N_23353,N_22677,N_22464);
or U23354 (N_23354,N_22706,N_22678);
or U23355 (N_23355,N_22458,N_22329);
or U23356 (N_23356,N_22430,N_22466);
nand U23357 (N_23357,N_22299,N_22594);
nand U23358 (N_23358,N_22753,N_22429);
nand U23359 (N_23359,N_22726,N_22322);
or U23360 (N_23360,N_22415,N_22584);
and U23361 (N_23361,N_22590,N_22612);
nand U23362 (N_23362,N_22652,N_22411);
nand U23363 (N_23363,N_22598,N_22525);
xor U23364 (N_23364,N_22519,N_22652);
and U23365 (N_23365,N_22254,N_22579);
or U23366 (N_23366,N_22480,N_22488);
nor U23367 (N_23367,N_22291,N_22367);
and U23368 (N_23368,N_22448,N_22340);
nand U23369 (N_23369,N_22389,N_22702);
and U23370 (N_23370,N_22336,N_22608);
nand U23371 (N_23371,N_22332,N_22334);
xnor U23372 (N_23372,N_22641,N_22626);
or U23373 (N_23373,N_22334,N_22248);
nand U23374 (N_23374,N_22729,N_22368);
and U23375 (N_23375,N_22557,N_22439);
or U23376 (N_23376,N_22558,N_22601);
nor U23377 (N_23377,N_22638,N_22693);
or U23378 (N_23378,N_22553,N_22501);
nand U23379 (N_23379,N_22349,N_22675);
xnor U23380 (N_23380,N_22319,N_22464);
nor U23381 (N_23381,N_22467,N_22349);
nor U23382 (N_23382,N_22266,N_22211);
nor U23383 (N_23383,N_22620,N_22360);
or U23384 (N_23384,N_22712,N_22597);
xnor U23385 (N_23385,N_22363,N_22304);
xor U23386 (N_23386,N_22218,N_22226);
nor U23387 (N_23387,N_22282,N_22786);
nor U23388 (N_23388,N_22561,N_22697);
nand U23389 (N_23389,N_22206,N_22429);
nand U23390 (N_23390,N_22480,N_22744);
and U23391 (N_23391,N_22784,N_22481);
nor U23392 (N_23392,N_22675,N_22316);
or U23393 (N_23393,N_22386,N_22281);
and U23394 (N_23394,N_22761,N_22397);
or U23395 (N_23395,N_22372,N_22589);
nand U23396 (N_23396,N_22558,N_22659);
nor U23397 (N_23397,N_22211,N_22373);
and U23398 (N_23398,N_22466,N_22547);
nor U23399 (N_23399,N_22282,N_22302);
xor U23400 (N_23400,N_23218,N_23142);
xor U23401 (N_23401,N_23055,N_23350);
nor U23402 (N_23402,N_23204,N_23390);
or U23403 (N_23403,N_23301,N_23287);
and U23404 (N_23404,N_23184,N_23334);
nor U23405 (N_23405,N_23082,N_23379);
nand U23406 (N_23406,N_23272,N_23393);
nor U23407 (N_23407,N_23199,N_23254);
or U23408 (N_23408,N_22893,N_23398);
nand U23409 (N_23409,N_22899,N_23126);
or U23410 (N_23410,N_23345,N_22977);
and U23411 (N_23411,N_23212,N_22842);
or U23412 (N_23412,N_22821,N_23361);
nand U23413 (N_23413,N_23356,N_23031);
xnor U23414 (N_23414,N_23009,N_23144);
nand U23415 (N_23415,N_23081,N_22817);
nor U23416 (N_23416,N_23170,N_23169);
or U23417 (N_23417,N_23022,N_23134);
or U23418 (N_23418,N_22960,N_23291);
nor U23419 (N_23419,N_23365,N_23303);
nand U23420 (N_23420,N_23122,N_23264);
nor U23421 (N_23421,N_22830,N_23066);
nand U23422 (N_23422,N_22945,N_23335);
or U23423 (N_23423,N_23226,N_22897);
nor U23424 (N_23424,N_23289,N_23056);
xnor U23425 (N_23425,N_22949,N_23131);
nand U23426 (N_23426,N_23186,N_22826);
and U23427 (N_23427,N_23174,N_23098);
and U23428 (N_23428,N_23239,N_22844);
or U23429 (N_23429,N_23075,N_23214);
nand U23430 (N_23430,N_23052,N_23331);
xnor U23431 (N_23431,N_22909,N_23358);
nand U23432 (N_23432,N_23112,N_22995);
nor U23433 (N_23433,N_23211,N_23215);
and U23434 (N_23434,N_22970,N_22981);
and U23435 (N_23435,N_23389,N_23093);
or U23436 (N_23436,N_22860,N_22916);
or U23437 (N_23437,N_23036,N_23300);
xor U23438 (N_23438,N_23103,N_23281);
nand U23439 (N_23439,N_23030,N_23258);
or U23440 (N_23440,N_23399,N_23090);
and U23441 (N_23441,N_22903,N_22965);
nor U23442 (N_23442,N_23124,N_23275);
nor U23443 (N_23443,N_22962,N_23306);
and U23444 (N_23444,N_22913,N_22998);
or U23445 (N_23445,N_22983,N_23140);
and U23446 (N_23446,N_22859,N_22801);
nor U23447 (N_23447,N_23241,N_23005);
nor U23448 (N_23448,N_22991,N_23373);
nand U23449 (N_23449,N_22939,N_23012);
or U23450 (N_23450,N_23385,N_23305);
xor U23451 (N_23451,N_23064,N_23282);
and U23452 (N_23452,N_22999,N_23027);
xnor U23453 (N_23453,N_22865,N_22959);
nor U23454 (N_23454,N_22871,N_23222);
or U23455 (N_23455,N_22941,N_23247);
nor U23456 (N_23456,N_22805,N_23260);
or U23457 (N_23457,N_23276,N_23020);
and U23458 (N_23458,N_23168,N_23352);
or U23459 (N_23459,N_23007,N_23245);
xnor U23460 (N_23460,N_23363,N_22819);
xor U23461 (N_23461,N_23357,N_23227);
nor U23462 (N_23462,N_22803,N_22831);
nand U23463 (N_23463,N_23203,N_23109);
nand U23464 (N_23464,N_23362,N_22815);
or U23465 (N_23465,N_23319,N_22809);
nor U23466 (N_23466,N_23173,N_23206);
or U23467 (N_23467,N_23375,N_23128);
xor U23468 (N_23468,N_22812,N_22984);
nor U23469 (N_23469,N_23015,N_23263);
xnor U23470 (N_23470,N_23394,N_23202);
nor U23471 (N_23471,N_23298,N_22902);
nor U23472 (N_23472,N_23296,N_23014);
and U23473 (N_23473,N_23327,N_23304);
nor U23474 (N_23474,N_22980,N_22832);
nand U23475 (N_23475,N_23002,N_23021);
or U23476 (N_23476,N_22943,N_22811);
xnor U23477 (N_23477,N_23072,N_23294);
nand U23478 (N_23478,N_23155,N_23129);
or U23479 (N_23479,N_22823,N_23164);
nor U23480 (N_23480,N_22979,N_23297);
nand U23481 (N_23481,N_23051,N_23384);
and U23482 (N_23482,N_22864,N_23091);
and U23483 (N_23483,N_23228,N_22892);
nand U23484 (N_23484,N_23286,N_23196);
nand U23485 (N_23485,N_23078,N_23299);
and U23486 (N_23486,N_23261,N_23382);
and U23487 (N_23487,N_23323,N_22907);
or U23488 (N_23488,N_22901,N_23154);
nor U23489 (N_23489,N_23029,N_22935);
nor U23490 (N_23490,N_23223,N_23339);
xor U23491 (N_23491,N_23079,N_23018);
or U23492 (N_23492,N_23201,N_23084);
nand U23493 (N_23493,N_23067,N_23285);
nor U23494 (N_23494,N_23351,N_22874);
and U23495 (N_23495,N_22967,N_23354);
nor U23496 (N_23496,N_23102,N_23086);
and U23497 (N_23497,N_23000,N_23041);
and U23498 (N_23498,N_23267,N_23376);
and U23499 (N_23499,N_22861,N_23355);
or U23500 (N_23500,N_23195,N_23006);
or U23501 (N_23501,N_22872,N_23187);
or U23502 (N_23502,N_23366,N_23225);
or U23503 (N_23503,N_22827,N_22848);
nand U23504 (N_23504,N_23085,N_23293);
nor U23505 (N_23505,N_23035,N_23185);
nand U23506 (N_23506,N_23229,N_23117);
nand U23507 (N_23507,N_23059,N_23312);
or U23508 (N_23508,N_22867,N_22870);
or U23509 (N_23509,N_22934,N_23388);
xor U23510 (N_23510,N_22988,N_23138);
xor U23511 (N_23511,N_22932,N_22822);
and U23512 (N_23512,N_22919,N_23116);
and U23513 (N_23513,N_22887,N_23065);
and U23514 (N_23514,N_23050,N_23324);
and U23515 (N_23515,N_22834,N_23364);
nand U23516 (N_23516,N_23274,N_23307);
nand U23517 (N_23517,N_22989,N_23045);
xnor U23518 (N_23518,N_23283,N_23244);
nand U23519 (N_23519,N_23161,N_22917);
nor U23520 (N_23520,N_23318,N_23231);
xnor U23521 (N_23521,N_23172,N_23210);
nand U23522 (N_23522,N_22938,N_22898);
and U23523 (N_23523,N_23205,N_23383);
or U23524 (N_23524,N_23233,N_22806);
nand U23525 (N_23525,N_23042,N_22888);
xor U23526 (N_23526,N_22966,N_23160);
xor U23527 (N_23527,N_23380,N_23137);
or U23528 (N_23528,N_23234,N_22845);
nand U23529 (N_23529,N_22857,N_23118);
or U23530 (N_23530,N_22851,N_23290);
nand U23531 (N_23531,N_23236,N_22863);
nand U23532 (N_23532,N_23209,N_23026);
or U23533 (N_23533,N_22884,N_23110);
nand U23534 (N_23534,N_22910,N_23265);
or U23535 (N_23535,N_22964,N_23353);
or U23536 (N_23536,N_22849,N_23177);
nor U23537 (N_23537,N_23284,N_23151);
xor U23538 (N_23538,N_23044,N_23280);
or U23539 (N_23539,N_22891,N_23068);
and U23540 (N_23540,N_22818,N_22882);
and U23541 (N_23541,N_22900,N_23370);
and U23542 (N_23542,N_23221,N_23054);
nand U23543 (N_23543,N_22956,N_23217);
or U23544 (N_23544,N_23266,N_23004);
nand U23545 (N_23545,N_23342,N_23381);
and U23546 (N_23546,N_23008,N_23387);
or U23547 (N_23547,N_22946,N_23347);
and U23548 (N_23548,N_22868,N_23270);
or U23549 (N_23549,N_23190,N_22914);
and U23550 (N_23550,N_23094,N_23251);
nor U23551 (N_23551,N_23073,N_23321);
and U23552 (N_23552,N_23048,N_22982);
xnor U23553 (N_23553,N_23273,N_23369);
nor U23554 (N_23554,N_23314,N_23242);
nor U23555 (N_23555,N_23145,N_23329);
nand U23556 (N_23556,N_22813,N_22931);
nand U23557 (N_23557,N_23250,N_23277);
xor U23558 (N_23558,N_22896,N_22974);
nand U23559 (N_23559,N_23011,N_23333);
xor U23560 (N_23560,N_23060,N_22918);
and U23561 (N_23561,N_22942,N_23038);
xor U23562 (N_23562,N_23188,N_23033);
or U23563 (N_23563,N_22824,N_22869);
nor U23564 (N_23564,N_23108,N_23371);
or U23565 (N_23565,N_23213,N_22958);
nor U23566 (N_23566,N_23087,N_22814);
and U23567 (N_23567,N_22883,N_23158);
xnor U23568 (N_23568,N_22856,N_23043);
nand U23569 (N_23569,N_22854,N_23180);
nor U23570 (N_23570,N_23183,N_23163);
or U23571 (N_23571,N_23189,N_22846);
and U23572 (N_23572,N_23175,N_23107);
xor U23573 (N_23573,N_23147,N_22866);
nand U23574 (N_23574,N_23097,N_23238);
or U23575 (N_23575,N_22880,N_23315);
nor U23576 (N_23576,N_23178,N_22937);
nor U23577 (N_23577,N_23113,N_23359);
and U23578 (N_23578,N_22972,N_23246);
or U23579 (N_23579,N_22894,N_22895);
nor U23580 (N_23580,N_22828,N_23368);
or U23581 (N_23581,N_23176,N_23136);
xor U23582 (N_23582,N_23132,N_23313);
xnor U23583 (N_23583,N_23083,N_23070);
nand U23584 (N_23584,N_23104,N_23232);
nor U23585 (N_23585,N_23088,N_22904);
nor U23586 (N_23586,N_23121,N_23336);
xor U23587 (N_23587,N_23243,N_22862);
nand U23588 (N_23588,N_22922,N_22853);
nor U23589 (N_23589,N_23235,N_22947);
and U23590 (N_23590,N_23058,N_23278);
xnor U23591 (N_23591,N_23023,N_22976);
nand U23592 (N_23592,N_23230,N_22825);
and U23593 (N_23593,N_23208,N_23099);
nor U23594 (N_23594,N_23332,N_23295);
xor U23595 (N_23595,N_23115,N_22843);
nand U23596 (N_23596,N_23193,N_22929);
nor U23597 (N_23597,N_22858,N_23240);
or U23598 (N_23598,N_22948,N_23325);
xor U23599 (N_23599,N_22920,N_22876);
xnor U23600 (N_23600,N_23157,N_23153);
nand U23601 (N_23601,N_23148,N_23292);
and U23602 (N_23602,N_23194,N_23089);
or U23603 (N_23603,N_23156,N_23063);
and U23604 (N_23604,N_23396,N_22975);
and U23605 (N_23605,N_22800,N_23092);
or U23606 (N_23606,N_22839,N_23077);
and U23607 (N_23607,N_22921,N_23360);
nor U23608 (N_23608,N_23047,N_23253);
and U23609 (N_23609,N_23271,N_22928);
xor U23610 (N_23610,N_23344,N_23025);
xor U23611 (N_23611,N_23224,N_22915);
and U23612 (N_23612,N_22997,N_23049);
or U23613 (N_23613,N_23057,N_23198);
and U23614 (N_23614,N_22993,N_23262);
xor U23615 (N_23615,N_23374,N_23237);
nor U23616 (N_23616,N_23395,N_23162);
or U23617 (N_23617,N_22940,N_23320);
xor U23618 (N_23618,N_22838,N_23001);
or U23619 (N_23619,N_23207,N_22875);
nand U23620 (N_23620,N_23053,N_23167);
xnor U23621 (N_23621,N_23181,N_22924);
and U23622 (N_23622,N_23034,N_22835);
nand U23623 (N_23623,N_23096,N_23219);
xor U23624 (N_23624,N_23200,N_23133);
nor U23625 (N_23625,N_23252,N_22837);
or U23626 (N_23626,N_23111,N_22930);
or U23627 (N_23627,N_22885,N_23119);
nor U23628 (N_23628,N_23003,N_23191);
nand U23629 (N_23629,N_22836,N_22911);
xnor U23630 (N_23630,N_22933,N_23114);
nor U23631 (N_23631,N_23037,N_23197);
nor U23632 (N_23632,N_22816,N_23143);
or U23633 (N_23633,N_22810,N_23372);
nor U23634 (N_23634,N_23269,N_22992);
xor U23635 (N_23635,N_22961,N_23159);
xnor U23636 (N_23636,N_23391,N_23309);
nor U23637 (N_23637,N_23182,N_23179);
xnor U23638 (N_23638,N_22936,N_22820);
nand U23639 (N_23639,N_23279,N_22829);
or U23640 (N_23640,N_23377,N_22886);
and U23641 (N_23641,N_23255,N_22881);
nand U23642 (N_23642,N_23046,N_23016);
nand U23643 (N_23643,N_23386,N_22802);
nor U23644 (N_23644,N_23248,N_22953);
xnor U23645 (N_23645,N_22878,N_23101);
nand U23646 (N_23646,N_23302,N_22952);
and U23647 (N_23647,N_22994,N_22879);
xnor U23648 (N_23648,N_23013,N_23216);
xor U23649 (N_23649,N_22906,N_23397);
and U23650 (N_23650,N_22890,N_23348);
or U23651 (N_23651,N_23328,N_22808);
and U23652 (N_23652,N_22850,N_22971);
nand U23653 (N_23653,N_23061,N_23139);
or U23654 (N_23654,N_22855,N_23076);
or U23655 (N_23655,N_23039,N_23322);
nor U23656 (N_23656,N_23257,N_23123);
nor U23657 (N_23657,N_23392,N_23316);
or U23658 (N_23658,N_22877,N_22873);
and U23659 (N_23659,N_23120,N_22950);
or U23660 (N_23660,N_23166,N_23171);
or U23661 (N_23661,N_23330,N_23141);
and U23662 (N_23662,N_22926,N_23268);
nor U23663 (N_23663,N_23311,N_23152);
and U23664 (N_23664,N_23080,N_23149);
xnor U23665 (N_23665,N_23337,N_23105);
and U23666 (N_23666,N_23074,N_23346);
and U23667 (N_23667,N_23349,N_23338);
xor U23668 (N_23668,N_22927,N_22908);
nor U23669 (N_23669,N_23317,N_23106);
or U23670 (N_23670,N_23032,N_23146);
xnor U23671 (N_23671,N_22963,N_22955);
xor U23672 (N_23672,N_23165,N_23130);
xnor U23673 (N_23673,N_23249,N_23259);
nor U23674 (N_23674,N_23100,N_23256);
xnor U23675 (N_23675,N_23343,N_22973);
xor U23676 (N_23676,N_23024,N_22852);
and U23677 (N_23677,N_22990,N_22986);
nand U23678 (N_23678,N_22957,N_22969);
or U23679 (N_23679,N_22951,N_23341);
nor U23680 (N_23680,N_23192,N_22923);
nand U23681 (N_23681,N_23378,N_22954);
nand U23682 (N_23682,N_23125,N_22804);
nor U23683 (N_23683,N_22996,N_23062);
xnor U23684 (N_23684,N_22987,N_23069);
xnor U23685 (N_23685,N_23095,N_23028);
or U23686 (N_23686,N_22944,N_23340);
and U23687 (N_23687,N_23071,N_23288);
and U23688 (N_23688,N_22807,N_23135);
nand U23689 (N_23689,N_22978,N_23019);
nor U23690 (N_23690,N_23040,N_22985);
nor U23691 (N_23691,N_22912,N_22841);
or U23692 (N_23692,N_23127,N_22889);
nor U23693 (N_23693,N_23367,N_22925);
or U23694 (N_23694,N_23017,N_23310);
nor U23695 (N_23695,N_23010,N_22905);
xnor U23696 (N_23696,N_23150,N_22847);
nor U23697 (N_23697,N_23326,N_23308);
nor U23698 (N_23698,N_23220,N_22840);
and U23699 (N_23699,N_22968,N_22833);
or U23700 (N_23700,N_23148,N_22957);
nand U23701 (N_23701,N_23140,N_22883);
xor U23702 (N_23702,N_23030,N_23105);
nor U23703 (N_23703,N_23310,N_23311);
nor U23704 (N_23704,N_23219,N_23217);
nor U23705 (N_23705,N_23369,N_23033);
xor U23706 (N_23706,N_23113,N_22822);
or U23707 (N_23707,N_23184,N_22971);
nand U23708 (N_23708,N_22864,N_22925);
nor U23709 (N_23709,N_23236,N_22868);
and U23710 (N_23710,N_23187,N_22843);
nand U23711 (N_23711,N_22881,N_23070);
nor U23712 (N_23712,N_22895,N_22885);
nand U23713 (N_23713,N_23068,N_23320);
xor U23714 (N_23714,N_22940,N_22840);
nand U23715 (N_23715,N_23119,N_22995);
xnor U23716 (N_23716,N_23228,N_23367);
or U23717 (N_23717,N_23348,N_23246);
nand U23718 (N_23718,N_23260,N_22833);
xor U23719 (N_23719,N_23207,N_23259);
or U23720 (N_23720,N_22988,N_23297);
xor U23721 (N_23721,N_23341,N_22822);
nor U23722 (N_23722,N_23326,N_23064);
or U23723 (N_23723,N_23171,N_23157);
or U23724 (N_23724,N_23150,N_22807);
nor U23725 (N_23725,N_23370,N_23327);
nand U23726 (N_23726,N_22930,N_23318);
xor U23727 (N_23727,N_23202,N_22887);
nor U23728 (N_23728,N_23229,N_23240);
or U23729 (N_23729,N_22836,N_23159);
nand U23730 (N_23730,N_22947,N_23074);
xnor U23731 (N_23731,N_22921,N_22876);
and U23732 (N_23732,N_23287,N_22938);
xor U23733 (N_23733,N_23223,N_23163);
or U23734 (N_23734,N_23231,N_22982);
nand U23735 (N_23735,N_23190,N_23117);
xor U23736 (N_23736,N_23132,N_23007);
or U23737 (N_23737,N_23180,N_23165);
xnor U23738 (N_23738,N_23013,N_23242);
or U23739 (N_23739,N_22971,N_23009);
nand U23740 (N_23740,N_23017,N_23233);
nand U23741 (N_23741,N_23075,N_22992);
or U23742 (N_23742,N_23046,N_22870);
nor U23743 (N_23743,N_23053,N_23023);
xnor U23744 (N_23744,N_23208,N_23239);
nand U23745 (N_23745,N_22950,N_23003);
xnor U23746 (N_23746,N_23249,N_23359);
xnor U23747 (N_23747,N_22885,N_22893);
nand U23748 (N_23748,N_23134,N_23285);
and U23749 (N_23749,N_22973,N_22920);
or U23750 (N_23750,N_23169,N_23014);
and U23751 (N_23751,N_23289,N_23117);
nand U23752 (N_23752,N_22912,N_23288);
or U23753 (N_23753,N_23180,N_23019);
and U23754 (N_23754,N_23149,N_23246);
or U23755 (N_23755,N_23351,N_23150);
or U23756 (N_23756,N_23225,N_23194);
nand U23757 (N_23757,N_23398,N_22833);
nor U23758 (N_23758,N_23274,N_22925);
or U23759 (N_23759,N_23197,N_23014);
nand U23760 (N_23760,N_23268,N_23265);
xor U23761 (N_23761,N_23078,N_23178);
and U23762 (N_23762,N_22945,N_23318);
nand U23763 (N_23763,N_23332,N_22888);
nand U23764 (N_23764,N_23180,N_22920);
nor U23765 (N_23765,N_22816,N_23102);
nand U23766 (N_23766,N_23021,N_23358);
nor U23767 (N_23767,N_23293,N_23259);
nor U23768 (N_23768,N_22890,N_23091);
nand U23769 (N_23769,N_23301,N_23230);
or U23770 (N_23770,N_23196,N_22804);
or U23771 (N_23771,N_23008,N_22857);
nor U23772 (N_23772,N_23038,N_23305);
nand U23773 (N_23773,N_23046,N_22913);
nor U23774 (N_23774,N_23277,N_22904);
nor U23775 (N_23775,N_23130,N_22956);
or U23776 (N_23776,N_23085,N_23390);
xnor U23777 (N_23777,N_23059,N_23304);
nand U23778 (N_23778,N_23325,N_22955);
nor U23779 (N_23779,N_23372,N_23245);
xnor U23780 (N_23780,N_23242,N_23370);
or U23781 (N_23781,N_23273,N_23209);
xor U23782 (N_23782,N_22937,N_23336);
xor U23783 (N_23783,N_23071,N_23126);
or U23784 (N_23784,N_22851,N_22995);
xor U23785 (N_23785,N_23119,N_22916);
nor U23786 (N_23786,N_23032,N_22812);
xor U23787 (N_23787,N_22806,N_22845);
or U23788 (N_23788,N_22996,N_23273);
xor U23789 (N_23789,N_23138,N_22936);
xnor U23790 (N_23790,N_23082,N_22832);
and U23791 (N_23791,N_23364,N_22914);
and U23792 (N_23792,N_22929,N_22802);
nor U23793 (N_23793,N_23196,N_23180);
nor U23794 (N_23794,N_23199,N_23237);
and U23795 (N_23795,N_23041,N_22901);
xnor U23796 (N_23796,N_23158,N_23051);
xor U23797 (N_23797,N_23195,N_23246);
or U23798 (N_23798,N_22877,N_23231);
and U23799 (N_23799,N_23065,N_23117);
and U23800 (N_23800,N_22878,N_22963);
nand U23801 (N_23801,N_23391,N_22876);
nor U23802 (N_23802,N_22801,N_23391);
nand U23803 (N_23803,N_23089,N_23195);
or U23804 (N_23804,N_22962,N_22915);
and U23805 (N_23805,N_23034,N_23136);
and U23806 (N_23806,N_23281,N_22888);
or U23807 (N_23807,N_23225,N_22919);
xor U23808 (N_23808,N_23011,N_22923);
and U23809 (N_23809,N_23236,N_23085);
nor U23810 (N_23810,N_23097,N_23155);
nor U23811 (N_23811,N_23328,N_22862);
or U23812 (N_23812,N_23118,N_23236);
or U23813 (N_23813,N_23261,N_23349);
or U23814 (N_23814,N_23327,N_23395);
or U23815 (N_23815,N_23284,N_23258);
nor U23816 (N_23816,N_23088,N_23058);
xor U23817 (N_23817,N_23074,N_23110);
nand U23818 (N_23818,N_22809,N_23086);
or U23819 (N_23819,N_23100,N_23060);
nand U23820 (N_23820,N_22968,N_23000);
nand U23821 (N_23821,N_23355,N_22872);
or U23822 (N_23822,N_23078,N_23090);
xnor U23823 (N_23823,N_22901,N_23305);
xnor U23824 (N_23824,N_23060,N_23058);
nand U23825 (N_23825,N_23298,N_22889);
nand U23826 (N_23826,N_23007,N_22857);
nor U23827 (N_23827,N_23356,N_23377);
and U23828 (N_23828,N_23159,N_22952);
xor U23829 (N_23829,N_22822,N_23338);
nor U23830 (N_23830,N_23109,N_23141);
nand U23831 (N_23831,N_22869,N_22800);
and U23832 (N_23832,N_22895,N_23044);
and U23833 (N_23833,N_23001,N_23311);
or U23834 (N_23834,N_22997,N_23108);
and U23835 (N_23835,N_23344,N_23178);
xor U23836 (N_23836,N_23017,N_23088);
or U23837 (N_23837,N_23218,N_23022);
nor U23838 (N_23838,N_23060,N_23081);
xnor U23839 (N_23839,N_23322,N_22970);
or U23840 (N_23840,N_22842,N_22811);
nand U23841 (N_23841,N_22989,N_22921);
and U23842 (N_23842,N_23387,N_23088);
or U23843 (N_23843,N_23393,N_22933);
and U23844 (N_23844,N_23268,N_22801);
xor U23845 (N_23845,N_23194,N_23069);
and U23846 (N_23846,N_22911,N_23164);
nand U23847 (N_23847,N_22837,N_23365);
and U23848 (N_23848,N_23130,N_23013);
or U23849 (N_23849,N_23283,N_23040);
xnor U23850 (N_23850,N_23389,N_22981);
or U23851 (N_23851,N_23236,N_23288);
nand U23852 (N_23852,N_23136,N_22807);
or U23853 (N_23853,N_22903,N_22837);
nor U23854 (N_23854,N_23170,N_23031);
or U23855 (N_23855,N_23172,N_22985);
xor U23856 (N_23856,N_23312,N_22815);
xnor U23857 (N_23857,N_22888,N_23144);
and U23858 (N_23858,N_22830,N_23331);
xor U23859 (N_23859,N_22911,N_23165);
or U23860 (N_23860,N_22994,N_23223);
and U23861 (N_23861,N_23253,N_22843);
and U23862 (N_23862,N_22831,N_23017);
nor U23863 (N_23863,N_22817,N_23200);
or U23864 (N_23864,N_23258,N_22936);
xor U23865 (N_23865,N_23229,N_23014);
xnor U23866 (N_23866,N_22896,N_23364);
nor U23867 (N_23867,N_23083,N_23146);
nand U23868 (N_23868,N_23310,N_22938);
nand U23869 (N_23869,N_23227,N_23314);
or U23870 (N_23870,N_23246,N_23141);
nor U23871 (N_23871,N_23148,N_22837);
nor U23872 (N_23872,N_23390,N_23249);
nand U23873 (N_23873,N_22961,N_23304);
nand U23874 (N_23874,N_22863,N_23193);
nand U23875 (N_23875,N_23205,N_23090);
and U23876 (N_23876,N_22902,N_23358);
or U23877 (N_23877,N_23329,N_23345);
nand U23878 (N_23878,N_22995,N_22970);
nand U23879 (N_23879,N_22883,N_23166);
xor U23880 (N_23880,N_22885,N_23005);
nor U23881 (N_23881,N_23048,N_23051);
nand U23882 (N_23882,N_23227,N_22911);
or U23883 (N_23883,N_23221,N_23044);
and U23884 (N_23884,N_23178,N_22902);
and U23885 (N_23885,N_23240,N_23121);
xor U23886 (N_23886,N_23096,N_23306);
or U23887 (N_23887,N_23315,N_22879);
xnor U23888 (N_23888,N_22808,N_22887);
nor U23889 (N_23889,N_22969,N_23095);
nor U23890 (N_23890,N_23389,N_23374);
xnor U23891 (N_23891,N_23308,N_23132);
nor U23892 (N_23892,N_23259,N_23130);
nor U23893 (N_23893,N_23102,N_22859);
nand U23894 (N_23894,N_22956,N_23202);
or U23895 (N_23895,N_23116,N_23051);
or U23896 (N_23896,N_22875,N_23240);
nor U23897 (N_23897,N_23141,N_23270);
nand U23898 (N_23898,N_22803,N_23265);
and U23899 (N_23899,N_22833,N_23361);
nand U23900 (N_23900,N_23002,N_23180);
and U23901 (N_23901,N_22837,N_23213);
xnor U23902 (N_23902,N_22950,N_23324);
xnor U23903 (N_23903,N_22940,N_22809);
nor U23904 (N_23904,N_22844,N_22816);
nor U23905 (N_23905,N_22931,N_22869);
nor U23906 (N_23906,N_23064,N_22818);
nor U23907 (N_23907,N_23324,N_23196);
and U23908 (N_23908,N_22937,N_22915);
and U23909 (N_23909,N_23047,N_23050);
and U23910 (N_23910,N_22911,N_23003);
and U23911 (N_23911,N_23239,N_23037);
or U23912 (N_23912,N_22993,N_23209);
nor U23913 (N_23913,N_23218,N_22907);
and U23914 (N_23914,N_23094,N_22937);
and U23915 (N_23915,N_23053,N_23080);
or U23916 (N_23916,N_23057,N_23040);
nor U23917 (N_23917,N_23330,N_23119);
nand U23918 (N_23918,N_22879,N_23189);
nor U23919 (N_23919,N_23214,N_22803);
nand U23920 (N_23920,N_23213,N_23101);
xor U23921 (N_23921,N_23391,N_22847);
and U23922 (N_23922,N_22902,N_22822);
nand U23923 (N_23923,N_23375,N_23279);
nand U23924 (N_23924,N_23209,N_22969);
and U23925 (N_23925,N_23165,N_23146);
nor U23926 (N_23926,N_23069,N_23380);
nand U23927 (N_23927,N_22809,N_23056);
or U23928 (N_23928,N_23119,N_22838);
xnor U23929 (N_23929,N_23296,N_23169);
nor U23930 (N_23930,N_22846,N_22870);
or U23931 (N_23931,N_23025,N_22993);
nand U23932 (N_23932,N_23205,N_23258);
nor U23933 (N_23933,N_23039,N_22901);
nand U23934 (N_23934,N_23330,N_23383);
and U23935 (N_23935,N_23039,N_23171);
nand U23936 (N_23936,N_23371,N_22859);
nor U23937 (N_23937,N_23035,N_23032);
and U23938 (N_23938,N_23347,N_22857);
xor U23939 (N_23939,N_23344,N_23061);
and U23940 (N_23940,N_23260,N_23369);
or U23941 (N_23941,N_23341,N_23086);
xor U23942 (N_23942,N_23275,N_23187);
nand U23943 (N_23943,N_23082,N_23247);
nand U23944 (N_23944,N_23167,N_22852);
nor U23945 (N_23945,N_23373,N_23122);
xnor U23946 (N_23946,N_23318,N_23155);
and U23947 (N_23947,N_23024,N_23059);
nor U23948 (N_23948,N_23163,N_23326);
nor U23949 (N_23949,N_23121,N_23291);
xor U23950 (N_23950,N_22950,N_22964);
or U23951 (N_23951,N_23195,N_23319);
nor U23952 (N_23952,N_22931,N_23263);
nand U23953 (N_23953,N_22988,N_23123);
nand U23954 (N_23954,N_22943,N_22929);
or U23955 (N_23955,N_23321,N_22826);
or U23956 (N_23956,N_23075,N_23228);
xnor U23957 (N_23957,N_23272,N_23168);
nand U23958 (N_23958,N_23339,N_23350);
xor U23959 (N_23959,N_23027,N_23043);
nor U23960 (N_23960,N_23310,N_23059);
nand U23961 (N_23961,N_23195,N_23242);
or U23962 (N_23962,N_23077,N_22908);
and U23963 (N_23963,N_23017,N_22821);
nand U23964 (N_23964,N_23017,N_22928);
xor U23965 (N_23965,N_23116,N_22921);
and U23966 (N_23966,N_23265,N_23206);
and U23967 (N_23967,N_23214,N_22814);
nor U23968 (N_23968,N_22910,N_23297);
nand U23969 (N_23969,N_22886,N_22806);
nor U23970 (N_23970,N_23391,N_23335);
nor U23971 (N_23971,N_22922,N_22962);
nor U23972 (N_23972,N_22946,N_23189);
nor U23973 (N_23973,N_23160,N_23351);
xnor U23974 (N_23974,N_23109,N_22910);
and U23975 (N_23975,N_23373,N_22850);
nand U23976 (N_23976,N_22935,N_23002);
nand U23977 (N_23977,N_22894,N_23133);
and U23978 (N_23978,N_23393,N_23145);
nand U23979 (N_23979,N_23031,N_22948);
nand U23980 (N_23980,N_22999,N_23120);
and U23981 (N_23981,N_23187,N_23335);
nand U23982 (N_23982,N_23155,N_23153);
or U23983 (N_23983,N_22981,N_23085);
nor U23984 (N_23984,N_23397,N_23187);
nor U23985 (N_23985,N_23182,N_23008);
nor U23986 (N_23986,N_23273,N_22926);
and U23987 (N_23987,N_23045,N_23144);
and U23988 (N_23988,N_23254,N_22933);
nand U23989 (N_23989,N_22963,N_23336);
xnor U23990 (N_23990,N_23317,N_23346);
nand U23991 (N_23991,N_23271,N_22837);
xnor U23992 (N_23992,N_22883,N_22879);
and U23993 (N_23993,N_23294,N_23066);
nor U23994 (N_23994,N_23302,N_22844);
xnor U23995 (N_23995,N_23392,N_22953);
or U23996 (N_23996,N_23204,N_23040);
and U23997 (N_23997,N_22947,N_23039);
nor U23998 (N_23998,N_22849,N_22807);
xnor U23999 (N_23999,N_23215,N_23332);
or U24000 (N_24000,N_23506,N_23975);
nand U24001 (N_24001,N_23861,N_23722);
and U24002 (N_24002,N_23782,N_23551);
xnor U24003 (N_24003,N_23442,N_23518);
nand U24004 (N_24004,N_23666,N_23915);
nor U24005 (N_24005,N_23553,N_23717);
nand U24006 (N_24006,N_23729,N_23826);
or U24007 (N_24007,N_23953,N_23626);
or U24008 (N_24008,N_23605,N_23445);
xor U24009 (N_24009,N_23471,N_23950);
and U24010 (N_24010,N_23929,N_23791);
nand U24011 (N_24011,N_23455,N_23721);
nand U24012 (N_24012,N_23832,N_23916);
and U24013 (N_24013,N_23744,N_23831);
nand U24014 (N_24014,N_23994,N_23519);
xnor U24015 (N_24015,N_23704,N_23575);
nor U24016 (N_24016,N_23673,N_23650);
nand U24017 (N_24017,N_23614,N_23503);
xnor U24018 (N_24018,N_23663,N_23612);
and U24019 (N_24019,N_23625,N_23909);
nor U24020 (N_24020,N_23576,N_23829);
xor U24021 (N_24021,N_23657,N_23680);
nor U24022 (N_24022,N_23429,N_23895);
nand U24023 (N_24023,N_23528,N_23745);
nand U24024 (N_24024,N_23815,N_23993);
nor U24025 (N_24025,N_23533,N_23646);
nor U24026 (N_24026,N_23858,N_23902);
nand U24027 (N_24027,N_23504,N_23874);
nor U24028 (N_24028,N_23498,N_23522);
nor U24029 (N_24029,N_23869,N_23784);
nor U24030 (N_24030,N_23502,N_23919);
nand U24031 (N_24031,N_23572,N_23496);
xor U24032 (N_24032,N_23427,N_23542);
xor U24033 (N_24033,N_23509,N_23788);
and U24034 (N_24034,N_23698,N_23821);
nor U24035 (N_24035,N_23860,N_23561);
nor U24036 (N_24036,N_23819,N_23571);
nand U24037 (N_24037,N_23403,N_23736);
xnor U24038 (N_24038,N_23598,N_23996);
and U24039 (N_24039,N_23497,N_23662);
nor U24040 (N_24040,N_23567,N_23664);
nor U24041 (N_24041,N_23412,N_23825);
and U24042 (N_24042,N_23488,N_23627);
nor U24043 (N_24043,N_23417,N_23456);
xor U24044 (N_24044,N_23921,N_23775);
xnor U24045 (N_24045,N_23402,N_23990);
nand U24046 (N_24046,N_23846,N_23405);
and U24047 (N_24047,N_23547,N_23521);
xor U24048 (N_24048,N_23726,N_23817);
xnor U24049 (N_24049,N_23885,N_23763);
or U24050 (N_24050,N_23751,N_23806);
and U24051 (N_24051,N_23952,N_23780);
or U24052 (N_24052,N_23678,N_23524);
nand U24053 (N_24053,N_23448,N_23894);
nor U24054 (N_24054,N_23684,N_23801);
nand U24055 (N_24055,N_23623,N_23406);
nand U24056 (N_24056,N_23688,N_23823);
and U24057 (N_24057,N_23499,N_23741);
nor U24058 (N_24058,N_23491,N_23712);
or U24059 (N_24059,N_23911,N_23809);
nor U24060 (N_24060,N_23987,N_23934);
or U24061 (N_24061,N_23495,N_23844);
or U24062 (N_24062,N_23527,N_23771);
and U24063 (N_24063,N_23776,N_23976);
and U24064 (N_24064,N_23848,N_23629);
nor U24065 (N_24065,N_23907,N_23563);
xor U24066 (N_24066,N_23798,N_23581);
xnor U24067 (N_24067,N_23743,N_23882);
or U24068 (N_24068,N_23834,N_23557);
xor U24069 (N_24069,N_23609,N_23449);
nand U24070 (N_24070,N_23638,N_23615);
nand U24071 (N_24071,N_23592,N_23492);
nor U24072 (N_24072,N_23989,N_23520);
xnor U24073 (N_24073,N_23415,N_23400);
or U24074 (N_24074,N_23851,N_23728);
nor U24075 (N_24075,N_23622,N_23774);
nor U24076 (N_24076,N_23749,N_23768);
or U24077 (N_24077,N_23924,N_23710);
nor U24078 (N_24078,N_23997,N_23893);
and U24079 (N_24079,N_23446,N_23683);
xnor U24080 (N_24080,N_23578,N_23886);
or U24081 (N_24081,N_23409,N_23473);
or U24082 (N_24082,N_23792,N_23946);
or U24083 (N_24083,N_23554,N_23912);
xor U24084 (N_24084,N_23984,N_23900);
nor U24085 (N_24085,N_23611,N_23787);
nor U24086 (N_24086,N_23765,N_23595);
or U24087 (N_24087,N_23873,N_23905);
xnor U24088 (N_24088,N_23640,N_23725);
and U24089 (N_24089,N_23936,N_23884);
or U24090 (N_24090,N_23670,N_23930);
nor U24091 (N_24091,N_23632,N_23720);
and U24092 (N_24092,N_23866,N_23980);
xor U24093 (N_24093,N_23805,N_23906);
or U24094 (N_24094,N_23653,N_23943);
and U24095 (N_24095,N_23904,N_23702);
xnor U24096 (N_24096,N_23671,N_23661);
xor U24097 (N_24097,N_23730,N_23515);
nor U24098 (N_24098,N_23843,N_23485);
xnor U24099 (N_24099,N_23480,N_23539);
or U24100 (N_24100,N_23752,N_23549);
nor U24101 (N_24101,N_23419,N_23922);
or U24102 (N_24102,N_23742,N_23878);
or U24103 (N_24103,N_23816,N_23418);
xnor U24104 (N_24104,N_23478,N_23501);
xor U24105 (N_24105,N_23458,N_23401);
and U24106 (N_24106,N_23476,N_23979);
nor U24107 (N_24107,N_23613,N_23773);
or U24108 (N_24108,N_23847,N_23457);
and U24109 (N_24109,N_23967,N_23735);
nor U24110 (N_24110,N_23971,N_23562);
or U24111 (N_24111,N_23525,N_23777);
xor U24112 (N_24112,N_23982,N_23969);
and U24113 (N_24113,N_23795,N_23530);
nor U24114 (N_24114,N_23838,N_23796);
nand U24115 (N_24115,N_23845,N_23948);
or U24116 (N_24116,N_23697,N_23414);
xor U24117 (N_24117,N_23477,N_23700);
and U24118 (N_24118,N_23966,N_23802);
or U24119 (N_24119,N_23510,N_23639);
xnor U24120 (N_24120,N_23746,N_23507);
xor U24121 (N_24121,N_23668,N_23451);
nor U24122 (N_24122,N_23674,N_23991);
nor U24123 (N_24123,N_23901,N_23514);
xor U24124 (N_24124,N_23660,N_23753);
or U24125 (N_24125,N_23600,N_23956);
nand U24126 (N_24126,N_23422,N_23596);
nor U24127 (N_24127,N_23871,N_23876);
xnor U24128 (N_24128,N_23459,N_23965);
or U24129 (N_24129,N_23694,N_23783);
nor U24130 (N_24130,N_23853,N_23913);
nand U24131 (N_24131,N_23636,N_23556);
or U24132 (N_24132,N_23849,N_23747);
xor U24133 (N_24133,N_23416,N_23460);
xnor U24134 (N_24134,N_23835,N_23691);
or U24135 (N_24135,N_23526,N_23941);
and U24136 (N_24136,N_23964,N_23610);
xor U24137 (N_24137,N_23441,N_23779);
xor U24138 (N_24138,N_23426,N_23590);
or U24139 (N_24139,N_23597,N_23675);
and U24140 (N_24140,N_23865,N_23789);
nand U24141 (N_24141,N_23814,N_23824);
or U24142 (N_24142,N_23651,N_23830);
nand U24143 (N_24143,N_23437,N_23920);
and U24144 (N_24144,N_23669,N_23642);
nand U24145 (N_24145,N_23641,N_23833);
or U24146 (N_24146,N_23879,N_23601);
nand U24147 (N_24147,N_23881,N_23617);
or U24148 (N_24148,N_23727,N_23404);
nand U24149 (N_24149,N_23750,N_23452);
and U24150 (N_24150,N_23568,N_23479);
nand U24151 (N_24151,N_23778,N_23564);
or U24152 (N_24152,N_23579,N_23433);
nor U24153 (N_24153,N_23794,N_23942);
xnor U24154 (N_24154,N_23544,N_23486);
xor U24155 (N_24155,N_23888,N_23555);
xnor U24156 (N_24156,N_23493,N_23469);
and U24157 (N_24157,N_23490,N_23608);
nor U24158 (N_24158,N_23864,N_23762);
nor U24159 (N_24159,N_23587,N_23465);
nor U24160 (N_24160,N_23511,N_23933);
xnor U24161 (N_24161,N_23820,N_23439);
nand U24162 (N_24162,N_23899,N_23961);
and U24163 (N_24163,N_23628,N_23450);
nand U24164 (N_24164,N_23890,N_23583);
xor U24165 (N_24165,N_23529,N_23467);
and U24166 (N_24166,N_23665,N_23548);
xor U24167 (N_24167,N_23654,N_23786);
and U24168 (N_24168,N_23803,N_23558);
nor U24169 (N_24169,N_23420,N_23538);
or U24170 (N_24170,N_23546,N_23925);
nor U24171 (N_24171,N_23444,N_23540);
xor U24172 (N_24172,N_23822,N_23755);
nand U24173 (N_24173,N_23594,N_23436);
nand U24174 (N_24174,N_23647,N_23903);
nand U24175 (N_24175,N_23602,N_23928);
nand U24176 (N_24176,N_23767,N_23580);
and U24177 (N_24177,N_23689,N_23701);
and U24178 (N_24178,N_23593,N_23523);
and U24179 (N_24179,N_23474,N_23868);
or U24180 (N_24180,N_23607,N_23644);
and U24181 (N_24181,N_23472,N_23734);
nand U24182 (N_24182,N_23937,N_23574);
or U24183 (N_24183,N_23740,N_23896);
xor U24184 (N_24184,N_23716,N_23897);
xor U24185 (N_24185,N_23986,N_23703);
nor U24186 (N_24186,N_23854,N_23807);
and U24187 (N_24187,N_23857,N_23944);
and U24188 (N_24188,N_23517,N_23483);
nor U24189 (N_24189,N_23962,N_23475);
xnor U24190 (N_24190,N_23758,N_23582);
xor U24191 (N_24191,N_23672,N_23793);
nor U24192 (N_24192,N_23978,N_23696);
xnor U24193 (N_24193,N_23938,N_23863);
xor U24194 (N_24194,N_23484,N_23923);
and U24195 (N_24195,N_23932,N_23959);
xor U24196 (N_24196,N_23659,N_23466);
and U24197 (N_24197,N_23705,N_23756);
nand U24198 (N_24198,N_23769,N_23431);
or U24199 (N_24199,N_23677,N_23761);
nand U24200 (N_24200,N_23588,N_23434);
and U24201 (N_24201,N_23898,N_23870);
nand U24202 (N_24202,N_23718,N_23839);
and U24203 (N_24203,N_23430,N_23685);
and U24204 (N_24204,N_23892,N_23828);
nand U24205 (N_24205,N_23440,N_23781);
xor U24206 (N_24206,N_23770,N_23604);
or U24207 (N_24207,N_23494,N_23958);
nor U24208 (N_24208,N_23827,N_23877);
and U24209 (N_24209,N_23655,N_23949);
nand U24210 (N_24210,N_23812,N_23424);
and U24211 (N_24211,N_23891,N_23408);
nand U24212 (N_24212,N_23957,N_23545);
and U24213 (N_24213,N_23453,N_23960);
nor U24214 (N_24214,N_23732,N_23852);
or U24215 (N_24215,N_23840,N_23482);
nor U24216 (N_24216,N_23800,N_23714);
and U24217 (N_24217,N_23589,N_23468);
and U24218 (N_24218,N_23463,N_23707);
nor U24219 (N_24219,N_23624,N_23713);
xor U24220 (N_24220,N_23676,N_23447);
xor U24221 (N_24221,N_23766,N_23813);
and U24222 (N_24222,N_23682,N_23918);
nor U24223 (N_24223,N_23799,N_23850);
nand U24224 (N_24224,N_23679,N_23591);
nor U24225 (N_24225,N_23737,N_23738);
nand U24226 (N_24226,N_23516,N_23648);
nor U24227 (N_24227,N_23867,N_23945);
and U24228 (N_24228,N_23470,N_23811);
nand U24229 (N_24229,N_23926,N_23724);
or U24230 (N_24230,N_23790,N_23739);
nor U24231 (N_24231,N_23837,N_23603);
xnor U24232 (N_24232,N_23706,N_23570);
and U24233 (N_24233,N_23686,N_23748);
nor U24234 (N_24234,N_23508,N_23972);
or U24235 (N_24235,N_23454,N_23500);
nand U24236 (N_24236,N_23637,N_23939);
and U24237 (N_24237,N_23534,N_23425);
xnor U24238 (N_24238,N_23645,N_23550);
nand U24239 (N_24239,N_23974,N_23772);
nor U24240 (N_24240,N_23955,N_23573);
or U24241 (N_24241,N_23977,N_23818);
nand U24242 (N_24242,N_23423,N_23649);
and U24243 (N_24243,N_23889,N_23487);
and U24244 (N_24244,N_23859,N_23887);
xor U24245 (N_24245,N_23631,N_23757);
or U24246 (N_24246,N_23428,N_23620);
nand U24247 (N_24247,N_23633,N_23692);
or U24248 (N_24248,N_23935,N_23875);
nor U24249 (N_24249,N_23566,N_23656);
and U24250 (N_24250,N_23658,N_23855);
and U24251 (N_24251,N_23585,N_23715);
nor U24252 (N_24252,N_23856,N_23764);
or U24253 (N_24253,N_23719,N_23759);
or U24254 (N_24254,N_23541,N_23513);
nand U24255 (N_24255,N_23917,N_23931);
xnor U24256 (N_24256,N_23634,N_23914);
and U24257 (N_24257,N_23543,N_23635);
nand U24258 (N_24258,N_23785,N_23970);
xnor U24259 (N_24259,N_23565,N_23995);
or U24260 (N_24260,N_23951,N_23973);
and U24261 (N_24261,N_23810,N_23586);
nand U24262 (N_24262,N_23532,N_23432);
nand U24263 (N_24263,N_23841,N_23940);
nor U24264 (N_24264,N_23733,N_23981);
and U24265 (N_24265,N_23968,N_23699);
nor U24266 (N_24266,N_23411,N_23693);
and U24267 (N_24267,N_23435,N_23687);
and U24268 (N_24268,N_23690,N_23992);
nand U24269 (N_24269,N_23711,N_23443);
and U24270 (N_24270,N_23535,N_23883);
or U24271 (N_24271,N_23695,N_23606);
or U24272 (N_24272,N_23808,N_23667);
nor U24273 (N_24273,N_23464,N_23862);
nor U24274 (N_24274,N_23407,N_23621);
and U24275 (N_24275,N_23618,N_23709);
nand U24276 (N_24276,N_23910,N_23512);
nand U24277 (N_24277,N_23998,N_23643);
or U24278 (N_24278,N_23954,N_23413);
xor U24279 (N_24279,N_23754,N_23531);
nor U24280 (N_24280,N_23481,N_23560);
and U24281 (N_24281,N_23630,N_23537);
nor U24282 (N_24282,N_23927,N_23908);
and U24283 (N_24283,N_23505,N_23797);
xnor U24284 (N_24284,N_23760,N_23681);
nand U24285 (N_24285,N_23880,N_23584);
nand U24286 (N_24286,N_23461,N_23804);
xnor U24287 (N_24287,N_23999,N_23462);
or U24288 (N_24288,N_23410,N_23872);
xor U24289 (N_24289,N_23489,N_23983);
xnor U24290 (N_24290,N_23731,N_23963);
or U24291 (N_24291,N_23988,N_23836);
nand U24292 (N_24292,N_23569,N_23438);
xnor U24293 (N_24293,N_23842,N_23619);
or U24294 (N_24294,N_23599,N_23616);
xor U24295 (N_24295,N_23559,N_23985);
nor U24296 (N_24296,N_23652,N_23723);
and U24297 (N_24297,N_23536,N_23708);
or U24298 (N_24298,N_23947,N_23552);
and U24299 (N_24299,N_23577,N_23421);
and U24300 (N_24300,N_23416,N_23607);
and U24301 (N_24301,N_23987,N_23707);
and U24302 (N_24302,N_23537,N_23886);
and U24303 (N_24303,N_23818,N_23420);
nor U24304 (N_24304,N_23695,N_23458);
and U24305 (N_24305,N_23990,N_23686);
nand U24306 (N_24306,N_23748,N_23852);
xnor U24307 (N_24307,N_23779,N_23910);
nor U24308 (N_24308,N_23483,N_23629);
or U24309 (N_24309,N_23877,N_23844);
and U24310 (N_24310,N_23693,N_23448);
and U24311 (N_24311,N_23990,N_23710);
and U24312 (N_24312,N_23777,N_23564);
xor U24313 (N_24313,N_23531,N_23781);
xor U24314 (N_24314,N_23895,N_23749);
and U24315 (N_24315,N_23879,N_23813);
or U24316 (N_24316,N_23995,N_23914);
xnor U24317 (N_24317,N_23670,N_23435);
nand U24318 (N_24318,N_23643,N_23646);
or U24319 (N_24319,N_23590,N_23696);
or U24320 (N_24320,N_23496,N_23810);
nor U24321 (N_24321,N_23877,N_23946);
and U24322 (N_24322,N_23750,N_23885);
and U24323 (N_24323,N_23763,N_23827);
nand U24324 (N_24324,N_23816,N_23540);
nor U24325 (N_24325,N_23687,N_23777);
xor U24326 (N_24326,N_23472,N_23502);
nand U24327 (N_24327,N_23448,N_23902);
nor U24328 (N_24328,N_23587,N_23737);
xnor U24329 (N_24329,N_23762,N_23834);
xor U24330 (N_24330,N_23624,N_23662);
xnor U24331 (N_24331,N_23403,N_23925);
and U24332 (N_24332,N_23887,N_23977);
or U24333 (N_24333,N_23614,N_23730);
xor U24334 (N_24334,N_23598,N_23556);
or U24335 (N_24335,N_23666,N_23839);
nor U24336 (N_24336,N_23510,N_23925);
or U24337 (N_24337,N_23558,N_23787);
xor U24338 (N_24338,N_23840,N_23887);
or U24339 (N_24339,N_23554,N_23955);
and U24340 (N_24340,N_23433,N_23839);
nand U24341 (N_24341,N_23792,N_23764);
nand U24342 (N_24342,N_23945,N_23730);
nand U24343 (N_24343,N_23575,N_23697);
nor U24344 (N_24344,N_23926,N_23955);
or U24345 (N_24345,N_23451,N_23743);
and U24346 (N_24346,N_23961,N_23971);
or U24347 (N_24347,N_23764,N_23409);
or U24348 (N_24348,N_23705,N_23732);
xor U24349 (N_24349,N_23693,N_23558);
xnor U24350 (N_24350,N_23500,N_23513);
nor U24351 (N_24351,N_23614,N_23677);
or U24352 (N_24352,N_23467,N_23553);
or U24353 (N_24353,N_23674,N_23681);
and U24354 (N_24354,N_23615,N_23746);
xor U24355 (N_24355,N_23484,N_23821);
or U24356 (N_24356,N_23479,N_23406);
and U24357 (N_24357,N_23409,N_23940);
or U24358 (N_24358,N_23487,N_23944);
xor U24359 (N_24359,N_23669,N_23412);
nor U24360 (N_24360,N_23778,N_23809);
nor U24361 (N_24361,N_23495,N_23742);
and U24362 (N_24362,N_23786,N_23697);
xor U24363 (N_24363,N_23851,N_23689);
nor U24364 (N_24364,N_23981,N_23980);
or U24365 (N_24365,N_23618,N_23830);
and U24366 (N_24366,N_23915,N_23605);
and U24367 (N_24367,N_23604,N_23809);
xnor U24368 (N_24368,N_23540,N_23956);
xnor U24369 (N_24369,N_23843,N_23774);
and U24370 (N_24370,N_23585,N_23872);
nor U24371 (N_24371,N_23943,N_23558);
nand U24372 (N_24372,N_23987,N_23692);
xor U24373 (N_24373,N_23536,N_23661);
nand U24374 (N_24374,N_23497,N_23893);
nand U24375 (N_24375,N_23542,N_23480);
xnor U24376 (N_24376,N_23452,N_23922);
nand U24377 (N_24377,N_23666,N_23884);
or U24378 (N_24378,N_23613,N_23562);
nor U24379 (N_24379,N_23942,N_23691);
or U24380 (N_24380,N_23811,N_23410);
and U24381 (N_24381,N_23785,N_23746);
and U24382 (N_24382,N_23601,N_23931);
and U24383 (N_24383,N_23730,N_23660);
xor U24384 (N_24384,N_23882,N_23788);
or U24385 (N_24385,N_23781,N_23819);
nand U24386 (N_24386,N_23598,N_23616);
or U24387 (N_24387,N_23682,N_23467);
nor U24388 (N_24388,N_23635,N_23416);
or U24389 (N_24389,N_23999,N_23979);
xor U24390 (N_24390,N_23483,N_23487);
nor U24391 (N_24391,N_23591,N_23917);
and U24392 (N_24392,N_23648,N_23551);
nand U24393 (N_24393,N_23713,N_23704);
or U24394 (N_24394,N_23990,N_23905);
xor U24395 (N_24395,N_23539,N_23705);
xor U24396 (N_24396,N_23950,N_23652);
and U24397 (N_24397,N_23510,N_23597);
or U24398 (N_24398,N_23645,N_23544);
and U24399 (N_24399,N_23493,N_23940);
nor U24400 (N_24400,N_23745,N_23436);
or U24401 (N_24401,N_23910,N_23709);
nand U24402 (N_24402,N_23474,N_23880);
nand U24403 (N_24403,N_23595,N_23599);
nor U24404 (N_24404,N_23651,N_23528);
and U24405 (N_24405,N_23821,N_23925);
nand U24406 (N_24406,N_23951,N_23671);
xor U24407 (N_24407,N_23914,N_23461);
and U24408 (N_24408,N_23730,N_23529);
nor U24409 (N_24409,N_23691,N_23839);
and U24410 (N_24410,N_23881,N_23994);
nor U24411 (N_24411,N_23555,N_23672);
and U24412 (N_24412,N_23646,N_23863);
nor U24413 (N_24413,N_23837,N_23628);
nor U24414 (N_24414,N_23560,N_23988);
or U24415 (N_24415,N_23854,N_23441);
nand U24416 (N_24416,N_23521,N_23749);
xnor U24417 (N_24417,N_23573,N_23999);
nand U24418 (N_24418,N_23743,N_23987);
and U24419 (N_24419,N_23952,N_23936);
xor U24420 (N_24420,N_23413,N_23706);
nand U24421 (N_24421,N_23797,N_23567);
nand U24422 (N_24422,N_23810,N_23688);
and U24423 (N_24423,N_23675,N_23486);
and U24424 (N_24424,N_23678,N_23854);
xnor U24425 (N_24425,N_23654,N_23627);
xor U24426 (N_24426,N_23529,N_23608);
xor U24427 (N_24427,N_23722,N_23652);
or U24428 (N_24428,N_23572,N_23847);
or U24429 (N_24429,N_23699,N_23510);
or U24430 (N_24430,N_23755,N_23617);
nand U24431 (N_24431,N_23844,N_23595);
xor U24432 (N_24432,N_23913,N_23652);
nand U24433 (N_24433,N_23747,N_23649);
nor U24434 (N_24434,N_23600,N_23837);
nand U24435 (N_24435,N_23721,N_23758);
and U24436 (N_24436,N_23862,N_23707);
and U24437 (N_24437,N_23716,N_23752);
nor U24438 (N_24438,N_23743,N_23669);
nand U24439 (N_24439,N_23512,N_23476);
nor U24440 (N_24440,N_23415,N_23425);
nor U24441 (N_24441,N_23716,N_23687);
and U24442 (N_24442,N_23760,N_23890);
or U24443 (N_24443,N_23835,N_23784);
and U24444 (N_24444,N_23880,N_23647);
nand U24445 (N_24445,N_23589,N_23550);
or U24446 (N_24446,N_23725,N_23678);
nor U24447 (N_24447,N_23446,N_23481);
nor U24448 (N_24448,N_23862,N_23417);
nor U24449 (N_24449,N_23706,N_23653);
xnor U24450 (N_24450,N_23915,N_23939);
nand U24451 (N_24451,N_23830,N_23837);
and U24452 (N_24452,N_23723,N_23900);
nand U24453 (N_24453,N_23683,N_23866);
and U24454 (N_24454,N_23543,N_23964);
xnor U24455 (N_24455,N_23721,N_23703);
xor U24456 (N_24456,N_23500,N_23614);
xor U24457 (N_24457,N_23409,N_23675);
nor U24458 (N_24458,N_23848,N_23809);
and U24459 (N_24459,N_23515,N_23908);
and U24460 (N_24460,N_23581,N_23401);
xor U24461 (N_24461,N_23951,N_23648);
nor U24462 (N_24462,N_23472,N_23424);
nor U24463 (N_24463,N_23532,N_23431);
and U24464 (N_24464,N_23554,N_23542);
xnor U24465 (N_24465,N_23497,N_23614);
nand U24466 (N_24466,N_23428,N_23821);
nor U24467 (N_24467,N_23499,N_23575);
xor U24468 (N_24468,N_23419,N_23499);
xnor U24469 (N_24469,N_23644,N_23695);
xor U24470 (N_24470,N_23721,N_23887);
nor U24471 (N_24471,N_23969,N_23501);
and U24472 (N_24472,N_23619,N_23520);
nand U24473 (N_24473,N_23408,N_23697);
nand U24474 (N_24474,N_23474,N_23679);
nor U24475 (N_24475,N_23914,N_23890);
or U24476 (N_24476,N_23453,N_23840);
xnor U24477 (N_24477,N_23997,N_23683);
nand U24478 (N_24478,N_23987,N_23416);
and U24479 (N_24479,N_23814,N_23503);
or U24480 (N_24480,N_23762,N_23774);
nor U24481 (N_24481,N_23651,N_23985);
and U24482 (N_24482,N_23542,N_23920);
or U24483 (N_24483,N_23858,N_23890);
nand U24484 (N_24484,N_23721,N_23648);
or U24485 (N_24485,N_23470,N_23905);
xor U24486 (N_24486,N_23935,N_23458);
and U24487 (N_24487,N_23848,N_23733);
nand U24488 (N_24488,N_23748,N_23408);
nor U24489 (N_24489,N_23421,N_23454);
or U24490 (N_24490,N_23854,N_23962);
nor U24491 (N_24491,N_23775,N_23769);
and U24492 (N_24492,N_23620,N_23539);
nand U24493 (N_24493,N_23655,N_23731);
nor U24494 (N_24494,N_23417,N_23827);
and U24495 (N_24495,N_23808,N_23638);
or U24496 (N_24496,N_23965,N_23423);
or U24497 (N_24497,N_23572,N_23581);
and U24498 (N_24498,N_23970,N_23617);
or U24499 (N_24499,N_23484,N_23464);
or U24500 (N_24500,N_23496,N_23593);
nand U24501 (N_24501,N_23970,N_23754);
nor U24502 (N_24502,N_23884,N_23493);
and U24503 (N_24503,N_23921,N_23455);
and U24504 (N_24504,N_23678,N_23567);
nor U24505 (N_24505,N_23774,N_23440);
or U24506 (N_24506,N_23799,N_23511);
and U24507 (N_24507,N_23673,N_23607);
nand U24508 (N_24508,N_23869,N_23546);
nand U24509 (N_24509,N_23887,N_23517);
nand U24510 (N_24510,N_23771,N_23959);
and U24511 (N_24511,N_23752,N_23758);
or U24512 (N_24512,N_23812,N_23504);
and U24513 (N_24513,N_23541,N_23530);
nand U24514 (N_24514,N_23888,N_23765);
or U24515 (N_24515,N_23463,N_23736);
xnor U24516 (N_24516,N_23648,N_23595);
xor U24517 (N_24517,N_23828,N_23884);
and U24518 (N_24518,N_23517,N_23864);
xnor U24519 (N_24519,N_23453,N_23792);
nor U24520 (N_24520,N_23916,N_23778);
or U24521 (N_24521,N_23869,N_23637);
nand U24522 (N_24522,N_23903,N_23682);
xnor U24523 (N_24523,N_23934,N_23900);
nor U24524 (N_24524,N_23895,N_23915);
and U24525 (N_24525,N_23803,N_23423);
nor U24526 (N_24526,N_23742,N_23617);
and U24527 (N_24527,N_23585,N_23833);
and U24528 (N_24528,N_23860,N_23684);
or U24529 (N_24529,N_23825,N_23821);
and U24530 (N_24530,N_23728,N_23418);
nand U24531 (N_24531,N_23528,N_23644);
nor U24532 (N_24532,N_23993,N_23529);
xnor U24533 (N_24533,N_23987,N_23818);
nand U24534 (N_24534,N_23855,N_23586);
xnor U24535 (N_24535,N_23803,N_23897);
nand U24536 (N_24536,N_23922,N_23875);
nor U24537 (N_24537,N_23523,N_23866);
nor U24538 (N_24538,N_23917,N_23418);
nor U24539 (N_24539,N_23579,N_23967);
and U24540 (N_24540,N_23944,N_23848);
or U24541 (N_24541,N_23536,N_23415);
or U24542 (N_24542,N_23552,N_23511);
or U24543 (N_24543,N_23447,N_23462);
nand U24544 (N_24544,N_23677,N_23833);
nand U24545 (N_24545,N_23894,N_23625);
nor U24546 (N_24546,N_23438,N_23972);
nand U24547 (N_24547,N_23966,N_23595);
nand U24548 (N_24548,N_23984,N_23723);
xnor U24549 (N_24549,N_23778,N_23851);
or U24550 (N_24550,N_23989,N_23598);
nor U24551 (N_24551,N_23921,N_23668);
nand U24552 (N_24552,N_23718,N_23550);
xor U24553 (N_24553,N_23988,N_23802);
or U24554 (N_24554,N_23598,N_23600);
and U24555 (N_24555,N_23903,N_23759);
and U24556 (N_24556,N_23643,N_23754);
nand U24557 (N_24557,N_23691,N_23626);
xor U24558 (N_24558,N_23487,N_23892);
nor U24559 (N_24559,N_23795,N_23655);
xor U24560 (N_24560,N_23732,N_23940);
nand U24561 (N_24561,N_23875,N_23700);
xnor U24562 (N_24562,N_23830,N_23984);
xnor U24563 (N_24563,N_23912,N_23752);
or U24564 (N_24564,N_23704,N_23404);
nor U24565 (N_24565,N_23718,N_23783);
and U24566 (N_24566,N_23621,N_23677);
nor U24567 (N_24567,N_23614,N_23458);
nand U24568 (N_24568,N_23501,N_23780);
xnor U24569 (N_24569,N_23992,N_23720);
or U24570 (N_24570,N_23511,N_23562);
xor U24571 (N_24571,N_23852,N_23725);
xor U24572 (N_24572,N_23494,N_23609);
and U24573 (N_24573,N_23814,N_23722);
and U24574 (N_24574,N_23541,N_23637);
nand U24575 (N_24575,N_23862,N_23532);
or U24576 (N_24576,N_23912,N_23568);
nand U24577 (N_24577,N_23457,N_23601);
and U24578 (N_24578,N_23410,N_23549);
nand U24579 (N_24579,N_23757,N_23592);
nor U24580 (N_24580,N_23818,N_23709);
nor U24581 (N_24581,N_23761,N_23445);
xnor U24582 (N_24582,N_23917,N_23516);
nor U24583 (N_24583,N_23865,N_23565);
xor U24584 (N_24584,N_23435,N_23433);
and U24585 (N_24585,N_23990,N_23494);
nand U24586 (N_24586,N_23498,N_23699);
xor U24587 (N_24587,N_23449,N_23736);
nor U24588 (N_24588,N_23403,N_23472);
nand U24589 (N_24589,N_23633,N_23642);
nand U24590 (N_24590,N_23447,N_23518);
nand U24591 (N_24591,N_23449,N_23581);
nor U24592 (N_24592,N_23610,N_23905);
nand U24593 (N_24593,N_23679,N_23484);
nand U24594 (N_24594,N_23706,N_23887);
nor U24595 (N_24595,N_23982,N_23400);
nand U24596 (N_24596,N_23473,N_23579);
or U24597 (N_24597,N_23513,N_23770);
and U24598 (N_24598,N_23649,N_23402);
nand U24599 (N_24599,N_23510,N_23908);
nand U24600 (N_24600,N_24525,N_24217);
nor U24601 (N_24601,N_24037,N_24385);
xnor U24602 (N_24602,N_24076,N_24289);
nand U24603 (N_24603,N_24365,N_24391);
xnor U24604 (N_24604,N_24084,N_24535);
or U24605 (N_24605,N_24098,N_24512);
nand U24606 (N_24606,N_24269,N_24077);
or U24607 (N_24607,N_24061,N_24344);
nor U24608 (N_24608,N_24260,N_24233);
or U24609 (N_24609,N_24250,N_24405);
nand U24610 (N_24610,N_24090,N_24430);
nor U24611 (N_24611,N_24219,N_24422);
nor U24612 (N_24612,N_24479,N_24075);
xnor U24613 (N_24613,N_24205,N_24304);
nor U24614 (N_24614,N_24068,N_24369);
nand U24615 (N_24615,N_24312,N_24243);
nor U24616 (N_24616,N_24033,N_24401);
or U24617 (N_24617,N_24332,N_24336);
or U24618 (N_24618,N_24018,N_24026);
nor U24619 (N_24619,N_24253,N_24297);
xor U24620 (N_24620,N_24557,N_24105);
nand U24621 (N_24621,N_24270,N_24381);
or U24622 (N_24622,N_24361,N_24360);
nand U24623 (N_24623,N_24490,N_24318);
or U24624 (N_24624,N_24393,N_24330);
nand U24625 (N_24625,N_24252,N_24514);
nand U24626 (N_24626,N_24131,N_24508);
and U24627 (N_24627,N_24325,N_24496);
nor U24628 (N_24628,N_24106,N_24346);
or U24629 (N_24629,N_24153,N_24129);
nand U24630 (N_24630,N_24211,N_24301);
or U24631 (N_24631,N_24409,N_24091);
nand U24632 (N_24632,N_24340,N_24449);
or U24633 (N_24633,N_24463,N_24442);
or U24634 (N_24634,N_24158,N_24287);
nor U24635 (N_24635,N_24335,N_24276);
and U24636 (N_24636,N_24014,N_24057);
and U24637 (N_24637,N_24394,N_24314);
nor U24638 (N_24638,N_24487,N_24049);
and U24639 (N_24639,N_24196,N_24238);
nor U24640 (N_24640,N_24371,N_24085);
nor U24641 (N_24641,N_24558,N_24109);
nor U24642 (N_24642,N_24152,N_24598);
nand U24643 (N_24643,N_24323,N_24311);
xnor U24644 (N_24644,N_24413,N_24310);
or U24645 (N_24645,N_24100,N_24114);
nor U24646 (N_24646,N_24221,N_24435);
nor U24647 (N_24647,N_24563,N_24599);
nor U24648 (N_24648,N_24283,N_24144);
or U24649 (N_24649,N_24454,N_24506);
and U24650 (N_24650,N_24389,N_24142);
or U24651 (N_24651,N_24458,N_24082);
and U24652 (N_24652,N_24171,N_24298);
nor U24653 (N_24653,N_24457,N_24333);
nand U24654 (N_24654,N_24583,N_24550);
nor U24655 (N_24655,N_24438,N_24482);
or U24656 (N_24656,N_24302,N_24559);
or U24657 (N_24657,N_24505,N_24532);
or U24658 (N_24658,N_24553,N_24414);
xnor U24659 (N_24659,N_24571,N_24154);
nor U24660 (N_24660,N_24198,N_24272);
nand U24661 (N_24661,N_24005,N_24140);
nand U24662 (N_24662,N_24516,N_24281);
nor U24663 (N_24663,N_24284,N_24519);
nand U24664 (N_24664,N_24088,N_24223);
or U24665 (N_24665,N_24426,N_24429);
nor U24666 (N_24666,N_24072,N_24275);
xor U24667 (N_24667,N_24596,N_24481);
or U24668 (N_24668,N_24296,N_24132);
xnor U24669 (N_24669,N_24498,N_24007);
nand U24670 (N_24670,N_24038,N_24578);
or U24671 (N_24671,N_24212,N_24143);
and U24672 (N_24672,N_24087,N_24161);
nor U24673 (N_24673,N_24273,N_24588);
xnor U24674 (N_24674,N_24064,N_24373);
nor U24675 (N_24675,N_24010,N_24130);
nor U24676 (N_24676,N_24338,N_24199);
xnor U24677 (N_24677,N_24056,N_24254);
and U24678 (N_24678,N_24006,N_24565);
nor U24679 (N_24679,N_24263,N_24448);
and U24680 (N_24680,N_24515,N_24227);
or U24681 (N_24681,N_24280,N_24025);
or U24682 (N_24682,N_24050,N_24177);
nor U24683 (N_24683,N_24122,N_24326);
nand U24684 (N_24684,N_24447,N_24124);
nand U24685 (N_24685,N_24424,N_24044);
nand U24686 (N_24686,N_24268,N_24180);
and U24687 (N_24687,N_24194,N_24101);
and U24688 (N_24688,N_24020,N_24561);
and U24689 (N_24689,N_24136,N_24059);
nor U24690 (N_24690,N_24523,N_24092);
xnor U24691 (N_24691,N_24484,N_24408);
xor U24692 (N_24692,N_24541,N_24475);
and U24693 (N_24693,N_24051,N_24230);
nand U24694 (N_24694,N_24264,N_24277);
xor U24695 (N_24695,N_24327,N_24045);
and U24696 (N_24696,N_24182,N_24539);
xor U24697 (N_24697,N_24237,N_24313);
and U24698 (N_24698,N_24288,N_24294);
nand U24699 (N_24699,N_24240,N_24507);
nor U24700 (N_24700,N_24522,N_24220);
xnor U24701 (N_24701,N_24444,N_24141);
and U24702 (N_24702,N_24489,N_24582);
nand U24703 (N_24703,N_24485,N_24570);
xnor U24704 (N_24704,N_24402,N_24537);
nor U24705 (N_24705,N_24041,N_24201);
nand U24706 (N_24706,N_24492,N_24104);
nor U24707 (N_24707,N_24034,N_24218);
and U24708 (N_24708,N_24128,N_24229);
and U24709 (N_24709,N_24504,N_24538);
nand U24710 (N_24710,N_24279,N_24554);
or U24711 (N_24711,N_24552,N_24231);
and U24712 (N_24712,N_24543,N_24095);
nand U24713 (N_24713,N_24247,N_24418);
or U24714 (N_24714,N_24303,N_24317);
and U24715 (N_24715,N_24116,N_24590);
or U24716 (N_24716,N_24580,N_24190);
or U24717 (N_24717,N_24255,N_24008);
nor U24718 (N_24718,N_24174,N_24183);
nor U24719 (N_24719,N_24001,N_24145);
nand U24720 (N_24720,N_24494,N_24189);
and U24721 (N_24721,N_24555,N_24094);
or U24722 (N_24722,N_24258,N_24581);
and U24723 (N_24723,N_24486,N_24023);
or U24724 (N_24724,N_24544,N_24052);
nand U24725 (N_24725,N_24388,N_24151);
xor U24726 (N_24726,N_24566,N_24358);
nand U24727 (N_24727,N_24450,N_24383);
nor U24728 (N_24728,N_24035,N_24376);
and U24729 (N_24729,N_24155,N_24356);
xor U24730 (N_24730,N_24173,N_24058);
and U24731 (N_24731,N_24123,N_24337);
nor U24732 (N_24732,N_24493,N_24146);
or U24733 (N_24733,N_24000,N_24043);
and U24734 (N_24734,N_24370,N_24319);
xor U24735 (N_24735,N_24245,N_24591);
xnor U24736 (N_24736,N_24355,N_24572);
or U24737 (N_24737,N_24546,N_24460);
nor U24738 (N_24738,N_24397,N_24593);
and U24739 (N_24739,N_24053,N_24187);
xor U24740 (N_24740,N_24046,N_24529);
nand U24741 (N_24741,N_24165,N_24597);
nand U24742 (N_24742,N_24549,N_24540);
nand U24743 (N_24743,N_24451,N_24455);
nor U24744 (N_24744,N_24467,N_24411);
nand U24745 (N_24745,N_24595,N_24320);
xor U24746 (N_24746,N_24226,N_24133);
nor U24747 (N_24747,N_24291,N_24399);
nor U24748 (N_24748,N_24322,N_24016);
or U24749 (N_24749,N_24178,N_24585);
and U24750 (N_24750,N_24334,N_24586);
and U24751 (N_24751,N_24307,N_24266);
xor U24752 (N_24752,N_24527,N_24465);
or U24753 (N_24753,N_24022,N_24491);
and U24754 (N_24754,N_24012,N_24070);
nand U24755 (N_24755,N_24074,N_24309);
or U24756 (N_24756,N_24040,N_24139);
nor U24757 (N_24757,N_24137,N_24015);
nor U24758 (N_24758,N_24257,N_24267);
xor U24759 (N_24759,N_24054,N_24420);
and U24760 (N_24760,N_24374,N_24531);
xor U24761 (N_24761,N_24021,N_24587);
and U24762 (N_24762,N_24466,N_24042);
or U24763 (N_24763,N_24521,N_24290);
nand U24764 (N_24764,N_24036,N_24501);
nor U24765 (N_24765,N_24511,N_24262);
nor U24766 (N_24766,N_24354,N_24428);
nand U24767 (N_24767,N_24188,N_24031);
or U24768 (N_24768,N_24300,N_24017);
nor U24769 (N_24769,N_24416,N_24500);
xnor U24770 (N_24770,N_24379,N_24019);
xnor U24771 (N_24771,N_24149,N_24147);
nor U24772 (N_24772,N_24202,N_24509);
nand U24773 (N_24773,N_24551,N_24380);
nand U24774 (N_24774,N_24060,N_24499);
or U24775 (N_24775,N_24461,N_24445);
and U24776 (N_24776,N_24436,N_24119);
xor U24777 (N_24777,N_24548,N_24066);
nand U24778 (N_24778,N_24536,N_24404);
and U24779 (N_24779,N_24589,N_24510);
and U24780 (N_24780,N_24160,N_24366);
or U24781 (N_24781,N_24259,N_24339);
xor U24782 (N_24782,N_24362,N_24185);
nor U24783 (N_24783,N_24286,N_24594);
or U24784 (N_24784,N_24179,N_24407);
xnor U24785 (N_24785,N_24278,N_24328);
xor U24786 (N_24786,N_24384,N_24568);
xnor U24787 (N_24787,N_24099,N_24200);
xnor U24788 (N_24788,N_24415,N_24534);
nand U24789 (N_24789,N_24443,N_24175);
or U24790 (N_24790,N_24324,N_24186);
or U24791 (N_24791,N_24047,N_24400);
xnor U24792 (N_24792,N_24004,N_24468);
xor U24793 (N_24793,N_24285,N_24193);
nand U24794 (N_24794,N_24039,N_24347);
xnor U24795 (N_24795,N_24584,N_24476);
nor U24796 (N_24796,N_24163,N_24431);
and U24797 (N_24797,N_24390,N_24156);
nand U24798 (N_24798,N_24111,N_24215);
xor U24799 (N_24799,N_24437,N_24472);
nand U24800 (N_24800,N_24069,N_24197);
nor U24801 (N_24801,N_24299,N_24097);
and U24802 (N_24802,N_24343,N_24392);
xor U24803 (N_24803,N_24209,N_24225);
nand U24804 (N_24804,N_24080,N_24439);
and U24805 (N_24805,N_24478,N_24592);
nand U24806 (N_24806,N_24524,N_24352);
xnor U24807 (N_24807,N_24562,N_24417);
nor U24808 (N_24808,N_24135,N_24192);
nand U24809 (N_24809,N_24024,N_24470);
xor U24810 (N_24810,N_24406,N_24432);
xnor U24811 (N_24811,N_24359,N_24027);
nand U24812 (N_24812,N_24434,N_24526);
xnor U24813 (N_24813,N_24127,N_24030);
nor U24814 (N_24814,N_24134,N_24009);
nand U24815 (N_24815,N_24256,N_24113);
or U24816 (N_24816,N_24533,N_24331);
nand U24817 (N_24817,N_24013,N_24363);
or U24818 (N_24818,N_24184,N_24086);
and U24819 (N_24819,N_24207,N_24028);
and U24820 (N_24820,N_24488,N_24305);
xnor U24821 (N_24821,N_24410,N_24248);
or U24822 (N_24822,N_24232,N_24115);
xor U24823 (N_24823,N_24222,N_24502);
nand U24824 (N_24824,N_24150,N_24452);
xor U24825 (N_24825,N_24308,N_24446);
nor U24826 (N_24826,N_24518,N_24067);
nand U24827 (N_24827,N_24169,N_24003);
or U24828 (N_24828,N_24236,N_24216);
and U24829 (N_24829,N_24469,N_24065);
nand U24830 (N_24830,N_24575,N_24375);
and U24831 (N_24831,N_24306,N_24372);
or U24832 (N_24832,N_24195,N_24377);
and U24833 (N_24833,N_24093,N_24121);
xor U24834 (N_24834,N_24357,N_24483);
xnor U24835 (N_24835,N_24295,N_24471);
xnor U24836 (N_24836,N_24517,N_24459);
and U24837 (N_24837,N_24441,N_24315);
or U24838 (N_24838,N_24118,N_24530);
nand U24839 (N_24839,N_24073,N_24574);
nor U24840 (N_24840,N_24528,N_24261);
nor U24841 (N_24841,N_24395,N_24112);
nand U24842 (N_24842,N_24569,N_24497);
nor U24843 (N_24843,N_24029,N_24235);
xnor U24844 (N_24844,N_24474,N_24148);
and U24845 (N_24845,N_24096,N_24176);
or U24846 (N_24846,N_24208,N_24556);
nor U24847 (N_24847,N_24078,N_24547);
xor U24848 (N_24848,N_24063,N_24398);
and U24849 (N_24849,N_24293,N_24117);
nand U24850 (N_24850,N_24480,N_24513);
or U24851 (N_24851,N_24503,N_24387);
nand U24852 (N_24852,N_24421,N_24079);
xnor U24853 (N_24853,N_24108,N_24081);
and U24854 (N_24854,N_24349,N_24242);
nand U24855 (N_24855,N_24214,N_24239);
xor U24856 (N_24856,N_24126,N_24341);
nor U24857 (N_24857,N_24168,N_24246);
and U24858 (N_24858,N_24321,N_24191);
nand U24859 (N_24859,N_24251,N_24567);
nand U24860 (N_24860,N_24292,N_24364);
or U24861 (N_24861,N_24329,N_24378);
nand U24862 (N_24862,N_24573,N_24213);
and U24863 (N_24863,N_24210,N_24244);
nor U24864 (N_24864,N_24427,N_24206);
nor U24865 (N_24865,N_24576,N_24520);
nor U24866 (N_24866,N_24453,N_24103);
nor U24867 (N_24867,N_24419,N_24167);
nand U24868 (N_24868,N_24159,N_24403);
nand U24869 (N_24869,N_24166,N_24412);
xor U24870 (N_24870,N_24473,N_24110);
nand U24871 (N_24871,N_24316,N_24224);
nor U24872 (N_24872,N_24351,N_24048);
nor U24873 (N_24873,N_24353,N_24120);
xnor U24874 (N_24874,N_24545,N_24440);
xnor U24875 (N_24875,N_24002,N_24579);
xnor U24876 (N_24876,N_24456,N_24350);
and U24877 (N_24877,N_24423,N_24367);
and U24878 (N_24878,N_24348,N_24138);
xor U24879 (N_24879,N_24464,N_24241);
nand U24880 (N_24880,N_24164,N_24560);
or U24881 (N_24881,N_24477,N_24228);
or U24882 (N_24882,N_24234,N_24433);
nor U24883 (N_24883,N_24386,N_24089);
nor U24884 (N_24884,N_24083,N_24382);
and U24885 (N_24885,N_24062,N_24564);
or U24886 (N_24886,N_24162,N_24107);
or U24887 (N_24887,N_24577,N_24368);
nor U24888 (N_24888,N_24011,N_24425);
or U24889 (N_24889,N_24032,N_24345);
nor U24890 (N_24890,N_24055,N_24102);
nand U24891 (N_24891,N_24274,N_24204);
nor U24892 (N_24892,N_24157,N_24396);
nand U24893 (N_24893,N_24542,N_24342);
xnor U24894 (N_24894,N_24495,N_24282);
or U24895 (N_24895,N_24170,N_24249);
or U24896 (N_24896,N_24462,N_24172);
nand U24897 (N_24897,N_24125,N_24181);
xor U24898 (N_24898,N_24265,N_24271);
or U24899 (N_24899,N_24203,N_24071);
nand U24900 (N_24900,N_24462,N_24594);
nor U24901 (N_24901,N_24487,N_24427);
nor U24902 (N_24902,N_24372,N_24106);
or U24903 (N_24903,N_24085,N_24198);
nand U24904 (N_24904,N_24165,N_24238);
nand U24905 (N_24905,N_24391,N_24045);
and U24906 (N_24906,N_24518,N_24388);
xnor U24907 (N_24907,N_24526,N_24510);
nor U24908 (N_24908,N_24040,N_24406);
nor U24909 (N_24909,N_24168,N_24027);
and U24910 (N_24910,N_24336,N_24526);
and U24911 (N_24911,N_24247,N_24503);
xnor U24912 (N_24912,N_24578,N_24076);
and U24913 (N_24913,N_24532,N_24225);
nand U24914 (N_24914,N_24173,N_24548);
xor U24915 (N_24915,N_24517,N_24191);
or U24916 (N_24916,N_24168,N_24325);
and U24917 (N_24917,N_24143,N_24317);
nand U24918 (N_24918,N_24357,N_24193);
nor U24919 (N_24919,N_24280,N_24353);
nor U24920 (N_24920,N_24559,N_24461);
or U24921 (N_24921,N_24049,N_24422);
or U24922 (N_24922,N_24458,N_24319);
nor U24923 (N_24923,N_24451,N_24146);
and U24924 (N_24924,N_24046,N_24458);
and U24925 (N_24925,N_24180,N_24008);
or U24926 (N_24926,N_24577,N_24228);
or U24927 (N_24927,N_24120,N_24181);
or U24928 (N_24928,N_24292,N_24380);
xor U24929 (N_24929,N_24285,N_24114);
nand U24930 (N_24930,N_24431,N_24320);
nor U24931 (N_24931,N_24306,N_24206);
nor U24932 (N_24932,N_24480,N_24542);
nor U24933 (N_24933,N_24263,N_24166);
xnor U24934 (N_24934,N_24434,N_24040);
nor U24935 (N_24935,N_24356,N_24208);
and U24936 (N_24936,N_24092,N_24060);
nand U24937 (N_24937,N_24182,N_24307);
nor U24938 (N_24938,N_24236,N_24304);
nand U24939 (N_24939,N_24464,N_24160);
and U24940 (N_24940,N_24495,N_24270);
or U24941 (N_24941,N_24562,N_24429);
xnor U24942 (N_24942,N_24031,N_24289);
or U24943 (N_24943,N_24440,N_24500);
nand U24944 (N_24944,N_24013,N_24414);
xor U24945 (N_24945,N_24563,N_24361);
xnor U24946 (N_24946,N_24518,N_24549);
nor U24947 (N_24947,N_24228,N_24536);
and U24948 (N_24948,N_24553,N_24550);
nand U24949 (N_24949,N_24520,N_24525);
or U24950 (N_24950,N_24303,N_24430);
xor U24951 (N_24951,N_24285,N_24198);
nor U24952 (N_24952,N_24132,N_24362);
nand U24953 (N_24953,N_24403,N_24532);
nand U24954 (N_24954,N_24192,N_24407);
nor U24955 (N_24955,N_24533,N_24121);
and U24956 (N_24956,N_24357,N_24531);
nor U24957 (N_24957,N_24326,N_24512);
and U24958 (N_24958,N_24468,N_24384);
or U24959 (N_24959,N_24140,N_24375);
and U24960 (N_24960,N_24530,N_24066);
and U24961 (N_24961,N_24145,N_24511);
nor U24962 (N_24962,N_24467,N_24049);
and U24963 (N_24963,N_24278,N_24289);
xor U24964 (N_24964,N_24527,N_24529);
or U24965 (N_24965,N_24188,N_24439);
and U24966 (N_24966,N_24505,N_24450);
nand U24967 (N_24967,N_24141,N_24575);
or U24968 (N_24968,N_24082,N_24216);
nor U24969 (N_24969,N_24153,N_24238);
xor U24970 (N_24970,N_24391,N_24281);
nand U24971 (N_24971,N_24141,N_24393);
and U24972 (N_24972,N_24414,N_24450);
nor U24973 (N_24973,N_24592,N_24090);
and U24974 (N_24974,N_24139,N_24571);
or U24975 (N_24975,N_24265,N_24202);
xor U24976 (N_24976,N_24453,N_24177);
nor U24977 (N_24977,N_24475,N_24110);
and U24978 (N_24978,N_24376,N_24126);
nand U24979 (N_24979,N_24252,N_24029);
or U24980 (N_24980,N_24282,N_24026);
nand U24981 (N_24981,N_24175,N_24575);
nand U24982 (N_24982,N_24474,N_24206);
xnor U24983 (N_24983,N_24261,N_24079);
nand U24984 (N_24984,N_24164,N_24208);
nand U24985 (N_24985,N_24255,N_24349);
and U24986 (N_24986,N_24369,N_24075);
nand U24987 (N_24987,N_24152,N_24050);
and U24988 (N_24988,N_24322,N_24142);
xnor U24989 (N_24989,N_24252,N_24523);
or U24990 (N_24990,N_24531,N_24274);
xnor U24991 (N_24991,N_24224,N_24471);
and U24992 (N_24992,N_24028,N_24316);
nor U24993 (N_24993,N_24492,N_24502);
xnor U24994 (N_24994,N_24383,N_24132);
nand U24995 (N_24995,N_24560,N_24504);
nor U24996 (N_24996,N_24004,N_24289);
nor U24997 (N_24997,N_24316,N_24396);
and U24998 (N_24998,N_24110,N_24451);
or U24999 (N_24999,N_24477,N_24219);
xor U25000 (N_25000,N_24331,N_24477);
and U25001 (N_25001,N_24232,N_24594);
and U25002 (N_25002,N_24524,N_24211);
nor U25003 (N_25003,N_24545,N_24084);
or U25004 (N_25004,N_24292,N_24152);
and U25005 (N_25005,N_24333,N_24489);
nand U25006 (N_25006,N_24124,N_24429);
xor U25007 (N_25007,N_24013,N_24273);
and U25008 (N_25008,N_24558,N_24242);
xor U25009 (N_25009,N_24042,N_24178);
nand U25010 (N_25010,N_24598,N_24353);
nor U25011 (N_25011,N_24073,N_24348);
nand U25012 (N_25012,N_24057,N_24425);
or U25013 (N_25013,N_24271,N_24238);
nor U25014 (N_25014,N_24544,N_24034);
or U25015 (N_25015,N_24495,N_24215);
and U25016 (N_25016,N_24552,N_24488);
and U25017 (N_25017,N_24338,N_24571);
nor U25018 (N_25018,N_24354,N_24254);
nand U25019 (N_25019,N_24503,N_24571);
nor U25020 (N_25020,N_24333,N_24563);
or U25021 (N_25021,N_24190,N_24392);
nor U25022 (N_25022,N_24431,N_24462);
nor U25023 (N_25023,N_24326,N_24218);
nand U25024 (N_25024,N_24287,N_24352);
or U25025 (N_25025,N_24301,N_24196);
or U25026 (N_25026,N_24107,N_24014);
xor U25027 (N_25027,N_24049,N_24316);
xnor U25028 (N_25028,N_24458,N_24339);
and U25029 (N_25029,N_24166,N_24394);
xnor U25030 (N_25030,N_24596,N_24284);
nand U25031 (N_25031,N_24062,N_24548);
or U25032 (N_25032,N_24311,N_24256);
nor U25033 (N_25033,N_24437,N_24350);
or U25034 (N_25034,N_24539,N_24286);
or U25035 (N_25035,N_24583,N_24555);
nor U25036 (N_25036,N_24238,N_24484);
xnor U25037 (N_25037,N_24052,N_24008);
nor U25038 (N_25038,N_24192,N_24282);
nand U25039 (N_25039,N_24336,N_24511);
nand U25040 (N_25040,N_24104,N_24447);
nand U25041 (N_25041,N_24186,N_24465);
or U25042 (N_25042,N_24162,N_24276);
nand U25043 (N_25043,N_24233,N_24546);
nand U25044 (N_25044,N_24540,N_24329);
and U25045 (N_25045,N_24290,N_24011);
and U25046 (N_25046,N_24277,N_24458);
and U25047 (N_25047,N_24156,N_24234);
xor U25048 (N_25048,N_24323,N_24270);
nor U25049 (N_25049,N_24429,N_24269);
or U25050 (N_25050,N_24006,N_24036);
xor U25051 (N_25051,N_24476,N_24306);
nand U25052 (N_25052,N_24540,N_24355);
or U25053 (N_25053,N_24304,N_24403);
or U25054 (N_25054,N_24010,N_24442);
nand U25055 (N_25055,N_24500,N_24314);
and U25056 (N_25056,N_24045,N_24309);
or U25057 (N_25057,N_24092,N_24172);
or U25058 (N_25058,N_24310,N_24280);
xor U25059 (N_25059,N_24338,N_24143);
nor U25060 (N_25060,N_24406,N_24529);
nand U25061 (N_25061,N_24504,N_24378);
and U25062 (N_25062,N_24093,N_24459);
xor U25063 (N_25063,N_24168,N_24346);
or U25064 (N_25064,N_24148,N_24582);
nor U25065 (N_25065,N_24510,N_24513);
or U25066 (N_25066,N_24483,N_24376);
xor U25067 (N_25067,N_24058,N_24469);
xor U25068 (N_25068,N_24502,N_24188);
nand U25069 (N_25069,N_24599,N_24218);
or U25070 (N_25070,N_24063,N_24387);
and U25071 (N_25071,N_24364,N_24159);
nor U25072 (N_25072,N_24464,N_24266);
xnor U25073 (N_25073,N_24565,N_24302);
and U25074 (N_25074,N_24040,N_24001);
and U25075 (N_25075,N_24071,N_24364);
or U25076 (N_25076,N_24250,N_24056);
nor U25077 (N_25077,N_24480,N_24113);
nand U25078 (N_25078,N_24460,N_24222);
and U25079 (N_25079,N_24386,N_24238);
nand U25080 (N_25080,N_24221,N_24544);
xor U25081 (N_25081,N_24092,N_24453);
or U25082 (N_25082,N_24364,N_24056);
and U25083 (N_25083,N_24272,N_24520);
and U25084 (N_25084,N_24283,N_24018);
nor U25085 (N_25085,N_24129,N_24590);
xnor U25086 (N_25086,N_24579,N_24158);
nand U25087 (N_25087,N_24254,N_24453);
and U25088 (N_25088,N_24088,N_24337);
nor U25089 (N_25089,N_24059,N_24407);
xnor U25090 (N_25090,N_24072,N_24176);
and U25091 (N_25091,N_24022,N_24588);
xnor U25092 (N_25092,N_24169,N_24311);
nor U25093 (N_25093,N_24314,N_24433);
or U25094 (N_25094,N_24091,N_24481);
nand U25095 (N_25095,N_24530,N_24177);
and U25096 (N_25096,N_24472,N_24162);
nor U25097 (N_25097,N_24259,N_24444);
or U25098 (N_25098,N_24493,N_24218);
nor U25099 (N_25099,N_24251,N_24508);
or U25100 (N_25100,N_24183,N_24037);
and U25101 (N_25101,N_24440,N_24576);
or U25102 (N_25102,N_24065,N_24320);
nand U25103 (N_25103,N_24180,N_24401);
nor U25104 (N_25104,N_24075,N_24316);
and U25105 (N_25105,N_24385,N_24152);
or U25106 (N_25106,N_24246,N_24461);
and U25107 (N_25107,N_24512,N_24393);
and U25108 (N_25108,N_24340,N_24332);
nand U25109 (N_25109,N_24491,N_24549);
nand U25110 (N_25110,N_24120,N_24030);
xnor U25111 (N_25111,N_24571,N_24465);
nand U25112 (N_25112,N_24236,N_24560);
nor U25113 (N_25113,N_24516,N_24353);
xor U25114 (N_25114,N_24081,N_24539);
xor U25115 (N_25115,N_24589,N_24535);
or U25116 (N_25116,N_24068,N_24295);
nand U25117 (N_25117,N_24450,N_24026);
xor U25118 (N_25118,N_24087,N_24451);
and U25119 (N_25119,N_24291,N_24008);
nand U25120 (N_25120,N_24030,N_24188);
or U25121 (N_25121,N_24392,N_24540);
xor U25122 (N_25122,N_24422,N_24168);
xor U25123 (N_25123,N_24584,N_24110);
and U25124 (N_25124,N_24109,N_24182);
and U25125 (N_25125,N_24207,N_24063);
xor U25126 (N_25126,N_24580,N_24076);
nor U25127 (N_25127,N_24581,N_24293);
nor U25128 (N_25128,N_24598,N_24092);
and U25129 (N_25129,N_24079,N_24438);
or U25130 (N_25130,N_24296,N_24078);
and U25131 (N_25131,N_24536,N_24263);
and U25132 (N_25132,N_24449,N_24187);
and U25133 (N_25133,N_24161,N_24422);
nand U25134 (N_25134,N_24234,N_24529);
xor U25135 (N_25135,N_24021,N_24361);
or U25136 (N_25136,N_24104,N_24041);
nand U25137 (N_25137,N_24006,N_24534);
nor U25138 (N_25138,N_24200,N_24374);
nand U25139 (N_25139,N_24151,N_24217);
xor U25140 (N_25140,N_24239,N_24162);
or U25141 (N_25141,N_24329,N_24364);
nand U25142 (N_25142,N_24282,N_24577);
nand U25143 (N_25143,N_24564,N_24502);
or U25144 (N_25144,N_24281,N_24304);
or U25145 (N_25145,N_24474,N_24335);
xnor U25146 (N_25146,N_24374,N_24248);
and U25147 (N_25147,N_24172,N_24082);
or U25148 (N_25148,N_24048,N_24165);
and U25149 (N_25149,N_24001,N_24141);
and U25150 (N_25150,N_24410,N_24454);
xnor U25151 (N_25151,N_24017,N_24453);
xor U25152 (N_25152,N_24226,N_24429);
or U25153 (N_25153,N_24245,N_24258);
and U25154 (N_25154,N_24299,N_24078);
and U25155 (N_25155,N_24332,N_24024);
xor U25156 (N_25156,N_24134,N_24133);
xnor U25157 (N_25157,N_24588,N_24514);
or U25158 (N_25158,N_24457,N_24181);
nand U25159 (N_25159,N_24220,N_24150);
nor U25160 (N_25160,N_24350,N_24439);
nor U25161 (N_25161,N_24555,N_24356);
nand U25162 (N_25162,N_24223,N_24312);
nor U25163 (N_25163,N_24421,N_24385);
xnor U25164 (N_25164,N_24090,N_24263);
and U25165 (N_25165,N_24303,N_24057);
xnor U25166 (N_25166,N_24205,N_24325);
nand U25167 (N_25167,N_24461,N_24515);
nand U25168 (N_25168,N_24317,N_24241);
xor U25169 (N_25169,N_24390,N_24087);
nand U25170 (N_25170,N_24317,N_24322);
xor U25171 (N_25171,N_24241,N_24021);
and U25172 (N_25172,N_24316,N_24549);
nand U25173 (N_25173,N_24289,N_24267);
xor U25174 (N_25174,N_24463,N_24375);
or U25175 (N_25175,N_24394,N_24554);
or U25176 (N_25176,N_24268,N_24428);
or U25177 (N_25177,N_24075,N_24241);
or U25178 (N_25178,N_24067,N_24048);
nand U25179 (N_25179,N_24141,N_24036);
and U25180 (N_25180,N_24477,N_24108);
xnor U25181 (N_25181,N_24088,N_24210);
and U25182 (N_25182,N_24303,N_24018);
or U25183 (N_25183,N_24232,N_24512);
nor U25184 (N_25184,N_24274,N_24483);
or U25185 (N_25185,N_24379,N_24076);
and U25186 (N_25186,N_24027,N_24544);
nand U25187 (N_25187,N_24157,N_24292);
xnor U25188 (N_25188,N_24465,N_24240);
or U25189 (N_25189,N_24103,N_24298);
nor U25190 (N_25190,N_24285,N_24438);
nand U25191 (N_25191,N_24195,N_24138);
xor U25192 (N_25192,N_24588,N_24161);
or U25193 (N_25193,N_24045,N_24171);
nor U25194 (N_25194,N_24517,N_24327);
xor U25195 (N_25195,N_24258,N_24595);
and U25196 (N_25196,N_24501,N_24071);
or U25197 (N_25197,N_24164,N_24111);
nand U25198 (N_25198,N_24224,N_24155);
or U25199 (N_25199,N_24415,N_24406);
nor U25200 (N_25200,N_24727,N_25108);
xnor U25201 (N_25201,N_24816,N_25128);
nand U25202 (N_25202,N_25176,N_24675);
nand U25203 (N_25203,N_25045,N_24858);
nor U25204 (N_25204,N_24879,N_24868);
xnor U25205 (N_25205,N_24708,N_24739);
or U25206 (N_25206,N_24789,N_24856);
and U25207 (N_25207,N_24688,N_25072);
nand U25208 (N_25208,N_25051,N_24793);
xor U25209 (N_25209,N_24875,N_24953);
and U25210 (N_25210,N_25162,N_24670);
and U25211 (N_25211,N_25174,N_24844);
xnor U25212 (N_25212,N_24831,N_24887);
or U25213 (N_25213,N_25075,N_24909);
xnor U25214 (N_25214,N_25151,N_24780);
nor U25215 (N_25215,N_24933,N_24796);
nand U25216 (N_25216,N_24797,N_24735);
and U25217 (N_25217,N_25018,N_24666);
or U25218 (N_25218,N_25147,N_25104);
xnor U25219 (N_25219,N_25066,N_25123);
xor U25220 (N_25220,N_24872,N_24608);
xor U25221 (N_25221,N_25120,N_24745);
and U25222 (N_25222,N_24792,N_24896);
xnor U25223 (N_25223,N_24852,N_25154);
nand U25224 (N_25224,N_24993,N_24799);
or U25225 (N_25225,N_24604,N_25191);
nand U25226 (N_25226,N_24818,N_24956);
xnor U25227 (N_25227,N_25171,N_24821);
nor U25228 (N_25228,N_25060,N_25166);
or U25229 (N_25229,N_24746,N_24683);
nand U25230 (N_25230,N_24696,N_25110);
nor U25231 (N_25231,N_24772,N_24864);
xor U25232 (N_25232,N_24658,N_25119);
nor U25233 (N_25233,N_25199,N_25161);
xnor U25234 (N_25234,N_24878,N_24988);
nor U25235 (N_25235,N_24918,N_25153);
and U25236 (N_25236,N_25041,N_25084);
nor U25237 (N_25237,N_24775,N_24890);
nor U25238 (N_25238,N_24718,N_25182);
nor U25239 (N_25239,N_25013,N_25136);
xnor U25240 (N_25240,N_24862,N_25054);
or U25241 (N_25241,N_24992,N_24968);
nor U25242 (N_25242,N_24954,N_24960);
or U25243 (N_25243,N_24689,N_24921);
nand U25244 (N_25244,N_24750,N_24805);
and U25245 (N_25245,N_24606,N_24810);
nor U25246 (N_25246,N_24659,N_24947);
or U25247 (N_25247,N_24945,N_24731);
and U25248 (N_25248,N_24903,N_24698);
nor U25249 (N_25249,N_24867,N_25003);
and U25250 (N_25250,N_24777,N_24702);
or U25251 (N_25251,N_25085,N_24725);
xnor U25252 (N_25252,N_24785,N_25062);
nand U25253 (N_25253,N_25142,N_24733);
xnor U25254 (N_25254,N_24663,N_25083);
nand U25255 (N_25255,N_24760,N_25036);
xor U25256 (N_25256,N_24850,N_25094);
and U25257 (N_25257,N_25179,N_24685);
nor U25258 (N_25258,N_24961,N_25076);
nand U25259 (N_25259,N_24815,N_24943);
and U25260 (N_25260,N_24619,N_25080);
nor U25261 (N_25261,N_25074,N_24631);
xor U25262 (N_25262,N_24749,N_24782);
nor U25263 (N_25263,N_25004,N_24932);
xnor U25264 (N_25264,N_24808,N_25052);
and U25265 (N_25265,N_24969,N_25073);
and U25266 (N_25266,N_24617,N_24964);
and U25267 (N_25267,N_24712,N_25088);
nor U25268 (N_25268,N_25126,N_25117);
nand U25269 (N_25269,N_25095,N_24625);
nand U25270 (N_25270,N_25158,N_24840);
and U25271 (N_25271,N_24835,N_25091);
xor U25272 (N_25272,N_25043,N_24916);
nand U25273 (N_25273,N_24755,N_25030);
nand U25274 (N_25274,N_25145,N_24700);
or U25275 (N_25275,N_25037,N_24703);
nand U25276 (N_25276,N_24829,N_24667);
nor U25277 (N_25277,N_24824,N_24940);
or U25278 (N_25278,N_25113,N_24929);
or U25279 (N_25279,N_24905,N_24788);
or U25280 (N_25280,N_24740,N_24966);
or U25281 (N_25281,N_24819,N_24915);
xnor U25282 (N_25282,N_24711,N_24763);
or U25283 (N_25283,N_24946,N_24889);
nand U25284 (N_25284,N_24853,N_24798);
xor U25285 (N_25285,N_25040,N_24978);
and U25286 (N_25286,N_25038,N_25170);
xor U25287 (N_25287,N_24690,N_24999);
nor U25288 (N_25288,N_24774,N_24776);
xnor U25289 (N_25289,N_24838,N_25102);
nor U25290 (N_25290,N_24734,N_24975);
nor U25291 (N_25291,N_24942,N_25061);
and U25292 (N_25292,N_24614,N_24633);
xnor U25293 (N_25293,N_24884,N_24672);
xnor U25294 (N_25294,N_24678,N_24795);
and U25295 (N_25295,N_24653,N_24847);
xor U25296 (N_25296,N_24985,N_24743);
nor U25297 (N_25297,N_24938,N_24710);
nand U25298 (N_25298,N_24822,N_24849);
and U25299 (N_25299,N_24923,N_24638);
or U25300 (N_25300,N_25134,N_24748);
nor U25301 (N_25301,N_25164,N_24935);
nor U25302 (N_25302,N_25109,N_24680);
or U25303 (N_25303,N_24976,N_25016);
and U25304 (N_25304,N_24699,N_24624);
nand U25305 (N_25305,N_24963,N_24610);
xnor U25306 (N_25306,N_24924,N_25141);
or U25307 (N_25307,N_24726,N_24769);
or U25308 (N_25308,N_24605,N_24626);
and U25309 (N_25309,N_25024,N_24973);
or U25310 (N_25310,N_25089,N_25168);
nor U25311 (N_25311,N_25068,N_24939);
and U25312 (N_25312,N_25114,N_24640);
nand U25313 (N_25313,N_24997,N_24691);
or U25314 (N_25314,N_25053,N_24803);
and U25315 (N_25315,N_25186,N_24627);
or U25316 (N_25316,N_25020,N_25106);
xnor U25317 (N_25317,N_24669,N_24836);
nand U25318 (N_25318,N_24860,N_24714);
and U25319 (N_25319,N_24671,N_25070);
xnor U25320 (N_25320,N_25196,N_25121);
xnor U25321 (N_25321,N_24650,N_24995);
nor U25322 (N_25322,N_25178,N_24637);
xor U25323 (N_25323,N_24888,N_24880);
or U25324 (N_25324,N_25099,N_24778);
xor U25325 (N_25325,N_24870,N_24828);
or U25326 (N_25326,N_25001,N_24830);
nor U25327 (N_25327,N_25077,N_24902);
nor U25328 (N_25328,N_24987,N_25194);
and U25329 (N_25329,N_25048,N_25044);
and U25330 (N_25330,N_24766,N_25148);
nor U25331 (N_25331,N_24720,N_25130);
nor U25332 (N_25332,N_24705,N_24756);
and U25333 (N_25333,N_25069,N_24704);
and U25334 (N_25334,N_25090,N_24645);
xnor U25335 (N_25335,N_24790,N_24959);
or U25336 (N_25336,N_24832,N_25014);
nor U25337 (N_25337,N_24899,N_24621);
or U25338 (N_25338,N_25193,N_24982);
and U25339 (N_25339,N_24842,N_24834);
and U25340 (N_25340,N_24767,N_25049);
nand U25341 (N_25341,N_24996,N_25175);
and U25342 (N_25342,N_24761,N_24732);
or U25343 (N_25343,N_24931,N_25096);
xor U25344 (N_25344,N_24794,N_24812);
nand U25345 (N_25345,N_24676,N_24859);
nand U25346 (N_25346,N_25185,N_25116);
or U25347 (N_25347,N_24764,N_24674);
nor U25348 (N_25348,N_24677,N_25046);
xnor U25349 (N_25349,N_24693,N_24679);
and U25350 (N_25350,N_24657,N_25167);
or U25351 (N_25351,N_24636,N_24930);
nor U25352 (N_25352,N_24607,N_24948);
xnor U25353 (N_25353,N_24613,N_24656);
nor U25354 (N_25354,N_24660,N_24773);
nand U25355 (N_25355,N_24919,N_25056);
nand U25356 (N_25356,N_24787,N_24781);
xor U25357 (N_25357,N_25086,N_24706);
or U25358 (N_25358,N_25042,N_25055);
nor U25359 (N_25359,N_24861,N_25137);
or U25360 (N_25360,N_24846,N_24717);
and U25361 (N_25361,N_25008,N_25047);
xnor U25362 (N_25362,N_24928,N_24723);
xnor U25363 (N_25363,N_24837,N_24759);
xnor U25364 (N_25364,N_24747,N_24786);
or U25365 (N_25365,N_25188,N_25146);
nor U25366 (N_25366,N_24986,N_24843);
or U25367 (N_25367,N_24715,N_25079);
nand U25368 (N_25368,N_25152,N_24673);
xnor U25369 (N_25369,N_25063,N_25101);
nand U25370 (N_25370,N_25189,N_25122);
nand U25371 (N_25371,N_25165,N_24904);
and U25372 (N_25372,N_24779,N_24970);
or U25373 (N_25373,N_24643,N_24998);
nand U25374 (N_25374,N_24967,N_24694);
nor U25375 (N_25375,N_24925,N_24983);
or U25376 (N_25376,N_24937,N_24791);
and U25377 (N_25377,N_24753,N_24883);
and U25378 (N_25378,N_24618,N_24817);
and U25379 (N_25379,N_25034,N_24994);
nand U25380 (N_25380,N_24655,N_25160);
nand U25381 (N_25381,N_24632,N_24800);
nand U25382 (N_25382,N_24603,N_24724);
nand U25383 (N_25383,N_25092,N_24941);
or U25384 (N_25384,N_24936,N_25125);
nor U25385 (N_25385,N_25118,N_25082);
xnor U25386 (N_25386,N_24742,N_24802);
and U25387 (N_25387,N_25180,N_24770);
nand U25388 (N_25388,N_24971,N_24885);
nand U25389 (N_25389,N_24713,N_24965);
nand U25390 (N_25390,N_25023,N_24913);
nand U25391 (N_25391,N_25028,N_25197);
and U25392 (N_25392,N_25112,N_24681);
nor U25393 (N_25393,N_24744,N_24820);
or U25394 (N_25394,N_24736,N_24922);
nand U25395 (N_25395,N_24665,N_25031);
xor U25396 (N_25396,N_24926,N_24651);
xor U25397 (N_25397,N_24991,N_25050);
or U25398 (N_25398,N_24845,N_24668);
or U25399 (N_25399,N_25124,N_24851);
or U25400 (N_25400,N_24962,N_25071);
or U25401 (N_25401,N_25032,N_24980);
or U25402 (N_25402,N_24757,N_24891);
or U25403 (N_25403,N_25025,N_24639);
nand U25404 (N_25404,N_24701,N_25057);
xor U25405 (N_25405,N_24754,N_25131);
nand U25406 (N_25406,N_25150,N_25012);
nand U25407 (N_25407,N_25035,N_25177);
or U25408 (N_25408,N_24752,N_25005);
xnor U25409 (N_25409,N_24839,N_24662);
nand U25410 (N_25410,N_25111,N_24762);
xnor U25411 (N_25411,N_24895,N_25100);
nand U25412 (N_25412,N_25187,N_24893);
or U25413 (N_25413,N_24897,N_25172);
or U25414 (N_25414,N_24981,N_25143);
xnor U25415 (N_25415,N_24811,N_24623);
xnor U25416 (N_25416,N_24881,N_24984);
and U25417 (N_25417,N_24951,N_24709);
xor U25418 (N_25418,N_24876,N_25163);
and U25419 (N_25419,N_24609,N_25002);
nor U25420 (N_25420,N_24801,N_25156);
and U25421 (N_25421,N_24911,N_24611);
and U25422 (N_25422,N_24661,N_24654);
and U25423 (N_25423,N_24866,N_24616);
nand U25424 (N_25424,N_24707,N_25144);
nand U25425 (N_25425,N_24634,N_25138);
nor U25426 (N_25426,N_24692,N_24871);
nand U25427 (N_25427,N_25169,N_25135);
nand U25428 (N_25428,N_24644,N_25019);
nand U25429 (N_25429,N_24944,N_24894);
xnor U25430 (N_25430,N_25097,N_24768);
nor U25431 (N_25431,N_24825,N_25006);
or U25432 (N_25432,N_24728,N_24814);
nor U25433 (N_25433,N_25132,N_24841);
xnor U25434 (N_25434,N_25159,N_24730);
or U25435 (N_25435,N_25022,N_25039);
and U25436 (N_25436,N_24920,N_24684);
or U25437 (N_25437,N_24642,N_24869);
and U25438 (N_25438,N_25067,N_24863);
nand U25439 (N_25439,N_24813,N_25017);
nor U25440 (N_25440,N_25181,N_25155);
nand U25441 (N_25441,N_25010,N_24927);
or U25442 (N_25442,N_24857,N_25064);
and U25443 (N_25443,N_25103,N_24729);
or U25444 (N_25444,N_25026,N_24807);
and U25445 (N_25445,N_25192,N_24912);
nand U25446 (N_25446,N_24664,N_25087);
nor U25447 (N_25447,N_24771,N_24827);
nand U25448 (N_25448,N_25000,N_24620);
xnor U25449 (N_25449,N_24641,N_24622);
and U25450 (N_25450,N_24635,N_24647);
or U25451 (N_25451,N_24865,N_25105);
nor U25452 (N_25452,N_24854,N_25198);
or U25453 (N_25453,N_24958,N_24615);
nand U25454 (N_25454,N_24906,N_25081);
nor U25455 (N_25455,N_25173,N_24758);
or U25456 (N_25456,N_25183,N_24914);
xnor U25457 (N_25457,N_24901,N_25009);
or U25458 (N_25458,N_24695,N_24601);
and U25459 (N_25459,N_25093,N_25139);
xnor U25460 (N_25460,N_24877,N_24649);
xnor U25461 (N_25461,N_24687,N_24977);
nor U25462 (N_25462,N_24721,N_24600);
nand U25463 (N_25463,N_25065,N_24949);
and U25464 (N_25464,N_24873,N_24629);
or U25465 (N_25465,N_24646,N_24612);
nor U25466 (N_25466,N_25190,N_24974);
nand U25467 (N_25467,N_25184,N_25027);
nand U25468 (N_25468,N_25115,N_25127);
nand U25469 (N_25469,N_24907,N_25129);
or U25470 (N_25470,N_25133,N_25021);
or U25471 (N_25471,N_24806,N_24874);
or U25472 (N_25472,N_24898,N_24784);
nor U25473 (N_25473,N_24722,N_24833);
and U25474 (N_25474,N_24751,N_24765);
nor U25475 (N_25475,N_24957,N_24716);
xor U25476 (N_25476,N_24823,N_25098);
or U25477 (N_25477,N_24910,N_24686);
xnor U25478 (N_25478,N_24682,N_25149);
nor U25479 (N_25479,N_24989,N_25033);
xor U25480 (N_25480,N_24648,N_25107);
nand U25481 (N_25481,N_24917,N_25011);
and U25482 (N_25482,N_25078,N_24934);
nor U25483 (N_25483,N_25195,N_24979);
or U25484 (N_25484,N_24848,N_24783);
xor U25485 (N_25485,N_24882,N_25007);
xnor U25486 (N_25486,N_24950,N_24652);
xnor U25487 (N_25487,N_24737,N_24892);
nand U25488 (N_25488,N_24955,N_24855);
nand U25489 (N_25489,N_25059,N_24900);
or U25490 (N_25490,N_25140,N_24741);
nand U25491 (N_25491,N_24697,N_24952);
nor U25492 (N_25492,N_24990,N_24630);
and U25493 (N_25493,N_24809,N_24908);
nor U25494 (N_25494,N_25029,N_24719);
or U25495 (N_25495,N_24602,N_24738);
and U25496 (N_25496,N_25058,N_25157);
and U25497 (N_25497,N_24972,N_24886);
xor U25498 (N_25498,N_25015,N_24628);
and U25499 (N_25499,N_24826,N_24804);
nor U25500 (N_25500,N_24868,N_24663);
xor U25501 (N_25501,N_24730,N_24998);
nand U25502 (N_25502,N_25163,N_25058);
or U25503 (N_25503,N_25025,N_24916);
and U25504 (N_25504,N_25070,N_24764);
nand U25505 (N_25505,N_25167,N_25098);
or U25506 (N_25506,N_25082,N_24816);
or U25507 (N_25507,N_24746,N_25145);
and U25508 (N_25508,N_25100,N_24627);
nand U25509 (N_25509,N_24952,N_24844);
xor U25510 (N_25510,N_24719,N_24712);
nand U25511 (N_25511,N_24668,N_25126);
or U25512 (N_25512,N_24850,N_25027);
nor U25513 (N_25513,N_24764,N_24680);
nand U25514 (N_25514,N_24745,N_24817);
or U25515 (N_25515,N_25159,N_24941);
nor U25516 (N_25516,N_25114,N_25158);
and U25517 (N_25517,N_24748,N_24786);
nand U25518 (N_25518,N_24606,N_24671);
nand U25519 (N_25519,N_24874,N_25037);
or U25520 (N_25520,N_25065,N_25090);
xnor U25521 (N_25521,N_24693,N_24787);
nand U25522 (N_25522,N_24689,N_24790);
nand U25523 (N_25523,N_25128,N_24731);
or U25524 (N_25524,N_25059,N_24615);
nor U25525 (N_25525,N_25190,N_25054);
xor U25526 (N_25526,N_24621,N_24893);
and U25527 (N_25527,N_24915,N_24817);
or U25528 (N_25528,N_24633,N_24982);
nand U25529 (N_25529,N_24698,N_25198);
or U25530 (N_25530,N_24989,N_24829);
or U25531 (N_25531,N_24634,N_25153);
xnor U25532 (N_25532,N_24664,N_25172);
nand U25533 (N_25533,N_25159,N_25121);
or U25534 (N_25534,N_24910,N_24845);
nand U25535 (N_25535,N_24847,N_25194);
nand U25536 (N_25536,N_25126,N_24684);
xnor U25537 (N_25537,N_24852,N_24652);
xnor U25538 (N_25538,N_25055,N_24950);
xor U25539 (N_25539,N_24697,N_24878);
and U25540 (N_25540,N_24976,N_24941);
or U25541 (N_25541,N_24935,N_24920);
and U25542 (N_25542,N_24950,N_25131);
xor U25543 (N_25543,N_25111,N_24667);
nor U25544 (N_25544,N_24751,N_24752);
and U25545 (N_25545,N_24790,N_25118);
xor U25546 (N_25546,N_25022,N_24909);
nand U25547 (N_25547,N_25016,N_25026);
nand U25548 (N_25548,N_24991,N_24803);
nand U25549 (N_25549,N_24909,N_25177);
nor U25550 (N_25550,N_24971,N_24757);
nor U25551 (N_25551,N_25139,N_25133);
and U25552 (N_25552,N_24628,N_24908);
and U25553 (N_25553,N_24722,N_24813);
nor U25554 (N_25554,N_25136,N_24810);
and U25555 (N_25555,N_25165,N_24716);
xor U25556 (N_25556,N_24732,N_24728);
xnor U25557 (N_25557,N_24920,N_24863);
nand U25558 (N_25558,N_24757,N_24818);
or U25559 (N_25559,N_24806,N_24876);
or U25560 (N_25560,N_24801,N_24666);
nand U25561 (N_25561,N_25087,N_24974);
nor U25562 (N_25562,N_24818,N_24800);
xor U25563 (N_25563,N_24962,N_24715);
nand U25564 (N_25564,N_25198,N_24940);
nor U25565 (N_25565,N_24616,N_24951);
and U25566 (N_25566,N_24698,N_24722);
nand U25567 (N_25567,N_25124,N_24655);
nand U25568 (N_25568,N_25161,N_25060);
nand U25569 (N_25569,N_24768,N_25079);
xor U25570 (N_25570,N_24962,N_24833);
or U25571 (N_25571,N_25004,N_24812);
xor U25572 (N_25572,N_25103,N_24800);
or U25573 (N_25573,N_24845,N_24858);
or U25574 (N_25574,N_24836,N_24638);
nand U25575 (N_25575,N_25192,N_25004);
xnor U25576 (N_25576,N_24909,N_25132);
xor U25577 (N_25577,N_25152,N_24951);
xor U25578 (N_25578,N_24865,N_24668);
and U25579 (N_25579,N_25196,N_24622);
nand U25580 (N_25580,N_25010,N_24865);
nor U25581 (N_25581,N_25065,N_24955);
and U25582 (N_25582,N_25078,N_24752);
nand U25583 (N_25583,N_25173,N_24830);
nor U25584 (N_25584,N_24825,N_24989);
xor U25585 (N_25585,N_24637,N_25060);
and U25586 (N_25586,N_24779,N_24620);
nor U25587 (N_25587,N_24749,N_25106);
or U25588 (N_25588,N_24752,N_24708);
nor U25589 (N_25589,N_24783,N_25155);
or U25590 (N_25590,N_24633,N_24872);
xnor U25591 (N_25591,N_24928,N_24719);
xnor U25592 (N_25592,N_24640,N_25002);
or U25593 (N_25593,N_25156,N_24845);
or U25594 (N_25594,N_25108,N_24624);
nand U25595 (N_25595,N_25068,N_25165);
and U25596 (N_25596,N_25195,N_24642);
and U25597 (N_25597,N_25059,N_24707);
or U25598 (N_25598,N_24688,N_25197);
xor U25599 (N_25599,N_24700,N_24857);
or U25600 (N_25600,N_24942,N_24644);
nor U25601 (N_25601,N_24982,N_25184);
or U25602 (N_25602,N_25179,N_24785);
or U25603 (N_25603,N_24991,N_25065);
and U25604 (N_25604,N_25107,N_24717);
or U25605 (N_25605,N_24662,N_24919);
and U25606 (N_25606,N_24762,N_24612);
and U25607 (N_25607,N_24987,N_25054);
xnor U25608 (N_25608,N_25075,N_24842);
nand U25609 (N_25609,N_24796,N_25159);
xor U25610 (N_25610,N_24826,N_25191);
nand U25611 (N_25611,N_24647,N_25187);
or U25612 (N_25612,N_24928,N_24732);
or U25613 (N_25613,N_25095,N_24885);
and U25614 (N_25614,N_25011,N_24740);
or U25615 (N_25615,N_24615,N_24915);
nand U25616 (N_25616,N_25013,N_25155);
or U25617 (N_25617,N_25042,N_25167);
xor U25618 (N_25618,N_24917,N_25147);
xnor U25619 (N_25619,N_24825,N_24714);
and U25620 (N_25620,N_24665,N_25033);
and U25621 (N_25621,N_24976,N_24958);
and U25622 (N_25622,N_24623,N_25008);
nand U25623 (N_25623,N_25048,N_25030);
xor U25624 (N_25624,N_25058,N_25160);
or U25625 (N_25625,N_24726,N_24956);
nand U25626 (N_25626,N_25177,N_25130);
xnor U25627 (N_25627,N_24857,N_25186);
or U25628 (N_25628,N_25010,N_25190);
or U25629 (N_25629,N_24782,N_24745);
and U25630 (N_25630,N_24779,N_24682);
nor U25631 (N_25631,N_24719,N_24618);
xnor U25632 (N_25632,N_24814,N_24669);
nand U25633 (N_25633,N_24705,N_24959);
xnor U25634 (N_25634,N_24662,N_24991);
nor U25635 (N_25635,N_25077,N_25024);
xnor U25636 (N_25636,N_25015,N_24716);
nor U25637 (N_25637,N_25064,N_24759);
xnor U25638 (N_25638,N_25191,N_24957);
and U25639 (N_25639,N_24821,N_25032);
nand U25640 (N_25640,N_24921,N_25023);
nor U25641 (N_25641,N_24636,N_25088);
nor U25642 (N_25642,N_25061,N_24867);
nand U25643 (N_25643,N_24731,N_24679);
nor U25644 (N_25644,N_24761,N_25014);
nor U25645 (N_25645,N_25168,N_25129);
and U25646 (N_25646,N_24722,N_24749);
and U25647 (N_25647,N_24815,N_24776);
xnor U25648 (N_25648,N_25007,N_25116);
nand U25649 (N_25649,N_25054,N_24842);
nand U25650 (N_25650,N_24954,N_24672);
xor U25651 (N_25651,N_25057,N_24990);
nor U25652 (N_25652,N_25108,N_24922);
and U25653 (N_25653,N_24692,N_24783);
xnor U25654 (N_25654,N_24753,N_24950);
xnor U25655 (N_25655,N_24675,N_24601);
xor U25656 (N_25656,N_24658,N_25071);
nand U25657 (N_25657,N_24713,N_25019);
nand U25658 (N_25658,N_24763,N_24869);
xor U25659 (N_25659,N_24702,N_25135);
and U25660 (N_25660,N_24958,N_24923);
xnor U25661 (N_25661,N_25197,N_25038);
and U25662 (N_25662,N_24975,N_24792);
and U25663 (N_25663,N_25146,N_24977);
xor U25664 (N_25664,N_24601,N_25198);
xnor U25665 (N_25665,N_25103,N_24970);
xor U25666 (N_25666,N_24671,N_25108);
or U25667 (N_25667,N_24844,N_24653);
and U25668 (N_25668,N_24808,N_24784);
xor U25669 (N_25669,N_25036,N_24826);
xor U25670 (N_25670,N_24853,N_25102);
nand U25671 (N_25671,N_24631,N_25125);
or U25672 (N_25672,N_24688,N_24967);
xor U25673 (N_25673,N_25027,N_24856);
nand U25674 (N_25674,N_24727,N_24881);
nor U25675 (N_25675,N_24779,N_24939);
xnor U25676 (N_25676,N_24908,N_24709);
nor U25677 (N_25677,N_25004,N_24616);
and U25678 (N_25678,N_25005,N_25054);
or U25679 (N_25679,N_24700,N_24996);
or U25680 (N_25680,N_24775,N_25030);
nand U25681 (N_25681,N_24630,N_24617);
nand U25682 (N_25682,N_25083,N_25181);
xor U25683 (N_25683,N_24732,N_25178);
nand U25684 (N_25684,N_24845,N_25170);
xor U25685 (N_25685,N_24946,N_25152);
and U25686 (N_25686,N_24688,N_25176);
nor U25687 (N_25687,N_25141,N_24721);
xnor U25688 (N_25688,N_25006,N_24779);
and U25689 (N_25689,N_24631,N_24655);
xor U25690 (N_25690,N_24760,N_24622);
or U25691 (N_25691,N_24768,N_25004);
nand U25692 (N_25692,N_25167,N_25129);
and U25693 (N_25693,N_24806,N_25159);
nand U25694 (N_25694,N_24604,N_24610);
or U25695 (N_25695,N_24854,N_24932);
xor U25696 (N_25696,N_25121,N_25082);
nor U25697 (N_25697,N_24741,N_25175);
xnor U25698 (N_25698,N_24679,N_25159);
xor U25699 (N_25699,N_24953,N_25009);
or U25700 (N_25700,N_24769,N_24992);
xnor U25701 (N_25701,N_24891,N_24924);
xnor U25702 (N_25702,N_24804,N_24907);
nand U25703 (N_25703,N_24912,N_25179);
or U25704 (N_25704,N_25012,N_25043);
or U25705 (N_25705,N_25051,N_24714);
and U25706 (N_25706,N_24922,N_24828);
nand U25707 (N_25707,N_25060,N_24958);
or U25708 (N_25708,N_25062,N_24610);
nand U25709 (N_25709,N_24811,N_24953);
nand U25710 (N_25710,N_24829,N_25057);
or U25711 (N_25711,N_24867,N_24641);
xnor U25712 (N_25712,N_24926,N_24908);
and U25713 (N_25713,N_24782,N_24951);
nor U25714 (N_25714,N_24700,N_25179);
nor U25715 (N_25715,N_24846,N_24690);
nor U25716 (N_25716,N_24774,N_24724);
xor U25717 (N_25717,N_24747,N_24714);
or U25718 (N_25718,N_24695,N_25136);
xnor U25719 (N_25719,N_25031,N_24795);
and U25720 (N_25720,N_24966,N_24967);
or U25721 (N_25721,N_25146,N_24756);
nor U25722 (N_25722,N_24871,N_25062);
and U25723 (N_25723,N_24699,N_24965);
xor U25724 (N_25724,N_24623,N_24630);
nand U25725 (N_25725,N_25189,N_25077);
nor U25726 (N_25726,N_24614,N_25159);
or U25727 (N_25727,N_25081,N_24731);
xnor U25728 (N_25728,N_25180,N_25064);
nor U25729 (N_25729,N_24714,N_25197);
and U25730 (N_25730,N_24631,N_24698);
nand U25731 (N_25731,N_24930,N_24668);
and U25732 (N_25732,N_25163,N_25112);
nand U25733 (N_25733,N_25068,N_24699);
or U25734 (N_25734,N_24600,N_24843);
or U25735 (N_25735,N_24806,N_24836);
nand U25736 (N_25736,N_25115,N_24676);
xor U25737 (N_25737,N_25140,N_24783);
nand U25738 (N_25738,N_24759,N_24854);
nor U25739 (N_25739,N_25189,N_25147);
and U25740 (N_25740,N_25006,N_24697);
nand U25741 (N_25741,N_24836,N_24779);
and U25742 (N_25742,N_25035,N_24792);
xor U25743 (N_25743,N_24627,N_24667);
xor U25744 (N_25744,N_24917,N_25010);
or U25745 (N_25745,N_24719,N_24840);
xor U25746 (N_25746,N_24865,N_24922);
xnor U25747 (N_25747,N_25083,N_24630);
and U25748 (N_25748,N_25157,N_25035);
and U25749 (N_25749,N_24885,N_25135);
xor U25750 (N_25750,N_25010,N_24899);
and U25751 (N_25751,N_24710,N_25080);
nand U25752 (N_25752,N_24631,N_24995);
nand U25753 (N_25753,N_25068,N_24701);
xnor U25754 (N_25754,N_25099,N_24998);
and U25755 (N_25755,N_25185,N_25022);
and U25756 (N_25756,N_25084,N_24950);
xor U25757 (N_25757,N_25171,N_24969);
xor U25758 (N_25758,N_24831,N_25182);
xor U25759 (N_25759,N_24670,N_25158);
or U25760 (N_25760,N_25128,N_25018);
and U25761 (N_25761,N_24682,N_24972);
nor U25762 (N_25762,N_24910,N_25060);
or U25763 (N_25763,N_24912,N_25122);
or U25764 (N_25764,N_24984,N_25160);
xnor U25765 (N_25765,N_24654,N_24645);
and U25766 (N_25766,N_24728,N_24727);
xor U25767 (N_25767,N_25120,N_25029);
and U25768 (N_25768,N_25027,N_25002);
nor U25769 (N_25769,N_24951,N_24913);
xnor U25770 (N_25770,N_24699,N_25059);
xnor U25771 (N_25771,N_24638,N_24741);
nor U25772 (N_25772,N_24913,N_25198);
or U25773 (N_25773,N_24673,N_24970);
nand U25774 (N_25774,N_25161,N_24725);
xor U25775 (N_25775,N_25048,N_24944);
nand U25776 (N_25776,N_25191,N_25004);
nand U25777 (N_25777,N_25013,N_24915);
xor U25778 (N_25778,N_24765,N_24683);
nor U25779 (N_25779,N_24603,N_24999);
nor U25780 (N_25780,N_25184,N_25196);
and U25781 (N_25781,N_25141,N_24870);
xnor U25782 (N_25782,N_25164,N_25194);
or U25783 (N_25783,N_24671,N_24662);
and U25784 (N_25784,N_25060,N_24697);
nand U25785 (N_25785,N_25076,N_25165);
xnor U25786 (N_25786,N_24896,N_25090);
and U25787 (N_25787,N_24622,N_24953);
xor U25788 (N_25788,N_25136,N_25077);
xor U25789 (N_25789,N_24630,N_24882);
nor U25790 (N_25790,N_25072,N_24908);
nor U25791 (N_25791,N_24628,N_25009);
nor U25792 (N_25792,N_24854,N_24818);
and U25793 (N_25793,N_24874,N_24939);
xnor U25794 (N_25794,N_24604,N_25029);
xnor U25795 (N_25795,N_24719,N_24813);
nand U25796 (N_25796,N_24805,N_24736);
nand U25797 (N_25797,N_24691,N_24778);
or U25798 (N_25798,N_24977,N_24743);
or U25799 (N_25799,N_24927,N_24817);
and U25800 (N_25800,N_25532,N_25242);
nand U25801 (N_25801,N_25456,N_25332);
or U25802 (N_25802,N_25607,N_25689);
nor U25803 (N_25803,N_25714,N_25270);
nand U25804 (N_25804,N_25454,N_25572);
or U25805 (N_25805,N_25288,N_25351);
nor U25806 (N_25806,N_25387,N_25752);
nand U25807 (N_25807,N_25558,N_25368);
nor U25808 (N_25808,N_25416,N_25415);
nor U25809 (N_25809,N_25372,N_25531);
nor U25810 (N_25810,N_25510,N_25629);
nor U25811 (N_25811,N_25243,N_25560);
or U25812 (N_25812,N_25796,N_25321);
and U25813 (N_25813,N_25487,N_25502);
and U25814 (N_25814,N_25644,N_25514);
or U25815 (N_25815,N_25413,N_25300);
or U25816 (N_25816,N_25423,N_25621);
nor U25817 (N_25817,N_25706,N_25587);
and U25818 (N_25818,N_25218,N_25669);
nand U25819 (N_25819,N_25488,N_25449);
and U25820 (N_25820,N_25590,N_25767);
nand U25821 (N_25821,N_25260,N_25484);
or U25822 (N_25822,N_25769,N_25268);
or U25823 (N_25823,N_25734,N_25690);
nor U25824 (N_25824,N_25469,N_25526);
xnor U25825 (N_25825,N_25329,N_25278);
nand U25826 (N_25826,N_25762,N_25744);
xnor U25827 (N_25827,N_25655,N_25201);
nand U25828 (N_25828,N_25557,N_25408);
nand U25829 (N_25829,N_25682,N_25320);
nor U25830 (N_25830,N_25404,N_25637);
or U25831 (N_25831,N_25652,N_25516);
nor U25832 (N_25832,N_25610,N_25505);
nand U25833 (N_25833,N_25569,N_25729);
nor U25834 (N_25834,N_25639,N_25792);
and U25835 (N_25835,N_25246,N_25458);
xnor U25836 (N_25836,N_25707,N_25631);
nand U25837 (N_25837,N_25605,N_25463);
and U25838 (N_25838,N_25399,N_25548);
or U25839 (N_25839,N_25700,N_25654);
xnor U25840 (N_25840,N_25537,N_25584);
and U25841 (N_25841,N_25642,N_25742);
xnor U25842 (N_25842,N_25518,N_25779);
or U25843 (N_25843,N_25713,N_25710);
xnor U25844 (N_25844,N_25692,N_25496);
nor U25845 (N_25845,N_25539,N_25726);
nand U25846 (N_25846,N_25377,N_25773);
nor U25847 (N_25847,N_25738,N_25468);
or U25848 (N_25848,N_25325,N_25214);
or U25849 (N_25849,N_25438,N_25294);
and U25850 (N_25850,N_25527,N_25202);
or U25851 (N_25851,N_25418,N_25576);
and U25852 (N_25852,N_25676,N_25684);
nor U25853 (N_25853,N_25793,N_25254);
or U25854 (N_25854,N_25464,N_25618);
and U25855 (N_25855,N_25213,N_25210);
and U25856 (N_25856,N_25436,N_25765);
nand U25857 (N_25857,N_25562,N_25670);
xor U25858 (N_25858,N_25442,N_25285);
and U25859 (N_25859,N_25543,N_25704);
nand U25860 (N_25860,N_25381,N_25656);
xor U25861 (N_25861,N_25389,N_25613);
or U25862 (N_25862,N_25480,N_25289);
and U25863 (N_25863,N_25597,N_25358);
nand U25864 (N_25864,N_25225,N_25638);
nor U25865 (N_25865,N_25217,N_25386);
and U25866 (N_25866,N_25643,N_25318);
and U25867 (N_25867,N_25553,N_25309);
or U25868 (N_25868,N_25252,N_25360);
nor U25869 (N_25869,N_25785,N_25570);
and U25870 (N_25870,N_25237,N_25273);
and U25871 (N_25871,N_25312,N_25256);
nor U25872 (N_25872,N_25478,N_25675);
xnor U25873 (N_25873,N_25298,N_25588);
nand U25874 (N_25874,N_25427,N_25661);
nor U25875 (N_25875,N_25574,N_25739);
nand U25876 (N_25876,N_25794,N_25296);
and U25877 (N_25877,N_25228,N_25719);
xor U25878 (N_25878,N_25405,N_25374);
nand U25879 (N_25879,N_25559,N_25444);
and U25880 (N_25880,N_25786,N_25552);
nor U25881 (N_25881,N_25781,N_25671);
and U25882 (N_25882,N_25678,N_25303);
nand U25883 (N_25883,N_25315,N_25705);
nor U25884 (N_25884,N_25319,N_25275);
nand U25885 (N_25885,N_25503,N_25366);
and U25886 (N_25886,N_25263,N_25208);
xor U25887 (N_25887,N_25411,N_25595);
nand U25888 (N_25888,N_25730,N_25554);
and U25889 (N_25889,N_25340,N_25251);
xnor U25890 (N_25890,N_25533,N_25258);
nor U25891 (N_25891,N_25205,N_25271);
and U25892 (N_25892,N_25585,N_25625);
xor U25893 (N_25893,N_25627,N_25662);
nor U25894 (N_25894,N_25596,N_25754);
or U25895 (N_25895,N_25437,N_25339);
xor U25896 (N_25896,N_25619,N_25239);
nor U25897 (N_25897,N_25513,N_25265);
and U25898 (N_25898,N_25326,N_25474);
or U25899 (N_25899,N_25221,N_25261);
and U25900 (N_25900,N_25626,N_25733);
nand U25901 (N_25901,N_25407,N_25216);
nor U25902 (N_25902,N_25486,N_25666);
xor U25903 (N_25903,N_25720,N_25534);
or U25904 (N_25904,N_25245,N_25743);
xnor U25905 (N_25905,N_25780,N_25353);
nor U25906 (N_25906,N_25400,N_25519);
nand U25907 (N_25907,N_25264,N_25341);
and U25908 (N_25908,N_25598,N_25711);
or U25909 (N_25909,N_25520,N_25230);
nor U25910 (N_25910,N_25499,N_25555);
and U25911 (N_25911,N_25435,N_25453);
nand U25912 (N_25912,N_25757,N_25299);
or U25913 (N_25913,N_25591,N_25760);
nor U25914 (N_25914,N_25538,N_25628);
nand U25915 (N_25915,N_25316,N_25508);
nand U25916 (N_25916,N_25380,N_25363);
or U25917 (N_25917,N_25266,N_25592);
and U25918 (N_25918,N_25434,N_25623);
or U25919 (N_25919,N_25650,N_25732);
and U25920 (N_25920,N_25223,N_25566);
or U25921 (N_25921,N_25723,N_25493);
xor U25922 (N_25922,N_25203,N_25219);
nand U25923 (N_25923,N_25515,N_25336);
nand U25924 (N_25924,N_25349,N_25630);
xor U25925 (N_25925,N_25426,N_25641);
nand U25926 (N_25926,N_25660,N_25291);
nor U25927 (N_25927,N_25346,N_25716);
nor U25928 (N_25928,N_25753,N_25445);
nor U25929 (N_25929,N_25234,N_25582);
and U25930 (N_25930,N_25200,N_25211);
or U25931 (N_25931,N_25751,N_25479);
xor U25932 (N_25932,N_25451,N_25787);
nand U25933 (N_25933,N_25241,N_25390);
and U25934 (N_25934,N_25282,N_25718);
nor U25935 (N_25935,N_25540,N_25209);
nor U25936 (N_25936,N_25746,N_25798);
and U25937 (N_25937,N_25788,N_25778);
or U25938 (N_25938,N_25724,N_25494);
or U25939 (N_25939,N_25460,N_25364);
nor U25940 (N_25940,N_25401,N_25524);
and U25941 (N_25941,N_25640,N_25616);
xnor U25942 (N_25942,N_25267,N_25440);
and U25943 (N_25943,N_25735,N_25335);
nor U25944 (N_25944,N_25337,N_25477);
nor U25945 (N_25945,N_25653,N_25215);
xnor U25946 (N_25946,N_25233,N_25248);
nor U25947 (N_25947,N_25425,N_25568);
and U25948 (N_25948,N_25378,N_25565);
or U25949 (N_25949,N_25471,N_25799);
or U25950 (N_25950,N_25370,N_25546);
and U25951 (N_25951,N_25651,N_25693);
or U25952 (N_25952,N_25317,N_25314);
xor U25953 (N_25953,N_25287,N_25433);
or U25954 (N_25954,N_25284,N_25365);
or U25955 (N_25955,N_25331,N_25721);
or U25956 (N_25956,N_25511,N_25634);
and U25957 (N_25957,N_25338,N_25717);
or U25958 (N_25958,N_25699,N_25367);
xor U25959 (N_25959,N_25361,N_25668);
nor U25960 (N_25960,N_25279,N_25269);
and U25961 (N_25961,N_25485,N_25283);
and U25962 (N_25962,N_25632,N_25465);
and U25963 (N_25963,N_25775,N_25521);
nand U25964 (N_25964,N_25672,N_25412);
and U25965 (N_25965,N_25509,N_25310);
and U25966 (N_25966,N_25611,N_25549);
nor U25967 (N_25967,N_25530,N_25715);
or U25968 (N_25968,N_25280,N_25617);
nor U25969 (N_25969,N_25448,N_25747);
xor U25970 (N_25970,N_25419,N_25347);
nor U25971 (N_25971,N_25357,N_25204);
and U25972 (N_25972,N_25475,N_25677);
nor U25973 (N_25973,N_25541,N_25523);
nand U25974 (N_25974,N_25281,N_25712);
xnor U25975 (N_25975,N_25455,N_25304);
xnor U25976 (N_25976,N_25497,N_25323);
nor U25977 (N_25977,N_25355,N_25687);
and U25978 (N_25978,N_25741,N_25740);
nand U25979 (N_25979,N_25342,N_25681);
nand U25980 (N_25980,N_25750,N_25648);
nand U25981 (N_25981,N_25615,N_25709);
or U25982 (N_25982,N_25255,N_25601);
xor U25983 (N_25983,N_25447,N_25536);
nand U25984 (N_25984,N_25686,N_25581);
nand U25985 (N_25985,N_25306,N_25446);
nand U25986 (N_25986,N_25286,N_25575);
and U25987 (N_25987,N_25385,N_25535);
or U25988 (N_25988,N_25428,N_25473);
nor U25989 (N_25989,N_25795,N_25352);
or U25990 (N_25990,N_25439,N_25772);
xnor U25991 (N_25991,N_25667,N_25249);
nand U25992 (N_25992,N_25229,N_25602);
and U25993 (N_25993,N_25774,N_25647);
or U25994 (N_25994,N_25745,N_25222);
xnor U25995 (N_25995,N_25371,N_25220);
or U25996 (N_25996,N_25529,N_25685);
nand U25997 (N_25997,N_25356,N_25589);
or U25998 (N_25998,N_25573,N_25550);
xnor U25999 (N_25999,N_25292,N_25736);
or U26000 (N_26000,N_25253,N_25756);
xor U26001 (N_26001,N_25334,N_25244);
nand U26002 (N_26002,N_25790,N_25698);
nand U26003 (N_26003,N_25702,N_25580);
xnor U26004 (N_26004,N_25410,N_25556);
and U26005 (N_26005,N_25461,N_25207);
and U26006 (N_26006,N_25766,N_25771);
and U26007 (N_26007,N_25697,N_25344);
or U26008 (N_26008,N_25350,N_25633);
nor U26009 (N_26009,N_25295,N_25379);
nand U26010 (N_26010,N_25659,N_25276);
and U26011 (N_26011,N_25783,N_25545);
or U26012 (N_26012,N_25674,N_25476);
and U26013 (N_26013,N_25506,N_25422);
xnor U26014 (N_26014,N_25231,N_25235);
xor U26015 (N_26015,N_25376,N_25459);
and U26016 (N_26016,N_25250,N_25578);
nand U26017 (N_26017,N_25432,N_25722);
xnor U26018 (N_26018,N_25236,N_25583);
or U26019 (N_26019,N_25564,N_25563);
nand U26020 (N_26020,N_25593,N_25491);
and U26021 (N_26021,N_25257,N_25409);
nor U26022 (N_26022,N_25791,N_25470);
nand U26023 (N_26023,N_25259,N_25301);
and U26024 (N_26024,N_25624,N_25688);
nor U26025 (N_26025,N_25343,N_25481);
nand U26026 (N_26026,N_25482,N_25450);
or U26027 (N_26027,N_25322,N_25224);
nor U26028 (N_26028,N_25430,N_25397);
or U26029 (N_26029,N_25330,N_25606);
xor U26030 (N_26030,N_25517,N_25594);
xnor U26031 (N_26031,N_25636,N_25274);
and U26032 (N_26032,N_25749,N_25784);
and U26033 (N_26033,N_25696,N_25608);
nor U26034 (N_26034,N_25302,N_25457);
xnor U26035 (N_26035,N_25777,N_25761);
and U26036 (N_26036,N_25797,N_25240);
nor U26037 (N_26037,N_25232,N_25311);
xor U26038 (N_26038,N_25369,N_25424);
nand U26039 (N_26039,N_25759,N_25414);
nand U26040 (N_26040,N_25421,N_25748);
and U26041 (N_26041,N_25467,N_25402);
nand U26042 (N_26042,N_25649,N_25395);
nand U26043 (N_26043,N_25737,N_25388);
nor U26044 (N_26044,N_25441,N_25525);
nor U26045 (N_26045,N_25507,N_25603);
xnor U26046 (N_26046,N_25212,N_25247);
nor U26047 (N_26047,N_25665,N_25614);
and U26048 (N_26048,N_25492,N_25645);
or U26049 (N_26049,N_25620,N_25417);
or U26050 (N_26050,N_25683,N_25764);
nor U26051 (N_26051,N_25420,N_25472);
xnor U26052 (N_26052,N_25551,N_25561);
nor U26053 (N_26053,N_25622,N_25727);
nand U26054 (N_26054,N_25373,N_25443);
nand U26055 (N_26055,N_25577,N_25272);
or U26056 (N_26056,N_25393,N_25206);
and U26057 (N_26057,N_25579,N_25586);
nor U26058 (N_26058,N_25701,N_25227);
nand U26059 (N_26059,N_25359,N_25333);
xnor U26060 (N_26060,N_25680,N_25768);
xnor U26061 (N_26061,N_25462,N_25567);
or U26062 (N_26062,N_25658,N_25763);
nor U26063 (N_26063,N_25646,N_25544);
nor U26064 (N_26064,N_25277,N_25663);
nor U26065 (N_26065,N_25694,N_25297);
or U26066 (N_26066,N_25728,N_25290);
nor U26067 (N_26067,N_25345,N_25758);
nor U26068 (N_26068,N_25305,N_25635);
and U26069 (N_26069,N_25512,N_25354);
nor U26070 (N_26070,N_25504,N_25452);
nand U26071 (N_26071,N_25522,N_25262);
or U26072 (N_26072,N_25362,N_25600);
nand U26073 (N_26073,N_25490,N_25547);
and U26074 (N_26074,N_25398,N_25695);
nor U26075 (N_26075,N_25599,N_25392);
nor U26076 (N_26076,N_25429,N_25776);
and U26077 (N_26077,N_25238,N_25483);
xor U26078 (N_26078,N_25528,N_25226);
nor U26079 (N_26079,N_25348,N_25770);
or U26080 (N_26080,N_25375,N_25501);
xnor U26081 (N_26081,N_25431,N_25394);
or U26082 (N_26082,N_25679,N_25403);
xor U26083 (N_26083,N_25782,N_25391);
and U26084 (N_26084,N_25308,N_25489);
and U26085 (N_26085,N_25466,N_25703);
xor U26086 (N_26086,N_25542,N_25664);
xnor U26087 (N_26087,N_25384,N_25327);
or U26088 (N_26088,N_25673,N_25604);
xnor U26089 (N_26089,N_25731,N_25612);
xnor U26090 (N_26090,N_25406,N_25383);
xnor U26091 (N_26091,N_25657,N_25328);
and U26092 (N_26092,N_25725,N_25313);
and U26093 (N_26093,N_25609,N_25571);
xor U26094 (N_26094,N_25382,N_25396);
nand U26095 (N_26095,N_25324,N_25708);
xnor U26096 (N_26096,N_25789,N_25293);
nand U26097 (N_26097,N_25691,N_25500);
or U26098 (N_26098,N_25307,N_25498);
and U26099 (N_26099,N_25495,N_25755);
nand U26100 (N_26100,N_25383,N_25630);
xor U26101 (N_26101,N_25386,N_25528);
nand U26102 (N_26102,N_25430,N_25332);
or U26103 (N_26103,N_25239,N_25407);
nor U26104 (N_26104,N_25397,N_25662);
xor U26105 (N_26105,N_25316,N_25473);
nor U26106 (N_26106,N_25263,N_25549);
xor U26107 (N_26107,N_25412,N_25512);
and U26108 (N_26108,N_25696,N_25550);
nor U26109 (N_26109,N_25716,N_25552);
nand U26110 (N_26110,N_25517,N_25722);
or U26111 (N_26111,N_25767,N_25397);
xnor U26112 (N_26112,N_25260,N_25642);
nand U26113 (N_26113,N_25622,N_25329);
nor U26114 (N_26114,N_25227,N_25285);
and U26115 (N_26115,N_25275,N_25228);
nor U26116 (N_26116,N_25413,N_25412);
nand U26117 (N_26117,N_25745,N_25449);
nor U26118 (N_26118,N_25666,N_25314);
or U26119 (N_26119,N_25551,N_25514);
or U26120 (N_26120,N_25205,N_25632);
and U26121 (N_26121,N_25251,N_25357);
nor U26122 (N_26122,N_25586,N_25238);
xor U26123 (N_26123,N_25629,N_25427);
nand U26124 (N_26124,N_25208,N_25503);
nor U26125 (N_26125,N_25286,N_25784);
nor U26126 (N_26126,N_25367,N_25688);
nand U26127 (N_26127,N_25679,N_25731);
and U26128 (N_26128,N_25730,N_25634);
and U26129 (N_26129,N_25367,N_25438);
and U26130 (N_26130,N_25209,N_25422);
xnor U26131 (N_26131,N_25274,N_25560);
or U26132 (N_26132,N_25552,N_25398);
xor U26133 (N_26133,N_25286,N_25248);
or U26134 (N_26134,N_25696,N_25202);
and U26135 (N_26135,N_25274,N_25494);
or U26136 (N_26136,N_25709,N_25442);
nor U26137 (N_26137,N_25243,N_25356);
xnor U26138 (N_26138,N_25518,N_25412);
xor U26139 (N_26139,N_25662,N_25682);
and U26140 (N_26140,N_25639,N_25573);
and U26141 (N_26141,N_25273,N_25277);
xnor U26142 (N_26142,N_25427,N_25340);
nand U26143 (N_26143,N_25309,N_25432);
and U26144 (N_26144,N_25347,N_25700);
nor U26145 (N_26145,N_25209,N_25796);
xnor U26146 (N_26146,N_25714,N_25648);
nor U26147 (N_26147,N_25463,N_25662);
and U26148 (N_26148,N_25476,N_25537);
nor U26149 (N_26149,N_25701,N_25266);
or U26150 (N_26150,N_25334,N_25637);
nor U26151 (N_26151,N_25239,N_25517);
nand U26152 (N_26152,N_25723,N_25483);
nor U26153 (N_26153,N_25487,N_25420);
xnor U26154 (N_26154,N_25473,N_25747);
nor U26155 (N_26155,N_25480,N_25721);
xnor U26156 (N_26156,N_25439,N_25580);
xnor U26157 (N_26157,N_25768,N_25431);
nor U26158 (N_26158,N_25337,N_25399);
nand U26159 (N_26159,N_25388,N_25428);
xnor U26160 (N_26160,N_25678,N_25593);
xor U26161 (N_26161,N_25593,N_25258);
xor U26162 (N_26162,N_25783,N_25339);
and U26163 (N_26163,N_25573,N_25218);
and U26164 (N_26164,N_25626,N_25260);
nor U26165 (N_26165,N_25397,N_25661);
or U26166 (N_26166,N_25390,N_25255);
xor U26167 (N_26167,N_25223,N_25278);
nand U26168 (N_26168,N_25351,N_25462);
and U26169 (N_26169,N_25723,N_25440);
or U26170 (N_26170,N_25447,N_25611);
and U26171 (N_26171,N_25743,N_25585);
nor U26172 (N_26172,N_25285,N_25723);
xor U26173 (N_26173,N_25782,N_25457);
xor U26174 (N_26174,N_25297,N_25634);
or U26175 (N_26175,N_25486,N_25226);
or U26176 (N_26176,N_25345,N_25383);
nand U26177 (N_26177,N_25667,N_25437);
or U26178 (N_26178,N_25233,N_25633);
nor U26179 (N_26179,N_25547,N_25749);
nand U26180 (N_26180,N_25794,N_25741);
xor U26181 (N_26181,N_25707,N_25380);
nand U26182 (N_26182,N_25232,N_25297);
or U26183 (N_26183,N_25607,N_25308);
xnor U26184 (N_26184,N_25602,N_25251);
nor U26185 (N_26185,N_25504,N_25662);
nor U26186 (N_26186,N_25200,N_25665);
or U26187 (N_26187,N_25408,N_25312);
nand U26188 (N_26188,N_25745,N_25445);
or U26189 (N_26189,N_25563,N_25269);
and U26190 (N_26190,N_25650,N_25481);
nor U26191 (N_26191,N_25537,N_25278);
xor U26192 (N_26192,N_25708,N_25565);
xnor U26193 (N_26193,N_25296,N_25729);
nand U26194 (N_26194,N_25791,N_25393);
xnor U26195 (N_26195,N_25673,N_25588);
and U26196 (N_26196,N_25622,N_25265);
or U26197 (N_26197,N_25360,N_25209);
and U26198 (N_26198,N_25263,N_25548);
nand U26199 (N_26199,N_25501,N_25229);
nand U26200 (N_26200,N_25363,N_25475);
and U26201 (N_26201,N_25464,N_25272);
and U26202 (N_26202,N_25322,N_25526);
and U26203 (N_26203,N_25761,N_25313);
or U26204 (N_26204,N_25703,N_25627);
or U26205 (N_26205,N_25597,N_25259);
nand U26206 (N_26206,N_25585,N_25322);
nor U26207 (N_26207,N_25698,N_25215);
nor U26208 (N_26208,N_25557,N_25517);
nor U26209 (N_26209,N_25387,N_25259);
xnor U26210 (N_26210,N_25508,N_25206);
and U26211 (N_26211,N_25409,N_25283);
nand U26212 (N_26212,N_25564,N_25603);
and U26213 (N_26213,N_25599,N_25344);
or U26214 (N_26214,N_25742,N_25246);
or U26215 (N_26215,N_25207,N_25344);
and U26216 (N_26216,N_25392,N_25417);
and U26217 (N_26217,N_25284,N_25790);
or U26218 (N_26218,N_25441,N_25309);
and U26219 (N_26219,N_25765,N_25268);
or U26220 (N_26220,N_25446,N_25497);
or U26221 (N_26221,N_25735,N_25650);
or U26222 (N_26222,N_25268,N_25431);
xnor U26223 (N_26223,N_25785,N_25340);
nor U26224 (N_26224,N_25489,N_25451);
xnor U26225 (N_26225,N_25294,N_25430);
nand U26226 (N_26226,N_25370,N_25774);
nand U26227 (N_26227,N_25466,N_25653);
nor U26228 (N_26228,N_25451,N_25211);
or U26229 (N_26229,N_25534,N_25516);
xor U26230 (N_26230,N_25294,N_25360);
and U26231 (N_26231,N_25779,N_25707);
nor U26232 (N_26232,N_25578,N_25411);
xor U26233 (N_26233,N_25252,N_25297);
and U26234 (N_26234,N_25478,N_25244);
xnor U26235 (N_26235,N_25459,N_25401);
xor U26236 (N_26236,N_25740,N_25440);
or U26237 (N_26237,N_25337,N_25657);
or U26238 (N_26238,N_25461,N_25409);
nor U26239 (N_26239,N_25558,N_25650);
xnor U26240 (N_26240,N_25357,N_25711);
and U26241 (N_26241,N_25576,N_25311);
xnor U26242 (N_26242,N_25371,N_25417);
or U26243 (N_26243,N_25784,N_25411);
xnor U26244 (N_26244,N_25700,N_25471);
nand U26245 (N_26245,N_25509,N_25690);
or U26246 (N_26246,N_25627,N_25229);
xnor U26247 (N_26247,N_25470,N_25216);
or U26248 (N_26248,N_25413,N_25711);
xnor U26249 (N_26249,N_25659,N_25339);
xor U26250 (N_26250,N_25725,N_25536);
nand U26251 (N_26251,N_25443,N_25389);
xnor U26252 (N_26252,N_25708,N_25694);
or U26253 (N_26253,N_25278,N_25553);
nor U26254 (N_26254,N_25351,N_25338);
nor U26255 (N_26255,N_25261,N_25299);
nand U26256 (N_26256,N_25588,N_25296);
nor U26257 (N_26257,N_25729,N_25742);
nand U26258 (N_26258,N_25436,N_25309);
or U26259 (N_26259,N_25338,N_25404);
or U26260 (N_26260,N_25543,N_25378);
or U26261 (N_26261,N_25645,N_25424);
nand U26262 (N_26262,N_25723,N_25350);
or U26263 (N_26263,N_25357,N_25660);
nor U26264 (N_26264,N_25557,N_25414);
or U26265 (N_26265,N_25664,N_25347);
or U26266 (N_26266,N_25369,N_25611);
nand U26267 (N_26267,N_25216,N_25465);
or U26268 (N_26268,N_25742,N_25295);
nor U26269 (N_26269,N_25775,N_25250);
and U26270 (N_26270,N_25378,N_25671);
and U26271 (N_26271,N_25556,N_25670);
and U26272 (N_26272,N_25259,N_25630);
and U26273 (N_26273,N_25473,N_25659);
nor U26274 (N_26274,N_25345,N_25426);
nor U26275 (N_26275,N_25493,N_25365);
xnor U26276 (N_26276,N_25425,N_25328);
nor U26277 (N_26277,N_25791,N_25602);
xor U26278 (N_26278,N_25249,N_25413);
and U26279 (N_26279,N_25791,N_25211);
nor U26280 (N_26280,N_25297,N_25340);
xor U26281 (N_26281,N_25420,N_25608);
and U26282 (N_26282,N_25249,N_25716);
nor U26283 (N_26283,N_25558,N_25285);
or U26284 (N_26284,N_25766,N_25763);
or U26285 (N_26285,N_25521,N_25588);
nor U26286 (N_26286,N_25615,N_25661);
or U26287 (N_26287,N_25268,N_25454);
nor U26288 (N_26288,N_25564,N_25681);
nand U26289 (N_26289,N_25458,N_25701);
nand U26290 (N_26290,N_25778,N_25453);
nand U26291 (N_26291,N_25642,N_25785);
nor U26292 (N_26292,N_25253,N_25502);
xor U26293 (N_26293,N_25710,N_25221);
and U26294 (N_26294,N_25711,N_25787);
and U26295 (N_26295,N_25363,N_25420);
or U26296 (N_26296,N_25346,N_25494);
and U26297 (N_26297,N_25688,N_25519);
or U26298 (N_26298,N_25330,N_25730);
nor U26299 (N_26299,N_25429,N_25681);
nand U26300 (N_26300,N_25451,N_25207);
and U26301 (N_26301,N_25769,N_25220);
nor U26302 (N_26302,N_25463,N_25448);
nor U26303 (N_26303,N_25401,N_25344);
and U26304 (N_26304,N_25625,N_25439);
or U26305 (N_26305,N_25714,N_25394);
xnor U26306 (N_26306,N_25782,N_25362);
nand U26307 (N_26307,N_25235,N_25498);
nand U26308 (N_26308,N_25667,N_25492);
or U26309 (N_26309,N_25333,N_25671);
xnor U26310 (N_26310,N_25607,N_25486);
nor U26311 (N_26311,N_25494,N_25221);
and U26312 (N_26312,N_25512,N_25205);
xor U26313 (N_26313,N_25726,N_25667);
nand U26314 (N_26314,N_25334,N_25422);
nand U26315 (N_26315,N_25210,N_25527);
xnor U26316 (N_26316,N_25578,N_25726);
nand U26317 (N_26317,N_25408,N_25285);
nor U26318 (N_26318,N_25794,N_25463);
nor U26319 (N_26319,N_25719,N_25650);
nor U26320 (N_26320,N_25751,N_25555);
nand U26321 (N_26321,N_25430,N_25704);
nor U26322 (N_26322,N_25759,N_25346);
or U26323 (N_26323,N_25735,N_25700);
nor U26324 (N_26324,N_25442,N_25433);
and U26325 (N_26325,N_25437,N_25433);
or U26326 (N_26326,N_25785,N_25501);
or U26327 (N_26327,N_25309,N_25507);
nand U26328 (N_26328,N_25591,N_25429);
xnor U26329 (N_26329,N_25674,N_25305);
and U26330 (N_26330,N_25464,N_25741);
or U26331 (N_26331,N_25434,N_25667);
xnor U26332 (N_26332,N_25644,N_25283);
nor U26333 (N_26333,N_25522,N_25342);
nor U26334 (N_26334,N_25462,N_25530);
nand U26335 (N_26335,N_25487,N_25354);
nor U26336 (N_26336,N_25200,N_25610);
nand U26337 (N_26337,N_25251,N_25413);
and U26338 (N_26338,N_25692,N_25202);
nand U26339 (N_26339,N_25396,N_25744);
or U26340 (N_26340,N_25557,N_25441);
xor U26341 (N_26341,N_25555,N_25722);
nor U26342 (N_26342,N_25304,N_25537);
nor U26343 (N_26343,N_25798,N_25704);
nand U26344 (N_26344,N_25274,N_25292);
nor U26345 (N_26345,N_25242,N_25715);
and U26346 (N_26346,N_25502,N_25364);
nor U26347 (N_26347,N_25774,N_25781);
and U26348 (N_26348,N_25450,N_25544);
or U26349 (N_26349,N_25756,N_25507);
nor U26350 (N_26350,N_25708,N_25521);
nor U26351 (N_26351,N_25714,N_25224);
and U26352 (N_26352,N_25471,N_25633);
xor U26353 (N_26353,N_25633,N_25318);
nand U26354 (N_26354,N_25404,N_25657);
or U26355 (N_26355,N_25295,N_25728);
nor U26356 (N_26356,N_25284,N_25230);
or U26357 (N_26357,N_25254,N_25294);
nor U26358 (N_26358,N_25422,N_25378);
nand U26359 (N_26359,N_25271,N_25765);
nand U26360 (N_26360,N_25599,N_25532);
and U26361 (N_26361,N_25774,N_25794);
or U26362 (N_26362,N_25537,N_25758);
nand U26363 (N_26363,N_25655,N_25544);
nor U26364 (N_26364,N_25722,N_25473);
nand U26365 (N_26365,N_25610,N_25411);
nor U26366 (N_26366,N_25301,N_25316);
or U26367 (N_26367,N_25314,N_25343);
or U26368 (N_26368,N_25613,N_25352);
and U26369 (N_26369,N_25255,N_25265);
nand U26370 (N_26370,N_25283,N_25357);
or U26371 (N_26371,N_25379,N_25373);
xnor U26372 (N_26372,N_25559,N_25529);
nand U26373 (N_26373,N_25226,N_25417);
or U26374 (N_26374,N_25520,N_25530);
and U26375 (N_26375,N_25341,N_25305);
or U26376 (N_26376,N_25359,N_25342);
xnor U26377 (N_26377,N_25527,N_25343);
or U26378 (N_26378,N_25607,N_25669);
or U26379 (N_26379,N_25308,N_25735);
nor U26380 (N_26380,N_25667,N_25469);
xor U26381 (N_26381,N_25254,N_25561);
and U26382 (N_26382,N_25482,N_25325);
xnor U26383 (N_26383,N_25787,N_25790);
nand U26384 (N_26384,N_25675,N_25793);
xor U26385 (N_26385,N_25266,N_25549);
nor U26386 (N_26386,N_25787,N_25486);
nor U26387 (N_26387,N_25222,N_25450);
nor U26388 (N_26388,N_25401,N_25741);
nand U26389 (N_26389,N_25284,N_25275);
or U26390 (N_26390,N_25613,N_25263);
nand U26391 (N_26391,N_25559,N_25774);
xor U26392 (N_26392,N_25632,N_25284);
nor U26393 (N_26393,N_25684,N_25715);
or U26394 (N_26394,N_25508,N_25284);
and U26395 (N_26395,N_25559,N_25578);
nand U26396 (N_26396,N_25229,N_25671);
and U26397 (N_26397,N_25700,N_25314);
nand U26398 (N_26398,N_25297,N_25720);
nor U26399 (N_26399,N_25788,N_25320);
nor U26400 (N_26400,N_26302,N_26043);
xnor U26401 (N_26401,N_26224,N_25986);
nor U26402 (N_26402,N_26367,N_25991);
and U26403 (N_26403,N_26132,N_26119);
and U26404 (N_26404,N_26351,N_25882);
nand U26405 (N_26405,N_26156,N_25983);
nor U26406 (N_26406,N_25917,N_25998);
nor U26407 (N_26407,N_26110,N_26262);
nor U26408 (N_26408,N_26317,N_26344);
and U26409 (N_26409,N_26244,N_26106);
nand U26410 (N_26410,N_26188,N_26009);
or U26411 (N_26411,N_26363,N_26255);
nand U26412 (N_26412,N_26118,N_25818);
and U26413 (N_26413,N_26096,N_25930);
and U26414 (N_26414,N_26207,N_25895);
nand U26415 (N_26415,N_26082,N_26340);
nor U26416 (N_26416,N_26274,N_25836);
xor U26417 (N_26417,N_25929,N_25832);
or U26418 (N_26418,N_26240,N_25972);
xor U26419 (N_26419,N_25827,N_25934);
nor U26420 (N_26420,N_25921,N_25888);
nor U26421 (N_26421,N_26375,N_26273);
xor U26422 (N_26422,N_25822,N_26296);
or U26423 (N_26423,N_26384,N_25813);
nand U26424 (N_26424,N_25865,N_25812);
and U26425 (N_26425,N_26270,N_26383);
nor U26426 (N_26426,N_26256,N_25871);
xor U26427 (N_26427,N_26216,N_26307);
nand U26428 (N_26428,N_26086,N_26194);
xnor U26429 (N_26429,N_26048,N_25966);
or U26430 (N_26430,N_26233,N_26231);
or U26431 (N_26431,N_26292,N_25840);
or U26432 (N_26432,N_26228,N_26271);
xnor U26433 (N_26433,N_25994,N_25869);
and U26434 (N_26434,N_26394,N_25946);
and U26435 (N_26435,N_25807,N_26331);
or U26436 (N_26436,N_26312,N_25941);
xnor U26437 (N_26437,N_25811,N_26095);
xor U26438 (N_26438,N_25896,N_25876);
nor U26439 (N_26439,N_25906,N_26018);
nand U26440 (N_26440,N_25849,N_25874);
and U26441 (N_26441,N_26191,N_25916);
nand U26442 (N_26442,N_26392,N_26362);
xnor U26443 (N_26443,N_26075,N_26254);
nor U26444 (N_26444,N_26301,N_26235);
nor U26445 (N_26445,N_26014,N_25846);
and U26446 (N_26446,N_26126,N_25875);
nand U26447 (N_26447,N_25988,N_26354);
or U26448 (N_26448,N_25961,N_25877);
nand U26449 (N_26449,N_25959,N_26315);
and U26450 (N_26450,N_25801,N_26068);
and U26451 (N_26451,N_26381,N_26136);
xnor U26452 (N_26452,N_25843,N_25945);
nor U26453 (N_26453,N_25937,N_25940);
xnor U26454 (N_26454,N_26109,N_26006);
and U26455 (N_26455,N_26389,N_25868);
nand U26456 (N_26456,N_25978,N_25815);
xor U26457 (N_26457,N_26275,N_26388);
or U26458 (N_26458,N_25808,N_26304);
and U26459 (N_26459,N_25954,N_25928);
nand U26460 (N_26460,N_25838,N_26376);
and U26461 (N_26461,N_26398,N_26158);
and U26462 (N_26462,N_26290,N_26115);
nor U26463 (N_26463,N_25873,N_26030);
or U26464 (N_26464,N_26034,N_26064);
and U26465 (N_26465,N_26140,N_26120);
nand U26466 (N_26466,N_25977,N_26121);
xor U26467 (N_26467,N_26349,N_26322);
nor U26468 (N_26468,N_26298,N_26316);
or U26469 (N_26469,N_25802,N_26143);
and U26470 (N_26470,N_26151,N_25913);
nand U26471 (N_26471,N_26090,N_25855);
xor U26472 (N_26472,N_26360,N_26092);
and U26473 (N_26473,N_26278,N_25830);
xnor U26474 (N_26474,N_25850,N_25953);
nor U26475 (N_26475,N_25950,N_26167);
nor U26476 (N_26476,N_26153,N_26159);
and U26477 (N_26477,N_26370,N_26016);
nor U26478 (N_26478,N_26348,N_26102);
and U26479 (N_26479,N_26027,N_26123);
xnor U26480 (N_26480,N_26220,N_26038);
or U26481 (N_26481,N_25984,N_26393);
xor U26482 (N_26482,N_26072,N_26071);
xnor U26483 (N_26483,N_25826,N_25975);
xnor U26484 (N_26484,N_26347,N_26020);
and U26485 (N_26485,N_26265,N_26236);
xnor U26486 (N_26486,N_26280,N_26223);
xnor U26487 (N_26487,N_25878,N_26077);
xor U26488 (N_26488,N_26341,N_26088);
and U26489 (N_26489,N_26085,N_26277);
xor U26490 (N_26490,N_26033,N_26154);
nand U26491 (N_26491,N_26229,N_25829);
xnor U26492 (N_26492,N_25870,N_25824);
and U26493 (N_26493,N_26365,N_26319);
and U26494 (N_26494,N_26287,N_26028);
nand U26495 (N_26495,N_26031,N_25881);
or U26496 (N_26496,N_26323,N_25823);
xor U26497 (N_26497,N_25989,N_26128);
or U26498 (N_26498,N_26380,N_25804);
or U26499 (N_26499,N_25938,N_26013);
or U26500 (N_26500,N_25819,N_26008);
xnor U26501 (N_26501,N_26172,N_26382);
xor U26502 (N_26502,N_26177,N_26239);
and U26503 (N_26503,N_26147,N_26232);
or U26504 (N_26504,N_26185,N_26299);
nand U26505 (N_26505,N_26378,N_26134);
and U26506 (N_26506,N_26142,N_26002);
nor U26507 (N_26507,N_26192,N_25885);
nand U26508 (N_26508,N_26345,N_26005);
and U26509 (N_26509,N_26163,N_26122);
nand U26510 (N_26510,N_25936,N_26133);
xnor U26511 (N_26511,N_26291,N_26141);
and U26512 (N_26512,N_26035,N_26368);
nand U26513 (N_26513,N_25920,N_25963);
or U26514 (N_26514,N_26117,N_25833);
nor U26515 (N_26515,N_25919,N_26385);
nand U26516 (N_26516,N_26197,N_26281);
nor U26517 (N_26517,N_26210,N_26359);
or U26518 (N_26518,N_26173,N_25842);
or U26519 (N_26519,N_25862,N_25814);
and U26520 (N_26520,N_26138,N_25837);
nand U26521 (N_26521,N_26250,N_26285);
xor U26522 (N_26522,N_25987,N_26337);
nor U26523 (N_26523,N_25912,N_26045);
or U26524 (N_26524,N_25944,N_26130);
and U26525 (N_26525,N_25957,N_25962);
nand U26526 (N_26526,N_26047,N_26333);
and U26527 (N_26527,N_25853,N_26000);
nand U26528 (N_26528,N_26076,N_25973);
nor U26529 (N_26529,N_25817,N_25828);
nor U26530 (N_26530,N_25904,N_26377);
and U26531 (N_26531,N_26361,N_26097);
nor U26532 (N_26532,N_26019,N_26248);
nor U26533 (N_26533,N_25816,N_26001);
or U26534 (N_26534,N_25982,N_26037);
nand U26535 (N_26535,N_26293,N_26079);
xor U26536 (N_26536,N_26314,N_26024);
or U26537 (N_26537,N_26352,N_25805);
or U26538 (N_26538,N_26335,N_26057);
and U26539 (N_26539,N_25861,N_26054);
nand U26540 (N_26540,N_26157,N_26003);
or U26541 (N_26541,N_25948,N_26330);
xnor U26542 (N_26542,N_26311,N_26198);
or U26543 (N_26543,N_26056,N_25935);
nand U26544 (N_26544,N_26284,N_26282);
or U26545 (N_26545,N_25859,N_25910);
xnor U26546 (N_26546,N_26036,N_26346);
and U26547 (N_26547,N_26395,N_26321);
xor U26548 (N_26548,N_26225,N_26084);
nand U26549 (N_26549,N_25883,N_26358);
and U26550 (N_26550,N_26234,N_25899);
nand U26551 (N_26551,N_26253,N_26397);
xor U26552 (N_26552,N_26227,N_26300);
xor U26553 (N_26553,N_26139,N_26135);
xnor U26554 (N_26554,N_26243,N_26066);
and U26555 (N_26555,N_26238,N_26325);
nor U26556 (N_26556,N_25857,N_26164);
and U26557 (N_26557,N_26053,N_26355);
nand U26558 (N_26558,N_26187,N_25890);
and U26559 (N_26559,N_26369,N_26241);
nor U26560 (N_26560,N_25858,N_26252);
and U26561 (N_26561,N_25851,N_26386);
and U26562 (N_26562,N_26218,N_26230);
nand U26563 (N_26563,N_26065,N_26182);
xnor U26564 (N_26564,N_26087,N_26204);
and U26565 (N_26565,N_26168,N_26012);
xor U26566 (N_26566,N_26171,N_26170);
or U26567 (N_26567,N_26372,N_25911);
xor U26568 (N_26568,N_26181,N_26101);
xnor U26569 (N_26569,N_26026,N_26387);
xor U26570 (N_26570,N_25803,N_25997);
nand U26571 (N_26571,N_26371,N_26129);
xor U26572 (N_26572,N_26144,N_25810);
or U26573 (N_26573,N_25974,N_26226);
nor U26574 (N_26574,N_25964,N_25951);
or U26575 (N_26575,N_25981,N_25947);
nor U26576 (N_26576,N_26112,N_26195);
and U26577 (N_26577,N_25864,N_26149);
nand U26578 (N_26578,N_26203,N_26089);
nand U26579 (N_26579,N_26334,N_26353);
nand U26580 (N_26580,N_26217,N_26247);
and U26581 (N_26581,N_26306,N_25893);
nand U26582 (N_26582,N_25965,N_26189);
or U26583 (N_26583,N_26070,N_25955);
xor U26584 (N_26584,N_26276,N_25927);
nor U26585 (N_26585,N_25902,N_25852);
xnor U26586 (N_26586,N_26391,N_26116);
xor U26587 (N_26587,N_26078,N_26124);
nor U26588 (N_26588,N_25900,N_26100);
xor U26589 (N_26589,N_26356,N_26327);
nor U26590 (N_26590,N_25915,N_26015);
or U26591 (N_26591,N_26329,N_26162);
and U26592 (N_26592,N_26199,N_25979);
nand U26593 (N_26593,N_26190,N_26039);
and U26594 (N_26594,N_26336,N_25926);
xor U26595 (N_26595,N_26127,N_26309);
nand U26596 (N_26596,N_26050,N_26041);
and U26597 (N_26597,N_26155,N_26399);
xor U26598 (N_26598,N_26152,N_26258);
or U26599 (N_26599,N_25990,N_26094);
nand U26600 (N_26600,N_26073,N_25939);
or U26601 (N_26601,N_25914,N_26104);
nor U26602 (N_26602,N_26193,N_25866);
and U26603 (N_26603,N_26267,N_26074);
and U26604 (N_26604,N_26011,N_26313);
or U26605 (N_26605,N_25847,N_26080);
nor U26606 (N_26606,N_25894,N_26214);
or U26607 (N_26607,N_25806,N_26205);
xor U26608 (N_26608,N_25886,N_26350);
and U26609 (N_26609,N_25903,N_26289);
nand U26610 (N_26610,N_26390,N_25845);
and U26611 (N_26611,N_25901,N_25943);
or U26612 (N_26612,N_26324,N_26251);
or U26613 (N_26613,N_26113,N_25854);
or U26614 (N_26614,N_26021,N_26206);
nor U26615 (N_26615,N_25985,N_26342);
and U26616 (N_26616,N_26175,N_26286);
nand U26617 (N_26617,N_26269,N_25992);
nand U26618 (N_26618,N_26111,N_25993);
and U26619 (N_26619,N_26176,N_25831);
or U26620 (N_26620,N_26046,N_26067);
or U26621 (N_26621,N_26137,N_25924);
nand U26622 (N_26622,N_25925,N_25970);
nor U26623 (N_26623,N_25967,N_25860);
and U26624 (N_26624,N_25949,N_26017);
nand U26625 (N_26625,N_26261,N_26029);
nor U26626 (N_26626,N_26328,N_25891);
nor U26627 (N_26627,N_26264,N_26108);
and U26628 (N_26628,N_25999,N_25848);
nand U26629 (N_26629,N_26186,N_25996);
or U26630 (N_26630,N_26055,N_26215);
nand U26631 (N_26631,N_26007,N_26366);
and U26632 (N_26632,N_26196,N_26211);
or U26633 (N_26633,N_25809,N_26069);
or U26634 (N_26634,N_26145,N_26081);
nand U26635 (N_26635,N_26212,N_26260);
nand U26636 (N_26636,N_25976,N_26279);
xor U26637 (N_26637,N_26059,N_26040);
nor U26638 (N_26638,N_26242,N_26326);
or U26639 (N_26639,N_26208,N_25905);
or U26640 (N_26640,N_25821,N_25909);
nor U26641 (N_26641,N_26297,N_26184);
nand U26642 (N_26642,N_26052,N_26310);
nor U26643 (N_26643,N_25907,N_26263);
xnor U26644 (N_26644,N_25971,N_25892);
nor U26645 (N_26645,N_26178,N_26219);
and U26646 (N_26646,N_26379,N_26098);
xnor U26647 (N_26647,N_25931,N_26245);
nand U26648 (N_26648,N_26374,N_25863);
nand U26649 (N_26649,N_25872,N_26103);
xnor U26650 (N_26650,N_26060,N_26396);
xnor U26651 (N_26651,N_26364,N_25800);
xor U26652 (N_26652,N_26022,N_25867);
nor U26653 (N_26653,N_26343,N_26161);
nor U26654 (N_26654,N_25880,N_26010);
nor U26655 (N_26655,N_26025,N_25995);
nor U26656 (N_26656,N_25889,N_26357);
nand U26657 (N_26657,N_26174,N_26042);
nand U26658 (N_26658,N_26166,N_26023);
xnor U26659 (N_26659,N_26051,N_26201);
nand U26660 (N_26660,N_25968,N_26107);
xor U26661 (N_26661,N_26202,N_25898);
xnor U26662 (N_26662,N_25908,N_26180);
and U26663 (N_26663,N_26288,N_26165);
xnor U26664 (N_26664,N_26318,N_26062);
xnor U26665 (N_26665,N_26179,N_25834);
and U26666 (N_26666,N_26338,N_25879);
xnor U26667 (N_26667,N_25844,N_25884);
nand U26668 (N_26668,N_26246,N_26004);
and U26669 (N_26669,N_26049,N_26266);
xor U26670 (N_26670,N_25918,N_26308);
and U26671 (N_26671,N_26063,N_25825);
nand U26672 (N_26672,N_26249,N_25969);
or U26673 (N_26673,N_26213,N_26294);
nand U26674 (N_26674,N_26125,N_26283);
and U26675 (N_26675,N_26268,N_25820);
or U26676 (N_26676,N_26131,N_26091);
nand U26677 (N_26677,N_25958,N_26339);
xor U26678 (N_26678,N_25922,N_26114);
nand U26679 (N_26679,N_25960,N_25897);
xor U26680 (N_26680,N_26200,N_26160);
nor U26681 (N_26681,N_26099,N_26332);
nor U26682 (N_26682,N_25952,N_26209);
nor U26683 (N_26683,N_25980,N_26105);
nand U26684 (N_26684,N_26061,N_26032);
nor U26685 (N_26685,N_26169,N_25856);
and U26686 (N_26686,N_26272,N_26295);
xnor U26687 (N_26687,N_26373,N_26058);
and U26688 (N_26688,N_26044,N_25933);
nor U26689 (N_26689,N_25956,N_26237);
xnor U26690 (N_26690,N_26222,N_26221);
and U26691 (N_26691,N_26146,N_26150);
nor U26692 (N_26692,N_26305,N_26148);
and U26693 (N_26693,N_25841,N_25932);
nor U26694 (N_26694,N_25839,N_26257);
nand U26695 (N_26695,N_26093,N_25835);
or U26696 (N_26696,N_26183,N_26320);
xor U26697 (N_26697,N_26083,N_25942);
nor U26698 (N_26698,N_25887,N_26259);
nand U26699 (N_26699,N_26303,N_25923);
or U26700 (N_26700,N_26111,N_25858);
nor U26701 (N_26701,N_25834,N_26399);
or U26702 (N_26702,N_26027,N_25831);
nand U26703 (N_26703,N_25800,N_25903);
and U26704 (N_26704,N_26314,N_26135);
nand U26705 (N_26705,N_25826,N_26296);
nor U26706 (N_26706,N_25906,N_26343);
nor U26707 (N_26707,N_26121,N_26090);
or U26708 (N_26708,N_26094,N_26366);
and U26709 (N_26709,N_25944,N_26140);
xor U26710 (N_26710,N_26306,N_26278);
and U26711 (N_26711,N_26249,N_25916);
nand U26712 (N_26712,N_26117,N_25906);
and U26713 (N_26713,N_26364,N_26044);
xor U26714 (N_26714,N_26028,N_26132);
or U26715 (N_26715,N_26387,N_25821);
or U26716 (N_26716,N_26036,N_26167);
or U26717 (N_26717,N_25851,N_26388);
nand U26718 (N_26718,N_26178,N_26199);
and U26719 (N_26719,N_26055,N_26059);
nand U26720 (N_26720,N_26252,N_25977);
nand U26721 (N_26721,N_26216,N_26093);
nand U26722 (N_26722,N_26296,N_26365);
nor U26723 (N_26723,N_25866,N_26158);
or U26724 (N_26724,N_26324,N_26170);
or U26725 (N_26725,N_25816,N_26356);
and U26726 (N_26726,N_26223,N_26020);
and U26727 (N_26727,N_26239,N_26373);
nor U26728 (N_26728,N_26149,N_26082);
or U26729 (N_26729,N_26138,N_25984);
and U26730 (N_26730,N_26271,N_26384);
and U26731 (N_26731,N_26196,N_26269);
nand U26732 (N_26732,N_25836,N_26200);
and U26733 (N_26733,N_25877,N_26032);
nor U26734 (N_26734,N_25861,N_26022);
or U26735 (N_26735,N_26276,N_26219);
or U26736 (N_26736,N_26049,N_25849);
nand U26737 (N_26737,N_26219,N_25937);
nor U26738 (N_26738,N_26052,N_26143);
and U26739 (N_26739,N_26220,N_26226);
xor U26740 (N_26740,N_26213,N_25956);
or U26741 (N_26741,N_26107,N_25844);
or U26742 (N_26742,N_26085,N_25879);
nor U26743 (N_26743,N_26041,N_26184);
or U26744 (N_26744,N_25843,N_25907);
or U26745 (N_26745,N_26074,N_26104);
and U26746 (N_26746,N_26202,N_26027);
and U26747 (N_26747,N_26228,N_26036);
nand U26748 (N_26748,N_25821,N_25891);
and U26749 (N_26749,N_26089,N_25932);
or U26750 (N_26750,N_25801,N_26042);
nor U26751 (N_26751,N_26089,N_26386);
or U26752 (N_26752,N_26309,N_26117);
and U26753 (N_26753,N_25903,N_26177);
or U26754 (N_26754,N_25960,N_26387);
and U26755 (N_26755,N_25819,N_26177);
nand U26756 (N_26756,N_26286,N_26035);
xnor U26757 (N_26757,N_26369,N_25873);
nand U26758 (N_26758,N_26102,N_25990);
nor U26759 (N_26759,N_26357,N_26325);
or U26760 (N_26760,N_25923,N_26183);
xnor U26761 (N_26761,N_25831,N_26226);
and U26762 (N_26762,N_26155,N_26054);
or U26763 (N_26763,N_25816,N_26216);
nor U26764 (N_26764,N_26115,N_26101);
xnor U26765 (N_26765,N_26149,N_25860);
and U26766 (N_26766,N_26051,N_26353);
or U26767 (N_26767,N_26383,N_25821);
and U26768 (N_26768,N_26262,N_26057);
nand U26769 (N_26769,N_26178,N_26277);
and U26770 (N_26770,N_26366,N_26134);
nor U26771 (N_26771,N_25902,N_26216);
nor U26772 (N_26772,N_26289,N_25972);
nor U26773 (N_26773,N_25804,N_25822);
xor U26774 (N_26774,N_26063,N_26382);
nor U26775 (N_26775,N_26176,N_26166);
xor U26776 (N_26776,N_26066,N_26283);
or U26777 (N_26777,N_26134,N_26303);
xnor U26778 (N_26778,N_25964,N_26161);
nor U26779 (N_26779,N_26098,N_26224);
nand U26780 (N_26780,N_26080,N_26354);
and U26781 (N_26781,N_25934,N_26015);
or U26782 (N_26782,N_26083,N_26087);
xor U26783 (N_26783,N_25946,N_26370);
nor U26784 (N_26784,N_26260,N_25955);
xnor U26785 (N_26785,N_26046,N_26374);
nor U26786 (N_26786,N_25965,N_26302);
and U26787 (N_26787,N_26201,N_26375);
nor U26788 (N_26788,N_26399,N_25974);
xnor U26789 (N_26789,N_25857,N_25936);
or U26790 (N_26790,N_26215,N_26212);
and U26791 (N_26791,N_25865,N_26331);
nor U26792 (N_26792,N_25954,N_26168);
nor U26793 (N_26793,N_26264,N_26019);
or U26794 (N_26794,N_25883,N_25864);
xor U26795 (N_26795,N_26165,N_25884);
xnor U26796 (N_26796,N_26344,N_26376);
xnor U26797 (N_26797,N_26390,N_26235);
and U26798 (N_26798,N_26158,N_25948);
nand U26799 (N_26799,N_26371,N_25823);
nand U26800 (N_26800,N_25993,N_25826);
nand U26801 (N_26801,N_26159,N_26323);
and U26802 (N_26802,N_25840,N_26372);
and U26803 (N_26803,N_26253,N_26027);
and U26804 (N_26804,N_25835,N_25930);
nor U26805 (N_26805,N_26128,N_26239);
nor U26806 (N_26806,N_26129,N_26128);
nand U26807 (N_26807,N_25874,N_26193);
nor U26808 (N_26808,N_26210,N_26156);
nor U26809 (N_26809,N_26155,N_26386);
nand U26810 (N_26810,N_26328,N_26076);
xor U26811 (N_26811,N_25940,N_26162);
nor U26812 (N_26812,N_26221,N_25917);
nor U26813 (N_26813,N_26209,N_25857);
nor U26814 (N_26814,N_26375,N_26129);
nand U26815 (N_26815,N_25874,N_26376);
nor U26816 (N_26816,N_26214,N_25837);
nor U26817 (N_26817,N_26275,N_25899);
or U26818 (N_26818,N_26008,N_26361);
nor U26819 (N_26819,N_26313,N_26063);
or U26820 (N_26820,N_25822,N_26186);
or U26821 (N_26821,N_26042,N_26311);
nor U26822 (N_26822,N_26380,N_26057);
and U26823 (N_26823,N_25931,N_25985);
nand U26824 (N_26824,N_26044,N_26365);
or U26825 (N_26825,N_25958,N_26146);
xor U26826 (N_26826,N_25827,N_25864);
nand U26827 (N_26827,N_26350,N_26005);
nor U26828 (N_26828,N_26358,N_26025);
or U26829 (N_26829,N_25917,N_26255);
xnor U26830 (N_26830,N_26362,N_26255);
xor U26831 (N_26831,N_26253,N_25972);
nor U26832 (N_26832,N_25909,N_26269);
or U26833 (N_26833,N_25951,N_25931);
and U26834 (N_26834,N_25904,N_26061);
xor U26835 (N_26835,N_26020,N_25933);
nand U26836 (N_26836,N_25940,N_26151);
nor U26837 (N_26837,N_26318,N_26197);
nor U26838 (N_26838,N_25893,N_26355);
nor U26839 (N_26839,N_26038,N_25863);
nor U26840 (N_26840,N_26014,N_26060);
nor U26841 (N_26841,N_25853,N_26072);
and U26842 (N_26842,N_26039,N_25887);
nand U26843 (N_26843,N_26170,N_26309);
nand U26844 (N_26844,N_25900,N_26379);
or U26845 (N_26845,N_26254,N_26356);
or U26846 (N_26846,N_26352,N_26369);
nor U26847 (N_26847,N_26033,N_26308);
xnor U26848 (N_26848,N_26207,N_25988);
and U26849 (N_26849,N_25986,N_25805);
nand U26850 (N_26850,N_26301,N_26088);
or U26851 (N_26851,N_25863,N_26020);
and U26852 (N_26852,N_25827,N_25933);
or U26853 (N_26853,N_25813,N_26263);
nand U26854 (N_26854,N_26360,N_26378);
nor U26855 (N_26855,N_26028,N_25829);
nand U26856 (N_26856,N_26235,N_25917);
nor U26857 (N_26857,N_26069,N_25851);
xor U26858 (N_26858,N_25835,N_26384);
and U26859 (N_26859,N_26182,N_26315);
and U26860 (N_26860,N_25954,N_25917);
nor U26861 (N_26861,N_25986,N_26206);
nor U26862 (N_26862,N_26004,N_26041);
nand U26863 (N_26863,N_25905,N_26119);
nand U26864 (N_26864,N_26247,N_25810);
nor U26865 (N_26865,N_26258,N_25895);
or U26866 (N_26866,N_25828,N_25857);
nor U26867 (N_26867,N_26211,N_26065);
or U26868 (N_26868,N_26213,N_26136);
nand U26869 (N_26869,N_26172,N_26267);
nor U26870 (N_26870,N_26203,N_25941);
nand U26871 (N_26871,N_25835,N_26239);
nand U26872 (N_26872,N_25964,N_25829);
or U26873 (N_26873,N_25841,N_25821);
and U26874 (N_26874,N_26072,N_26158);
and U26875 (N_26875,N_25934,N_26123);
xnor U26876 (N_26876,N_26178,N_26134);
xnor U26877 (N_26877,N_25911,N_26030);
nand U26878 (N_26878,N_25996,N_26295);
or U26879 (N_26879,N_25993,N_26057);
and U26880 (N_26880,N_26185,N_26171);
nand U26881 (N_26881,N_26150,N_26367);
nor U26882 (N_26882,N_26185,N_25904);
nand U26883 (N_26883,N_26081,N_26334);
or U26884 (N_26884,N_26079,N_26191);
or U26885 (N_26885,N_26351,N_26016);
nand U26886 (N_26886,N_26053,N_26269);
nand U26887 (N_26887,N_26272,N_26354);
xnor U26888 (N_26888,N_26199,N_26004);
nand U26889 (N_26889,N_26270,N_26212);
and U26890 (N_26890,N_25817,N_25831);
or U26891 (N_26891,N_26345,N_25802);
or U26892 (N_26892,N_25987,N_26318);
nand U26893 (N_26893,N_26073,N_26017);
or U26894 (N_26894,N_25888,N_26093);
and U26895 (N_26895,N_26166,N_26077);
and U26896 (N_26896,N_26264,N_25990);
and U26897 (N_26897,N_26262,N_26249);
nand U26898 (N_26898,N_26071,N_26225);
nor U26899 (N_26899,N_26000,N_25887);
or U26900 (N_26900,N_26330,N_25842);
nor U26901 (N_26901,N_26312,N_26336);
or U26902 (N_26902,N_25877,N_26350);
nand U26903 (N_26903,N_26299,N_26308);
or U26904 (N_26904,N_26319,N_26041);
nor U26905 (N_26905,N_26378,N_26293);
nand U26906 (N_26906,N_26315,N_26039);
nand U26907 (N_26907,N_26337,N_26399);
xnor U26908 (N_26908,N_25807,N_25830);
nor U26909 (N_26909,N_26340,N_26026);
or U26910 (N_26910,N_26080,N_26246);
nand U26911 (N_26911,N_25891,N_26135);
xnor U26912 (N_26912,N_25953,N_26340);
and U26913 (N_26913,N_26015,N_26288);
xnor U26914 (N_26914,N_25809,N_25832);
and U26915 (N_26915,N_26079,N_26368);
nand U26916 (N_26916,N_25848,N_26311);
and U26917 (N_26917,N_26341,N_26362);
nand U26918 (N_26918,N_26284,N_26088);
xor U26919 (N_26919,N_26098,N_25951);
or U26920 (N_26920,N_26245,N_26283);
and U26921 (N_26921,N_25980,N_26093);
nand U26922 (N_26922,N_26201,N_25935);
and U26923 (N_26923,N_25945,N_25859);
nor U26924 (N_26924,N_26304,N_26058);
nand U26925 (N_26925,N_25837,N_26018);
and U26926 (N_26926,N_26166,N_26365);
nor U26927 (N_26927,N_26363,N_26325);
nand U26928 (N_26928,N_26000,N_26201);
nand U26929 (N_26929,N_26064,N_26054);
nand U26930 (N_26930,N_26151,N_26077);
xnor U26931 (N_26931,N_26349,N_26045);
or U26932 (N_26932,N_25814,N_25995);
or U26933 (N_26933,N_26291,N_25983);
nor U26934 (N_26934,N_25950,N_26308);
xnor U26935 (N_26935,N_26219,N_25924);
xor U26936 (N_26936,N_26271,N_25903);
or U26937 (N_26937,N_26241,N_25980);
xnor U26938 (N_26938,N_25806,N_26171);
and U26939 (N_26939,N_26334,N_26269);
xor U26940 (N_26940,N_25814,N_26073);
nor U26941 (N_26941,N_26111,N_26091);
or U26942 (N_26942,N_26286,N_25850);
and U26943 (N_26943,N_26210,N_26326);
nand U26944 (N_26944,N_25924,N_25826);
and U26945 (N_26945,N_26053,N_26145);
xnor U26946 (N_26946,N_25925,N_26313);
nand U26947 (N_26947,N_26269,N_26055);
nor U26948 (N_26948,N_25969,N_25987);
xor U26949 (N_26949,N_25924,N_25993);
and U26950 (N_26950,N_25803,N_26279);
nor U26951 (N_26951,N_26352,N_26136);
nor U26952 (N_26952,N_26235,N_26170);
or U26953 (N_26953,N_26386,N_26119);
and U26954 (N_26954,N_25864,N_26061);
nand U26955 (N_26955,N_26242,N_26337);
xor U26956 (N_26956,N_26138,N_26373);
or U26957 (N_26957,N_26236,N_26371);
or U26958 (N_26958,N_26357,N_26371);
and U26959 (N_26959,N_26306,N_25943);
and U26960 (N_26960,N_26274,N_25987);
or U26961 (N_26961,N_25819,N_26162);
xnor U26962 (N_26962,N_26185,N_26065);
nor U26963 (N_26963,N_26000,N_26276);
and U26964 (N_26964,N_25971,N_26385);
and U26965 (N_26965,N_26244,N_26393);
or U26966 (N_26966,N_25968,N_25883);
or U26967 (N_26967,N_25968,N_25998);
and U26968 (N_26968,N_26312,N_26126);
and U26969 (N_26969,N_26321,N_25927);
xnor U26970 (N_26970,N_26371,N_25808);
nand U26971 (N_26971,N_26241,N_26175);
nor U26972 (N_26972,N_26075,N_26044);
nand U26973 (N_26973,N_26312,N_25838);
nand U26974 (N_26974,N_26159,N_26283);
xor U26975 (N_26975,N_26398,N_26389);
and U26976 (N_26976,N_26279,N_26182);
or U26977 (N_26977,N_26277,N_26149);
xnor U26978 (N_26978,N_26249,N_25826);
nor U26979 (N_26979,N_26317,N_26198);
nand U26980 (N_26980,N_26300,N_26309);
and U26981 (N_26981,N_25961,N_26276);
xnor U26982 (N_26982,N_26011,N_25849);
or U26983 (N_26983,N_25961,N_26107);
nor U26984 (N_26984,N_26353,N_26315);
and U26985 (N_26985,N_26272,N_25930);
and U26986 (N_26986,N_25907,N_26354);
nand U26987 (N_26987,N_26353,N_25980);
nand U26988 (N_26988,N_26330,N_26364);
xnor U26989 (N_26989,N_26018,N_26209);
nand U26990 (N_26990,N_26164,N_25864);
and U26991 (N_26991,N_26375,N_26119);
xor U26992 (N_26992,N_25924,N_25969);
and U26993 (N_26993,N_26184,N_25933);
nand U26994 (N_26994,N_25989,N_26024);
and U26995 (N_26995,N_26224,N_26284);
and U26996 (N_26996,N_26156,N_26177);
nand U26997 (N_26997,N_26381,N_26338);
and U26998 (N_26998,N_25967,N_26263);
nand U26999 (N_26999,N_26056,N_25909);
nor U27000 (N_27000,N_26710,N_26812);
nand U27001 (N_27001,N_26897,N_26889);
nor U27002 (N_27002,N_26850,N_26949);
and U27003 (N_27003,N_26456,N_26938);
xnor U27004 (N_27004,N_26730,N_26828);
xor U27005 (N_27005,N_26965,N_26997);
nor U27006 (N_27006,N_26943,N_26811);
and U27007 (N_27007,N_26624,N_26603);
nor U27008 (N_27008,N_26962,N_26857);
nor U27009 (N_27009,N_26805,N_26854);
nor U27010 (N_27010,N_26879,N_26475);
nor U27011 (N_27011,N_26676,N_26816);
nand U27012 (N_27012,N_26584,N_26588);
xor U27013 (N_27013,N_26903,N_26551);
nand U27014 (N_27014,N_26982,N_26736);
and U27015 (N_27015,N_26958,N_26634);
or U27016 (N_27016,N_26685,N_26426);
or U27017 (N_27017,N_26725,N_26462);
xnor U27018 (N_27018,N_26771,N_26498);
or U27019 (N_27019,N_26919,N_26683);
or U27020 (N_27020,N_26450,N_26993);
and U27021 (N_27021,N_26642,N_26891);
xnor U27022 (N_27022,N_26988,N_26820);
nand U27023 (N_27023,N_26627,N_26984);
and U27024 (N_27024,N_26513,N_26434);
or U27025 (N_27025,N_26774,N_26468);
xnor U27026 (N_27026,N_26636,N_26616);
or U27027 (N_27027,N_26901,N_26872);
and U27028 (N_27028,N_26478,N_26795);
nor U27029 (N_27029,N_26966,N_26680);
nand U27030 (N_27030,N_26449,N_26444);
nand U27031 (N_27031,N_26959,N_26835);
or U27032 (N_27032,N_26998,N_26622);
xor U27033 (N_27033,N_26731,N_26798);
nor U27034 (N_27034,N_26803,N_26825);
xor U27035 (N_27035,N_26884,N_26840);
nor U27036 (N_27036,N_26712,N_26611);
and U27037 (N_27037,N_26418,N_26686);
or U27038 (N_27038,N_26651,N_26600);
or U27039 (N_27039,N_26987,N_26429);
xor U27040 (N_27040,N_26473,N_26727);
or U27041 (N_27041,N_26996,N_26869);
xor U27042 (N_27042,N_26920,N_26442);
or U27043 (N_27043,N_26635,N_26671);
and U27044 (N_27044,N_26494,N_26639);
xor U27045 (N_27045,N_26753,N_26930);
nor U27046 (N_27046,N_26519,N_26955);
xnor U27047 (N_27047,N_26660,N_26437);
and U27048 (N_27048,N_26617,N_26817);
or U27049 (N_27049,N_26488,N_26914);
or U27050 (N_27050,N_26575,N_26976);
nor U27051 (N_27051,N_26734,N_26907);
or U27052 (N_27052,N_26717,N_26654);
nor U27053 (N_27053,N_26610,N_26657);
nand U27054 (N_27054,N_26514,N_26496);
xnor U27055 (N_27055,N_26824,N_26497);
and U27056 (N_27056,N_26621,N_26916);
and U27057 (N_27057,N_26581,N_26947);
xnor U27058 (N_27058,N_26802,N_26793);
xnor U27059 (N_27059,N_26792,N_26438);
and U27060 (N_27060,N_26412,N_26750);
nand U27061 (N_27061,N_26618,N_26403);
and U27062 (N_27062,N_26841,N_26596);
nand U27063 (N_27063,N_26466,N_26928);
or U27064 (N_27064,N_26602,N_26439);
xor U27065 (N_27065,N_26870,N_26737);
xnor U27066 (N_27066,N_26667,N_26815);
xor U27067 (N_27067,N_26826,N_26855);
or U27068 (N_27068,N_26577,N_26886);
nor U27069 (N_27069,N_26760,N_26415);
nor U27070 (N_27070,N_26700,N_26784);
nor U27071 (N_27071,N_26493,N_26446);
nor U27072 (N_27072,N_26591,N_26791);
and U27073 (N_27073,N_26483,N_26648);
xor U27074 (N_27074,N_26666,N_26659);
or U27075 (N_27075,N_26451,N_26661);
and U27076 (N_27076,N_26909,N_26777);
nor U27077 (N_27077,N_26781,N_26650);
xnor U27078 (N_27078,N_26929,N_26945);
xor U27079 (N_27079,N_26923,N_26881);
or U27080 (N_27080,N_26453,N_26876);
nand U27081 (N_27081,N_26873,N_26709);
nand U27082 (N_27082,N_26428,N_26821);
or U27083 (N_27083,N_26833,N_26948);
and U27084 (N_27084,N_26590,N_26770);
or U27085 (N_27085,N_26754,N_26643);
xnor U27086 (N_27086,N_26932,N_26423);
xor U27087 (N_27087,N_26665,N_26492);
nand U27088 (N_27088,N_26924,N_26529);
or U27089 (N_27089,N_26527,N_26836);
nand U27090 (N_27090,N_26458,N_26986);
nand U27091 (N_27091,N_26677,N_26829);
and U27092 (N_27092,N_26411,N_26564);
and U27093 (N_27093,N_26888,N_26560);
nor U27094 (N_27094,N_26764,N_26799);
nand U27095 (N_27095,N_26539,N_26674);
nand U27096 (N_27096,N_26517,N_26559);
nand U27097 (N_27097,N_26556,N_26838);
nand U27098 (N_27098,N_26904,N_26406);
xnor U27099 (N_27099,N_26443,N_26510);
xor U27100 (N_27100,N_26804,N_26447);
xor U27101 (N_27101,N_26834,N_26892);
or U27102 (N_27102,N_26956,N_26688);
xnor U27103 (N_27103,N_26787,N_26819);
or U27104 (N_27104,N_26626,N_26578);
nor U27105 (N_27105,N_26615,N_26548);
nand U27106 (N_27106,N_26555,N_26504);
nand U27107 (N_27107,N_26663,N_26757);
nand U27108 (N_27108,N_26452,N_26655);
nand U27109 (N_27109,N_26552,N_26952);
and U27110 (N_27110,N_26946,N_26632);
xnor U27111 (N_27111,N_26936,N_26525);
or U27112 (N_27112,N_26613,N_26761);
xor U27113 (N_27113,N_26922,N_26703);
and U27114 (N_27114,N_26913,N_26720);
or U27115 (N_27115,N_26940,N_26668);
and U27116 (N_27116,N_26530,N_26574);
and U27117 (N_27117,N_26521,N_26482);
nor U27118 (N_27118,N_26424,N_26858);
and U27119 (N_27119,N_26404,N_26606);
or U27120 (N_27120,N_26441,N_26506);
or U27121 (N_27121,N_26706,N_26832);
or U27122 (N_27122,N_26601,N_26699);
nor U27123 (N_27123,N_26813,N_26417);
nand U27124 (N_27124,N_26557,N_26927);
nand U27125 (N_27125,N_26561,N_26973);
nor U27126 (N_27126,N_26896,N_26915);
nand U27127 (N_27127,N_26673,N_26522);
and U27128 (N_27128,N_26844,N_26895);
nor U27129 (N_27129,N_26851,N_26582);
and U27130 (N_27130,N_26520,N_26448);
and U27131 (N_27131,N_26689,N_26547);
xnor U27132 (N_27132,N_26465,N_26818);
and U27133 (N_27133,N_26431,N_26918);
nand U27134 (N_27134,N_26630,N_26460);
or U27135 (N_27135,N_26545,N_26868);
and U27136 (N_27136,N_26810,N_26741);
xor U27137 (N_27137,N_26491,N_26474);
xor U27138 (N_27138,N_26432,N_26528);
or U27139 (N_27139,N_26652,N_26427);
or U27140 (N_27140,N_26887,N_26692);
xor U27141 (N_27141,N_26598,N_26461);
and U27142 (N_27142,N_26806,N_26842);
nor U27143 (N_27143,N_26776,N_26664);
and U27144 (N_27144,N_26637,N_26723);
xor U27145 (N_27145,N_26587,N_26985);
nor U27146 (N_27146,N_26516,N_26779);
and U27147 (N_27147,N_26782,N_26569);
nor U27148 (N_27148,N_26524,N_26523);
nand U27149 (N_27149,N_26902,N_26526);
and U27150 (N_27150,N_26565,N_26794);
xnor U27151 (N_27151,N_26990,N_26535);
nand U27152 (N_27152,N_26808,N_26537);
and U27153 (N_27153,N_26682,N_26638);
nand U27154 (N_27154,N_26848,N_26900);
nor U27155 (N_27155,N_26463,N_26459);
nor U27156 (N_27156,N_26662,N_26540);
xnor U27157 (N_27157,N_26407,N_26687);
nand U27158 (N_27158,N_26963,N_26809);
nor U27159 (N_27159,N_26421,N_26908);
xnor U27160 (N_27160,N_26573,N_26653);
and U27161 (N_27161,N_26647,N_26981);
nand U27162 (N_27162,N_26935,N_26503);
xor U27163 (N_27163,N_26472,N_26684);
nor U27164 (N_27164,N_26735,N_26971);
xnor U27165 (N_27165,N_26464,N_26631);
nand U27166 (N_27166,N_26977,N_26675);
xor U27167 (N_27167,N_26999,N_26576);
nand U27168 (N_27168,N_26745,N_26430);
nand U27169 (N_27169,N_26856,N_26690);
nand U27170 (N_27170,N_26899,N_26845);
xnor U27171 (N_27171,N_26983,N_26501);
and U27172 (N_27172,N_26457,N_26507);
and U27173 (N_27173,N_26944,N_26589);
nor U27174 (N_27174,N_26558,N_26882);
and U27175 (N_27175,N_26477,N_26479);
nand U27176 (N_27176,N_26747,N_26553);
and U27177 (N_27177,N_26485,N_26486);
and U27178 (N_27178,N_26695,N_26681);
and U27179 (N_27179,N_26445,N_26738);
xnor U27180 (N_27180,N_26933,N_26402);
xor U27181 (N_27181,N_26612,N_26436);
nor U27182 (N_27182,N_26669,N_26707);
and U27183 (N_27183,N_26964,N_26866);
xor U27184 (N_27184,N_26954,N_26562);
nand U27185 (N_27185,N_26549,N_26495);
nand U27186 (N_27186,N_26619,N_26780);
nor U27187 (N_27187,N_26941,N_26629);
nand U27188 (N_27188,N_26672,N_26925);
nor U27189 (N_27189,N_26778,N_26785);
xor U27190 (N_27190,N_26843,N_26715);
and U27191 (N_27191,N_26583,N_26454);
nor U27192 (N_27192,N_26697,N_26801);
nor U27193 (N_27193,N_26620,N_26645);
nand U27194 (N_27194,N_26796,N_26623);
or U27195 (N_27195,N_26515,N_26509);
xor U27196 (N_27196,N_26847,N_26470);
nor U27197 (N_27197,N_26762,N_26679);
nand U27198 (N_27198,N_26566,N_26970);
and U27199 (N_27199,N_26658,N_26975);
or U27200 (N_27200,N_26786,N_26992);
xor U27201 (N_27201,N_26440,N_26435);
nand U27202 (N_27202,N_26512,N_26489);
xor U27203 (N_27203,N_26713,N_26740);
or U27204 (N_27204,N_26937,N_26532);
nor U27205 (N_27205,N_26580,N_26957);
and U27206 (N_27206,N_26646,N_26724);
and U27207 (N_27207,N_26701,N_26994);
or U27208 (N_27208,N_26849,N_26563);
xor U27209 (N_27209,N_26797,N_26921);
nor U27210 (N_27210,N_26862,N_26678);
nor U27211 (N_27211,N_26531,N_26773);
nor U27212 (N_27212,N_26830,N_26867);
nand U27213 (N_27213,N_26533,N_26865);
or U27214 (N_27214,N_26743,N_26732);
and U27215 (N_27215,N_26425,N_26972);
and U27216 (N_27216,N_26518,N_26586);
or U27217 (N_27217,N_26739,N_26550);
nor U27218 (N_27218,N_26728,N_26733);
and U27219 (N_27219,N_26831,N_26863);
xnor U27220 (N_27220,N_26894,N_26656);
and U27221 (N_27221,N_26538,N_26942);
xor U27222 (N_27222,N_26694,N_26505);
xor U27223 (N_27223,N_26726,N_26814);
xor U27224 (N_27224,N_26883,N_26716);
and U27225 (N_27225,N_26419,N_26481);
and U27226 (N_27226,N_26625,N_26934);
nor U27227 (N_27227,N_26742,N_26766);
nor U27228 (N_27228,N_26693,N_26570);
or U27229 (N_27229,N_26758,N_26974);
and U27230 (N_27230,N_26953,N_26641);
nand U27231 (N_27231,N_26413,N_26961);
nand U27232 (N_27232,N_26579,N_26544);
xor U27233 (N_27233,N_26400,N_26585);
xor U27234 (N_27234,N_26572,N_26871);
xnor U27235 (N_27235,N_26480,N_26765);
xor U27236 (N_27236,N_26751,N_26875);
or U27237 (N_27237,N_26846,N_26536);
and U27238 (N_27238,N_26749,N_26905);
xnor U27239 (N_27239,N_26542,N_26768);
or U27240 (N_27240,N_26752,N_26691);
or U27241 (N_27241,N_26410,N_26420);
xnor U27242 (N_27242,N_26860,N_26416);
or U27243 (N_27243,N_26789,N_26951);
or U27244 (N_27244,N_26877,N_26978);
nand U27245 (N_27245,N_26670,N_26790);
nand U27246 (N_27246,N_26769,N_26989);
or U27247 (N_27247,N_26775,N_26837);
xnor U27248 (N_27248,N_26960,N_26853);
and U27249 (N_27249,N_26729,N_26711);
nand U27250 (N_27250,N_26772,N_26939);
and U27251 (N_27251,N_26604,N_26609);
nor U27252 (N_27252,N_26823,N_26500);
nor U27253 (N_27253,N_26614,N_26783);
and U27254 (N_27254,N_26800,N_26696);
and U27255 (N_27255,N_26748,N_26911);
nor U27256 (N_27256,N_26718,N_26546);
nand U27257 (N_27257,N_26979,N_26839);
nand U27258 (N_27258,N_26893,N_26605);
nand U27259 (N_27259,N_26874,N_26788);
nor U27260 (N_27260,N_26405,N_26467);
xnor U27261 (N_27261,N_26571,N_26827);
nand U27262 (N_27262,N_26511,N_26926);
or U27263 (N_27263,N_26592,N_26422);
or U27264 (N_27264,N_26607,N_26859);
nand U27265 (N_27265,N_26471,N_26628);
xor U27266 (N_27266,N_26543,N_26567);
or U27267 (N_27267,N_26433,N_26499);
xnor U27268 (N_27268,N_26490,N_26597);
and U27269 (N_27269,N_26917,N_26755);
or U27270 (N_27270,N_26508,N_26608);
nor U27271 (N_27271,N_26861,N_26931);
nor U27272 (N_27272,N_26759,N_26991);
and U27273 (N_27273,N_26721,N_26950);
nand U27274 (N_27274,N_26714,N_26807);
or U27275 (N_27275,N_26640,N_26968);
nand U27276 (N_27276,N_26967,N_26649);
or U27277 (N_27277,N_26633,N_26593);
and U27278 (N_27278,N_26878,N_26704);
and U27279 (N_27279,N_26864,N_26408);
nor U27280 (N_27280,N_26469,N_26719);
or U27281 (N_27281,N_26906,N_26822);
nand U27282 (N_27282,N_26885,N_26409);
nand U27283 (N_27283,N_26910,N_26484);
nand U27284 (N_27284,N_26502,N_26969);
and U27285 (N_27285,N_26980,N_26487);
xnor U27286 (N_27286,N_26554,N_26595);
nand U27287 (N_27287,N_26705,N_26722);
nor U27288 (N_27288,N_26476,N_26746);
nor U27289 (N_27289,N_26401,N_26744);
and U27290 (N_27290,N_26455,N_26594);
or U27291 (N_27291,N_26912,N_26599);
or U27292 (N_27292,N_26708,N_26644);
or U27293 (N_27293,N_26414,N_26702);
nand U27294 (N_27294,N_26995,N_26767);
nand U27295 (N_27295,N_26756,N_26880);
xnor U27296 (N_27296,N_26890,N_26898);
xor U27297 (N_27297,N_26698,N_26534);
or U27298 (N_27298,N_26763,N_26852);
xor U27299 (N_27299,N_26568,N_26541);
xor U27300 (N_27300,N_26932,N_26907);
nand U27301 (N_27301,N_26754,N_26698);
xor U27302 (N_27302,N_26533,N_26821);
nand U27303 (N_27303,N_26718,N_26604);
and U27304 (N_27304,N_26928,N_26552);
and U27305 (N_27305,N_26460,N_26921);
xor U27306 (N_27306,N_26895,N_26717);
nand U27307 (N_27307,N_26665,N_26400);
xnor U27308 (N_27308,N_26976,N_26522);
or U27309 (N_27309,N_26676,N_26897);
xnor U27310 (N_27310,N_26941,N_26508);
nor U27311 (N_27311,N_26977,N_26516);
nor U27312 (N_27312,N_26875,N_26819);
nand U27313 (N_27313,N_26411,N_26696);
nor U27314 (N_27314,N_26564,N_26880);
or U27315 (N_27315,N_26838,N_26721);
and U27316 (N_27316,N_26620,N_26769);
nor U27317 (N_27317,N_26952,N_26586);
nand U27318 (N_27318,N_26666,N_26870);
and U27319 (N_27319,N_26696,N_26748);
nor U27320 (N_27320,N_26730,N_26658);
and U27321 (N_27321,N_26648,N_26596);
and U27322 (N_27322,N_26801,N_26466);
and U27323 (N_27323,N_26982,N_26730);
nor U27324 (N_27324,N_26708,N_26939);
or U27325 (N_27325,N_26894,N_26435);
nand U27326 (N_27326,N_26802,N_26684);
xor U27327 (N_27327,N_26953,N_26666);
or U27328 (N_27328,N_26768,N_26451);
nand U27329 (N_27329,N_26465,N_26646);
and U27330 (N_27330,N_26967,N_26443);
and U27331 (N_27331,N_26748,N_26708);
nor U27332 (N_27332,N_26914,N_26503);
xor U27333 (N_27333,N_26826,N_26617);
and U27334 (N_27334,N_26565,N_26833);
nand U27335 (N_27335,N_26951,N_26731);
xnor U27336 (N_27336,N_26539,N_26502);
nand U27337 (N_27337,N_26457,N_26854);
xnor U27338 (N_27338,N_26665,N_26990);
xor U27339 (N_27339,N_26755,N_26908);
or U27340 (N_27340,N_26544,N_26554);
and U27341 (N_27341,N_26683,N_26690);
nor U27342 (N_27342,N_26539,N_26948);
or U27343 (N_27343,N_26529,N_26704);
or U27344 (N_27344,N_26582,N_26688);
and U27345 (N_27345,N_26441,N_26892);
and U27346 (N_27346,N_26941,N_26418);
nand U27347 (N_27347,N_26909,N_26938);
and U27348 (N_27348,N_26919,N_26655);
and U27349 (N_27349,N_26416,N_26869);
nor U27350 (N_27350,N_26683,N_26691);
or U27351 (N_27351,N_26545,N_26926);
xor U27352 (N_27352,N_26563,N_26474);
or U27353 (N_27353,N_26873,N_26648);
xnor U27354 (N_27354,N_26986,N_26605);
nor U27355 (N_27355,N_26993,N_26905);
xor U27356 (N_27356,N_26572,N_26811);
nand U27357 (N_27357,N_26571,N_26946);
nor U27358 (N_27358,N_26552,N_26869);
or U27359 (N_27359,N_26640,N_26984);
or U27360 (N_27360,N_26993,N_26585);
nand U27361 (N_27361,N_26560,N_26639);
nand U27362 (N_27362,N_26909,N_26480);
and U27363 (N_27363,N_26463,N_26573);
xnor U27364 (N_27364,N_26854,N_26492);
and U27365 (N_27365,N_26915,N_26549);
nand U27366 (N_27366,N_26606,N_26892);
xnor U27367 (N_27367,N_26652,N_26475);
xnor U27368 (N_27368,N_26523,N_26543);
nor U27369 (N_27369,N_26958,N_26696);
or U27370 (N_27370,N_26844,N_26455);
xnor U27371 (N_27371,N_26646,N_26657);
nand U27372 (N_27372,N_26729,N_26611);
nor U27373 (N_27373,N_26707,N_26500);
and U27374 (N_27374,N_26537,N_26983);
nor U27375 (N_27375,N_26665,N_26830);
xor U27376 (N_27376,N_26971,N_26910);
nand U27377 (N_27377,N_26699,N_26606);
nor U27378 (N_27378,N_26814,N_26616);
or U27379 (N_27379,N_26521,N_26444);
and U27380 (N_27380,N_26504,N_26900);
nand U27381 (N_27381,N_26569,N_26452);
or U27382 (N_27382,N_26729,N_26928);
nand U27383 (N_27383,N_26805,N_26959);
xor U27384 (N_27384,N_26857,N_26533);
xor U27385 (N_27385,N_26985,N_26617);
xnor U27386 (N_27386,N_26684,N_26651);
nand U27387 (N_27387,N_26617,N_26883);
and U27388 (N_27388,N_26918,N_26417);
nand U27389 (N_27389,N_26780,N_26669);
nand U27390 (N_27390,N_26986,N_26478);
or U27391 (N_27391,N_26650,N_26776);
or U27392 (N_27392,N_26837,N_26485);
xnor U27393 (N_27393,N_26959,N_26775);
or U27394 (N_27394,N_26791,N_26874);
or U27395 (N_27395,N_26445,N_26730);
or U27396 (N_27396,N_26518,N_26830);
nor U27397 (N_27397,N_26557,N_26543);
nand U27398 (N_27398,N_26497,N_26714);
nand U27399 (N_27399,N_26812,N_26451);
xnor U27400 (N_27400,N_26725,N_26727);
xor U27401 (N_27401,N_26502,N_26703);
or U27402 (N_27402,N_26627,N_26890);
xor U27403 (N_27403,N_26558,N_26814);
and U27404 (N_27404,N_26767,N_26655);
xor U27405 (N_27405,N_26758,N_26921);
nand U27406 (N_27406,N_26939,N_26454);
nand U27407 (N_27407,N_26745,N_26897);
nor U27408 (N_27408,N_26887,N_26792);
and U27409 (N_27409,N_26854,N_26491);
or U27410 (N_27410,N_26920,N_26935);
nand U27411 (N_27411,N_26716,N_26843);
or U27412 (N_27412,N_26439,N_26777);
and U27413 (N_27413,N_26477,N_26668);
nor U27414 (N_27414,N_26759,N_26610);
xnor U27415 (N_27415,N_26829,N_26401);
xor U27416 (N_27416,N_26496,N_26775);
nand U27417 (N_27417,N_26885,N_26768);
nand U27418 (N_27418,N_26436,N_26564);
or U27419 (N_27419,N_26594,N_26631);
nor U27420 (N_27420,N_26565,N_26797);
or U27421 (N_27421,N_26884,N_26601);
nor U27422 (N_27422,N_26564,N_26924);
nand U27423 (N_27423,N_26888,N_26931);
and U27424 (N_27424,N_26685,N_26636);
xnor U27425 (N_27425,N_26421,N_26787);
and U27426 (N_27426,N_26751,N_26678);
nand U27427 (N_27427,N_26866,N_26635);
nand U27428 (N_27428,N_26564,N_26845);
xnor U27429 (N_27429,N_26427,N_26582);
xor U27430 (N_27430,N_26995,N_26430);
nand U27431 (N_27431,N_26946,N_26878);
or U27432 (N_27432,N_26799,N_26809);
or U27433 (N_27433,N_26648,N_26750);
nor U27434 (N_27434,N_26614,N_26558);
nand U27435 (N_27435,N_26632,N_26654);
xor U27436 (N_27436,N_26457,N_26847);
xor U27437 (N_27437,N_26446,N_26781);
or U27438 (N_27438,N_26828,N_26817);
nor U27439 (N_27439,N_26718,N_26486);
nand U27440 (N_27440,N_26629,N_26878);
and U27441 (N_27441,N_26935,N_26506);
nand U27442 (N_27442,N_26569,N_26541);
nor U27443 (N_27443,N_26435,N_26959);
and U27444 (N_27444,N_26774,N_26440);
nand U27445 (N_27445,N_26963,N_26665);
nand U27446 (N_27446,N_26808,N_26427);
or U27447 (N_27447,N_26953,N_26856);
nor U27448 (N_27448,N_26796,N_26776);
nand U27449 (N_27449,N_26475,N_26623);
nor U27450 (N_27450,N_26517,N_26927);
nand U27451 (N_27451,N_26949,N_26812);
and U27452 (N_27452,N_26945,N_26889);
or U27453 (N_27453,N_26424,N_26600);
and U27454 (N_27454,N_26898,N_26439);
or U27455 (N_27455,N_26858,N_26684);
nand U27456 (N_27456,N_26988,N_26853);
nor U27457 (N_27457,N_26610,N_26837);
nor U27458 (N_27458,N_26545,N_26456);
or U27459 (N_27459,N_26524,N_26670);
nand U27460 (N_27460,N_26831,N_26451);
or U27461 (N_27461,N_26724,N_26447);
nand U27462 (N_27462,N_26783,N_26732);
and U27463 (N_27463,N_26578,N_26715);
xor U27464 (N_27464,N_26959,N_26930);
or U27465 (N_27465,N_26486,N_26760);
nor U27466 (N_27466,N_26599,N_26528);
or U27467 (N_27467,N_26881,N_26732);
nor U27468 (N_27468,N_26552,N_26892);
xor U27469 (N_27469,N_26644,N_26487);
nand U27470 (N_27470,N_26533,N_26656);
nand U27471 (N_27471,N_26663,N_26494);
xor U27472 (N_27472,N_26780,N_26649);
and U27473 (N_27473,N_26927,N_26719);
nand U27474 (N_27474,N_26603,N_26777);
or U27475 (N_27475,N_26905,N_26450);
nor U27476 (N_27476,N_26640,N_26691);
or U27477 (N_27477,N_26743,N_26902);
or U27478 (N_27478,N_26753,N_26756);
and U27479 (N_27479,N_26901,N_26589);
nand U27480 (N_27480,N_26503,N_26539);
nor U27481 (N_27481,N_26865,N_26828);
or U27482 (N_27482,N_26490,N_26881);
nand U27483 (N_27483,N_26419,N_26571);
and U27484 (N_27484,N_26411,N_26717);
nand U27485 (N_27485,N_26533,N_26405);
nand U27486 (N_27486,N_26838,N_26421);
xor U27487 (N_27487,N_26730,N_26944);
xnor U27488 (N_27488,N_26591,N_26474);
xor U27489 (N_27489,N_26789,N_26746);
xor U27490 (N_27490,N_26463,N_26794);
nand U27491 (N_27491,N_26465,N_26403);
nor U27492 (N_27492,N_26965,N_26881);
or U27493 (N_27493,N_26467,N_26654);
xnor U27494 (N_27494,N_26424,N_26595);
nand U27495 (N_27495,N_26597,N_26892);
or U27496 (N_27496,N_26537,N_26749);
nand U27497 (N_27497,N_26750,N_26509);
or U27498 (N_27498,N_26411,N_26700);
xor U27499 (N_27499,N_26536,N_26686);
nand U27500 (N_27500,N_26741,N_26993);
or U27501 (N_27501,N_26803,N_26844);
nor U27502 (N_27502,N_26977,N_26774);
nand U27503 (N_27503,N_26435,N_26810);
nand U27504 (N_27504,N_26778,N_26521);
nor U27505 (N_27505,N_26838,N_26695);
or U27506 (N_27506,N_26866,N_26970);
xnor U27507 (N_27507,N_26754,N_26436);
and U27508 (N_27508,N_26508,N_26926);
or U27509 (N_27509,N_26705,N_26508);
or U27510 (N_27510,N_26993,N_26962);
xor U27511 (N_27511,N_26914,N_26622);
nor U27512 (N_27512,N_26785,N_26534);
or U27513 (N_27513,N_26816,N_26635);
nor U27514 (N_27514,N_26648,N_26604);
or U27515 (N_27515,N_26851,N_26940);
nor U27516 (N_27516,N_26502,N_26441);
or U27517 (N_27517,N_26937,N_26551);
nand U27518 (N_27518,N_26411,N_26458);
or U27519 (N_27519,N_26918,N_26644);
or U27520 (N_27520,N_26761,N_26587);
nor U27521 (N_27521,N_26434,N_26751);
nand U27522 (N_27522,N_26603,N_26728);
nand U27523 (N_27523,N_26763,N_26818);
and U27524 (N_27524,N_26520,N_26403);
and U27525 (N_27525,N_26631,N_26865);
xor U27526 (N_27526,N_26691,N_26401);
and U27527 (N_27527,N_26651,N_26901);
nand U27528 (N_27528,N_26973,N_26471);
nor U27529 (N_27529,N_26730,N_26964);
nand U27530 (N_27530,N_26978,N_26614);
nor U27531 (N_27531,N_26613,N_26708);
and U27532 (N_27532,N_26467,N_26475);
nor U27533 (N_27533,N_26608,N_26430);
xor U27534 (N_27534,N_26619,N_26491);
nand U27535 (N_27535,N_26761,N_26878);
and U27536 (N_27536,N_26731,N_26662);
and U27537 (N_27537,N_26842,N_26589);
nand U27538 (N_27538,N_26670,N_26445);
or U27539 (N_27539,N_26513,N_26956);
nand U27540 (N_27540,N_26957,N_26523);
nor U27541 (N_27541,N_26993,N_26735);
xor U27542 (N_27542,N_26703,N_26538);
or U27543 (N_27543,N_26984,N_26951);
nor U27544 (N_27544,N_26786,N_26780);
xor U27545 (N_27545,N_26437,N_26721);
xnor U27546 (N_27546,N_26566,N_26446);
or U27547 (N_27547,N_26606,N_26834);
xnor U27548 (N_27548,N_26994,N_26883);
or U27549 (N_27549,N_26527,N_26560);
and U27550 (N_27550,N_26475,N_26827);
nor U27551 (N_27551,N_26596,N_26443);
nor U27552 (N_27552,N_26730,N_26599);
or U27553 (N_27553,N_26567,N_26719);
nand U27554 (N_27554,N_26923,N_26468);
xor U27555 (N_27555,N_26499,N_26436);
and U27556 (N_27556,N_26917,N_26453);
and U27557 (N_27557,N_26663,N_26487);
nor U27558 (N_27558,N_26900,N_26602);
and U27559 (N_27559,N_26553,N_26496);
nor U27560 (N_27560,N_26491,N_26984);
or U27561 (N_27561,N_26800,N_26531);
xnor U27562 (N_27562,N_26815,N_26781);
nand U27563 (N_27563,N_26862,N_26505);
xor U27564 (N_27564,N_26555,N_26462);
xor U27565 (N_27565,N_26880,N_26595);
nand U27566 (N_27566,N_26531,N_26496);
xnor U27567 (N_27567,N_26660,N_26533);
or U27568 (N_27568,N_26525,N_26473);
or U27569 (N_27569,N_26514,N_26590);
or U27570 (N_27570,N_26931,N_26612);
nand U27571 (N_27571,N_26981,N_26620);
or U27572 (N_27572,N_26875,N_26557);
nand U27573 (N_27573,N_26746,N_26598);
nand U27574 (N_27574,N_26693,N_26639);
xor U27575 (N_27575,N_26758,N_26715);
nand U27576 (N_27576,N_26542,N_26776);
nor U27577 (N_27577,N_26974,N_26569);
or U27578 (N_27578,N_26803,N_26966);
xor U27579 (N_27579,N_26923,N_26874);
or U27580 (N_27580,N_26796,N_26901);
nand U27581 (N_27581,N_26649,N_26442);
xnor U27582 (N_27582,N_26987,N_26404);
nand U27583 (N_27583,N_26935,N_26805);
xor U27584 (N_27584,N_26808,N_26749);
and U27585 (N_27585,N_26928,N_26786);
and U27586 (N_27586,N_26817,N_26995);
nand U27587 (N_27587,N_26854,N_26556);
xor U27588 (N_27588,N_26819,N_26611);
and U27589 (N_27589,N_26715,N_26680);
and U27590 (N_27590,N_26975,N_26716);
nand U27591 (N_27591,N_26578,N_26720);
or U27592 (N_27592,N_26798,N_26639);
xor U27593 (N_27593,N_26537,N_26621);
or U27594 (N_27594,N_26846,N_26512);
nand U27595 (N_27595,N_26631,N_26701);
and U27596 (N_27596,N_26405,N_26625);
and U27597 (N_27597,N_26606,N_26443);
nand U27598 (N_27598,N_26468,N_26936);
and U27599 (N_27599,N_26844,N_26533);
xnor U27600 (N_27600,N_27032,N_27114);
and U27601 (N_27601,N_27170,N_27250);
xor U27602 (N_27602,N_27290,N_27314);
or U27603 (N_27603,N_27262,N_27404);
nor U27604 (N_27604,N_27111,N_27279);
or U27605 (N_27605,N_27365,N_27096);
and U27606 (N_27606,N_27068,N_27287);
or U27607 (N_27607,N_27004,N_27196);
nor U27608 (N_27608,N_27014,N_27309);
nand U27609 (N_27609,N_27077,N_27083);
or U27610 (N_27610,N_27289,N_27478);
and U27611 (N_27611,N_27393,N_27218);
nand U27612 (N_27612,N_27100,N_27126);
xor U27613 (N_27613,N_27230,N_27491);
or U27614 (N_27614,N_27240,N_27121);
nand U27615 (N_27615,N_27277,N_27324);
and U27616 (N_27616,N_27310,N_27165);
nor U27617 (N_27617,N_27430,N_27294);
nand U27618 (N_27618,N_27179,N_27398);
nand U27619 (N_27619,N_27358,N_27442);
or U27620 (N_27620,N_27207,N_27137);
or U27621 (N_27621,N_27496,N_27595);
or U27622 (N_27622,N_27475,N_27204);
nor U27623 (N_27623,N_27097,N_27331);
nand U27624 (N_27624,N_27092,N_27584);
nor U27625 (N_27625,N_27446,N_27009);
nor U27626 (N_27626,N_27284,N_27282);
and U27627 (N_27627,N_27188,N_27167);
and U27628 (N_27628,N_27265,N_27192);
or U27629 (N_27629,N_27316,N_27039);
or U27630 (N_27630,N_27185,N_27254);
nor U27631 (N_27631,N_27276,N_27258);
or U27632 (N_27632,N_27460,N_27055);
or U27633 (N_27633,N_27356,N_27351);
nand U27634 (N_27634,N_27163,N_27295);
and U27635 (N_27635,N_27427,N_27132);
nand U27636 (N_27636,N_27221,N_27182);
nor U27637 (N_27637,N_27539,N_27286);
or U27638 (N_27638,N_27283,N_27368);
or U27639 (N_27639,N_27171,N_27473);
and U27640 (N_27640,N_27134,N_27555);
xor U27641 (N_27641,N_27005,N_27317);
and U27642 (N_27642,N_27047,N_27244);
and U27643 (N_27643,N_27523,N_27572);
or U27644 (N_27644,N_27166,N_27236);
xnor U27645 (N_27645,N_27469,N_27548);
and U27646 (N_27646,N_27220,N_27502);
or U27647 (N_27647,N_27383,N_27044);
xor U27648 (N_27648,N_27151,N_27482);
nand U27649 (N_27649,N_27110,N_27519);
xnor U27650 (N_27650,N_27078,N_27147);
or U27651 (N_27651,N_27041,N_27328);
nor U27652 (N_27652,N_27193,N_27264);
nand U27653 (N_27653,N_27545,N_27015);
nor U27654 (N_27654,N_27088,N_27000);
and U27655 (N_27655,N_27191,N_27468);
nand U27656 (N_27656,N_27497,N_27259);
xor U27657 (N_27657,N_27367,N_27085);
nand U27658 (N_27658,N_27586,N_27072);
and U27659 (N_27659,N_27190,N_27387);
nand U27660 (N_27660,N_27094,N_27023);
and U27661 (N_27661,N_27483,N_27037);
and U27662 (N_27662,N_27210,N_27579);
xnor U27663 (N_27663,N_27474,N_27175);
xor U27664 (N_27664,N_27566,N_27411);
and U27665 (N_27665,N_27285,N_27256);
or U27666 (N_27666,N_27599,N_27026);
xnor U27667 (N_27667,N_27061,N_27139);
and U27668 (N_27668,N_27433,N_27526);
and U27669 (N_27669,N_27381,N_27101);
nand U27670 (N_27670,N_27223,N_27150);
xnor U27671 (N_27671,N_27124,N_27071);
nor U27672 (N_27672,N_27326,N_27148);
nand U27673 (N_27673,N_27457,N_27048);
nand U27674 (N_27674,N_27544,N_27470);
nand U27675 (N_27675,N_27552,N_27081);
and U27676 (N_27676,N_27325,N_27213);
and U27677 (N_27677,N_27117,N_27030);
and U27678 (N_27678,N_27522,N_27127);
or U27679 (N_27679,N_27378,N_27530);
nand U27680 (N_27680,N_27487,N_27480);
xnor U27681 (N_27681,N_27027,N_27202);
nor U27682 (N_27682,N_27180,N_27518);
nand U27683 (N_27683,N_27389,N_27375);
nand U27684 (N_27684,N_27371,N_27436);
or U27685 (N_27685,N_27059,N_27532);
xnor U27686 (N_27686,N_27456,N_27403);
or U27687 (N_27687,N_27575,N_27510);
nand U27688 (N_27688,N_27341,N_27141);
nand U27689 (N_27689,N_27238,N_27099);
xor U27690 (N_27690,N_27146,N_27297);
nor U27691 (N_27691,N_27489,N_27020);
or U27692 (N_27692,N_27205,N_27402);
nand U27693 (N_27693,N_27329,N_27057);
xor U27694 (N_27694,N_27400,N_27012);
nand U27695 (N_27695,N_27394,N_27098);
and U27696 (N_27696,N_27525,N_27506);
or U27697 (N_27697,N_27063,N_27155);
and U27698 (N_27698,N_27422,N_27299);
xor U27699 (N_27699,N_27149,N_27407);
and U27700 (N_27700,N_27248,N_27231);
xor U27701 (N_27701,N_27273,N_27354);
or U27702 (N_27702,N_27449,N_27472);
nor U27703 (N_27703,N_27247,N_27076);
nand U27704 (N_27704,N_27567,N_27206);
and U27705 (N_27705,N_27554,N_27194);
and U27706 (N_27706,N_27217,N_27355);
or U27707 (N_27707,N_27122,N_27500);
nor U27708 (N_27708,N_27542,N_27578);
and U27709 (N_27709,N_27533,N_27538);
nand U27710 (N_27710,N_27024,N_27168);
nand U27711 (N_27711,N_27476,N_27018);
nor U27712 (N_27712,N_27156,N_27342);
or U27713 (N_27713,N_27275,N_27327);
nor U27714 (N_27714,N_27219,N_27298);
xnor U27715 (N_27715,N_27235,N_27036);
and U27716 (N_27716,N_27103,N_27452);
or U27717 (N_27717,N_27490,N_27471);
or U27718 (N_27718,N_27498,N_27379);
xor U27719 (N_27719,N_27089,N_27215);
xor U27720 (N_27720,N_27271,N_27073);
xnor U27721 (N_27721,N_27019,N_27527);
nand U27722 (N_27722,N_27348,N_27549);
nor U27723 (N_27723,N_27591,N_27302);
or U27724 (N_27724,N_27531,N_27455);
and U27725 (N_27725,N_27153,N_27115);
nor U27726 (N_27726,N_27107,N_27561);
or U27727 (N_27727,N_27105,N_27189);
nor U27728 (N_27728,N_27070,N_27435);
and U27729 (N_27729,N_27082,N_27292);
xor U27730 (N_27730,N_27125,N_27176);
nand U27731 (N_27731,N_27187,N_27138);
or U27732 (N_27732,N_27420,N_27161);
and U27733 (N_27733,N_27415,N_27528);
xor U27734 (N_27734,N_27512,N_27479);
nor U27735 (N_27735,N_27459,N_27577);
and U27736 (N_27736,N_27425,N_27065);
nor U27737 (N_27737,N_27514,N_27142);
xnor U27738 (N_27738,N_27080,N_27501);
and U27739 (N_27739,N_27597,N_27405);
nand U27740 (N_27740,N_27598,N_27164);
and U27741 (N_27741,N_27260,N_27521);
nor U27742 (N_27742,N_27056,N_27390);
nand U27743 (N_27743,N_27136,N_27488);
and U27744 (N_27744,N_27051,N_27344);
and U27745 (N_27745,N_27408,N_27253);
nand U27746 (N_27746,N_27364,N_27492);
nor U27747 (N_27747,N_27308,N_27395);
and U27748 (N_27748,N_27226,N_27133);
or U27749 (N_27749,N_27128,N_27347);
xor U27750 (N_27750,N_27551,N_27440);
or U27751 (N_27751,N_27064,N_27054);
nor U27752 (N_27752,N_27546,N_27323);
or U27753 (N_27753,N_27090,N_27537);
xnor U27754 (N_27754,N_27143,N_27162);
xnor U27755 (N_27755,N_27046,N_27432);
and U27756 (N_27756,N_27493,N_27588);
xor U27757 (N_27757,N_27335,N_27031);
or U27758 (N_27758,N_27516,N_27252);
xnor U27759 (N_27759,N_27560,N_27507);
and U27760 (N_27760,N_27450,N_27222);
nor U27761 (N_27761,N_27203,N_27332);
nor U27762 (N_27762,N_27319,N_27573);
and U27763 (N_27763,N_27372,N_27304);
xor U27764 (N_27764,N_27352,N_27465);
or U27765 (N_27765,N_27382,N_27257);
nor U27766 (N_27766,N_27087,N_27246);
nand U27767 (N_27767,N_27233,N_27200);
xor U27768 (N_27768,N_27003,N_27412);
and U27769 (N_27769,N_27343,N_27401);
and U27770 (N_27770,N_27001,N_27119);
nand U27771 (N_27771,N_27086,N_27447);
or U27772 (N_27772,N_27249,N_27157);
or U27773 (N_27773,N_27118,N_27458);
nand U27774 (N_27774,N_27587,N_27216);
and U27775 (N_27775,N_27414,N_27330);
and U27776 (N_27776,N_27373,N_27034);
xnor U27777 (N_27777,N_27035,N_27583);
and U27778 (N_27778,N_27195,N_27423);
nor U27779 (N_27779,N_27592,N_27208);
or U27780 (N_27780,N_27008,N_27568);
nor U27781 (N_27781,N_27232,N_27384);
or U27782 (N_27782,N_27464,N_27120);
xnor U27783 (N_27783,N_27535,N_27011);
nor U27784 (N_27784,N_27198,N_27154);
nand U27785 (N_27785,N_27439,N_27060);
nor U27786 (N_27786,N_27333,N_27511);
nand U27787 (N_27787,N_27558,N_27376);
xor U27788 (N_27788,N_27495,N_27543);
xnor U27789 (N_27789,N_27123,N_27234);
nand U27790 (N_27790,N_27569,N_27564);
xnor U27791 (N_27791,N_27069,N_27209);
nor U27792 (N_27792,N_27385,N_27485);
nor U27793 (N_27793,N_27438,N_27013);
xnor U27794 (N_27794,N_27370,N_27291);
nand U27795 (N_27795,N_27444,N_27504);
xnor U27796 (N_27796,N_27010,N_27093);
or U27797 (N_27797,N_27074,N_27261);
or U27798 (N_27798,N_27278,N_27296);
nand U27799 (N_27799,N_27269,N_27050);
nand U27800 (N_27800,N_27006,N_27428);
nor U27801 (N_27801,N_27448,N_27116);
nand U27802 (N_27802,N_27225,N_27300);
nand U27803 (N_27803,N_27270,N_27321);
and U27804 (N_27804,N_27245,N_27353);
and U27805 (N_27805,N_27361,N_27241);
xnor U27806 (N_27806,N_27349,N_27534);
and U27807 (N_27807,N_27434,N_27517);
xor U27808 (N_27808,N_27437,N_27315);
or U27809 (N_27809,N_27075,N_27547);
nand U27810 (N_27810,N_27380,N_27084);
and U27811 (N_27811,N_27145,N_27007);
and U27812 (N_27812,N_27536,N_27158);
nor U27813 (N_27813,N_27513,N_27021);
nor U27814 (N_27814,N_27529,N_27392);
nand U27815 (N_27815,N_27274,N_27388);
nand U27816 (N_27816,N_27453,N_27183);
and U27817 (N_27817,N_27441,N_27002);
nand U27818 (N_27818,N_27419,N_27267);
and U27819 (N_27819,N_27224,N_27463);
nand U27820 (N_27820,N_27102,N_27307);
nand U27821 (N_27821,N_27280,N_27106);
nand U27822 (N_27822,N_27045,N_27494);
nor U27823 (N_27823,N_27152,N_27160);
and U27824 (N_27824,N_27509,N_27505);
and U27825 (N_27825,N_27229,N_27243);
nor U27826 (N_27826,N_27172,N_27550);
xor U27827 (N_27827,N_27112,N_27184);
or U27828 (N_27828,N_27268,N_27186);
nor U27829 (N_27829,N_27058,N_27357);
and U27830 (N_27830,N_27445,N_27091);
xor U27831 (N_27831,N_27016,N_27462);
and U27832 (N_27832,N_27318,N_27320);
nor U27833 (N_27833,N_27066,N_27052);
xnor U27834 (N_27834,N_27574,N_27255);
and U27835 (N_27835,N_27337,N_27466);
or U27836 (N_27836,N_27350,N_27360);
and U27837 (N_27837,N_27589,N_27239);
nand U27838 (N_27838,N_27557,N_27374);
nand U27839 (N_27839,N_27177,N_27028);
and U27840 (N_27840,N_27563,N_27042);
xnor U27841 (N_27841,N_27340,N_27429);
or U27842 (N_27842,N_27593,N_27359);
nand U27843 (N_27843,N_27140,N_27369);
nor U27844 (N_27844,N_27301,N_27406);
and U27845 (N_27845,N_27334,N_27212);
nor U27846 (N_27846,N_27396,N_27391);
nand U27847 (N_27847,N_27040,N_27556);
or U27848 (N_27848,N_27339,N_27017);
or U27849 (N_27849,N_27594,N_27251);
xor U27850 (N_27850,N_27311,N_27053);
or U27851 (N_27851,N_27113,N_27362);
xnor U27852 (N_27852,N_27033,N_27197);
and U27853 (N_27853,N_27467,N_27443);
nand U27854 (N_27854,N_27227,N_27590);
nor U27855 (N_27855,N_27173,N_27174);
nor U27856 (N_27856,N_27303,N_27477);
and U27857 (N_27857,N_27363,N_27263);
or U27858 (N_27858,N_27410,N_27043);
xnor U27859 (N_27859,N_27022,N_27520);
nand U27860 (N_27860,N_27237,N_27062);
xor U27861 (N_27861,N_27426,N_27305);
nand U27862 (N_27862,N_27580,N_27159);
xor U27863 (N_27863,N_27386,N_27499);
and U27864 (N_27864,N_27366,N_27129);
or U27865 (N_27865,N_27508,N_27038);
and U27866 (N_27866,N_27481,N_27541);
or U27867 (N_27867,N_27416,N_27029);
nand U27868 (N_27868,N_27562,N_27109);
and U27869 (N_27869,N_27228,N_27293);
and U27870 (N_27870,N_27211,N_27135);
nand U27871 (N_27871,N_27553,N_27418);
xnor U27872 (N_27872,N_27559,N_27025);
xnor U27873 (N_27873,N_27486,N_27272);
or U27874 (N_27874,N_27131,N_27581);
nor U27875 (N_27875,N_27346,N_27306);
and U27876 (N_27876,N_27322,N_27095);
and U27877 (N_27877,N_27571,N_27409);
nor U27878 (N_27878,N_27130,N_27144);
and U27879 (N_27879,N_27281,N_27336);
nand U27880 (N_27880,N_27417,N_27178);
or U27881 (N_27881,N_27079,N_27451);
nand U27882 (N_27882,N_27565,N_27461);
and U27883 (N_27883,N_27582,N_27596);
or U27884 (N_27884,N_27524,N_27431);
xnor U27885 (N_27885,N_27345,N_27312);
or U27886 (N_27886,N_27338,N_27454);
or U27887 (N_27887,N_27515,N_27169);
nor U27888 (N_27888,N_27288,N_27540);
xnor U27889 (N_27889,N_27067,N_27585);
xor U27890 (N_27890,N_27503,N_27377);
and U27891 (N_27891,N_27199,N_27397);
nor U27892 (N_27892,N_27421,N_27484);
nor U27893 (N_27893,N_27399,N_27214);
nor U27894 (N_27894,N_27266,N_27313);
nor U27895 (N_27895,N_27242,N_27104);
or U27896 (N_27896,N_27424,N_27570);
nor U27897 (N_27897,N_27413,N_27201);
or U27898 (N_27898,N_27108,N_27181);
nand U27899 (N_27899,N_27576,N_27049);
or U27900 (N_27900,N_27076,N_27504);
and U27901 (N_27901,N_27036,N_27503);
xnor U27902 (N_27902,N_27122,N_27378);
and U27903 (N_27903,N_27296,N_27514);
nand U27904 (N_27904,N_27256,N_27191);
xor U27905 (N_27905,N_27477,N_27208);
nor U27906 (N_27906,N_27182,N_27186);
nand U27907 (N_27907,N_27068,N_27501);
or U27908 (N_27908,N_27230,N_27463);
nand U27909 (N_27909,N_27212,N_27526);
or U27910 (N_27910,N_27014,N_27560);
xor U27911 (N_27911,N_27300,N_27064);
xnor U27912 (N_27912,N_27152,N_27097);
or U27913 (N_27913,N_27564,N_27068);
or U27914 (N_27914,N_27248,N_27491);
nor U27915 (N_27915,N_27598,N_27575);
or U27916 (N_27916,N_27579,N_27272);
xnor U27917 (N_27917,N_27453,N_27347);
or U27918 (N_27918,N_27479,N_27013);
and U27919 (N_27919,N_27205,N_27283);
nor U27920 (N_27920,N_27448,N_27335);
nand U27921 (N_27921,N_27323,N_27191);
nand U27922 (N_27922,N_27037,N_27049);
nor U27923 (N_27923,N_27229,N_27525);
and U27924 (N_27924,N_27194,N_27501);
or U27925 (N_27925,N_27396,N_27338);
nor U27926 (N_27926,N_27286,N_27592);
or U27927 (N_27927,N_27494,N_27222);
nor U27928 (N_27928,N_27237,N_27165);
and U27929 (N_27929,N_27005,N_27560);
nand U27930 (N_27930,N_27556,N_27432);
xor U27931 (N_27931,N_27462,N_27390);
xnor U27932 (N_27932,N_27324,N_27535);
xnor U27933 (N_27933,N_27328,N_27272);
xnor U27934 (N_27934,N_27331,N_27094);
or U27935 (N_27935,N_27575,N_27231);
nor U27936 (N_27936,N_27539,N_27567);
or U27937 (N_27937,N_27495,N_27417);
and U27938 (N_27938,N_27524,N_27214);
or U27939 (N_27939,N_27320,N_27442);
xnor U27940 (N_27940,N_27288,N_27257);
or U27941 (N_27941,N_27115,N_27034);
or U27942 (N_27942,N_27239,N_27203);
and U27943 (N_27943,N_27241,N_27078);
and U27944 (N_27944,N_27435,N_27024);
nor U27945 (N_27945,N_27150,N_27231);
nand U27946 (N_27946,N_27210,N_27190);
or U27947 (N_27947,N_27216,N_27000);
nor U27948 (N_27948,N_27473,N_27338);
nand U27949 (N_27949,N_27314,N_27007);
nand U27950 (N_27950,N_27336,N_27409);
and U27951 (N_27951,N_27071,N_27023);
xnor U27952 (N_27952,N_27485,N_27156);
xor U27953 (N_27953,N_27224,N_27110);
xnor U27954 (N_27954,N_27448,N_27443);
and U27955 (N_27955,N_27412,N_27076);
or U27956 (N_27956,N_27003,N_27428);
nor U27957 (N_27957,N_27449,N_27029);
nor U27958 (N_27958,N_27308,N_27130);
nand U27959 (N_27959,N_27071,N_27057);
or U27960 (N_27960,N_27221,N_27522);
xnor U27961 (N_27961,N_27455,N_27026);
or U27962 (N_27962,N_27506,N_27057);
nand U27963 (N_27963,N_27288,N_27318);
nand U27964 (N_27964,N_27235,N_27160);
nor U27965 (N_27965,N_27000,N_27473);
or U27966 (N_27966,N_27106,N_27474);
xor U27967 (N_27967,N_27198,N_27543);
nor U27968 (N_27968,N_27363,N_27198);
nor U27969 (N_27969,N_27088,N_27080);
and U27970 (N_27970,N_27271,N_27330);
nor U27971 (N_27971,N_27449,N_27414);
xnor U27972 (N_27972,N_27420,N_27030);
nor U27973 (N_27973,N_27465,N_27448);
and U27974 (N_27974,N_27007,N_27294);
or U27975 (N_27975,N_27496,N_27038);
nand U27976 (N_27976,N_27487,N_27224);
nor U27977 (N_27977,N_27549,N_27361);
nor U27978 (N_27978,N_27348,N_27439);
nor U27979 (N_27979,N_27500,N_27440);
or U27980 (N_27980,N_27077,N_27390);
nor U27981 (N_27981,N_27141,N_27444);
xor U27982 (N_27982,N_27133,N_27190);
nand U27983 (N_27983,N_27384,N_27317);
xor U27984 (N_27984,N_27447,N_27146);
xnor U27985 (N_27985,N_27142,N_27194);
xor U27986 (N_27986,N_27392,N_27108);
and U27987 (N_27987,N_27574,N_27474);
nand U27988 (N_27988,N_27248,N_27107);
xnor U27989 (N_27989,N_27019,N_27529);
and U27990 (N_27990,N_27147,N_27575);
nor U27991 (N_27991,N_27208,N_27111);
xor U27992 (N_27992,N_27062,N_27422);
nor U27993 (N_27993,N_27519,N_27227);
xor U27994 (N_27994,N_27190,N_27584);
nand U27995 (N_27995,N_27046,N_27040);
xnor U27996 (N_27996,N_27061,N_27346);
or U27997 (N_27997,N_27458,N_27328);
nor U27998 (N_27998,N_27561,N_27082);
or U27999 (N_27999,N_27503,N_27332);
nand U28000 (N_28000,N_27015,N_27580);
or U28001 (N_28001,N_27022,N_27309);
or U28002 (N_28002,N_27047,N_27501);
or U28003 (N_28003,N_27181,N_27543);
xor U28004 (N_28004,N_27246,N_27478);
xnor U28005 (N_28005,N_27095,N_27266);
and U28006 (N_28006,N_27502,N_27459);
xor U28007 (N_28007,N_27232,N_27477);
and U28008 (N_28008,N_27383,N_27167);
or U28009 (N_28009,N_27347,N_27016);
nand U28010 (N_28010,N_27448,N_27231);
or U28011 (N_28011,N_27377,N_27066);
xor U28012 (N_28012,N_27145,N_27511);
nor U28013 (N_28013,N_27311,N_27548);
or U28014 (N_28014,N_27052,N_27524);
or U28015 (N_28015,N_27517,N_27338);
or U28016 (N_28016,N_27016,N_27582);
nand U28017 (N_28017,N_27559,N_27377);
and U28018 (N_28018,N_27401,N_27109);
nor U28019 (N_28019,N_27304,N_27477);
xnor U28020 (N_28020,N_27589,N_27356);
and U28021 (N_28021,N_27199,N_27230);
nand U28022 (N_28022,N_27244,N_27483);
or U28023 (N_28023,N_27566,N_27095);
nand U28024 (N_28024,N_27597,N_27286);
nand U28025 (N_28025,N_27123,N_27125);
nor U28026 (N_28026,N_27435,N_27369);
nand U28027 (N_28027,N_27589,N_27514);
nand U28028 (N_28028,N_27498,N_27133);
nand U28029 (N_28029,N_27444,N_27016);
nand U28030 (N_28030,N_27416,N_27114);
xnor U28031 (N_28031,N_27302,N_27464);
nand U28032 (N_28032,N_27073,N_27395);
nor U28033 (N_28033,N_27094,N_27095);
nor U28034 (N_28034,N_27473,N_27523);
nand U28035 (N_28035,N_27445,N_27018);
nor U28036 (N_28036,N_27565,N_27431);
nand U28037 (N_28037,N_27462,N_27467);
xor U28038 (N_28038,N_27564,N_27200);
nand U28039 (N_28039,N_27455,N_27512);
xnor U28040 (N_28040,N_27403,N_27330);
nand U28041 (N_28041,N_27425,N_27151);
or U28042 (N_28042,N_27129,N_27101);
and U28043 (N_28043,N_27393,N_27366);
and U28044 (N_28044,N_27034,N_27529);
nand U28045 (N_28045,N_27139,N_27447);
nand U28046 (N_28046,N_27502,N_27450);
and U28047 (N_28047,N_27106,N_27490);
xnor U28048 (N_28048,N_27349,N_27055);
nand U28049 (N_28049,N_27177,N_27446);
nor U28050 (N_28050,N_27311,N_27458);
nand U28051 (N_28051,N_27250,N_27511);
nor U28052 (N_28052,N_27210,N_27192);
nand U28053 (N_28053,N_27310,N_27088);
and U28054 (N_28054,N_27056,N_27575);
or U28055 (N_28055,N_27140,N_27078);
xnor U28056 (N_28056,N_27064,N_27584);
or U28057 (N_28057,N_27479,N_27007);
or U28058 (N_28058,N_27177,N_27245);
nor U28059 (N_28059,N_27248,N_27261);
or U28060 (N_28060,N_27130,N_27336);
or U28061 (N_28061,N_27294,N_27035);
and U28062 (N_28062,N_27117,N_27177);
nor U28063 (N_28063,N_27405,N_27070);
nor U28064 (N_28064,N_27026,N_27001);
xor U28065 (N_28065,N_27001,N_27090);
or U28066 (N_28066,N_27422,N_27416);
nand U28067 (N_28067,N_27530,N_27343);
nor U28068 (N_28068,N_27047,N_27450);
nor U28069 (N_28069,N_27481,N_27023);
xor U28070 (N_28070,N_27473,N_27035);
nand U28071 (N_28071,N_27149,N_27460);
nor U28072 (N_28072,N_27025,N_27380);
xor U28073 (N_28073,N_27423,N_27339);
or U28074 (N_28074,N_27452,N_27217);
xor U28075 (N_28075,N_27446,N_27219);
or U28076 (N_28076,N_27116,N_27109);
xnor U28077 (N_28077,N_27203,N_27088);
nand U28078 (N_28078,N_27409,N_27518);
nor U28079 (N_28079,N_27575,N_27296);
nor U28080 (N_28080,N_27047,N_27522);
and U28081 (N_28081,N_27151,N_27437);
and U28082 (N_28082,N_27425,N_27328);
and U28083 (N_28083,N_27026,N_27301);
xor U28084 (N_28084,N_27198,N_27202);
nor U28085 (N_28085,N_27189,N_27520);
xor U28086 (N_28086,N_27306,N_27064);
xor U28087 (N_28087,N_27208,N_27533);
and U28088 (N_28088,N_27598,N_27027);
and U28089 (N_28089,N_27531,N_27033);
or U28090 (N_28090,N_27214,N_27379);
xnor U28091 (N_28091,N_27504,N_27404);
xnor U28092 (N_28092,N_27058,N_27511);
nand U28093 (N_28093,N_27313,N_27529);
xnor U28094 (N_28094,N_27484,N_27475);
or U28095 (N_28095,N_27248,N_27402);
nand U28096 (N_28096,N_27129,N_27396);
nor U28097 (N_28097,N_27064,N_27404);
and U28098 (N_28098,N_27015,N_27389);
and U28099 (N_28099,N_27503,N_27228);
or U28100 (N_28100,N_27211,N_27345);
nand U28101 (N_28101,N_27059,N_27099);
or U28102 (N_28102,N_27522,N_27158);
nand U28103 (N_28103,N_27420,N_27339);
nand U28104 (N_28104,N_27343,N_27539);
xor U28105 (N_28105,N_27529,N_27179);
or U28106 (N_28106,N_27213,N_27492);
or U28107 (N_28107,N_27441,N_27551);
and U28108 (N_28108,N_27063,N_27519);
or U28109 (N_28109,N_27582,N_27223);
and U28110 (N_28110,N_27375,N_27502);
nor U28111 (N_28111,N_27000,N_27053);
nor U28112 (N_28112,N_27381,N_27013);
and U28113 (N_28113,N_27424,N_27262);
xnor U28114 (N_28114,N_27467,N_27324);
xor U28115 (N_28115,N_27485,N_27136);
or U28116 (N_28116,N_27141,N_27307);
nand U28117 (N_28117,N_27216,N_27434);
xor U28118 (N_28118,N_27483,N_27589);
and U28119 (N_28119,N_27095,N_27458);
nor U28120 (N_28120,N_27356,N_27577);
nand U28121 (N_28121,N_27133,N_27225);
xor U28122 (N_28122,N_27214,N_27453);
xnor U28123 (N_28123,N_27322,N_27297);
xor U28124 (N_28124,N_27499,N_27180);
or U28125 (N_28125,N_27269,N_27037);
nand U28126 (N_28126,N_27355,N_27452);
nor U28127 (N_28127,N_27588,N_27249);
and U28128 (N_28128,N_27260,N_27302);
nand U28129 (N_28129,N_27368,N_27575);
and U28130 (N_28130,N_27187,N_27533);
or U28131 (N_28131,N_27188,N_27332);
nor U28132 (N_28132,N_27263,N_27279);
nor U28133 (N_28133,N_27314,N_27031);
and U28134 (N_28134,N_27551,N_27517);
nor U28135 (N_28135,N_27023,N_27461);
xor U28136 (N_28136,N_27381,N_27014);
nand U28137 (N_28137,N_27361,N_27511);
nor U28138 (N_28138,N_27016,N_27391);
or U28139 (N_28139,N_27334,N_27058);
nand U28140 (N_28140,N_27479,N_27218);
nand U28141 (N_28141,N_27252,N_27118);
nand U28142 (N_28142,N_27012,N_27468);
nor U28143 (N_28143,N_27399,N_27354);
xor U28144 (N_28144,N_27021,N_27189);
nand U28145 (N_28145,N_27298,N_27209);
and U28146 (N_28146,N_27039,N_27187);
xor U28147 (N_28147,N_27060,N_27264);
or U28148 (N_28148,N_27316,N_27537);
or U28149 (N_28149,N_27353,N_27006);
or U28150 (N_28150,N_27127,N_27565);
xor U28151 (N_28151,N_27410,N_27535);
or U28152 (N_28152,N_27133,N_27284);
nand U28153 (N_28153,N_27146,N_27008);
or U28154 (N_28154,N_27506,N_27337);
nand U28155 (N_28155,N_27171,N_27085);
or U28156 (N_28156,N_27511,N_27388);
xnor U28157 (N_28157,N_27494,N_27411);
nand U28158 (N_28158,N_27240,N_27034);
or U28159 (N_28159,N_27473,N_27405);
or U28160 (N_28160,N_27290,N_27530);
and U28161 (N_28161,N_27373,N_27508);
nand U28162 (N_28162,N_27097,N_27308);
and U28163 (N_28163,N_27496,N_27015);
and U28164 (N_28164,N_27398,N_27185);
xor U28165 (N_28165,N_27423,N_27479);
nor U28166 (N_28166,N_27155,N_27175);
xnor U28167 (N_28167,N_27511,N_27135);
or U28168 (N_28168,N_27479,N_27055);
nor U28169 (N_28169,N_27384,N_27010);
nand U28170 (N_28170,N_27356,N_27075);
and U28171 (N_28171,N_27298,N_27030);
and U28172 (N_28172,N_27205,N_27539);
and U28173 (N_28173,N_27553,N_27258);
nor U28174 (N_28174,N_27042,N_27031);
nor U28175 (N_28175,N_27274,N_27519);
or U28176 (N_28176,N_27387,N_27092);
or U28177 (N_28177,N_27064,N_27235);
and U28178 (N_28178,N_27426,N_27221);
nand U28179 (N_28179,N_27217,N_27376);
nand U28180 (N_28180,N_27157,N_27535);
nor U28181 (N_28181,N_27381,N_27008);
or U28182 (N_28182,N_27494,N_27543);
xnor U28183 (N_28183,N_27093,N_27300);
and U28184 (N_28184,N_27438,N_27598);
and U28185 (N_28185,N_27154,N_27356);
xor U28186 (N_28186,N_27408,N_27068);
and U28187 (N_28187,N_27374,N_27467);
and U28188 (N_28188,N_27540,N_27476);
xor U28189 (N_28189,N_27471,N_27408);
or U28190 (N_28190,N_27501,N_27234);
nor U28191 (N_28191,N_27370,N_27209);
nand U28192 (N_28192,N_27020,N_27463);
xnor U28193 (N_28193,N_27301,N_27194);
nor U28194 (N_28194,N_27463,N_27514);
nand U28195 (N_28195,N_27025,N_27427);
nor U28196 (N_28196,N_27269,N_27107);
xnor U28197 (N_28197,N_27156,N_27007);
or U28198 (N_28198,N_27250,N_27428);
and U28199 (N_28199,N_27119,N_27576);
nand U28200 (N_28200,N_27623,N_28128);
nand U28201 (N_28201,N_27989,N_28179);
or U28202 (N_28202,N_27627,N_27991);
or U28203 (N_28203,N_28074,N_28014);
xnor U28204 (N_28204,N_27718,N_27935);
or U28205 (N_28205,N_27689,N_27653);
nand U28206 (N_28206,N_28133,N_27751);
xnor U28207 (N_28207,N_27695,N_28170);
nand U28208 (N_28208,N_27803,N_28083);
nor U28209 (N_28209,N_28071,N_27605);
xnor U28210 (N_28210,N_27643,N_27774);
or U28211 (N_28211,N_27773,N_28106);
xor U28212 (N_28212,N_27887,N_27811);
nor U28213 (N_28213,N_27668,N_27913);
and U28214 (N_28214,N_27859,N_27785);
xnor U28215 (N_28215,N_28099,N_27816);
and U28216 (N_28216,N_28173,N_27841);
nor U28217 (N_28217,N_27888,N_27618);
nor U28218 (N_28218,N_28078,N_27684);
and U28219 (N_28219,N_27647,N_27606);
nor U28220 (N_28220,N_27798,N_27840);
or U28221 (N_28221,N_27789,N_28108);
and U28222 (N_28222,N_27716,N_27719);
nor U28223 (N_28223,N_28116,N_27874);
and U28224 (N_28224,N_27973,N_27780);
or U28225 (N_28225,N_28144,N_27865);
xnor U28226 (N_28226,N_28080,N_28127);
nor U28227 (N_28227,N_27827,N_27796);
xor U28228 (N_28228,N_28183,N_28076);
xor U28229 (N_28229,N_28089,N_27748);
or U28230 (N_28230,N_27876,N_27686);
or U28231 (N_28231,N_27609,N_28160);
or U28232 (N_28232,N_28098,N_28045);
and U28233 (N_28233,N_27782,N_27885);
and U28234 (N_28234,N_28149,N_27934);
nor U28235 (N_28235,N_27897,N_27866);
nand U28236 (N_28236,N_27784,N_28015);
nand U28237 (N_28237,N_28181,N_28115);
nor U28238 (N_28238,N_27617,N_28086);
or U28239 (N_28239,N_27758,N_27725);
and U28240 (N_28240,N_27645,N_27769);
nand U28241 (N_28241,N_28085,N_27752);
nand U28242 (N_28242,N_27965,N_27633);
or U28243 (N_28243,N_27677,N_27616);
xnor U28244 (N_28244,N_27906,N_28152);
and U28245 (N_28245,N_27649,N_28069);
and U28246 (N_28246,N_27821,N_28130);
nand U28247 (N_28247,N_27786,N_27676);
nand U28248 (N_28248,N_27992,N_27799);
or U28249 (N_28249,N_27704,N_27914);
and U28250 (N_28250,N_27978,N_27928);
nand U28251 (N_28251,N_28112,N_27920);
nor U28252 (N_28252,N_27931,N_27851);
and U28253 (N_28253,N_27958,N_27937);
xnor U28254 (N_28254,N_28172,N_27714);
or U28255 (N_28255,N_27720,N_27967);
or U28256 (N_28256,N_27860,N_27947);
nor U28257 (N_28257,N_27916,N_28059);
nor U28258 (N_28258,N_27954,N_27926);
or U28259 (N_28259,N_27942,N_27619);
nor U28260 (N_28260,N_28138,N_27955);
nand U28261 (N_28261,N_28146,N_27766);
nand U28262 (N_28262,N_27895,N_27604);
nor U28263 (N_28263,N_27849,N_28122);
nor U28264 (N_28264,N_28189,N_27801);
and U28265 (N_28265,N_27857,N_27754);
and U28266 (N_28266,N_28066,N_28151);
and U28267 (N_28267,N_28162,N_27679);
nand U28268 (N_28268,N_27940,N_27834);
nand U28269 (N_28269,N_27662,N_27855);
and U28270 (N_28270,N_27731,N_27724);
xor U28271 (N_28271,N_27862,N_27950);
xnor U28272 (N_28272,N_27999,N_27659);
and U28273 (N_28273,N_27656,N_27912);
xor U28274 (N_28274,N_28140,N_27858);
and U28275 (N_28275,N_27867,N_27666);
nor U28276 (N_28276,N_28011,N_28057);
xnor U28277 (N_28277,N_28003,N_28020);
and U28278 (N_28278,N_27658,N_28145);
or U28279 (N_28279,N_28065,N_28126);
xnor U28280 (N_28280,N_27839,N_27744);
xor U28281 (N_28281,N_28185,N_28052);
or U28282 (N_28282,N_27702,N_27630);
and U28283 (N_28283,N_27750,N_28043);
and U28284 (N_28284,N_27898,N_27925);
nor U28285 (N_28285,N_28167,N_27815);
nor U28286 (N_28286,N_28018,N_27698);
nor U28287 (N_28287,N_27843,N_27753);
and U28288 (N_28288,N_27611,N_27878);
nor U28289 (N_28289,N_27673,N_28064);
nand U28290 (N_28290,N_27975,N_27995);
nor U28291 (N_28291,N_27621,N_27699);
nand U28292 (N_28292,N_28178,N_27941);
nor U28293 (N_28293,N_28087,N_27700);
or U28294 (N_28294,N_27644,N_28055);
nand U28295 (N_28295,N_28024,N_27842);
nand U28296 (N_28296,N_27688,N_27615);
and U28297 (N_28297,N_27831,N_27632);
or U28298 (N_28298,N_28072,N_28001);
nor U28299 (N_28299,N_27870,N_27911);
xnor U28300 (N_28300,N_28180,N_28171);
or U28301 (N_28301,N_27943,N_27997);
xnor U28302 (N_28302,N_27959,N_27655);
or U28303 (N_28303,N_28190,N_28082);
nor U28304 (N_28304,N_28104,N_28021);
nor U28305 (N_28305,N_27661,N_28168);
nand U28306 (N_28306,N_28081,N_27635);
nor U28307 (N_28307,N_27886,N_27850);
nor U28308 (N_28308,N_28034,N_27848);
xnor U28309 (N_28309,N_27740,N_27736);
nand U28310 (N_28310,N_27678,N_28118);
and U28311 (N_28311,N_27749,N_28051);
and U28312 (N_28312,N_27810,N_28060);
and U28313 (N_28313,N_27813,N_27902);
and U28314 (N_28314,N_27923,N_27838);
and U28315 (N_28315,N_27901,N_28123);
nand U28316 (N_28316,N_27880,N_27904);
nand U28317 (N_28317,N_28196,N_28134);
xnor U28318 (N_28318,N_28006,N_27847);
nand U28319 (N_28319,N_27809,N_27930);
xor U28320 (N_28320,N_27908,N_27951);
nor U28321 (N_28321,N_27891,N_27663);
or U28322 (N_28322,N_28025,N_28022);
and U28323 (N_28323,N_28191,N_27949);
nor U28324 (N_28324,N_27828,N_28046);
and U28325 (N_28325,N_27960,N_28166);
nand U28326 (N_28326,N_27979,N_27957);
and U28327 (N_28327,N_27833,N_27781);
nand U28328 (N_28328,N_27853,N_28120);
and U28329 (N_28329,N_27890,N_28195);
and U28330 (N_28330,N_27733,N_28016);
nand U28331 (N_28331,N_28163,N_27819);
and U28332 (N_28332,N_27685,N_27622);
and U28333 (N_28333,N_28048,N_27844);
and U28334 (N_28334,N_28062,N_28063);
or U28335 (N_28335,N_28174,N_28169);
xnor U28336 (N_28336,N_27936,N_27905);
nor U28337 (N_28337,N_28079,N_27787);
and U28338 (N_28338,N_28019,N_27835);
or U28339 (N_28339,N_27804,N_28027);
xnor U28340 (N_28340,N_27657,N_27963);
xnor U28341 (N_28341,N_27994,N_28036);
nand U28342 (N_28342,N_27654,N_27864);
and U28343 (N_28343,N_28142,N_27739);
nor U28344 (N_28344,N_27823,N_27756);
xor U28345 (N_28345,N_27800,N_27620);
nand U28346 (N_28346,N_28032,N_27927);
or U28347 (N_28347,N_28047,N_28092);
nand U28348 (N_28348,N_27812,N_28154);
and U28349 (N_28349,N_28070,N_27708);
nand U28350 (N_28350,N_28113,N_27696);
xnor U28351 (N_28351,N_27755,N_28155);
xnor U28352 (N_28352,N_27938,N_27778);
nor U28353 (N_28353,N_27712,N_27729);
xor U28354 (N_28354,N_27776,N_27875);
nor U28355 (N_28355,N_27775,N_28009);
and U28356 (N_28356,N_27741,N_27646);
and U28357 (N_28357,N_27993,N_28050);
and U28358 (N_28358,N_27721,N_27650);
and U28359 (N_28359,N_27939,N_27952);
nor U28360 (N_28360,N_27976,N_27956);
nand U28361 (N_28361,N_28007,N_27660);
nor U28362 (N_28362,N_28187,N_28157);
nand U28363 (N_28363,N_27665,N_28177);
or U28364 (N_28364,N_27770,N_27818);
or U28365 (N_28365,N_27760,N_27625);
or U28366 (N_28366,N_27613,N_27869);
xor U28367 (N_28367,N_28165,N_27889);
nand U28368 (N_28368,N_27664,N_27974);
nor U28369 (N_28369,N_27996,N_28010);
nor U28370 (N_28370,N_27987,N_28023);
nor U28371 (N_28371,N_28176,N_27814);
nand U28372 (N_28372,N_27624,N_28143);
nand U28373 (N_28373,N_28114,N_28041);
xor U28374 (N_28374,N_27797,N_27675);
nand U28375 (N_28375,N_28111,N_28061);
and U28376 (N_28376,N_27899,N_28198);
nor U28377 (N_28377,N_27612,N_28091);
or U28378 (N_28378,N_27610,N_28029);
or U28379 (N_28379,N_27919,N_28026);
or U28380 (N_28380,N_27948,N_27737);
and U28381 (N_28381,N_27969,N_27639);
nor U28382 (N_28382,N_27953,N_27795);
nor U28383 (N_28383,N_28199,N_27707);
or U28384 (N_28384,N_28049,N_27681);
and U28385 (N_28385,N_27907,N_27896);
or U28386 (N_28386,N_27998,N_28068);
or U28387 (N_28387,N_27697,N_27894);
nand U28388 (N_28388,N_27972,N_28073);
or U28389 (N_28389,N_28136,N_28004);
or U28390 (N_28390,N_27735,N_27674);
xor U28391 (N_28391,N_27817,N_28037);
or U28392 (N_28392,N_27881,N_27711);
or U28393 (N_28393,N_28175,N_27966);
nor U28394 (N_28394,N_27723,N_27691);
and U28395 (N_28395,N_27980,N_27832);
xor U28396 (N_28396,N_27727,N_27683);
xor U28397 (N_28397,N_27877,N_28186);
nor U28398 (N_28398,N_28161,N_28094);
xor U28399 (N_28399,N_27946,N_27682);
nand U28400 (N_28400,N_28139,N_28153);
nand U28401 (N_28401,N_27924,N_28054);
xnor U28402 (N_28402,N_28097,N_28058);
and U28403 (N_28403,N_28135,N_27779);
xor U28404 (N_28404,N_27767,N_27763);
xnor U28405 (N_28405,N_27693,N_28013);
or U28406 (N_28406,N_28192,N_27667);
and U28407 (N_28407,N_27694,N_28141);
nor U28408 (N_28408,N_28184,N_27670);
and U28409 (N_28409,N_27820,N_27873);
nor U28410 (N_28410,N_27636,N_27961);
nand U28411 (N_28411,N_27964,N_27764);
and U28412 (N_28412,N_27692,N_28148);
xnor U28413 (N_28413,N_27970,N_28008);
xor U28414 (N_28414,N_27824,N_27761);
xor U28415 (N_28415,N_28000,N_28084);
nor U28416 (N_28416,N_27822,N_27868);
xnor U28417 (N_28417,N_27871,N_27802);
nand U28418 (N_28418,N_27709,N_27757);
xor U28419 (N_28419,N_27984,N_27637);
xor U28420 (N_28420,N_28030,N_27672);
nand U28421 (N_28421,N_28090,N_27705);
xnor U28422 (N_28422,N_28125,N_27829);
nand U28423 (N_28423,N_28067,N_27900);
or U28424 (N_28424,N_27642,N_27701);
nand U28425 (N_28425,N_28044,N_27882);
or U28426 (N_28426,N_27845,N_27903);
or U28427 (N_28427,N_27768,N_27614);
or U28428 (N_28428,N_28005,N_28182);
or U28429 (N_28429,N_28102,N_27759);
nand U28430 (N_28430,N_27687,N_27745);
or U28431 (N_28431,N_27747,N_28194);
xor U28432 (N_28432,N_27772,N_27805);
xnor U28433 (N_28433,N_27634,N_27641);
and U28434 (N_28434,N_28156,N_27986);
or U28435 (N_28435,N_27791,N_28103);
nand U28436 (N_28436,N_28040,N_28053);
nor U28437 (N_28437,N_28002,N_28105);
nand U28438 (N_28438,N_27962,N_27893);
or U28439 (N_28439,N_28095,N_27713);
or U28440 (N_28440,N_27628,N_28131);
and U28441 (N_28441,N_27710,N_28110);
and U28442 (N_28442,N_27825,N_27730);
or U28443 (N_28443,N_27792,N_27602);
and U28444 (N_28444,N_27981,N_27790);
and U28445 (N_28445,N_27626,N_27917);
xor U28446 (N_28446,N_27807,N_27728);
and U28447 (N_28447,N_27783,N_28017);
nand U28448 (N_28448,N_27794,N_27703);
nor U28449 (N_28449,N_27884,N_27863);
xnor U28450 (N_28450,N_27892,N_28035);
xnor U28451 (N_28451,N_27746,N_28039);
and U28452 (N_28452,N_27856,N_27837);
and U28453 (N_28453,N_28033,N_27765);
nor U28454 (N_28454,N_28164,N_27717);
nor U28455 (N_28455,N_27680,N_27846);
nor U28456 (N_28456,N_28124,N_28137);
nor U28457 (N_28457,N_27910,N_27883);
or U28458 (N_28458,N_27671,N_27607);
or U28459 (N_28459,N_28147,N_27738);
nand U28460 (N_28460,N_27945,N_27706);
xnor U28461 (N_28461,N_27777,N_27944);
nand U28462 (N_28462,N_28042,N_27806);
nor U28463 (N_28463,N_27600,N_27861);
or U28464 (N_28464,N_27771,N_28075);
xor U28465 (N_28465,N_28197,N_27872);
and U28466 (N_28466,N_27985,N_28031);
nor U28467 (N_28467,N_28158,N_27742);
xnor U28468 (N_28468,N_27732,N_27879);
xnor U28469 (N_28469,N_27631,N_27601);
or U28470 (N_28470,N_27743,N_27968);
nand U28471 (N_28471,N_27652,N_28117);
xor U28472 (N_28472,N_27762,N_27629);
or U28473 (N_28473,N_27932,N_28088);
xor U28474 (N_28474,N_27722,N_28193);
and U28475 (N_28475,N_28129,N_27929);
nand U28476 (N_28476,N_27669,N_28188);
or U28477 (N_28477,N_27977,N_27734);
nand U28478 (N_28478,N_27651,N_27603);
or U28479 (N_28479,N_27971,N_28096);
nand U28480 (N_28480,N_27690,N_27648);
xnor U28481 (N_28481,N_27638,N_28121);
or U28482 (N_28482,N_27852,N_27808);
nand U28483 (N_28483,N_27854,N_27793);
or U28484 (N_28484,N_27836,N_28132);
xor U28485 (N_28485,N_27608,N_27909);
xnor U28486 (N_28486,N_27922,N_28038);
nor U28487 (N_28487,N_27826,N_28119);
xnor U28488 (N_28488,N_28077,N_27921);
nand U28489 (N_28489,N_27983,N_27982);
nor U28490 (N_28490,N_27788,N_27830);
nor U28491 (N_28491,N_27915,N_27726);
xnor U28492 (N_28492,N_28012,N_28028);
xnor U28493 (N_28493,N_27990,N_27933);
or U28494 (N_28494,N_28101,N_28150);
or U28495 (N_28495,N_27640,N_28100);
xnor U28496 (N_28496,N_28107,N_28056);
or U28497 (N_28497,N_27715,N_27918);
or U28498 (N_28498,N_27988,N_28093);
xor U28499 (N_28499,N_28159,N_28109);
nor U28500 (N_28500,N_27690,N_27637);
xor U28501 (N_28501,N_27794,N_27795);
nor U28502 (N_28502,N_27608,N_28138);
xnor U28503 (N_28503,N_27725,N_27907);
or U28504 (N_28504,N_28001,N_27664);
and U28505 (N_28505,N_27969,N_28121);
xor U28506 (N_28506,N_27900,N_27945);
nand U28507 (N_28507,N_27898,N_28086);
or U28508 (N_28508,N_27848,N_27815);
nand U28509 (N_28509,N_28169,N_27902);
and U28510 (N_28510,N_27923,N_28107);
nor U28511 (N_28511,N_27741,N_28024);
and U28512 (N_28512,N_27906,N_28149);
xnor U28513 (N_28513,N_27636,N_27615);
xor U28514 (N_28514,N_27941,N_27936);
nor U28515 (N_28515,N_28157,N_27702);
or U28516 (N_28516,N_27882,N_28086);
and U28517 (N_28517,N_27881,N_27936);
and U28518 (N_28518,N_27755,N_27639);
nand U28519 (N_28519,N_27785,N_27978);
or U28520 (N_28520,N_27626,N_27662);
nor U28521 (N_28521,N_27954,N_27631);
xor U28522 (N_28522,N_27802,N_27983);
nand U28523 (N_28523,N_27827,N_28040);
nor U28524 (N_28524,N_27773,N_27670);
and U28525 (N_28525,N_27867,N_27611);
nor U28526 (N_28526,N_27682,N_27888);
nand U28527 (N_28527,N_27618,N_27641);
and U28528 (N_28528,N_28120,N_27679);
nor U28529 (N_28529,N_27836,N_27731);
xor U28530 (N_28530,N_28143,N_27786);
xnor U28531 (N_28531,N_28144,N_27928);
or U28532 (N_28532,N_28131,N_27967);
nor U28533 (N_28533,N_28100,N_27879);
and U28534 (N_28534,N_28018,N_27612);
and U28535 (N_28535,N_27687,N_27668);
nand U28536 (N_28536,N_28124,N_27750);
or U28537 (N_28537,N_28040,N_27666);
and U28538 (N_28538,N_27830,N_27802);
xnor U28539 (N_28539,N_27913,N_27804);
nand U28540 (N_28540,N_27648,N_27861);
nor U28541 (N_28541,N_27923,N_28003);
nor U28542 (N_28542,N_27773,N_27758);
or U28543 (N_28543,N_27626,N_27853);
or U28544 (N_28544,N_27839,N_27940);
xor U28545 (N_28545,N_27889,N_28169);
and U28546 (N_28546,N_27895,N_28164);
nor U28547 (N_28547,N_28026,N_27776);
xnor U28548 (N_28548,N_27676,N_28000);
and U28549 (N_28549,N_28078,N_27789);
xnor U28550 (N_28550,N_27858,N_28023);
nor U28551 (N_28551,N_27886,N_27961);
xnor U28552 (N_28552,N_27756,N_28158);
xnor U28553 (N_28553,N_27904,N_27743);
nand U28554 (N_28554,N_27794,N_27717);
or U28555 (N_28555,N_28091,N_27886);
nor U28556 (N_28556,N_27655,N_27653);
nor U28557 (N_28557,N_27791,N_27848);
or U28558 (N_28558,N_27818,N_28143);
or U28559 (N_28559,N_27783,N_27624);
nand U28560 (N_28560,N_27786,N_28021);
or U28561 (N_28561,N_27798,N_28037);
nor U28562 (N_28562,N_27954,N_28106);
and U28563 (N_28563,N_28151,N_28188);
nor U28564 (N_28564,N_27655,N_27602);
xor U28565 (N_28565,N_27987,N_28073);
nor U28566 (N_28566,N_28071,N_28179);
nor U28567 (N_28567,N_28001,N_27701);
and U28568 (N_28568,N_27804,N_28123);
nand U28569 (N_28569,N_27731,N_28148);
and U28570 (N_28570,N_28096,N_28152);
nand U28571 (N_28571,N_27968,N_28128);
or U28572 (N_28572,N_28167,N_27866);
xor U28573 (N_28573,N_28155,N_28176);
or U28574 (N_28574,N_27660,N_27925);
and U28575 (N_28575,N_27806,N_27886);
xnor U28576 (N_28576,N_27761,N_27917);
and U28577 (N_28577,N_28127,N_27780);
nand U28578 (N_28578,N_27770,N_27734);
nand U28579 (N_28579,N_28000,N_28042);
xnor U28580 (N_28580,N_27998,N_27942);
and U28581 (N_28581,N_27700,N_28119);
nor U28582 (N_28582,N_27832,N_27932);
or U28583 (N_28583,N_28156,N_27925);
nor U28584 (N_28584,N_28082,N_27689);
and U28585 (N_28585,N_27688,N_28138);
nand U28586 (N_28586,N_27738,N_27731);
nor U28587 (N_28587,N_27656,N_27773);
and U28588 (N_28588,N_28031,N_28197);
xor U28589 (N_28589,N_28177,N_27642);
or U28590 (N_28590,N_27749,N_27878);
nor U28591 (N_28591,N_27918,N_27919);
xnor U28592 (N_28592,N_27746,N_27817);
xor U28593 (N_28593,N_28122,N_28080);
nor U28594 (N_28594,N_28066,N_28191);
or U28595 (N_28595,N_28061,N_27609);
nand U28596 (N_28596,N_27813,N_28146);
or U28597 (N_28597,N_27771,N_27923);
nor U28598 (N_28598,N_27979,N_27912);
nand U28599 (N_28599,N_27645,N_27743);
and U28600 (N_28600,N_27955,N_28167);
xor U28601 (N_28601,N_27710,N_27749);
nor U28602 (N_28602,N_28150,N_28170);
or U28603 (N_28603,N_27834,N_27620);
or U28604 (N_28604,N_28007,N_27771);
nand U28605 (N_28605,N_27965,N_27856);
and U28606 (N_28606,N_27689,N_27926);
nor U28607 (N_28607,N_27912,N_28139);
and U28608 (N_28608,N_27710,N_27640);
nor U28609 (N_28609,N_27807,N_27911);
nand U28610 (N_28610,N_27755,N_27706);
nand U28611 (N_28611,N_27811,N_28180);
nand U28612 (N_28612,N_28171,N_27732);
nand U28613 (N_28613,N_28031,N_28021);
nand U28614 (N_28614,N_28111,N_28051);
or U28615 (N_28615,N_28077,N_28081);
nor U28616 (N_28616,N_27752,N_28198);
xor U28617 (N_28617,N_28190,N_27807);
nand U28618 (N_28618,N_28053,N_28162);
and U28619 (N_28619,N_28139,N_28085);
or U28620 (N_28620,N_28005,N_27914);
or U28621 (N_28621,N_28127,N_28150);
nand U28622 (N_28622,N_28001,N_28144);
or U28623 (N_28623,N_27881,N_27878);
or U28624 (N_28624,N_27706,N_27786);
or U28625 (N_28625,N_27606,N_28164);
or U28626 (N_28626,N_28190,N_27709);
xnor U28627 (N_28627,N_27739,N_27806);
or U28628 (N_28628,N_27804,N_27925);
xnor U28629 (N_28629,N_27840,N_27865);
nor U28630 (N_28630,N_27721,N_27781);
or U28631 (N_28631,N_28164,N_28090);
nand U28632 (N_28632,N_28152,N_28070);
nor U28633 (N_28633,N_27980,N_28091);
nor U28634 (N_28634,N_27706,N_28127);
nor U28635 (N_28635,N_28074,N_27677);
and U28636 (N_28636,N_27799,N_27739);
or U28637 (N_28637,N_27895,N_28119);
or U28638 (N_28638,N_28051,N_27854);
or U28639 (N_28639,N_28092,N_27763);
xor U28640 (N_28640,N_28079,N_28102);
or U28641 (N_28641,N_28115,N_28139);
xnor U28642 (N_28642,N_27896,N_28061);
or U28643 (N_28643,N_27981,N_27632);
or U28644 (N_28644,N_27907,N_27903);
xor U28645 (N_28645,N_27989,N_27906);
nand U28646 (N_28646,N_28189,N_27770);
xnor U28647 (N_28647,N_27799,N_27842);
nor U28648 (N_28648,N_27651,N_28015);
or U28649 (N_28649,N_28026,N_28159);
nand U28650 (N_28650,N_28145,N_28059);
nor U28651 (N_28651,N_27789,N_28091);
xor U28652 (N_28652,N_28090,N_28036);
nand U28653 (N_28653,N_27604,N_28000);
nand U28654 (N_28654,N_28012,N_27875);
xnor U28655 (N_28655,N_28019,N_27764);
xnor U28656 (N_28656,N_27902,N_28078);
nor U28657 (N_28657,N_28153,N_27670);
xnor U28658 (N_28658,N_27800,N_27601);
nor U28659 (N_28659,N_28053,N_27771);
or U28660 (N_28660,N_28016,N_28123);
and U28661 (N_28661,N_27769,N_27643);
xor U28662 (N_28662,N_28156,N_27995);
or U28663 (N_28663,N_27787,N_28093);
nand U28664 (N_28664,N_27678,N_27962);
and U28665 (N_28665,N_27895,N_28128);
or U28666 (N_28666,N_27619,N_27985);
xor U28667 (N_28667,N_27675,N_27643);
or U28668 (N_28668,N_28135,N_28009);
or U28669 (N_28669,N_27792,N_27695);
or U28670 (N_28670,N_27997,N_27702);
nor U28671 (N_28671,N_27665,N_27981);
xnor U28672 (N_28672,N_27909,N_27712);
xnor U28673 (N_28673,N_27730,N_28132);
or U28674 (N_28674,N_27973,N_27691);
and U28675 (N_28675,N_27804,N_27996);
xnor U28676 (N_28676,N_28146,N_27838);
nand U28677 (N_28677,N_27935,N_27736);
nor U28678 (N_28678,N_27912,N_28034);
and U28679 (N_28679,N_27895,N_27736);
nand U28680 (N_28680,N_27903,N_28078);
nor U28681 (N_28681,N_27746,N_27982);
nand U28682 (N_28682,N_27761,N_28037);
xor U28683 (N_28683,N_27971,N_27802);
xnor U28684 (N_28684,N_27711,N_27937);
or U28685 (N_28685,N_28054,N_27830);
nand U28686 (N_28686,N_27702,N_27965);
and U28687 (N_28687,N_27616,N_28062);
or U28688 (N_28688,N_27810,N_27644);
xor U28689 (N_28689,N_27655,N_27876);
or U28690 (N_28690,N_28180,N_28187);
nor U28691 (N_28691,N_28021,N_28162);
nor U28692 (N_28692,N_27790,N_27806);
or U28693 (N_28693,N_27718,N_27944);
nand U28694 (N_28694,N_27870,N_27839);
and U28695 (N_28695,N_27813,N_28199);
and U28696 (N_28696,N_27750,N_28042);
nor U28697 (N_28697,N_28038,N_27842);
or U28698 (N_28698,N_27825,N_27646);
and U28699 (N_28699,N_27782,N_28147);
nand U28700 (N_28700,N_28165,N_27923);
nor U28701 (N_28701,N_27901,N_27845);
or U28702 (N_28702,N_27609,N_27897);
xnor U28703 (N_28703,N_27703,N_27942);
xnor U28704 (N_28704,N_27811,N_27837);
and U28705 (N_28705,N_28143,N_28040);
or U28706 (N_28706,N_27754,N_27886);
nand U28707 (N_28707,N_27847,N_28075);
or U28708 (N_28708,N_27932,N_28043);
xor U28709 (N_28709,N_28177,N_27879);
xor U28710 (N_28710,N_28170,N_27927);
and U28711 (N_28711,N_27613,N_28008);
and U28712 (N_28712,N_28075,N_27748);
or U28713 (N_28713,N_27924,N_27952);
or U28714 (N_28714,N_28057,N_27872);
nand U28715 (N_28715,N_27839,N_28065);
or U28716 (N_28716,N_27700,N_27761);
nand U28717 (N_28717,N_27654,N_27956);
xor U28718 (N_28718,N_28150,N_27715);
nand U28719 (N_28719,N_27731,N_28167);
nand U28720 (N_28720,N_27720,N_28116);
and U28721 (N_28721,N_28148,N_27702);
nand U28722 (N_28722,N_27773,N_28178);
nand U28723 (N_28723,N_27822,N_27834);
or U28724 (N_28724,N_27865,N_27710);
nor U28725 (N_28725,N_27764,N_28036);
nand U28726 (N_28726,N_27687,N_27728);
nor U28727 (N_28727,N_27898,N_28062);
nor U28728 (N_28728,N_27696,N_28182);
nand U28729 (N_28729,N_28110,N_27625);
xnor U28730 (N_28730,N_28029,N_28071);
xnor U28731 (N_28731,N_28116,N_27661);
and U28732 (N_28732,N_27680,N_27891);
or U28733 (N_28733,N_28024,N_27921);
nand U28734 (N_28734,N_27616,N_27893);
or U28735 (N_28735,N_27790,N_27966);
xor U28736 (N_28736,N_27874,N_28049);
or U28737 (N_28737,N_28010,N_28154);
and U28738 (N_28738,N_28159,N_27818);
nor U28739 (N_28739,N_28178,N_27899);
nand U28740 (N_28740,N_28177,N_27958);
nand U28741 (N_28741,N_27829,N_28189);
nor U28742 (N_28742,N_27706,N_27653);
nor U28743 (N_28743,N_27861,N_27912);
or U28744 (N_28744,N_28035,N_27652);
nor U28745 (N_28745,N_27652,N_28039);
nor U28746 (N_28746,N_27978,N_28062);
or U28747 (N_28747,N_28052,N_28091);
nor U28748 (N_28748,N_27775,N_28085);
or U28749 (N_28749,N_28184,N_27657);
or U28750 (N_28750,N_27646,N_27857);
nor U28751 (N_28751,N_27616,N_27684);
xor U28752 (N_28752,N_27848,N_27708);
nor U28753 (N_28753,N_28138,N_27711);
xor U28754 (N_28754,N_27970,N_28145);
nand U28755 (N_28755,N_27998,N_28002);
or U28756 (N_28756,N_28019,N_27948);
nand U28757 (N_28757,N_28039,N_27653);
xor U28758 (N_28758,N_27986,N_28017);
nand U28759 (N_28759,N_27917,N_28183);
xor U28760 (N_28760,N_28084,N_27810);
nand U28761 (N_28761,N_27943,N_27648);
or U28762 (N_28762,N_27649,N_27971);
xor U28763 (N_28763,N_28038,N_27675);
nor U28764 (N_28764,N_27881,N_27746);
xor U28765 (N_28765,N_27948,N_28007);
xor U28766 (N_28766,N_27896,N_27979);
nor U28767 (N_28767,N_27960,N_28155);
and U28768 (N_28768,N_27885,N_27680);
xnor U28769 (N_28769,N_28096,N_27633);
nand U28770 (N_28770,N_27882,N_28148);
and U28771 (N_28771,N_27988,N_27966);
xnor U28772 (N_28772,N_27856,N_28066);
nor U28773 (N_28773,N_27604,N_27888);
and U28774 (N_28774,N_27808,N_27785);
and U28775 (N_28775,N_27783,N_28193);
and U28776 (N_28776,N_28187,N_27797);
nor U28777 (N_28777,N_27651,N_27895);
or U28778 (N_28778,N_28179,N_28009);
xor U28779 (N_28779,N_27769,N_27931);
nand U28780 (N_28780,N_27956,N_28054);
nand U28781 (N_28781,N_27784,N_27768);
nand U28782 (N_28782,N_27751,N_27942);
nor U28783 (N_28783,N_27619,N_27998);
xor U28784 (N_28784,N_27732,N_27623);
nor U28785 (N_28785,N_27752,N_27976);
xor U28786 (N_28786,N_27635,N_28146);
xor U28787 (N_28787,N_27753,N_27754);
and U28788 (N_28788,N_27791,N_28044);
nor U28789 (N_28789,N_27740,N_27687);
nor U28790 (N_28790,N_28101,N_27689);
or U28791 (N_28791,N_28064,N_28083);
xnor U28792 (N_28792,N_27679,N_27718);
or U28793 (N_28793,N_27937,N_27823);
nand U28794 (N_28794,N_28057,N_27624);
nor U28795 (N_28795,N_28087,N_27858);
and U28796 (N_28796,N_28075,N_27933);
xor U28797 (N_28797,N_27719,N_27858);
nor U28798 (N_28798,N_27985,N_27927);
and U28799 (N_28799,N_27781,N_28010);
or U28800 (N_28800,N_28365,N_28399);
xnor U28801 (N_28801,N_28412,N_28648);
and U28802 (N_28802,N_28600,N_28368);
xor U28803 (N_28803,N_28567,N_28263);
and U28804 (N_28804,N_28764,N_28446);
xor U28805 (N_28805,N_28409,N_28612);
xor U28806 (N_28806,N_28233,N_28715);
and U28807 (N_28807,N_28675,N_28563);
nand U28808 (N_28808,N_28571,N_28492);
nand U28809 (N_28809,N_28255,N_28654);
and U28810 (N_28810,N_28331,N_28423);
nand U28811 (N_28811,N_28302,N_28433);
or U28812 (N_28812,N_28538,N_28685);
xnor U28813 (N_28813,N_28531,N_28754);
or U28814 (N_28814,N_28630,N_28551);
nand U28815 (N_28815,N_28617,N_28561);
xnor U28816 (N_28816,N_28311,N_28496);
xor U28817 (N_28817,N_28213,N_28592);
or U28818 (N_28818,N_28658,N_28320);
nor U28819 (N_28819,N_28798,N_28204);
nand U28820 (N_28820,N_28393,N_28521);
nand U28821 (N_28821,N_28436,N_28580);
and U28822 (N_28822,N_28757,N_28363);
xnor U28823 (N_28823,N_28301,N_28208);
nand U28824 (N_28824,N_28625,N_28408);
and U28825 (N_28825,N_28540,N_28297);
nand U28826 (N_28826,N_28400,N_28366);
or U28827 (N_28827,N_28513,N_28488);
and U28828 (N_28828,N_28618,N_28799);
or U28829 (N_28829,N_28598,N_28464);
or U28830 (N_28830,N_28495,N_28448);
xnor U28831 (N_28831,N_28265,N_28307);
or U28832 (N_28832,N_28471,N_28383);
nor U28833 (N_28833,N_28766,N_28321);
nand U28834 (N_28834,N_28609,N_28639);
nor U28835 (N_28835,N_28678,N_28437);
nor U28836 (N_28836,N_28696,N_28793);
or U28837 (N_28837,N_28681,N_28278);
nand U28838 (N_28838,N_28646,N_28699);
or U28839 (N_28839,N_28355,N_28276);
and U28840 (N_28840,N_28642,N_28740);
and U28841 (N_28841,N_28586,N_28629);
nor U28842 (N_28842,N_28419,N_28323);
and U28843 (N_28843,N_28362,N_28677);
or U28844 (N_28844,N_28673,N_28640);
and U28845 (N_28845,N_28421,N_28207);
or U28846 (N_28846,N_28761,N_28398);
nor U28847 (N_28847,N_28657,N_28282);
xnor U28848 (N_28848,N_28522,N_28294);
and U28849 (N_28849,N_28298,N_28367);
and U28850 (N_28850,N_28728,N_28432);
and U28851 (N_28851,N_28337,N_28425);
or U28852 (N_28852,N_28403,N_28281);
nand U28853 (N_28853,N_28482,N_28529);
xor U28854 (N_28854,N_28442,N_28633);
nor U28855 (N_28855,N_28410,N_28303);
nor U28856 (N_28856,N_28634,N_28315);
nor U28857 (N_28857,N_28792,N_28309);
xor U28858 (N_28858,N_28552,N_28268);
and U28859 (N_28859,N_28553,N_28261);
and U28860 (N_28860,N_28631,N_28287);
or U28861 (N_28861,N_28656,N_28645);
xor U28862 (N_28862,N_28735,N_28486);
nor U28863 (N_28863,N_28568,N_28418);
xor U28864 (N_28864,N_28209,N_28379);
and U28865 (N_28865,N_28576,N_28284);
nand U28866 (N_28866,N_28716,N_28719);
nor U28867 (N_28867,N_28259,N_28542);
or U28868 (N_28868,N_28463,N_28245);
xnor U28869 (N_28869,N_28416,N_28733);
nand U28870 (N_28870,N_28290,N_28304);
xor U28871 (N_28871,N_28653,N_28435);
nand U28872 (N_28872,N_28546,N_28539);
xnor U28873 (N_28873,N_28777,N_28732);
nand U28874 (N_28874,N_28701,N_28756);
nand U28875 (N_28875,N_28234,N_28385);
or U28876 (N_28876,N_28246,N_28687);
and U28877 (N_28877,N_28288,N_28790);
xnor U28878 (N_28878,N_28316,N_28344);
nor U28879 (N_28879,N_28623,N_28351);
and U28880 (N_28880,N_28594,N_28588);
or U28881 (N_28881,N_28326,N_28229);
nand U28882 (N_28882,N_28387,N_28606);
nor U28883 (N_28883,N_28396,N_28490);
nand U28884 (N_28884,N_28342,N_28671);
nand U28885 (N_28885,N_28724,N_28478);
nor U28886 (N_28886,N_28256,N_28784);
or U28887 (N_28887,N_28796,N_28370);
xor U28888 (N_28888,N_28781,N_28550);
or U28889 (N_28889,N_28565,N_28655);
nand U28890 (N_28890,N_28610,N_28575);
xor U28891 (N_28891,N_28557,N_28258);
nand U28892 (N_28892,N_28200,N_28688);
or U28893 (N_28893,N_28498,N_28750);
nand U28894 (N_28894,N_28212,N_28447);
nor U28895 (N_28895,N_28686,N_28374);
and U28896 (N_28896,N_28534,N_28581);
xor U28897 (N_28897,N_28264,N_28573);
nor U28898 (N_28898,N_28248,N_28267);
and U28899 (N_28899,N_28720,N_28202);
nand U28900 (N_28900,N_28308,N_28242);
nor U28901 (N_28901,N_28704,N_28449);
xor U28902 (N_28902,N_28520,N_28438);
xor U28903 (N_28903,N_28599,N_28584);
and U28904 (N_28904,N_28455,N_28462);
nor U28905 (N_28905,N_28613,N_28417);
or U28906 (N_28906,N_28397,N_28273);
nor U28907 (N_28907,N_28205,N_28707);
xor U28908 (N_28908,N_28661,N_28743);
nor U28909 (N_28909,N_28774,N_28348);
nand U28910 (N_28910,N_28649,N_28601);
or U28911 (N_28911,N_28770,N_28730);
nor U28912 (N_28912,N_28663,N_28558);
and U28913 (N_28913,N_28439,N_28786);
nor U28914 (N_28914,N_28747,N_28411);
xnor U28915 (N_28915,N_28477,N_28289);
xnor U28916 (N_28916,N_28611,N_28357);
and U28917 (N_28917,N_28221,N_28660);
and U28918 (N_28918,N_28505,N_28746);
xor U28919 (N_28919,N_28440,N_28773);
nor U28920 (N_28920,N_28783,N_28672);
nand U28921 (N_28921,N_28401,N_28238);
nor U28922 (N_28922,N_28483,N_28252);
xor U28923 (N_28923,N_28624,N_28347);
or U28924 (N_28924,N_28314,N_28748);
nor U28925 (N_28925,N_28578,N_28525);
nand U28926 (N_28926,N_28335,N_28402);
nand U28927 (N_28927,N_28420,N_28532);
xor U28928 (N_28928,N_28758,N_28726);
xor U28929 (N_28929,N_28262,N_28605);
and U28930 (N_28930,N_28241,N_28484);
nor U28931 (N_28931,N_28591,N_28349);
or U28932 (N_28932,N_28797,N_28459);
nand U28933 (N_28933,N_28710,N_28514);
or U28934 (N_28934,N_28547,N_28723);
xor U28935 (N_28935,N_28371,N_28493);
nand U28936 (N_28936,N_28216,N_28711);
nor U28937 (N_28937,N_28583,N_28380);
nand U28938 (N_28938,N_28451,N_28562);
nand U28939 (N_28939,N_28251,N_28406);
and U28940 (N_28940,N_28293,N_28690);
nand U28941 (N_28941,N_28560,N_28407);
xor U28942 (N_28942,N_28731,N_28249);
or U28943 (N_28943,N_28239,N_28501);
xor U28944 (N_28944,N_28373,N_28377);
xor U28945 (N_28945,N_28668,N_28266);
nand U28946 (N_28946,N_28689,N_28779);
nand U28947 (N_28947,N_28306,N_28339);
or U28948 (N_28948,N_28322,N_28595);
and U28949 (N_28949,N_28776,N_28780);
nand U28950 (N_28950,N_28674,N_28280);
nor U28951 (N_28951,N_28340,N_28622);
nor U28952 (N_28952,N_28211,N_28788);
nor U28953 (N_28953,N_28507,N_28745);
and U28954 (N_28954,N_28332,N_28669);
nor U28955 (N_28955,N_28523,N_28620);
and U28956 (N_28956,N_28555,N_28712);
nor U28957 (N_28957,N_28222,N_28574);
or U28958 (N_28958,N_28452,N_28358);
and U28959 (N_28959,N_28424,N_28789);
xnor U28960 (N_28960,N_28260,N_28607);
nor U28961 (N_28961,N_28794,N_28369);
or U28962 (N_28962,N_28736,N_28299);
and U28963 (N_28963,N_28354,N_28384);
and U28964 (N_28964,N_28670,N_28577);
xnor U28965 (N_28965,N_28422,N_28215);
xor U28966 (N_28966,N_28392,N_28231);
and U28967 (N_28967,N_28643,N_28705);
or U28968 (N_28968,N_28738,N_28760);
nand U28969 (N_28969,N_28537,N_28388);
or U28970 (N_28970,N_28458,N_28692);
xnor U28971 (N_28971,N_28635,N_28706);
xnor U28972 (N_28972,N_28698,N_28697);
nor U28973 (N_28973,N_28503,N_28554);
nor U28974 (N_28974,N_28556,N_28253);
and U28975 (N_28975,N_28772,N_28785);
xor U28976 (N_28976,N_28721,N_28404);
or U28977 (N_28977,N_28381,N_28206);
xnor U28978 (N_28978,N_28460,N_28637);
nand U28979 (N_28979,N_28694,N_28257);
nor U28980 (N_28980,N_28317,N_28682);
xor U28981 (N_28981,N_28389,N_28566);
or U28982 (N_28982,N_28450,N_28667);
nor U28983 (N_28983,N_28765,N_28327);
xnor U28984 (N_28984,N_28286,N_28312);
xnor U28985 (N_28985,N_28214,N_28352);
and U28986 (N_28986,N_28430,N_28596);
xnor U28987 (N_28987,N_28627,N_28338);
and U28988 (N_28988,N_28664,N_28666);
or U28989 (N_28989,N_28269,N_28545);
and U28990 (N_28990,N_28579,N_28644);
or U28991 (N_28991,N_28376,N_28589);
or U28992 (N_28992,N_28517,N_28227);
or U28993 (N_28993,N_28481,N_28519);
xor U28994 (N_28994,N_28461,N_28472);
or U28995 (N_28995,N_28230,N_28465);
xor U28996 (N_28996,N_28378,N_28441);
or U28997 (N_28997,N_28457,N_28203);
and U28998 (N_28998,N_28585,N_28787);
and U28999 (N_28999,N_28235,N_28469);
nor U29000 (N_29000,N_28386,N_28341);
and U29001 (N_29001,N_28359,N_28489);
nand U29002 (N_29002,N_28751,N_28722);
nor U29003 (N_29003,N_28587,N_28621);
nand U29004 (N_29004,N_28626,N_28744);
or U29005 (N_29005,N_28602,N_28665);
or U29006 (N_29006,N_28528,N_28375);
xor U29007 (N_29007,N_28703,N_28691);
and U29008 (N_29008,N_28454,N_28564);
nand U29009 (N_29009,N_28527,N_28742);
and U29010 (N_29010,N_28487,N_28778);
or U29011 (N_29011,N_28467,N_28695);
xnor U29012 (N_29012,N_28572,N_28608);
xnor U29013 (N_29013,N_28508,N_28725);
nand U29014 (N_29014,N_28453,N_28782);
nor U29015 (N_29015,N_28524,N_28734);
nor U29016 (N_29016,N_28479,N_28346);
and U29017 (N_29017,N_28741,N_28313);
nor U29018 (N_29018,N_28714,N_28755);
xnor U29019 (N_29019,N_28718,N_28510);
or U29020 (N_29020,N_28391,N_28717);
xor U29021 (N_29021,N_28739,N_28499);
and U29022 (N_29022,N_28291,N_28456);
nor U29023 (N_29023,N_28651,N_28659);
and U29024 (N_29024,N_28218,N_28413);
nand U29025 (N_29025,N_28769,N_28762);
xnor U29026 (N_29026,N_28541,N_28274);
xnor U29027 (N_29027,N_28570,N_28443);
nor U29028 (N_29028,N_28559,N_28597);
nand U29029 (N_29029,N_28619,N_28791);
nand U29030 (N_29030,N_28243,N_28217);
nand U29031 (N_29031,N_28353,N_28533);
and U29032 (N_29032,N_28727,N_28210);
nand U29033 (N_29033,N_28426,N_28300);
or U29034 (N_29034,N_28614,N_28350);
nand U29035 (N_29035,N_28535,N_28641);
nand U29036 (N_29036,N_28247,N_28737);
and U29037 (N_29037,N_28593,N_28476);
nand U29038 (N_29038,N_28271,N_28237);
xor U29039 (N_29039,N_28431,N_28530);
xor U29040 (N_29040,N_28310,N_28636);
xnor U29041 (N_29041,N_28676,N_28662);
nand U29042 (N_29042,N_28753,N_28395);
nand U29043 (N_29043,N_28473,N_28650);
nand U29044 (N_29044,N_28232,N_28224);
or U29045 (N_29045,N_28356,N_28485);
and U29046 (N_29046,N_28445,N_28491);
or U29047 (N_29047,N_28709,N_28292);
nand U29048 (N_29048,N_28394,N_28516);
and U29049 (N_29049,N_28604,N_28512);
nand U29050 (N_29050,N_28228,N_28647);
nor U29051 (N_29051,N_28763,N_28548);
nand U29052 (N_29052,N_28223,N_28480);
nor U29053 (N_29053,N_28285,N_28504);
and U29054 (N_29054,N_28468,N_28713);
nor U29055 (N_29055,N_28767,N_28582);
nand U29056 (N_29056,N_28771,N_28325);
or U29057 (N_29057,N_28240,N_28225);
and U29058 (N_29058,N_28795,N_28700);
or U29059 (N_29059,N_28506,N_28768);
and U29060 (N_29060,N_28277,N_28270);
and U29061 (N_29061,N_28638,N_28345);
xnor U29062 (N_29062,N_28749,N_28708);
nor U29063 (N_29063,N_28543,N_28759);
nor U29064 (N_29064,N_28318,N_28500);
xor U29065 (N_29065,N_28511,N_28679);
nor U29066 (N_29066,N_28680,N_28549);
nand U29067 (N_29067,N_28272,N_28336);
or U29068 (N_29068,N_28615,N_28693);
or U29069 (N_29069,N_28497,N_28683);
nor U29070 (N_29070,N_28390,N_28360);
nor U29071 (N_29071,N_28515,N_28474);
xor U29072 (N_29072,N_28415,N_28382);
nand U29073 (N_29073,N_28329,N_28466);
nor U29074 (N_29074,N_28279,N_28428);
nor U29075 (N_29075,N_28405,N_28319);
xor U29076 (N_29076,N_28632,N_28470);
xor U29077 (N_29077,N_28334,N_28226);
xor U29078 (N_29078,N_28444,N_28429);
and U29079 (N_29079,N_28250,N_28729);
or U29080 (N_29080,N_28364,N_28333);
nor U29081 (N_29081,N_28414,N_28244);
xnor U29082 (N_29082,N_28343,N_28361);
and U29083 (N_29083,N_28518,N_28502);
or U29084 (N_29084,N_28702,N_28590);
nor U29085 (N_29085,N_28569,N_28544);
nor U29086 (N_29086,N_28427,N_28434);
nand U29087 (N_29087,N_28628,N_28219);
nand U29088 (N_29088,N_28526,N_28254);
nand U29089 (N_29089,N_28305,N_28752);
nor U29090 (N_29090,N_28372,N_28330);
or U29091 (N_29091,N_28220,N_28775);
xnor U29092 (N_29092,N_28536,N_28494);
or U29093 (N_29093,N_28475,N_28283);
and U29094 (N_29094,N_28616,N_28603);
nor U29095 (N_29095,N_28652,N_28275);
xnor U29096 (N_29096,N_28509,N_28296);
or U29097 (N_29097,N_28684,N_28236);
xor U29098 (N_29098,N_28324,N_28295);
xor U29099 (N_29099,N_28201,N_28328);
or U29100 (N_29100,N_28564,N_28642);
xor U29101 (N_29101,N_28637,N_28581);
or U29102 (N_29102,N_28321,N_28507);
nor U29103 (N_29103,N_28715,N_28788);
nor U29104 (N_29104,N_28782,N_28444);
nor U29105 (N_29105,N_28307,N_28647);
nand U29106 (N_29106,N_28527,N_28650);
nor U29107 (N_29107,N_28318,N_28592);
xor U29108 (N_29108,N_28498,N_28669);
nand U29109 (N_29109,N_28737,N_28524);
and U29110 (N_29110,N_28625,N_28243);
nand U29111 (N_29111,N_28778,N_28498);
nand U29112 (N_29112,N_28570,N_28358);
nor U29113 (N_29113,N_28796,N_28619);
or U29114 (N_29114,N_28681,N_28341);
xnor U29115 (N_29115,N_28565,N_28223);
or U29116 (N_29116,N_28360,N_28309);
xnor U29117 (N_29117,N_28797,N_28687);
nand U29118 (N_29118,N_28766,N_28524);
and U29119 (N_29119,N_28268,N_28696);
or U29120 (N_29120,N_28737,N_28428);
and U29121 (N_29121,N_28426,N_28470);
and U29122 (N_29122,N_28775,N_28426);
or U29123 (N_29123,N_28324,N_28770);
nor U29124 (N_29124,N_28673,N_28420);
nor U29125 (N_29125,N_28256,N_28632);
or U29126 (N_29126,N_28786,N_28793);
or U29127 (N_29127,N_28235,N_28679);
or U29128 (N_29128,N_28401,N_28435);
xor U29129 (N_29129,N_28341,N_28221);
xor U29130 (N_29130,N_28607,N_28438);
nor U29131 (N_29131,N_28292,N_28477);
and U29132 (N_29132,N_28273,N_28712);
xnor U29133 (N_29133,N_28793,N_28407);
nor U29134 (N_29134,N_28657,N_28204);
or U29135 (N_29135,N_28428,N_28476);
xnor U29136 (N_29136,N_28764,N_28531);
or U29137 (N_29137,N_28798,N_28221);
or U29138 (N_29138,N_28404,N_28372);
nor U29139 (N_29139,N_28521,N_28341);
xnor U29140 (N_29140,N_28573,N_28254);
xnor U29141 (N_29141,N_28539,N_28487);
or U29142 (N_29142,N_28483,N_28216);
nor U29143 (N_29143,N_28552,N_28271);
or U29144 (N_29144,N_28565,N_28392);
or U29145 (N_29145,N_28374,N_28615);
nand U29146 (N_29146,N_28660,N_28533);
nor U29147 (N_29147,N_28476,N_28791);
xor U29148 (N_29148,N_28213,N_28572);
and U29149 (N_29149,N_28315,N_28507);
nor U29150 (N_29150,N_28415,N_28424);
xor U29151 (N_29151,N_28709,N_28291);
xnor U29152 (N_29152,N_28736,N_28379);
or U29153 (N_29153,N_28235,N_28724);
or U29154 (N_29154,N_28687,N_28540);
and U29155 (N_29155,N_28532,N_28727);
xor U29156 (N_29156,N_28418,N_28411);
nand U29157 (N_29157,N_28543,N_28459);
nor U29158 (N_29158,N_28231,N_28203);
and U29159 (N_29159,N_28242,N_28576);
or U29160 (N_29160,N_28420,N_28236);
nand U29161 (N_29161,N_28322,N_28481);
xor U29162 (N_29162,N_28403,N_28792);
nand U29163 (N_29163,N_28221,N_28784);
xnor U29164 (N_29164,N_28346,N_28568);
or U29165 (N_29165,N_28744,N_28316);
xor U29166 (N_29166,N_28764,N_28684);
or U29167 (N_29167,N_28508,N_28545);
and U29168 (N_29168,N_28647,N_28419);
nand U29169 (N_29169,N_28309,N_28641);
nand U29170 (N_29170,N_28394,N_28501);
xor U29171 (N_29171,N_28569,N_28457);
or U29172 (N_29172,N_28767,N_28298);
and U29173 (N_29173,N_28664,N_28728);
or U29174 (N_29174,N_28662,N_28244);
and U29175 (N_29175,N_28467,N_28582);
nor U29176 (N_29176,N_28674,N_28618);
nand U29177 (N_29177,N_28525,N_28638);
nor U29178 (N_29178,N_28302,N_28660);
nor U29179 (N_29179,N_28681,N_28326);
and U29180 (N_29180,N_28487,N_28668);
nand U29181 (N_29181,N_28451,N_28495);
and U29182 (N_29182,N_28470,N_28322);
nand U29183 (N_29183,N_28441,N_28355);
or U29184 (N_29184,N_28512,N_28769);
or U29185 (N_29185,N_28324,N_28347);
and U29186 (N_29186,N_28299,N_28652);
and U29187 (N_29187,N_28597,N_28782);
or U29188 (N_29188,N_28382,N_28246);
or U29189 (N_29189,N_28592,N_28566);
or U29190 (N_29190,N_28385,N_28245);
nor U29191 (N_29191,N_28569,N_28436);
and U29192 (N_29192,N_28527,N_28463);
nor U29193 (N_29193,N_28712,N_28562);
nand U29194 (N_29194,N_28660,N_28680);
nor U29195 (N_29195,N_28513,N_28501);
and U29196 (N_29196,N_28798,N_28506);
and U29197 (N_29197,N_28350,N_28698);
nand U29198 (N_29198,N_28744,N_28605);
or U29199 (N_29199,N_28458,N_28748);
or U29200 (N_29200,N_28529,N_28574);
xnor U29201 (N_29201,N_28310,N_28536);
and U29202 (N_29202,N_28403,N_28724);
or U29203 (N_29203,N_28609,N_28388);
nor U29204 (N_29204,N_28510,N_28779);
nand U29205 (N_29205,N_28305,N_28527);
nand U29206 (N_29206,N_28259,N_28338);
nand U29207 (N_29207,N_28688,N_28292);
and U29208 (N_29208,N_28422,N_28720);
nor U29209 (N_29209,N_28509,N_28568);
and U29210 (N_29210,N_28260,N_28737);
and U29211 (N_29211,N_28479,N_28278);
and U29212 (N_29212,N_28661,N_28449);
nand U29213 (N_29213,N_28492,N_28581);
xnor U29214 (N_29214,N_28786,N_28481);
nor U29215 (N_29215,N_28762,N_28336);
and U29216 (N_29216,N_28484,N_28645);
nor U29217 (N_29217,N_28555,N_28556);
xnor U29218 (N_29218,N_28455,N_28702);
or U29219 (N_29219,N_28513,N_28369);
or U29220 (N_29220,N_28315,N_28240);
or U29221 (N_29221,N_28452,N_28226);
nand U29222 (N_29222,N_28683,N_28279);
xnor U29223 (N_29223,N_28436,N_28624);
and U29224 (N_29224,N_28715,N_28680);
xnor U29225 (N_29225,N_28546,N_28390);
or U29226 (N_29226,N_28742,N_28451);
nand U29227 (N_29227,N_28603,N_28674);
nor U29228 (N_29228,N_28371,N_28441);
or U29229 (N_29229,N_28226,N_28577);
nor U29230 (N_29230,N_28630,N_28596);
and U29231 (N_29231,N_28565,N_28204);
and U29232 (N_29232,N_28757,N_28403);
or U29233 (N_29233,N_28699,N_28264);
xor U29234 (N_29234,N_28425,N_28599);
nor U29235 (N_29235,N_28247,N_28779);
xor U29236 (N_29236,N_28392,N_28498);
or U29237 (N_29237,N_28471,N_28360);
nand U29238 (N_29238,N_28637,N_28663);
nand U29239 (N_29239,N_28282,N_28524);
xor U29240 (N_29240,N_28750,N_28553);
xor U29241 (N_29241,N_28356,N_28794);
and U29242 (N_29242,N_28657,N_28541);
or U29243 (N_29243,N_28515,N_28209);
nand U29244 (N_29244,N_28504,N_28463);
xnor U29245 (N_29245,N_28315,N_28753);
or U29246 (N_29246,N_28785,N_28363);
or U29247 (N_29247,N_28356,N_28439);
nand U29248 (N_29248,N_28613,N_28243);
or U29249 (N_29249,N_28458,N_28417);
nand U29250 (N_29250,N_28609,N_28641);
nor U29251 (N_29251,N_28283,N_28604);
and U29252 (N_29252,N_28294,N_28494);
nor U29253 (N_29253,N_28441,N_28543);
or U29254 (N_29254,N_28648,N_28604);
nand U29255 (N_29255,N_28221,N_28236);
nor U29256 (N_29256,N_28334,N_28529);
xor U29257 (N_29257,N_28713,N_28674);
and U29258 (N_29258,N_28793,N_28451);
nor U29259 (N_29259,N_28690,N_28653);
nor U29260 (N_29260,N_28338,N_28375);
and U29261 (N_29261,N_28691,N_28693);
and U29262 (N_29262,N_28506,N_28610);
or U29263 (N_29263,N_28437,N_28475);
and U29264 (N_29264,N_28462,N_28314);
or U29265 (N_29265,N_28415,N_28258);
xor U29266 (N_29266,N_28241,N_28478);
xnor U29267 (N_29267,N_28597,N_28533);
and U29268 (N_29268,N_28537,N_28657);
nand U29269 (N_29269,N_28627,N_28301);
nand U29270 (N_29270,N_28643,N_28653);
and U29271 (N_29271,N_28414,N_28372);
nor U29272 (N_29272,N_28484,N_28554);
nand U29273 (N_29273,N_28632,N_28700);
or U29274 (N_29274,N_28564,N_28539);
nand U29275 (N_29275,N_28369,N_28609);
nand U29276 (N_29276,N_28373,N_28482);
xnor U29277 (N_29277,N_28308,N_28696);
or U29278 (N_29278,N_28280,N_28692);
xnor U29279 (N_29279,N_28696,N_28239);
and U29280 (N_29280,N_28793,N_28584);
or U29281 (N_29281,N_28329,N_28202);
nand U29282 (N_29282,N_28277,N_28362);
xor U29283 (N_29283,N_28353,N_28253);
nor U29284 (N_29284,N_28753,N_28469);
nor U29285 (N_29285,N_28313,N_28424);
nand U29286 (N_29286,N_28535,N_28384);
xor U29287 (N_29287,N_28260,N_28679);
and U29288 (N_29288,N_28578,N_28328);
or U29289 (N_29289,N_28604,N_28441);
and U29290 (N_29290,N_28694,N_28716);
nor U29291 (N_29291,N_28653,N_28446);
nor U29292 (N_29292,N_28381,N_28274);
nor U29293 (N_29293,N_28356,N_28778);
or U29294 (N_29294,N_28729,N_28271);
or U29295 (N_29295,N_28222,N_28352);
or U29296 (N_29296,N_28414,N_28201);
nand U29297 (N_29297,N_28482,N_28412);
and U29298 (N_29298,N_28642,N_28686);
nor U29299 (N_29299,N_28329,N_28204);
nand U29300 (N_29300,N_28632,N_28593);
nand U29301 (N_29301,N_28305,N_28592);
xor U29302 (N_29302,N_28657,N_28697);
nor U29303 (N_29303,N_28704,N_28500);
xor U29304 (N_29304,N_28264,N_28245);
xnor U29305 (N_29305,N_28467,N_28346);
nand U29306 (N_29306,N_28395,N_28478);
and U29307 (N_29307,N_28794,N_28517);
nor U29308 (N_29308,N_28478,N_28570);
or U29309 (N_29309,N_28675,N_28369);
nor U29310 (N_29310,N_28631,N_28311);
xnor U29311 (N_29311,N_28433,N_28689);
and U29312 (N_29312,N_28338,N_28699);
nand U29313 (N_29313,N_28419,N_28356);
nand U29314 (N_29314,N_28679,N_28522);
or U29315 (N_29315,N_28672,N_28665);
xor U29316 (N_29316,N_28246,N_28309);
xor U29317 (N_29317,N_28606,N_28353);
or U29318 (N_29318,N_28428,N_28245);
or U29319 (N_29319,N_28569,N_28437);
nor U29320 (N_29320,N_28217,N_28263);
xnor U29321 (N_29321,N_28767,N_28258);
nor U29322 (N_29322,N_28270,N_28454);
xnor U29323 (N_29323,N_28251,N_28451);
or U29324 (N_29324,N_28795,N_28562);
and U29325 (N_29325,N_28647,N_28659);
and U29326 (N_29326,N_28213,N_28331);
xnor U29327 (N_29327,N_28417,N_28572);
and U29328 (N_29328,N_28595,N_28225);
nand U29329 (N_29329,N_28595,N_28608);
nand U29330 (N_29330,N_28600,N_28338);
nand U29331 (N_29331,N_28545,N_28275);
and U29332 (N_29332,N_28278,N_28568);
and U29333 (N_29333,N_28724,N_28634);
xor U29334 (N_29334,N_28658,N_28450);
nand U29335 (N_29335,N_28778,N_28529);
nor U29336 (N_29336,N_28753,N_28277);
xnor U29337 (N_29337,N_28512,N_28754);
nand U29338 (N_29338,N_28432,N_28250);
xor U29339 (N_29339,N_28628,N_28648);
xnor U29340 (N_29340,N_28781,N_28689);
xnor U29341 (N_29341,N_28434,N_28432);
or U29342 (N_29342,N_28735,N_28769);
xor U29343 (N_29343,N_28402,N_28734);
xnor U29344 (N_29344,N_28647,N_28277);
xnor U29345 (N_29345,N_28432,N_28403);
or U29346 (N_29346,N_28583,N_28643);
nand U29347 (N_29347,N_28450,N_28267);
or U29348 (N_29348,N_28702,N_28388);
nor U29349 (N_29349,N_28462,N_28407);
nand U29350 (N_29350,N_28230,N_28543);
or U29351 (N_29351,N_28612,N_28594);
nand U29352 (N_29352,N_28431,N_28393);
nand U29353 (N_29353,N_28352,N_28782);
and U29354 (N_29354,N_28237,N_28207);
nand U29355 (N_29355,N_28758,N_28784);
or U29356 (N_29356,N_28407,N_28552);
xor U29357 (N_29357,N_28643,N_28270);
nor U29358 (N_29358,N_28302,N_28376);
nor U29359 (N_29359,N_28479,N_28297);
or U29360 (N_29360,N_28475,N_28385);
and U29361 (N_29361,N_28388,N_28264);
nand U29362 (N_29362,N_28549,N_28712);
xor U29363 (N_29363,N_28595,N_28665);
xnor U29364 (N_29364,N_28409,N_28629);
nor U29365 (N_29365,N_28438,N_28491);
nand U29366 (N_29366,N_28303,N_28521);
nand U29367 (N_29367,N_28226,N_28620);
and U29368 (N_29368,N_28484,N_28378);
xor U29369 (N_29369,N_28514,N_28642);
nor U29370 (N_29370,N_28489,N_28561);
nor U29371 (N_29371,N_28599,N_28753);
nor U29372 (N_29372,N_28483,N_28316);
xnor U29373 (N_29373,N_28540,N_28586);
xnor U29374 (N_29374,N_28323,N_28674);
and U29375 (N_29375,N_28427,N_28580);
nand U29376 (N_29376,N_28794,N_28432);
or U29377 (N_29377,N_28704,N_28437);
or U29378 (N_29378,N_28634,N_28292);
nor U29379 (N_29379,N_28698,N_28542);
and U29380 (N_29380,N_28729,N_28534);
and U29381 (N_29381,N_28568,N_28218);
xor U29382 (N_29382,N_28368,N_28675);
xor U29383 (N_29383,N_28662,N_28680);
nor U29384 (N_29384,N_28409,N_28399);
xor U29385 (N_29385,N_28498,N_28627);
nor U29386 (N_29386,N_28451,N_28593);
nor U29387 (N_29387,N_28327,N_28500);
or U29388 (N_29388,N_28223,N_28552);
xor U29389 (N_29389,N_28479,N_28215);
and U29390 (N_29390,N_28201,N_28650);
or U29391 (N_29391,N_28610,N_28238);
and U29392 (N_29392,N_28319,N_28210);
nand U29393 (N_29393,N_28661,N_28467);
nand U29394 (N_29394,N_28246,N_28284);
or U29395 (N_29395,N_28390,N_28438);
xnor U29396 (N_29396,N_28603,N_28544);
xnor U29397 (N_29397,N_28254,N_28259);
nor U29398 (N_29398,N_28529,N_28799);
xor U29399 (N_29399,N_28737,N_28531);
nand U29400 (N_29400,N_29110,N_29123);
and U29401 (N_29401,N_28848,N_29296);
and U29402 (N_29402,N_29099,N_29298);
and U29403 (N_29403,N_29030,N_29297);
and U29404 (N_29404,N_29245,N_29368);
nor U29405 (N_29405,N_28804,N_29131);
or U29406 (N_29406,N_29201,N_28948);
xor U29407 (N_29407,N_28806,N_29086);
or U29408 (N_29408,N_28920,N_28902);
nand U29409 (N_29409,N_29292,N_28976);
or U29410 (N_29410,N_29170,N_29080);
nand U29411 (N_29411,N_29087,N_29209);
and U29412 (N_29412,N_29204,N_29098);
nand U29413 (N_29413,N_28901,N_28905);
nand U29414 (N_29414,N_29338,N_29067);
nor U29415 (N_29415,N_28864,N_29358);
and U29416 (N_29416,N_29044,N_29304);
or U29417 (N_29417,N_29130,N_28906);
and U29418 (N_29418,N_29257,N_28816);
xor U29419 (N_29419,N_28968,N_29140);
and U29420 (N_29420,N_29236,N_29356);
and U29421 (N_29421,N_29047,N_28965);
and U29422 (N_29422,N_28904,N_28871);
nor U29423 (N_29423,N_29395,N_29271);
nor U29424 (N_29424,N_28865,N_29061);
and U29425 (N_29425,N_28808,N_29021);
xor U29426 (N_29426,N_29185,N_29012);
xor U29427 (N_29427,N_28837,N_28887);
and U29428 (N_29428,N_28999,N_29128);
xnor U29429 (N_29429,N_29006,N_29325);
nor U29430 (N_29430,N_29235,N_29380);
xor U29431 (N_29431,N_29238,N_29057);
xnor U29432 (N_29432,N_28841,N_29393);
nor U29433 (N_29433,N_28981,N_28891);
and U29434 (N_29434,N_29052,N_28972);
or U29435 (N_29435,N_28859,N_28953);
or U29436 (N_29436,N_29142,N_29295);
or U29437 (N_29437,N_29253,N_29303);
nor U29438 (N_29438,N_29028,N_28979);
or U29439 (N_29439,N_29008,N_29045);
or U29440 (N_29440,N_28938,N_29068);
nor U29441 (N_29441,N_28944,N_28923);
or U29442 (N_29442,N_28880,N_28826);
or U29443 (N_29443,N_29120,N_28955);
xor U29444 (N_29444,N_29191,N_28984);
nand U29445 (N_29445,N_29166,N_29314);
xnor U29446 (N_29446,N_28827,N_29063);
and U29447 (N_29447,N_29171,N_29137);
and U29448 (N_29448,N_28819,N_29102);
nand U29449 (N_29449,N_29108,N_28863);
or U29450 (N_29450,N_29095,N_28980);
nor U29451 (N_29451,N_28959,N_28829);
nor U29452 (N_29452,N_28861,N_28843);
or U29453 (N_29453,N_28978,N_29058);
xnor U29454 (N_29454,N_29059,N_29233);
nor U29455 (N_29455,N_29306,N_29225);
nand U29456 (N_29456,N_29211,N_29266);
xnor U29457 (N_29457,N_29139,N_28877);
and U29458 (N_29458,N_29391,N_29039);
and U29459 (N_29459,N_28846,N_29144);
nor U29460 (N_29460,N_29373,N_28860);
nor U29461 (N_29461,N_29180,N_29291);
or U29462 (N_29462,N_29312,N_28915);
and U29463 (N_29463,N_29136,N_29256);
nand U29464 (N_29464,N_29398,N_29165);
nand U29465 (N_29465,N_29284,N_29268);
xnor U29466 (N_29466,N_28935,N_29188);
nand U29467 (N_29467,N_28857,N_29060);
or U29468 (N_29468,N_28815,N_29074);
nand U29469 (N_29469,N_29392,N_28987);
or U29470 (N_29470,N_29056,N_29357);
xor U29471 (N_29471,N_29249,N_29153);
nand U29472 (N_29472,N_29133,N_28921);
nand U29473 (N_29473,N_29109,N_29082);
xor U29474 (N_29474,N_29277,N_28872);
or U29475 (N_29475,N_29182,N_29365);
or U29476 (N_29476,N_29138,N_28890);
xor U29477 (N_29477,N_29332,N_29203);
or U29478 (N_29478,N_29263,N_28867);
or U29479 (N_29479,N_29145,N_28844);
xnor U29480 (N_29480,N_29319,N_29321);
and U29481 (N_29481,N_29343,N_28840);
xor U29482 (N_29482,N_29169,N_29024);
or U29483 (N_29483,N_29383,N_28991);
nand U29484 (N_29484,N_28961,N_29017);
or U29485 (N_29485,N_29230,N_28866);
and U29486 (N_29486,N_28936,N_28943);
or U29487 (N_29487,N_29183,N_29157);
or U29488 (N_29488,N_29324,N_28810);
or U29489 (N_29489,N_28894,N_28822);
xor U29490 (N_29490,N_29156,N_29200);
or U29491 (N_29491,N_29223,N_29290);
or U29492 (N_29492,N_29029,N_29009);
nor U29493 (N_29493,N_28913,N_28853);
xnor U29494 (N_29494,N_29122,N_29041);
or U29495 (N_29495,N_29375,N_28952);
nor U29496 (N_29496,N_29261,N_29175);
and U29497 (N_29497,N_29388,N_29331);
nand U29498 (N_29498,N_28962,N_29001);
or U29499 (N_29499,N_29033,N_29300);
nand U29500 (N_29500,N_29196,N_29042);
or U29501 (N_29501,N_28832,N_29349);
and U29502 (N_29502,N_29119,N_28946);
and U29503 (N_29503,N_28849,N_29330);
nor U29504 (N_29504,N_29112,N_29316);
and U29505 (N_29505,N_29107,N_29281);
or U29506 (N_29506,N_29382,N_28812);
xor U29507 (N_29507,N_29282,N_29014);
nand U29508 (N_29508,N_29081,N_28818);
or U29509 (N_29509,N_29089,N_29333);
nand U29510 (N_29510,N_29083,N_29232);
nor U29511 (N_29511,N_29315,N_29305);
or U29512 (N_29512,N_28879,N_28817);
and U29513 (N_29513,N_28856,N_29317);
xnor U29514 (N_29514,N_29226,N_29097);
nand U29515 (N_29515,N_29072,N_29342);
nor U29516 (N_29516,N_29092,N_29351);
and U29517 (N_29517,N_29376,N_29251);
nand U29518 (N_29518,N_29397,N_29246);
and U29519 (N_29519,N_29101,N_29287);
nand U29520 (N_29520,N_29124,N_28949);
or U29521 (N_29521,N_29354,N_29346);
nor U29522 (N_29522,N_29371,N_28967);
nand U29523 (N_29523,N_29259,N_29071);
nor U29524 (N_29524,N_29055,N_28855);
or U29525 (N_29525,N_29250,N_28800);
nand U29526 (N_29526,N_28995,N_28996);
or U29527 (N_29527,N_29301,N_28868);
nand U29528 (N_29528,N_29005,N_29270);
nand U29529 (N_29529,N_29218,N_29224);
xnor U29530 (N_29530,N_29255,N_28809);
and U29531 (N_29531,N_28954,N_29036);
and U29532 (N_29532,N_29004,N_29289);
nand U29533 (N_29533,N_29049,N_29173);
or U29534 (N_29534,N_29276,N_28807);
or U29535 (N_29535,N_28912,N_28825);
nand U29536 (N_29536,N_29073,N_29384);
xnor U29537 (N_29537,N_29066,N_28966);
xor U29538 (N_29538,N_29031,N_29229);
nor U29539 (N_29539,N_29025,N_29372);
nor U29540 (N_29540,N_29146,N_28886);
and U29541 (N_29541,N_29339,N_29105);
or U29542 (N_29542,N_29126,N_29329);
nor U29543 (N_29543,N_29378,N_29274);
or U29544 (N_29544,N_28934,N_29077);
nor U29545 (N_29545,N_28878,N_29093);
xor U29546 (N_29546,N_29396,N_29186);
and U29547 (N_29547,N_28895,N_29187);
nor U29548 (N_29548,N_29007,N_29335);
and U29549 (N_29549,N_29337,N_29248);
nand U29550 (N_29550,N_28884,N_28924);
or U29551 (N_29551,N_29189,N_28942);
nand U29552 (N_29552,N_28925,N_28903);
nor U29553 (N_29553,N_28830,N_29264);
nor U29554 (N_29554,N_29190,N_29205);
xnor U29555 (N_29555,N_29283,N_29090);
nand U29556 (N_29556,N_29159,N_29370);
nor U29557 (N_29557,N_29269,N_29158);
xor U29558 (N_29558,N_29194,N_29010);
nand U29559 (N_29559,N_28852,N_29070);
or U29560 (N_29560,N_29364,N_29034);
xnor U29561 (N_29561,N_28892,N_28882);
xnor U29562 (N_29562,N_28986,N_28919);
or U29563 (N_29563,N_28824,N_29336);
or U29564 (N_29564,N_28910,N_29216);
xnor U29565 (N_29565,N_28811,N_29309);
nor U29566 (N_29566,N_29000,N_29374);
nor U29567 (N_29567,N_28963,N_29275);
nor U29568 (N_29568,N_28951,N_28833);
xnor U29569 (N_29569,N_29195,N_28922);
nor U29570 (N_29570,N_28940,N_29177);
nand U29571 (N_29571,N_28989,N_28862);
or U29572 (N_29572,N_29091,N_29192);
xnor U29573 (N_29573,N_29132,N_28881);
and U29574 (N_29574,N_29310,N_29207);
or U29575 (N_29575,N_29286,N_28939);
nand U29576 (N_29576,N_29019,N_29143);
and U29577 (N_29577,N_28813,N_29085);
nor U29578 (N_29578,N_29273,N_29328);
xnor U29579 (N_29579,N_29125,N_29168);
or U29580 (N_29580,N_29212,N_29234);
and U29581 (N_29581,N_29172,N_28874);
xor U29582 (N_29582,N_28997,N_29228);
and U29583 (N_29583,N_28900,N_29043);
xor U29584 (N_29584,N_29299,N_29242);
nor U29585 (N_29585,N_28831,N_29272);
nand U29586 (N_29586,N_29096,N_29178);
nor U29587 (N_29587,N_29320,N_29239);
nand U29588 (N_29588,N_29174,N_28932);
nor U29589 (N_29589,N_29053,N_28928);
nand U29590 (N_29590,N_29064,N_29240);
or U29591 (N_29591,N_29149,N_29241);
or U29592 (N_29592,N_29114,N_29160);
nand U29593 (N_29593,N_28985,N_29147);
nand U29594 (N_29594,N_29161,N_29322);
xnor U29595 (N_29595,N_28916,N_29244);
nand U29596 (N_29596,N_28893,N_28970);
xnor U29597 (N_29597,N_29046,N_29237);
and U29598 (N_29598,N_29345,N_28836);
and U29599 (N_29599,N_28911,N_28918);
nor U29600 (N_29600,N_29113,N_28909);
nor U29601 (N_29601,N_28931,N_29214);
and U29602 (N_29602,N_29152,N_29386);
or U29603 (N_29603,N_28982,N_28998);
nor U29604 (N_29604,N_29037,N_29103);
nand U29605 (N_29605,N_29381,N_29260);
or U29606 (N_29606,N_29258,N_29134);
nand U29607 (N_29607,N_28888,N_28956);
nor U29608 (N_29608,N_29387,N_29106);
and U29609 (N_29609,N_28896,N_28838);
xor U29610 (N_29610,N_29088,N_28941);
and U29611 (N_29611,N_28801,N_29334);
xnor U29612 (N_29612,N_28828,N_29350);
nor U29613 (N_29613,N_28823,N_29385);
xor U29614 (N_29614,N_28834,N_28845);
and U29615 (N_29615,N_29323,N_28803);
and U29616 (N_29616,N_29111,N_29279);
and U29617 (N_29617,N_29293,N_28858);
or U29618 (N_29618,N_29075,N_28847);
or U29619 (N_29619,N_29394,N_28958);
nand U29620 (N_29620,N_29078,N_29361);
xor U29621 (N_29621,N_28937,N_28917);
nand U29622 (N_29622,N_28875,N_29151);
nor U29623 (N_29623,N_29227,N_29231);
nand U29624 (N_29624,N_29018,N_29206);
or U29625 (N_29625,N_29288,N_29176);
or U29626 (N_29626,N_29362,N_29117);
or U29627 (N_29627,N_29220,N_29366);
nor U29628 (N_29628,N_29094,N_29184);
nand U29629 (N_29629,N_29352,N_29210);
nand U29630 (N_29630,N_29127,N_29208);
nor U29631 (N_29631,N_28820,N_28850);
xor U29632 (N_29632,N_29154,N_29353);
nor U29633 (N_29633,N_29141,N_28992);
nor U29634 (N_29634,N_28908,N_29032);
xnor U29635 (N_29635,N_28930,N_28945);
xnor U29636 (N_29636,N_29359,N_29222);
nor U29637 (N_29637,N_28805,N_29026);
nor U29638 (N_29638,N_29003,N_29079);
nand U29639 (N_29639,N_29217,N_29015);
xor U29640 (N_29640,N_28814,N_28873);
nand U29641 (N_29641,N_29318,N_29023);
nand U29642 (N_29642,N_29104,N_29162);
and U29643 (N_29643,N_29307,N_29002);
and U29644 (N_29644,N_28876,N_29344);
and U29645 (N_29645,N_28974,N_28957);
or U29646 (N_29646,N_29311,N_28914);
nor U29647 (N_29647,N_28869,N_28854);
nor U29648 (N_29648,N_29115,N_29129);
xor U29649 (N_29649,N_29198,N_28802);
or U29650 (N_29650,N_28933,N_29065);
and U29651 (N_29651,N_28835,N_28947);
and U29652 (N_29652,N_29116,N_28950);
or U29653 (N_29653,N_28851,N_28990);
xnor U29654 (N_29654,N_29181,N_28993);
nand U29655 (N_29655,N_29084,N_29179);
nand U29656 (N_29656,N_28975,N_29118);
xnor U29657 (N_29657,N_29377,N_29197);
xor U29658 (N_29658,N_29262,N_29050);
and U29659 (N_29659,N_29265,N_28977);
and U29660 (N_29660,N_29011,N_29252);
nor U29661 (N_29661,N_29150,N_29360);
or U29662 (N_29662,N_29100,N_28994);
and U29663 (N_29663,N_28883,N_28821);
or U29664 (N_29664,N_29035,N_29294);
nor U29665 (N_29665,N_28897,N_29348);
xnor U29666 (N_29666,N_29221,N_29193);
xnor U29667 (N_29667,N_28842,N_29163);
nor U29668 (N_29668,N_29254,N_28870);
and U29669 (N_29669,N_28889,N_29062);
xor U29670 (N_29670,N_29038,N_29135);
xor U29671 (N_29671,N_29013,N_29347);
and U29672 (N_29672,N_29247,N_29327);
xnor U29673 (N_29673,N_28839,N_29363);
and U29674 (N_29674,N_28929,N_28988);
or U29675 (N_29675,N_28983,N_29355);
and U29676 (N_29676,N_29040,N_29076);
or U29677 (N_29677,N_29148,N_29369);
nor U29678 (N_29678,N_29399,N_29367);
or U29679 (N_29679,N_29313,N_28885);
nand U29680 (N_29680,N_29164,N_28898);
or U29681 (N_29681,N_29308,N_28926);
nand U29682 (N_29682,N_29280,N_28927);
xor U29683 (N_29683,N_29390,N_29016);
or U29684 (N_29684,N_29267,N_29167);
nand U29685 (N_29685,N_29048,N_29389);
nor U29686 (N_29686,N_29219,N_29215);
nor U29687 (N_29687,N_29278,N_29243);
nor U29688 (N_29688,N_29051,N_29027);
nor U29689 (N_29689,N_29022,N_29155);
and U29690 (N_29690,N_28960,N_29341);
xor U29691 (N_29691,N_28971,N_29326);
nor U29692 (N_29692,N_29302,N_28973);
xor U29693 (N_29693,N_29340,N_29202);
xor U29694 (N_29694,N_28907,N_29285);
nand U29695 (N_29695,N_29199,N_29121);
nand U29696 (N_29696,N_28899,N_28969);
nand U29697 (N_29697,N_29213,N_29020);
xnor U29698 (N_29698,N_28964,N_29054);
xnor U29699 (N_29699,N_29069,N_29379);
or U29700 (N_29700,N_29069,N_28830);
and U29701 (N_29701,N_29313,N_29106);
and U29702 (N_29702,N_29363,N_29253);
and U29703 (N_29703,N_29056,N_29004);
nand U29704 (N_29704,N_29066,N_28847);
nor U29705 (N_29705,N_29072,N_29164);
nor U29706 (N_29706,N_28996,N_29184);
xnor U29707 (N_29707,N_28994,N_28877);
nor U29708 (N_29708,N_29040,N_28865);
and U29709 (N_29709,N_29121,N_29313);
or U29710 (N_29710,N_29188,N_28947);
nor U29711 (N_29711,N_29184,N_29296);
nor U29712 (N_29712,N_28948,N_29316);
or U29713 (N_29713,N_28823,N_29216);
xor U29714 (N_29714,N_29371,N_29087);
xnor U29715 (N_29715,N_28830,N_28913);
nand U29716 (N_29716,N_29336,N_29003);
nor U29717 (N_29717,N_29045,N_28834);
and U29718 (N_29718,N_29000,N_29059);
nand U29719 (N_29719,N_29126,N_29339);
or U29720 (N_29720,N_29231,N_29320);
or U29721 (N_29721,N_28902,N_29012);
nand U29722 (N_29722,N_29097,N_28868);
xnor U29723 (N_29723,N_29393,N_29248);
nor U29724 (N_29724,N_28903,N_28808);
xnor U29725 (N_29725,N_29082,N_28801);
xor U29726 (N_29726,N_28925,N_28866);
nand U29727 (N_29727,N_29012,N_29211);
or U29728 (N_29728,N_29033,N_28896);
nand U29729 (N_29729,N_29397,N_28821);
xnor U29730 (N_29730,N_29225,N_29222);
or U29731 (N_29731,N_29135,N_28959);
nand U29732 (N_29732,N_29032,N_28926);
or U29733 (N_29733,N_29207,N_29086);
nor U29734 (N_29734,N_28857,N_29328);
or U29735 (N_29735,N_29068,N_29327);
or U29736 (N_29736,N_29267,N_29114);
xnor U29737 (N_29737,N_29068,N_29112);
xor U29738 (N_29738,N_28804,N_29374);
and U29739 (N_29739,N_29065,N_29172);
xnor U29740 (N_29740,N_29098,N_28991);
or U29741 (N_29741,N_29133,N_29242);
and U29742 (N_29742,N_28932,N_28891);
xor U29743 (N_29743,N_28923,N_29061);
and U29744 (N_29744,N_28810,N_28928);
and U29745 (N_29745,N_29057,N_29069);
xor U29746 (N_29746,N_28842,N_29109);
or U29747 (N_29747,N_29137,N_28811);
and U29748 (N_29748,N_29085,N_29019);
or U29749 (N_29749,N_29315,N_28870);
nand U29750 (N_29750,N_29160,N_29193);
and U29751 (N_29751,N_29385,N_29383);
or U29752 (N_29752,N_29092,N_29090);
or U29753 (N_29753,N_29311,N_28936);
nand U29754 (N_29754,N_29186,N_28913);
nand U29755 (N_29755,N_28956,N_29030);
or U29756 (N_29756,N_28869,N_29316);
nand U29757 (N_29757,N_29063,N_29201);
xnor U29758 (N_29758,N_28877,N_28860);
xor U29759 (N_29759,N_28901,N_29090);
and U29760 (N_29760,N_29003,N_29392);
nor U29761 (N_29761,N_29273,N_29224);
xor U29762 (N_29762,N_29049,N_29256);
xor U29763 (N_29763,N_29186,N_28951);
nand U29764 (N_29764,N_29105,N_29353);
nand U29765 (N_29765,N_29251,N_28893);
nor U29766 (N_29766,N_29251,N_29146);
or U29767 (N_29767,N_29208,N_29189);
and U29768 (N_29768,N_29283,N_29271);
and U29769 (N_29769,N_28972,N_29001);
xnor U29770 (N_29770,N_29380,N_28831);
nor U29771 (N_29771,N_28939,N_29272);
xnor U29772 (N_29772,N_28871,N_29201);
nor U29773 (N_29773,N_28922,N_29185);
and U29774 (N_29774,N_29388,N_29232);
nor U29775 (N_29775,N_29012,N_29370);
nand U29776 (N_29776,N_29046,N_29206);
xor U29777 (N_29777,N_29004,N_29173);
or U29778 (N_29778,N_28922,N_28985);
nand U29779 (N_29779,N_29318,N_28967);
nand U29780 (N_29780,N_29240,N_29269);
nand U29781 (N_29781,N_29154,N_29230);
and U29782 (N_29782,N_28819,N_29305);
nor U29783 (N_29783,N_29314,N_29056);
xnor U29784 (N_29784,N_28928,N_28955);
nand U29785 (N_29785,N_29293,N_29097);
and U29786 (N_29786,N_29029,N_28874);
nand U29787 (N_29787,N_29091,N_29145);
nand U29788 (N_29788,N_29329,N_28977);
nor U29789 (N_29789,N_29019,N_29051);
nand U29790 (N_29790,N_29195,N_29014);
xor U29791 (N_29791,N_29023,N_28823);
xnor U29792 (N_29792,N_28865,N_29101);
nor U29793 (N_29793,N_29306,N_28937);
nand U29794 (N_29794,N_28989,N_28917);
nand U29795 (N_29795,N_29178,N_28870);
nand U29796 (N_29796,N_28927,N_28942);
and U29797 (N_29797,N_28921,N_29336);
nor U29798 (N_29798,N_29240,N_29394);
xnor U29799 (N_29799,N_29257,N_28845);
nand U29800 (N_29800,N_29120,N_29175);
nand U29801 (N_29801,N_29313,N_28974);
nor U29802 (N_29802,N_28851,N_28975);
xnor U29803 (N_29803,N_28855,N_29275);
nand U29804 (N_29804,N_28871,N_28954);
nor U29805 (N_29805,N_29233,N_29370);
and U29806 (N_29806,N_29026,N_29134);
and U29807 (N_29807,N_28996,N_29135);
nor U29808 (N_29808,N_29078,N_28831);
nand U29809 (N_29809,N_29206,N_28903);
nor U29810 (N_29810,N_29399,N_29268);
nand U29811 (N_29811,N_29294,N_29306);
nor U29812 (N_29812,N_29251,N_28855);
xnor U29813 (N_29813,N_28840,N_28924);
and U29814 (N_29814,N_28803,N_29270);
or U29815 (N_29815,N_29252,N_28970);
nor U29816 (N_29816,N_28976,N_29100);
and U29817 (N_29817,N_28855,N_28857);
xnor U29818 (N_29818,N_29333,N_28890);
nor U29819 (N_29819,N_29204,N_29340);
nand U29820 (N_29820,N_29103,N_28842);
nand U29821 (N_29821,N_28815,N_29002);
nor U29822 (N_29822,N_29024,N_29080);
nand U29823 (N_29823,N_29146,N_28924);
nor U29824 (N_29824,N_29126,N_29112);
nand U29825 (N_29825,N_28899,N_28954);
nand U29826 (N_29826,N_28935,N_28966);
xnor U29827 (N_29827,N_29338,N_29255);
nand U29828 (N_29828,N_29109,N_28808);
and U29829 (N_29829,N_29060,N_28975);
xor U29830 (N_29830,N_28954,N_29313);
nor U29831 (N_29831,N_29358,N_28874);
or U29832 (N_29832,N_28933,N_29226);
nor U29833 (N_29833,N_29043,N_29251);
and U29834 (N_29834,N_29180,N_29189);
nand U29835 (N_29835,N_29099,N_28810);
nand U29836 (N_29836,N_28976,N_28820);
xnor U29837 (N_29837,N_28939,N_29269);
nand U29838 (N_29838,N_28999,N_29361);
and U29839 (N_29839,N_28824,N_28817);
or U29840 (N_29840,N_29057,N_29343);
nor U29841 (N_29841,N_28961,N_28823);
nand U29842 (N_29842,N_29275,N_29139);
nor U29843 (N_29843,N_28910,N_29185);
nand U29844 (N_29844,N_29265,N_29354);
xnor U29845 (N_29845,N_29269,N_29387);
xnor U29846 (N_29846,N_29018,N_28985);
nand U29847 (N_29847,N_29370,N_29148);
nor U29848 (N_29848,N_29205,N_29152);
or U29849 (N_29849,N_29020,N_29100);
nor U29850 (N_29850,N_28881,N_29255);
nand U29851 (N_29851,N_29260,N_29184);
nand U29852 (N_29852,N_29113,N_28925);
nand U29853 (N_29853,N_29396,N_29397);
nand U29854 (N_29854,N_29135,N_29216);
nand U29855 (N_29855,N_29297,N_29000);
or U29856 (N_29856,N_29324,N_29122);
and U29857 (N_29857,N_28988,N_29196);
xor U29858 (N_29858,N_29106,N_29062);
nor U29859 (N_29859,N_29060,N_29126);
nand U29860 (N_29860,N_29020,N_29018);
xor U29861 (N_29861,N_29112,N_28951);
nand U29862 (N_29862,N_28960,N_28980);
xnor U29863 (N_29863,N_28880,N_29225);
and U29864 (N_29864,N_29041,N_29172);
nor U29865 (N_29865,N_28859,N_28962);
and U29866 (N_29866,N_29192,N_29399);
and U29867 (N_29867,N_29023,N_28845);
or U29868 (N_29868,N_28969,N_29157);
xnor U29869 (N_29869,N_29170,N_28918);
nor U29870 (N_29870,N_29244,N_29311);
or U29871 (N_29871,N_28977,N_29282);
nand U29872 (N_29872,N_28957,N_28886);
nand U29873 (N_29873,N_29380,N_28896);
or U29874 (N_29874,N_28870,N_29179);
nand U29875 (N_29875,N_28973,N_28893);
and U29876 (N_29876,N_28953,N_29373);
xor U29877 (N_29877,N_28996,N_28910);
nor U29878 (N_29878,N_29140,N_28951);
or U29879 (N_29879,N_29070,N_29125);
or U29880 (N_29880,N_29011,N_29151);
nand U29881 (N_29881,N_29043,N_29307);
nor U29882 (N_29882,N_29031,N_29376);
xor U29883 (N_29883,N_29310,N_29232);
xor U29884 (N_29884,N_29094,N_28939);
nor U29885 (N_29885,N_28934,N_28944);
nor U29886 (N_29886,N_29228,N_28870);
and U29887 (N_29887,N_28977,N_29292);
nand U29888 (N_29888,N_28886,N_29034);
or U29889 (N_29889,N_28927,N_29147);
and U29890 (N_29890,N_29338,N_28800);
xnor U29891 (N_29891,N_29237,N_28957);
nor U29892 (N_29892,N_28946,N_29059);
and U29893 (N_29893,N_29176,N_29095);
nor U29894 (N_29894,N_28891,N_29199);
or U29895 (N_29895,N_28895,N_29194);
nand U29896 (N_29896,N_29228,N_29238);
nor U29897 (N_29897,N_29230,N_29266);
or U29898 (N_29898,N_29330,N_29214);
or U29899 (N_29899,N_29026,N_28828);
nor U29900 (N_29900,N_28926,N_29184);
or U29901 (N_29901,N_28829,N_28998);
and U29902 (N_29902,N_28941,N_29371);
or U29903 (N_29903,N_28914,N_28819);
and U29904 (N_29904,N_29289,N_29150);
nand U29905 (N_29905,N_28905,N_29092);
xor U29906 (N_29906,N_29196,N_29141);
xor U29907 (N_29907,N_28833,N_28837);
xor U29908 (N_29908,N_28807,N_29175);
xor U29909 (N_29909,N_29329,N_29254);
xor U29910 (N_29910,N_28944,N_28860);
xor U29911 (N_29911,N_29110,N_28829);
nand U29912 (N_29912,N_28973,N_28885);
nor U29913 (N_29913,N_28886,N_29027);
xnor U29914 (N_29914,N_29283,N_29329);
and U29915 (N_29915,N_29007,N_29224);
nor U29916 (N_29916,N_28861,N_28927);
or U29917 (N_29917,N_29287,N_28843);
nor U29918 (N_29918,N_28907,N_29091);
xor U29919 (N_29919,N_29355,N_29334);
nand U29920 (N_29920,N_29140,N_29389);
and U29921 (N_29921,N_29029,N_28828);
and U29922 (N_29922,N_28936,N_29315);
or U29923 (N_29923,N_28899,N_29183);
or U29924 (N_29924,N_29343,N_29399);
and U29925 (N_29925,N_29058,N_29052);
nand U29926 (N_29926,N_28970,N_29288);
nor U29927 (N_29927,N_29355,N_29138);
xnor U29928 (N_29928,N_29320,N_29013);
nor U29929 (N_29929,N_29315,N_29104);
xnor U29930 (N_29930,N_29217,N_29231);
nand U29931 (N_29931,N_29091,N_29302);
nand U29932 (N_29932,N_29106,N_28951);
nand U29933 (N_29933,N_29158,N_29347);
or U29934 (N_29934,N_29268,N_29322);
nor U29935 (N_29935,N_29286,N_28871);
nor U29936 (N_29936,N_29136,N_29134);
or U29937 (N_29937,N_29371,N_29073);
xor U29938 (N_29938,N_28818,N_29064);
nor U29939 (N_29939,N_28836,N_29120);
nand U29940 (N_29940,N_29132,N_28867);
and U29941 (N_29941,N_29059,N_29265);
and U29942 (N_29942,N_28938,N_29077);
nor U29943 (N_29943,N_28808,N_29342);
nor U29944 (N_29944,N_28988,N_29067);
and U29945 (N_29945,N_29204,N_28934);
or U29946 (N_29946,N_28872,N_28845);
or U29947 (N_29947,N_29066,N_29392);
and U29948 (N_29948,N_29167,N_29117);
nand U29949 (N_29949,N_29207,N_29325);
or U29950 (N_29950,N_29268,N_29120);
nor U29951 (N_29951,N_29133,N_29217);
or U29952 (N_29952,N_28803,N_29200);
or U29953 (N_29953,N_29098,N_28851);
nor U29954 (N_29954,N_29145,N_29274);
or U29955 (N_29955,N_28863,N_29010);
nor U29956 (N_29956,N_29229,N_28885);
xor U29957 (N_29957,N_28837,N_29035);
and U29958 (N_29958,N_29258,N_29038);
and U29959 (N_29959,N_29127,N_29100);
nor U29960 (N_29960,N_29262,N_29320);
nand U29961 (N_29961,N_29183,N_29209);
nand U29962 (N_29962,N_29117,N_28981);
or U29963 (N_29963,N_29105,N_29192);
nor U29964 (N_29964,N_28942,N_29134);
nor U29965 (N_29965,N_29130,N_28900);
or U29966 (N_29966,N_29191,N_29208);
nor U29967 (N_29967,N_28972,N_29073);
nand U29968 (N_29968,N_29340,N_28890);
or U29969 (N_29969,N_28823,N_29144);
nand U29970 (N_29970,N_28907,N_28979);
nor U29971 (N_29971,N_29050,N_28980);
nor U29972 (N_29972,N_28934,N_29112);
nor U29973 (N_29973,N_28842,N_28889);
or U29974 (N_29974,N_29327,N_28940);
or U29975 (N_29975,N_29354,N_29070);
xnor U29976 (N_29976,N_29054,N_29357);
and U29977 (N_29977,N_28985,N_29348);
xnor U29978 (N_29978,N_28931,N_29291);
nand U29979 (N_29979,N_29184,N_29304);
xnor U29980 (N_29980,N_29038,N_29121);
and U29981 (N_29981,N_29384,N_29310);
or U29982 (N_29982,N_28935,N_28811);
or U29983 (N_29983,N_29142,N_28913);
nor U29984 (N_29984,N_29077,N_28862);
and U29985 (N_29985,N_29154,N_29026);
or U29986 (N_29986,N_29200,N_28919);
and U29987 (N_29987,N_29014,N_29393);
or U29988 (N_29988,N_29186,N_29224);
and U29989 (N_29989,N_28910,N_28990);
or U29990 (N_29990,N_29377,N_28845);
nand U29991 (N_29991,N_29157,N_28939);
nand U29992 (N_29992,N_29324,N_29206);
nor U29993 (N_29993,N_29122,N_29001);
nor U29994 (N_29994,N_28805,N_29256);
and U29995 (N_29995,N_29380,N_28853);
and U29996 (N_29996,N_29272,N_29032);
nor U29997 (N_29997,N_29218,N_29171);
xnor U29998 (N_29998,N_29020,N_29277);
nor U29999 (N_29999,N_28881,N_29168);
xor UO_0 (O_0,N_29784,N_29911);
nor UO_1 (O_1,N_29558,N_29456);
or UO_2 (O_2,N_29413,N_29457);
nor UO_3 (O_3,N_29451,N_29735);
or UO_4 (O_4,N_29710,N_29483);
nand UO_5 (O_5,N_29706,N_29926);
xnor UO_6 (O_6,N_29914,N_29793);
or UO_7 (O_7,N_29465,N_29832);
or UO_8 (O_8,N_29750,N_29595);
xnor UO_9 (O_9,N_29461,N_29920);
xor UO_10 (O_10,N_29912,N_29455);
xor UO_11 (O_11,N_29661,N_29765);
and UO_12 (O_12,N_29759,N_29788);
or UO_13 (O_13,N_29825,N_29437);
nor UO_14 (O_14,N_29683,N_29726);
nand UO_15 (O_15,N_29538,N_29981);
and UO_16 (O_16,N_29831,N_29688);
or UO_17 (O_17,N_29858,N_29887);
and UO_18 (O_18,N_29962,N_29527);
xnor UO_19 (O_19,N_29497,N_29725);
or UO_20 (O_20,N_29507,N_29857);
or UO_21 (O_21,N_29877,N_29939);
xor UO_22 (O_22,N_29980,N_29739);
nor UO_23 (O_23,N_29593,N_29448);
and UO_24 (O_24,N_29771,N_29740);
nand UO_25 (O_25,N_29879,N_29623);
or UO_26 (O_26,N_29770,N_29466);
nand UO_27 (O_27,N_29910,N_29473);
nand UO_28 (O_28,N_29500,N_29947);
xor UO_29 (O_29,N_29731,N_29572);
and UO_30 (O_30,N_29485,N_29961);
nor UO_31 (O_31,N_29417,N_29443);
and UO_32 (O_32,N_29848,N_29976);
or UO_33 (O_33,N_29892,N_29699);
nand UO_34 (O_34,N_29612,N_29607);
nor UO_35 (O_35,N_29539,N_29563);
nand UO_36 (O_36,N_29732,N_29436);
nor UO_37 (O_37,N_29493,N_29773);
nor UO_38 (O_38,N_29797,N_29542);
and UO_39 (O_39,N_29954,N_29772);
or UO_40 (O_40,N_29746,N_29968);
nor UO_41 (O_41,N_29988,N_29641);
nand UO_42 (O_42,N_29600,N_29479);
xor UO_43 (O_43,N_29960,N_29843);
or UO_44 (O_44,N_29841,N_29511);
or UO_45 (O_45,N_29454,N_29444);
nand UO_46 (O_46,N_29452,N_29591);
xor UO_47 (O_47,N_29575,N_29907);
nor UO_48 (O_48,N_29780,N_29551);
or UO_49 (O_49,N_29894,N_29628);
nand UO_50 (O_50,N_29696,N_29760);
xor UO_51 (O_51,N_29526,N_29668);
and UO_52 (O_52,N_29667,N_29653);
nor UO_53 (O_53,N_29897,N_29973);
or UO_54 (O_54,N_29613,N_29734);
nor UO_55 (O_55,N_29932,N_29764);
or UO_56 (O_56,N_29634,N_29811);
nand UO_57 (O_57,N_29953,N_29785);
or UO_58 (O_58,N_29618,N_29700);
xor UO_59 (O_59,N_29669,N_29547);
nor UO_60 (O_60,N_29581,N_29895);
nand UO_61 (O_61,N_29923,N_29498);
and UO_62 (O_62,N_29453,N_29676);
or UO_63 (O_63,N_29549,N_29899);
or UO_64 (O_64,N_29862,N_29602);
xnor UO_65 (O_65,N_29543,N_29475);
nor UO_66 (O_66,N_29643,N_29698);
or UO_67 (O_67,N_29930,N_29477);
xnor UO_68 (O_68,N_29738,N_29870);
or UO_69 (O_69,N_29809,N_29412);
or UO_70 (O_70,N_29918,N_29824);
and UO_71 (O_71,N_29971,N_29402);
xnor UO_72 (O_72,N_29422,N_29712);
nor UO_73 (O_73,N_29666,N_29671);
nor UO_74 (O_74,N_29817,N_29404);
or UO_75 (O_75,N_29790,N_29847);
nand UO_76 (O_76,N_29680,N_29938);
or UO_77 (O_77,N_29723,N_29830);
nor UO_78 (O_78,N_29482,N_29576);
nor UO_79 (O_79,N_29946,N_29878);
xnor UO_80 (O_80,N_29645,N_29521);
and UO_81 (O_81,N_29836,N_29516);
xor UO_82 (O_82,N_29820,N_29950);
nand UO_83 (O_83,N_29484,N_29619);
or UO_84 (O_84,N_29405,N_29761);
nand UO_85 (O_85,N_29503,N_29424);
nor UO_86 (O_86,N_29873,N_29801);
and UO_87 (O_87,N_29789,N_29640);
nand UO_88 (O_88,N_29693,N_29625);
or UO_89 (O_89,N_29604,N_29467);
nor UO_90 (O_90,N_29999,N_29664);
or UO_91 (O_91,N_29917,N_29719);
xor UO_92 (O_92,N_29989,N_29967);
and UO_93 (O_93,N_29942,N_29798);
xnor UO_94 (O_94,N_29983,N_29545);
xor UO_95 (O_95,N_29481,N_29684);
nand UO_96 (O_96,N_29646,N_29502);
nand UO_97 (O_97,N_29695,N_29990);
xnor UO_98 (O_98,N_29506,N_29766);
nor UO_99 (O_99,N_29733,N_29865);
nor UO_100 (O_100,N_29838,N_29852);
or UO_101 (O_101,N_29615,N_29845);
nand UO_102 (O_102,N_29494,N_29569);
and UO_103 (O_103,N_29590,N_29863);
nor UO_104 (O_104,N_29963,N_29508);
nor UO_105 (O_105,N_29903,N_29501);
nor UO_106 (O_106,N_29587,N_29513);
nand UO_107 (O_107,N_29639,N_29745);
or UO_108 (O_108,N_29450,N_29837);
nor UO_109 (O_109,N_29647,N_29660);
or UO_110 (O_110,N_29802,N_29753);
and UO_111 (O_111,N_29742,N_29617);
or UO_112 (O_112,N_29889,N_29974);
nand UO_113 (O_113,N_29702,N_29560);
nand UO_114 (O_114,N_29685,N_29977);
and UO_115 (O_115,N_29985,N_29626);
xor UO_116 (O_116,N_29658,N_29557);
nor UO_117 (O_117,N_29813,N_29534);
nor UO_118 (O_118,N_29565,N_29902);
nand UO_119 (O_119,N_29420,N_29823);
and UO_120 (O_120,N_29975,N_29470);
nor UO_121 (O_121,N_29499,N_29401);
nor UO_122 (O_122,N_29979,N_29901);
nor UO_123 (O_123,N_29927,N_29559);
nand UO_124 (O_124,N_29919,N_29803);
nand UO_125 (O_125,N_29808,N_29799);
and UO_126 (O_126,N_29921,N_29654);
nand UO_127 (O_127,N_29578,N_29655);
and UO_128 (O_128,N_29864,N_29818);
or UO_129 (O_129,N_29426,N_29574);
nor UO_130 (O_130,N_29906,N_29540);
nand UO_131 (O_131,N_29629,N_29792);
and UO_132 (O_132,N_29851,N_29544);
xnor UO_133 (O_133,N_29495,N_29636);
nand UO_134 (O_134,N_29925,N_29632);
xnor UO_135 (O_135,N_29682,N_29867);
nor UO_136 (O_136,N_29692,N_29550);
nor UO_137 (O_137,N_29987,N_29638);
or UO_138 (O_138,N_29714,N_29828);
xnor UO_139 (O_139,N_29582,N_29969);
and UO_140 (O_140,N_29909,N_29440);
or UO_141 (O_141,N_29812,N_29767);
nor UO_142 (O_142,N_29517,N_29815);
nand UO_143 (O_143,N_29562,N_29986);
nor UO_144 (O_144,N_29561,N_29447);
and UO_145 (O_145,N_29425,N_29880);
nand UO_146 (O_146,N_29642,N_29694);
xor UO_147 (O_147,N_29594,N_29995);
or UO_148 (O_148,N_29536,N_29614);
nand UO_149 (O_149,N_29997,N_29535);
and UO_150 (O_150,N_29896,N_29786);
nand UO_151 (O_151,N_29672,N_29621);
or UO_152 (O_152,N_29755,N_29428);
xor UO_153 (O_153,N_29566,N_29480);
or UO_154 (O_154,N_29966,N_29598);
nor UO_155 (O_155,N_29728,N_29603);
or UO_156 (O_156,N_29414,N_29711);
or UO_157 (O_157,N_29774,N_29807);
xnor UO_158 (O_158,N_29573,N_29984);
xnor UO_159 (O_159,N_29842,N_29609);
xnor UO_160 (O_160,N_29652,N_29757);
nor UO_161 (O_161,N_29514,N_29644);
xor UO_162 (O_162,N_29724,N_29687);
xor UO_163 (O_163,N_29537,N_29616);
nor UO_164 (O_164,N_29935,N_29421);
and UO_165 (O_165,N_29721,N_29541);
nand UO_166 (O_166,N_29662,N_29522);
xor UO_167 (O_167,N_29934,N_29675);
nor UO_168 (O_168,N_29430,N_29601);
and UO_169 (O_169,N_29528,N_29637);
nand UO_170 (O_170,N_29720,N_29861);
and UO_171 (O_171,N_29936,N_29596);
or UO_172 (O_172,N_29474,N_29471);
and UO_173 (O_173,N_29821,N_29915);
nor UO_174 (O_174,N_29834,N_29835);
nand UO_175 (O_175,N_29605,N_29610);
and UO_176 (O_176,N_29805,N_29580);
xor UO_177 (O_177,N_29872,N_29588);
and UO_178 (O_178,N_29442,N_29577);
nor UO_179 (O_179,N_29679,N_29743);
or UO_180 (O_180,N_29592,N_29881);
xor UO_181 (O_181,N_29476,N_29568);
nor UO_182 (O_182,N_29904,N_29427);
or UO_183 (O_183,N_29648,N_29875);
nor UO_184 (O_184,N_29690,N_29972);
nand UO_185 (O_185,N_29762,N_29869);
or UO_186 (O_186,N_29599,N_29491);
nor UO_187 (O_187,N_29955,N_29890);
or UO_188 (O_188,N_29717,N_29620);
or UO_189 (O_189,N_29900,N_29518);
xnor UO_190 (O_190,N_29589,N_29747);
and UO_191 (O_191,N_29978,N_29438);
or UO_192 (O_192,N_29718,N_29931);
nor UO_193 (O_193,N_29776,N_29781);
xor UO_194 (O_194,N_29850,N_29853);
and UO_195 (O_195,N_29597,N_29713);
and UO_196 (O_196,N_29553,N_29663);
nor UO_197 (O_197,N_29703,N_29673);
nor UO_198 (O_198,N_29439,N_29727);
xor UO_199 (O_199,N_29697,N_29525);
xnor UO_200 (O_200,N_29775,N_29940);
nand UO_201 (O_201,N_29678,N_29548);
or UO_202 (O_202,N_29691,N_29844);
nand UO_203 (O_203,N_29937,N_29729);
nand UO_204 (O_204,N_29686,N_29716);
and UO_205 (O_205,N_29994,N_29464);
or UO_206 (O_206,N_29840,N_29949);
xor UO_207 (O_207,N_29856,N_29783);
nand UO_208 (O_208,N_29886,N_29556);
nand UO_209 (O_209,N_29749,N_29606);
or UO_210 (O_210,N_29519,N_29410);
nor UO_211 (O_211,N_29419,N_29496);
xor UO_212 (O_212,N_29933,N_29860);
nand UO_213 (O_213,N_29488,N_29406);
or UO_214 (O_214,N_29744,N_29631);
or UO_215 (O_215,N_29871,N_29650);
and UO_216 (O_216,N_29891,N_29701);
nor UO_217 (O_217,N_29800,N_29510);
xor UO_218 (O_218,N_29996,N_29445);
xor UO_219 (O_219,N_29893,N_29751);
nand UO_220 (O_220,N_29570,N_29492);
nor UO_221 (O_221,N_29630,N_29504);
or UO_222 (O_222,N_29787,N_29957);
and UO_223 (O_223,N_29552,N_29737);
nor UO_224 (O_224,N_29777,N_29884);
or UO_225 (O_225,N_29585,N_29400);
or UO_226 (O_226,N_29964,N_29730);
nor UO_227 (O_227,N_29418,N_29458);
nor UO_228 (O_228,N_29463,N_29991);
or UO_229 (O_229,N_29584,N_29722);
xor UO_230 (O_230,N_29965,N_29833);
or UO_231 (O_231,N_29674,N_29433);
xor UO_232 (O_232,N_29622,N_29822);
and UO_233 (O_233,N_29469,N_29681);
or UO_234 (O_234,N_29952,N_29411);
xnor UO_235 (O_235,N_29959,N_29707);
or UO_236 (O_236,N_29806,N_29791);
nor UO_237 (O_237,N_29778,N_29533);
and UO_238 (O_238,N_29407,N_29478);
or UO_239 (O_239,N_29882,N_29929);
or UO_240 (O_240,N_29656,N_29754);
nor UO_241 (O_241,N_29489,N_29705);
and UO_242 (O_242,N_29758,N_29768);
nor UO_243 (O_243,N_29462,N_29846);
or UO_244 (O_244,N_29423,N_29571);
nand UO_245 (O_245,N_29992,N_29736);
xnor UO_246 (O_246,N_29659,N_29429);
xnor UO_247 (O_247,N_29715,N_29922);
or UO_248 (O_248,N_29564,N_29855);
or UO_249 (O_249,N_29472,N_29866);
nand UO_250 (O_250,N_29839,N_29416);
nor UO_251 (O_251,N_29819,N_29515);
nand UO_252 (O_252,N_29948,N_29868);
and UO_253 (O_253,N_29409,N_29532);
nand UO_254 (O_254,N_29804,N_29898);
and UO_255 (O_255,N_29885,N_29859);
or UO_256 (O_256,N_29849,N_29982);
nor UO_257 (O_257,N_29524,N_29509);
and UO_258 (O_258,N_29708,N_29567);
or UO_259 (O_259,N_29993,N_29794);
and UO_260 (O_260,N_29970,N_29709);
nor UO_261 (O_261,N_29633,N_29814);
and UO_262 (O_262,N_29958,N_29829);
nand UO_263 (O_263,N_29649,N_29651);
xnor UO_264 (O_264,N_29554,N_29795);
and UO_265 (O_265,N_29468,N_29512);
nor UO_266 (O_266,N_29432,N_29555);
and UO_267 (O_267,N_29916,N_29435);
nor UO_268 (O_268,N_29941,N_29769);
nor UO_269 (O_269,N_29928,N_29956);
nand UO_270 (O_270,N_29403,N_29810);
nor UO_271 (O_271,N_29827,N_29529);
xnor UO_272 (O_272,N_29951,N_29490);
nor UO_273 (O_273,N_29756,N_29624);
nand UO_274 (O_274,N_29816,N_29883);
nand UO_275 (O_275,N_29505,N_29908);
nor UO_276 (O_276,N_29446,N_29449);
or UO_277 (O_277,N_29874,N_29748);
or UO_278 (O_278,N_29531,N_29796);
xnor UO_279 (O_279,N_29945,N_29741);
and UO_280 (O_280,N_29998,N_29459);
xnor UO_281 (O_281,N_29408,N_29689);
nor UO_282 (O_282,N_29854,N_29586);
nor UO_283 (O_283,N_29826,N_29752);
xor UO_284 (O_284,N_29530,N_29924);
xor UO_285 (O_285,N_29943,N_29677);
and UO_286 (O_286,N_29431,N_29441);
and UO_287 (O_287,N_29434,N_29763);
xnor UO_288 (O_288,N_29579,N_29460);
xnor UO_289 (O_289,N_29665,N_29704);
xnor UO_290 (O_290,N_29635,N_29913);
or UO_291 (O_291,N_29888,N_29627);
or UO_292 (O_292,N_29611,N_29657);
and UO_293 (O_293,N_29876,N_29546);
nor UO_294 (O_294,N_29944,N_29487);
xor UO_295 (O_295,N_29608,N_29779);
and UO_296 (O_296,N_29583,N_29520);
nor UO_297 (O_297,N_29670,N_29523);
nand UO_298 (O_298,N_29782,N_29415);
nor UO_299 (O_299,N_29905,N_29486);
or UO_300 (O_300,N_29768,N_29706);
xnor UO_301 (O_301,N_29954,N_29557);
or UO_302 (O_302,N_29834,N_29494);
nor UO_303 (O_303,N_29564,N_29827);
nor UO_304 (O_304,N_29423,N_29641);
or UO_305 (O_305,N_29683,N_29997);
nand UO_306 (O_306,N_29828,N_29919);
nand UO_307 (O_307,N_29561,N_29983);
or UO_308 (O_308,N_29996,N_29884);
nor UO_309 (O_309,N_29851,N_29453);
and UO_310 (O_310,N_29552,N_29753);
nor UO_311 (O_311,N_29864,N_29903);
xor UO_312 (O_312,N_29527,N_29971);
or UO_313 (O_313,N_29785,N_29801);
nor UO_314 (O_314,N_29685,N_29738);
xor UO_315 (O_315,N_29751,N_29581);
nor UO_316 (O_316,N_29536,N_29521);
nor UO_317 (O_317,N_29945,N_29577);
and UO_318 (O_318,N_29429,N_29496);
xnor UO_319 (O_319,N_29592,N_29760);
nand UO_320 (O_320,N_29695,N_29856);
and UO_321 (O_321,N_29805,N_29879);
or UO_322 (O_322,N_29669,N_29751);
or UO_323 (O_323,N_29638,N_29452);
nor UO_324 (O_324,N_29904,N_29554);
or UO_325 (O_325,N_29825,N_29620);
and UO_326 (O_326,N_29654,N_29764);
nor UO_327 (O_327,N_29875,N_29426);
xor UO_328 (O_328,N_29858,N_29851);
or UO_329 (O_329,N_29944,N_29819);
nor UO_330 (O_330,N_29986,N_29439);
or UO_331 (O_331,N_29439,N_29562);
and UO_332 (O_332,N_29736,N_29737);
or UO_333 (O_333,N_29514,N_29862);
or UO_334 (O_334,N_29426,N_29732);
nor UO_335 (O_335,N_29837,N_29419);
or UO_336 (O_336,N_29656,N_29454);
nand UO_337 (O_337,N_29705,N_29571);
nand UO_338 (O_338,N_29589,N_29480);
xnor UO_339 (O_339,N_29708,N_29741);
nand UO_340 (O_340,N_29702,N_29524);
or UO_341 (O_341,N_29594,N_29630);
or UO_342 (O_342,N_29671,N_29762);
or UO_343 (O_343,N_29973,N_29796);
and UO_344 (O_344,N_29718,N_29729);
nand UO_345 (O_345,N_29776,N_29674);
and UO_346 (O_346,N_29716,N_29931);
or UO_347 (O_347,N_29505,N_29980);
and UO_348 (O_348,N_29903,N_29922);
nand UO_349 (O_349,N_29880,N_29825);
or UO_350 (O_350,N_29474,N_29626);
or UO_351 (O_351,N_29955,N_29800);
xor UO_352 (O_352,N_29955,N_29699);
nor UO_353 (O_353,N_29521,N_29418);
or UO_354 (O_354,N_29641,N_29539);
nand UO_355 (O_355,N_29456,N_29476);
xor UO_356 (O_356,N_29492,N_29664);
and UO_357 (O_357,N_29783,N_29878);
nor UO_358 (O_358,N_29711,N_29751);
or UO_359 (O_359,N_29418,N_29513);
nor UO_360 (O_360,N_29738,N_29416);
nor UO_361 (O_361,N_29655,N_29413);
xnor UO_362 (O_362,N_29685,N_29833);
or UO_363 (O_363,N_29684,N_29681);
xnor UO_364 (O_364,N_29603,N_29552);
and UO_365 (O_365,N_29818,N_29965);
or UO_366 (O_366,N_29550,N_29455);
nand UO_367 (O_367,N_29896,N_29619);
xor UO_368 (O_368,N_29430,N_29873);
xor UO_369 (O_369,N_29535,N_29450);
or UO_370 (O_370,N_29794,N_29983);
and UO_371 (O_371,N_29714,N_29969);
nand UO_372 (O_372,N_29963,N_29957);
or UO_373 (O_373,N_29493,N_29934);
and UO_374 (O_374,N_29403,N_29998);
or UO_375 (O_375,N_29507,N_29818);
nand UO_376 (O_376,N_29782,N_29437);
nor UO_377 (O_377,N_29651,N_29761);
xnor UO_378 (O_378,N_29600,N_29672);
or UO_379 (O_379,N_29909,N_29584);
or UO_380 (O_380,N_29680,N_29847);
nor UO_381 (O_381,N_29716,N_29937);
and UO_382 (O_382,N_29763,N_29483);
xnor UO_383 (O_383,N_29523,N_29839);
or UO_384 (O_384,N_29415,N_29667);
xor UO_385 (O_385,N_29872,N_29509);
or UO_386 (O_386,N_29691,N_29922);
xor UO_387 (O_387,N_29655,N_29780);
nand UO_388 (O_388,N_29544,N_29947);
or UO_389 (O_389,N_29758,N_29460);
or UO_390 (O_390,N_29950,N_29602);
nand UO_391 (O_391,N_29974,N_29951);
and UO_392 (O_392,N_29784,N_29707);
nand UO_393 (O_393,N_29774,N_29944);
nor UO_394 (O_394,N_29812,N_29835);
and UO_395 (O_395,N_29847,N_29904);
and UO_396 (O_396,N_29928,N_29578);
or UO_397 (O_397,N_29698,N_29863);
xor UO_398 (O_398,N_29747,N_29868);
or UO_399 (O_399,N_29546,N_29855);
and UO_400 (O_400,N_29760,N_29993);
nand UO_401 (O_401,N_29585,N_29950);
or UO_402 (O_402,N_29967,N_29920);
nand UO_403 (O_403,N_29805,N_29440);
or UO_404 (O_404,N_29508,N_29501);
and UO_405 (O_405,N_29517,N_29947);
nand UO_406 (O_406,N_29950,N_29555);
nand UO_407 (O_407,N_29444,N_29757);
nor UO_408 (O_408,N_29692,N_29702);
xor UO_409 (O_409,N_29494,N_29986);
nor UO_410 (O_410,N_29422,N_29765);
xnor UO_411 (O_411,N_29612,N_29549);
nand UO_412 (O_412,N_29711,N_29561);
or UO_413 (O_413,N_29889,N_29493);
nor UO_414 (O_414,N_29598,N_29437);
or UO_415 (O_415,N_29978,N_29666);
xnor UO_416 (O_416,N_29621,N_29999);
nand UO_417 (O_417,N_29994,N_29748);
xor UO_418 (O_418,N_29921,N_29704);
nor UO_419 (O_419,N_29415,N_29825);
xnor UO_420 (O_420,N_29863,N_29880);
or UO_421 (O_421,N_29841,N_29937);
nor UO_422 (O_422,N_29462,N_29767);
and UO_423 (O_423,N_29558,N_29419);
xor UO_424 (O_424,N_29684,N_29410);
or UO_425 (O_425,N_29561,N_29531);
and UO_426 (O_426,N_29731,N_29702);
xnor UO_427 (O_427,N_29604,N_29959);
nor UO_428 (O_428,N_29774,N_29409);
and UO_429 (O_429,N_29606,N_29938);
nor UO_430 (O_430,N_29466,N_29896);
xnor UO_431 (O_431,N_29452,N_29721);
or UO_432 (O_432,N_29862,N_29819);
xnor UO_433 (O_433,N_29818,N_29953);
nor UO_434 (O_434,N_29566,N_29782);
nor UO_435 (O_435,N_29752,N_29840);
or UO_436 (O_436,N_29872,N_29855);
or UO_437 (O_437,N_29487,N_29824);
and UO_438 (O_438,N_29979,N_29914);
nor UO_439 (O_439,N_29530,N_29804);
nor UO_440 (O_440,N_29745,N_29580);
nand UO_441 (O_441,N_29856,N_29550);
or UO_442 (O_442,N_29404,N_29666);
and UO_443 (O_443,N_29947,N_29721);
and UO_444 (O_444,N_29964,N_29734);
and UO_445 (O_445,N_29801,N_29619);
nor UO_446 (O_446,N_29652,N_29554);
or UO_447 (O_447,N_29819,N_29826);
xnor UO_448 (O_448,N_29559,N_29658);
xor UO_449 (O_449,N_29624,N_29442);
nand UO_450 (O_450,N_29498,N_29666);
and UO_451 (O_451,N_29641,N_29601);
and UO_452 (O_452,N_29946,N_29701);
xor UO_453 (O_453,N_29437,N_29682);
nor UO_454 (O_454,N_29804,N_29713);
and UO_455 (O_455,N_29404,N_29697);
nor UO_456 (O_456,N_29835,N_29731);
xor UO_457 (O_457,N_29598,N_29896);
or UO_458 (O_458,N_29491,N_29764);
nor UO_459 (O_459,N_29662,N_29430);
nand UO_460 (O_460,N_29475,N_29937);
nor UO_461 (O_461,N_29738,N_29793);
xor UO_462 (O_462,N_29786,N_29956);
or UO_463 (O_463,N_29554,N_29925);
and UO_464 (O_464,N_29917,N_29728);
or UO_465 (O_465,N_29766,N_29534);
xnor UO_466 (O_466,N_29673,N_29681);
nor UO_467 (O_467,N_29702,N_29464);
xor UO_468 (O_468,N_29857,N_29557);
xnor UO_469 (O_469,N_29891,N_29772);
nand UO_470 (O_470,N_29431,N_29673);
or UO_471 (O_471,N_29883,N_29722);
nor UO_472 (O_472,N_29531,N_29547);
nor UO_473 (O_473,N_29764,N_29817);
and UO_474 (O_474,N_29834,N_29519);
nand UO_475 (O_475,N_29813,N_29941);
xnor UO_476 (O_476,N_29743,N_29658);
xor UO_477 (O_477,N_29546,N_29988);
or UO_478 (O_478,N_29652,N_29807);
and UO_479 (O_479,N_29993,N_29615);
nor UO_480 (O_480,N_29546,N_29787);
nor UO_481 (O_481,N_29746,N_29846);
nand UO_482 (O_482,N_29457,N_29815);
and UO_483 (O_483,N_29709,N_29809);
or UO_484 (O_484,N_29457,N_29478);
and UO_485 (O_485,N_29989,N_29947);
xnor UO_486 (O_486,N_29957,N_29509);
or UO_487 (O_487,N_29474,N_29686);
and UO_488 (O_488,N_29960,N_29538);
nand UO_489 (O_489,N_29497,N_29469);
or UO_490 (O_490,N_29617,N_29674);
nor UO_491 (O_491,N_29511,N_29636);
and UO_492 (O_492,N_29619,N_29751);
and UO_493 (O_493,N_29648,N_29612);
nor UO_494 (O_494,N_29961,N_29533);
or UO_495 (O_495,N_29822,N_29558);
nor UO_496 (O_496,N_29706,N_29921);
and UO_497 (O_497,N_29555,N_29452);
nand UO_498 (O_498,N_29495,N_29583);
and UO_499 (O_499,N_29560,N_29979);
and UO_500 (O_500,N_29411,N_29570);
nor UO_501 (O_501,N_29462,N_29526);
xor UO_502 (O_502,N_29511,N_29792);
xor UO_503 (O_503,N_29871,N_29531);
and UO_504 (O_504,N_29850,N_29420);
nor UO_505 (O_505,N_29871,N_29533);
xor UO_506 (O_506,N_29842,N_29458);
xnor UO_507 (O_507,N_29743,N_29462);
and UO_508 (O_508,N_29802,N_29828);
xnor UO_509 (O_509,N_29858,N_29962);
or UO_510 (O_510,N_29886,N_29797);
or UO_511 (O_511,N_29691,N_29896);
nor UO_512 (O_512,N_29636,N_29540);
nand UO_513 (O_513,N_29585,N_29739);
nand UO_514 (O_514,N_29675,N_29851);
nor UO_515 (O_515,N_29630,N_29569);
nand UO_516 (O_516,N_29547,N_29580);
nand UO_517 (O_517,N_29849,N_29614);
and UO_518 (O_518,N_29775,N_29430);
and UO_519 (O_519,N_29904,N_29950);
nor UO_520 (O_520,N_29445,N_29816);
nor UO_521 (O_521,N_29481,N_29850);
nand UO_522 (O_522,N_29834,N_29433);
and UO_523 (O_523,N_29657,N_29793);
xor UO_524 (O_524,N_29407,N_29919);
and UO_525 (O_525,N_29490,N_29468);
xnor UO_526 (O_526,N_29610,N_29658);
or UO_527 (O_527,N_29841,N_29788);
nand UO_528 (O_528,N_29642,N_29931);
or UO_529 (O_529,N_29522,N_29815);
nand UO_530 (O_530,N_29906,N_29729);
xor UO_531 (O_531,N_29450,N_29561);
and UO_532 (O_532,N_29552,N_29657);
or UO_533 (O_533,N_29402,N_29702);
nor UO_534 (O_534,N_29945,N_29578);
and UO_535 (O_535,N_29999,N_29618);
and UO_536 (O_536,N_29595,N_29978);
nor UO_537 (O_537,N_29468,N_29569);
xnor UO_538 (O_538,N_29742,N_29773);
xor UO_539 (O_539,N_29829,N_29929);
nand UO_540 (O_540,N_29786,N_29429);
xnor UO_541 (O_541,N_29688,N_29755);
xor UO_542 (O_542,N_29599,N_29405);
nor UO_543 (O_543,N_29980,N_29765);
xnor UO_544 (O_544,N_29955,N_29403);
nand UO_545 (O_545,N_29892,N_29783);
or UO_546 (O_546,N_29587,N_29628);
or UO_547 (O_547,N_29623,N_29580);
and UO_548 (O_548,N_29606,N_29755);
xor UO_549 (O_549,N_29982,N_29857);
xor UO_550 (O_550,N_29491,N_29913);
and UO_551 (O_551,N_29610,N_29909);
or UO_552 (O_552,N_29669,N_29774);
or UO_553 (O_553,N_29710,N_29752);
or UO_554 (O_554,N_29550,N_29706);
xor UO_555 (O_555,N_29922,N_29633);
nand UO_556 (O_556,N_29959,N_29784);
nand UO_557 (O_557,N_29604,N_29620);
or UO_558 (O_558,N_29828,N_29477);
nand UO_559 (O_559,N_29626,N_29733);
or UO_560 (O_560,N_29785,N_29617);
and UO_561 (O_561,N_29531,N_29660);
nand UO_562 (O_562,N_29755,N_29454);
xnor UO_563 (O_563,N_29420,N_29472);
nor UO_564 (O_564,N_29900,N_29446);
nand UO_565 (O_565,N_29450,N_29708);
and UO_566 (O_566,N_29627,N_29417);
nor UO_567 (O_567,N_29676,N_29460);
nor UO_568 (O_568,N_29568,N_29723);
nor UO_569 (O_569,N_29852,N_29600);
xnor UO_570 (O_570,N_29904,N_29466);
nand UO_571 (O_571,N_29540,N_29658);
nand UO_572 (O_572,N_29993,N_29744);
and UO_573 (O_573,N_29622,N_29679);
and UO_574 (O_574,N_29918,N_29838);
and UO_575 (O_575,N_29679,N_29558);
xnor UO_576 (O_576,N_29472,N_29715);
or UO_577 (O_577,N_29682,N_29575);
nor UO_578 (O_578,N_29833,N_29827);
nor UO_579 (O_579,N_29961,N_29768);
nand UO_580 (O_580,N_29800,N_29458);
xnor UO_581 (O_581,N_29892,N_29839);
and UO_582 (O_582,N_29942,N_29656);
and UO_583 (O_583,N_29817,N_29662);
nor UO_584 (O_584,N_29817,N_29462);
or UO_585 (O_585,N_29787,N_29797);
and UO_586 (O_586,N_29763,N_29958);
nand UO_587 (O_587,N_29656,N_29991);
nor UO_588 (O_588,N_29815,N_29996);
nor UO_589 (O_589,N_29864,N_29931);
xnor UO_590 (O_590,N_29513,N_29645);
nand UO_591 (O_591,N_29705,N_29491);
and UO_592 (O_592,N_29486,N_29933);
xnor UO_593 (O_593,N_29692,N_29928);
and UO_594 (O_594,N_29817,N_29876);
nor UO_595 (O_595,N_29757,N_29996);
nand UO_596 (O_596,N_29953,N_29636);
nor UO_597 (O_597,N_29576,N_29660);
nand UO_598 (O_598,N_29681,N_29971);
and UO_599 (O_599,N_29819,N_29677);
xnor UO_600 (O_600,N_29902,N_29883);
and UO_601 (O_601,N_29460,N_29825);
nor UO_602 (O_602,N_29427,N_29855);
and UO_603 (O_603,N_29482,N_29905);
nand UO_604 (O_604,N_29909,N_29604);
nand UO_605 (O_605,N_29797,N_29916);
and UO_606 (O_606,N_29676,N_29952);
or UO_607 (O_607,N_29646,N_29932);
nor UO_608 (O_608,N_29426,N_29887);
nand UO_609 (O_609,N_29602,N_29467);
xnor UO_610 (O_610,N_29969,N_29776);
and UO_611 (O_611,N_29449,N_29441);
and UO_612 (O_612,N_29980,N_29687);
nor UO_613 (O_613,N_29705,N_29898);
or UO_614 (O_614,N_29451,N_29403);
or UO_615 (O_615,N_29741,N_29929);
xnor UO_616 (O_616,N_29844,N_29819);
xor UO_617 (O_617,N_29672,N_29837);
xnor UO_618 (O_618,N_29932,N_29607);
and UO_619 (O_619,N_29739,N_29990);
and UO_620 (O_620,N_29548,N_29712);
or UO_621 (O_621,N_29477,N_29954);
nor UO_622 (O_622,N_29641,N_29628);
and UO_623 (O_623,N_29901,N_29537);
nand UO_624 (O_624,N_29505,N_29515);
xnor UO_625 (O_625,N_29985,N_29652);
and UO_626 (O_626,N_29541,N_29640);
or UO_627 (O_627,N_29580,N_29688);
nor UO_628 (O_628,N_29698,N_29403);
or UO_629 (O_629,N_29643,N_29672);
and UO_630 (O_630,N_29845,N_29878);
nand UO_631 (O_631,N_29890,N_29782);
and UO_632 (O_632,N_29474,N_29458);
or UO_633 (O_633,N_29909,N_29532);
xor UO_634 (O_634,N_29770,N_29419);
xor UO_635 (O_635,N_29690,N_29696);
and UO_636 (O_636,N_29809,N_29473);
nand UO_637 (O_637,N_29661,N_29964);
nand UO_638 (O_638,N_29869,N_29413);
nor UO_639 (O_639,N_29533,N_29624);
nand UO_640 (O_640,N_29725,N_29893);
nand UO_641 (O_641,N_29675,N_29577);
or UO_642 (O_642,N_29992,N_29883);
or UO_643 (O_643,N_29571,N_29663);
nor UO_644 (O_644,N_29830,N_29518);
nand UO_645 (O_645,N_29646,N_29957);
nand UO_646 (O_646,N_29564,N_29874);
nand UO_647 (O_647,N_29829,N_29523);
or UO_648 (O_648,N_29553,N_29984);
xor UO_649 (O_649,N_29976,N_29565);
and UO_650 (O_650,N_29403,N_29687);
nand UO_651 (O_651,N_29654,N_29766);
xor UO_652 (O_652,N_29905,N_29551);
nor UO_653 (O_653,N_29797,N_29794);
or UO_654 (O_654,N_29680,N_29481);
nor UO_655 (O_655,N_29606,N_29535);
nand UO_656 (O_656,N_29802,N_29966);
and UO_657 (O_657,N_29770,N_29556);
nand UO_658 (O_658,N_29677,N_29955);
nor UO_659 (O_659,N_29506,N_29662);
or UO_660 (O_660,N_29402,N_29816);
xnor UO_661 (O_661,N_29833,N_29519);
and UO_662 (O_662,N_29538,N_29861);
or UO_663 (O_663,N_29498,N_29891);
xor UO_664 (O_664,N_29932,N_29407);
xnor UO_665 (O_665,N_29942,N_29606);
nor UO_666 (O_666,N_29562,N_29919);
or UO_667 (O_667,N_29755,N_29744);
and UO_668 (O_668,N_29631,N_29928);
xnor UO_669 (O_669,N_29575,N_29624);
nand UO_670 (O_670,N_29925,N_29558);
xor UO_671 (O_671,N_29580,N_29861);
nor UO_672 (O_672,N_29725,N_29755);
and UO_673 (O_673,N_29653,N_29569);
nor UO_674 (O_674,N_29676,N_29464);
nand UO_675 (O_675,N_29994,N_29896);
and UO_676 (O_676,N_29607,N_29986);
nor UO_677 (O_677,N_29674,N_29567);
nand UO_678 (O_678,N_29497,N_29638);
xnor UO_679 (O_679,N_29693,N_29797);
nand UO_680 (O_680,N_29706,N_29685);
or UO_681 (O_681,N_29619,N_29875);
or UO_682 (O_682,N_29441,N_29874);
xnor UO_683 (O_683,N_29665,N_29874);
and UO_684 (O_684,N_29502,N_29782);
xnor UO_685 (O_685,N_29743,N_29993);
xor UO_686 (O_686,N_29494,N_29824);
or UO_687 (O_687,N_29651,N_29456);
xor UO_688 (O_688,N_29870,N_29685);
nand UO_689 (O_689,N_29449,N_29499);
xnor UO_690 (O_690,N_29761,N_29861);
nand UO_691 (O_691,N_29994,N_29571);
nor UO_692 (O_692,N_29777,N_29728);
nor UO_693 (O_693,N_29814,N_29567);
or UO_694 (O_694,N_29806,N_29814);
or UO_695 (O_695,N_29783,N_29704);
nand UO_696 (O_696,N_29917,N_29461);
nand UO_697 (O_697,N_29763,N_29706);
nor UO_698 (O_698,N_29910,N_29649);
xnor UO_699 (O_699,N_29452,N_29811);
and UO_700 (O_700,N_29530,N_29960);
xor UO_701 (O_701,N_29904,N_29582);
or UO_702 (O_702,N_29411,N_29808);
or UO_703 (O_703,N_29405,N_29461);
or UO_704 (O_704,N_29922,N_29575);
xor UO_705 (O_705,N_29760,N_29879);
nor UO_706 (O_706,N_29985,N_29750);
xor UO_707 (O_707,N_29432,N_29939);
or UO_708 (O_708,N_29696,N_29703);
nor UO_709 (O_709,N_29849,N_29502);
nand UO_710 (O_710,N_29660,N_29672);
nand UO_711 (O_711,N_29780,N_29613);
nor UO_712 (O_712,N_29863,N_29756);
or UO_713 (O_713,N_29505,N_29937);
nor UO_714 (O_714,N_29632,N_29879);
xnor UO_715 (O_715,N_29886,N_29602);
or UO_716 (O_716,N_29418,N_29959);
nand UO_717 (O_717,N_29418,N_29949);
and UO_718 (O_718,N_29665,N_29851);
nor UO_719 (O_719,N_29735,N_29657);
nand UO_720 (O_720,N_29830,N_29822);
nand UO_721 (O_721,N_29451,N_29763);
and UO_722 (O_722,N_29896,N_29590);
nor UO_723 (O_723,N_29664,N_29728);
or UO_724 (O_724,N_29437,N_29963);
xor UO_725 (O_725,N_29890,N_29478);
nand UO_726 (O_726,N_29454,N_29671);
or UO_727 (O_727,N_29652,N_29441);
nor UO_728 (O_728,N_29474,N_29832);
nand UO_729 (O_729,N_29523,N_29966);
or UO_730 (O_730,N_29903,N_29895);
or UO_731 (O_731,N_29905,N_29668);
and UO_732 (O_732,N_29962,N_29953);
and UO_733 (O_733,N_29921,N_29875);
nand UO_734 (O_734,N_29970,N_29594);
and UO_735 (O_735,N_29891,N_29744);
nor UO_736 (O_736,N_29455,N_29444);
nand UO_737 (O_737,N_29836,N_29573);
or UO_738 (O_738,N_29788,N_29504);
and UO_739 (O_739,N_29854,N_29856);
or UO_740 (O_740,N_29705,N_29518);
or UO_741 (O_741,N_29806,N_29616);
nor UO_742 (O_742,N_29746,N_29792);
or UO_743 (O_743,N_29944,N_29754);
and UO_744 (O_744,N_29648,N_29512);
xor UO_745 (O_745,N_29507,N_29481);
nand UO_746 (O_746,N_29648,N_29743);
xnor UO_747 (O_747,N_29514,N_29863);
xnor UO_748 (O_748,N_29732,N_29439);
or UO_749 (O_749,N_29789,N_29575);
and UO_750 (O_750,N_29472,N_29761);
or UO_751 (O_751,N_29475,N_29897);
nor UO_752 (O_752,N_29921,N_29942);
and UO_753 (O_753,N_29943,N_29435);
xnor UO_754 (O_754,N_29640,N_29662);
and UO_755 (O_755,N_29557,N_29466);
nand UO_756 (O_756,N_29859,N_29585);
xor UO_757 (O_757,N_29877,N_29458);
xor UO_758 (O_758,N_29435,N_29751);
xnor UO_759 (O_759,N_29560,N_29452);
nand UO_760 (O_760,N_29647,N_29888);
and UO_761 (O_761,N_29613,N_29996);
nor UO_762 (O_762,N_29752,N_29440);
or UO_763 (O_763,N_29932,N_29714);
and UO_764 (O_764,N_29523,N_29562);
nand UO_765 (O_765,N_29472,N_29910);
and UO_766 (O_766,N_29843,N_29524);
or UO_767 (O_767,N_29565,N_29844);
xor UO_768 (O_768,N_29929,N_29616);
or UO_769 (O_769,N_29651,N_29962);
and UO_770 (O_770,N_29583,N_29949);
and UO_771 (O_771,N_29834,N_29486);
xnor UO_772 (O_772,N_29853,N_29773);
nor UO_773 (O_773,N_29752,N_29590);
nand UO_774 (O_774,N_29567,N_29685);
or UO_775 (O_775,N_29618,N_29909);
and UO_776 (O_776,N_29436,N_29481);
xnor UO_777 (O_777,N_29698,N_29752);
nor UO_778 (O_778,N_29923,N_29744);
and UO_779 (O_779,N_29801,N_29520);
or UO_780 (O_780,N_29969,N_29611);
or UO_781 (O_781,N_29903,N_29554);
nor UO_782 (O_782,N_29905,N_29724);
nand UO_783 (O_783,N_29433,N_29752);
nand UO_784 (O_784,N_29954,N_29479);
xor UO_785 (O_785,N_29589,N_29915);
nor UO_786 (O_786,N_29915,N_29703);
or UO_787 (O_787,N_29672,N_29685);
and UO_788 (O_788,N_29556,N_29949);
nand UO_789 (O_789,N_29444,N_29580);
or UO_790 (O_790,N_29574,N_29590);
nor UO_791 (O_791,N_29822,N_29705);
xnor UO_792 (O_792,N_29765,N_29445);
and UO_793 (O_793,N_29867,N_29631);
and UO_794 (O_794,N_29656,N_29965);
nand UO_795 (O_795,N_29456,N_29857);
nand UO_796 (O_796,N_29638,N_29456);
nand UO_797 (O_797,N_29970,N_29684);
nand UO_798 (O_798,N_29848,N_29887);
nand UO_799 (O_799,N_29562,N_29464);
nor UO_800 (O_800,N_29500,N_29699);
xnor UO_801 (O_801,N_29802,N_29649);
nor UO_802 (O_802,N_29742,N_29974);
nand UO_803 (O_803,N_29716,N_29943);
nand UO_804 (O_804,N_29607,N_29674);
and UO_805 (O_805,N_29616,N_29663);
nand UO_806 (O_806,N_29954,N_29940);
and UO_807 (O_807,N_29526,N_29783);
or UO_808 (O_808,N_29569,N_29627);
and UO_809 (O_809,N_29418,N_29811);
or UO_810 (O_810,N_29589,N_29663);
nor UO_811 (O_811,N_29909,N_29849);
and UO_812 (O_812,N_29799,N_29723);
xnor UO_813 (O_813,N_29818,N_29524);
nand UO_814 (O_814,N_29770,N_29495);
nand UO_815 (O_815,N_29567,N_29869);
or UO_816 (O_816,N_29700,N_29909);
or UO_817 (O_817,N_29636,N_29654);
xnor UO_818 (O_818,N_29479,N_29957);
and UO_819 (O_819,N_29441,N_29726);
and UO_820 (O_820,N_29477,N_29674);
and UO_821 (O_821,N_29870,N_29500);
nand UO_822 (O_822,N_29586,N_29440);
or UO_823 (O_823,N_29733,N_29927);
and UO_824 (O_824,N_29629,N_29469);
nand UO_825 (O_825,N_29796,N_29479);
nand UO_826 (O_826,N_29576,N_29601);
nand UO_827 (O_827,N_29441,N_29885);
nand UO_828 (O_828,N_29910,N_29979);
xor UO_829 (O_829,N_29932,N_29687);
xnor UO_830 (O_830,N_29973,N_29630);
nor UO_831 (O_831,N_29627,N_29922);
and UO_832 (O_832,N_29556,N_29831);
nor UO_833 (O_833,N_29412,N_29646);
or UO_834 (O_834,N_29598,N_29484);
nor UO_835 (O_835,N_29952,N_29979);
and UO_836 (O_836,N_29636,N_29453);
or UO_837 (O_837,N_29715,N_29505);
xor UO_838 (O_838,N_29660,N_29775);
and UO_839 (O_839,N_29879,N_29482);
nand UO_840 (O_840,N_29740,N_29809);
nor UO_841 (O_841,N_29607,N_29542);
nor UO_842 (O_842,N_29683,N_29676);
and UO_843 (O_843,N_29768,N_29989);
nor UO_844 (O_844,N_29522,N_29884);
nor UO_845 (O_845,N_29893,N_29678);
xor UO_846 (O_846,N_29603,N_29498);
nor UO_847 (O_847,N_29729,N_29798);
and UO_848 (O_848,N_29847,N_29768);
and UO_849 (O_849,N_29540,N_29414);
nand UO_850 (O_850,N_29883,N_29799);
xnor UO_851 (O_851,N_29945,N_29986);
or UO_852 (O_852,N_29684,N_29589);
nand UO_853 (O_853,N_29440,N_29665);
or UO_854 (O_854,N_29421,N_29986);
nand UO_855 (O_855,N_29767,N_29595);
nor UO_856 (O_856,N_29402,N_29774);
xor UO_857 (O_857,N_29934,N_29632);
and UO_858 (O_858,N_29703,N_29949);
xor UO_859 (O_859,N_29407,N_29425);
nor UO_860 (O_860,N_29637,N_29430);
nand UO_861 (O_861,N_29772,N_29463);
or UO_862 (O_862,N_29751,N_29844);
and UO_863 (O_863,N_29789,N_29464);
or UO_864 (O_864,N_29471,N_29731);
nand UO_865 (O_865,N_29878,N_29607);
and UO_866 (O_866,N_29864,N_29708);
or UO_867 (O_867,N_29845,N_29917);
and UO_868 (O_868,N_29961,N_29972);
nor UO_869 (O_869,N_29766,N_29433);
or UO_870 (O_870,N_29445,N_29815);
nor UO_871 (O_871,N_29504,N_29464);
nor UO_872 (O_872,N_29772,N_29485);
nand UO_873 (O_873,N_29494,N_29970);
and UO_874 (O_874,N_29659,N_29700);
and UO_875 (O_875,N_29920,N_29844);
nand UO_876 (O_876,N_29528,N_29978);
or UO_877 (O_877,N_29610,N_29768);
nand UO_878 (O_878,N_29557,N_29991);
and UO_879 (O_879,N_29440,N_29847);
nor UO_880 (O_880,N_29447,N_29481);
nand UO_881 (O_881,N_29738,N_29428);
nand UO_882 (O_882,N_29903,N_29882);
xnor UO_883 (O_883,N_29841,N_29979);
or UO_884 (O_884,N_29785,N_29836);
nand UO_885 (O_885,N_29807,N_29625);
and UO_886 (O_886,N_29846,N_29677);
and UO_887 (O_887,N_29835,N_29992);
or UO_888 (O_888,N_29541,N_29736);
xnor UO_889 (O_889,N_29466,N_29874);
nand UO_890 (O_890,N_29958,N_29826);
nand UO_891 (O_891,N_29569,N_29503);
and UO_892 (O_892,N_29795,N_29968);
or UO_893 (O_893,N_29514,N_29707);
nand UO_894 (O_894,N_29680,N_29632);
nor UO_895 (O_895,N_29707,N_29564);
xnor UO_896 (O_896,N_29827,N_29657);
and UO_897 (O_897,N_29737,N_29773);
and UO_898 (O_898,N_29710,N_29780);
nand UO_899 (O_899,N_29584,N_29769);
or UO_900 (O_900,N_29649,N_29788);
and UO_901 (O_901,N_29774,N_29698);
and UO_902 (O_902,N_29663,N_29711);
xor UO_903 (O_903,N_29435,N_29445);
nor UO_904 (O_904,N_29644,N_29676);
and UO_905 (O_905,N_29864,N_29921);
xnor UO_906 (O_906,N_29576,N_29506);
nor UO_907 (O_907,N_29492,N_29568);
nor UO_908 (O_908,N_29548,N_29513);
xor UO_909 (O_909,N_29688,N_29494);
nand UO_910 (O_910,N_29695,N_29407);
or UO_911 (O_911,N_29996,N_29505);
nand UO_912 (O_912,N_29591,N_29460);
xnor UO_913 (O_913,N_29511,N_29402);
or UO_914 (O_914,N_29516,N_29719);
nand UO_915 (O_915,N_29632,N_29998);
nand UO_916 (O_916,N_29977,N_29630);
nand UO_917 (O_917,N_29890,N_29690);
and UO_918 (O_918,N_29483,N_29762);
or UO_919 (O_919,N_29461,N_29987);
and UO_920 (O_920,N_29648,N_29912);
or UO_921 (O_921,N_29944,N_29879);
nor UO_922 (O_922,N_29404,N_29721);
nand UO_923 (O_923,N_29953,N_29765);
nand UO_924 (O_924,N_29899,N_29617);
or UO_925 (O_925,N_29628,N_29560);
nor UO_926 (O_926,N_29481,N_29456);
or UO_927 (O_927,N_29944,N_29993);
xor UO_928 (O_928,N_29468,N_29942);
and UO_929 (O_929,N_29578,N_29936);
nor UO_930 (O_930,N_29719,N_29880);
nand UO_931 (O_931,N_29698,N_29427);
nor UO_932 (O_932,N_29671,N_29831);
nand UO_933 (O_933,N_29670,N_29553);
or UO_934 (O_934,N_29991,N_29761);
or UO_935 (O_935,N_29777,N_29987);
xor UO_936 (O_936,N_29803,N_29788);
nand UO_937 (O_937,N_29515,N_29496);
or UO_938 (O_938,N_29726,N_29524);
xnor UO_939 (O_939,N_29862,N_29783);
xnor UO_940 (O_940,N_29515,N_29817);
and UO_941 (O_941,N_29490,N_29482);
or UO_942 (O_942,N_29982,N_29492);
nor UO_943 (O_943,N_29980,N_29625);
and UO_944 (O_944,N_29423,N_29844);
nand UO_945 (O_945,N_29422,N_29718);
xor UO_946 (O_946,N_29409,N_29907);
nand UO_947 (O_947,N_29791,N_29709);
nand UO_948 (O_948,N_29462,N_29447);
or UO_949 (O_949,N_29563,N_29771);
nand UO_950 (O_950,N_29865,N_29574);
and UO_951 (O_951,N_29870,N_29903);
or UO_952 (O_952,N_29978,N_29961);
and UO_953 (O_953,N_29868,N_29446);
nand UO_954 (O_954,N_29727,N_29674);
or UO_955 (O_955,N_29675,N_29530);
and UO_956 (O_956,N_29494,N_29718);
nor UO_957 (O_957,N_29404,N_29629);
or UO_958 (O_958,N_29598,N_29580);
or UO_959 (O_959,N_29595,N_29711);
or UO_960 (O_960,N_29699,N_29923);
xnor UO_961 (O_961,N_29691,N_29950);
xor UO_962 (O_962,N_29467,N_29526);
nor UO_963 (O_963,N_29578,N_29730);
and UO_964 (O_964,N_29536,N_29539);
xor UO_965 (O_965,N_29414,N_29439);
and UO_966 (O_966,N_29980,N_29740);
and UO_967 (O_967,N_29842,N_29833);
nor UO_968 (O_968,N_29553,N_29734);
nor UO_969 (O_969,N_29985,N_29861);
or UO_970 (O_970,N_29806,N_29676);
and UO_971 (O_971,N_29413,N_29776);
and UO_972 (O_972,N_29989,N_29956);
nand UO_973 (O_973,N_29884,N_29726);
or UO_974 (O_974,N_29919,N_29855);
xor UO_975 (O_975,N_29495,N_29505);
xnor UO_976 (O_976,N_29589,N_29981);
or UO_977 (O_977,N_29834,N_29707);
or UO_978 (O_978,N_29945,N_29780);
and UO_979 (O_979,N_29686,N_29999);
and UO_980 (O_980,N_29808,N_29523);
and UO_981 (O_981,N_29522,N_29974);
xnor UO_982 (O_982,N_29715,N_29622);
nor UO_983 (O_983,N_29868,N_29721);
xnor UO_984 (O_984,N_29661,N_29881);
or UO_985 (O_985,N_29775,N_29943);
nand UO_986 (O_986,N_29498,N_29924);
nor UO_987 (O_987,N_29612,N_29742);
nand UO_988 (O_988,N_29545,N_29618);
and UO_989 (O_989,N_29401,N_29849);
nor UO_990 (O_990,N_29878,N_29819);
and UO_991 (O_991,N_29573,N_29506);
xnor UO_992 (O_992,N_29906,N_29938);
nand UO_993 (O_993,N_29975,N_29920);
or UO_994 (O_994,N_29730,N_29610);
and UO_995 (O_995,N_29615,N_29423);
nand UO_996 (O_996,N_29755,N_29662);
nand UO_997 (O_997,N_29809,N_29664);
xor UO_998 (O_998,N_29467,N_29953);
nor UO_999 (O_999,N_29900,N_29976);
and UO_1000 (O_1000,N_29690,N_29551);
nor UO_1001 (O_1001,N_29709,N_29735);
nand UO_1002 (O_1002,N_29901,N_29926);
nand UO_1003 (O_1003,N_29504,N_29635);
and UO_1004 (O_1004,N_29514,N_29616);
and UO_1005 (O_1005,N_29844,N_29870);
and UO_1006 (O_1006,N_29611,N_29840);
or UO_1007 (O_1007,N_29561,N_29537);
nor UO_1008 (O_1008,N_29688,N_29668);
xor UO_1009 (O_1009,N_29633,N_29410);
xnor UO_1010 (O_1010,N_29836,N_29929);
nor UO_1011 (O_1011,N_29554,N_29451);
or UO_1012 (O_1012,N_29992,N_29661);
nor UO_1013 (O_1013,N_29919,N_29534);
nand UO_1014 (O_1014,N_29930,N_29664);
and UO_1015 (O_1015,N_29510,N_29707);
and UO_1016 (O_1016,N_29588,N_29993);
nor UO_1017 (O_1017,N_29412,N_29624);
or UO_1018 (O_1018,N_29811,N_29905);
nor UO_1019 (O_1019,N_29972,N_29967);
or UO_1020 (O_1020,N_29783,N_29904);
and UO_1021 (O_1021,N_29647,N_29788);
xnor UO_1022 (O_1022,N_29560,N_29916);
or UO_1023 (O_1023,N_29468,N_29814);
xor UO_1024 (O_1024,N_29492,N_29589);
nand UO_1025 (O_1025,N_29414,N_29484);
xnor UO_1026 (O_1026,N_29471,N_29846);
xor UO_1027 (O_1027,N_29630,N_29616);
and UO_1028 (O_1028,N_29610,N_29698);
xnor UO_1029 (O_1029,N_29543,N_29451);
or UO_1030 (O_1030,N_29756,N_29550);
or UO_1031 (O_1031,N_29461,N_29471);
xnor UO_1032 (O_1032,N_29775,N_29842);
nand UO_1033 (O_1033,N_29965,N_29681);
xor UO_1034 (O_1034,N_29420,N_29523);
and UO_1035 (O_1035,N_29426,N_29825);
and UO_1036 (O_1036,N_29624,N_29605);
nor UO_1037 (O_1037,N_29888,N_29882);
and UO_1038 (O_1038,N_29400,N_29536);
or UO_1039 (O_1039,N_29493,N_29991);
or UO_1040 (O_1040,N_29740,N_29914);
xor UO_1041 (O_1041,N_29937,N_29552);
nor UO_1042 (O_1042,N_29900,N_29682);
nor UO_1043 (O_1043,N_29410,N_29769);
xnor UO_1044 (O_1044,N_29581,N_29856);
xor UO_1045 (O_1045,N_29508,N_29625);
and UO_1046 (O_1046,N_29797,N_29449);
nand UO_1047 (O_1047,N_29848,N_29475);
or UO_1048 (O_1048,N_29839,N_29940);
xnor UO_1049 (O_1049,N_29826,N_29970);
nor UO_1050 (O_1050,N_29881,N_29913);
nor UO_1051 (O_1051,N_29703,N_29683);
xor UO_1052 (O_1052,N_29968,N_29454);
xor UO_1053 (O_1053,N_29936,N_29754);
nand UO_1054 (O_1054,N_29475,N_29882);
and UO_1055 (O_1055,N_29718,N_29701);
nor UO_1056 (O_1056,N_29600,N_29466);
and UO_1057 (O_1057,N_29759,N_29997);
xnor UO_1058 (O_1058,N_29717,N_29965);
and UO_1059 (O_1059,N_29693,N_29657);
and UO_1060 (O_1060,N_29981,N_29845);
nor UO_1061 (O_1061,N_29640,N_29457);
or UO_1062 (O_1062,N_29725,N_29596);
or UO_1063 (O_1063,N_29571,N_29680);
nor UO_1064 (O_1064,N_29610,N_29870);
nand UO_1065 (O_1065,N_29744,N_29895);
xor UO_1066 (O_1066,N_29829,N_29844);
or UO_1067 (O_1067,N_29791,N_29532);
nand UO_1068 (O_1068,N_29811,N_29458);
xnor UO_1069 (O_1069,N_29559,N_29796);
nand UO_1070 (O_1070,N_29412,N_29926);
or UO_1071 (O_1071,N_29810,N_29478);
nand UO_1072 (O_1072,N_29720,N_29764);
and UO_1073 (O_1073,N_29891,N_29642);
xor UO_1074 (O_1074,N_29666,N_29935);
and UO_1075 (O_1075,N_29801,N_29943);
nor UO_1076 (O_1076,N_29466,N_29854);
nand UO_1077 (O_1077,N_29689,N_29493);
and UO_1078 (O_1078,N_29882,N_29405);
or UO_1079 (O_1079,N_29558,N_29657);
nand UO_1080 (O_1080,N_29942,N_29529);
nand UO_1081 (O_1081,N_29665,N_29420);
nor UO_1082 (O_1082,N_29459,N_29903);
nor UO_1083 (O_1083,N_29946,N_29875);
xor UO_1084 (O_1084,N_29963,N_29943);
or UO_1085 (O_1085,N_29955,N_29993);
or UO_1086 (O_1086,N_29735,N_29794);
or UO_1087 (O_1087,N_29974,N_29538);
xnor UO_1088 (O_1088,N_29548,N_29825);
nor UO_1089 (O_1089,N_29609,N_29532);
nand UO_1090 (O_1090,N_29764,N_29950);
or UO_1091 (O_1091,N_29769,N_29648);
xor UO_1092 (O_1092,N_29632,N_29525);
or UO_1093 (O_1093,N_29420,N_29966);
nand UO_1094 (O_1094,N_29501,N_29866);
and UO_1095 (O_1095,N_29553,N_29748);
and UO_1096 (O_1096,N_29489,N_29732);
or UO_1097 (O_1097,N_29893,N_29806);
nor UO_1098 (O_1098,N_29410,N_29439);
or UO_1099 (O_1099,N_29956,N_29825);
nand UO_1100 (O_1100,N_29408,N_29875);
or UO_1101 (O_1101,N_29757,N_29581);
nand UO_1102 (O_1102,N_29732,N_29929);
and UO_1103 (O_1103,N_29827,N_29877);
xnor UO_1104 (O_1104,N_29776,N_29497);
or UO_1105 (O_1105,N_29889,N_29726);
nor UO_1106 (O_1106,N_29527,N_29894);
and UO_1107 (O_1107,N_29561,N_29845);
and UO_1108 (O_1108,N_29668,N_29857);
nand UO_1109 (O_1109,N_29752,N_29680);
nor UO_1110 (O_1110,N_29431,N_29543);
nor UO_1111 (O_1111,N_29777,N_29717);
xnor UO_1112 (O_1112,N_29525,N_29535);
nand UO_1113 (O_1113,N_29512,N_29616);
or UO_1114 (O_1114,N_29470,N_29896);
xnor UO_1115 (O_1115,N_29955,N_29417);
nor UO_1116 (O_1116,N_29445,N_29522);
or UO_1117 (O_1117,N_29710,N_29814);
or UO_1118 (O_1118,N_29770,N_29971);
nor UO_1119 (O_1119,N_29508,N_29769);
xnor UO_1120 (O_1120,N_29787,N_29510);
or UO_1121 (O_1121,N_29487,N_29516);
and UO_1122 (O_1122,N_29668,N_29574);
nand UO_1123 (O_1123,N_29973,N_29810);
and UO_1124 (O_1124,N_29864,N_29723);
nand UO_1125 (O_1125,N_29917,N_29441);
nand UO_1126 (O_1126,N_29474,N_29802);
xor UO_1127 (O_1127,N_29660,N_29532);
and UO_1128 (O_1128,N_29933,N_29876);
and UO_1129 (O_1129,N_29527,N_29758);
or UO_1130 (O_1130,N_29914,N_29959);
nand UO_1131 (O_1131,N_29991,N_29671);
and UO_1132 (O_1132,N_29426,N_29660);
nor UO_1133 (O_1133,N_29514,N_29434);
nor UO_1134 (O_1134,N_29968,N_29676);
or UO_1135 (O_1135,N_29691,N_29981);
or UO_1136 (O_1136,N_29500,N_29443);
nand UO_1137 (O_1137,N_29493,N_29710);
nor UO_1138 (O_1138,N_29926,N_29456);
or UO_1139 (O_1139,N_29800,N_29793);
nand UO_1140 (O_1140,N_29712,N_29928);
nor UO_1141 (O_1141,N_29614,N_29784);
xor UO_1142 (O_1142,N_29767,N_29986);
nand UO_1143 (O_1143,N_29497,N_29756);
xor UO_1144 (O_1144,N_29688,N_29611);
and UO_1145 (O_1145,N_29793,N_29638);
nand UO_1146 (O_1146,N_29646,N_29799);
xnor UO_1147 (O_1147,N_29577,N_29660);
nor UO_1148 (O_1148,N_29474,N_29788);
or UO_1149 (O_1149,N_29929,N_29866);
nor UO_1150 (O_1150,N_29616,N_29720);
and UO_1151 (O_1151,N_29723,N_29415);
and UO_1152 (O_1152,N_29425,N_29801);
xnor UO_1153 (O_1153,N_29974,N_29882);
nand UO_1154 (O_1154,N_29767,N_29575);
and UO_1155 (O_1155,N_29448,N_29662);
and UO_1156 (O_1156,N_29499,N_29746);
nand UO_1157 (O_1157,N_29605,N_29985);
and UO_1158 (O_1158,N_29406,N_29834);
xnor UO_1159 (O_1159,N_29799,N_29667);
xnor UO_1160 (O_1160,N_29995,N_29763);
nor UO_1161 (O_1161,N_29570,N_29808);
nand UO_1162 (O_1162,N_29532,N_29655);
nand UO_1163 (O_1163,N_29464,N_29929);
nand UO_1164 (O_1164,N_29596,N_29877);
nand UO_1165 (O_1165,N_29753,N_29554);
nand UO_1166 (O_1166,N_29741,N_29993);
nand UO_1167 (O_1167,N_29574,N_29759);
nor UO_1168 (O_1168,N_29595,N_29636);
nand UO_1169 (O_1169,N_29994,N_29413);
or UO_1170 (O_1170,N_29872,N_29817);
or UO_1171 (O_1171,N_29805,N_29713);
nor UO_1172 (O_1172,N_29933,N_29520);
nand UO_1173 (O_1173,N_29449,N_29858);
nand UO_1174 (O_1174,N_29980,N_29519);
and UO_1175 (O_1175,N_29983,N_29619);
or UO_1176 (O_1176,N_29797,N_29860);
xnor UO_1177 (O_1177,N_29417,N_29477);
or UO_1178 (O_1178,N_29790,N_29624);
and UO_1179 (O_1179,N_29848,N_29904);
and UO_1180 (O_1180,N_29587,N_29570);
and UO_1181 (O_1181,N_29716,N_29979);
xor UO_1182 (O_1182,N_29996,N_29913);
and UO_1183 (O_1183,N_29602,N_29489);
or UO_1184 (O_1184,N_29842,N_29468);
and UO_1185 (O_1185,N_29457,N_29824);
nor UO_1186 (O_1186,N_29970,N_29435);
and UO_1187 (O_1187,N_29690,N_29513);
and UO_1188 (O_1188,N_29741,N_29745);
nor UO_1189 (O_1189,N_29640,N_29976);
and UO_1190 (O_1190,N_29408,N_29995);
and UO_1191 (O_1191,N_29550,N_29541);
and UO_1192 (O_1192,N_29424,N_29832);
xor UO_1193 (O_1193,N_29485,N_29537);
and UO_1194 (O_1194,N_29547,N_29787);
nor UO_1195 (O_1195,N_29591,N_29798);
xor UO_1196 (O_1196,N_29705,N_29693);
and UO_1197 (O_1197,N_29764,N_29887);
nand UO_1198 (O_1198,N_29459,N_29406);
xor UO_1199 (O_1199,N_29777,N_29720);
nor UO_1200 (O_1200,N_29685,N_29850);
nor UO_1201 (O_1201,N_29489,N_29755);
or UO_1202 (O_1202,N_29684,N_29758);
or UO_1203 (O_1203,N_29737,N_29503);
xor UO_1204 (O_1204,N_29744,N_29806);
nand UO_1205 (O_1205,N_29735,N_29644);
nor UO_1206 (O_1206,N_29447,N_29785);
nand UO_1207 (O_1207,N_29850,N_29955);
and UO_1208 (O_1208,N_29891,N_29485);
and UO_1209 (O_1209,N_29554,N_29525);
or UO_1210 (O_1210,N_29532,N_29917);
nand UO_1211 (O_1211,N_29576,N_29514);
nand UO_1212 (O_1212,N_29858,N_29838);
or UO_1213 (O_1213,N_29736,N_29873);
xnor UO_1214 (O_1214,N_29508,N_29807);
nor UO_1215 (O_1215,N_29453,N_29468);
xnor UO_1216 (O_1216,N_29629,N_29852);
and UO_1217 (O_1217,N_29512,N_29961);
or UO_1218 (O_1218,N_29713,N_29894);
nand UO_1219 (O_1219,N_29934,N_29979);
and UO_1220 (O_1220,N_29793,N_29879);
xnor UO_1221 (O_1221,N_29943,N_29718);
and UO_1222 (O_1222,N_29513,N_29542);
or UO_1223 (O_1223,N_29579,N_29818);
or UO_1224 (O_1224,N_29793,N_29861);
or UO_1225 (O_1225,N_29716,N_29577);
or UO_1226 (O_1226,N_29572,N_29609);
xnor UO_1227 (O_1227,N_29503,N_29516);
nand UO_1228 (O_1228,N_29457,N_29797);
nor UO_1229 (O_1229,N_29487,N_29901);
xor UO_1230 (O_1230,N_29990,N_29553);
xnor UO_1231 (O_1231,N_29804,N_29544);
and UO_1232 (O_1232,N_29470,N_29587);
nor UO_1233 (O_1233,N_29877,N_29811);
xnor UO_1234 (O_1234,N_29438,N_29822);
or UO_1235 (O_1235,N_29468,N_29434);
nor UO_1236 (O_1236,N_29412,N_29567);
or UO_1237 (O_1237,N_29819,N_29871);
or UO_1238 (O_1238,N_29920,N_29522);
nor UO_1239 (O_1239,N_29914,N_29984);
or UO_1240 (O_1240,N_29943,N_29831);
xor UO_1241 (O_1241,N_29725,N_29468);
or UO_1242 (O_1242,N_29868,N_29814);
nor UO_1243 (O_1243,N_29681,N_29457);
nand UO_1244 (O_1244,N_29462,N_29911);
xnor UO_1245 (O_1245,N_29936,N_29473);
xnor UO_1246 (O_1246,N_29998,N_29930);
nand UO_1247 (O_1247,N_29689,N_29492);
and UO_1248 (O_1248,N_29513,N_29448);
nand UO_1249 (O_1249,N_29554,N_29958);
and UO_1250 (O_1250,N_29986,N_29989);
xnor UO_1251 (O_1251,N_29927,N_29998);
xnor UO_1252 (O_1252,N_29777,N_29850);
and UO_1253 (O_1253,N_29889,N_29830);
or UO_1254 (O_1254,N_29572,N_29626);
or UO_1255 (O_1255,N_29783,N_29930);
nand UO_1256 (O_1256,N_29767,N_29446);
nand UO_1257 (O_1257,N_29718,N_29416);
nand UO_1258 (O_1258,N_29590,N_29791);
nand UO_1259 (O_1259,N_29551,N_29854);
and UO_1260 (O_1260,N_29825,N_29949);
or UO_1261 (O_1261,N_29689,N_29723);
and UO_1262 (O_1262,N_29402,N_29649);
or UO_1263 (O_1263,N_29658,N_29699);
nor UO_1264 (O_1264,N_29936,N_29997);
xor UO_1265 (O_1265,N_29567,N_29542);
xor UO_1266 (O_1266,N_29826,N_29944);
nor UO_1267 (O_1267,N_29885,N_29967);
or UO_1268 (O_1268,N_29896,N_29942);
and UO_1269 (O_1269,N_29776,N_29694);
and UO_1270 (O_1270,N_29913,N_29442);
xor UO_1271 (O_1271,N_29734,N_29911);
or UO_1272 (O_1272,N_29775,N_29814);
xnor UO_1273 (O_1273,N_29675,N_29623);
xor UO_1274 (O_1274,N_29410,N_29831);
nand UO_1275 (O_1275,N_29446,N_29591);
xor UO_1276 (O_1276,N_29459,N_29411);
and UO_1277 (O_1277,N_29864,N_29619);
nand UO_1278 (O_1278,N_29594,N_29894);
nor UO_1279 (O_1279,N_29876,N_29645);
and UO_1280 (O_1280,N_29894,N_29935);
and UO_1281 (O_1281,N_29635,N_29800);
and UO_1282 (O_1282,N_29523,N_29680);
nand UO_1283 (O_1283,N_29775,N_29993);
and UO_1284 (O_1284,N_29795,N_29574);
nand UO_1285 (O_1285,N_29553,N_29837);
nor UO_1286 (O_1286,N_29413,N_29722);
and UO_1287 (O_1287,N_29617,N_29692);
nor UO_1288 (O_1288,N_29666,N_29591);
nand UO_1289 (O_1289,N_29476,N_29520);
or UO_1290 (O_1290,N_29946,N_29794);
and UO_1291 (O_1291,N_29901,N_29921);
and UO_1292 (O_1292,N_29947,N_29424);
and UO_1293 (O_1293,N_29800,N_29657);
and UO_1294 (O_1294,N_29994,N_29880);
xnor UO_1295 (O_1295,N_29965,N_29777);
nand UO_1296 (O_1296,N_29413,N_29500);
and UO_1297 (O_1297,N_29842,N_29973);
nand UO_1298 (O_1298,N_29496,N_29905);
nor UO_1299 (O_1299,N_29569,N_29675);
nor UO_1300 (O_1300,N_29991,N_29614);
nor UO_1301 (O_1301,N_29540,N_29895);
and UO_1302 (O_1302,N_29559,N_29986);
nor UO_1303 (O_1303,N_29994,N_29682);
and UO_1304 (O_1304,N_29857,N_29578);
or UO_1305 (O_1305,N_29674,N_29997);
xnor UO_1306 (O_1306,N_29557,N_29465);
nor UO_1307 (O_1307,N_29979,N_29896);
xor UO_1308 (O_1308,N_29638,N_29537);
xor UO_1309 (O_1309,N_29454,N_29604);
or UO_1310 (O_1310,N_29809,N_29691);
or UO_1311 (O_1311,N_29771,N_29854);
nor UO_1312 (O_1312,N_29729,N_29660);
nand UO_1313 (O_1313,N_29469,N_29891);
xor UO_1314 (O_1314,N_29849,N_29891);
and UO_1315 (O_1315,N_29822,N_29540);
xor UO_1316 (O_1316,N_29422,N_29664);
or UO_1317 (O_1317,N_29968,N_29757);
nand UO_1318 (O_1318,N_29568,N_29878);
or UO_1319 (O_1319,N_29499,N_29542);
xor UO_1320 (O_1320,N_29594,N_29770);
and UO_1321 (O_1321,N_29579,N_29471);
or UO_1322 (O_1322,N_29404,N_29756);
nand UO_1323 (O_1323,N_29842,N_29800);
and UO_1324 (O_1324,N_29751,N_29745);
nor UO_1325 (O_1325,N_29736,N_29828);
and UO_1326 (O_1326,N_29949,N_29736);
xor UO_1327 (O_1327,N_29637,N_29898);
or UO_1328 (O_1328,N_29986,N_29756);
xnor UO_1329 (O_1329,N_29604,N_29891);
nand UO_1330 (O_1330,N_29598,N_29619);
and UO_1331 (O_1331,N_29768,N_29753);
nor UO_1332 (O_1332,N_29552,N_29900);
or UO_1333 (O_1333,N_29919,N_29921);
or UO_1334 (O_1334,N_29495,N_29536);
nor UO_1335 (O_1335,N_29412,N_29850);
and UO_1336 (O_1336,N_29587,N_29968);
nor UO_1337 (O_1337,N_29486,N_29553);
or UO_1338 (O_1338,N_29404,N_29528);
and UO_1339 (O_1339,N_29430,N_29871);
nor UO_1340 (O_1340,N_29811,N_29568);
or UO_1341 (O_1341,N_29954,N_29597);
nor UO_1342 (O_1342,N_29664,N_29406);
xor UO_1343 (O_1343,N_29479,N_29483);
nor UO_1344 (O_1344,N_29854,N_29665);
and UO_1345 (O_1345,N_29410,N_29912);
nor UO_1346 (O_1346,N_29780,N_29433);
nand UO_1347 (O_1347,N_29514,N_29494);
or UO_1348 (O_1348,N_29484,N_29952);
nand UO_1349 (O_1349,N_29615,N_29544);
nor UO_1350 (O_1350,N_29471,N_29510);
and UO_1351 (O_1351,N_29449,N_29585);
nand UO_1352 (O_1352,N_29738,N_29657);
nand UO_1353 (O_1353,N_29625,N_29536);
or UO_1354 (O_1354,N_29511,N_29679);
or UO_1355 (O_1355,N_29427,N_29914);
or UO_1356 (O_1356,N_29898,N_29877);
xor UO_1357 (O_1357,N_29758,N_29931);
nand UO_1358 (O_1358,N_29416,N_29415);
xor UO_1359 (O_1359,N_29691,N_29689);
and UO_1360 (O_1360,N_29639,N_29862);
nor UO_1361 (O_1361,N_29764,N_29951);
nand UO_1362 (O_1362,N_29952,N_29428);
and UO_1363 (O_1363,N_29870,N_29531);
nor UO_1364 (O_1364,N_29697,N_29608);
xnor UO_1365 (O_1365,N_29466,N_29542);
nand UO_1366 (O_1366,N_29416,N_29496);
nand UO_1367 (O_1367,N_29419,N_29534);
nand UO_1368 (O_1368,N_29528,N_29409);
or UO_1369 (O_1369,N_29754,N_29854);
or UO_1370 (O_1370,N_29583,N_29857);
or UO_1371 (O_1371,N_29541,N_29639);
xnor UO_1372 (O_1372,N_29774,N_29463);
and UO_1373 (O_1373,N_29642,N_29864);
and UO_1374 (O_1374,N_29986,N_29795);
nand UO_1375 (O_1375,N_29839,N_29740);
or UO_1376 (O_1376,N_29500,N_29415);
and UO_1377 (O_1377,N_29960,N_29811);
or UO_1378 (O_1378,N_29478,N_29794);
nor UO_1379 (O_1379,N_29968,N_29481);
and UO_1380 (O_1380,N_29520,N_29470);
xor UO_1381 (O_1381,N_29481,N_29641);
nand UO_1382 (O_1382,N_29995,N_29936);
nor UO_1383 (O_1383,N_29603,N_29831);
xnor UO_1384 (O_1384,N_29817,N_29629);
xnor UO_1385 (O_1385,N_29569,N_29416);
or UO_1386 (O_1386,N_29685,N_29865);
and UO_1387 (O_1387,N_29712,N_29580);
nand UO_1388 (O_1388,N_29982,N_29924);
and UO_1389 (O_1389,N_29709,N_29649);
or UO_1390 (O_1390,N_29788,N_29607);
xnor UO_1391 (O_1391,N_29946,N_29950);
xnor UO_1392 (O_1392,N_29598,N_29927);
and UO_1393 (O_1393,N_29951,N_29750);
nand UO_1394 (O_1394,N_29880,N_29662);
or UO_1395 (O_1395,N_29827,N_29517);
xor UO_1396 (O_1396,N_29466,N_29865);
nand UO_1397 (O_1397,N_29594,N_29426);
and UO_1398 (O_1398,N_29949,N_29620);
nand UO_1399 (O_1399,N_29552,N_29454);
or UO_1400 (O_1400,N_29839,N_29643);
and UO_1401 (O_1401,N_29669,N_29634);
nor UO_1402 (O_1402,N_29911,N_29425);
and UO_1403 (O_1403,N_29743,N_29967);
nand UO_1404 (O_1404,N_29908,N_29755);
nand UO_1405 (O_1405,N_29499,N_29898);
nand UO_1406 (O_1406,N_29414,N_29923);
xor UO_1407 (O_1407,N_29414,N_29927);
or UO_1408 (O_1408,N_29574,N_29812);
nor UO_1409 (O_1409,N_29421,N_29809);
and UO_1410 (O_1410,N_29719,N_29639);
xor UO_1411 (O_1411,N_29526,N_29869);
xor UO_1412 (O_1412,N_29700,N_29695);
xnor UO_1413 (O_1413,N_29604,N_29739);
nor UO_1414 (O_1414,N_29458,N_29496);
nor UO_1415 (O_1415,N_29740,N_29922);
or UO_1416 (O_1416,N_29943,N_29603);
xor UO_1417 (O_1417,N_29960,N_29493);
nand UO_1418 (O_1418,N_29554,N_29702);
or UO_1419 (O_1419,N_29750,N_29557);
xor UO_1420 (O_1420,N_29641,N_29964);
nand UO_1421 (O_1421,N_29672,N_29639);
or UO_1422 (O_1422,N_29912,N_29683);
nand UO_1423 (O_1423,N_29768,N_29618);
and UO_1424 (O_1424,N_29990,N_29427);
xor UO_1425 (O_1425,N_29831,N_29800);
nand UO_1426 (O_1426,N_29447,N_29506);
xnor UO_1427 (O_1427,N_29709,N_29514);
and UO_1428 (O_1428,N_29905,N_29732);
or UO_1429 (O_1429,N_29846,N_29786);
and UO_1430 (O_1430,N_29614,N_29970);
and UO_1431 (O_1431,N_29715,N_29864);
and UO_1432 (O_1432,N_29789,N_29573);
nand UO_1433 (O_1433,N_29988,N_29438);
nand UO_1434 (O_1434,N_29402,N_29420);
xnor UO_1435 (O_1435,N_29927,N_29530);
or UO_1436 (O_1436,N_29414,N_29837);
xnor UO_1437 (O_1437,N_29563,N_29773);
and UO_1438 (O_1438,N_29634,N_29868);
and UO_1439 (O_1439,N_29877,N_29656);
or UO_1440 (O_1440,N_29512,N_29999);
nor UO_1441 (O_1441,N_29661,N_29788);
nand UO_1442 (O_1442,N_29566,N_29685);
or UO_1443 (O_1443,N_29838,N_29418);
nand UO_1444 (O_1444,N_29448,N_29630);
nor UO_1445 (O_1445,N_29972,N_29535);
and UO_1446 (O_1446,N_29982,N_29669);
xor UO_1447 (O_1447,N_29546,N_29996);
or UO_1448 (O_1448,N_29771,N_29418);
and UO_1449 (O_1449,N_29454,N_29708);
nor UO_1450 (O_1450,N_29904,N_29769);
and UO_1451 (O_1451,N_29427,N_29632);
and UO_1452 (O_1452,N_29603,N_29437);
nor UO_1453 (O_1453,N_29577,N_29624);
nor UO_1454 (O_1454,N_29958,N_29775);
nand UO_1455 (O_1455,N_29728,N_29649);
and UO_1456 (O_1456,N_29892,N_29579);
xnor UO_1457 (O_1457,N_29928,N_29970);
or UO_1458 (O_1458,N_29976,N_29751);
nor UO_1459 (O_1459,N_29888,N_29728);
xnor UO_1460 (O_1460,N_29980,N_29895);
nand UO_1461 (O_1461,N_29569,N_29686);
nand UO_1462 (O_1462,N_29730,N_29881);
or UO_1463 (O_1463,N_29467,N_29610);
xnor UO_1464 (O_1464,N_29803,N_29862);
nand UO_1465 (O_1465,N_29921,N_29480);
nand UO_1466 (O_1466,N_29806,N_29865);
or UO_1467 (O_1467,N_29579,N_29470);
xor UO_1468 (O_1468,N_29416,N_29731);
nor UO_1469 (O_1469,N_29865,N_29711);
nor UO_1470 (O_1470,N_29583,N_29489);
or UO_1471 (O_1471,N_29485,N_29732);
xor UO_1472 (O_1472,N_29448,N_29693);
and UO_1473 (O_1473,N_29621,N_29598);
nand UO_1474 (O_1474,N_29512,N_29564);
xnor UO_1475 (O_1475,N_29935,N_29855);
and UO_1476 (O_1476,N_29584,N_29710);
or UO_1477 (O_1477,N_29834,N_29541);
or UO_1478 (O_1478,N_29466,N_29471);
nor UO_1479 (O_1479,N_29567,N_29773);
nor UO_1480 (O_1480,N_29509,N_29405);
or UO_1481 (O_1481,N_29670,N_29920);
or UO_1482 (O_1482,N_29607,N_29782);
or UO_1483 (O_1483,N_29681,N_29714);
nand UO_1484 (O_1484,N_29597,N_29460);
xnor UO_1485 (O_1485,N_29712,N_29516);
or UO_1486 (O_1486,N_29586,N_29748);
xnor UO_1487 (O_1487,N_29958,N_29922);
xor UO_1488 (O_1488,N_29667,N_29942);
or UO_1489 (O_1489,N_29458,N_29751);
and UO_1490 (O_1490,N_29469,N_29921);
nor UO_1491 (O_1491,N_29685,N_29963);
nor UO_1492 (O_1492,N_29794,N_29835);
nand UO_1493 (O_1493,N_29802,N_29691);
or UO_1494 (O_1494,N_29764,N_29832);
nand UO_1495 (O_1495,N_29682,N_29730);
and UO_1496 (O_1496,N_29575,N_29934);
and UO_1497 (O_1497,N_29411,N_29437);
xor UO_1498 (O_1498,N_29761,N_29503);
xnor UO_1499 (O_1499,N_29690,N_29830);
nor UO_1500 (O_1500,N_29626,N_29852);
xnor UO_1501 (O_1501,N_29918,N_29949);
xnor UO_1502 (O_1502,N_29513,N_29601);
nand UO_1503 (O_1503,N_29913,N_29919);
nor UO_1504 (O_1504,N_29818,N_29421);
xnor UO_1505 (O_1505,N_29836,N_29684);
or UO_1506 (O_1506,N_29601,N_29831);
nand UO_1507 (O_1507,N_29802,N_29517);
nand UO_1508 (O_1508,N_29412,N_29431);
nand UO_1509 (O_1509,N_29799,N_29480);
xnor UO_1510 (O_1510,N_29677,N_29453);
and UO_1511 (O_1511,N_29808,N_29757);
xor UO_1512 (O_1512,N_29925,N_29949);
or UO_1513 (O_1513,N_29607,N_29719);
or UO_1514 (O_1514,N_29443,N_29664);
nand UO_1515 (O_1515,N_29499,N_29427);
nor UO_1516 (O_1516,N_29715,N_29797);
xor UO_1517 (O_1517,N_29777,N_29773);
and UO_1518 (O_1518,N_29669,N_29679);
or UO_1519 (O_1519,N_29723,N_29874);
nand UO_1520 (O_1520,N_29474,N_29910);
nand UO_1521 (O_1521,N_29936,N_29410);
nand UO_1522 (O_1522,N_29841,N_29568);
nand UO_1523 (O_1523,N_29709,N_29794);
nand UO_1524 (O_1524,N_29421,N_29644);
nand UO_1525 (O_1525,N_29562,N_29747);
and UO_1526 (O_1526,N_29950,N_29769);
and UO_1527 (O_1527,N_29747,N_29649);
nor UO_1528 (O_1528,N_29581,N_29738);
and UO_1529 (O_1529,N_29691,N_29511);
xnor UO_1530 (O_1530,N_29495,N_29621);
or UO_1531 (O_1531,N_29876,N_29596);
nand UO_1532 (O_1532,N_29469,N_29411);
nand UO_1533 (O_1533,N_29646,N_29755);
and UO_1534 (O_1534,N_29784,N_29534);
and UO_1535 (O_1535,N_29813,N_29482);
or UO_1536 (O_1536,N_29776,N_29454);
xnor UO_1537 (O_1537,N_29539,N_29684);
nand UO_1538 (O_1538,N_29547,N_29429);
and UO_1539 (O_1539,N_29971,N_29690);
or UO_1540 (O_1540,N_29869,N_29782);
xnor UO_1541 (O_1541,N_29875,N_29823);
nor UO_1542 (O_1542,N_29923,N_29806);
or UO_1543 (O_1543,N_29438,N_29775);
nor UO_1544 (O_1544,N_29640,N_29429);
xnor UO_1545 (O_1545,N_29499,N_29789);
xnor UO_1546 (O_1546,N_29933,N_29801);
nand UO_1547 (O_1547,N_29441,N_29913);
nor UO_1548 (O_1548,N_29863,N_29534);
and UO_1549 (O_1549,N_29712,N_29477);
nor UO_1550 (O_1550,N_29520,N_29648);
nand UO_1551 (O_1551,N_29590,N_29983);
nor UO_1552 (O_1552,N_29687,N_29668);
and UO_1553 (O_1553,N_29970,N_29621);
nand UO_1554 (O_1554,N_29495,N_29946);
nand UO_1555 (O_1555,N_29625,N_29687);
and UO_1556 (O_1556,N_29860,N_29573);
xor UO_1557 (O_1557,N_29996,N_29871);
xnor UO_1558 (O_1558,N_29571,N_29632);
or UO_1559 (O_1559,N_29558,N_29743);
or UO_1560 (O_1560,N_29499,N_29484);
xnor UO_1561 (O_1561,N_29839,N_29921);
nor UO_1562 (O_1562,N_29958,N_29649);
xnor UO_1563 (O_1563,N_29864,N_29926);
nor UO_1564 (O_1564,N_29516,N_29701);
or UO_1565 (O_1565,N_29823,N_29614);
or UO_1566 (O_1566,N_29527,N_29425);
or UO_1567 (O_1567,N_29608,N_29542);
xnor UO_1568 (O_1568,N_29465,N_29747);
or UO_1569 (O_1569,N_29620,N_29869);
nor UO_1570 (O_1570,N_29622,N_29703);
nor UO_1571 (O_1571,N_29758,N_29712);
xor UO_1572 (O_1572,N_29688,N_29407);
nand UO_1573 (O_1573,N_29757,N_29724);
nor UO_1574 (O_1574,N_29630,N_29836);
xnor UO_1575 (O_1575,N_29693,N_29894);
xnor UO_1576 (O_1576,N_29782,N_29954);
xor UO_1577 (O_1577,N_29916,N_29783);
nand UO_1578 (O_1578,N_29966,N_29457);
or UO_1579 (O_1579,N_29424,N_29582);
nand UO_1580 (O_1580,N_29641,N_29892);
xnor UO_1581 (O_1581,N_29747,N_29915);
xnor UO_1582 (O_1582,N_29826,N_29803);
or UO_1583 (O_1583,N_29516,N_29525);
xor UO_1584 (O_1584,N_29963,N_29997);
or UO_1585 (O_1585,N_29410,N_29513);
nor UO_1586 (O_1586,N_29814,N_29498);
or UO_1587 (O_1587,N_29866,N_29432);
or UO_1588 (O_1588,N_29435,N_29791);
or UO_1589 (O_1589,N_29895,N_29707);
nor UO_1590 (O_1590,N_29471,N_29581);
xnor UO_1591 (O_1591,N_29558,N_29856);
nand UO_1592 (O_1592,N_29403,N_29966);
or UO_1593 (O_1593,N_29806,N_29862);
nor UO_1594 (O_1594,N_29611,N_29436);
nand UO_1595 (O_1595,N_29901,N_29714);
and UO_1596 (O_1596,N_29502,N_29415);
nor UO_1597 (O_1597,N_29886,N_29967);
nor UO_1598 (O_1598,N_29643,N_29618);
and UO_1599 (O_1599,N_29954,N_29512);
nand UO_1600 (O_1600,N_29531,N_29981);
and UO_1601 (O_1601,N_29922,N_29496);
or UO_1602 (O_1602,N_29634,N_29544);
and UO_1603 (O_1603,N_29630,N_29988);
xnor UO_1604 (O_1604,N_29876,N_29700);
or UO_1605 (O_1605,N_29464,N_29603);
xnor UO_1606 (O_1606,N_29473,N_29757);
xor UO_1607 (O_1607,N_29872,N_29937);
xor UO_1608 (O_1608,N_29714,N_29657);
or UO_1609 (O_1609,N_29606,N_29717);
nor UO_1610 (O_1610,N_29570,N_29555);
nor UO_1611 (O_1611,N_29765,N_29526);
xor UO_1612 (O_1612,N_29925,N_29785);
or UO_1613 (O_1613,N_29981,N_29718);
or UO_1614 (O_1614,N_29855,N_29557);
nor UO_1615 (O_1615,N_29960,N_29877);
or UO_1616 (O_1616,N_29477,N_29590);
and UO_1617 (O_1617,N_29414,N_29794);
nand UO_1618 (O_1618,N_29876,N_29966);
nand UO_1619 (O_1619,N_29746,N_29626);
or UO_1620 (O_1620,N_29776,N_29689);
or UO_1621 (O_1621,N_29597,N_29773);
nand UO_1622 (O_1622,N_29868,N_29763);
nor UO_1623 (O_1623,N_29479,N_29750);
and UO_1624 (O_1624,N_29471,N_29938);
nor UO_1625 (O_1625,N_29424,N_29750);
and UO_1626 (O_1626,N_29429,N_29471);
xnor UO_1627 (O_1627,N_29763,N_29838);
nand UO_1628 (O_1628,N_29779,N_29771);
and UO_1629 (O_1629,N_29428,N_29996);
nand UO_1630 (O_1630,N_29891,N_29657);
xnor UO_1631 (O_1631,N_29441,N_29487);
nor UO_1632 (O_1632,N_29940,N_29948);
and UO_1633 (O_1633,N_29693,N_29908);
xnor UO_1634 (O_1634,N_29958,N_29691);
or UO_1635 (O_1635,N_29599,N_29705);
and UO_1636 (O_1636,N_29804,N_29604);
xnor UO_1637 (O_1637,N_29823,N_29719);
nor UO_1638 (O_1638,N_29675,N_29920);
or UO_1639 (O_1639,N_29676,N_29712);
nor UO_1640 (O_1640,N_29688,N_29681);
nand UO_1641 (O_1641,N_29435,N_29964);
and UO_1642 (O_1642,N_29866,N_29430);
or UO_1643 (O_1643,N_29503,N_29426);
and UO_1644 (O_1644,N_29591,N_29777);
or UO_1645 (O_1645,N_29969,N_29464);
and UO_1646 (O_1646,N_29649,N_29587);
or UO_1647 (O_1647,N_29993,N_29723);
and UO_1648 (O_1648,N_29656,N_29709);
xnor UO_1649 (O_1649,N_29749,N_29491);
or UO_1650 (O_1650,N_29479,N_29901);
or UO_1651 (O_1651,N_29504,N_29571);
nand UO_1652 (O_1652,N_29558,N_29735);
nand UO_1653 (O_1653,N_29479,N_29584);
or UO_1654 (O_1654,N_29787,N_29620);
nor UO_1655 (O_1655,N_29755,N_29976);
nand UO_1656 (O_1656,N_29809,N_29984);
nand UO_1657 (O_1657,N_29578,N_29697);
and UO_1658 (O_1658,N_29669,N_29689);
nor UO_1659 (O_1659,N_29903,N_29779);
nand UO_1660 (O_1660,N_29748,N_29428);
nor UO_1661 (O_1661,N_29823,N_29779);
nor UO_1662 (O_1662,N_29644,N_29581);
xor UO_1663 (O_1663,N_29659,N_29715);
or UO_1664 (O_1664,N_29530,N_29700);
nand UO_1665 (O_1665,N_29411,N_29666);
nor UO_1666 (O_1666,N_29742,N_29433);
or UO_1667 (O_1667,N_29737,N_29548);
and UO_1668 (O_1668,N_29527,N_29497);
xor UO_1669 (O_1669,N_29675,N_29490);
xor UO_1670 (O_1670,N_29943,N_29475);
or UO_1671 (O_1671,N_29773,N_29634);
and UO_1672 (O_1672,N_29755,N_29536);
nand UO_1673 (O_1673,N_29988,N_29587);
nand UO_1674 (O_1674,N_29812,N_29808);
xor UO_1675 (O_1675,N_29959,N_29708);
xor UO_1676 (O_1676,N_29845,N_29658);
or UO_1677 (O_1677,N_29993,N_29419);
and UO_1678 (O_1678,N_29517,N_29424);
or UO_1679 (O_1679,N_29525,N_29895);
xor UO_1680 (O_1680,N_29433,N_29963);
and UO_1681 (O_1681,N_29731,N_29716);
nand UO_1682 (O_1682,N_29798,N_29904);
or UO_1683 (O_1683,N_29762,N_29527);
and UO_1684 (O_1684,N_29922,N_29563);
nor UO_1685 (O_1685,N_29862,N_29440);
and UO_1686 (O_1686,N_29644,N_29907);
nand UO_1687 (O_1687,N_29483,N_29964);
xor UO_1688 (O_1688,N_29738,N_29780);
nand UO_1689 (O_1689,N_29840,N_29775);
nor UO_1690 (O_1690,N_29854,N_29966);
and UO_1691 (O_1691,N_29457,N_29526);
and UO_1692 (O_1692,N_29430,N_29642);
nor UO_1693 (O_1693,N_29717,N_29412);
and UO_1694 (O_1694,N_29508,N_29962);
nor UO_1695 (O_1695,N_29832,N_29942);
or UO_1696 (O_1696,N_29561,N_29908);
and UO_1697 (O_1697,N_29631,N_29501);
or UO_1698 (O_1698,N_29450,N_29911);
or UO_1699 (O_1699,N_29860,N_29782);
and UO_1700 (O_1700,N_29590,N_29767);
xnor UO_1701 (O_1701,N_29502,N_29692);
and UO_1702 (O_1702,N_29958,N_29743);
nor UO_1703 (O_1703,N_29775,N_29459);
xnor UO_1704 (O_1704,N_29744,N_29884);
nor UO_1705 (O_1705,N_29428,N_29747);
and UO_1706 (O_1706,N_29769,N_29929);
and UO_1707 (O_1707,N_29869,N_29528);
or UO_1708 (O_1708,N_29997,N_29993);
or UO_1709 (O_1709,N_29400,N_29842);
nand UO_1710 (O_1710,N_29485,N_29421);
nor UO_1711 (O_1711,N_29805,N_29702);
or UO_1712 (O_1712,N_29792,N_29408);
xnor UO_1713 (O_1713,N_29584,N_29524);
nand UO_1714 (O_1714,N_29722,N_29672);
xor UO_1715 (O_1715,N_29636,N_29588);
or UO_1716 (O_1716,N_29933,N_29694);
nand UO_1717 (O_1717,N_29931,N_29573);
or UO_1718 (O_1718,N_29543,N_29787);
nor UO_1719 (O_1719,N_29725,N_29760);
xor UO_1720 (O_1720,N_29760,N_29572);
or UO_1721 (O_1721,N_29497,N_29767);
nor UO_1722 (O_1722,N_29507,N_29654);
nand UO_1723 (O_1723,N_29870,N_29914);
nand UO_1724 (O_1724,N_29425,N_29813);
nor UO_1725 (O_1725,N_29649,N_29546);
nor UO_1726 (O_1726,N_29880,N_29653);
or UO_1727 (O_1727,N_29631,N_29695);
and UO_1728 (O_1728,N_29482,N_29434);
and UO_1729 (O_1729,N_29810,N_29792);
nor UO_1730 (O_1730,N_29601,N_29699);
nand UO_1731 (O_1731,N_29465,N_29561);
nand UO_1732 (O_1732,N_29962,N_29465);
and UO_1733 (O_1733,N_29739,N_29508);
and UO_1734 (O_1734,N_29837,N_29914);
or UO_1735 (O_1735,N_29418,N_29819);
xnor UO_1736 (O_1736,N_29446,N_29785);
xnor UO_1737 (O_1737,N_29702,N_29649);
and UO_1738 (O_1738,N_29947,N_29567);
and UO_1739 (O_1739,N_29782,N_29471);
xor UO_1740 (O_1740,N_29768,N_29650);
nor UO_1741 (O_1741,N_29763,N_29944);
nand UO_1742 (O_1742,N_29971,N_29777);
and UO_1743 (O_1743,N_29917,N_29925);
or UO_1744 (O_1744,N_29617,N_29748);
xor UO_1745 (O_1745,N_29669,N_29778);
nand UO_1746 (O_1746,N_29424,N_29571);
or UO_1747 (O_1747,N_29504,N_29723);
and UO_1748 (O_1748,N_29944,N_29717);
or UO_1749 (O_1749,N_29598,N_29955);
nand UO_1750 (O_1750,N_29840,N_29858);
xor UO_1751 (O_1751,N_29829,N_29541);
xor UO_1752 (O_1752,N_29869,N_29875);
nand UO_1753 (O_1753,N_29779,N_29822);
nand UO_1754 (O_1754,N_29841,N_29637);
or UO_1755 (O_1755,N_29751,N_29716);
nand UO_1756 (O_1756,N_29436,N_29847);
or UO_1757 (O_1757,N_29879,N_29987);
xor UO_1758 (O_1758,N_29938,N_29838);
nand UO_1759 (O_1759,N_29839,N_29876);
nor UO_1760 (O_1760,N_29824,N_29618);
or UO_1761 (O_1761,N_29479,N_29619);
nand UO_1762 (O_1762,N_29603,N_29709);
nor UO_1763 (O_1763,N_29667,N_29714);
nor UO_1764 (O_1764,N_29427,N_29410);
xnor UO_1765 (O_1765,N_29769,N_29436);
and UO_1766 (O_1766,N_29997,N_29797);
nand UO_1767 (O_1767,N_29680,N_29966);
nor UO_1768 (O_1768,N_29883,N_29680);
xnor UO_1769 (O_1769,N_29728,N_29893);
and UO_1770 (O_1770,N_29596,N_29889);
and UO_1771 (O_1771,N_29709,N_29871);
or UO_1772 (O_1772,N_29916,N_29404);
xor UO_1773 (O_1773,N_29460,N_29435);
and UO_1774 (O_1774,N_29672,N_29655);
and UO_1775 (O_1775,N_29584,N_29606);
or UO_1776 (O_1776,N_29696,N_29868);
or UO_1777 (O_1777,N_29453,N_29953);
and UO_1778 (O_1778,N_29771,N_29695);
xor UO_1779 (O_1779,N_29423,N_29502);
nand UO_1780 (O_1780,N_29435,N_29730);
nor UO_1781 (O_1781,N_29750,N_29720);
and UO_1782 (O_1782,N_29844,N_29610);
or UO_1783 (O_1783,N_29921,N_29860);
xnor UO_1784 (O_1784,N_29870,N_29660);
nand UO_1785 (O_1785,N_29575,N_29574);
or UO_1786 (O_1786,N_29529,N_29540);
nand UO_1787 (O_1787,N_29557,N_29510);
or UO_1788 (O_1788,N_29633,N_29710);
or UO_1789 (O_1789,N_29554,N_29679);
and UO_1790 (O_1790,N_29828,N_29753);
nor UO_1791 (O_1791,N_29629,N_29845);
xnor UO_1792 (O_1792,N_29972,N_29659);
nor UO_1793 (O_1793,N_29545,N_29895);
xnor UO_1794 (O_1794,N_29415,N_29974);
xnor UO_1795 (O_1795,N_29984,N_29661);
nor UO_1796 (O_1796,N_29694,N_29594);
nand UO_1797 (O_1797,N_29938,N_29833);
nor UO_1798 (O_1798,N_29661,N_29547);
and UO_1799 (O_1799,N_29618,N_29521);
nor UO_1800 (O_1800,N_29883,N_29615);
nand UO_1801 (O_1801,N_29458,N_29940);
nor UO_1802 (O_1802,N_29775,N_29781);
or UO_1803 (O_1803,N_29550,N_29969);
nand UO_1804 (O_1804,N_29892,N_29741);
xnor UO_1805 (O_1805,N_29537,N_29778);
nand UO_1806 (O_1806,N_29769,N_29816);
nor UO_1807 (O_1807,N_29716,N_29417);
xor UO_1808 (O_1808,N_29987,N_29933);
or UO_1809 (O_1809,N_29408,N_29552);
and UO_1810 (O_1810,N_29559,N_29472);
nor UO_1811 (O_1811,N_29768,N_29709);
and UO_1812 (O_1812,N_29515,N_29606);
nor UO_1813 (O_1813,N_29767,N_29969);
nand UO_1814 (O_1814,N_29543,N_29821);
or UO_1815 (O_1815,N_29554,N_29986);
nor UO_1816 (O_1816,N_29464,N_29450);
nand UO_1817 (O_1817,N_29669,N_29969);
xor UO_1818 (O_1818,N_29726,N_29406);
nand UO_1819 (O_1819,N_29896,N_29974);
and UO_1820 (O_1820,N_29722,N_29748);
nand UO_1821 (O_1821,N_29536,N_29442);
and UO_1822 (O_1822,N_29771,N_29896);
nand UO_1823 (O_1823,N_29909,N_29636);
xor UO_1824 (O_1824,N_29997,N_29757);
nand UO_1825 (O_1825,N_29935,N_29487);
or UO_1826 (O_1826,N_29743,N_29416);
nand UO_1827 (O_1827,N_29672,N_29923);
or UO_1828 (O_1828,N_29528,N_29454);
or UO_1829 (O_1829,N_29508,N_29652);
nand UO_1830 (O_1830,N_29923,N_29735);
and UO_1831 (O_1831,N_29798,N_29974);
or UO_1832 (O_1832,N_29761,N_29852);
nand UO_1833 (O_1833,N_29451,N_29919);
nand UO_1834 (O_1834,N_29744,N_29835);
and UO_1835 (O_1835,N_29878,N_29589);
or UO_1836 (O_1836,N_29785,N_29875);
or UO_1837 (O_1837,N_29697,N_29974);
or UO_1838 (O_1838,N_29795,N_29670);
nand UO_1839 (O_1839,N_29835,N_29927);
xnor UO_1840 (O_1840,N_29499,N_29815);
and UO_1841 (O_1841,N_29569,N_29778);
xor UO_1842 (O_1842,N_29753,N_29483);
nand UO_1843 (O_1843,N_29899,N_29605);
or UO_1844 (O_1844,N_29594,N_29607);
xor UO_1845 (O_1845,N_29885,N_29692);
nand UO_1846 (O_1846,N_29874,N_29718);
nand UO_1847 (O_1847,N_29801,N_29589);
nand UO_1848 (O_1848,N_29792,N_29806);
xnor UO_1849 (O_1849,N_29536,N_29516);
and UO_1850 (O_1850,N_29538,N_29546);
nor UO_1851 (O_1851,N_29984,N_29974);
nor UO_1852 (O_1852,N_29412,N_29731);
nand UO_1853 (O_1853,N_29819,N_29631);
nor UO_1854 (O_1854,N_29721,N_29928);
or UO_1855 (O_1855,N_29654,N_29853);
xor UO_1856 (O_1856,N_29847,N_29711);
nand UO_1857 (O_1857,N_29578,N_29930);
and UO_1858 (O_1858,N_29428,N_29608);
xnor UO_1859 (O_1859,N_29877,N_29977);
and UO_1860 (O_1860,N_29435,N_29776);
xnor UO_1861 (O_1861,N_29903,N_29651);
and UO_1862 (O_1862,N_29858,N_29570);
or UO_1863 (O_1863,N_29864,N_29879);
and UO_1864 (O_1864,N_29880,N_29809);
or UO_1865 (O_1865,N_29870,N_29922);
xor UO_1866 (O_1866,N_29989,N_29857);
xnor UO_1867 (O_1867,N_29603,N_29620);
nand UO_1868 (O_1868,N_29678,N_29826);
xnor UO_1869 (O_1869,N_29736,N_29669);
xor UO_1870 (O_1870,N_29881,N_29973);
xor UO_1871 (O_1871,N_29599,N_29630);
or UO_1872 (O_1872,N_29626,N_29740);
and UO_1873 (O_1873,N_29743,N_29741);
and UO_1874 (O_1874,N_29675,N_29911);
nor UO_1875 (O_1875,N_29596,N_29600);
or UO_1876 (O_1876,N_29998,N_29597);
nand UO_1877 (O_1877,N_29434,N_29921);
nand UO_1878 (O_1878,N_29818,N_29584);
or UO_1879 (O_1879,N_29820,N_29961);
xnor UO_1880 (O_1880,N_29544,N_29916);
and UO_1881 (O_1881,N_29490,N_29440);
or UO_1882 (O_1882,N_29950,N_29614);
nor UO_1883 (O_1883,N_29702,N_29700);
xor UO_1884 (O_1884,N_29977,N_29454);
and UO_1885 (O_1885,N_29545,N_29701);
xor UO_1886 (O_1886,N_29803,N_29775);
nor UO_1887 (O_1887,N_29872,N_29500);
nand UO_1888 (O_1888,N_29865,N_29873);
nand UO_1889 (O_1889,N_29828,N_29418);
xor UO_1890 (O_1890,N_29802,N_29804);
and UO_1891 (O_1891,N_29850,N_29753);
nand UO_1892 (O_1892,N_29434,N_29499);
or UO_1893 (O_1893,N_29623,N_29730);
nand UO_1894 (O_1894,N_29734,N_29593);
nor UO_1895 (O_1895,N_29534,N_29958);
and UO_1896 (O_1896,N_29877,N_29704);
nand UO_1897 (O_1897,N_29968,N_29886);
nand UO_1898 (O_1898,N_29779,N_29631);
nor UO_1899 (O_1899,N_29998,N_29648);
nand UO_1900 (O_1900,N_29922,N_29670);
nand UO_1901 (O_1901,N_29832,N_29828);
or UO_1902 (O_1902,N_29714,N_29867);
nand UO_1903 (O_1903,N_29790,N_29832);
nor UO_1904 (O_1904,N_29423,N_29427);
nor UO_1905 (O_1905,N_29418,N_29877);
and UO_1906 (O_1906,N_29777,N_29660);
nor UO_1907 (O_1907,N_29673,N_29995);
nor UO_1908 (O_1908,N_29835,N_29475);
or UO_1909 (O_1909,N_29707,N_29678);
nand UO_1910 (O_1910,N_29847,N_29584);
xnor UO_1911 (O_1911,N_29705,N_29856);
nand UO_1912 (O_1912,N_29829,N_29787);
nor UO_1913 (O_1913,N_29928,N_29621);
nor UO_1914 (O_1914,N_29653,N_29794);
or UO_1915 (O_1915,N_29516,N_29869);
xor UO_1916 (O_1916,N_29431,N_29481);
nor UO_1917 (O_1917,N_29587,N_29651);
nand UO_1918 (O_1918,N_29533,N_29654);
or UO_1919 (O_1919,N_29455,N_29959);
or UO_1920 (O_1920,N_29845,N_29948);
nor UO_1921 (O_1921,N_29516,N_29598);
nor UO_1922 (O_1922,N_29931,N_29502);
xor UO_1923 (O_1923,N_29766,N_29906);
or UO_1924 (O_1924,N_29610,N_29543);
and UO_1925 (O_1925,N_29872,N_29714);
nor UO_1926 (O_1926,N_29639,N_29521);
nor UO_1927 (O_1927,N_29665,N_29934);
and UO_1928 (O_1928,N_29821,N_29801);
xor UO_1929 (O_1929,N_29655,N_29682);
nand UO_1930 (O_1930,N_29965,N_29700);
nor UO_1931 (O_1931,N_29895,N_29657);
and UO_1932 (O_1932,N_29699,N_29430);
nand UO_1933 (O_1933,N_29678,N_29697);
and UO_1934 (O_1934,N_29980,N_29894);
or UO_1935 (O_1935,N_29933,N_29409);
nor UO_1936 (O_1936,N_29566,N_29728);
nor UO_1937 (O_1937,N_29833,N_29521);
or UO_1938 (O_1938,N_29643,N_29657);
xor UO_1939 (O_1939,N_29548,N_29702);
nand UO_1940 (O_1940,N_29815,N_29809);
and UO_1941 (O_1941,N_29944,N_29942);
xor UO_1942 (O_1942,N_29628,N_29469);
or UO_1943 (O_1943,N_29947,N_29888);
nand UO_1944 (O_1944,N_29771,N_29593);
xor UO_1945 (O_1945,N_29602,N_29752);
nor UO_1946 (O_1946,N_29526,N_29816);
and UO_1947 (O_1947,N_29567,N_29471);
or UO_1948 (O_1948,N_29678,N_29525);
and UO_1949 (O_1949,N_29977,N_29515);
xor UO_1950 (O_1950,N_29917,N_29962);
nor UO_1951 (O_1951,N_29739,N_29511);
and UO_1952 (O_1952,N_29506,N_29489);
and UO_1953 (O_1953,N_29503,N_29941);
nand UO_1954 (O_1954,N_29840,N_29563);
or UO_1955 (O_1955,N_29786,N_29419);
or UO_1956 (O_1956,N_29930,N_29852);
nor UO_1957 (O_1957,N_29653,N_29846);
xor UO_1958 (O_1958,N_29414,N_29779);
or UO_1959 (O_1959,N_29683,N_29511);
and UO_1960 (O_1960,N_29796,N_29409);
or UO_1961 (O_1961,N_29743,N_29784);
or UO_1962 (O_1962,N_29951,N_29881);
nand UO_1963 (O_1963,N_29932,N_29781);
or UO_1964 (O_1964,N_29892,N_29452);
or UO_1965 (O_1965,N_29658,N_29491);
and UO_1966 (O_1966,N_29741,N_29712);
and UO_1967 (O_1967,N_29534,N_29712);
nor UO_1968 (O_1968,N_29951,N_29929);
or UO_1969 (O_1969,N_29704,N_29812);
xor UO_1970 (O_1970,N_29891,N_29544);
and UO_1971 (O_1971,N_29417,N_29781);
and UO_1972 (O_1972,N_29811,N_29921);
or UO_1973 (O_1973,N_29928,N_29668);
or UO_1974 (O_1974,N_29595,N_29572);
or UO_1975 (O_1975,N_29833,N_29483);
or UO_1976 (O_1976,N_29489,N_29779);
nor UO_1977 (O_1977,N_29965,N_29534);
xor UO_1978 (O_1978,N_29920,N_29700);
xor UO_1979 (O_1979,N_29786,N_29951);
or UO_1980 (O_1980,N_29850,N_29570);
xnor UO_1981 (O_1981,N_29454,N_29998);
xor UO_1982 (O_1982,N_29670,N_29708);
and UO_1983 (O_1983,N_29826,N_29737);
nand UO_1984 (O_1984,N_29964,N_29625);
nand UO_1985 (O_1985,N_29867,N_29686);
or UO_1986 (O_1986,N_29639,N_29886);
xor UO_1987 (O_1987,N_29827,N_29673);
nor UO_1988 (O_1988,N_29489,N_29884);
nand UO_1989 (O_1989,N_29941,N_29865);
xnor UO_1990 (O_1990,N_29661,N_29995);
or UO_1991 (O_1991,N_29816,N_29403);
nand UO_1992 (O_1992,N_29517,N_29840);
or UO_1993 (O_1993,N_29836,N_29590);
and UO_1994 (O_1994,N_29681,N_29417);
or UO_1995 (O_1995,N_29955,N_29500);
nand UO_1996 (O_1996,N_29598,N_29529);
nand UO_1997 (O_1997,N_29818,N_29685);
nor UO_1998 (O_1998,N_29797,N_29827);
or UO_1999 (O_1999,N_29403,N_29730);
nor UO_2000 (O_2000,N_29449,N_29522);
and UO_2001 (O_2001,N_29525,N_29499);
nand UO_2002 (O_2002,N_29663,N_29786);
and UO_2003 (O_2003,N_29458,N_29654);
nor UO_2004 (O_2004,N_29567,N_29826);
and UO_2005 (O_2005,N_29615,N_29795);
and UO_2006 (O_2006,N_29610,N_29719);
nand UO_2007 (O_2007,N_29508,N_29559);
xor UO_2008 (O_2008,N_29799,N_29696);
xor UO_2009 (O_2009,N_29452,N_29751);
nor UO_2010 (O_2010,N_29736,N_29575);
nand UO_2011 (O_2011,N_29780,N_29910);
or UO_2012 (O_2012,N_29866,N_29757);
nand UO_2013 (O_2013,N_29988,N_29595);
xor UO_2014 (O_2014,N_29411,N_29460);
nand UO_2015 (O_2015,N_29818,N_29438);
and UO_2016 (O_2016,N_29944,N_29668);
nor UO_2017 (O_2017,N_29439,N_29459);
and UO_2018 (O_2018,N_29644,N_29614);
nand UO_2019 (O_2019,N_29680,N_29907);
xor UO_2020 (O_2020,N_29852,N_29449);
or UO_2021 (O_2021,N_29563,N_29500);
nor UO_2022 (O_2022,N_29918,N_29583);
xor UO_2023 (O_2023,N_29824,N_29712);
or UO_2024 (O_2024,N_29462,N_29407);
nor UO_2025 (O_2025,N_29506,N_29408);
nand UO_2026 (O_2026,N_29555,N_29970);
nand UO_2027 (O_2027,N_29507,N_29815);
xnor UO_2028 (O_2028,N_29810,N_29549);
xor UO_2029 (O_2029,N_29743,N_29684);
or UO_2030 (O_2030,N_29693,N_29415);
or UO_2031 (O_2031,N_29532,N_29944);
nand UO_2032 (O_2032,N_29458,N_29573);
xor UO_2033 (O_2033,N_29469,N_29679);
nand UO_2034 (O_2034,N_29711,N_29891);
xnor UO_2035 (O_2035,N_29905,N_29695);
nand UO_2036 (O_2036,N_29445,N_29465);
and UO_2037 (O_2037,N_29973,N_29793);
nand UO_2038 (O_2038,N_29976,N_29620);
or UO_2039 (O_2039,N_29994,N_29561);
nand UO_2040 (O_2040,N_29588,N_29571);
or UO_2041 (O_2041,N_29895,N_29878);
nor UO_2042 (O_2042,N_29867,N_29855);
and UO_2043 (O_2043,N_29933,N_29492);
and UO_2044 (O_2044,N_29777,N_29885);
and UO_2045 (O_2045,N_29438,N_29716);
or UO_2046 (O_2046,N_29956,N_29822);
or UO_2047 (O_2047,N_29535,N_29616);
nor UO_2048 (O_2048,N_29565,N_29904);
and UO_2049 (O_2049,N_29481,N_29721);
and UO_2050 (O_2050,N_29445,N_29512);
xor UO_2051 (O_2051,N_29656,N_29908);
xnor UO_2052 (O_2052,N_29430,N_29920);
xnor UO_2053 (O_2053,N_29842,N_29449);
and UO_2054 (O_2054,N_29733,N_29516);
nor UO_2055 (O_2055,N_29922,N_29914);
and UO_2056 (O_2056,N_29635,N_29626);
nor UO_2057 (O_2057,N_29978,N_29462);
and UO_2058 (O_2058,N_29818,N_29937);
nor UO_2059 (O_2059,N_29846,N_29992);
nor UO_2060 (O_2060,N_29537,N_29569);
and UO_2061 (O_2061,N_29537,N_29750);
nor UO_2062 (O_2062,N_29610,N_29583);
or UO_2063 (O_2063,N_29461,N_29973);
nor UO_2064 (O_2064,N_29701,N_29436);
and UO_2065 (O_2065,N_29760,N_29927);
or UO_2066 (O_2066,N_29829,N_29531);
or UO_2067 (O_2067,N_29768,N_29832);
or UO_2068 (O_2068,N_29539,N_29949);
nor UO_2069 (O_2069,N_29789,N_29729);
nor UO_2070 (O_2070,N_29656,N_29907);
xnor UO_2071 (O_2071,N_29977,N_29431);
xor UO_2072 (O_2072,N_29913,N_29452);
and UO_2073 (O_2073,N_29778,N_29525);
or UO_2074 (O_2074,N_29505,N_29851);
nor UO_2075 (O_2075,N_29764,N_29689);
nor UO_2076 (O_2076,N_29875,N_29715);
xor UO_2077 (O_2077,N_29460,N_29731);
or UO_2078 (O_2078,N_29871,N_29836);
and UO_2079 (O_2079,N_29405,N_29416);
and UO_2080 (O_2080,N_29870,N_29669);
or UO_2081 (O_2081,N_29725,N_29558);
nand UO_2082 (O_2082,N_29696,N_29614);
xnor UO_2083 (O_2083,N_29715,N_29610);
or UO_2084 (O_2084,N_29401,N_29650);
xor UO_2085 (O_2085,N_29876,N_29785);
nand UO_2086 (O_2086,N_29533,N_29403);
or UO_2087 (O_2087,N_29765,N_29642);
and UO_2088 (O_2088,N_29741,N_29861);
nor UO_2089 (O_2089,N_29880,N_29609);
or UO_2090 (O_2090,N_29565,N_29664);
nor UO_2091 (O_2091,N_29938,N_29867);
xnor UO_2092 (O_2092,N_29432,N_29649);
xnor UO_2093 (O_2093,N_29452,N_29958);
or UO_2094 (O_2094,N_29735,N_29425);
nor UO_2095 (O_2095,N_29477,N_29750);
nand UO_2096 (O_2096,N_29879,N_29863);
nand UO_2097 (O_2097,N_29919,N_29633);
or UO_2098 (O_2098,N_29527,N_29760);
xor UO_2099 (O_2099,N_29838,N_29939);
nand UO_2100 (O_2100,N_29474,N_29782);
or UO_2101 (O_2101,N_29810,N_29947);
nor UO_2102 (O_2102,N_29665,N_29999);
nand UO_2103 (O_2103,N_29538,N_29744);
nand UO_2104 (O_2104,N_29671,N_29664);
or UO_2105 (O_2105,N_29656,N_29961);
and UO_2106 (O_2106,N_29458,N_29491);
or UO_2107 (O_2107,N_29644,N_29973);
nand UO_2108 (O_2108,N_29504,N_29530);
nand UO_2109 (O_2109,N_29633,N_29567);
xor UO_2110 (O_2110,N_29793,N_29997);
nor UO_2111 (O_2111,N_29748,N_29938);
or UO_2112 (O_2112,N_29438,N_29571);
nor UO_2113 (O_2113,N_29432,N_29613);
or UO_2114 (O_2114,N_29662,N_29516);
or UO_2115 (O_2115,N_29695,N_29578);
nor UO_2116 (O_2116,N_29408,N_29990);
and UO_2117 (O_2117,N_29707,N_29536);
and UO_2118 (O_2118,N_29782,N_29917);
nor UO_2119 (O_2119,N_29608,N_29613);
or UO_2120 (O_2120,N_29543,N_29493);
nor UO_2121 (O_2121,N_29800,N_29871);
xnor UO_2122 (O_2122,N_29824,N_29543);
xnor UO_2123 (O_2123,N_29942,N_29812);
xor UO_2124 (O_2124,N_29808,N_29494);
xnor UO_2125 (O_2125,N_29408,N_29881);
or UO_2126 (O_2126,N_29906,N_29464);
nand UO_2127 (O_2127,N_29553,N_29626);
nor UO_2128 (O_2128,N_29846,N_29943);
and UO_2129 (O_2129,N_29688,N_29857);
xnor UO_2130 (O_2130,N_29801,N_29761);
xnor UO_2131 (O_2131,N_29713,N_29521);
or UO_2132 (O_2132,N_29691,N_29637);
or UO_2133 (O_2133,N_29690,N_29927);
nor UO_2134 (O_2134,N_29772,N_29778);
nand UO_2135 (O_2135,N_29549,N_29794);
nand UO_2136 (O_2136,N_29819,N_29437);
nor UO_2137 (O_2137,N_29844,N_29930);
nor UO_2138 (O_2138,N_29725,N_29444);
and UO_2139 (O_2139,N_29562,N_29429);
or UO_2140 (O_2140,N_29765,N_29906);
or UO_2141 (O_2141,N_29653,N_29433);
xnor UO_2142 (O_2142,N_29891,N_29465);
or UO_2143 (O_2143,N_29586,N_29847);
or UO_2144 (O_2144,N_29931,N_29559);
nand UO_2145 (O_2145,N_29434,N_29732);
or UO_2146 (O_2146,N_29539,N_29735);
nor UO_2147 (O_2147,N_29632,N_29549);
and UO_2148 (O_2148,N_29990,N_29416);
nand UO_2149 (O_2149,N_29511,N_29502);
or UO_2150 (O_2150,N_29942,N_29953);
xor UO_2151 (O_2151,N_29428,N_29986);
and UO_2152 (O_2152,N_29540,N_29469);
xnor UO_2153 (O_2153,N_29416,N_29540);
or UO_2154 (O_2154,N_29989,N_29744);
xnor UO_2155 (O_2155,N_29426,N_29894);
nand UO_2156 (O_2156,N_29806,N_29972);
or UO_2157 (O_2157,N_29455,N_29717);
nand UO_2158 (O_2158,N_29882,N_29674);
xnor UO_2159 (O_2159,N_29534,N_29401);
nand UO_2160 (O_2160,N_29980,N_29442);
xor UO_2161 (O_2161,N_29474,N_29882);
or UO_2162 (O_2162,N_29535,N_29675);
or UO_2163 (O_2163,N_29903,N_29836);
nor UO_2164 (O_2164,N_29712,N_29568);
and UO_2165 (O_2165,N_29989,N_29537);
and UO_2166 (O_2166,N_29452,N_29995);
and UO_2167 (O_2167,N_29480,N_29513);
nor UO_2168 (O_2168,N_29591,N_29461);
or UO_2169 (O_2169,N_29427,N_29675);
nor UO_2170 (O_2170,N_29461,N_29769);
nand UO_2171 (O_2171,N_29813,N_29860);
nor UO_2172 (O_2172,N_29615,N_29987);
and UO_2173 (O_2173,N_29550,N_29403);
and UO_2174 (O_2174,N_29561,N_29918);
or UO_2175 (O_2175,N_29628,N_29614);
and UO_2176 (O_2176,N_29404,N_29748);
xor UO_2177 (O_2177,N_29779,N_29756);
xnor UO_2178 (O_2178,N_29598,N_29498);
and UO_2179 (O_2179,N_29484,N_29823);
and UO_2180 (O_2180,N_29661,N_29702);
or UO_2181 (O_2181,N_29857,N_29414);
or UO_2182 (O_2182,N_29506,N_29886);
and UO_2183 (O_2183,N_29601,N_29978);
nand UO_2184 (O_2184,N_29773,N_29945);
or UO_2185 (O_2185,N_29883,N_29938);
and UO_2186 (O_2186,N_29867,N_29419);
and UO_2187 (O_2187,N_29633,N_29558);
and UO_2188 (O_2188,N_29672,N_29590);
nand UO_2189 (O_2189,N_29701,N_29429);
or UO_2190 (O_2190,N_29478,N_29825);
nor UO_2191 (O_2191,N_29813,N_29912);
or UO_2192 (O_2192,N_29631,N_29673);
nand UO_2193 (O_2193,N_29972,N_29914);
nand UO_2194 (O_2194,N_29423,N_29821);
or UO_2195 (O_2195,N_29794,N_29693);
xor UO_2196 (O_2196,N_29994,N_29517);
nand UO_2197 (O_2197,N_29691,N_29562);
nor UO_2198 (O_2198,N_29476,N_29784);
or UO_2199 (O_2199,N_29613,N_29615);
nand UO_2200 (O_2200,N_29605,N_29795);
and UO_2201 (O_2201,N_29908,N_29659);
nand UO_2202 (O_2202,N_29765,N_29789);
and UO_2203 (O_2203,N_29531,N_29599);
nand UO_2204 (O_2204,N_29653,N_29901);
nand UO_2205 (O_2205,N_29780,N_29888);
nor UO_2206 (O_2206,N_29530,N_29518);
xor UO_2207 (O_2207,N_29746,N_29515);
nand UO_2208 (O_2208,N_29735,N_29949);
and UO_2209 (O_2209,N_29402,N_29809);
or UO_2210 (O_2210,N_29523,N_29492);
xor UO_2211 (O_2211,N_29957,N_29775);
nand UO_2212 (O_2212,N_29999,N_29635);
or UO_2213 (O_2213,N_29646,N_29594);
or UO_2214 (O_2214,N_29640,N_29692);
nor UO_2215 (O_2215,N_29492,N_29674);
or UO_2216 (O_2216,N_29475,N_29751);
nor UO_2217 (O_2217,N_29710,N_29646);
nor UO_2218 (O_2218,N_29647,N_29564);
or UO_2219 (O_2219,N_29781,N_29686);
and UO_2220 (O_2220,N_29838,N_29952);
or UO_2221 (O_2221,N_29631,N_29420);
or UO_2222 (O_2222,N_29658,N_29930);
and UO_2223 (O_2223,N_29533,N_29424);
nand UO_2224 (O_2224,N_29751,N_29554);
nor UO_2225 (O_2225,N_29914,N_29916);
nand UO_2226 (O_2226,N_29854,N_29706);
nand UO_2227 (O_2227,N_29808,N_29871);
or UO_2228 (O_2228,N_29754,N_29757);
nor UO_2229 (O_2229,N_29901,N_29896);
nand UO_2230 (O_2230,N_29911,N_29849);
or UO_2231 (O_2231,N_29895,N_29689);
or UO_2232 (O_2232,N_29427,N_29680);
or UO_2233 (O_2233,N_29629,N_29602);
xor UO_2234 (O_2234,N_29479,N_29880);
nand UO_2235 (O_2235,N_29609,N_29894);
xor UO_2236 (O_2236,N_29551,N_29588);
xnor UO_2237 (O_2237,N_29585,N_29827);
and UO_2238 (O_2238,N_29697,N_29411);
and UO_2239 (O_2239,N_29876,N_29881);
nand UO_2240 (O_2240,N_29712,N_29909);
or UO_2241 (O_2241,N_29780,N_29591);
nor UO_2242 (O_2242,N_29798,N_29919);
nand UO_2243 (O_2243,N_29721,N_29909);
and UO_2244 (O_2244,N_29560,N_29911);
xor UO_2245 (O_2245,N_29785,N_29867);
and UO_2246 (O_2246,N_29800,N_29592);
nand UO_2247 (O_2247,N_29676,N_29628);
and UO_2248 (O_2248,N_29817,N_29824);
nor UO_2249 (O_2249,N_29568,N_29534);
and UO_2250 (O_2250,N_29995,N_29906);
and UO_2251 (O_2251,N_29903,N_29766);
or UO_2252 (O_2252,N_29538,N_29751);
nor UO_2253 (O_2253,N_29614,N_29773);
nor UO_2254 (O_2254,N_29636,N_29400);
nand UO_2255 (O_2255,N_29752,N_29404);
nor UO_2256 (O_2256,N_29785,N_29636);
nor UO_2257 (O_2257,N_29732,N_29675);
xnor UO_2258 (O_2258,N_29817,N_29491);
or UO_2259 (O_2259,N_29937,N_29867);
nand UO_2260 (O_2260,N_29698,N_29410);
xor UO_2261 (O_2261,N_29811,N_29723);
and UO_2262 (O_2262,N_29644,N_29534);
nand UO_2263 (O_2263,N_29895,N_29477);
nor UO_2264 (O_2264,N_29717,N_29866);
or UO_2265 (O_2265,N_29692,N_29567);
nand UO_2266 (O_2266,N_29786,N_29405);
and UO_2267 (O_2267,N_29798,N_29663);
and UO_2268 (O_2268,N_29597,N_29879);
nor UO_2269 (O_2269,N_29570,N_29678);
nand UO_2270 (O_2270,N_29547,N_29944);
xor UO_2271 (O_2271,N_29979,N_29862);
nand UO_2272 (O_2272,N_29697,N_29911);
and UO_2273 (O_2273,N_29668,N_29733);
nand UO_2274 (O_2274,N_29535,N_29412);
nand UO_2275 (O_2275,N_29963,N_29811);
xor UO_2276 (O_2276,N_29463,N_29864);
xor UO_2277 (O_2277,N_29538,N_29641);
nand UO_2278 (O_2278,N_29919,N_29735);
xnor UO_2279 (O_2279,N_29758,N_29418);
xor UO_2280 (O_2280,N_29931,N_29452);
nand UO_2281 (O_2281,N_29538,N_29596);
nand UO_2282 (O_2282,N_29728,N_29994);
and UO_2283 (O_2283,N_29917,N_29937);
and UO_2284 (O_2284,N_29994,N_29931);
or UO_2285 (O_2285,N_29662,N_29540);
nand UO_2286 (O_2286,N_29549,N_29789);
xor UO_2287 (O_2287,N_29891,N_29764);
nand UO_2288 (O_2288,N_29868,N_29857);
nand UO_2289 (O_2289,N_29407,N_29985);
nor UO_2290 (O_2290,N_29489,N_29825);
or UO_2291 (O_2291,N_29426,N_29519);
xnor UO_2292 (O_2292,N_29967,N_29660);
nand UO_2293 (O_2293,N_29692,N_29531);
or UO_2294 (O_2294,N_29721,N_29792);
or UO_2295 (O_2295,N_29982,N_29997);
nand UO_2296 (O_2296,N_29481,N_29602);
nor UO_2297 (O_2297,N_29622,N_29680);
and UO_2298 (O_2298,N_29476,N_29941);
nor UO_2299 (O_2299,N_29438,N_29770);
and UO_2300 (O_2300,N_29759,N_29982);
and UO_2301 (O_2301,N_29646,N_29782);
nand UO_2302 (O_2302,N_29659,N_29899);
nand UO_2303 (O_2303,N_29748,N_29801);
xor UO_2304 (O_2304,N_29946,N_29802);
xor UO_2305 (O_2305,N_29790,N_29869);
nand UO_2306 (O_2306,N_29425,N_29452);
or UO_2307 (O_2307,N_29521,N_29441);
nor UO_2308 (O_2308,N_29900,N_29711);
and UO_2309 (O_2309,N_29796,N_29774);
and UO_2310 (O_2310,N_29436,N_29926);
nor UO_2311 (O_2311,N_29918,N_29673);
nand UO_2312 (O_2312,N_29417,N_29924);
nor UO_2313 (O_2313,N_29540,N_29561);
xor UO_2314 (O_2314,N_29453,N_29922);
nor UO_2315 (O_2315,N_29464,N_29443);
nor UO_2316 (O_2316,N_29668,N_29673);
or UO_2317 (O_2317,N_29745,N_29485);
and UO_2318 (O_2318,N_29782,N_29576);
or UO_2319 (O_2319,N_29927,N_29677);
nand UO_2320 (O_2320,N_29701,N_29460);
nor UO_2321 (O_2321,N_29558,N_29860);
nor UO_2322 (O_2322,N_29907,N_29784);
nand UO_2323 (O_2323,N_29597,N_29808);
xnor UO_2324 (O_2324,N_29840,N_29495);
nor UO_2325 (O_2325,N_29951,N_29497);
nor UO_2326 (O_2326,N_29609,N_29926);
nand UO_2327 (O_2327,N_29584,N_29610);
or UO_2328 (O_2328,N_29919,N_29800);
nor UO_2329 (O_2329,N_29970,N_29503);
or UO_2330 (O_2330,N_29527,N_29846);
nand UO_2331 (O_2331,N_29817,N_29621);
or UO_2332 (O_2332,N_29649,N_29769);
nand UO_2333 (O_2333,N_29527,N_29942);
and UO_2334 (O_2334,N_29666,N_29641);
nor UO_2335 (O_2335,N_29792,N_29976);
nand UO_2336 (O_2336,N_29670,N_29579);
nand UO_2337 (O_2337,N_29939,N_29933);
nand UO_2338 (O_2338,N_29668,N_29865);
nand UO_2339 (O_2339,N_29684,N_29867);
and UO_2340 (O_2340,N_29937,N_29584);
and UO_2341 (O_2341,N_29937,N_29418);
nor UO_2342 (O_2342,N_29913,N_29470);
xnor UO_2343 (O_2343,N_29845,N_29818);
and UO_2344 (O_2344,N_29769,N_29699);
or UO_2345 (O_2345,N_29871,N_29884);
and UO_2346 (O_2346,N_29985,N_29469);
and UO_2347 (O_2347,N_29761,N_29505);
and UO_2348 (O_2348,N_29692,N_29991);
xnor UO_2349 (O_2349,N_29914,N_29453);
nor UO_2350 (O_2350,N_29495,N_29401);
and UO_2351 (O_2351,N_29466,N_29724);
nand UO_2352 (O_2352,N_29646,N_29775);
nand UO_2353 (O_2353,N_29909,N_29955);
nand UO_2354 (O_2354,N_29888,N_29870);
or UO_2355 (O_2355,N_29525,N_29620);
nand UO_2356 (O_2356,N_29687,N_29977);
nand UO_2357 (O_2357,N_29966,N_29847);
or UO_2358 (O_2358,N_29474,N_29446);
or UO_2359 (O_2359,N_29730,N_29453);
or UO_2360 (O_2360,N_29609,N_29595);
and UO_2361 (O_2361,N_29466,N_29736);
or UO_2362 (O_2362,N_29466,N_29731);
and UO_2363 (O_2363,N_29814,N_29669);
or UO_2364 (O_2364,N_29848,N_29664);
and UO_2365 (O_2365,N_29863,N_29629);
nor UO_2366 (O_2366,N_29713,N_29935);
or UO_2367 (O_2367,N_29925,N_29832);
and UO_2368 (O_2368,N_29410,N_29834);
and UO_2369 (O_2369,N_29666,N_29577);
nand UO_2370 (O_2370,N_29681,N_29446);
or UO_2371 (O_2371,N_29815,N_29664);
and UO_2372 (O_2372,N_29599,N_29436);
nor UO_2373 (O_2373,N_29629,N_29791);
or UO_2374 (O_2374,N_29780,N_29896);
xnor UO_2375 (O_2375,N_29520,N_29439);
xnor UO_2376 (O_2376,N_29905,N_29948);
and UO_2377 (O_2377,N_29877,N_29882);
and UO_2378 (O_2378,N_29915,N_29857);
and UO_2379 (O_2379,N_29613,N_29551);
and UO_2380 (O_2380,N_29676,N_29672);
and UO_2381 (O_2381,N_29478,N_29400);
or UO_2382 (O_2382,N_29522,N_29462);
xor UO_2383 (O_2383,N_29818,N_29413);
nand UO_2384 (O_2384,N_29709,N_29795);
xnor UO_2385 (O_2385,N_29559,N_29906);
xnor UO_2386 (O_2386,N_29993,N_29690);
nor UO_2387 (O_2387,N_29993,N_29755);
xnor UO_2388 (O_2388,N_29813,N_29959);
nor UO_2389 (O_2389,N_29996,N_29805);
and UO_2390 (O_2390,N_29699,N_29961);
and UO_2391 (O_2391,N_29502,N_29425);
or UO_2392 (O_2392,N_29760,N_29434);
nand UO_2393 (O_2393,N_29468,N_29780);
xnor UO_2394 (O_2394,N_29592,N_29759);
nand UO_2395 (O_2395,N_29818,N_29831);
or UO_2396 (O_2396,N_29411,N_29571);
and UO_2397 (O_2397,N_29441,N_29664);
nor UO_2398 (O_2398,N_29797,N_29857);
nor UO_2399 (O_2399,N_29726,N_29849);
nor UO_2400 (O_2400,N_29846,N_29499);
and UO_2401 (O_2401,N_29477,N_29534);
nand UO_2402 (O_2402,N_29692,N_29833);
nand UO_2403 (O_2403,N_29702,N_29922);
xnor UO_2404 (O_2404,N_29742,N_29695);
or UO_2405 (O_2405,N_29610,N_29598);
nand UO_2406 (O_2406,N_29727,N_29569);
nand UO_2407 (O_2407,N_29938,N_29474);
xnor UO_2408 (O_2408,N_29481,N_29878);
and UO_2409 (O_2409,N_29838,N_29427);
xnor UO_2410 (O_2410,N_29726,N_29470);
nand UO_2411 (O_2411,N_29608,N_29768);
nand UO_2412 (O_2412,N_29571,N_29885);
and UO_2413 (O_2413,N_29558,N_29717);
and UO_2414 (O_2414,N_29889,N_29526);
and UO_2415 (O_2415,N_29790,N_29451);
nand UO_2416 (O_2416,N_29894,N_29984);
xnor UO_2417 (O_2417,N_29718,N_29546);
xor UO_2418 (O_2418,N_29754,N_29842);
xor UO_2419 (O_2419,N_29443,N_29591);
and UO_2420 (O_2420,N_29621,N_29541);
xnor UO_2421 (O_2421,N_29629,N_29798);
or UO_2422 (O_2422,N_29868,N_29972);
nor UO_2423 (O_2423,N_29410,N_29917);
xnor UO_2424 (O_2424,N_29500,N_29743);
xnor UO_2425 (O_2425,N_29831,N_29779);
or UO_2426 (O_2426,N_29871,N_29977);
xnor UO_2427 (O_2427,N_29631,N_29725);
and UO_2428 (O_2428,N_29912,N_29592);
and UO_2429 (O_2429,N_29835,N_29574);
nand UO_2430 (O_2430,N_29958,N_29519);
nor UO_2431 (O_2431,N_29730,N_29529);
nand UO_2432 (O_2432,N_29941,N_29976);
nor UO_2433 (O_2433,N_29861,N_29661);
and UO_2434 (O_2434,N_29920,N_29779);
or UO_2435 (O_2435,N_29646,N_29447);
or UO_2436 (O_2436,N_29676,N_29955);
nand UO_2437 (O_2437,N_29771,N_29832);
nand UO_2438 (O_2438,N_29887,N_29706);
nor UO_2439 (O_2439,N_29579,N_29915);
and UO_2440 (O_2440,N_29922,N_29960);
nor UO_2441 (O_2441,N_29552,N_29562);
xnor UO_2442 (O_2442,N_29419,N_29641);
nor UO_2443 (O_2443,N_29419,N_29861);
or UO_2444 (O_2444,N_29681,N_29599);
or UO_2445 (O_2445,N_29915,N_29597);
nand UO_2446 (O_2446,N_29913,N_29400);
or UO_2447 (O_2447,N_29600,N_29581);
nor UO_2448 (O_2448,N_29459,N_29462);
nand UO_2449 (O_2449,N_29615,N_29955);
nand UO_2450 (O_2450,N_29682,N_29617);
and UO_2451 (O_2451,N_29995,N_29584);
xor UO_2452 (O_2452,N_29625,N_29530);
xor UO_2453 (O_2453,N_29954,N_29560);
and UO_2454 (O_2454,N_29496,N_29690);
xnor UO_2455 (O_2455,N_29886,N_29806);
or UO_2456 (O_2456,N_29520,N_29650);
xnor UO_2457 (O_2457,N_29504,N_29455);
nand UO_2458 (O_2458,N_29997,N_29441);
or UO_2459 (O_2459,N_29557,N_29650);
xnor UO_2460 (O_2460,N_29465,N_29581);
and UO_2461 (O_2461,N_29969,N_29595);
xor UO_2462 (O_2462,N_29706,N_29402);
and UO_2463 (O_2463,N_29600,N_29772);
nor UO_2464 (O_2464,N_29884,N_29423);
and UO_2465 (O_2465,N_29474,N_29497);
and UO_2466 (O_2466,N_29476,N_29439);
or UO_2467 (O_2467,N_29879,N_29767);
xor UO_2468 (O_2468,N_29749,N_29627);
xor UO_2469 (O_2469,N_29565,N_29614);
nor UO_2470 (O_2470,N_29912,N_29792);
or UO_2471 (O_2471,N_29491,N_29438);
nand UO_2472 (O_2472,N_29511,N_29877);
xnor UO_2473 (O_2473,N_29903,N_29866);
nor UO_2474 (O_2474,N_29944,N_29834);
and UO_2475 (O_2475,N_29460,N_29482);
or UO_2476 (O_2476,N_29692,N_29883);
nor UO_2477 (O_2477,N_29879,N_29526);
nor UO_2478 (O_2478,N_29554,N_29608);
xnor UO_2479 (O_2479,N_29772,N_29685);
or UO_2480 (O_2480,N_29770,N_29877);
nor UO_2481 (O_2481,N_29443,N_29609);
nor UO_2482 (O_2482,N_29974,N_29529);
or UO_2483 (O_2483,N_29726,N_29784);
and UO_2484 (O_2484,N_29505,N_29636);
or UO_2485 (O_2485,N_29404,N_29879);
nand UO_2486 (O_2486,N_29904,N_29583);
xor UO_2487 (O_2487,N_29790,N_29641);
or UO_2488 (O_2488,N_29645,N_29864);
nor UO_2489 (O_2489,N_29591,N_29932);
or UO_2490 (O_2490,N_29564,N_29536);
nor UO_2491 (O_2491,N_29671,N_29790);
and UO_2492 (O_2492,N_29502,N_29754);
nor UO_2493 (O_2493,N_29517,N_29558);
xnor UO_2494 (O_2494,N_29515,N_29461);
and UO_2495 (O_2495,N_29629,N_29411);
xnor UO_2496 (O_2496,N_29625,N_29720);
nand UO_2497 (O_2497,N_29695,N_29609);
nand UO_2498 (O_2498,N_29495,N_29470);
nand UO_2499 (O_2499,N_29650,N_29486);
nor UO_2500 (O_2500,N_29861,N_29407);
nor UO_2501 (O_2501,N_29781,N_29888);
and UO_2502 (O_2502,N_29854,N_29600);
or UO_2503 (O_2503,N_29671,N_29729);
nor UO_2504 (O_2504,N_29485,N_29894);
nand UO_2505 (O_2505,N_29621,N_29745);
nor UO_2506 (O_2506,N_29548,N_29789);
nor UO_2507 (O_2507,N_29473,N_29446);
xor UO_2508 (O_2508,N_29606,N_29726);
nand UO_2509 (O_2509,N_29794,N_29479);
nand UO_2510 (O_2510,N_29727,N_29622);
or UO_2511 (O_2511,N_29922,N_29884);
nor UO_2512 (O_2512,N_29786,N_29799);
or UO_2513 (O_2513,N_29745,N_29425);
or UO_2514 (O_2514,N_29586,N_29497);
nor UO_2515 (O_2515,N_29711,N_29750);
xor UO_2516 (O_2516,N_29760,N_29897);
nor UO_2517 (O_2517,N_29579,N_29838);
or UO_2518 (O_2518,N_29711,N_29626);
and UO_2519 (O_2519,N_29761,N_29653);
and UO_2520 (O_2520,N_29462,N_29742);
nor UO_2521 (O_2521,N_29673,N_29812);
or UO_2522 (O_2522,N_29644,N_29956);
xor UO_2523 (O_2523,N_29699,N_29705);
and UO_2524 (O_2524,N_29815,N_29470);
nand UO_2525 (O_2525,N_29821,N_29724);
nand UO_2526 (O_2526,N_29577,N_29563);
xnor UO_2527 (O_2527,N_29658,N_29919);
or UO_2528 (O_2528,N_29771,N_29680);
and UO_2529 (O_2529,N_29568,N_29707);
nor UO_2530 (O_2530,N_29941,N_29950);
nand UO_2531 (O_2531,N_29939,N_29822);
nand UO_2532 (O_2532,N_29513,N_29893);
and UO_2533 (O_2533,N_29458,N_29757);
and UO_2534 (O_2534,N_29645,N_29861);
or UO_2535 (O_2535,N_29849,N_29809);
nand UO_2536 (O_2536,N_29504,N_29747);
nor UO_2537 (O_2537,N_29952,N_29470);
nand UO_2538 (O_2538,N_29489,N_29446);
nor UO_2539 (O_2539,N_29726,N_29509);
or UO_2540 (O_2540,N_29909,N_29482);
nand UO_2541 (O_2541,N_29906,N_29552);
nor UO_2542 (O_2542,N_29824,N_29656);
and UO_2543 (O_2543,N_29876,N_29736);
nor UO_2544 (O_2544,N_29932,N_29490);
or UO_2545 (O_2545,N_29999,N_29639);
or UO_2546 (O_2546,N_29614,N_29568);
or UO_2547 (O_2547,N_29940,N_29566);
xnor UO_2548 (O_2548,N_29807,N_29465);
xor UO_2549 (O_2549,N_29591,N_29631);
and UO_2550 (O_2550,N_29417,N_29943);
or UO_2551 (O_2551,N_29555,N_29577);
nand UO_2552 (O_2552,N_29698,N_29859);
xor UO_2553 (O_2553,N_29907,N_29943);
and UO_2554 (O_2554,N_29723,N_29538);
and UO_2555 (O_2555,N_29796,N_29977);
or UO_2556 (O_2556,N_29806,N_29975);
nor UO_2557 (O_2557,N_29951,N_29785);
and UO_2558 (O_2558,N_29990,N_29991);
and UO_2559 (O_2559,N_29886,N_29655);
or UO_2560 (O_2560,N_29655,N_29625);
nand UO_2561 (O_2561,N_29419,N_29809);
or UO_2562 (O_2562,N_29430,N_29458);
nand UO_2563 (O_2563,N_29654,N_29467);
xor UO_2564 (O_2564,N_29477,N_29436);
xor UO_2565 (O_2565,N_29467,N_29755);
nand UO_2566 (O_2566,N_29662,N_29676);
or UO_2567 (O_2567,N_29481,N_29413);
and UO_2568 (O_2568,N_29605,N_29971);
or UO_2569 (O_2569,N_29405,N_29626);
xor UO_2570 (O_2570,N_29787,N_29863);
nand UO_2571 (O_2571,N_29756,N_29864);
and UO_2572 (O_2572,N_29494,N_29558);
xor UO_2573 (O_2573,N_29942,N_29512);
and UO_2574 (O_2574,N_29452,N_29691);
or UO_2575 (O_2575,N_29867,N_29718);
nor UO_2576 (O_2576,N_29926,N_29655);
nor UO_2577 (O_2577,N_29937,N_29713);
xor UO_2578 (O_2578,N_29839,N_29402);
or UO_2579 (O_2579,N_29718,N_29884);
nand UO_2580 (O_2580,N_29928,N_29874);
or UO_2581 (O_2581,N_29683,N_29446);
xor UO_2582 (O_2582,N_29683,N_29607);
nand UO_2583 (O_2583,N_29852,N_29830);
nand UO_2584 (O_2584,N_29407,N_29579);
xnor UO_2585 (O_2585,N_29986,N_29894);
xnor UO_2586 (O_2586,N_29610,N_29862);
nand UO_2587 (O_2587,N_29833,N_29491);
xor UO_2588 (O_2588,N_29915,N_29663);
nor UO_2589 (O_2589,N_29863,N_29731);
xnor UO_2590 (O_2590,N_29971,N_29986);
and UO_2591 (O_2591,N_29809,N_29803);
nor UO_2592 (O_2592,N_29738,N_29505);
and UO_2593 (O_2593,N_29709,N_29655);
nor UO_2594 (O_2594,N_29915,N_29428);
and UO_2595 (O_2595,N_29948,N_29775);
nand UO_2596 (O_2596,N_29884,N_29702);
and UO_2597 (O_2597,N_29457,N_29451);
and UO_2598 (O_2598,N_29931,N_29441);
or UO_2599 (O_2599,N_29877,N_29445);
nor UO_2600 (O_2600,N_29997,N_29616);
nand UO_2601 (O_2601,N_29441,N_29631);
nand UO_2602 (O_2602,N_29623,N_29781);
and UO_2603 (O_2603,N_29712,N_29983);
xnor UO_2604 (O_2604,N_29567,N_29860);
xnor UO_2605 (O_2605,N_29755,N_29938);
or UO_2606 (O_2606,N_29845,N_29882);
or UO_2607 (O_2607,N_29682,N_29600);
nor UO_2608 (O_2608,N_29780,N_29497);
or UO_2609 (O_2609,N_29611,N_29477);
nand UO_2610 (O_2610,N_29944,N_29428);
nand UO_2611 (O_2611,N_29815,N_29573);
or UO_2612 (O_2612,N_29418,N_29527);
nor UO_2613 (O_2613,N_29925,N_29438);
nand UO_2614 (O_2614,N_29728,N_29989);
xor UO_2615 (O_2615,N_29551,N_29578);
and UO_2616 (O_2616,N_29918,N_29455);
or UO_2617 (O_2617,N_29817,N_29444);
nor UO_2618 (O_2618,N_29564,N_29879);
and UO_2619 (O_2619,N_29890,N_29455);
xnor UO_2620 (O_2620,N_29428,N_29972);
nor UO_2621 (O_2621,N_29646,N_29811);
nand UO_2622 (O_2622,N_29887,N_29400);
xnor UO_2623 (O_2623,N_29585,N_29545);
nand UO_2624 (O_2624,N_29712,N_29976);
and UO_2625 (O_2625,N_29632,N_29446);
nor UO_2626 (O_2626,N_29475,N_29464);
or UO_2627 (O_2627,N_29406,N_29872);
and UO_2628 (O_2628,N_29991,N_29856);
or UO_2629 (O_2629,N_29801,N_29588);
xnor UO_2630 (O_2630,N_29569,N_29737);
and UO_2631 (O_2631,N_29546,N_29867);
xor UO_2632 (O_2632,N_29451,N_29920);
or UO_2633 (O_2633,N_29778,N_29482);
nand UO_2634 (O_2634,N_29479,N_29819);
and UO_2635 (O_2635,N_29856,N_29619);
or UO_2636 (O_2636,N_29447,N_29469);
nor UO_2637 (O_2637,N_29800,N_29689);
nor UO_2638 (O_2638,N_29874,N_29910);
or UO_2639 (O_2639,N_29904,N_29618);
nand UO_2640 (O_2640,N_29422,N_29473);
nand UO_2641 (O_2641,N_29852,N_29818);
nor UO_2642 (O_2642,N_29521,N_29554);
xnor UO_2643 (O_2643,N_29627,N_29654);
and UO_2644 (O_2644,N_29489,N_29412);
or UO_2645 (O_2645,N_29790,N_29520);
xnor UO_2646 (O_2646,N_29486,N_29779);
xnor UO_2647 (O_2647,N_29985,N_29571);
and UO_2648 (O_2648,N_29759,N_29535);
nand UO_2649 (O_2649,N_29595,N_29628);
nor UO_2650 (O_2650,N_29771,N_29528);
nor UO_2651 (O_2651,N_29723,N_29556);
nand UO_2652 (O_2652,N_29733,N_29918);
nand UO_2653 (O_2653,N_29868,N_29584);
and UO_2654 (O_2654,N_29640,N_29480);
xor UO_2655 (O_2655,N_29792,N_29655);
xor UO_2656 (O_2656,N_29826,N_29497);
or UO_2657 (O_2657,N_29668,N_29473);
xnor UO_2658 (O_2658,N_29678,N_29504);
nor UO_2659 (O_2659,N_29678,N_29945);
and UO_2660 (O_2660,N_29485,N_29949);
xor UO_2661 (O_2661,N_29541,N_29615);
and UO_2662 (O_2662,N_29759,N_29481);
and UO_2663 (O_2663,N_29943,N_29912);
nand UO_2664 (O_2664,N_29914,N_29770);
xnor UO_2665 (O_2665,N_29544,N_29819);
or UO_2666 (O_2666,N_29863,N_29872);
xnor UO_2667 (O_2667,N_29746,N_29546);
and UO_2668 (O_2668,N_29639,N_29755);
or UO_2669 (O_2669,N_29669,N_29864);
or UO_2670 (O_2670,N_29655,N_29783);
nand UO_2671 (O_2671,N_29627,N_29956);
xor UO_2672 (O_2672,N_29448,N_29832);
and UO_2673 (O_2673,N_29684,N_29472);
nor UO_2674 (O_2674,N_29550,N_29901);
nand UO_2675 (O_2675,N_29935,N_29810);
nand UO_2676 (O_2676,N_29825,N_29679);
nand UO_2677 (O_2677,N_29993,N_29995);
nand UO_2678 (O_2678,N_29532,N_29794);
and UO_2679 (O_2679,N_29839,N_29752);
nand UO_2680 (O_2680,N_29522,N_29410);
xor UO_2681 (O_2681,N_29918,N_29756);
nor UO_2682 (O_2682,N_29990,N_29633);
nor UO_2683 (O_2683,N_29671,N_29953);
nor UO_2684 (O_2684,N_29912,N_29606);
and UO_2685 (O_2685,N_29561,N_29757);
or UO_2686 (O_2686,N_29712,N_29813);
nor UO_2687 (O_2687,N_29997,N_29598);
xor UO_2688 (O_2688,N_29803,N_29998);
or UO_2689 (O_2689,N_29723,N_29685);
xor UO_2690 (O_2690,N_29607,N_29415);
xnor UO_2691 (O_2691,N_29476,N_29951);
nand UO_2692 (O_2692,N_29997,N_29967);
and UO_2693 (O_2693,N_29526,N_29582);
nand UO_2694 (O_2694,N_29518,N_29761);
or UO_2695 (O_2695,N_29856,N_29869);
or UO_2696 (O_2696,N_29508,N_29497);
nor UO_2697 (O_2697,N_29414,N_29534);
xnor UO_2698 (O_2698,N_29594,N_29602);
xor UO_2699 (O_2699,N_29501,N_29426);
and UO_2700 (O_2700,N_29742,N_29452);
nor UO_2701 (O_2701,N_29688,N_29684);
xnor UO_2702 (O_2702,N_29702,N_29741);
and UO_2703 (O_2703,N_29721,N_29693);
nand UO_2704 (O_2704,N_29518,N_29945);
nand UO_2705 (O_2705,N_29708,N_29934);
nor UO_2706 (O_2706,N_29987,N_29853);
nand UO_2707 (O_2707,N_29934,N_29491);
nand UO_2708 (O_2708,N_29402,N_29972);
nand UO_2709 (O_2709,N_29941,N_29484);
and UO_2710 (O_2710,N_29547,N_29643);
or UO_2711 (O_2711,N_29465,N_29617);
or UO_2712 (O_2712,N_29948,N_29726);
and UO_2713 (O_2713,N_29426,N_29943);
and UO_2714 (O_2714,N_29509,N_29662);
nor UO_2715 (O_2715,N_29770,N_29966);
or UO_2716 (O_2716,N_29444,N_29942);
nand UO_2717 (O_2717,N_29503,N_29423);
xnor UO_2718 (O_2718,N_29751,N_29530);
nand UO_2719 (O_2719,N_29461,N_29838);
nor UO_2720 (O_2720,N_29841,N_29853);
nor UO_2721 (O_2721,N_29835,N_29801);
and UO_2722 (O_2722,N_29681,N_29936);
or UO_2723 (O_2723,N_29621,N_29499);
nor UO_2724 (O_2724,N_29888,N_29449);
nand UO_2725 (O_2725,N_29772,N_29797);
nand UO_2726 (O_2726,N_29991,N_29753);
xor UO_2727 (O_2727,N_29433,N_29496);
nand UO_2728 (O_2728,N_29887,N_29777);
xor UO_2729 (O_2729,N_29631,N_29432);
xor UO_2730 (O_2730,N_29900,N_29738);
xor UO_2731 (O_2731,N_29680,N_29990);
and UO_2732 (O_2732,N_29805,N_29491);
nor UO_2733 (O_2733,N_29929,N_29473);
or UO_2734 (O_2734,N_29988,N_29969);
nor UO_2735 (O_2735,N_29583,N_29766);
nand UO_2736 (O_2736,N_29645,N_29603);
nor UO_2737 (O_2737,N_29910,N_29748);
nor UO_2738 (O_2738,N_29886,N_29769);
nor UO_2739 (O_2739,N_29687,N_29826);
nand UO_2740 (O_2740,N_29820,N_29768);
and UO_2741 (O_2741,N_29890,N_29544);
nor UO_2742 (O_2742,N_29884,N_29422);
nor UO_2743 (O_2743,N_29414,N_29778);
or UO_2744 (O_2744,N_29735,N_29414);
xor UO_2745 (O_2745,N_29535,N_29600);
or UO_2746 (O_2746,N_29718,N_29542);
xor UO_2747 (O_2747,N_29668,N_29431);
xnor UO_2748 (O_2748,N_29638,N_29460);
nor UO_2749 (O_2749,N_29742,N_29941);
and UO_2750 (O_2750,N_29556,N_29586);
or UO_2751 (O_2751,N_29666,N_29890);
xnor UO_2752 (O_2752,N_29829,N_29818);
and UO_2753 (O_2753,N_29708,N_29725);
xor UO_2754 (O_2754,N_29993,N_29737);
nand UO_2755 (O_2755,N_29946,N_29743);
nand UO_2756 (O_2756,N_29894,N_29711);
and UO_2757 (O_2757,N_29888,N_29550);
nand UO_2758 (O_2758,N_29800,N_29802);
xnor UO_2759 (O_2759,N_29941,N_29438);
nor UO_2760 (O_2760,N_29892,N_29631);
or UO_2761 (O_2761,N_29472,N_29947);
or UO_2762 (O_2762,N_29585,N_29875);
xor UO_2763 (O_2763,N_29542,N_29668);
and UO_2764 (O_2764,N_29885,N_29587);
xor UO_2765 (O_2765,N_29695,N_29795);
nor UO_2766 (O_2766,N_29749,N_29840);
nor UO_2767 (O_2767,N_29566,N_29964);
nor UO_2768 (O_2768,N_29609,N_29560);
or UO_2769 (O_2769,N_29856,N_29559);
nand UO_2770 (O_2770,N_29691,N_29628);
and UO_2771 (O_2771,N_29985,N_29419);
xnor UO_2772 (O_2772,N_29990,N_29554);
nor UO_2773 (O_2773,N_29587,N_29488);
or UO_2774 (O_2774,N_29839,N_29805);
and UO_2775 (O_2775,N_29762,N_29549);
nand UO_2776 (O_2776,N_29920,N_29638);
and UO_2777 (O_2777,N_29989,N_29605);
and UO_2778 (O_2778,N_29531,N_29600);
nor UO_2779 (O_2779,N_29644,N_29998);
nand UO_2780 (O_2780,N_29413,N_29470);
nor UO_2781 (O_2781,N_29716,N_29690);
xnor UO_2782 (O_2782,N_29701,N_29613);
or UO_2783 (O_2783,N_29837,N_29473);
xor UO_2784 (O_2784,N_29591,N_29453);
or UO_2785 (O_2785,N_29736,N_29747);
nand UO_2786 (O_2786,N_29624,N_29745);
nand UO_2787 (O_2787,N_29793,N_29942);
and UO_2788 (O_2788,N_29722,N_29834);
nor UO_2789 (O_2789,N_29743,N_29646);
nor UO_2790 (O_2790,N_29786,N_29579);
nor UO_2791 (O_2791,N_29707,N_29558);
nand UO_2792 (O_2792,N_29614,N_29478);
xor UO_2793 (O_2793,N_29410,N_29437);
xor UO_2794 (O_2794,N_29527,N_29511);
nor UO_2795 (O_2795,N_29736,N_29844);
or UO_2796 (O_2796,N_29989,N_29906);
or UO_2797 (O_2797,N_29539,N_29656);
and UO_2798 (O_2798,N_29651,N_29593);
nand UO_2799 (O_2799,N_29614,N_29558);
or UO_2800 (O_2800,N_29477,N_29600);
xor UO_2801 (O_2801,N_29837,N_29503);
nor UO_2802 (O_2802,N_29636,N_29639);
or UO_2803 (O_2803,N_29897,N_29987);
and UO_2804 (O_2804,N_29527,N_29874);
xor UO_2805 (O_2805,N_29993,N_29531);
or UO_2806 (O_2806,N_29411,N_29528);
or UO_2807 (O_2807,N_29989,N_29431);
or UO_2808 (O_2808,N_29632,N_29860);
nand UO_2809 (O_2809,N_29953,N_29927);
or UO_2810 (O_2810,N_29783,N_29828);
nand UO_2811 (O_2811,N_29479,N_29643);
nand UO_2812 (O_2812,N_29766,N_29720);
nand UO_2813 (O_2813,N_29988,N_29672);
or UO_2814 (O_2814,N_29605,N_29792);
xnor UO_2815 (O_2815,N_29787,N_29480);
or UO_2816 (O_2816,N_29516,N_29555);
nor UO_2817 (O_2817,N_29839,N_29840);
nand UO_2818 (O_2818,N_29635,N_29843);
nor UO_2819 (O_2819,N_29474,N_29728);
and UO_2820 (O_2820,N_29751,N_29528);
xnor UO_2821 (O_2821,N_29849,N_29798);
or UO_2822 (O_2822,N_29845,N_29847);
or UO_2823 (O_2823,N_29484,N_29555);
nor UO_2824 (O_2824,N_29632,N_29981);
nor UO_2825 (O_2825,N_29796,N_29957);
nand UO_2826 (O_2826,N_29608,N_29806);
nor UO_2827 (O_2827,N_29899,N_29440);
xnor UO_2828 (O_2828,N_29574,N_29605);
nor UO_2829 (O_2829,N_29885,N_29689);
xor UO_2830 (O_2830,N_29818,N_29611);
or UO_2831 (O_2831,N_29965,N_29894);
nor UO_2832 (O_2832,N_29487,N_29458);
and UO_2833 (O_2833,N_29889,N_29445);
and UO_2834 (O_2834,N_29935,N_29456);
xor UO_2835 (O_2835,N_29754,N_29549);
or UO_2836 (O_2836,N_29511,N_29742);
nor UO_2837 (O_2837,N_29588,N_29773);
or UO_2838 (O_2838,N_29502,N_29774);
nand UO_2839 (O_2839,N_29826,N_29640);
nand UO_2840 (O_2840,N_29516,N_29415);
nand UO_2841 (O_2841,N_29905,N_29884);
and UO_2842 (O_2842,N_29609,N_29589);
or UO_2843 (O_2843,N_29988,N_29981);
nand UO_2844 (O_2844,N_29427,N_29757);
and UO_2845 (O_2845,N_29834,N_29466);
and UO_2846 (O_2846,N_29407,N_29543);
nand UO_2847 (O_2847,N_29992,N_29919);
xnor UO_2848 (O_2848,N_29890,N_29649);
nor UO_2849 (O_2849,N_29919,N_29694);
nor UO_2850 (O_2850,N_29683,N_29695);
nor UO_2851 (O_2851,N_29843,N_29461);
xor UO_2852 (O_2852,N_29633,N_29564);
and UO_2853 (O_2853,N_29577,N_29794);
and UO_2854 (O_2854,N_29757,N_29538);
nor UO_2855 (O_2855,N_29794,N_29578);
xor UO_2856 (O_2856,N_29803,N_29762);
nand UO_2857 (O_2857,N_29407,N_29886);
xnor UO_2858 (O_2858,N_29420,N_29672);
or UO_2859 (O_2859,N_29995,N_29652);
nor UO_2860 (O_2860,N_29629,N_29813);
and UO_2861 (O_2861,N_29453,N_29479);
or UO_2862 (O_2862,N_29982,N_29916);
xnor UO_2863 (O_2863,N_29416,N_29504);
and UO_2864 (O_2864,N_29489,N_29487);
nor UO_2865 (O_2865,N_29946,N_29478);
or UO_2866 (O_2866,N_29663,N_29830);
nor UO_2867 (O_2867,N_29433,N_29840);
or UO_2868 (O_2868,N_29511,N_29541);
and UO_2869 (O_2869,N_29817,N_29898);
nor UO_2870 (O_2870,N_29930,N_29804);
or UO_2871 (O_2871,N_29631,N_29449);
or UO_2872 (O_2872,N_29435,N_29654);
xor UO_2873 (O_2873,N_29742,N_29962);
nand UO_2874 (O_2874,N_29581,N_29702);
nor UO_2875 (O_2875,N_29705,N_29632);
and UO_2876 (O_2876,N_29775,N_29414);
nand UO_2877 (O_2877,N_29659,N_29654);
xor UO_2878 (O_2878,N_29402,N_29731);
nand UO_2879 (O_2879,N_29706,N_29418);
nand UO_2880 (O_2880,N_29984,N_29803);
or UO_2881 (O_2881,N_29602,N_29718);
and UO_2882 (O_2882,N_29529,N_29620);
or UO_2883 (O_2883,N_29881,N_29453);
nor UO_2884 (O_2884,N_29739,N_29683);
or UO_2885 (O_2885,N_29709,N_29841);
xnor UO_2886 (O_2886,N_29640,N_29519);
nand UO_2887 (O_2887,N_29496,N_29613);
nand UO_2888 (O_2888,N_29652,N_29940);
nand UO_2889 (O_2889,N_29524,N_29438);
nand UO_2890 (O_2890,N_29761,N_29926);
nor UO_2891 (O_2891,N_29705,N_29753);
and UO_2892 (O_2892,N_29740,N_29431);
nor UO_2893 (O_2893,N_29612,N_29716);
nand UO_2894 (O_2894,N_29914,N_29760);
or UO_2895 (O_2895,N_29431,N_29656);
nor UO_2896 (O_2896,N_29771,N_29793);
or UO_2897 (O_2897,N_29404,N_29880);
nor UO_2898 (O_2898,N_29558,N_29990);
nor UO_2899 (O_2899,N_29680,N_29426);
or UO_2900 (O_2900,N_29928,N_29649);
nor UO_2901 (O_2901,N_29698,N_29987);
or UO_2902 (O_2902,N_29616,N_29771);
or UO_2903 (O_2903,N_29412,N_29912);
nand UO_2904 (O_2904,N_29502,N_29640);
nand UO_2905 (O_2905,N_29653,N_29811);
xnor UO_2906 (O_2906,N_29630,N_29482);
nor UO_2907 (O_2907,N_29457,N_29916);
and UO_2908 (O_2908,N_29991,N_29868);
nand UO_2909 (O_2909,N_29815,N_29498);
xnor UO_2910 (O_2910,N_29568,N_29697);
xnor UO_2911 (O_2911,N_29431,N_29976);
xnor UO_2912 (O_2912,N_29459,N_29769);
and UO_2913 (O_2913,N_29417,N_29516);
and UO_2914 (O_2914,N_29518,N_29635);
nand UO_2915 (O_2915,N_29558,N_29923);
xor UO_2916 (O_2916,N_29766,N_29941);
xor UO_2917 (O_2917,N_29925,N_29789);
and UO_2918 (O_2918,N_29987,N_29466);
nor UO_2919 (O_2919,N_29760,N_29558);
or UO_2920 (O_2920,N_29909,N_29862);
or UO_2921 (O_2921,N_29595,N_29400);
or UO_2922 (O_2922,N_29662,N_29827);
nor UO_2923 (O_2923,N_29687,N_29947);
xor UO_2924 (O_2924,N_29663,N_29669);
and UO_2925 (O_2925,N_29879,N_29790);
or UO_2926 (O_2926,N_29871,N_29880);
nor UO_2927 (O_2927,N_29616,N_29744);
nand UO_2928 (O_2928,N_29473,N_29645);
and UO_2929 (O_2929,N_29722,N_29604);
nor UO_2930 (O_2930,N_29719,N_29469);
nor UO_2931 (O_2931,N_29490,N_29744);
and UO_2932 (O_2932,N_29449,N_29518);
nor UO_2933 (O_2933,N_29584,N_29755);
nand UO_2934 (O_2934,N_29942,N_29828);
nor UO_2935 (O_2935,N_29890,N_29427);
nor UO_2936 (O_2936,N_29942,N_29989);
nor UO_2937 (O_2937,N_29643,N_29741);
xor UO_2938 (O_2938,N_29598,N_29721);
xor UO_2939 (O_2939,N_29763,N_29840);
or UO_2940 (O_2940,N_29609,N_29416);
and UO_2941 (O_2941,N_29646,N_29946);
nor UO_2942 (O_2942,N_29983,N_29478);
or UO_2943 (O_2943,N_29889,N_29741);
and UO_2944 (O_2944,N_29424,N_29630);
nand UO_2945 (O_2945,N_29433,N_29577);
nor UO_2946 (O_2946,N_29898,N_29709);
nand UO_2947 (O_2947,N_29598,N_29470);
nor UO_2948 (O_2948,N_29541,N_29481);
or UO_2949 (O_2949,N_29619,N_29977);
nand UO_2950 (O_2950,N_29822,N_29503);
nor UO_2951 (O_2951,N_29622,N_29677);
xor UO_2952 (O_2952,N_29634,N_29458);
and UO_2953 (O_2953,N_29633,N_29487);
and UO_2954 (O_2954,N_29984,N_29982);
and UO_2955 (O_2955,N_29748,N_29585);
xor UO_2956 (O_2956,N_29942,N_29489);
nand UO_2957 (O_2957,N_29809,N_29599);
nand UO_2958 (O_2958,N_29696,N_29506);
nor UO_2959 (O_2959,N_29813,N_29571);
nand UO_2960 (O_2960,N_29921,N_29601);
or UO_2961 (O_2961,N_29838,N_29945);
xnor UO_2962 (O_2962,N_29765,N_29691);
or UO_2963 (O_2963,N_29983,N_29818);
and UO_2964 (O_2964,N_29737,N_29401);
and UO_2965 (O_2965,N_29910,N_29914);
xor UO_2966 (O_2966,N_29960,N_29414);
xnor UO_2967 (O_2967,N_29774,N_29434);
nor UO_2968 (O_2968,N_29873,N_29915);
nor UO_2969 (O_2969,N_29835,N_29696);
or UO_2970 (O_2970,N_29507,N_29590);
and UO_2971 (O_2971,N_29811,N_29680);
nor UO_2972 (O_2972,N_29745,N_29672);
xor UO_2973 (O_2973,N_29628,N_29864);
xor UO_2974 (O_2974,N_29614,N_29791);
nor UO_2975 (O_2975,N_29715,N_29744);
nor UO_2976 (O_2976,N_29563,N_29404);
xor UO_2977 (O_2977,N_29416,N_29869);
nor UO_2978 (O_2978,N_29783,N_29687);
nand UO_2979 (O_2979,N_29794,N_29542);
or UO_2980 (O_2980,N_29893,N_29417);
xor UO_2981 (O_2981,N_29494,N_29892);
nand UO_2982 (O_2982,N_29697,N_29462);
nand UO_2983 (O_2983,N_29873,N_29767);
or UO_2984 (O_2984,N_29488,N_29937);
and UO_2985 (O_2985,N_29991,N_29829);
and UO_2986 (O_2986,N_29835,N_29679);
xnor UO_2987 (O_2987,N_29629,N_29461);
or UO_2988 (O_2988,N_29602,N_29814);
or UO_2989 (O_2989,N_29475,N_29433);
xor UO_2990 (O_2990,N_29480,N_29532);
or UO_2991 (O_2991,N_29640,N_29419);
or UO_2992 (O_2992,N_29836,N_29551);
or UO_2993 (O_2993,N_29488,N_29993);
nand UO_2994 (O_2994,N_29818,N_29928);
xor UO_2995 (O_2995,N_29823,N_29439);
nand UO_2996 (O_2996,N_29847,N_29580);
and UO_2997 (O_2997,N_29964,N_29786);
nand UO_2998 (O_2998,N_29581,N_29794);
nand UO_2999 (O_2999,N_29548,N_29632);
nor UO_3000 (O_3000,N_29750,N_29776);
nor UO_3001 (O_3001,N_29994,N_29617);
or UO_3002 (O_3002,N_29975,N_29722);
and UO_3003 (O_3003,N_29659,N_29542);
nand UO_3004 (O_3004,N_29933,N_29779);
nand UO_3005 (O_3005,N_29943,N_29605);
xor UO_3006 (O_3006,N_29594,N_29640);
and UO_3007 (O_3007,N_29872,N_29462);
or UO_3008 (O_3008,N_29805,N_29657);
nand UO_3009 (O_3009,N_29498,N_29878);
nand UO_3010 (O_3010,N_29852,N_29820);
nor UO_3011 (O_3011,N_29769,N_29845);
or UO_3012 (O_3012,N_29614,N_29463);
or UO_3013 (O_3013,N_29572,N_29799);
and UO_3014 (O_3014,N_29654,N_29811);
nand UO_3015 (O_3015,N_29511,N_29887);
nor UO_3016 (O_3016,N_29954,N_29475);
xnor UO_3017 (O_3017,N_29625,N_29798);
or UO_3018 (O_3018,N_29424,N_29499);
and UO_3019 (O_3019,N_29728,N_29499);
or UO_3020 (O_3020,N_29612,N_29924);
or UO_3021 (O_3021,N_29728,N_29434);
and UO_3022 (O_3022,N_29620,N_29743);
or UO_3023 (O_3023,N_29524,N_29403);
or UO_3024 (O_3024,N_29493,N_29624);
nor UO_3025 (O_3025,N_29420,N_29975);
nand UO_3026 (O_3026,N_29707,N_29745);
nor UO_3027 (O_3027,N_29484,N_29754);
nor UO_3028 (O_3028,N_29924,N_29589);
nor UO_3029 (O_3029,N_29691,N_29473);
nand UO_3030 (O_3030,N_29661,N_29407);
or UO_3031 (O_3031,N_29564,N_29837);
and UO_3032 (O_3032,N_29937,N_29649);
and UO_3033 (O_3033,N_29842,N_29784);
and UO_3034 (O_3034,N_29741,N_29412);
or UO_3035 (O_3035,N_29725,N_29553);
xnor UO_3036 (O_3036,N_29858,N_29494);
xnor UO_3037 (O_3037,N_29998,N_29663);
nor UO_3038 (O_3038,N_29821,N_29847);
nor UO_3039 (O_3039,N_29800,N_29967);
xnor UO_3040 (O_3040,N_29541,N_29755);
xor UO_3041 (O_3041,N_29925,N_29462);
xnor UO_3042 (O_3042,N_29626,N_29607);
nand UO_3043 (O_3043,N_29845,N_29511);
and UO_3044 (O_3044,N_29708,N_29462);
nand UO_3045 (O_3045,N_29835,N_29588);
or UO_3046 (O_3046,N_29488,N_29694);
xor UO_3047 (O_3047,N_29536,N_29717);
nor UO_3048 (O_3048,N_29806,N_29981);
xnor UO_3049 (O_3049,N_29826,N_29634);
xnor UO_3050 (O_3050,N_29950,N_29805);
or UO_3051 (O_3051,N_29610,N_29533);
nor UO_3052 (O_3052,N_29824,N_29897);
and UO_3053 (O_3053,N_29795,N_29546);
or UO_3054 (O_3054,N_29808,N_29723);
nand UO_3055 (O_3055,N_29686,N_29698);
and UO_3056 (O_3056,N_29404,N_29401);
nand UO_3057 (O_3057,N_29811,N_29616);
or UO_3058 (O_3058,N_29926,N_29632);
xnor UO_3059 (O_3059,N_29630,N_29592);
nor UO_3060 (O_3060,N_29572,N_29521);
or UO_3061 (O_3061,N_29549,N_29802);
or UO_3062 (O_3062,N_29475,N_29657);
and UO_3063 (O_3063,N_29897,N_29685);
or UO_3064 (O_3064,N_29900,N_29582);
and UO_3065 (O_3065,N_29597,N_29419);
nor UO_3066 (O_3066,N_29963,N_29547);
xnor UO_3067 (O_3067,N_29964,N_29753);
and UO_3068 (O_3068,N_29624,N_29965);
nor UO_3069 (O_3069,N_29658,N_29465);
nor UO_3070 (O_3070,N_29930,N_29757);
xor UO_3071 (O_3071,N_29926,N_29664);
nand UO_3072 (O_3072,N_29419,N_29599);
xnor UO_3073 (O_3073,N_29982,N_29722);
nand UO_3074 (O_3074,N_29850,N_29959);
xnor UO_3075 (O_3075,N_29679,N_29667);
or UO_3076 (O_3076,N_29800,N_29756);
nor UO_3077 (O_3077,N_29787,N_29886);
or UO_3078 (O_3078,N_29834,N_29849);
and UO_3079 (O_3079,N_29865,N_29781);
nor UO_3080 (O_3080,N_29816,N_29483);
xor UO_3081 (O_3081,N_29839,N_29898);
and UO_3082 (O_3082,N_29860,N_29656);
nor UO_3083 (O_3083,N_29691,N_29449);
or UO_3084 (O_3084,N_29436,N_29917);
nand UO_3085 (O_3085,N_29682,N_29996);
nor UO_3086 (O_3086,N_29873,N_29954);
or UO_3087 (O_3087,N_29899,N_29822);
xor UO_3088 (O_3088,N_29706,N_29558);
nor UO_3089 (O_3089,N_29645,N_29988);
and UO_3090 (O_3090,N_29508,N_29604);
xnor UO_3091 (O_3091,N_29732,N_29806);
nor UO_3092 (O_3092,N_29405,N_29946);
nand UO_3093 (O_3093,N_29992,N_29513);
xnor UO_3094 (O_3094,N_29999,N_29727);
xor UO_3095 (O_3095,N_29515,N_29783);
nor UO_3096 (O_3096,N_29876,N_29742);
or UO_3097 (O_3097,N_29644,N_29424);
xor UO_3098 (O_3098,N_29929,N_29937);
nand UO_3099 (O_3099,N_29853,N_29738);
and UO_3100 (O_3100,N_29728,N_29436);
or UO_3101 (O_3101,N_29860,N_29635);
nor UO_3102 (O_3102,N_29771,N_29512);
or UO_3103 (O_3103,N_29684,N_29468);
xnor UO_3104 (O_3104,N_29959,N_29974);
or UO_3105 (O_3105,N_29476,N_29712);
nand UO_3106 (O_3106,N_29481,N_29929);
and UO_3107 (O_3107,N_29735,N_29668);
xnor UO_3108 (O_3108,N_29710,N_29714);
or UO_3109 (O_3109,N_29980,N_29717);
nand UO_3110 (O_3110,N_29756,N_29623);
or UO_3111 (O_3111,N_29830,N_29457);
nand UO_3112 (O_3112,N_29513,N_29471);
or UO_3113 (O_3113,N_29812,N_29806);
or UO_3114 (O_3114,N_29750,N_29961);
xor UO_3115 (O_3115,N_29583,N_29900);
nand UO_3116 (O_3116,N_29614,N_29574);
nor UO_3117 (O_3117,N_29699,N_29848);
nor UO_3118 (O_3118,N_29836,N_29911);
or UO_3119 (O_3119,N_29408,N_29945);
nand UO_3120 (O_3120,N_29720,N_29479);
or UO_3121 (O_3121,N_29566,N_29753);
and UO_3122 (O_3122,N_29458,N_29911);
nand UO_3123 (O_3123,N_29585,N_29991);
nor UO_3124 (O_3124,N_29554,N_29839);
nor UO_3125 (O_3125,N_29978,N_29802);
and UO_3126 (O_3126,N_29415,N_29919);
nor UO_3127 (O_3127,N_29996,N_29412);
or UO_3128 (O_3128,N_29448,N_29751);
or UO_3129 (O_3129,N_29530,N_29780);
or UO_3130 (O_3130,N_29455,N_29553);
xnor UO_3131 (O_3131,N_29466,N_29528);
nand UO_3132 (O_3132,N_29726,N_29950);
xnor UO_3133 (O_3133,N_29778,N_29513);
nand UO_3134 (O_3134,N_29695,N_29733);
xnor UO_3135 (O_3135,N_29457,N_29657);
nand UO_3136 (O_3136,N_29669,N_29892);
nand UO_3137 (O_3137,N_29468,N_29415);
or UO_3138 (O_3138,N_29954,N_29510);
and UO_3139 (O_3139,N_29852,N_29558);
nand UO_3140 (O_3140,N_29589,N_29713);
xor UO_3141 (O_3141,N_29668,N_29564);
xor UO_3142 (O_3142,N_29886,N_29837);
or UO_3143 (O_3143,N_29934,N_29444);
xnor UO_3144 (O_3144,N_29900,N_29929);
xor UO_3145 (O_3145,N_29809,N_29716);
or UO_3146 (O_3146,N_29524,N_29476);
or UO_3147 (O_3147,N_29815,N_29455);
nand UO_3148 (O_3148,N_29699,N_29713);
or UO_3149 (O_3149,N_29911,N_29897);
nand UO_3150 (O_3150,N_29845,N_29763);
nand UO_3151 (O_3151,N_29444,N_29458);
or UO_3152 (O_3152,N_29696,N_29889);
and UO_3153 (O_3153,N_29676,N_29856);
or UO_3154 (O_3154,N_29570,N_29968);
or UO_3155 (O_3155,N_29957,N_29712);
nand UO_3156 (O_3156,N_29467,N_29554);
nand UO_3157 (O_3157,N_29962,N_29463);
xnor UO_3158 (O_3158,N_29624,N_29834);
xnor UO_3159 (O_3159,N_29793,N_29685);
nand UO_3160 (O_3160,N_29993,N_29709);
and UO_3161 (O_3161,N_29843,N_29532);
nor UO_3162 (O_3162,N_29733,N_29696);
nor UO_3163 (O_3163,N_29788,N_29838);
nand UO_3164 (O_3164,N_29417,N_29593);
or UO_3165 (O_3165,N_29990,N_29915);
and UO_3166 (O_3166,N_29560,N_29643);
xnor UO_3167 (O_3167,N_29637,N_29401);
and UO_3168 (O_3168,N_29428,N_29731);
nor UO_3169 (O_3169,N_29734,N_29635);
and UO_3170 (O_3170,N_29565,N_29962);
nand UO_3171 (O_3171,N_29429,N_29947);
and UO_3172 (O_3172,N_29564,N_29598);
nor UO_3173 (O_3173,N_29855,N_29719);
or UO_3174 (O_3174,N_29667,N_29440);
nand UO_3175 (O_3175,N_29681,N_29466);
nor UO_3176 (O_3176,N_29980,N_29591);
and UO_3177 (O_3177,N_29675,N_29815);
nor UO_3178 (O_3178,N_29948,N_29704);
nor UO_3179 (O_3179,N_29623,N_29661);
nor UO_3180 (O_3180,N_29772,N_29721);
xor UO_3181 (O_3181,N_29812,N_29799);
nand UO_3182 (O_3182,N_29932,N_29577);
xor UO_3183 (O_3183,N_29695,N_29696);
xnor UO_3184 (O_3184,N_29670,N_29407);
or UO_3185 (O_3185,N_29945,N_29940);
nor UO_3186 (O_3186,N_29631,N_29427);
xor UO_3187 (O_3187,N_29424,N_29978);
xnor UO_3188 (O_3188,N_29498,N_29642);
and UO_3189 (O_3189,N_29575,N_29425);
nor UO_3190 (O_3190,N_29885,N_29584);
xnor UO_3191 (O_3191,N_29782,N_29960);
nor UO_3192 (O_3192,N_29805,N_29746);
xor UO_3193 (O_3193,N_29841,N_29958);
nor UO_3194 (O_3194,N_29511,N_29954);
or UO_3195 (O_3195,N_29910,N_29601);
and UO_3196 (O_3196,N_29476,N_29425);
xor UO_3197 (O_3197,N_29842,N_29546);
xor UO_3198 (O_3198,N_29465,N_29537);
xnor UO_3199 (O_3199,N_29941,N_29610);
xnor UO_3200 (O_3200,N_29621,N_29553);
or UO_3201 (O_3201,N_29423,N_29853);
xor UO_3202 (O_3202,N_29836,N_29540);
and UO_3203 (O_3203,N_29641,N_29531);
xor UO_3204 (O_3204,N_29792,N_29563);
nor UO_3205 (O_3205,N_29630,N_29457);
nor UO_3206 (O_3206,N_29814,N_29815);
nor UO_3207 (O_3207,N_29515,N_29614);
and UO_3208 (O_3208,N_29510,N_29802);
nor UO_3209 (O_3209,N_29829,N_29428);
or UO_3210 (O_3210,N_29464,N_29670);
nand UO_3211 (O_3211,N_29984,N_29875);
xor UO_3212 (O_3212,N_29485,N_29554);
xor UO_3213 (O_3213,N_29893,N_29413);
xnor UO_3214 (O_3214,N_29859,N_29740);
nand UO_3215 (O_3215,N_29865,N_29734);
xnor UO_3216 (O_3216,N_29646,N_29841);
nor UO_3217 (O_3217,N_29418,N_29814);
nor UO_3218 (O_3218,N_29420,N_29463);
xnor UO_3219 (O_3219,N_29592,N_29485);
and UO_3220 (O_3220,N_29622,N_29468);
nor UO_3221 (O_3221,N_29762,N_29522);
xnor UO_3222 (O_3222,N_29596,N_29405);
nor UO_3223 (O_3223,N_29844,N_29784);
nor UO_3224 (O_3224,N_29546,N_29635);
nor UO_3225 (O_3225,N_29710,N_29597);
and UO_3226 (O_3226,N_29751,N_29789);
nor UO_3227 (O_3227,N_29773,N_29966);
and UO_3228 (O_3228,N_29822,N_29988);
or UO_3229 (O_3229,N_29778,N_29970);
nor UO_3230 (O_3230,N_29829,N_29749);
xor UO_3231 (O_3231,N_29709,N_29776);
xnor UO_3232 (O_3232,N_29802,N_29963);
xnor UO_3233 (O_3233,N_29839,N_29902);
and UO_3234 (O_3234,N_29777,N_29823);
xnor UO_3235 (O_3235,N_29433,N_29730);
xnor UO_3236 (O_3236,N_29829,N_29936);
nand UO_3237 (O_3237,N_29419,N_29858);
nor UO_3238 (O_3238,N_29445,N_29545);
xor UO_3239 (O_3239,N_29680,N_29739);
xnor UO_3240 (O_3240,N_29992,N_29912);
and UO_3241 (O_3241,N_29576,N_29409);
nand UO_3242 (O_3242,N_29746,N_29570);
nor UO_3243 (O_3243,N_29553,N_29970);
nand UO_3244 (O_3244,N_29596,N_29557);
xor UO_3245 (O_3245,N_29557,N_29485);
or UO_3246 (O_3246,N_29612,N_29595);
or UO_3247 (O_3247,N_29997,N_29574);
and UO_3248 (O_3248,N_29846,N_29750);
xnor UO_3249 (O_3249,N_29862,N_29696);
nor UO_3250 (O_3250,N_29741,N_29694);
xnor UO_3251 (O_3251,N_29563,N_29682);
nand UO_3252 (O_3252,N_29843,N_29967);
nor UO_3253 (O_3253,N_29513,N_29510);
xor UO_3254 (O_3254,N_29609,N_29627);
and UO_3255 (O_3255,N_29516,N_29844);
nor UO_3256 (O_3256,N_29611,N_29659);
xnor UO_3257 (O_3257,N_29427,N_29493);
nand UO_3258 (O_3258,N_29502,N_29892);
xor UO_3259 (O_3259,N_29550,N_29564);
nand UO_3260 (O_3260,N_29778,N_29664);
and UO_3261 (O_3261,N_29422,N_29630);
xnor UO_3262 (O_3262,N_29918,N_29744);
nand UO_3263 (O_3263,N_29913,N_29455);
and UO_3264 (O_3264,N_29842,N_29523);
nand UO_3265 (O_3265,N_29980,N_29672);
nand UO_3266 (O_3266,N_29748,N_29777);
and UO_3267 (O_3267,N_29408,N_29633);
xnor UO_3268 (O_3268,N_29975,N_29896);
or UO_3269 (O_3269,N_29713,N_29496);
nor UO_3270 (O_3270,N_29581,N_29669);
nor UO_3271 (O_3271,N_29816,N_29890);
and UO_3272 (O_3272,N_29627,N_29928);
or UO_3273 (O_3273,N_29605,N_29770);
nor UO_3274 (O_3274,N_29583,N_29424);
and UO_3275 (O_3275,N_29577,N_29757);
nand UO_3276 (O_3276,N_29879,N_29761);
nor UO_3277 (O_3277,N_29788,N_29415);
xnor UO_3278 (O_3278,N_29806,N_29778);
and UO_3279 (O_3279,N_29765,N_29990);
nor UO_3280 (O_3280,N_29930,N_29875);
and UO_3281 (O_3281,N_29828,N_29733);
nor UO_3282 (O_3282,N_29442,N_29921);
or UO_3283 (O_3283,N_29688,N_29967);
nand UO_3284 (O_3284,N_29595,N_29474);
xor UO_3285 (O_3285,N_29418,N_29416);
xor UO_3286 (O_3286,N_29675,N_29646);
and UO_3287 (O_3287,N_29495,N_29624);
xnor UO_3288 (O_3288,N_29489,N_29437);
xnor UO_3289 (O_3289,N_29495,N_29404);
or UO_3290 (O_3290,N_29564,N_29430);
xnor UO_3291 (O_3291,N_29512,N_29700);
nand UO_3292 (O_3292,N_29823,N_29559);
xnor UO_3293 (O_3293,N_29761,N_29785);
and UO_3294 (O_3294,N_29445,N_29850);
nand UO_3295 (O_3295,N_29436,N_29859);
xnor UO_3296 (O_3296,N_29622,N_29730);
nor UO_3297 (O_3297,N_29683,N_29963);
and UO_3298 (O_3298,N_29432,N_29648);
nor UO_3299 (O_3299,N_29767,N_29666);
nand UO_3300 (O_3300,N_29660,N_29771);
nor UO_3301 (O_3301,N_29920,N_29971);
nand UO_3302 (O_3302,N_29891,N_29689);
xnor UO_3303 (O_3303,N_29823,N_29432);
and UO_3304 (O_3304,N_29919,N_29522);
xor UO_3305 (O_3305,N_29847,N_29952);
nand UO_3306 (O_3306,N_29555,N_29413);
and UO_3307 (O_3307,N_29796,N_29979);
or UO_3308 (O_3308,N_29893,N_29759);
or UO_3309 (O_3309,N_29920,N_29679);
or UO_3310 (O_3310,N_29637,N_29706);
or UO_3311 (O_3311,N_29567,N_29776);
or UO_3312 (O_3312,N_29897,N_29989);
xor UO_3313 (O_3313,N_29756,N_29673);
xor UO_3314 (O_3314,N_29772,N_29936);
xor UO_3315 (O_3315,N_29403,N_29620);
nor UO_3316 (O_3316,N_29973,N_29665);
nand UO_3317 (O_3317,N_29772,N_29735);
nor UO_3318 (O_3318,N_29449,N_29617);
nor UO_3319 (O_3319,N_29719,N_29852);
nor UO_3320 (O_3320,N_29748,N_29525);
and UO_3321 (O_3321,N_29403,N_29802);
xnor UO_3322 (O_3322,N_29652,N_29839);
or UO_3323 (O_3323,N_29866,N_29419);
xnor UO_3324 (O_3324,N_29931,N_29625);
and UO_3325 (O_3325,N_29903,N_29439);
xor UO_3326 (O_3326,N_29973,N_29860);
nand UO_3327 (O_3327,N_29624,N_29569);
nor UO_3328 (O_3328,N_29984,N_29981);
nor UO_3329 (O_3329,N_29912,N_29922);
and UO_3330 (O_3330,N_29998,N_29771);
nand UO_3331 (O_3331,N_29886,N_29457);
or UO_3332 (O_3332,N_29637,N_29631);
xor UO_3333 (O_3333,N_29652,N_29894);
nor UO_3334 (O_3334,N_29932,N_29457);
xor UO_3335 (O_3335,N_29834,N_29734);
nor UO_3336 (O_3336,N_29990,N_29851);
nor UO_3337 (O_3337,N_29618,N_29539);
and UO_3338 (O_3338,N_29934,N_29876);
or UO_3339 (O_3339,N_29495,N_29448);
or UO_3340 (O_3340,N_29607,N_29715);
and UO_3341 (O_3341,N_29777,N_29672);
xnor UO_3342 (O_3342,N_29648,N_29441);
xnor UO_3343 (O_3343,N_29614,N_29427);
nand UO_3344 (O_3344,N_29830,N_29612);
or UO_3345 (O_3345,N_29732,N_29815);
xnor UO_3346 (O_3346,N_29715,N_29780);
or UO_3347 (O_3347,N_29758,N_29991);
nor UO_3348 (O_3348,N_29626,N_29441);
nand UO_3349 (O_3349,N_29680,N_29979);
and UO_3350 (O_3350,N_29731,N_29439);
nand UO_3351 (O_3351,N_29571,N_29793);
nand UO_3352 (O_3352,N_29631,N_29922);
nand UO_3353 (O_3353,N_29527,N_29989);
or UO_3354 (O_3354,N_29936,N_29974);
nand UO_3355 (O_3355,N_29673,N_29461);
nor UO_3356 (O_3356,N_29994,N_29726);
xnor UO_3357 (O_3357,N_29819,N_29845);
or UO_3358 (O_3358,N_29872,N_29463);
and UO_3359 (O_3359,N_29479,N_29400);
or UO_3360 (O_3360,N_29418,N_29857);
nand UO_3361 (O_3361,N_29857,N_29922);
or UO_3362 (O_3362,N_29836,N_29717);
or UO_3363 (O_3363,N_29556,N_29847);
xnor UO_3364 (O_3364,N_29482,N_29569);
nor UO_3365 (O_3365,N_29623,N_29792);
or UO_3366 (O_3366,N_29976,N_29752);
xor UO_3367 (O_3367,N_29926,N_29643);
or UO_3368 (O_3368,N_29989,N_29979);
or UO_3369 (O_3369,N_29977,N_29745);
nand UO_3370 (O_3370,N_29819,N_29867);
or UO_3371 (O_3371,N_29655,N_29510);
xnor UO_3372 (O_3372,N_29499,N_29854);
xnor UO_3373 (O_3373,N_29590,N_29425);
nor UO_3374 (O_3374,N_29497,N_29965);
and UO_3375 (O_3375,N_29777,N_29985);
xnor UO_3376 (O_3376,N_29920,N_29869);
xnor UO_3377 (O_3377,N_29939,N_29409);
nor UO_3378 (O_3378,N_29821,N_29875);
nand UO_3379 (O_3379,N_29911,N_29775);
or UO_3380 (O_3380,N_29547,N_29676);
or UO_3381 (O_3381,N_29516,N_29494);
xnor UO_3382 (O_3382,N_29515,N_29667);
and UO_3383 (O_3383,N_29802,N_29443);
or UO_3384 (O_3384,N_29407,N_29792);
nand UO_3385 (O_3385,N_29725,N_29848);
nand UO_3386 (O_3386,N_29937,N_29553);
or UO_3387 (O_3387,N_29716,N_29869);
nand UO_3388 (O_3388,N_29493,N_29847);
nand UO_3389 (O_3389,N_29743,N_29403);
nor UO_3390 (O_3390,N_29660,N_29450);
or UO_3391 (O_3391,N_29574,N_29745);
xor UO_3392 (O_3392,N_29431,N_29528);
nand UO_3393 (O_3393,N_29658,N_29769);
or UO_3394 (O_3394,N_29503,N_29504);
xor UO_3395 (O_3395,N_29644,N_29986);
and UO_3396 (O_3396,N_29986,N_29748);
or UO_3397 (O_3397,N_29741,N_29423);
or UO_3398 (O_3398,N_29589,N_29569);
nand UO_3399 (O_3399,N_29443,N_29629);
xor UO_3400 (O_3400,N_29456,N_29775);
nor UO_3401 (O_3401,N_29819,N_29900);
nor UO_3402 (O_3402,N_29730,N_29451);
and UO_3403 (O_3403,N_29846,N_29953);
and UO_3404 (O_3404,N_29473,N_29481);
xor UO_3405 (O_3405,N_29949,N_29908);
nand UO_3406 (O_3406,N_29782,N_29484);
xor UO_3407 (O_3407,N_29560,N_29703);
or UO_3408 (O_3408,N_29786,N_29566);
or UO_3409 (O_3409,N_29852,N_29936);
nor UO_3410 (O_3410,N_29437,N_29418);
and UO_3411 (O_3411,N_29414,N_29672);
xnor UO_3412 (O_3412,N_29765,N_29675);
nor UO_3413 (O_3413,N_29994,N_29443);
or UO_3414 (O_3414,N_29600,N_29612);
xor UO_3415 (O_3415,N_29617,N_29997);
xnor UO_3416 (O_3416,N_29922,N_29565);
nand UO_3417 (O_3417,N_29846,N_29546);
or UO_3418 (O_3418,N_29619,N_29907);
nor UO_3419 (O_3419,N_29998,N_29657);
xor UO_3420 (O_3420,N_29591,N_29991);
and UO_3421 (O_3421,N_29487,N_29694);
nand UO_3422 (O_3422,N_29763,N_29779);
and UO_3423 (O_3423,N_29814,N_29880);
nor UO_3424 (O_3424,N_29442,N_29621);
nor UO_3425 (O_3425,N_29987,N_29669);
or UO_3426 (O_3426,N_29931,N_29646);
and UO_3427 (O_3427,N_29481,N_29746);
nor UO_3428 (O_3428,N_29668,N_29552);
xor UO_3429 (O_3429,N_29554,N_29493);
nand UO_3430 (O_3430,N_29462,N_29871);
or UO_3431 (O_3431,N_29870,N_29458);
xor UO_3432 (O_3432,N_29596,N_29800);
and UO_3433 (O_3433,N_29407,N_29526);
nor UO_3434 (O_3434,N_29726,N_29610);
nor UO_3435 (O_3435,N_29465,N_29433);
xnor UO_3436 (O_3436,N_29424,N_29719);
nor UO_3437 (O_3437,N_29697,N_29888);
or UO_3438 (O_3438,N_29710,N_29566);
and UO_3439 (O_3439,N_29926,N_29461);
xor UO_3440 (O_3440,N_29953,N_29571);
nor UO_3441 (O_3441,N_29510,N_29729);
xnor UO_3442 (O_3442,N_29637,N_29667);
and UO_3443 (O_3443,N_29592,N_29873);
or UO_3444 (O_3444,N_29680,N_29838);
and UO_3445 (O_3445,N_29851,N_29537);
xor UO_3446 (O_3446,N_29781,N_29549);
and UO_3447 (O_3447,N_29766,N_29429);
or UO_3448 (O_3448,N_29830,N_29817);
xor UO_3449 (O_3449,N_29657,N_29781);
or UO_3450 (O_3450,N_29966,N_29755);
xor UO_3451 (O_3451,N_29643,N_29911);
or UO_3452 (O_3452,N_29522,N_29932);
and UO_3453 (O_3453,N_29465,N_29705);
or UO_3454 (O_3454,N_29843,N_29530);
and UO_3455 (O_3455,N_29454,N_29700);
xnor UO_3456 (O_3456,N_29985,N_29755);
and UO_3457 (O_3457,N_29490,N_29683);
xor UO_3458 (O_3458,N_29726,N_29480);
or UO_3459 (O_3459,N_29885,N_29454);
or UO_3460 (O_3460,N_29522,N_29523);
nand UO_3461 (O_3461,N_29574,N_29703);
nand UO_3462 (O_3462,N_29598,N_29829);
nand UO_3463 (O_3463,N_29621,N_29526);
xor UO_3464 (O_3464,N_29531,N_29667);
nand UO_3465 (O_3465,N_29430,N_29615);
or UO_3466 (O_3466,N_29532,N_29886);
and UO_3467 (O_3467,N_29954,N_29459);
nor UO_3468 (O_3468,N_29984,N_29800);
and UO_3469 (O_3469,N_29770,N_29815);
or UO_3470 (O_3470,N_29737,N_29878);
or UO_3471 (O_3471,N_29962,N_29736);
nor UO_3472 (O_3472,N_29701,N_29494);
nor UO_3473 (O_3473,N_29844,N_29616);
nor UO_3474 (O_3474,N_29824,N_29957);
or UO_3475 (O_3475,N_29616,N_29746);
xnor UO_3476 (O_3476,N_29837,N_29724);
or UO_3477 (O_3477,N_29915,N_29994);
nor UO_3478 (O_3478,N_29590,N_29479);
xor UO_3479 (O_3479,N_29984,N_29764);
and UO_3480 (O_3480,N_29627,N_29623);
or UO_3481 (O_3481,N_29775,N_29515);
xor UO_3482 (O_3482,N_29868,N_29587);
and UO_3483 (O_3483,N_29675,N_29919);
nand UO_3484 (O_3484,N_29500,N_29909);
nand UO_3485 (O_3485,N_29452,N_29801);
xor UO_3486 (O_3486,N_29572,N_29981);
and UO_3487 (O_3487,N_29974,N_29731);
xnor UO_3488 (O_3488,N_29493,N_29641);
and UO_3489 (O_3489,N_29717,N_29780);
nand UO_3490 (O_3490,N_29784,N_29514);
and UO_3491 (O_3491,N_29767,N_29444);
nor UO_3492 (O_3492,N_29976,N_29942);
nor UO_3493 (O_3493,N_29436,N_29524);
xor UO_3494 (O_3494,N_29687,N_29689);
nand UO_3495 (O_3495,N_29954,N_29919);
nor UO_3496 (O_3496,N_29875,N_29628);
nor UO_3497 (O_3497,N_29953,N_29904);
nand UO_3498 (O_3498,N_29496,N_29880);
xnor UO_3499 (O_3499,N_29451,N_29580);
endmodule