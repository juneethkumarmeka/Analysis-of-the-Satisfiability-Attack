module basic_3000_30000_3500_20_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2415,In_2464);
and U1 (N_1,In_2651,In_1142);
xor U2 (N_2,In_2525,In_1978);
xor U3 (N_3,In_496,In_2609);
xor U4 (N_4,In_1992,In_272);
nor U5 (N_5,In_1257,In_1459);
or U6 (N_6,In_1860,In_167);
nand U7 (N_7,In_2985,In_2532);
nor U8 (N_8,In_1116,In_2219);
xor U9 (N_9,In_824,In_1621);
nand U10 (N_10,In_2167,In_2437);
nor U11 (N_11,In_829,In_1668);
and U12 (N_12,In_2090,In_90);
xnor U13 (N_13,In_1593,In_2519);
nor U14 (N_14,In_1895,In_1087);
nor U15 (N_15,In_1080,In_1383);
xor U16 (N_16,In_2199,In_2150);
xor U17 (N_17,In_1690,In_2014);
nand U18 (N_18,In_2121,In_1039);
or U19 (N_19,In_83,In_1029);
or U20 (N_20,In_1477,In_2367);
xor U21 (N_21,In_528,In_1340);
nand U22 (N_22,In_371,In_2189);
or U23 (N_23,In_361,In_970);
nor U24 (N_24,In_2620,In_2416);
and U25 (N_25,In_2796,In_1289);
xor U26 (N_26,In_1034,In_20);
or U27 (N_27,In_2716,In_2473);
and U28 (N_28,In_1191,In_1872);
or U29 (N_29,In_240,In_2173);
xnor U30 (N_30,In_750,In_2029);
and U31 (N_31,In_2541,In_2535);
nand U32 (N_32,In_165,In_980);
nand U33 (N_33,In_955,In_1336);
and U34 (N_34,In_954,In_300);
nand U35 (N_35,In_435,In_1238);
nand U36 (N_36,In_1792,In_2152);
and U37 (N_37,In_2075,In_2583);
nor U38 (N_38,In_1414,In_1758);
nand U39 (N_39,In_781,In_357);
nor U40 (N_40,In_2952,In_879);
and U41 (N_41,In_376,In_506);
xor U42 (N_42,In_410,In_1879);
xnor U43 (N_43,In_2986,In_2607);
xnor U44 (N_44,In_1045,In_2166);
xnor U45 (N_45,In_2487,In_893);
xor U46 (N_46,In_1568,In_2310);
nor U47 (N_47,In_859,In_2264);
or U48 (N_48,In_951,In_734);
and U49 (N_49,In_624,In_2270);
nand U50 (N_50,In_1762,In_2263);
or U51 (N_51,In_2844,In_521);
nor U52 (N_52,In_1181,In_1741);
or U53 (N_53,In_906,In_1436);
xnor U54 (N_54,In_1241,In_1352);
or U55 (N_55,In_424,In_749);
xor U56 (N_56,In_1102,In_1749);
xor U57 (N_57,In_159,In_2703);
nand U58 (N_58,In_2035,In_321);
nor U59 (N_59,In_867,In_996);
xor U60 (N_60,In_2718,In_785);
nor U61 (N_61,In_229,In_2223);
or U62 (N_62,In_2436,In_2808);
or U63 (N_63,In_1986,In_641);
or U64 (N_64,In_2559,In_655);
and U65 (N_65,In_2929,In_1524);
nand U66 (N_66,In_1864,In_1255);
xnor U67 (N_67,In_1491,In_369);
and U68 (N_68,In_1313,In_2771);
nand U69 (N_69,In_2863,In_149);
nand U70 (N_70,In_2504,In_80);
nor U71 (N_71,In_929,In_1398);
nor U72 (N_72,In_504,In_467);
and U73 (N_73,In_2719,In_2721);
xnor U74 (N_74,In_349,In_1458);
and U75 (N_75,In_779,In_1595);
nand U76 (N_76,In_2474,In_112);
and U77 (N_77,In_2755,In_739);
or U78 (N_78,In_1721,In_2048);
nor U79 (N_79,In_869,In_2563);
and U80 (N_80,In_1615,In_604);
nand U81 (N_81,In_2763,In_156);
nand U82 (N_82,In_2632,In_146);
nor U83 (N_83,In_1553,In_1552);
nand U84 (N_84,In_2873,In_65);
or U85 (N_85,In_2492,In_1789);
nor U86 (N_86,In_1780,In_2480);
nor U87 (N_87,In_1226,In_1334);
or U88 (N_88,In_1567,In_1331);
or U89 (N_89,In_1820,In_1058);
nand U90 (N_90,In_2656,In_540);
nand U91 (N_91,In_350,In_1307);
nor U92 (N_92,In_2300,In_302);
nand U93 (N_93,In_441,In_1966);
nor U94 (N_94,In_1543,In_2281);
nor U95 (N_95,In_649,In_132);
nor U96 (N_96,In_296,In_2979);
or U97 (N_97,In_2700,In_2671);
or U98 (N_98,In_714,In_2936);
and U99 (N_99,In_1400,In_2477);
nor U100 (N_100,In_2858,In_284);
xor U101 (N_101,In_987,In_21);
or U102 (N_102,In_831,In_2241);
and U103 (N_103,In_194,In_2764);
nand U104 (N_104,In_742,In_2829);
or U105 (N_105,In_1127,In_2137);
xnor U106 (N_106,In_2413,In_2289);
or U107 (N_107,In_861,In_1017);
nor U108 (N_108,In_1756,In_481);
or U109 (N_109,In_1627,In_319);
nor U110 (N_110,In_1773,In_351);
or U111 (N_111,In_1151,In_418);
xor U112 (N_112,In_1107,In_2951);
and U113 (N_113,In_2694,In_2809);
nor U114 (N_114,In_193,In_2811);
or U115 (N_115,In_1246,In_2548);
nor U116 (N_116,In_1767,In_1369);
and U117 (N_117,In_1139,In_2142);
nor U118 (N_118,In_1440,In_2795);
or U119 (N_119,In_2455,In_1924);
nor U120 (N_120,In_2364,In_1394);
nor U121 (N_121,In_735,In_1382);
nor U122 (N_122,In_2186,In_2523);
nand U123 (N_123,In_1551,In_1222);
and U124 (N_124,In_2080,In_698);
nor U125 (N_125,In_775,In_1613);
nor U126 (N_126,In_2328,In_2370);
nand U127 (N_127,In_2698,In_32);
and U128 (N_128,In_2648,In_140);
nand U129 (N_129,In_1363,In_1884);
nand U130 (N_130,In_1731,In_789);
or U131 (N_131,In_1434,In_2418);
or U132 (N_132,In_258,In_2557);
nand U133 (N_133,In_2439,In_2115);
or U134 (N_134,In_2044,In_638);
xor U135 (N_135,In_283,In_646);
nor U136 (N_136,In_513,In_458);
xor U137 (N_137,In_2383,In_2365);
nor U138 (N_138,In_1694,In_2999);
or U139 (N_139,In_1625,In_898);
xnor U140 (N_140,In_1735,In_1566);
and U141 (N_141,In_2012,In_1512);
or U142 (N_142,In_1252,In_1957);
xnor U143 (N_143,In_2200,In_2468);
nor U144 (N_144,In_1371,In_2513);
nand U145 (N_145,In_1299,In_1320);
nand U146 (N_146,In_2720,In_812);
and U147 (N_147,In_1120,In_2807);
nand U148 (N_148,In_1947,In_1486);
or U149 (N_149,In_56,In_2838);
nor U150 (N_150,In_2560,In_2944);
nand U151 (N_151,In_1411,In_596);
and U152 (N_152,In_2256,In_787);
xor U153 (N_153,In_1189,In_515);
nor U154 (N_154,In_2091,In_136);
nor U155 (N_155,In_1955,In_1048);
nand U156 (N_156,In_423,In_723);
or U157 (N_157,In_1559,In_1921);
or U158 (N_158,In_877,In_1215);
nor U159 (N_159,In_1739,In_172);
xor U160 (N_160,In_2537,In_1023);
nor U161 (N_161,In_1090,In_634);
or U162 (N_162,In_1798,In_1545);
nor U163 (N_163,In_2063,In_607);
xor U164 (N_164,In_2987,In_1304);
or U165 (N_165,In_2258,In_1272);
nand U166 (N_166,In_1032,In_1072);
xnor U167 (N_167,In_2597,In_131);
nand U168 (N_168,In_177,In_2023);
and U169 (N_169,In_1790,In_2351);
nor U170 (N_170,In_91,In_1569);
xnor U171 (N_171,In_2687,In_1496);
nand U172 (N_172,In_2736,In_820);
nand U173 (N_173,In_87,In_2382);
nor U174 (N_174,In_2295,In_1687);
nand U175 (N_175,In_364,In_1135);
or U176 (N_176,In_817,In_765);
nor U177 (N_177,In_1943,In_1963);
or U178 (N_178,In_2613,In_1609);
xnor U179 (N_179,In_2627,In_1092);
nand U180 (N_180,In_1168,In_348);
and U181 (N_181,In_1649,In_2884);
nor U182 (N_182,In_2950,In_1285);
nor U183 (N_183,In_1244,In_2512);
or U184 (N_184,In_1404,In_2376);
nor U185 (N_185,In_850,In_1532);
nor U186 (N_186,In_1565,In_1103);
nand U187 (N_187,In_2830,In_715);
nor U188 (N_188,In_1323,In_292);
and U189 (N_189,In_205,In_168);
nand U190 (N_190,In_1097,In_262);
or U191 (N_191,In_1817,In_2397);
nand U192 (N_192,In_1281,In_1204);
nor U193 (N_193,In_1321,In_2545);
nor U194 (N_194,In_2742,In_2184);
and U195 (N_195,In_2686,In_396);
or U196 (N_196,In_2068,In_1347);
xor U197 (N_197,In_1044,In_397);
xnor U198 (N_198,In_1522,In_1732);
nand U199 (N_199,In_1852,In_203);
nand U200 (N_200,In_678,In_39);
nand U201 (N_201,In_886,In_1647);
and U202 (N_202,In_1905,In_416);
xor U203 (N_203,In_2488,In_2723);
and U204 (N_204,In_1046,In_2888);
xnor U205 (N_205,In_2288,In_625);
or U206 (N_206,In_958,In_1010);
xor U207 (N_207,In_2959,In_677);
xor U208 (N_208,In_1591,In_2814);
xnor U209 (N_209,In_1855,In_552);
and U210 (N_210,In_2840,In_1501);
nand U211 (N_211,In_2566,In_238);
nand U212 (N_212,In_1209,In_2816);
nand U213 (N_213,In_2965,In_64);
nand U214 (N_214,In_2362,In_1482);
nand U215 (N_215,In_531,In_1502);
nor U216 (N_216,In_2041,In_2308);
and U217 (N_217,In_2089,In_1796);
and U218 (N_218,In_58,In_395);
nor U219 (N_219,In_598,In_2332);
nand U220 (N_220,In_135,In_720);
and U221 (N_221,In_2336,In_3);
and U222 (N_222,In_702,In_2193);
xor U223 (N_223,In_1348,In_1799);
nand U224 (N_224,In_1013,In_414);
or U225 (N_225,In_727,In_2253);
nor U226 (N_226,In_288,In_1920);
nand U227 (N_227,In_1991,In_476);
or U228 (N_228,In_2564,In_672);
xor U229 (N_229,In_780,In_161);
xor U230 (N_230,In_196,In_553);
and U231 (N_231,In_1133,In_2805);
xor U232 (N_232,In_470,In_1717);
nand U233 (N_233,In_2653,In_926);
xnor U234 (N_234,In_1406,In_991);
or U235 (N_235,In_557,In_1607);
nand U236 (N_236,In_1779,In_129);
nor U237 (N_237,In_108,In_1385);
nand U238 (N_238,In_24,In_1787);
xor U239 (N_239,In_276,In_2096);
or U240 (N_240,In_1936,In_2897);
and U241 (N_241,In_2502,In_1112);
and U242 (N_242,In_2003,In_662);
nand U243 (N_243,In_643,In_1068);
or U244 (N_244,In_1581,In_2961);
or U245 (N_245,In_335,In_851);
xnor U246 (N_246,In_706,In_964);
or U247 (N_247,In_2753,In_2976);
nand U248 (N_248,In_2759,In_2886);
nor U249 (N_249,In_1182,In_884);
xor U250 (N_250,In_793,In_2921);
nand U251 (N_251,In_1498,In_2550);
xor U252 (N_252,In_2461,In_2274);
xnor U253 (N_253,In_47,In_1675);
or U254 (N_254,In_2702,In_2409);
and U255 (N_255,In_1001,In_979);
nor U256 (N_256,In_60,In_1818);
and U257 (N_257,In_2645,In_1974);
xnor U258 (N_258,In_323,In_2267);
and U259 (N_259,In_2879,In_1078);
nand U260 (N_260,In_2785,In_2304);
or U261 (N_261,In_636,In_1402);
nand U262 (N_262,In_2923,In_1804);
and U263 (N_263,In_2154,In_593);
nor U264 (N_264,In_2010,In_2801);
or U265 (N_265,In_523,In_1297);
nor U266 (N_266,In_1165,In_2478);
nand U267 (N_267,In_2528,In_2989);
xor U268 (N_268,In_766,In_1490);
nand U269 (N_269,In_1768,In_1227);
or U270 (N_270,In_1998,In_1169);
xnor U271 (N_271,In_541,In_2963);
nor U272 (N_272,In_1225,In_2083);
and U273 (N_273,In_184,In_626);
and U274 (N_274,In_2770,In_1248);
and U275 (N_275,In_921,In_101);
nor U276 (N_276,In_532,In_1918);
nor U277 (N_277,In_2427,In_848);
and U278 (N_278,In_1691,In_764);
xor U279 (N_279,In_1563,In_1865);
xnor U280 (N_280,In_670,In_1995);
xnor U281 (N_281,In_1574,In_2107);
or U282 (N_282,In_825,In_409);
nor U283 (N_283,In_2856,In_651);
xor U284 (N_284,In_2244,In_322);
and U285 (N_285,In_2065,In_2922);
and U286 (N_286,In_1765,In_282);
and U287 (N_287,In_1948,In_2210);
or U288 (N_288,In_1934,In_1471);
or U289 (N_289,In_2329,In_790);
nor U290 (N_290,In_471,In_1637);
xor U291 (N_291,In_2230,In_2220);
nor U292 (N_292,In_485,In_147);
xor U293 (N_293,In_1906,In_2740);
nor U294 (N_294,In_1005,In_1843);
nand U295 (N_295,In_2011,In_1977);
xor U296 (N_296,In_2162,In_1324);
and U297 (N_297,In_2465,In_1831);
and U298 (N_298,In_2261,In_54);
or U299 (N_299,In_337,In_667);
and U300 (N_300,In_1040,In_1750);
nor U301 (N_301,In_1973,In_1784);
xnor U302 (N_302,In_48,In_1152);
nand U303 (N_303,In_2767,In_963);
nor U304 (N_304,In_2820,In_2099);
and U305 (N_305,In_1951,In_2992);
xnor U306 (N_306,In_2273,In_202);
or U307 (N_307,In_1064,In_1081);
nand U308 (N_308,In_1075,In_255);
nand U309 (N_309,In_800,In_353);
nand U310 (N_310,In_1344,In_2791);
or U311 (N_311,In_2835,In_1518);
nand U312 (N_312,In_993,In_227);
xor U313 (N_313,In_1540,In_547);
and U314 (N_314,In_2917,In_1031);
xnor U315 (N_315,In_602,In_2576);
nor U316 (N_316,In_1823,In_1827);
or U317 (N_317,In_1970,In_1442);
nor U318 (N_318,In_2337,In_730);
nor U319 (N_319,In_2452,In_663);
nand U320 (N_320,In_2112,In_2260);
nor U321 (N_321,In_405,In_1021);
nand U322 (N_322,In_1003,In_2290);
nor U323 (N_323,In_1199,In_1156);
nor U324 (N_324,In_1328,In_280);
nor U325 (N_325,In_2297,In_374);
and U326 (N_326,In_837,In_45);
and U327 (N_327,In_1186,In_2388);
or U328 (N_328,In_806,In_310);
or U329 (N_329,In_606,In_1071);
nand U330 (N_330,In_2788,In_2129);
nand U331 (N_331,In_591,In_2713);
nor U332 (N_332,In_2892,In_2417);
or U333 (N_333,In_726,In_1258);
or U334 (N_334,In_784,In_2546);
or U335 (N_335,In_1890,In_586);
xor U336 (N_336,In_2305,In_2630);
nor U337 (N_337,In_1546,In_2691);
nand U338 (N_338,In_1488,In_997);
or U339 (N_339,In_95,In_472);
and U340 (N_340,In_2428,In_630);
nand U341 (N_341,In_2891,In_512);
nor U342 (N_342,In_1990,In_1124);
and U343 (N_343,In_673,In_889);
xor U344 (N_344,In_740,In_1100);
xor U345 (N_345,In_786,In_2715);
or U346 (N_346,In_2489,In_2187);
or U347 (N_347,In_1560,In_1202);
nand U348 (N_348,In_1698,In_2458);
and U349 (N_349,In_1365,In_771);
nand U350 (N_350,In_1016,In_1723);
xor U351 (N_351,In_2920,In_975);
or U352 (N_352,In_2070,In_245);
or U353 (N_353,In_1700,In_2857);
nand U354 (N_354,In_1250,In_1194);
nor U355 (N_355,In_912,In_2466);
xnor U356 (N_356,In_2265,In_1819);
or U357 (N_357,In_477,In_535);
nand U358 (N_358,In_1337,In_2616);
or U359 (N_359,In_543,In_1999);
nor U360 (N_360,In_1249,In_1764);
xnor U361 (N_361,In_1975,In_1867);
xor U362 (N_362,In_295,In_18);
nor U363 (N_363,In_2600,In_2198);
nand U364 (N_364,In_1054,In_2553);
nor U365 (N_365,In_2093,In_762);
and U366 (N_366,In_2284,In_334);
or U367 (N_367,In_1751,In_1826);
or U368 (N_368,In_590,In_1984);
or U369 (N_369,In_248,In_1210);
xor U370 (N_370,In_2454,In_1662);
or U371 (N_371,In_1134,In_428);
or U372 (N_372,In_241,In_1310);
xor U373 (N_373,In_653,In_75);
xnor U374 (N_374,In_916,In_2972);
nor U375 (N_375,In_1318,In_327);
nor U376 (N_376,In_2578,In_534);
or U377 (N_377,In_2650,In_1129);
nor U378 (N_378,In_2393,In_2524);
xor U379 (N_379,In_1038,In_1508);
nand U380 (N_380,In_971,In_2743);
or U381 (N_381,In_2475,In_1067);
xor U382 (N_382,In_2677,In_1851);
xnor U383 (N_383,In_747,In_2237);
nor U384 (N_384,In_1161,In_2539);
nand U385 (N_385,In_708,In_632);
nor U386 (N_386,In_2350,In_913);
nand U387 (N_387,In_454,In_2619);
nand U388 (N_388,In_2860,In_338);
xor U389 (N_389,In_12,In_841);
nand U390 (N_390,In_1600,In_2710);
or U391 (N_391,In_2993,In_1830);
or U392 (N_392,In_1744,In_170);
nor U393 (N_393,In_2847,In_1163);
or U394 (N_394,In_1678,In_961);
and U395 (N_395,In_1505,In_2157);
nand U396 (N_396,In_2185,In_2009);
nand U397 (N_397,In_171,In_367);
nor U398 (N_398,In_2580,In_1418);
xnor U399 (N_399,In_1093,In_451);
or U400 (N_400,In_1341,In_473);
nand U401 (N_401,In_2681,In_1096);
or U402 (N_402,In_1526,In_597);
nand U403 (N_403,In_516,In_758);
and U404 (N_404,In_1420,In_565);
and U405 (N_405,In_2957,In_328);
nor U406 (N_406,In_1828,In_967);
nand U407 (N_407,In_391,In_2148);
and U408 (N_408,In_1917,In_2051);
and U409 (N_409,In_2655,In_668);
or U410 (N_410,In_2937,In_1665);
or U411 (N_411,In_696,In_316);
nand U412 (N_412,In_1469,In_2614);
nand U413 (N_413,In_285,In_885);
or U414 (N_414,In_1683,In_2194);
or U415 (N_415,In_2153,In_264);
nor U416 (N_416,In_330,In_144);
xor U417 (N_417,In_2554,In_2867);
and U418 (N_418,In_1262,In_2047);
and U419 (N_419,In_1136,In_2479);
xnor U420 (N_420,In_826,In_1208);
xnor U421 (N_421,In_1801,In_299);
nand U422 (N_422,In_840,In_2109);
xor U423 (N_423,In_1309,In_1919);
nand U424 (N_424,In_2854,In_445);
or U425 (N_425,In_2299,In_254);
or U426 (N_426,In_1870,In_2776);
nor U427 (N_427,In_2889,In_718);
xnor U428 (N_428,In_1586,In_1618);
or U429 (N_429,In_453,In_2218);
or U430 (N_430,In_407,In_305);
and U431 (N_431,In_2022,In_1295);
or U432 (N_432,In_911,In_77);
nand U433 (N_433,In_1927,In_2916);
nor U434 (N_434,In_2410,In_844);
nand U435 (N_435,In_1314,In_691);
xnor U436 (N_436,In_974,In_2195);
or U437 (N_437,In_2943,In_705);
nand U438 (N_438,In_936,In_1554);
xor U439 (N_439,In_2931,In_1390);
nor U440 (N_440,In_157,In_545);
xnor U441 (N_441,In_313,In_459);
nor U442 (N_442,In_1640,In_2207);
and U443 (N_443,In_549,In_320);
and U444 (N_444,In_1104,In_2732);
nand U445 (N_445,In_744,In_994);
or U446 (N_446,In_2384,In_365);
xor U447 (N_447,In_493,In_2180);
or U448 (N_448,In_1461,In_403);
or U449 (N_449,In_2354,In_2666);
and U450 (N_450,In_2629,In_1467);
xnor U451 (N_451,In_402,In_2201);
and U452 (N_452,In_1535,In_2968);
or U453 (N_453,In_1858,In_615);
nor U454 (N_454,In_988,In_1614);
or U455 (N_455,In_2024,In_658);
or U456 (N_456,In_2927,In_2138);
nor U457 (N_457,In_959,In_1897);
nand U458 (N_458,In_2983,In_2778);
nor U459 (N_459,In_2568,In_2604);
or U460 (N_460,In_518,In_2596);
xor U461 (N_461,In_2733,In_2673);
and U462 (N_462,In_2448,In_2587);
xor U463 (N_463,In_13,In_645);
nand U464 (N_464,In_1624,In_1479);
nor U465 (N_465,In_1386,In_2188);
xor U466 (N_466,In_2034,In_289);
nor U467 (N_467,In_931,In_411);
xnor U468 (N_468,In_1084,In_1118);
or U469 (N_469,In_188,In_263);
or U470 (N_470,In_977,In_1421);
and U471 (N_471,In_82,In_2626);
and U472 (N_472,In_738,In_432);
nor U473 (N_473,In_1577,In_2303);
nand U474 (N_474,In_2240,In_2839);
and U475 (N_475,In_582,In_2599);
and U476 (N_476,In_2903,In_1125);
and U477 (N_477,In_922,In_266);
nand U478 (N_478,In_1141,In_2737);
nor U479 (N_479,In_968,In_440);
and U480 (N_480,In_1126,In_497);
nor U481 (N_481,In_1833,In_1771);
xnor U482 (N_482,In_937,In_1747);
xor U483 (N_483,In_2386,In_579);
xnor U484 (N_484,In_125,In_1176);
nor U485 (N_485,In_2092,In_1909);
nand U486 (N_486,In_2555,In_124);
and U487 (N_487,In_176,In_1745);
and U488 (N_488,In_2110,In_488);
nor U489 (N_489,In_1521,In_2144);
xor U490 (N_490,In_53,In_1473);
nor U491 (N_491,In_1841,In_2085);
nand U492 (N_492,In_989,In_1280);
nand U493 (N_493,In_2482,In_200);
xnor U494 (N_494,In_237,In_594);
and U495 (N_495,In_0,In_116);
or U496 (N_496,In_1769,In_166);
xor U497 (N_497,In_2558,In_2421);
or U498 (N_498,In_475,In_110);
and U499 (N_499,In_616,In_621);
nor U500 (N_500,In_823,In_148);
nor U501 (N_501,In_2717,In_2000);
and U502 (N_502,In_86,In_1415);
or U503 (N_503,In_2738,In_433);
and U504 (N_504,In_2007,In_225);
nand U505 (N_505,In_1785,In_957);
nor U506 (N_506,In_1416,In_2756);
nand U507 (N_507,In_1525,In_1572);
or U508 (N_508,In_2649,In_1503);
nand U509 (N_509,In_179,In_2538);
or U510 (N_510,In_420,In_2777);
xor U511 (N_511,In_1338,In_1410);
xor U512 (N_512,In_1696,In_2757);
or U513 (N_513,In_1873,In_2394);
xnor U514 (N_514,In_2822,In_1251);
nor U515 (N_515,In_1290,In_1881);
xor U516 (N_516,In_1140,In_1329);
nor U517 (N_517,In_1025,In_2216);
xnor U518 (N_518,In_2761,In_2078);
xor U519 (N_519,In_1433,In_347);
or U520 (N_520,In_1903,In_17);
or U521 (N_521,In_2974,In_2734);
or U522 (N_522,In_63,In_1846);
and U523 (N_523,In_1688,In_941);
nor U524 (N_524,In_390,In_1076);
and U525 (N_525,In_2327,In_1938);
nor U526 (N_526,In_796,In_293);
nand U527 (N_527,In_930,In_1200);
xnor U528 (N_528,In_2171,In_2102);
and U529 (N_529,In_1437,In_550);
nor U530 (N_530,In_1681,In_2585);
xnor U531 (N_531,In_1449,In_983);
or U532 (N_532,In_878,In_2894);
or U533 (N_533,In_2690,In_2859);
nand U534 (N_534,In_1274,In_1060);
nand U535 (N_535,In_219,In_2977);
or U536 (N_536,In_1850,In_962);
nand U537 (N_537,In_1693,In_1802);
and U538 (N_538,In_924,In_1253);
and U539 (N_539,In_628,In_1339);
nand U540 (N_540,In_386,In_746);
and U541 (N_541,In_1550,In_2088);
and U542 (N_542,In_483,In_1598);
and U543 (N_543,In_2995,In_567);
or U544 (N_544,In_1370,In_1777);
nand U545 (N_545,In_1154,In_753);
nand U546 (N_546,In_2291,In_1298);
or U547 (N_547,In_2652,In_1783);
xor U548 (N_548,In_2443,In_783);
or U549 (N_549,In_2663,In_2094);
nor U550 (N_550,In_1931,In_308);
xnor U551 (N_551,In_1184,In_2202);
xnor U552 (N_552,In_1530,In_1901);
or U553 (N_553,In_2781,In_1822);
nor U554 (N_554,In_1912,In_2097);
xor U555 (N_555,In_1077,In_128);
xor U556 (N_556,In_681,In_2914);
and U557 (N_557,In_1122,In_2956);
and U558 (N_558,In_539,In_1217);
and U559 (N_559,In_2392,In_2813);
xnor U560 (N_560,In_947,In_2053);
and U561 (N_561,In_2817,In_1111);
xnor U562 (N_562,In_2909,In_1057);
nor U563 (N_563,In_2298,In_2570);
or U564 (N_564,In_1177,In_1088);
and U565 (N_565,In_2398,In_2056);
nand U566 (N_566,In_380,In_2045);
and U567 (N_567,In_1465,In_2864);
or U568 (N_568,In_757,In_1011);
xor U569 (N_569,In_1438,In_1218);
and U570 (N_570,In_1407,In_1132);
and U571 (N_571,In_2368,In_244);
xnor U572 (N_572,In_2908,In_2292);
nand U573 (N_573,In_111,In_2038);
nand U574 (N_574,In_438,In_2257);
or U575 (N_575,In_2659,In_1742);
and U576 (N_576,In_2707,In_1940);
or U577 (N_577,In_2405,In_1429);
xor U578 (N_578,In_688,In_1463);
nor U579 (N_579,In_2435,In_1179);
and U580 (N_580,In_940,In_1811);
nor U581 (N_581,In_2958,In_1149);
and U582 (N_582,In_1715,In_1781);
xnor U583 (N_583,In_2170,In_2824);
xor U584 (N_584,In_729,In_2271);
nand U585 (N_585,In_2633,In_2918);
xor U586 (N_586,In_1597,In_2792);
nor U587 (N_587,In_1474,In_2798);
nand U588 (N_588,In_1778,In_1667);
xnor U589 (N_589,In_1188,In_311);
nor U590 (N_590,In_1119,In_286);
nor U591 (N_591,In_406,In_588);
nor U592 (N_592,In_2197,In_2975);
xnor U593 (N_593,In_1480,In_1944);
nand U594 (N_594,In_871,In_1892);
or U595 (N_595,In_1875,In_1267);
nor U596 (N_596,In_2212,In_1266);
or U597 (N_597,In_2574,In_2363);
nor U598 (N_598,In_537,In_1305);
and U599 (N_599,In_798,In_1454);
nor U600 (N_600,In_982,In_2158);
or U601 (N_601,In_2789,In_1757);
or U602 (N_602,In_162,In_2815);
nor U603 (N_603,In_2459,In_1335);
xor U604 (N_604,In_2991,In_1286);
or U605 (N_605,In_425,In_1237);
xnor U606 (N_606,In_2882,In_1558);
or U607 (N_607,In_1604,In_443);
or U608 (N_608,In_1902,In_2819);
nand U609 (N_609,In_398,In_1929);
nor U610 (N_610,In_1475,In_1430);
nand U611 (N_611,In_2377,In_2247);
nand U612 (N_612,In_1772,In_1599);
or U613 (N_613,In_2684,In_1896);
and U614 (N_614,In_2463,In_635);
xor U615 (N_615,In_2869,In_2229);
and U616 (N_616,In_2353,In_2748);
and U617 (N_617,In_858,In_1049);
nand U618 (N_618,In_160,In_1981);
xor U619 (N_619,In_1345,In_502);
nand U620 (N_620,In_1725,In_1391);
or U621 (N_621,In_2953,In_1000);
nor U622 (N_622,In_478,In_2275);
and U623 (N_623,In_2486,In_1886);
or U624 (N_624,In_637,In_1050);
nand U625 (N_625,In_1620,In_985);
nand U626 (N_626,In_2311,In_2654);
xnor U627 (N_627,In_1709,In_1516);
or U628 (N_628,In_31,In_949);
nand U629 (N_629,In_174,In_883);
and U630 (N_630,In_902,In_442);
xor U631 (N_631,In_230,In_526);
and U632 (N_632,In_1956,In_2852);
nand U633 (N_633,In_525,In_1412);
nand U634 (N_634,In_1891,In_1008);
nor U635 (N_635,In_2206,In_873);
or U636 (N_636,In_1294,In_1746);
and U637 (N_637,In_2611,In_589);
and U638 (N_638,In_221,In_16);
or U639 (N_639,In_1795,In_1594);
nand U640 (N_640,In_2954,In_1704);
nand U641 (N_641,In_2940,In_89);
nand U642 (N_642,In_900,In_2127);
and U643 (N_643,In_2880,In_2324);
xor U644 (N_644,In_707,In_1874);
xor U645 (N_645,In_2543,In_1610);
nor U646 (N_646,In_548,In_2227);
nand U647 (N_647,In_37,In_1066);
nand U648 (N_648,In_984,In_278);
and U649 (N_649,In_1601,In_2730);
and U650 (N_650,In_142,In_1355);
xnor U651 (N_651,In_2997,In_304);
or U652 (N_652,In_1839,In_1937);
and U653 (N_653,In_1528,In_1115);
or U654 (N_654,In_2372,In_2125);
and U655 (N_655,In_96,In_1736);
nand U656 (N_656,In_828,In_1734);
and U657 (N_657,In_2301,In_659);
or U658 (N_658,In_1020,In_2470);
and U659 (N_659,In_2870,In_2317);
and U660 (N_660,In_2027,In_2025);
xor U661 (N_661,In_1882,In_270);
nand U662 (N_662,In_2875,In_1452);
nor U663 (N_663,In_2982,In_2924);
nand U664 (N_664,In_1333,In_2401);
or U665 (N_665,In_1446,In_2973);
nand U666 (N_666,In_1123,In_1061);
nor U667 (N_667,In_2912,In_1470);
or U668 (N_668,In_1231,In_1056);
nor U669 (N_669,In_560,In_269);
nand U670 (N_670,In_660,In_1590);
xnor U671 (N_671,In_854,In_1425);
xnor U672 (N_672,In_890,In_1388);
nor U673 (N_673,In_1014,In_109);
xor U674 (N_674,In_2725,In_1171);
and U675 (N_675,In_2680,In_2147);
and U676 (N_676,In_1300,In_2828);
or U677 (N_677,In_2095,In_2084);
nand U678 (N_678,In_791,In_2904);
nor U679 (N_679,In_1012,In_716);
nor U680 (N_680,In_42,In_55);
xnor U681 (N_681,In_2522,In_2783);
nand U682 (N_682,In_8,In_417);
nor U683 (N_683,In_2926,In_1303);
nand U684 (N_684,In_2161,In_556);
xnor U685 (N_685,In_577,In_1296);
nand U686 (N_686,In_257,In_2374);
or U687 (N_687,In_2196,In_777);
or U688 (N_688,In_2899,In_2536);
nor U689 (N_689,In_25,In_2402);
nand U690 (N_690,In_1201,In_2245);
and U691 (N_691,In_2565,In_1423);
nor U692 (N_692,In_676,In_2890);
or U693 (N_693,In_164,In_1302);
nand U694 (N_694,In_2572,In_2132);
and U695 (N_695,In_2391,In_114);
xor U696 (N_696,In_972,In_2446);
xnor U697 (N_697,In_2215,In_748);
and U698 (N_698,In_1573,In_1871);
and U699 (N_699,In_2262,In_1806);
and U700 (N_700,In_2772,In_2316);
and U701 (N_701,In_1711,In_2874);
xnor U702 (N_702,In_1971,In_2727);
xnor U703 (N_703,In_1,In_426);
and U704 (N_704,In_2119,In_1108);
or U705 (N_705,In_1497,In_1466);
or U706 (N_706,In_1868,In_1234);
xnor U707 (N_707,In_392,In_599);
xor U708 (N_708,In_2637,In_2925);
and U709 (N_709,In_1537,In_2693);
or U710 (N_710,In_794,In_326);
nor U711 (N_711,In_1489,In_2457);
xnor U712 (N_712,In_511,In_2662);
nand U713 (N_713,In_2160,In_2672);
nand U714 (N_714,In_1740,In_2573);
and U715 (N_715,In_2082,In_1556);
xnor U716 (N_716,In_743,In_1834);
and U717 (N_717,In_2204,In_1254);
nand U718 (N_718,In_1847,In_575);
or U719 (N_719,In_2547,In_2222);
nor U720 (N_720,In_359,In_1026);
nor U721 (N_721,In_2111,In_769);
nor U722 (N_722,In_1994,In_1243);
nand U723 (N_723,In_499,In_2823);
and U724 (N_724,In_613,In_189);
nand U725 (N_725,In_2371,In_2683);
nor U726 (N_726,In_1192,In_115);
and U727 (N_727,In_2594,In_932);
nand U728 (N_728,In_2434,In_2800);
and U729 (N_729,In_19,In_1997);
xnor U730 (N_730,In_1657,In_2877);
xnor U731 (N_731,In_2534,In_928);
xnor U732 (N_732,In_1213,In_935);
and U733 (N_733,In_760,In_2087);
or U734 (N_734,In_2603,In_1825);
and U735 (N_735,In_1987,In_2067);
xor U736 (N_736,In_2674,In_208);
xnor U737 (N_737,In_899,In_745);
or U738 (N_738,In_2701,In_2848);
nand U739 (N_739,In_2323,In_68);
or U740 (N_740,In_815,In_752);
nor U741 (N_741,In_281,In_104);
xor U742 (N_742,In_2794,In_1373);
xor U743 (N_743,In_2887,In_533);
or U744 (N_744,In_1923,In_684);
and U745 (N_745,In_2667,In_368);
or U746 (N_746,In_2499,In_2131);
nand U747 (N_747,In_2521,In_1053);
or U748 (N_748,In_956,In_2179);
xnor U749 (N_749,In_699,In_1579);
nor U750 (N_750,In_2049,In_1101);
nand U751 (N_751,In_943,In_2028);
nor U752 (N_752,In_595,In_2059);
and U753 (N_753,In_500,In_2407);
nand U754 (N_754,In_1018,In_1529);
nor U755 (N_755,In_2177,In_2895);
nor U756 (N_756,In_1095,In_2678);
nand U757 (N_757,In_1327,In_759);
and U758 (N_758,In_1612,In_450);
or U759 (N_759,In_152,In_1315);
and U760 (N_760,In_201,In_1085);
or U761 (N_761,In_379,In_447);
xor U762 (N_762,In_408,In_2113);
nor U763 (N_763,In_462,In_1580);
nor U764 (N_764,In_2338,In_43);
or U765 (N_765,In_2932,In_2622);
and U766 (N_766,In_495,In_999);
nor U767 (N_767,In_145,In_1576);
xor U768 (N_768,In_250,In_2483);
xor U769 (N_769,In_1712,In_2079);
nand U770 (N_770,In_623,In_1708);
nand U771 (N_771,In_2834,In_249);
nand U772 (N_772,In_1926,In_1603);
nand U773 (N_773,In_801,In_1639);
xnor U774 (N_774,In_1958,In_686);
and U775 (N_775,In_856,In_2708);
nand U776 (N_776,In_811,In_1247);
xnor U777 (N_777,In_1002,In_446);
or U778 (N_778,In_2074,In_857);
and U779 (N_779,In_2326,In_2726);
and U780 (N_780,In_197,In_1173);
or U781 (N_781,In_1619,In_2978);
and U782 (N_782,In_2871,In_141);
nor U783 (N_783,In_1342,In_1074);
xnor U784 (N_784,In_375,In_2062);
and U785 (N_785,In_788,In_933);
nor U786 (N_786,In_1261,In_226);
nand U787 (N_787,In_1028,In_1147);
xor U788 (N_788,In_1880,In_1190);
xor U789 (N_789,In_239,In_1138);
xnor U790 (N_790,In_1533,In_1232);
nand U791 (N_791,In_2598,In_2530);
nor U792 (N_792,In_1268,In_1626);
nor U793 (N_793,In_1148,In_897);
or U794 (N_794,In_692,In_400);
and U795 (N_795,In_2450,In_584);
xnor U796 (N_796,In_2933,In_2124);
nor U797 (N_797,In_333,In_2915);
and U798 (N_798,In_1083,In_1652);
and U799 (N_799,In_1183,In_291);
nor U800 (N_800,In_2309,In_2949);
nor U801 (N_801,In_2804,In_2319);
nand U802 (N_802,In_1114,In_2540);
xnor U803 (N_803,In_72,In_559);
nand U804 (N_804,In_1350,In_876);
and U805 (N_805,In_1571,In_914);
nor U806 (N_806,In_1810,In_1651);
or U807 (N_807,In_2249,In_1223);
and U808 (N_808,In_1493,In_1353);
nand U809 (N_809,In_2531,In_1367);
nor U810 (N_810,In_732,In_1131);
nand U811 (N_811,In_33,In_1701);
nor U812 (N_812,In_627,In_2352);
xor U813 (N_813,In_2242,In_761);
xnor U814 (N_814,In_207,In_1719);
or U815 (N_815,In_2026,In_352);
nand U816 (N_816,In_2699,In_2621);
and U817 (N_817,In_690,In_2339);
nand U818 (N_818,In_1888,In_1677);
nand U819 (N_819,In_1144,In_741);
or U820 (N_820,In_1349,In_2505);
nand U821 (N_821,In_2503,In_436);
and U822 (N_822,In_301,In_1354);
and U823 (N_823,In_945,In_1376);
nor U824 (N_824,In_127,In_2064);
xor U825 (N_825,In_2039,In_2825);
or U826 (N_826,In_773,In_1898);
xnor U827 (N_827,In_1893,In_2561);
xor U828 (N_828,In_2741,In_2251);
xor U829 (N_829,In_1259,In_2361);
nor U830 (N_830,In_2669,In_874);
nand U831 (N_831,In_1401,In_2928);
nor U832 (N_832,In_2081,In_360);
nand U833 (N_833,In_669,In_382);
nand U834 (N_834,In_1396,In_2590);
or U835 (N_835,In_343,In_839);
nor U836 (N_836,In_701,In_412);
nor U837 (N_837,In_2334,In_81);
xnor U838 (N_838,In_728,In_855);
xnor U839 (N_839,In_2472,In_389);
xor U840 (N_840,In_274,In_803);
nand U841 (N_841,In_2469,In_1976);
and U842 (N_842,In_1794,In_120);
and U843 (N_843,In_2641,In_888);
nor U844 (N_844,In_2254,In_2518);
nand U845 (N_845,In_920,In_1311);
nand U846 (N_846,In_816,In_2582);
or U847 (N_847,In_619,In_2238);
and U848 (N_848,In_1643,In_2340);
nor U849 (N_849,In_1448,In_1840);
and U850 (N_850,In_211,In_2168);
xor U851 (N_851,In_2872,In_1589);
and U852 (N_852,In_2108,In_1939);
nor U853 (N_853,In_26,In_1813);
and U854 (N_854,In_639,In_907);
or U855 (N_855,In_2250,In_314);
and U856 (N_856,In_832,In_1377);
or U857 (N_857,In_1679,In_1379);
nor U858 (N_858,In_2843,In_307);
or U859 (N_859,In_2769,In_2176);
and U860 (N_860,In_675,In_215);
or U861 (N_861,In_981,In_2001);
nand U862 (N_862,In_2294,In_505);
and U863 (N_863,In_2766,In_2774);
xor U864 (N_864,In_1635,In_703);
or U865 (N_865,In_2938,In_419);
or U866 (N_866,In_242,In_881);
nand U867 (N_867,In_2898,In_1669);
or U868 (N_868,In_1648,In_113);
xor U869 (N_869,In_2225,In_763);
xnor U870 (N_870,In_1389,In_1445);
nand U871 (N_871,In_6,In_998);
nor U872 (N_872,In_566,In_102);
nor U873 (N_873,In_1633,In_2476);
nor U874 (N_874,In_363,In_563);
xor U875 (N_875,In_461,In_486);
xnor U876 (N_876,In_1062,In_2057);
or U877 (N_877,In_1094,In_1838);
xor U878 (N_878,In_2135,In_1608);
nand U879 (N_879,In_2355,In_1786);
and U880 (N_880,In_1548,In_1275);
or U881 (N_881,In_1180,In_1816);
xnor U882 (N_882,In_7,In_2279);
and U883 (N_883,In_2181,In_2306);
or U884 (N_884,In_2462,In_915);
xnor U885 (N_885,In_2679,In_1628);
nor U886 (N_886,In_1228,In_2101);
and U887 (N_887,In_340,In_770);
or U888 (N_888,In_995,In_2128);
and U889 (N_889,In_355,In_1945);
xnor U890 (N_890,In_2467,In_2623);
xnor U891 (N_891,In_990,In_1128);
or U892 (N_892,In_2744,In_2426);
nand U893 (N_893,In_2037,In_1366);
nand U894 (N_894,In_1146,In_650);
xor U895 (N_895,In_2373,In_2507);
nand U896 (N_896,In_362,In_1842);
xnor U897 (N_897,In_1814,In_1866);
xor U898 (N_898,In_2865,In_1022);
xor U899 (N_899,In_2404,In_206);
xor U900 (N_900,In_1728,In_1063);
xor U901 (N_901,In_1236,In_387);
xnor U902 (N_902,In_1292,In_273);
nor U903 (N_903,In_685,In_622);
nor U904 (N_904,In_1506,In_797);
xor U905 (N_905,In_2456,In_862);
or U906 (N_906,In_2685,In_1514);
and U907 (N_907,In_2712,In_2268);
nor U908 (N_908,In_2605,In_2213);
nand U909 (N_909,In_1178,In_1343);
and U910 (N_910,In_1968,In_94);
and U911 (N_911,In_950,In_2485);
xnor U912 (N_912,In_1375,In_904);
and U913 (N_913,In_2802,In_2190);
nand U914 (N_914,In_2779,In_2624);
xnor U915 (N_915,In_1174,In_558);
nand U916 (N_916,In_1646,In_2086);
xor U917 (N_917,In_712,In_1686);
and U918 (N_918,In_356,In_813);
nor U919 (N_919,In_2420,In_1660);
or U920 (N_920,In_2018,In_2747);
xor U921 (N_921,In_2224,In_2549);
and U922 (N_922,In_847,In_455);
nor U923 (N_923,In_1288,In_2935);
nor U924 (N_924,In_1245,In_544);
and U925 (N_925,In_1672,In_767);
xor U926 (N_926,In_546,In_1583);
nor U927 (N_927,In_2881,In_819);
xor U928 (N_928,In_810,In_966);
xnor U929 (N_929,In_2019,In_315);
nand U930 (N_930,In_67,In_1485);
or U931 (N_931,In_647,In_809);
and U932 (N_932,In_277,In_1004);
nor U933 (N_933,In_2315,In_1575);
or U934 (N_934,In_2496,In_1523);
nand U935 (N_935,In_2515,In_1426);
or U936 (N_936,In_2739,In_2658);
xnor U937 (N_937,In_865,In_183);
and U938 (N_938,In_905,In_1928);
nand U939 (N_939,In_1211,In_2172);
nor U940 (N_940,In_2841,In_2052);
nor U941 (N_941,In_2211,In_303);
or U942 (N_942,In_246,In_2682);
nor U943 (N_943,In_2866,In_342);
or U944 (N_944,In_464,In_2169);
or U945 (N_945,In_578,In_2235);
nor U946 (N_946,In_2758,In_1037);
xor U947 (N_947,In_267,In_2849);
nor U948 (N_948,In_1972,In_2893);
xor U949 (N_949,In_1517,In_287);
xnor U950 (N_950,In_2661,In_1059);
nor U951 (N_951,In_2617,In_1848);
and U952 (N_952,In_1547,In_1755);
or U953 (N_953,In_2960,In_2203);
nand U954 (N_954,In_2422,In_1036);
xnor U955 (N_955,In_231,In_1399);
nand U956 (N_956,In_934,In_1697);
and U957 (N_957,In_603,In_2347);
and U958 (N_958,In_223,In_1444);
nor U959 (N_959,In_1562,In_1726);
xor U960 (N_960,In_838,In_69);
nor U961 (N_961,In_1876,In_896);
xor U962 (N_962,In_1748,In_1230);
xnor U963 (N_963,In_2853,In_76);
nand U964 (N_964,In_1638,In_895);
nor U965 (N_965,In_2058,In_700);
nand U966 (N_966,In_2066,In_2634);
xnor U967 (N_967,In_354,In_50);
nand U968 (N_968,In_460,In_1706);
nor U969 (N_969,In_510,In_2577);
nor U970 (N_970,In_2990,In_1889);
or U971 (N_971,In_2408,In_2643);
or U972 (N_972,In_1361,In_2517);
nor U973 (N_973,In_2277,In_413);
nand U974 (N_974,In_198,In_422);
xnor U975 (N_975,In_1317,In_1264);
nand U976 (N_976,In_1419,In_79);
xor U977 (N_977,In_1051,In_754);
or U978 (N_978,In_1441,In_2106);
or U979 (N_979,In_2098,In_551);
and U980 (N_980,In_2787,In_868);
nand U981 (N_981,In_252,In_2276);
nor U982 (N_982,In_332,In_1293);
xnor U983 (N_983,In_1949,In_2321);
nor U984 (N_984,In_1824,In_778);
or U985 (N_985,In_711,In_1006);
and U986 (N_986,In_1160,In_9);
xnor U987 (N_987,In_1641,In_774);
and U988 (N_988,In_1510,In_1240);
xnor U989 (N_989,In_2272,In_2900);
xor U990 (N_990,In_554,In_228);
xnor U991 (N_991,In_318,In_265);
and U992 (N_992,In_2731,In_799);
nor U993 (N_993,In_2980,In_268);
and U994 (N_994,In_2330,In_2356);
nor U995 (N_995,In_1207,In_1106);
nor U996 (N_996,In_1372,In_2998);
nand U997 (N_997,In_680,In_2883);
or U998 (N_998,In_2579,In_98);
or U999 (N_999,In_1685,In_2638);
nor U1000 (N_1000,In_2036,In_2149);
or U1001 (N_1001,In_1159,In_1024);
nand U1002 (N_1002,In_2390,In_2100);
nor U1003 (N_1003,In_62,In_1570);
and U1004 (N_1004,In_1495,In_2762);
or U1005 (N_1005,In_2544,In_2331);
xnor U1006 (N_1006,In_925,In_704);
or U1007 (N_1007,In_2939,In_1952);
xnor U1008 (N_1008,In_1117,In_1332);
nand U1009 (N_1009,In_2602,In_1427);
nand U1010 (N_1010,In_1766,In_2285);
and U1011 (N_1011,In_1561,In_2994);
and U1012 (N_1012,In_143,In_1907);
nor U1013 (N_1013,In_1961,In_2833);
and U1014 (N_1014,In_2259,In_2610);
or U1015 (N_1015,In_2907,In_694);
or U1016 (N_1016,In_74,In_2008);
nor U1017 (N_1017,In_2236,In_2375);
nor U1018 (N_1018,In_1642,In_2941);
xor U1019 (N_1019,In_1674,In_2697);
nor U1020 (N_1020,In_126,In_2631);
xor U1021 (N_1021,In_2567,In_204);
and U1022 (N_1022,In_1162,In_1239);
and U1023 (N_1023,In_366,In_1464);
nand U1024 (N_1024,In_1431,In_1960);
nor U1025 (N_1025,In_1689,In_2286);
and U1026 (N_1026,In_1428,In_2810);
or U1027 (N_1027,In_2711,In_232);
and U1028 (N_1028,In_2786,In_2136);
nor U1029 (N_1029,In_1157,In_1967);
xnor U1030 (N_1030,In_1499,In_498);
xnor U1031 (N_1031,In_2657,In_2320);
nand U1032 (N_1032,In_119,In_610);
nand U1033 (N_1033,In_2033,In_381);
nor U1034 (N_1034,In_927,In_2913);
or U1035 (N_1035,In_1707,In_1483);
nand U1036 (N_1036,In_2812,In_2307);
and U1037 (N_1037,In_2803,In_2625);
nor U1038 (N_1038,In_520,In_1815);
nand U1039 (N_1039,In_1395,In_469);
or U1040 (N_1040,In_59,In_1405);
xnor U1041 (N_1041,In_946,In_341);
nand U1042 (N_1042,In_640,In_2232);
and U1043 (N_1043,In_1797,In_1435);
or U1044 (N_1044,In_1710,In_306);
nor U1045 (N_1045,In_1043,In_191);
nor U1046 (N_1046,In_151,In_468);
or U1047 (N_1047,In_2192,In_180);
nor U1048 (N_1048,In_2312,In_1602);
nand U1049 (N_1049,In_492,In_2423);
xor U1050 (N_1050,In_2345,In_1716);
xnor U1051 (N_1051,In_2359,In_731);
xnor U1052 (N_1052,In_1494,In_399);
xnor U1053 (N_1053,In_833,In_992);
nand U1054 (N_1054,In_2460,In_457);
xnor U1055 (N_1055,In_1284,In_2615);
and U1056 (N_1056,In_1844,In_1282);
or U1057 (N_1057,In_103,In_1364);
nor U1058 (N_1058,In_1143,In_1507);
nand U1059 (N_1059,In_404,In_1047);
or U1060 (N_1060,In_1256,In_1812);
nor U1061 (N_1061,In_1915,In_1392);
and U1062 (N_1062,In_388,In_618);
nand U1063 (N_1063,In_260,In_1894);
nand U1064 (N_1064,In_122,In_2775);
nor U1065 (N_1065,In_1041,In_491);
and U1066 (N_1066,In_99,In_1932);
nor U1067 (N_1067,In_117,In_592);
nand U1068 (N_1068,In_309,In_918);
and U1069 (N_1069,In_92,In_1319);
and U1070 (N_1070,In_5,In_41);
xor U1071 (N_1071,In_11,In_2424);
and U1072 (N_1072,In_2491,In_1205);
and U1073 (N_1073,In_2601,In_1279);
nand U1074 (N_1074,In_1703,In_1233);
and U1075 (N_1075,In_1478,In_2378);
nand U1076 (N_1076,In_2930,In_2163);
and U1077 (N_1077,In_137,In_2396);
and U1078 (N_1078,In_1219,In_2780);
xor U1079 (N_1079,In_1203,In_2140);
xnor U1080 (N_1080,In_2016,In_2964);
and U1081 (N_1081,In_1007,In_509);
xor U1082 (N_1082,In_346,In_2706);
nor U1083 (N_1083,In_199,In_1763);
and U1084 (N_1084,In_97,In_1042);
or U1085 (N_1085,In_633,In_683);
xnor U1086 (N_1086,In_724,In_608);
nor U1087 (N_1087,In_948,In_617);
and U1088 (N_1088,In_721,In_1033);
nand U1089 (N_1089,In_253,In_217);
nor U1090 (N_1090,In_1541,In_555);
and U1091 (N_1091,In_1996,In_2231);
nand U1092 (N_1092,In_1242,In_2228);
nor U1093 (N_1093,In_1983,In_2552);
and U1094 (N_1094,In_1800,In_1175);
or U1095 (N_1095,In_564,In_2314);
nor U1096 (N_1096,In_2670,In_2333);
xnor U1097 (N_1097,In_2984,In_2050);
or U1098 (N_1098,In_378,In_344);
or U1099 (N_1099,In_863,In_2842);
nor U1100 (N_1100,In_1082,In_1511);
nor U1101 (N_1101,In_2696,In_1500);
nand U1102 (N_1102,In_2252,In_1137);
nor U1103 (N_1103,In_1509,In_275);
xnor U1104 (N_1104,In_804,In_1539);
and U1105 (N_1105,In_118,In_1650);
nand U1106 (N_1106,In_1578,In_2280);
and U1107 (N_1107,In_965,In_1484);
or U1108 (N_1108,In_2433,In_1167);
xnor U1109 (N_1109,In_654,In_614);
nor U1110 (N_1110,In_2043,In_1837);
nor U1111 (N_1111,In_1098,In_1684);
and U1112 (N_1112,In_2527,In_452);
nor U1113 (N_1113,In_2282,In_133);
and U1114 (N_1114,In_358,In_439);
and U1115 (N_1115,In_1455,In_792);
nor U1116 (N_1116,In_1793,In_1761);
nand U1117 (N_1117,In_261,In_489);
nand U1118 (N_1118,In_2511,In_580);
xnor U1119 (N_1119,In_2344,In_1089);
and U1120 (N_1120,In_163,In_1862);
xnor U1121 (N_1121,In_2139,In_1277);
nand U1122 (N_1122,In_2342,In_30);
and U1123 (N_1123,In_571,In_1910);
xor U1124 (N_1124,In_2494,In_2283);
or U1125 (N_1125,In_631,In_710);
nor U1126 (N_1126,In_1699,In_2440);
nand U1127 (N_1127,In_1055,In_1775);
or U1128 (N_1128,In_2425,In_782);
nand U1129 (N_1129,In_1979,In_1629);
xnor U1130 (N_1130,In_1930,In_2826);
xor U1131 (N_1131,In_903,In_2484);
and U1132 (N_1132,In_892,In_713);
and U1133 (N_1133,In_449,In_2749);
or U1134 (N_1134,In_2571,In_1105);
and U1135 (N_1135,In_576,In_1753);
and U1136 (N_1136,In_2071,In_40);
and U1137 (N_1137,In_2134,In_695);
nor U1138 (N_1138,In_2133,In_298);
or U1139 (N_1139,In_1468,In_1663);
nor U1140 (N_1140,In_1854,In_185);
xnor U1141 (N_1141,In_2754,In_2178);
or U1142 (N_1142,In_1121,In_1271);
nor U1143 (N_1143,In_1456,In_1291);
and U1144 (N_1144,In_1954,In_427);
xnor U1145 (N_1145,In_1397,In_2901);
nor U1146 (N_1146,In_1754,In_1659);
or U1147 (N_1147,In_569,In_2105);
xor U1148 (N_1148,In_2335,In_190);
nor U1149 (N_1149,In_2589,In_1720);
nor U1150 (N_1150,In_336,In_1611);
xor U1151 (N_1151,In_1462,In_2591);
xor U1152 (N_1152,In_384,In_2752);
nand U1153 (N_1153,In_1914,In_139);
nand U1154 (N_1154,In_2750,In_2243);
or U1155 (N_1155,In_908,In_466);
nor U1156 (N_1156,In_1729,In_2208);
nand U1157 (N_1157,In_507,In_2431);
and U1158 (N_1158,In_581,In_2453);
nor U1159 (N_1159,In_1935,In_2017);
and U1160 (N_1160,In_1351,In_1432);
and U1161 (N_1161,In_2318,In_2896);
xor U1162 (N_1162,In_2919,In_138);
xor U1163 (N_1163,In_1592,In_2006);
or U1164 (N_1164,In_1368,In_2313);
nor U1165 (N_1165,In_181,In_2246);
and U1166 (N_1166,In_717,In_2595);
or U1167 (N_1167,In_233,In_944);
xor U1168 (N_1168,In_501,In_370);
nor U1169 (N_1169,In_1185,In_2380);
or U1170 (N_1170,In_1899,In_866);
nor U1171 (N_1171,In_2471,In_1803);
or U1172 (N_1172,In_612,In_1166);
or U1173 (N_1173,In_939,In_1630);
nor U1174 (N_1174,In_2073,In_860);
or U1175 (N_1175,In_297,In_2542);
xor U1176 (N_1176,In_214,In_1661);
xnor U1177 (N_1177,In_1682,In_536);
nand U1178 (N_1178,In_1555,In_2556);
or U1179 (N_1179,In_679,In_736);
and U1180 (N_1180,In_1322,In_574);
or U1181 (N_1181,In_1287,In_345);
xor U1182 (N_1182,In_187,In_1492);
nor U1183 (N_1183,In_1065,In_2293);
nand U1184 (N_1184,In_891,In_2366);
nor U1185 (N_1185,In_1316,In_1904);
or U1186 (N_1186,In_1596,In_1451);
xor U1187 (N_1187,In_1695,In_2832);
or U1188 (N_1188,In_882,In_236);
nor U1189 (N_1189,In_1557,In_2054);
nor U1190 (N_1190,In_689,In_2174);
nand U1191 (N_1191,In_1805,In_2145);
and U1192 (N_1192,In_2042,In_733);
nor U1193 (N_1193,In_2688,In_2514);
xor U1194 (N_1194,In_434,In_822);
xor U1195 (N_1195,In_836,In_1276);
or U1196 (N_1196,In_2061,In_173);
xor U1197 (N_1197,In_2325,In_1357);
or U1198 (N_1198,In_2040,In_2444);
xor U1199 (N_1199,In_78,In_1714);
or U1200 (N_1200,In_2934,In_709);
nor U1201 (N_1201,In_887,In_1821);
nand U1202 (N_1202,In_1265,In_2117);
nor U1203 (N_1203,In_22,In_2784);
nor U1204 (N_1204,In_755,In_827);
and U1205 (N_1205,In_1656,In_2676);
or U1206 (N_1206,In_648,In_2628);
or U1207 (N_1207,In_35,In_2745);
xor U1208 (N_1208,In_953,In_1450);
and U1209 (N_1209,In_1724,In_1849);
xor U1210 (N_1210,In_843,In_2902);
or U1211 (N_1211,In_480,In_1911);
and U1212 (N_1212,In_2412,In_2876);
and U1213 (N_1213,In_1953,In_2481);
nor U1214 (N_1214,In_28,In_383);
xor U1215 (N_1215,In_2429,In_1269);
and U1216 (N_1216,In_1836,In_2031);
nor U1217 (N_1217,In_2322,In_1713);
nor U1218 (N_1218,In_1631,In_1422);
nor U1219 (N_1219,In_1380,In_1632);
nand U1220 (N_1220,In_1153,In_2818);
or U1221 (N_1221,In_1531,In_2414);
or U1222 (N_1222,In_2060,In_2709);
nor U1223 (N_1223,In_2646,In_756);
xor U1224 (N_1224,In_2729,In_952);
nor U1225 (N_1225,In_880,In_2248);
xnor U1226 (N_1226,In_1206,In_243);
and U1227 (N_1227,In_1925,In_2606);
nand U1228 (N_1228,In_1069,In_222);
nand U1229 (N_1229,In_1722,In_938);
nor U1230 (N_1230,In_2217,In_1273);
or U1231 (N_1231,In_429,In_2827);
and U1232 (N_1232,In_393,In_2126);
nand U1233 (N_1233,In_2971,In_220);
or U1234 (N_1234,In_2831,In_1549);
or U1235 (N_1235,In_697,In_1198);
nand U1236 (N_1236,In_2506,In_256);
xnor U1237 (N_1237,In_1980,In_1195);
nor U1238 (N_1238,In_2358,In_2122);
and U1239 (N_1239,In_2945,In_1170);
nor U1240 (N_1240,In_2668,In_1235);
and U1241 (N_1241,In_524,In_1481);
xor U1242 (N_1242,In_2782,In_1417);
xor U1243 (N_1243,In_2845,In_1965);
nor U1244 (N_1244,In_312,In_84);
and U1245 (N_1245,In_842,In_1673);
nor U1246 (N_1246,In_1052,In_1409);
nand U1247 (N_1247,In_2966,In_814);
nor U1248 (N_1248,In_2508,In_1776);
xor U1249 (N_1249,In_849,In_1378);
or U1250 (N_1250,In_1788,In_1900);
nor U1251 (N_1251,In_2905,In_2529);
nor U1252 (N_1252,In_121,In_802);
and U1253 (N_1253,In_973,In_1356);
xor U1254 (N_1254,In_2013,In_1150);
and U1255 (N_1255,In_2836,In_251);
nand U1256 (N_1256,In_154,In_1913);
xor U1257 (N_1257,In_2946,In_2055);
nor U1258 (N_1258,In_986,In_2773);
or U1259 (N_1259,In_2988,In_2072);
and U1260 (N_1260,In_2151,In_2175);
nor U1261 (N_1261,In_2120,In_271);
and U1262 (N_1262,In_561,In_503);
nor U1263 (N_1263,In_2296,In_1680);
and U1264 (N_1264,In_2911,In_482);
nor U1265 (N_1265,In_2255,In_2955);
and U1266 (N_1266,In_818,In_1306);
xor U1267 (N_1267,In_107,In_57);
nor U1268 (N_1268,In_1443,In_1616);
or U1269 (N_1269,In_657,In_212);
and U1270 (N_1270,In_1520,In_517);
nand U1271 (N_1271,In_29,In_1229);
xnor U1272 (N_1272,In_2501,In_2728);
nor U1273 (N_1273,In_875,In_186);
and U1274 (N_1274,In_2969,In_61);
nor U1275 (N_1275,In_1737,In_1099);
nand U1276 (N_1276,In_1346,In_2665);
or U1277 (N_1277,In_2593,In_629);
xnor U1278 (N_1278,In_1519,In_213);
and U1279 (N_1279,In_978,In_1460);
xor U1280 (N_1280,In_2664,In_2032);
xnor U1281 (N_1281,In_456,In_1933);
nor U1282 (N_1282,In_100,In_2389);
nand U1283 (N_1283,In_85,In_27);
xnor U1284 (N_1284,In_2449,In_620);
nand U1285 (N_1285,In_1158,In_611);
xnor U1286 (N_1286,In_2069,In_2287);
nand U1287 (N_1287,In_294,In_674);
or U1288 (N_1288,In_2588,In_2020);
or U1289 (N_1289,In_1384,In_562);
nor U1290 (N_1290,In_830,In_134);
or U1291 (N_1291,In_1950,In_1988);
nand U1292 (N_1292,In_2551,In_609);
xor U1293 (N_1293,In_106,In_2642);
nand U1294 (N_1294,In_2165,In_372);
or U1295 (N_1295,In_474,In_2768);
and U1296 (N_1296,In_529,In_1738);
nor U1297 (N_1297,In_530,In_1857);
nor U1298 (N_1298,In_2509,In_2432);
or U1299 (N_1299,In_1424,In_870);
or U1300 (N_1300,In_2403,In_585);
xnor U1301 (N_1301,In_845,In_1942);
nor U1302 (N_1302,In_2226,In_1527);
nor U1303 (N_1303,In_1664,In_235);
xnor U1304 (N_1304,In_1155,In_70);
nand U1305 (N_1305,In_656,In_2793);
and U1306 (N_1306,In_1670,In_317);
or U1307 (N_1307,In_1622,In_2612);
or U1308 (N_1308,In_329,In_2967);
nor U1309 (N_1309,In_2942,In_2266);
or U1310 (N_1310,In_909,In_394);
nor U1311 (N_1311,In_431,In_494);
nand U1312 (N_1312,In_2182,In_1636);
xor U1313 (N_1313,In_2948,In_2695);
xnor U1314 (N_1314,In_2406,In_2520);
or U1315 (N_1315,In_1542,In_23);
nand U1316 (N_1316,In_2269,In_2751);
and U1317 (N_1317,In_1326,In_1212);
xor U1318 (N_1318,In_216,In_976);
nor U1319 (N_1319,In_385,In_2821);
and U1320 (N_1320,In_2861,In_821);
nand U1321 (N_1321,In_1214,In_1718);
nor U1322 (N_1322,In_2906,In_1538);
xor U1323 (N_1323,In_1197,In_209);
or U1324 (N_1324,In_51,In_1845);
and U1325 (N_1325,In_430,In_1584);
nand U1326 (N_1326,In_1634,In_527);
nand U1327 (N_1327,In_1623,In_969);
and U1328 (N_1328,In_2015,In_2806);
or U1329 (N_1329,In_2,In_1922);
nor U1330 (N_1330,In_1861,In_666);
xnor U1331 (N_1331,In_38,In_175);
nor U1332 (N_1332,In_2640,In_737);
nand U1333 (N_1333,In_772,In_2855);
xnor U1334 (N_1334,In_542,In_259);
and U1335 (N_1335,In_224,In_2103);
nor U1336 (N_1336,In_169,In_2644);
or U1337 (N_1337,In_105,In_722);
nand U1338 (N_1338,In_1439,In_1959);
xor U1339 (N_1339,In_1534,In_2143);
nand U1340 (N_1340,In_14,In_2104);
or U1341 (N_1341,In_2575,In_479);
nand U1342 (N_1342,In_1671,In_587);
and U1343 (N_1343,In_1692,In_642);
nand U1344 (N_1344,In_2395,In_1791);
and U1345 (N_1345,In_15,In_325);
nand U1346 (N_1346,In_2495,In_1885);
and U1347 (N_1347,In_2510,In_2234);
or U1348 (N_1348,In_1869,In_2005);
nor U1349 (N_1349,In_671,In_10);
nand U1350 (N_1350,In_1654,In_2500);
and U1351 (N_1351,In_1130,In_2155);
nand U1352 (N_1352,In_130,In_570);
nand U1353 (N_1353,In_1393,In_324);
and U1354 (N_1354,In_463,In_2790);
or U1355 (N_1355,In_919,In_421);
nor U1356 (N_1356,In_1172,In_1070);
xnor U1357 (N_1357,In_2348,In_1374);
xor U1358 (N_1358,In_1702,In_1582);
nand U1359 (N_1359,In_1676,In_665);
and U1360 (N_1360,In_1587,In_519);
nor U1361 (N_1361,In_2379,In_158);
or U1362 (N_1362,In_1015,In_853);
nand U1363 (N_1363,In_1969,In_1260);
and U1364 (N_1364,In_2862,In_1782);
xor U1365 (N_1365,In_195,In_901);
xor U1366 (N_1366,In_1941,In_4);
nand U1367 (N_1367,In_1009,In_2981);
or U1368 (N_1368,In_661,In_1658);
and U1369 (N_1369,In_1829,In_1993);
nand U1370 (N_1370,In_1859,In_1835);
xor U1371 (N_1371,In_2490,In_1585);
xor U1372 (N_1372,In_2996,In_2430);
xor U1373 (N_1373,In_1387,In_401);
nand U1374 (N_1374,In_234,In_923);
and U1375 (N_1375,In_768,In_2660);
nor U1376 (N_1376,In_2851,In_834);
nand U1377 (N_1377,In_1312,In_2850);
nand U1378 (N_1378,In_2399,In_1887);
or U1379 (N_1379,In_1270,In_1962);
nor U1380 (N_1380,In_155,In_1606);
and U1381 (N_1381,In_687,In_1644);
or U1382 (N_1382,In_1808,In_444);
xnor U1383 (N_1383,In_2618,In_2302);
or U1384 (N_1384,In_1964,In_2636);
xnor U1385 (N_1385,In_2400,In_1408);
nor U1386 (N_1386,In_776,In_1358);
nand U1387 (N_1387,In_52,In_2493);
xnor U1388 (N_1388,In_218,In_1362);
and U1389 (N_1389,In_872,In_2214);
nand U1390 (N_1390,In_835,In_484);
or U1391 (N_1391,In_2021,In_2704);
xor U1392 (N_1392,In_572,In_1301);
xor U1393 (N_1393,In_2962,In_1617);
nor U1394 (N_1394,In_1325,In_2387);
nand U1395 (N_1395,In_2878,In_600);
and U1396 (N_1396,In_1705,In_290);
and U1397 (N_1397,In_1308,In_2123);
and U1398 (N_1398,In_2146,In_1476);
nand U1399 (N_1399,In_2438,In_2692);
or U1400 (N_1400,In_1220,In_2357);
nor U1401 (N_1401,In_1645,In_1278);
nand U1402 (N_1402,In_1216,In_2076);
and U1403 (N_1403,In_2608,In_1982);
and U1404 (N_1404,In_2797,In_2164);
or U1405 (N_1405,In_2209,In_1946);
nand U1406 (N_1406,In_1457,In_1653);
or U1407 (N_1407,In_1743,In_2910);
nor U1408 (N_1408,In_2349,In_182);
xor U1409 (N_1409,In_2765,In_2343);
or U1410 (N_1410,In_508,In_2360);
nor U1411 (N_1411,In_1113,In_2586);
nor U1412 (N_1412,In_49,In_1666);
nor U1413 (N_1413,In_1086,In_2156);
nand U1414 (N_1414,In_2116,In_1878);
nand U1415 (N_1415,In_2114,In_1515);
and U1416 (N_1416,In_2516,In_1330);
and U1417 (N_1417,In_2592,In_1035);
nor U1418 (N_1418,In_247,In_2885);
nand U1419 (N_1419,In_1863,In_1916);
nor U1420 (N_1420,In_2191,In_1985);
and U1421 (N_1421,In_1588,In_1109);
or U1422 (N_1422,In_583,In_2341);
xor U1423 (N_1423,In_377,In_894);
and U1424 (N_1424,In_2346,In_2533);
and U1425 (N_1425,In_373,In_2584);
and U1426 (N_1426,In_1110,In_605);
nand U1427 (N_1427,In_693,In_1187);
or U1428 (N_1428,In_2724,In_864);
xor U1429 (N_1429,In_910,In_1544);
nor U1430 (N_1430,In_1883,In_2581);
nand U1431 (N_1431,In_1774,In_448);
and U1432 (N_1432,In_1030,In_415);
nor U1433 (N_1433,In_1196,In_1853);
or U1434 (N_1434,In_1908,In_1536);
and U1435 (N_1435,In_1224,In_2445);
xor U1436 (N_1436,In_1760,In_1359);
or U1437 (N_1437,In_2278,In_1605);
nor U1438 (N_1438,In_1360,In_1472);
nand U1439 (N_1439,In_652,In_1079);
xnor U1440 (N_1440,In_36,In_2947);
nor U1441 (N_1441,In_514,In_2183);
or U1442 (N_1442,In_2118,In_34);
xnor U1443 (N_1443,In_795,In_2233);
and U1444 (N_1444,In_2868,In_1809);
and U1445 (N_1445,In_73,In_2451);
xor U1446 (N_1446,In_807,In_2046);
nor U1447 (N_1447,In_942,In_846);
or U1448 (N_1448,In_2159,In_279);
nand U1449 (N_1449,In_2030,In_339);
xor U1450 (N_1450,In_2385,In_1145);
nand U1451 (N_1451,In_2562,In_1770);
and U1452 (N_1452,In_2002,In_2837);
nand U1453 (N_1453,In_2846,In_1193);
and U1454 (N_1454,In_568,In_2799);
and U1455 (N_1455,In_960,In_2441);
and U1456 (N_1456,In_2635,In_123);
or U1457 (N_1457,In_88,In_719);
xnor U1458 (N_1458,In_1073,In_538);
xnor U1459 (N_1459,In_437,In_2221);
nor U1460 (N_1460,In_1221,In_487);
and U1461 (N_1461,In_1164,In_1832);
or U1462 (N_1462,In_2526,In_2411);
nand U1463 (N_1463,In_808,In_1263);
nor U1464 (N_1464,In_2689,In_2970);
and U1465 (N_1465,In_150,In_1733);
nand U1466 (N_1466,In_1727,In_2735);
xnor U1467 (N_1467,In_2497,In_2705);
xor U1468 (N_1468,In_1447,In_1807);
xor U1469 (N_1469,In_1381,In_1019);
nand U1470 (N_1470,In_331,In_751);
nor U1471 (N_1471,In_644,In_852);
xor U1472 (N_1472,In_2447,In_2077);
nand U1473 (N_1473,In_1403,In_2746);
or U1474 (N_1474,In_522,In_2419);
nor U1475 (N_1475,In_66,In_1453);
or U1476 (N_1476,In_1752,In_2141);
or U1477 (N_1477,In_601,In_1513);
nand U1478 (N_1478,In_573,In_44);
and U1479 (N_1479,In_1413,In_664);
xnor U1480 (N_1480,In_153,In_178);
nor U1481 (N_1481,In_2130,In_2381);
or U1482 (N_1482,In_917,In_210);
or U1483 (N_1483,In_2239,In_2760);
xor U1484 (N_1484,In_2639,In_465);
or U1485 (N_1485,In_2647,In_2004);
nor U1486 (N_1486,In_2498,In_1487);
nand U1487 (N_1487,In_1655,In_1856);
or U1488 (N_1488,In_2714,In_1504);
nor U1489 (N_1489,In_1027,In_192);
and U1490 (N_1490,In_1989,In_1759);
or U1491 (N_1491,In_682,In_93);
xor U1492 (N_1492,In_2205,In_2675);
or U1493 (N_1493,In_1877,In_1564);
nand U1494 (N_1494,In_71,In_2569);
or U1495 (N_1495,In_46,In_1730);
and U1496 (N_1496,In_1283,In_805);
or U1497 (N_1497,In_2369,In_1091);
nor U1498 (N_1498,In_2722,In_2442);
nor U1499 (N_1499,In_490,In_725);
nor U1500 (N_1500,N_183,N_511);
nand U1501 (N_1501,N_367,N_508);
xor U1502 (N_1502,N_485,N_223);
and U1503 (N_1503,N_1263,N_233);
xnor U1504 (N_1504,N_703,N_495);
xor U1505 (N_1505,N_738,N_1451);
and U1506 (N_1506,N_1269,N_527);
nand U1507 (N_1507,N_1435,N_1192);
nand U1508 (N_1508,N_373,N_726);
xor U1509 (N_1509,N_486,N_901);
xor U1510 (N_1510,N_1027,N_1406);
and U1511 (N_1511,N_547,N_53);
and U1512 (N_1512,N_1215,N_1409);
nor U1513 (N_1513,N_739,N_883);
nor U1514 (N_1514,N_431,N_942);
nor U1515 (N_1515,N_1219,N_470);
xnor U1516 (N_1516,N_1172,N_1092);
nand U1517 (N_1517,N_410,N_1495);
or U1518 (N_1518,N_647,N_1209);
xnor U1519 (N_1519,N_1227,N_1397);
xnor U1520 (N_1520,N_1132,N_175);
nand U1521 (N_1521,N_323,N_1370);
xnor U1522 (N_1522,N_1041,N_697);
nand U1523 (N_1523,N_787,N_1031);
nand U1524 (N_1524,N_819,N_960);
nand U1525 (N_1525,N_1111,N_272);
nor U1526 (N_1526,N_565,N_1106);
nand U1527 (N_1527,N_1144,N_891);
xnor U1528 (N_1528,N_657,N_610);
nand U1529 (N_1529,N_328,N_658);
nor U1530 (N_1530,N_59,N_928);
nor U1531 (N_1531,N_1290,N_354);
and U1532 (N_1532,N_1175,N_1422);
and U1533 (N_1533,N_690,N_832);
xnor U1534 (N_1534,N_1196,N_1496);
nor U1535 (N_1535,N_673,N_445);
nand U1536 (N_1536,N_1375,N_1321);
and U1537 (N_1537,N_775,N_839);
or U1538 (N_1538,N_366,N_8);
nand U1539 (N_1539,N_1083,N_1373);
and U1540 (N_1540,N_39,N_818);
and U1541 (N_1541,N_81,N_1418);
and U1542 (N_1542,N_1080,N_758);
or U1543 (N_1543,N_321,N_423);
xnor U1544 (N_1544,N_737,N_468);
and U1545 (N_1545,N_299,N_668);
or U1546 (N_1546,N_1363,N_885);
or U1547 (N_1547,N_1024,N_1183);
or U1548 (N_1548,N_1143,N_221);
and U1549 (N_1549,N_72,N_219);
or U1550 (N_1550,N_642,N_718);
nand U1551 (N_1551,N_362,N_415);
xnor U1552 (N_1552,N_904,N_1484);
and U1553 (N_1553,N_44,N_636);
or U1554 (N_1554,N_1464,N_1009);
nand U1555 (N_1555,N_207,N_191);
nand U1556 (N_1556,N_988,N_1051);
nand U1557 (N_1557,N_80,N_779);
nand U1558 (N_1558,N_654,N_553);
xnor U1559 (N_1559,N_246,N_424);
nor U1560 (N_1560,N_56,N_561);
nor U1561 (N_1561,N_194,N_898);
xnor U1562 (N_1562,N_377,N_734);
nand U1563 (N_1563,N_1214,N_753);
and U1564 (N_1564,N_811,N_580);
or U1565 (N_1565,N_286,N_780);
nor U1566 (N_1566,N_778,N_551);
or U1567 (N_1567,N_736,N_593);
xor U1568 (N_1568,N_1071,N_253);
nor U1569 (N_1569,N_1493,N_1008);
and U1570 (N_1570,N_555,N_683);
nand U1571 (N_1571,N_949,N_651);
and U1572 (N_1572,N_187,N_1304);
xnor U1573 (N_1573,N_1120,N_215);
nand U1574 (N_1574,N_135,N_628);
and U1575 (N_1575,N_550,N_777);
or U1576 (N_1576,N_948,N_999);
nor U1577 (N_1577,N_101,N_240);
nor U1578 (N_1578,N_976,N_613);
nor U1579 (N_1579,N_788,N_66);
nand U1580 (N_1580,N_863,N_688);
or U1581 (N_1581,N_270,N_1360);
nand U1582 (N_1582,N_1037,N_1243);
and U1583 (N_1583,N_318,N_766);
or U1584 (N_1584,N_1331,N_413);
xnor U1585 (N_1585,N_230,N_1249);
or U1586 (N_1586,N_1320,N_51);
and U1587 (N_1587,N_1049,N_465);
xor U1588 (N_1588,N_1486,N_1429);
and U1589 (N_1589,N_119,N_212);
and U1590 (N_1590,N_1157,N_98);
nor U1591 (N_1591,N_1184,N_902);
nor U1592 (N_1592,N_521,N_977);
xnor U1593 (N_1593,N_57,N_991);
xor U1594 (N_1594,N_265,N_608);
nand U1595 (N_1595,N_162,N_1152);
nand U1596 (N_1596,N_24,N_1354);
xnor U1597 (N_1597,N_786,N_97);
and U1598 (N_1598,N_528,N_829);
nor U1599 (N_1599,N_498,N_124);
xnor U1600 (N_1600,N_469,N_582);
nand U1601 (N_1601,N_1283,N_419);
nand U1602 (N_1602,N_1217,N_810);
and U1603 (N_1603,N_42,N_1436);
xnor U1604 (N_1604,N_634,N_1458);
or U1605 (N_1605,N_251,N_138);
nor U1606 (N_1606,N_368,N_952);
xnor U1607 (N_1607,N_311,N_1294);
nor U1608 (N_1608,N_517,N_1424);
nor U1609 (N_1609,N_992,N_1467);
nor U1610 (N_1610,N_1362,N_395);
and U1611 (N_1611,N_916,N_155);
or U1612 (N_1612,N_696,N_980);
xor U1613 (N_1613,N_963,N_1232);
xor U1614 (N_1614,N_292,N_306);
nand U1615 (N_1615,N_1153,N_1292);
nor U1616 (N_1616,N_386,N_978);
or U1617 (N_1617,N_447,N_1186);
and U1618 (N_1618,N_1161,N_914);
nand U1619 (N_1619,N_1056,N_574);
xnor U1620 (N_1620,N_947,N_332);
nor U1621 (N_1621,N_721,N_600);
xnor U1622 (N_1622,N_982,N_1385);
or U1623 (N_1623,N_1337,N_615);
and U1624 (N_1624,N_1229,N_861);
nand U1625 (N_1625,N_454,N_152);
nand U1626 (N_1626,N_1468,N_132);
nand U1627 (N_1627,N_78,N_1223);
and U1628 (N_1628,N_241,N_560);
or U1629 (N_1629,N_62,N_1343);
and U1630 (N_1630,N_1123,N_526);
or U1631 (N_1631,N_765,N_938);
xor U1632 (N_1632,N_1187,N_964);
nor U1633 (N_1633,N_64,N_704);
nand U1634 (N_1634,N_794,N_1282);
xnor U1635 (N_1635,N_283,N_562);
nor U1636 (N_1636,N_370,N_702);
or U1637 (N_1637,N_438,N_348);
nand U1638 (N_1638,N_1444,N_1043);
and U1639 (N_1639,N_1014,N_452);
or U1640 (N_1640,N_248,N_63);
or U1641 (N_1641,N_588,N_372);
nand U1642 (N_1642,N_1439,N_1115);
nand U1643 (N_1643,N_443,N_1159);
or U1644 (N_1644,N_958,N_147);
or U1645 (N_1645,N_1154,N_163);
nor U1646 (N_1646,N_403,N_1449);
and U1647 (N_1647,N_676,N_1303);
nand U1648 (N_1648,N_672,N_1440);
or U1649 (N_1649,N_385,N_873);
nor U1650 (N_1650,N_71,N_1118);
xor U1651 (N_1651,N_394,N_327);
nor U1652 (N_1652,N_22,N_484);
nand U1653 (N_1653,N_536,N_817);
xnor U1654 (N_1654,N_473,N_381);
nor U1655 (N_1655,N_520,N_1039);
xor U1656 (N_1656,N_455,N_1177);
and U1657 (N_1657,N_337,N_1279);
or U1658 (N_1658,N_356,N_1126);
and U1659 (N_1659,N_1270,N_353);
and U1660 (N_1660,N_854,N_481);
and U1661 (N_1661,N_1150,N_320);
nand U1662 (N_1662,N_317,N_396);
nand U1663 (N_1663,N_173,N_308);
xnor U1664 (N_1664,N_420,N_349);
or U1665 (N_1665,N_502,N_1368);
and U1666 (N_1666,N_745,N_1066);
nand U1667 (N_1667,N_1256,N_603);
or U1668 (N_1668,N_1365,N_558);
and U1669 (N_1669,N_1151,N_945);
or U1670 (N_1670,N_1046,N_1233);
xor U1671 (N_1671,N_1133,N_931);
or U1672 (N_1672,N_1237,N_759);
or U1673 (N_1673,N_875,N_1275);
nor U1674 (N_1674,N_789,N_235);
nand U1675 (N_1675,N_973,N_1193);
nor U1676 (N_1676,N_933,N_1179);
nand U1677 (N_1677,N_1463,N_1348);
or U1678 (N_1678,N_18,N_1421);
nand U1679 (N_1679,N_375,N_1178);
nand U1680 (N_1680,N_974,N_518);
and U1681 (N_1681,N_214,N_1280);
nand U1682 (N_1682,N_158,N_193);
and U1683 (N_1683,N_1206,N_369);
and U1684 (N_1684,N_257,N_939);
and U1685 (N_1685,N_886,N_1403);
nor U1686 (N_1686,N_453,N_442);
or U1687 (N_1687,N_247,N_434);
or U1688 (N_1688,N_679,N_1019);
or U1689 (N_1689,N_1202,N_165);
xor U1690 (N_1690,N_1061,N_355);
nand U1691 (N_1691,N_1399,N_1417);
or U1692 (N_1692,N_1076,N_869);
or U1693 (N_1693,N_1318,N_1366);
xor U1694 (N_1694,N_1253,N_416);
or U1695 (N_1695,N_1338,N_1313);
or U1696 (N_1696,N_6,N_1333);
nor U1697 (N_1697,N_514,N_316);
nor U1698 (N_1698,N_180,N_1125);
nand U1699 (N_1699,N_1021,N_995);
xnor U1700 (N_1700,N_260,N_113);
nor U1701 (N_1701,N_597,N_459);
or U1702 (N_1702,N_189,N_380);
nor U1703 (N_1703,N_1203,N_347);
and U1704 (N_1704,N_868,N_464);
or U1705 (N_1705,N_809,N_120);
or U1706 (N_1706,N_1479,N_218);
and U1707 (N_1707,N_1470,N_491);
xor U1708 (N_1708,N_500,N_531);
xnor U1709 (N_1709,N_14,N_92);
xnor U1710 (N_1710,N_289,N_534);
xor U1711 (N_1711,N_1136,N_4);
and U1712 (N_1712,N_767,N_448);
nand U1713 (N_1713,N_1453,N_252);
or U1714 (N_1714,N_576,N_796);
and U1715 (N_1715,N_709,N_569);
xnor U1716 (N_1716,N_1221,N_401);
nand U1717 (N_1717,N_1346,N_913);
nor U1718 (N_1718,N_649,N_856);
xor U1719 (N_1719,N_674,N_782);
or U1720 (N_1720,N_1460,N_1089);
xor U1721 (N_1721,N_213,N_1386);
and U1722 (N_1722,N_1314,N_1431);
or U1723 (N_1723,N_532,N_1259);
xor U1724 (N_1724,N_1176,N_621);
or U1725 (N_1725,N_1180,N_728);
or U1726 (N_1726,N_524,N_890);
xnor U1727 (N_1727,N_645,N_1430);
and U1728 (N_1728,N_409,N_346);
nor U1729 (N_1729,N_732,N_1419);
nor U1730 (N_1730,N_263,N_88);
nor U1731 (N_1731,N_123,N_427);
or U1732 (N_1732,N_1015,N_671);
nor U1733 (N_1733,N_1393,N_89);
xor U1734 (N_1734,N_1442,N_730);
and U1735 (N_1735,N_590,N_1077);
or U1736 (N_1736,N_40,N_1312);
nor U1737 (N_1737,N_461,N_754);
nor U1738 (N_1738,N_1218,N_107);
xnor U1739 (N_1739,N_1065,N_1257);
and U1740 (N_1740,N_710,N_584);
or U1741 (N_1741,N_178,N_694);
and U1742 (N_1742,N_271,N_538);
or U1743 (N_1743,N_1028,N_55);
and U1744 (N_1744,N_859,N_157);
nand U1745 (N_1745,N_930,N_1171);
and U1746 (N_1746,N_1389,N_1254);
nand U1747 (N_1747,N_1491,N_224);
or U1748 (N_1748,N_979,N_823);
and U1749 (N_1749,N_1480,N_1335);
nor U1750 (N_1750,N_29,N_393);
or U1751 (N_1751,N_993,N_865);
or U1752 (N_1752,N_382,N_1384);
nand U1753 (N_1753,N_35,N_879);
nor U1754 (N_1754,N_336,N_1247);
or U1755 (N_1755,N_1369,N_882);
nor U1756 (N_1756,N_1059,N_352);
and U1757 (N_1757,N_975,N_457);
nor U1758 (N_1758,N_609,N_851);
nand U1759 (N_1759,N_926,N_1322);
xor U1760 (N_1760,N_1459,N_125);
and U1761 (N_1761,N_262,N_677);
and U1762 (N_1762,N_1305,N_894);
and U1763 (N_1763,N_203,N_1473);
nand U1764 (N_1764,N_707,N_535);
nand U1765 (N_1765,N_855,N_79);
xor U1766 (N_1766,N_681,N_48);
or U1767 (N_1767,N_717,N_1446);
and U1768 (N_1768,N_340,N_1230);
or U1769 (N_1769,N_411,N_852);
xnor U1770 (N_1770,N_1287,N_121);
and U1771 (N_1771,N_392,N_548);
nand U1772 (N_1772,N_1396,N_1357);
and U1773 (N_1773,N_141,N_480);
nand U1774 (N_1774,N_813,N_429);
or U1775 (N_1775,N_236,N_282);
nand U1776 (N_1776,N_1383,N_1388);
nor U1777 (N_1777,N_705,N_763);
xor U1778 (N_1778,N_335,N_623);
xor U1779 (N_1779,N_781,N_1057);
nand U1780 (N_1780,N_446,N_1265);
and U1781 (N_1781,N_820,N_563);
nand U1782 (N_1782,N_573,N_860);
nand U1783 (N_1783,N_1053,N_1104);
and U1784 (N_1784,N_893,N_492);
or U1785 (N_1785,N_806,N_1211);
or U1786 (N_1786,N_1489,N_1286);
and U1787 (N_1787,N_1355,N_624);
nand U1788 (N_1788,N_1058,N_1);
nand U1789 (N_1789,N_25,N_720);
nand U1790 (N_1790,N_1340,N_334);
nor U1791 (N_1791,N_606,N_96);
and U1792 (N_1792,N_635,N_406);
or U1793 (N_1793,N_1235,N_1310);
or U1794 (N_1794,N_801,N_670);
nand U1795 (N_1795,N_12,N_379);
and U1796 (N_1796,N_644,N_871);
nand U1797 (N_1797,N_1328,N_274);
xnor U1798 (N_1798,N_250,N_1207);
xnor U1799 (N_1799,N_567,N_268);
nand U1800 (N_1800,N_1478,N_1345);
or U1801 (N_1801,N_1062,N_307);
and U1802 (N_1802,N_962,N_1007);
nand U1803 (N_1803,N_577,N_921);
xnor U1804 (N_1804,N_37,N_675);
or U1805 (N_1805,N_1213,N_1351);
and U1806 (N_1806,N_1163,N_772);
nand U1807 (N_1807,N_1438,N_444);
or U1808 (N_1808,N_36,N_1376);
or U1809 (N_1809,N_371,N_1117);
or U1810 (N_1810,N_46,N_1488);
nand U1811 (N_1811,N_1274,N_1352);
nor U1812 (N_1812,N_1086,N_0);
nand U1813 (N_1813,N_1364,N_877);
nand U1814 (N_1814,N_546,N_267);
nand U1815 (N_1815,N_1003,N_731);
nor U1816 (N_1816,N_225,N_60);
or U1817 (N_1817,N_1216,N_1324);
and U1818 (N_1818,N_329,N_166);
nand U1819 (N_1819,N_544,N_428);
xnor U1820 (N_1820,N_439,N_983);
or U1821 (N_1821,N_2,N_1073);
and U1822 (N_1822,N_769,N_1447);
xor U1823 (N_1823,N_460,N_872);
or U1824 (N_1824,N_5,N_1110);
and U1825 (N_1825,N_506,N_554);
xnor U1826 (N_1826,N_903,N_1006);
or U1827 (N_1827,N_640,N_83);
or U1828 (N_1828,N_757,N_325);
or U1829 (N_1829,N_106,N_1017);
or U1830 (N_1830,N_1450,N_50);
xnor U1831 (N_1831,N_404,N_1455);
xnor U1832 (N_1832,N_1428,N_493);
xnor U1833 (N_1833,N_803,N_475);
nand U1834 (N_1834,N_599,N_1099);
or U1835 (N_1835,N_1420,N_1081);
or U1836 (N_1836,N_598,N_515);
nor U1837 (N_1837,N_279,N_1063);
xor U1838 (N_1838,N_456,N_587);
nand U1839 (N_1839,N_1139,N_1330);
xnor U1840 (N_1840,N_751,N_1038);
xnor U1841 (N_1841,N_1413,N_1317);
nand U1842 (N_1842,N_1296,N_857);
or U1843 (N_1843,N_943,N_844);
nand U1844 (N_1844,N_525,N_111);
xnor U1845 (N_1845,N_907,N_579);
or U1846 (N_1846,N_174,N_682);
nand U1847 (N_1847,N_1128,N_1145);
and U1848 (N_1848,N_989,N_1045);
nand U1849 (N_1849,N_1372,N_510);
nand U1850 (N_1850,N_950,N_228);
nor U1851 (N_1851,N_586,N_1140);
nor U1852 (N_1852,N_302,N_1166);
nor U1853 (N_1853,N_816,N_896);
xor U1854 (N_1854,N_1020,N_650);
and U1855 (N_1855,N_216,N_1239);
and U1856 (N_1856,N_7,N_350);
nor U1857 (N_1857,N_1005,N_652);
nor U1858 (N_1858,N_1130,N_1261);
xor U1859 (N_1859,N_612,N_222);
or U1860 (N_1860,N_1390,N_1361);
and U1861 (N_1861,N_1064,N_516);
or U1862 (N_1862,N_591,N_1094);
xor U1863 (N_1863,N_105,N_1142);
or U1864 (N_1864,N_729,N_946);
or U1865 (N_1865,N_830,N_984);
xor U1866 (N_1866,N_227,N_1129);
and U1867 (N_1867,N_244,N_405);
nand U1868 (N_1868,N_1238,N_791);
and U1869 (N_1869,N_231,N_1252);
nand U1870 (N_1870,N_944,N_1212);
xor U1871 (N_1871,N_1173,N_981);
nor U1872 (N_1872,N_114,N_542);
xor U1873 (N_1873,N_1341,N_666);
or U1874 (N_1874,N_1068,N_773);
xor U1875 (N_1875,N_85,N_1079);
xnor U1876 (N_1876,N_680,N_229);
or U1877 (N_1877,N_1082,N_1339);
xor U1878 (N_1878,N_238,N_314);
and U1879 (N_1879,N_627,N_848);
and U1880 (N_1880,N_474,N_1298);
and U1881 (N_1881,N_1042,N_156);
or U1882 (N_1882,N_169,N_312);
and U1883 (N_1883,N_618,N_743);
nand U1884 (N_1884,N_632,N_1427);
nor U1885 (N_1885,N_287,N_1316);
nand U1886 (N_1886,N_450,N_815);
xor U1887 (N_1887,N_638,N_298);
or U1888 (N_1888,N_458,N_708);
and U1889 (N_1889,N_828,N_259);
nor U1890 (N_1890,N_559,N_77);
nor U1891 (N_1891,N_1168,N_47);
nand U1892 (N_1892,N_1072,N_874);
nand U1893 (N_1893,N_1359,N_82);
nor U1894 (N_1894,N_742,N_954);
nand U1895 (N_1895,N_522,N_571);
or U1896 (N_1896,N_835,N_1411);
nand U1897 (N_1897,N_834,N_17);
nand U1898 (N_1898,N_716,N_254);
nor U1899 (N_1899,N_825,N_1197);
and U1900 (N_1900,N_805,N_32);
and U1901 (N_1901,N_243,N_198);
nand U1902 (N_1902,N_210,N_842);
nor U1903 (N_1903,N_566,N_205);
and U1904 (N_1904,N_324,N_1010);
and U1905 (N_1905,N_1044,N_276);
or U1906 (N_1906,N_827,N_740);
nor U1907 (N_1907,N_714,N_698);
and U1908 (N_1908,N_1302,N_43);
nand U1909 (N_1909,N_1469,N_291);
or U1910 (N_1910,N_389,N_1169);
xor U1911 (N_1911,N_237,N_1022);
nand U1912 (N_1912,N_261,N_1069);
nor U1913 (N_1913,N_1210,N_539);
nand U1914 (N_1914,N_1398,N_333);
nand U1915 (N_1915,N_797,N_1378);
and U1916 (N_1916,N_1122,N_1085);
nand U1917 (N_1917,N_607,N_326);
xor U1918 (N_1918,N_1349,N_1162);
xor U1919 (N_1919,N_208,N_837);
or U1920 (N_1920,N_432,N_339);
and U1921 (N_1921,N_596,N_866);
nand U1922 (N_1922,N_653,N_19);
nor U1923 (N_1923,N_750,N_530);
xor U1924 (N_1924,N_139,N_16);
nor U1925 (N_1925,N_784,N_1474);
nand U1926 (N_1926,N_1060,N_126);
and U1927 (N_1927,N_552,N_422);
or U1928 (N_1928,N_987,N_1311);
and U1929 (N_1929,N_1107,N_853);
nor U1930 (N_1930,N_1148,N_887);
nor U1931 (N_1931,N_503,N_1164);
xor U1932 (N_1932,N_115,N_1358);
and U1933 (N_1933,N_204,N_614);
xor U1934 (N_1934,N_619,N_1258);
nor U1935 (N_1935,N_1100,N_13);
or U1936 (N_1936,N_1138,N_1033);
xor U1937 (N_1937,N_118,N_1097);
and U1938 (N_1938,N_545,N_391);
nand U1939 (N_1939,N_74,N_1475);
nor U1940 (N_1940,N_1412,N_1262);
xnor U1941 (N_1941,N_192,N_1228);
nor U1942 (N_1942,N_384,N_34);
nor U1943 (N_1943,N_1102,N_1105);
nor U1944 (N_1944,N_1147,N_112);
or U1945 (N_1945,N_1353,N_611);
nand U1946 (N_1946,N_1395,N_1408);
or U1947 (N_1947,N_418,N_641);
and U1948 (N_1948,N_1319,N_440);
nor U1949 (N_1949,N_1032,N_1181);
xnor U1950 (N_1950,N_840,N_70);
or U1951 (N_1951,N_585,N_906);
and U1952 (N_1952,N_275,N_924);
nand U1953 (N_1953,N_908,N_145);
or U1954 (N_1954,N_655,N_578);
xor U1955 (N_1955,N_153,N_604);
nand U1956 (N_1956,N_793,N_84);
and U1957 (N_1957,N_1476,N_1295);
xor U1958 (N_1958,N_996,N_1426);
xnor U1959 (N_1959,N_1267,N_541);
nand U1960 (N_1960,N_927,N_722);
or U1961 (N_1961,N_1090,N_665);
xor U1962 (N_1962,N_170,N_199);
nor U1963 (N_1963,N_1067,N_1371);
and U1964 (N_1964,N_303,N_581);
xnor U1965 (N_1965,N_300,N_998);
xnor U1966 (N_1966,N_1327,N_1158);
or U1967 (N_1967,N_188,N_1201);
or U1968 (N_1968,N_1289,N_833);
or U1969 (N_1969,N_31,N_637);
and U1970 (N_1970,N_463,N_537);
nor U1971 (N_1971,N_184,N_482);
xnor U1972 (N_1972,N_479,N_669);
xor U1973 (N_1973,N_488,N_951);
or U1974 (N_1974,N_363,N_1036);
nand U1975 (N_1975,N_836,N_1407);
xor U1976 (N_1976,N_790,N_1098);
nor U1977 (N_1977,N_102,N_109);
or U1978 (N_1978,N_1342,N_167);
nand U1979 (N_1979,N_255,N_1297);
xor U1980 (N_1980,N_295,N_804);
or U1981 (N_1981,N_1185,N_667);
xnor U1982 (N_1982,N_1461,N_912);
nand U1983 (N_1983,N_1160,N_864);
xor U1984 (N_1984,N_1276,N_509);
xnor U1985 (N_1985,N_845,N_313);
or U1986 (N_1986,N_747,N_990);
or U1987 (N_1987,N_646,N_626);
nand U1988 (N_1988,N_831,N_151);
or U1989 (N_1989,N_899,N_1101);
and U1990 (N_1990,N_21,N_967);
nor U1991 (N_1991,N_269,N_1155);
nor U1992 (N_1992,N_1198,N_3);
xor U1993 (N_1993,N_881,N_41);
nor U1994 (N_1994,N_661,N_760);
xnor U1995 (N_1995,N_1255,N_1167);
or U1996 (N_1996,N_1200,N_812);
nor U1997 (N_1997,N_195,N_1273);
xor U1998 (N_1998,N_807,N_376);
nor U1999 (N_1999,N_220,N_95);
or U2000 (N_2000,N_1481,N_388);
nand U2001 (N_2001,N_744,N_733);
xor U2002 (N_2002,N_1096,N_201);
xor U2003 (N_2003,N_847,N_630);
and U2004 (N_2004,N_91,N_1284);
and U2005 (N_2005,N_937,N_643);
nor U2006 (N_2006,N_497,N_1301);
nand U2007 (N_2007,N_1236,N_28);
nor U2008 (N_2008,N_1445,N_1124);
nor U2009 (N_2009,N_245,N_1109);
nand U2010 (N_2010,N_746,N_471);
nand U2011 (N_2011,N_1288,N_490);
nand U2012 (N_2012,N_1103,N_159);
xor U2013 (N_2013,N_905,N_1382);
xnor U2014 (N_2014,N_1307,N_1332);
and U2015 (N_2015,N_1108,N_687);
and U2016 (N_2016,N_997,N_862);
nor U2017 (N_2017,N_1182,N_685);
and U2018 (N_2018,N_602,N_122);
or U2019 (N_2019,N_1146,N_691);
or U2020 (N_2020,N_1050,N_656);
or U2021 (N_2021,N_1047,N_338);
or U2022 (N_2022,N_93,N_1278);
or U2023 (N_2023,N_986,N_1281);
or U2024 (N_2024,N_1456,N_1091);
nor U2025 (N_2025,N_1114,N_1016);
xor U2026 (N_2026,N_76,N_878);
nor U2027 (N_2027,N_592,N_1119);
xnor U2028 (N_2028,N_1483,N_1400);
and U2029 (N_2029,N_724,N_489);
or U2030 (N_2030,N_1350,N_897);
nor U2031 (N_2031,N_200,N_504);
nand U2032 (N_2032,N_1002,N_956);
or U2033 (N_2033,N_985,N_273);
nand U2034 (N_2034,N_774,N_768);
xor U2035 (N_2035,N_400,N_900);
nand U2036 (N_2036,N_822,N_589);
nand U2037 (N_2037,N_543,N_568);
and U2038 (N_2038,N_176,N_390);
nand U2039 (N_2039,N_69,N_172);
nor U2040 (N_2040,N_969,N_294);
nand U2041 (N_2041,N_293,N_850);
nand U2042 (N_2042,N_1308,N_629);
or U2043 (N_2043,N_761,N_181);
xor U2044 (N_2044,N_752,N_892);
nand U2045 (N_2045,N_430,N_575);
nand U2046 (N_2046,N_1194,N_1113);
xor U2047 (N_2047,N_9,N_330);
xor U2048 (N_2048,N_472,N_1087);
nor U2049 (N_2049,N_1405,N_1204);
nand U2050 (N_2050,N_1433,N_549);
xor U2051 (N_2051,N_972,N_65);
nor U2052 (N_2052,N_186,N_128);
and U2053 (N_2053,N_1048,N_935);
nand U2054 (N_2054,N_1011,N_712);
xnor U2055 (N_2055,N_715,N_1380);
nand U2056 (N_2056,N_1462,N_631);
nand U2057 (N_2057,N_206,N_570);
and U2058 (N_2058,N_483,N_756);
and U2059 (N_2059,N_1141,N_1300);
xor U2060 (N_2060,N_285,N_880);
and U2061 (N_2061,N_143,N_1241);
nor U2062 (N_2062,N_134,N_1121);
and U2063 (N_2063,N_1245,N_117);
xnor U2064 (N_2064,N_659,N_776);
nand U2065 (N_2065,N_795,N_378);
nor U2066 (N_2066,N_73,N_487);
nand U2067 (N_2067,N_741,N_920);
xor U2068 (N_2068,N_1457,N_1199);
xnor U2069 (N_2069,N_146,N_182);
or U2070 (N_2070,N_494,N_711);
nand U2071 (N_2071,N_288,N_1379);
nor U2072 (N_2072,N_678,N_466);
nor U2073 (N_2073,N_315,N_249);
nor U2074 (N_2074,N_217,N_1013);
nand U2075 (N_2075,N_1000,N_1084);
and U2076 (N_2076,N_99,N_1466);
nor U2077 (N_2077,N_915,N_953);
or U2078 (N_2078,N_27,N_1174);
xor U2079 (N_2079,N_595,N_918);
or U2080 (N_2080,N_360,N_1134);
and U2081 (N_2081,N_1205,N_876);
and U2082 (N_2082,N_137,N_1208);
nor U2083 (N_2083,N_280,N_1448);
nor U2084 (N_2084,N_399,N_284);
nand U2085 (N_2085,N_94,N_923);
xor U2086 (N_2086,N_513,N_1401);
xnor U2087 (N_2087,N_414,N_505);
nor U2088 (N_2088,N_1443,N_1437);
and U2089 (N_2089,N_594,N_1034);
xor U2090 (N_2090,N_639,N_889);
nand U2091 (N_2091,N_1299,N_116);
nor U2092 (N_2092,N_67,N_1190);
nor U2093 (N_2093,N_383,N_686);
xnor U2094 (N_2094,N_1250,N_695);
xor U2095 (N_2095,N_1452,N_932);
nand U2096 (N_2096,N_934,N_1415);
xnor U2097 (N_2097,N_449,N_358);
and U2098 (N_2098,N_1381,N_197);
xor U2099 (N_2099,N_451,N_735);
and U2100 (N_2100,N_1356,N_1135);
and U2101 (N_2101,N_802,N_1291);
xnor U2102 (N_2102,N_501,N_168);
and U2103 (N_2103,N_959,N_664);
nand U2104 (N_2104,N_1001,N_961);
and U2105 (N_2105,N_1285,N_800);
xnor U2106 (N_2106,N_1165,N_1242);
xnor U2107 (N_2107,N_1189,N_917);
xor U2108 (N_2108,N_177,N_1078);
nand U2109 (N_2109,N_20,N_1023);
nand U2110 (N_2110,N_1029,N_966);
nor U2111 (N_2111,N_719,N_1477);
or U2112 (N_2112,N_127,N_1487);
and U2113 (N_2113,N_149,N_33);
or U2114 (N_2114,N_994,N_911);
and U2115 (N_2115,N_925,N_1432);
and U2116 (N_2116,N_660,N_605);
or U2117 (N_2117,N_281,N_341);
xor U2118 (N_2118,N_1454,N_140);
xnor U2119 (N_2119,N_1367,N_23);
and U2120 (N_2120,N_799,N_755);
xnor U2121 (N_2121,N_684,N_499);
xnor U2122 (N_2122,N_846,N_929);
or U2123 (N_2123,N_1244,N_15);
and U2124 (N_2124,N_239,N_1329);
nor U2125 (N_2125,N_1485,N_345);
nand U2126 (N_2126,N_421,N_910);
nand U2127 (N_2127,N_1026,N_387);
or U2128 (N_2128,N_1035,N_1423);
nand U2129 (N_2129,N_304,N_625);
xor U2130 (N_2130,N_232,N_936);
nand U2131 (N_2131,N_1293,N_305);
nand U2132 (N_2132,N_196,N_412);
nand U2133 (N_2133,N_940,N_1306);
xor U2134 (N_2134,N_441,N_895);
nor U2135 (N_2135,N_264,N_343);
nand U2136 (N_2136,N_1272,N_557);
nand U2137 (N_2137,N_110,N_54);
or U2138 (N_2138,N_258,N_1344);
and U2139 (N_2139,N_838,N_202);
nand U2140 (N_2140,N_821,N_398);
xnor U2141 (N_2141,N_540,N_1497);
or U2142 (N_2142,N_179,N_1004);
nand U2143 (N_2143,N_601,N_154);
and U2144 (N_2144,N_1494,N_814);
or U2145 (N_2145,N_519,N_58);
and U2146 (N_2146,N_171,N_75);
or U2147 (N_2147,N_617,N_620);
nand U2148 (N_2148,N_1325,N_858);
or U2149 (N_2149,N_142,N_1315);
xnor U2150 (N_2150,N_310,N_148);
and U2151 (N_2151,N_1156,N_1025);
xor U2152 (N_2152,N_849,N_296);
or U2153 (N_2153,N_957,N_290);
nand U2154 (N_2154,N_1266,N_968);
and U2155 (N_2155,N_1416,N_462);
nand U2156 (N_2156,N_278,N_762);
nor U2157 (N_2157,N_319,N_417);
and U2158 (N_2158,N_512,N_90);
xor U2159 (N_2159,N_1387,N_86);
nor U2160 (N_2160,N_433,N_1018);
nor U2161 (N_2161,N_622,N_1277);
and U2162 (N_2162,N_365,N_426);
nand U2163 (N_2163,N_700,N_103);
nand U2164 (N_2164,N_161,N_87);
nor U2165 (N_2165,N_507,N_1095);
nor U2166 (N_2166,N_234,N_884);
nor U2167 (N_2167,N_572,N_841);
xor U2168 (N_2168,N_1271,N_129);
xnor U2169 (N_2169,N_30,N_1264);
nand U2170 (N_2170,N_843,N_1323);
xor U2171 (N_2171,N_1188,N_1191);
or U2172 (N_2172,N_798,N_496);
nor U2173 (N_2173,N_1404,N_1231);
xnor U2174 (N_2174,N_1030,N_662);
and U2175 (N_2175,N_309,N_1465);
and U2176 (N_2176,N_266,N_1472);
xnor U2177 (N_2177,N_1391,N_38);
or U2178 (N_2178,N_523,N_226);
nand U2179 (N_2179,N_61,N_130);
and U2180 (N_2180,N_408,N_1093);
nor U2181 (N_2181,N_1490,N_699);
and U2182 (N_2182,N_211,N_748);
or U2183 (N_2183,N_164,N_100);
nor U2184 (N_2184,N_1234,N_1492);
xor U2185 (N_2185,N_1222,N_1441);
nor U2186 (N_2186,N_185,N_1392);
and U2187 (N_2187,N_648,N_764);
xor U2188 (N_2188,N_256,N_478);
and U2189 (N_2189,N_1248,N_785);
nand U2190 (N_2190,N_965,N_1414);
or U2191 (N_2191,N_1482,N_1336);
nor U2192 (N_2192,N_1226,N_407);
nand U2193 (N_2193,N_1127,N_556);
nor U2194 (N_2194,N_351,N_436);
nor U2195 (N_2195,N_1137,N_52);
nor U2196 (N_2196,N_402,N_1410);
and U2197 (N_2197,N_209,N_397);
and U2198 (N_2198,N_1074,N_144);
and U2199 (N_2199,N_331,N_693);
xnor U2200 (N_2200,N_533,N_1052);
and U2201 (N_2201,N_1309,N_771);
or U2202 (N_2202,N_359,N_437);
xnor U2203 (N_2203,N_1374,N_45);
nor U2204 (N_2204,N_374,N_1251);
nor U2205 (N_2205,N_713,N_476);
or U2206 (N_2206,N_870,N_357);
nor U2207 (N_2207,N_692,N_1225);
xnor U2208 (N_2208,N_867,N_26);
xnor U2209 (N_2209,N_277,N_826);
and U2210 (N_2210,N_583,N_1260);
nand U2211 (N_2211,N_633,N_242);
nor U2212 (N_2212,N_477,N_529);
nand U2213 (N_2213,N_1240,N_301);
and U2214 (N_2214,N_808,N_909);
nor U2215 (N_2215,N_616,N_971);
nand U2216 (N_2216,N_344,N_1131);
xnor U2217 (N_2217,N_11,N_1394);
or U2218 (N_2218,N_104,N_783);
nor U2219 (N_2219,N_1112,N_689);
xnor U2220 (N_2220,N_919,N_663);
and U2221 (N_2221,N_1149,N_706);
nand U2222 (N_2222,N_1070,N_150);
and U2223 (N_2223,N_322,N_723);
nor U2224 (N_2224,N_49,N_955);
xnor U2225 (N_2225,N_1402,N_970);
xor U2226 (N_2226,N_1224,N_1012);
and U2227 (N_2227,N_1040,N_1471);
xnor U2228 (N_2228,N_888,N_1377);
and U2229 (N_2229,N_1347,N_364);
and U2230 (N_2230,N_792,N_425);
nor U2231 (N_2231,N_1434,N_701);
xor U2232 (N_2232,N_1075,N_1268);
or U2233 (N_2233,N_108,N_1054);
and U2234 (N_2234,N_133,N_1499);
nor U2235 (N_2235,N_1170,N_727);
or U2236 (N_2236,N_297,N_131);
xor U2237 (N_2237,N_564,N_1116);
nor U2238 (N_2238,N_467,N_136);
and U2239 (N_2239,N_941,N_10);
and U2240 (N_2240,N_1326,N_435);
nand U2241 (N_2241,N_770,N_1425);
nor U2242 (N_2242,N_1195,N_922);
or U2243 (N_2243,N_160,N_1220);
and U2244 (N_2244,N_749,N_1055);
nor U2245 (N_2245,N_725,N_361);
nor U2246 (N_2246,N_68,N_1334);
nor U2247 (N_2247,N_1498,N_1088);
or U2248 (N_2248,N_342,N_824);
xor U2249 (N_2249,N_190,N_1246);
and U2250 (N_2250,N_431,N_1047);
xor U2251 (N_2251,N_891,N_61);
nor U2252 (N_2252,N_1017,N_453);
xnor U2253 (N_2253,N_657,N_520);
nand U2254 (N_2254,N_1289,N_1174);
nor U2255 (N_2255,N_235,N_410);
and U2256 (N_2256,N_680,N_198);
xor U2257 (N_2257,N_1197,N_114);
nand U2258 (N_2258,N_1294,N_707);
nor U2259 (N_2259,N_1462,N_379);
nor U2260 (N_2260,N_500,N_1047);
nand U2261 (N_2261,N_1398,N_257);
nand U2262 (N_2262,N_943,N_1187);
nor U2263 (N_2263,N_363,N_155);
or U2264 (N_2264,N_1446,N_524);
nor U2265 (N_2265,N_772,N_582);
or U2266 (N_2266,N_1436,N_227);
or U2267 (N_2267,N_953,N_601);
and U2268 (N_2268,N_161,N_410);
xor U2269 (N_2269,N_1478,N_772);
nand U2270 (N_2270,N_804,N_621);
and U2271 (N_2271,N_42,N_214);
nor U2272 (N_2272,N_913,N_790);
xor U2273 (N_2273,N_541,N_921);
xor U2274 (N_2274,N_20,N_1357);
xor U2275 (N_2275,N_608,N_1371);
and U2276 (N_2276,N_1367,N_563);
and U2277 (N_2277,N_957,N_1343);
or U2278 (N_2278,N_525,N_611);
xor U2279 (N_2279,N_428,N_155);
nor U2280 (N_2280,N_1446,N_856);
nor U2281 (N_2281,N_1325,N_461);
and U2282 (N_2282,N_1445,N_1221);
and U2283 (N_2283,N_597,N_775);
and U2284 (N_2284,N_1297,N_1451);
and U2285 (N_2285,N_810,N_1494);
nand U2286 (N_2286,N_1474,N_555);
xor U2287 (N_2287,N_789,N_1306);
and U2288 (N_2288,N_1093,N_195);
nand U2289 (N_2289,N_750,N_170);
or U2290 (N_2290,N_1150,N_941);
xor U2291 (N_2291,N_1179,N_916);
xor U2292 (N_2292,N_1200,N_695);
nor U2293 (N_2293,N_699,N_750);
nand U2294 (N_2294,N_907,N_964);
nand U2295 (N_2295,N_288,N_88);
and U2296 (N_2296,N_728,N_799);
nand U2297 (N_2297,N_572,N_453);
and U2298 (N_2298,N_934,N_391);
nand U2299 (N_2299,N_1075,N_861);
and U2300 (N_2300,N_207,N_683);
and U2301 (N_2301,N_900,N_743);
and U2302 (N_2302,N_1197,N_839);
or U2303 (N_2303,N_391,N_1063);
xnor U2304 (N_2304,N_474,N_82);
nand U2305 (N_2305,N_1282,N_141);
xor U2306 (N_2306,N_1308,N_976);
nor U2307 (N_2307,N_209,N_1162);
and U2308 (N_2308,N_455,N_374);
and U2309 (N_2309,N_1164,N_575);
nor U2310 (N_2310,N_833,N_809);
nor U2311 (N_2311,N_1406,N_1150);
xor U2312 (N_2312,N_1298,N_75);
nand U2313 (N_2313,N_1377,N_38);
nor U2314 (N_2314,N_486,N_539);
or U2315 (N_2315,N_991,N_1401);
nand U2316 (N_2316,N_796,N_206);
nor U2317 (N_2317,N_1273,N_70);
or U2318 (N_2318,N_1096,N_1356);
nor U2319 (N_2319,N_1455,N_1387);
nor U2320 (N_2320,N_79,N_522);
and U2321 (N_2321,N_397,N_523);
or U2322 (N_2322,N_70,N_1033);
and U2323 (N_2323,N_239,N_636);
and U2324 (N_2324,N_1294,N_201);
or U2325 (N_2325,N_990,N_751);
nand U2326 (N_2326,N_1312,N_340);
nand U2327 (N_2327,N_1102,N_1494);
nand U2328 (N_2328,N_1343,N_539);
or U2329 (N_2329,N_1076,N_1372);
xor U2330 (N_2330,N_1482,N_1015);
or U2331 (N_2331,N_654,N_1420);
xnor U2332 (N_2332,N_659,N_943);
or U2333 (N_2333,N_1373,N_631);
xor U2334 (N_2334,N_486,N_295);
and U2335 (N_2335,N_196,N_743);
nand U2336 (N_2336,N_1062,N_263);
or U2337 (N_2337,N_120,N_715);
nor U2338 (N_2338,N_1044,N_703);
xnor U2339 (N_2339,N_493,N_91);
or U2340 (N_2340,N_880,N_1176);
and U2341 (N_2341,N_13,N_1046);
and U2342 (N_2342,N_1298,N_978);
nor U2343 (N_2343,N_1073,N_1344);
and U2344 (N_2344,N_1276,N_1485);
nand U2345 (N_2345,N_1098,N_908);
nor U2346 (N_2346,N_1147,N_262);
or U2347 (N_2347,N_1282,N_1380);
and U2348 (N_2348,N_1263,N_211);
or U2349 (N_2349,N_668,N_17);
nand U2350 (N_2350,N_139,N_1491);
xnor U2351 (N_2351,N_713,N_145);
or U2352 (N_2352,N_907,N_75);
xor U2353 (N_2353,N_1179,N_1281);
or U2354 (N_2354,N_480,N_1449);
or U2355 (N_2355,N_602,N_1115);
nand U2356 (N_2356,N_1257,N_905);
xor U2357 (N_2357,N_502,N_941);
or U2358 (N_2358,N_290,N_1334);
or U2359 (N_2359,N_109,N_648);
or U2360 (N_2360,N_215,N_323);
or U2361 (N_2361,N_206,N_1418);
and U2362 (N_2362,N_1052,N_527);
nand U2363 (N_2363,N_336,N_521);
and U2364 (N_2364,N_108,N_757);
and U2365 (N_2365,N_262,N_453);
and U2366 (N_2366,N_1437,N_1345);
or U2367 (N_2367,N_221,N_52);
or U2368 (N_2368,N_359,N_750);
and U2369 (N_2369,N_546,N_1353);
or U2370 (N_2370,N_1213,N_710);
nor U2371 (N_2371,N_855,N_241);
nand U2372 (N_2372,N_739,N_1163);
nand U2373 (N_2373,N_262,N_1268);
nor U2374 (N_2374,N_22,N_584);
or U2375 (N_2375,N_1428,N_945);
nand U2376 (N_2376,N_164,N_1354);
and U2377 (N_2377,N_335,N_815);
or U2378 (N_2378,N_602,N_978);
and U2379 (N_2379,N_840,N_918);
nor U2380 (N_2380,N_617,N_761);
nand U2381 (N_2381,N_1052,N_995);
and U2382 (N_2382,N_598,N_886);
xnor U2383 (N_2383,N_61,N_1044);
and U2384 (N_2384,N_193,N_1133);
and U2385 (N_2385,N_1493,N_1026);
and U2386 (N_2386,N_592,N_84);
and U2387 (N_2387,N_1087,N_1104);
or U2388 (N_2388,N_11,N_460);
and U2389 (N_2389,N_698,N_541);
nand U2390 (N_2390,N_374,N_619);
nand U2391 (N_2391,N_821,N_99);
xnor U2392 (N_2392,N_691,N_744);
nand U2393 (N_2393,N_597,N_803);
or U2394 (N_2394,N_140,N_218);
nor U2395 (N_2395,N_1378,N_16);
and U2396 (N_2396,N_1346,N_1452);
nand U2397 (N_2397,N_375,N_292);
and U2398 (N_2398,N_520,N_1482);
and U2399 (N_2399,N_51,N_989);
xnor U2400 (N_2400,N_1254,N_413);
nor U2401 (N_2401,N_1089,N_1129);
or U2402 (N_2402,N_1334,N_967);
and U2403 (N_2403,N_1289,N_1469);
nand U2404 (N_2404,N_1097,N_718);
nand U2405 (N_2405,N_357,N_986);
and U2406 (N_2406,N_737,N_1204);
and U2407 (N_2407,N_214,N_336);
and U2408 (N_2408,N_895,N_605);
or U2409 (N_2409,N_746,N_1116);
nor U2410 (N_2410,N_1027,N_354);
or U2411 (N_2411,N_1036,N_630);
and U2412 (N_2412,N_1322,N_808);
and U2413 (N_2413,N_283,N_1246);
nand U2414 (N_2414,N_85,N_195);
and U2415 (N_2415,N_387,N_1111);
and U2416 (N_2416,N_1417,N_1048);
xnor U2417 (N_2417,N_1307,N_109);
xnor U2418 (N_2418,N_282,N_589);
or U2419 (N_2419,N_940,N_592);
and U2420 (N_2420,N_818,N_1430);
and U2421 (N_2421,N_47,N_311);
or U2422 (N_2422,N_1491,N_644);
nand U2423 (N_2423,N_735,N_515);
nor U2424 (N_2424,N_950,N_590);
xnor U2425 (N_2425,N_1059,N_1438);
and U2426 (N_2426,N_466,N_123);
nand U2427 (N_2427,N_1207,N_1330);
nand U2428 (N_2428,N_1426,N_1451);
xnor U2429 (N_2429,N_1301,N_422);
nand U2430 (N_2430,N_1380,N_1031);
xor U2431 (N_2431,N_911,N_824);
or U2432 (N_2432,N_1213,N_1198);
and U2433 (N_2433,N_979,N_716);
or U2434 (N_2434,N_929,N_483);
or U2435 (N_2435,N_242,N_1083);
xor U2436 (N_2436,N_292,N_390);
xor U2437 (N_2437,N_1456,N_1408);
xnor U2438 (N_2438,N_1120,N_329);
nor U2439 (N_2439,N_810,N_608);
nor U2440 (N_2440,N_567,N_1081);
nand U2441 (N_2441,N_699,N_709);
nand U2442 (N_2442,N_615,N_790);
xor U2443 (N_2443,N_1036,N_565);
xnor U2444 (N_2444,N_956,N_33);
xnor U2445 (N_2445,N_1404,N_1376);
nand U2446 (N_2446,N_684,N_815);
or U2447 (N_2447,N_286,N_213);
and U2448 (N_2448,N_214,N_1383);
nand U2449 (N_2449,N_407,N_1204);
xnor U2450 (N_2450,N_770,N_484);
nor U2451 (N_2451,N_843,N_217);
nor U2452 (N_2452,N_694,N_888);
and U2453 (N_2453,N_368,N_563);
xnor U2454 (N_2454,N_790,N_1175);
nor U2455 (N_2455,N_515,N_163);
or U2456 (N_2456,N_511,N_1367);
xnor U2457 (N_2457,N_814,N_1205);
xnor U2458 (N_2458,N_465,N_557);
nand U2459 (N_2459,N_1181,N_798);
nor U2460 (N_2460,N_185,N_1072);
nor U2461 (N_2461,N_334,N_13);
nand U2462 (N_2462,N_651,N_661);
nand U2463 (N_2463,N_912,N_445);
xnor U2464 (N_2464,N_295,N_610);
and U2465 (N_2465,N_822,N_342);
xnor U2466 (N_2466,N_1410,N_908);
and U2467 (N_2467,N_759,N_798);
nand U2468 (N_2468,N_1447,N_798);
and U2469 (N_2469,N_451,N_995);
nand U2470 (N_2470,N_702,N_862);
and U2471 (N_2471,N_925,N_767);
or U2472 (N_2472,N_403,N_252);
nand U2473 (N_2473,N_961,N_1084);
nor U2474 (N_2474,N_813,N_791);
xnor U2475 (N_2475,N_504,N_1352);
xnor U2476 (N_2476,N_1117,N_1299);
and U2477 (N_2477,N_1122,N_12);
or U2478 (N_2478,N_220,N_410);
nor U2479 (N_2479,N_449,N_839);
nand U2480 (N_2480,N_1101,N_573);
and U2481 (N_2481,N_1485,N_18);
nand U2482 (N_2482,N_1412,N_1156);
nor U2483 (N_2483,N_146,N_367);
nor U2484 (N_2484,N_1396,N_132);
nor U2485 (N_2485,N_290,N_1446);
xor U2486 (N_2486,N_1452,N_182);
xor U2487 (N_2487,N_117,N_1122);
xnor U2488 (N_2488,N_1078,N_746);
xnor U2489 (N_2489,N_1215,N_1255);
and U2490 (N_2490,N_1331,N_431);
or U2491 (N_2491,N_958,N_1402);
nand U2492 (N_2492,N_918,N_458);
or U2493 (N_2493,N_1128,N_966);
or U2494 (N_2494,N_1177,N_666);
nand U2495 (N_2495,N_1251,N_1334);
nor U2496 (N_2496,N_51,N_836);
nand U2497 (N_2497,N_1483,N_308);
xnor U2498 (N_2498,N_944,N_158);
and U2499 (N_2499,N_6,N_909);
xnor U2500 (N_2500,N_861,N_1479);
nor U2501 (N_2501,N_1093,N_1320);
or U2502 (N_2502,N_415,N_756);
xor U2503 (N_2503,N_912,N_1088);
or U2504 (N_2504,N_655,N_1441);
or U2505 (N_2505,N_1277,N_1293);
nand U2506 (N_2506,N_489,N_1353);
nor U2507 (N_2507,N_1055,N_112);
nand U2508 (N_2508,N_916,N_749);
nand U2509 (N_2509,N_585,N_52);
or U2510 (N_2510,N_1093,N_401);
nor U2511 (N_2511,N_914,N_297);
and U2512 (N_2512,N_1375,N_621);
or U2513 (N_2513,N_931,N_612);
and U2514 (N_2514,N_637,N_783);
xor U2515 (N_2515,N_1450,N_1489);
and U2516 (N_2516,N_455,N_1347);
or U2517 (N_2517,N_1195,N_491);
and U2518 (N_2518,N_708,N_338);
and U2519 (N_2519,N_351,N_651);
nor U2520 (N_2520,N_117,N_609);
xnor U2521 (N_2521,N_1157,N_836);
nand U2522 (N_2522,N_917,N_1148);
nor U2523 (N_2523,N_924,N_1055);
nor U2524 (N_2524,N_1329,N_898);
nand U2525 (N_2525,N_609,N_380);
nor U2526 (N_2526,N_951,N_87);
nor U2527 (N_2527,N_27,N_1385);
and U2528 (N_2528,N_1293,N_802);
and U2529 (N_2529,N_1347,N_1213);
and U2530 (N_2530,N_346,N_905);
xnor U2531 (N_2531,N_986,N_343);
xnor U2532 (N_2532,N_1311,N_1247);
nor U2533 (N_2533,N_1149,N_758);
xor U2534 (N_2534,N_1441,N_1433);
or U2535 (N_2535,N_614,N_1274);
nor U2536 (N_2536,N_1317,N_1190);
xor U2537 (N_2537,N_839,N_274);
and U2538 (N_2538,N_970,N_1201);
xnor U2539 (N_2539,N_497,N_1214);
and U2540 (N_2540,N_251,N_621);
or U2541 (N_2541,N_360,N_645);
nor U2542 (N_2542,N_254,N_1354);
xor U2543 (N_2543,N_1050,N_1402);
nor U2544 (N_2544,N_1470,N_235);
nand U2545 (N_2545,N_801,N_857);
nor U2546 (N_2546,N_986,N_743);
and U2547 (N_2547,N_1125,N_738);
nand U2548 (N_2548,N_506,N_1048);
and U2549 (N_2549,N_184,N_1346);
nor U2550 (N_2550,N_248,N_22);
and U2551 (N_2551,N_229,N_740);
nor U2552 (N_2552,N_331,N_109);
xor U2553 (N_2553,N_49,N_89);
and U2554 (N_2554,N_347,N_194);
and U2555 (N_2555,N_567,N_590);
nand U2556 (N_2556,N_647,N_1125);
or U2557 (N_2557,N_28,N_227);
and U2558 (N_2558,N_14,N_140);
or U2559 (N_2559,N_445,N_437);
nor U2560 (N_2560,N_1069,N_678);
xor U2561 (N_2561,N_1431,N_911);
or U2562 (N_2562,N_1434,N_27);
nand U2563 (N_2563,N_1399,N_1249);
nand U2564 (N_2564,N_1132,N_926);
nor U2565 (N_2565,N_78,N_236);
or U2566 (N_2566,N_1075,N_58);
xnor U2567 (N_2567,N_468,N_553);
and U2568 (N_2568,N_1192,N_953);
nor U2569 (N_2569,N_378,N_1089);
nand U2570 (N_2570,N_387,N_513);
xnor U2571 (N_2571,N_1056,N_1251);
xnor U2572 (N_2572,N_788,N_121);
nand U2573 (N_2573,N_792,N_1157);
nand U2574 (N_2574,N_372,N_1182);
nand U2575 (N_2575,N_359,N_610);
xnor U2576 (N_2576,N_105,N_1136);
nand U2577 (N_2577,N_1345,N_507);
or U2578 (N_2578,N_89,N_90);
or U2579 (N_2579,N_1026,N_1329);
and U2580 (N_2580,N_545,N_1372);
nor U2581 (N_2581,N_1190,N_723);
and U2582 (N_2582,N_375,N_822);
or U2583 (N_2583,N_84,N_908);
nor U2584 (N_2584,N_1147,N_841);
nand U2585 (N_2585,N_735,N_692);
or U2586 (N_2586,N_176,N_640);
or U2587 (N_2587,N_1105,N_416);
xnor U2588 (N_2588,N_949,N_109);
or U2589 (N_2589,N_130,N_167);
nand U2590 (N_2590,N_496,N_458);
and U2591 (N_2591,N_1461,N_1490);
nor U2592 (N_2592,N_1479,N_431);
or U2593 (N_2593,N_790,N_873);
or U2594 (N_2594,N_388,N_1282);
xor U2595 (N_2595,N_205,N_387);
and U2596 (N_2596,N_1002,N_362);
or U2597 (N_2597,N_1387,N_1220);
and U2598 (N_2598,N_663,N_731);
xor U2599 (N_2599,N_501,N_406);
or U2600 (N_2600,N_157,N_1160);
nand U2601 (N_2601,N_998,N_676);
nand U2602 (N_2602,N_1189,N_69);
nand U2603 (N_2603,N_779,N_1154);
or U2604 (N_2604,N_1327,N_494);
or U2605 (N_2605,N_11,N_857);
or U2606 (N_2606,N_1428,N_793);
nand U2607 (N_2607,N_594,N_560);
and U2608 (N_2608,N_1412,N_1240);
xnor U2609 (N_2609,N_236,N_1290);
or U2610 (N_2610,N_1086,N_791);
and U2611 (N_2611,N_377,N_752);
nand U2612 (N_2612,N_856,N_250);
xnor U2613 (N_2613,N_965,N_916);
nor U2614 (N_2614,N_1043,N_126);
nor U2615 (N_2615,N_39,N_1006);
or U2616 (N_2616,N_335,N_383);
nand U2617 (N_2617,N_1338,N_472);
and U2618 (N_2618,N_1247,N_593);
and U2619 (N_2619,N_570,N_72);
nand U2620 (N_2620,N_932,N_1272);
or U2621 (N_2621,N_1450,N_1173);
xnor U2622 (N_2622,N_405,N_49);
nor U2623 (N_2623,N_407,N_154);
xnor U2624 (N_2624,N_569,N_1193);
xnor U2625 (N_2625,N_1150,N_444);
nand U2626 (N_2626,N_877,N_442);
nand U2627 (N_2627,N_882,N_635);
or U2628 (N_2628,N_1126,N_750);
nand U2629 (N_2629,N_1381,N_1152);
nand U2630 (N_2630,N_412,N_909);
nor U2631 (N_2631,N_915,N_836);
nor U2632 (N_2632,N_1098,N_1323);
xnor U2633 (N_2633,N_1236,N_172);
xnor U2634 (N_2634,N_405,N_583);
and U2635 (N_2635,N_1107,N_1409);
or U2636 (N_2636,N_881,N_1299);
xor U2637 (N_2637,N_1499,N_1036);
xnor U2638 (N_2638,N_473,N_273);
and U2639 (N_2639,N_1447,N_414);
xnor U2640 (N_2640,N_536,N_1117);
nor U2641 (N_2641,N_255,N_879);
and U2642 (N_2642,N_1347,N_712);
nand U2643 (N_2643,N_274,N_1279);
and U2644 (N_2644,N_824,N_1293);
nand U2645 (N_2645,N_1444,N_569);
xnor U2646 (N_2646,N_1238,N_961);
and U2647 (N_2647,N_376,N_757);
or U2648 (N_2648,N_956,N_1027);
nand U2649 (N_2649,N_141,N_1486);
nor U2650 (N_2650,N_591,N_1081);
nand U2651 (N_2651,N_253,N_1326);
and U2652 (N_2652,N_903,N_255);
nor U2653 (N_2653,N_393,N_980);
nor U2654 (N_2654,N_1027,N_916);
nand U2655 (N_2655,N_1181,N_1285);
nor U2656 (N_2656,N_19,N_1249);
nor U2657 (N_2657,N_128,N_863);
and U2658 (N_2658,N_862,N_976);
or U2659 (N_2659,N_398,N_1332);
or U2660 (N_2660,N_426,N_1049);
or U2661 (N_2661,N_312,N_135);
nand U2662 (N_2662,N_426,N_55);
nor U2663 (N_2663,N_1006,N_630);
nor U2664 (N_2664,N_654,N_758);
nand U2665 (N_2665,N_818,N_993);
nand U2666 (N_2666,N_810,N_118);
or U2667 (N_2667,N_40,N_234);
or U2668 (N_2668,N_1313,N_922);
and U2669 (N_2669,N_435,N_910);
xor U2670 (N_2670,N_218,N_657);
or U2671 (N_2671,N_1047,N_193);
nand U2672 (N_2672,N_1015,N_265);
nand U2673 (N_2673,N_119,N_903);
nor U2674 (N_2674,N_1432,N_180);
and U2675 (N_2675,N_295,N_968);
or U2676 (N_2676,N_577,N_1077);
nand U2677 (N_2677,N_296,N_179);
or U2678 (N_2678,N_127,N_1172);
and U2679 (N_2679,N_216,N_5);
and U2680 (N_2680,N_817,N_1227);
nor U2681 (N_2681,N_341,N_559);
nand U2682 (N_2682,N_1401,N_131);
and U2683 (N_2683,N_1232,N_149);
nor U2684 (N_2684,N_460,N_598);
nor U2685 (N_2685,N_1464,N_736);
nand U2686 (N_2686,N_496,N_1478);
and U2687 (N_2687,N_1168,N_949);
or U2688 (N_2688,N_978,N_480);
xnor U2689 (N_2689,N_527,N_1443);
nor U2690 (N_2690,N_626,N_991);
and U2691 (N_2691,N_653,N_545);
or U2692 (N_2692,N_227,N_441);
or U2693 (N_2693,N_131,N_1119);
or U2694 (N_2694,N_352,N_127);
or U2695 (N_2695,N_1097,N_1176);
nand U2696 (N_2696,N_1360,N_1058);
xor U2697 (N_2697,N_1034,N_1153);
or U2698 (N_2698,N_1479,N_647);
and U2699 (N_2699,N_401,N_427);
and U2700 (N_2700,N_1418,N_1381);
xor U2701 (N_2701,N_364,N_919);
or U2702 (N_2702,N_1418,N_812);
or U2703 (N_2703,N_637,N_1195);
and U2704 (N_2704,N_435,N_458);
or U2705 (N_2705,N_145,N_61);
and U2706 (N_2706,N_389,N_240);
nand U2707 (N_2707,N_1352,N_411);
nand U2708 (N_2708,N_27,N_1169);
or U2709 (N_2709,N_438,N_82);
or U2710 (N_2710,N_563,N_125);
nand U2711 (N_2711,N_225,N_431);
nor U2712 (N_2712,N_760,N_1338);
and U2713 (N_2713,N_645,N_1150);
or U2714 (N_2714,N_217,N_618);
or U2715 (N_2715,N_1471,N_187);
and U2716 (N_2716,N_291,N_617);
nor U2717 (N_2717,N_193,N_310);
nand U2718 (N_2718,N_1441,N_855);
nand U2719 (N_2719,N_774,N_570);
nor U2720 (N_2720,N_685,N_1404);
and U2721 (N_2721,N_1151,N_894);
nand U2722 (N_2722,N_835,N_396);
and U2723 (N_2723,N_226,N_961);
nor U2724 (N_2724,N_651,N_898);
nor U2725 (N_2725,N_1298,N_158);
and U2726 (N_2726,N_342,N_1236);
nand U2727 (N_2727,N_47,N_920);
xnor U2728 (N_2728,N_1090,N_797);
and U2729 (N_2729,N_243,N_1442);
nand U2730 (N_2730,N_694,N_1430);
nor U2731 (N_2731,N_759,N_318);
nor U2732 (N_2732,N_706,N_1346);
xnor U2733 (N_2733,N_120,N_1339);
and U2734 (N_2734,N_1418,N_968);
and U2735 (N_2735,N_612,N_563);
nor U2736 (N_2736,N_1154,N_1234);
nand U2737 (N_2737,N_1157,N_776);
nand U2738 (N_2738,N_139,N_1039);
or U2739 (N_2739,N_1377,N_354);
or U2740 (N_2740,N_642,N_29);
and U2741 (N_2741,N_620,N_326);
xor U2742 (N_2742,N_401,N_1340);
or U2743 (N_2743,N_58,N_1001);
and U2744 (N_2744,N_1060,N_618);
nor U2745 (N_2745,N_968,N_1432);
nor U2746 (N_2746,N_167,N_1340);
and U2747 (N_2747,N_999,N_1276);
xor U2748 (N_2748,N_505,N_294);
xor U2749 (N_2749,N_878,N_925);
nor U2750 (N_2750,N_85,N_730);
xor U2751 (N_2751,N_475,N_54);
nand U2752 (N_2752,N_94,N_746);
xor U2753 (N_2753,N_167,N_259);
nor U2754 (N_2754,N_376,N_507);
xnor U2755 (N_2755,N_134,N_205);
and U2756 (N_2756,N_90,N_1496);
nor U2757 (N_2757,N_432,N_592);
or U2758 (N_2758,N_1448,N_810);
nor U2759 (N_2759,N_478,N_960);
nand U2760 (N_2760,N_271,N_537);
xnor U2761 (N_2761,N_361,N_94);
and U2762 (N_2762,N_1236,N_1279);
nand U2763 (N_2763,N_190,N_604);
or U2764 (N_2764,N_1007,N_1283);
nor U2765 (N_2765,N_826,N_625);
nor U2766 (N_2766,N_1482,N_81);
xnor U2767 (N_2767,N_869,N_1489);
nand U2768 (N_2768,N_105,N_1330);
xor U2769 (N_2769,N_204,N_1183);
or U2770 (N_2770,N_678,N_837);
nand U2771 (N_2771,N_247,N_343);
and U2772 (N_2772,N_1265,N_995);
and U2773 (N_2773,N_397,N_622);
nor U2774 (N_2774,N_557,N_796);
nor U2775 (N_2775,N_582,N_1490);
nand U2776 (N_2776,N_1350,N_761);
nand U2777 (N_2777,N_1174,N_1469);
and U2778 (N_2778,N_126,N_1087);
and U2779 (N_2779,N_1014,N_627);
or U2780 (N_2780,N_1299,N_795);
xor U2781 (N_2781,N_338,N_379);
nand U2782 (N_2782,N_1383,N_1001);
nor U2783 (N_2783,N_192,N_126);
nand U2784 (N_2784,N_124,N_866);
and U2785 (N_2785,N_76,N_1222);
and U2786 (N_2786,N_1226,N_162);
or U2787 (N_2787,N_156,N_46);
nand U2788 (N_2788,N_1109,N_493);
and U2789 (N_2789,N_687,N_938);
xnor U2790 (N_2790,N_239,N_475);
or U2791 (N_2791,N_802,N_548);
or U2792 (N_2792,N_582,N_850);
and U2793 (N_2793,N_1115,N_1297);
xnor U2794 (N_2794,N_1454,N_888);
xor U2795 (N_2795,N_321,N_221);
xor U2796 (N_2796,N_1223,N_366);
nand U2797 (N_2797,N_920,N_1392);
or U2798 (N_2798,N_1296,N_219);
nor U2799 (N_2799,N_1327,N_172);
nand U2800 (N_2800,N_1477,N_714);
xnor U2801 (N_2801,N_1211,N_1147);
nand U2802 (N_2802,N_503,N_619);
nand U2803 (N_2803,N_1112,N_1209);
or U2804 (N_2804,N_1274,N_126);
nor U2805 (N_2805,N_159,N_264);
nand U2806 (N_2806,N_874,N_1093);
nor U2807 (N_2807,N_93,N_894);
xnor U2808 (N_2808,N_755,N_647);
nor U2809 (N_2809,N_126,N_729);
xnor U2810 (N_2810,N_15,N_262);
nor U2811 (N_2811,N_1055,N_317);
nor U2812 (N_2812,N_1343,N_755);
xnor U2813 (N_2813,N_504,N_432);
nor U2814 (N_2814,N_1165,N_1287);
or U2815 (N_2815,N_986,N_662);
and U2816 (N_2816,N_261,N_564);
and U2817 (N_2817,N_887,N_551);
nand U2818 (N_2818,N_1251,N_318);
xnor U2819 (N_2819,N_503,N_775);
nor U2820 (N_2820,N_966,N_1093);
or U2821 (N_2821,N_1479,N_898);
xnor U2822 (N_2822,N_68,N_397);
xor U2823 (N_2823,N_232,N_96);
xnor U2824 (N_2824,N_1432,N_541);
or U2825 (N_2825,N_604,N_844);
nor U2826 (N_2826,N_135,N_1314);
xor U2827 (N_2827,N_144,N_314);
and U2828 (N_2828,N_893,N_1435);
or U2829 (N_2829,N_761,N_662);
and U2830 (N_2830,N_465,N_284);
nor U2831 (N_2831,N_358,N_92);
or U2832 (N_2832,N_837,N_1308);
nand U2833 (N_2833,N_182,N_338);
or U2834 (N_2834,N_83,N_458);
or U2835 (N_2835,N_1365,N_1336);
xor U2836 (N_2836,N_568,N_421);
nand U2837 (N_2837,N_574,N_893);
or U2838 (N_2838,N_1394,N_1477);
or U2839 (N_2839,N_1010,N_1396);
and U2840 (N_2840,N_1354,N_915);
nor U2841 (N_2841,N_226,N_933);
nand U2842 (N_2842,N_747,N_545);
xnor U2843 (N_2843,N_1054,N_706);
nand U2844 (N_2844,N_684,N_1194);
nand U2845 (N_2845,N_788,N_1229);
nor U2846 (N_2846,N_710,N_361);
xnor U2847 (N_2847,N_924,N_516);
nor U2848 (N_2848,N_1215,N_660);
nand U2849 (N_2849,N_740,N_189);
xor U2850 (N_2850,N_769,N_1058);
and U2851 (N_2851,N_923,N_192);
and U2852 (N_2852,N_1002,N_122);
nand U2853 (N_2853,N_1232,N_202);
nor U2854 (N_2854,N_283,N_1491);
and U2855 (N_2855,N_920,N_220);
and U2856 (N_2856,N_1239,N_792);
nor U2857 (N_2857,N_1132,N_508);
and U2858 (N_2858,N_1222,N_561);
nand U2859 (N_2859,N_486,N_887);
nor U2860 (N_2860,N_57,N_132);
xor U2861 (N_2861,N_625,N_28);
and U2862 (N_2862,N_441,N_336);
or U2863 (N_2863,N_306,N_327);
xor U2864 (N_2864,N_347,N_1452);
nor U2865 (N_2865,N_93,N_242);
nand U2866 (N_2866,N_1450,N_1251);
or U2867 (N_2867,N_177,N_224);
or U2868 (N_2868,N_1406,N_902);
nand U2869 (N_2869,N_877,N_270);
nor U2870 (N_2870,N_1223,N_391);
and U2871 (N_2871,N_233,N_619);
xnor U2872 (N_2872,N_1334,N_697);
and U2873 (N_2873,N_1407,N_823);
xnor U2874 (N_2874,N_715,N_678);
nand U2875 (N_2875,N_1224,N_1381);
xnor U2876 (N_2876,N_674,N_885);
nor U2877 (N_2877,N_1396,N_26);
or U2878 (N_2878,N_1349,N_1122);
or U2879 (N_2879,N_1295,N_990);
nand U2880 (N_2880,N_301,N_1146);
xnor U2881 (N_2881,N_391,N_657);
nor U2882 (N_2882,N_290,N_1201);
xor U2883 (N_2883,N_786,N_1023);
xor U2884 (N_2884,N_696,N_773);
nor U2885 (N_2885,N_1239,N_1408);
nor U2886 (N_2886,N_1260,N_1020);
and U2887 (N_2887,N_975,N_1494);
nor U2888 (N_2888,N_1054,N_1286);
or U2889 (N_2889,N_893,N_364);
and U2890 (N_2890,N_435,N_580);
nor U2891 (N_2891,N_1325,N_561);
nor U2892 (N_2892,N_1352,N_547);
nand U2893 (N_2893,N_834,N_339);
nor U2894 (N_2894,N_1180,N_758);
xor U2895 (N_2895,N_412,N_5);
or U2896 (N_2896,N_33,N_866);
and U2897 (N_2897,N_786,N_437);
xor U2898 (N_2898,N_549,N_494);
and U2899 (N_2899,N_21,N_1098);
nor U2900 (N_2900,N_979,N_536);
or U2901 (N_2901,N_591,N_535);
or U2902 (N_2902,N_309,N_653);
nor U2903 (N_2903,N_944,N_37);
xnor U2904 (N_2904,N_596,N_1131);
xor U2905 (N_2905,N_631,N_1226);
xor U2906 (N_2906,N_1088,N_194);
or U2907 (N_2907,N_642,N_522);
or U2908 (N_2908,N_1151,N_1246);
xnor U2909 (N_2909,N_992,N_454);
or U2910 (N_2910,N_173,N_757);
xnor U2911 (N_2911,N_695,N_101);
nor U2912 (N_2912,N_731,N_219);
nand U2913 (N_2913,N_965,N_527);
and U2914 (N_2914,N_105,N_468);
and U2915 (N_2915,N_600,N_1052);
nand U2916 (N_2916,N_1064,N_1383);
or U2917 (N_2917,N_1099,N_373);
nand U2918 (N_2918,N_72,N_717);
and U2919 (N_2919,N_233,N_1024);
nand U2920 (N_2920,N_1403,N_396);
nand U2921 (N_2921,N_760,N_129);
nor U2922 (N_2922,N_1224,N_108);
and U2923 (N_2923,N_936,N_863);
nor U2924 (N_2924,N_441,N_1037);
or U2925 (N_2925,N_687,N_660);
or U2926 (N_2926,N_360,N_66);
xnor U2927 (N_2927,N_1190,N_660);
or U2928 (N_2928,N_460,N_984);
nor U2929 (N_2929,N_126,N_804);
or U2930 (N_2930,N_928,N_156);
nand U2931 (N_2931,N_812,N_338);
nand U2932 (N_2932,N_204,N_1284);
nor U2933 (N_2933,N_360,N_333);
and U2934 (N_2934,N_1174,N_1497);
or U2935 (N_2935,N_1307,N_878);
or U2936 (N_2936,N_926,N_1454);
and U2937 (N_2937,N_946,N_299);
xor U2938 (N_2938,N_1299,N_47);
nand U2939 (N_2939,N_1388,N_462);
nor U2940 (N_2940,N_1471,N_418);
or U2941 (N_2941,N_1015,N_1430);
or U2942 (N_2942,N_391,N_205);
xor U2943 (N_2943,N_480,N_673);
nand U2944 (N_2944,N_619,N_795);
or U2945 (N_2945,N_1349,N_559);
or U2946 (N_2946,N_959,N_1236);
and U2947 (N_2947,N_84,N_1438);
nand U2948 (N_2948,N_1038,N_1274);
xor U2949 (N_2949,N_792,N_603);
xnor U2950 (N_2950,N_880,N_753);
and U2951 (N_2951,N_813,N_1172);
xnor U2952 (N_2952,N_1265,N_1028);
and U2953 (N_2953,N_838,N_883);
or U2954 (N_2954,N_652,N_669);
and U2955 (N_2955,N_38,N_647);
or U2956 (N_2956,N_1039,N_1228);
xor U2957 (N_2957,N_824,N_1229);
xnor U2958 (N_2958,N_18,N_591);
xor U2959 (N_2959,N_776,N_514);
and U2960 (N_2960,N_1414,N_1335);
nor U2961 (N_2961,N_578,N_1407);
or U2962 (N_2962,N_1193,N_1254);
nor U2963 (N_2963,N_226,N_416);
and U2964 (N_2964,N_995,N_809);
or U2965 (N_2965,N_52,N_856);
nand U2966 (N_2966,N_445,N_212);
nor U2967 (N_2967,N_966,N_670);
or U2968 (N_2968,N_0,N_262);
xor U2969 (N_2969,N_824,N_927);
and U2970 (N_2970,N_541,N_239);
nor U2971 (N_2971,N_870,N_934);
or U2972 (N_2972,N_1160,N_1313);
nor U2973 (N_2973,N_1410,N_1248);
and U2974 (N_2974,N_995,N_556);
xor U2975 (N_2975,N_760,N_636);
xnor U2976 (N_2976,N_1413,N_412);
or U2977 (N_2977,N_1091,N_128);
and U2978 (N_2978,N_895,N_225);
xnor U2979 (N_2979,N_1475,N_318);
and U2980 (N_2980,N_83,N_1475);
xnor U2981 (N_2981,N_1065,N_243);
or U2982 (N_2982,N_27,N_766);
nand U2983 (N_2983,N_877,N_134);
nand U2984 (N_2984,N_899,N_1035);
nand U2985 (N_2985,N_328,N_157);
xnor U2986 (N_2986,N_289,N_1227);
nand U2987 (N_2987,N_744,N_373);
or U2988 (N_2988,N_340,N_1255);
or U2989 (N_2989,N_64,N_1417);
and U2990 (N_2990,N_795,N_1138);
and U2991 (N_2991,N_154,N_608);
xor U2992 (N_2992,N_1159,N_239);
nor U2993 (N_2993,N_450,N_928);
nor U2994 (N_2994,N_820,N_1464);
and U2995 (N_2995,N_149,N_162);
or U2996 (N_2996,N_923,N_882);
nor U2997 (N_2997,N_414,N_96);
nand U2998 (N_2998,N_748,N_573);
xnor U2999 (N_2999,N_1,N_1136);
nor U3000 (N_3000,N_2337,N_1749);
or U3001 (N_3001,N_1942,N_2516);
and U3002 (N_3002,N_2169,N_2472);
nor U3003 (N_3003,N_1500,N_2870);
nor U3004 (N_3004,N_2596,N_2595);
and U3005 (N_3005,N_1554,N_2469);
nand U3006 (N_3006,N_2957,N_2612);
or U3007 (N_3007,N_1722,N_1599);
xnor U3008 (N_3008,N_2001,N_2043);
and U3009 (N_3009,N_2526,N_2937);
and U3010 (N_3010,N_1777,N_1565);
or U3011 (N_3011,N_1947,N_1587);
nor U3012 (N_3012,N_2886,N_2325);
xnor U3013 (N_3013,N_2745,N_2108);
nor U3014 (N_3014,N_2319,N_1630);
nor U3015 (N_3015,N_2124,N_2012);
nor U3016 (N_3016,N_1629,N_2266);
nor U3017 (N_3017,N_2307,N_2106);
nand U3018 (N_3018,N_2630,N_2240);
or U3019 (N_3019,N_2386,N_1569);
or U3020 (N_3020,N_1862,N_2770);
xor U3021 (N_3021,N_1919,N_2268);
or U3022 (N_3022,N_1937,N_1639);
nor U3023 (N_3023,N_1971,N_2393);
nand U3024 (N_3024,N_2763,N_2663);
or U3025 (N_3025,N_2423,N_2771);
and U3026 (N_3026,N_1939,N_1622);
or U3027 (N_3027,N_1757,N_2315);
xor U3028 (N_3028,N_2285,N_2738);
xnor U3029 (N_3029,N_2326,N_2015);
xor U3030 (N_3030,N_2267,N_2504);
or U3031 (N_3031,N_2802,N_2027);
xor U3032 (N_3032,N_2543,N_2830);
and U3033 (N_3033,N_1710,N_2844);
xnor U3034 (N_3034,N_1957,N_2238);
nor U3035 (N_3035,N_2548,N_2571);
nand U3036 (N_3036,N_2500,N_1663);
or U3037 (N_3037,N_1697,N_2977);
nand U3038 (N_3038,N_2785,N_2212);
nand U3039 (N_3039,N_2247,N_1611);
nand U3040 (N_3040,N_2030,N_1782);
and U3041 (N_3041,N_2921,N_2308);
and U3042 (N_3042,N_2783,N_2601);
nand U3043 (N_3043,N_2780,N_1578);
xor U3044 (N_3044,N_1938,N_2406);
nand U3045 (N_3045,N_2803,N_2503);
or U3046 (N_3046,N_1640,N_1933);
and U3047 (N_3047,N_2557,N_2814);
nand U3048 (N_3048,N_1529,N_1868);
nor U3049 (N_3049,N_2560,N_2019);
nand U3050 (N_3050,N_2271,N_2322);
xor U3051 (N_3051,N_1901,N_2301);
or U3052 (N_3052,N_2400,N_2946);
xnor U3053 (N_3053,N_2729,N_2436);
or U3054 (N_3054,N_1527,N_1955);
nor U3055 (N_3055,N_2453,N_2750);
nor U3056 (N_3056,N_1582,N_1817);
xnor U3057 (N_3057,N_2736,N_1983);
xnor U3058 (N_3058,N_1752,N_1794);
nor U3059 (N_3059,N_2887,N_2664);
nor U3060 (N_3060,N_2576,N_1732);
or U3061 (N_3061,N_2579,N_2330);
xor U3062 (N_3062,N_2165,N_1535);
or U3063 (N_3063,N_2602,N_2687);
xnor U3064 (N_3064,N_1992,N_1678);
nor U3065 (N_3065,N_1515,N_2422);
and U3066 (N_3066,N_2537,N_1783);
nor U3067 (N_3067,N_1759,N_1709);
or U3068 (N_3068,N_2032,N_2950);
nor U3069 (N_3069,N_2339,N_2376);
nor U3070 (N_3070,N_2264,N_1606);
nand U3071 (N_3071,N_1597,N_2819);
or U3072 (N_3072,N_2539,N_2311);
nand U3073 (N_3073,N_2163,N_2631);
and U3074 (N_3074,N_1716,N_1665);
and U3075 (N_3075,N_2789,N_2833);
nor U3076 (N_3076,N_2935,N_2892);
nand U3077 (N_3077,N_2269,N_1895);
nand U3078 (N_3078,N_2829,N_2774);
nor U3079 (N_3079,N_1959,N_1613);
xnor U3080 (N_3080,N_2545,N_2765);
nand U3081 (N_3081,N_1674,N_1791);
or U3082 (N_3082,N_2943,N_1614);
or U3083 (N_3083,N_2440,N_2512);
and U3084 (N_3084,N_2359,N_2242);
or U3085 (N_3085,N_1830,N_1687);
nor U3086 (N_3086,N_2431,N_1666);
nand U3087 (N_3087,N_1949,N_1812);
or U3088 (N_3088,N_1680,N_2104);
or U3089 (N_3089,N_1656,N_1650);
and U3090 (N_3090,N_2712,N_1811);
xnor U3091 (N_3091,N_2689,N_1878);
or U3092 (N_3092,N_1774,N_1702);
nand U3093 (N_3093,N_2906,N_2270);
and U3094 (N_3094,N_2160,N_2197);
or U3095 (N_3095,N_1536,N_1815);
and U3096 (N_3096,N_2605,N_2798);
or U3097 (N_3097,N_2639,N_2928);
nand U3098 (N_3098,N_2973,N_2591);
or U3099 (N_3099,N_1882,N_1814);
and U3100 (N_3100,N_1564,N_2129);
xor U3101 (N_3101,N_2262,N_2984);
nor U3102 (N_3102,N_2228,N_1738);
or U3103 (N_3103,N_1690,N_2751);
nand U3104 (N_3104,N_1907,N_2583);
nand U3105 (N_3105,N_2904,N_2296);
nand U3106 (N_3106,N_2219,N_2580);
or U3107 (N_3107,N_1575,N_2684);
nor U3108 (N_3108,N_2233,N_1556);
and U3109 (N_3109,N_1841,N_2227);
xnor U3110 (N_3110,N_2794,N_2075);
nand U3111 (N_3111,N_1744,N_2413);
nor U3112 (N_3112,N_1728,N_2283);
nand U3113 (N_3113,N_2052,N_2125);
nand U3114 (N_3114,N_2320,N_2425);
nand U3115 (N_3115,N_1864,N_1906);
xor U3116 (N_3116,N_1638,N_2334);
nand U3117 (N_3117,N_1605,N_2788);
or U3118 (N_3118,N_1908,N_1623);
and U3119 (N_3119,N_2292,N_1813);
xor U3120 (N_3120,N_1528,N_2378);
nand U3121 (N_3121,N_2225,N_2737);
xnor U3122 (N_3122,N_1544,N_1632);
or U3123 (N_3123,N_2725,N_1828);
nor U3124 (N_3124,N_2498,N_2641);
nor U3125 (N_3125,N_2114,N_2151);
nand U3126 (N_3126,N_1988,N_2649);
nand U3127 (N_3127,N_1934,N_2969);
and U3128 (N_3128,N_2693,N_2380);
and U3129 (N_3129,N_2587,N_2620);
nand U3130 (N_3130,N_1979,N_2743);
or U3131 (N_3131,N_1795,N_1917);
nand U3132 (N_3132,N_1560,N_2009);
and U3133 (N_3133,N_1712,N_2593);
nand U3134 (N_3134,N_2069,N_2879);
nand U3135 (N_3135,N_2006,N_2700);
and U3136 (N_3136,N_1987,N_2575);
xor U3137 (N_3137,N_1966,N_1720);
xor U3138 (N_3138,N_2618,N_2561);
nor U3139 (N_3139,N_2170,N_1977);
xnor U3140 (N_3140,N_2056,N_2880);
or U3141 (N_3141,N_2975,N_2230);
or U3142 (N_3142,N_2517,N_2171);
xor U3143 (N_3143,N_1576,N_1771);
nor U3144 (N_3144,N_2885,N_2874);
and U3145 (N_3145,N_1888,N_2505);
and U3146 (N_3146,N_1603,N_1944);
and U3147 (N_3147,N_2848,N_2218);
nor U3148 (N_3148,N_2065,N_2187);
nor U3149 (N_3149,N_2377,N_2385);
nand U3150 (N_3150,N_1773,N_1809);
nand U3151 (N_3151,N_2179,N_2024);
and U3152 (N_3152,N_2724,N_2572);
nand U3153 (N_3153,N_2913,N_2749);
nand U3154 (N_3154,N_2760,N_2023);
nand U3155 (N_3155,N_2988,N_2925);
nand U3156 (N_3156,N_1974,N_2471);
nand U3157 (N_3157,N_1634,N_2932);
and U3158 (N_3158,N_2746,N_2507);
nor U3159 (N_3159,N_1790,N_1775);
nor U3160 (N_3160,N_2529,N_1677);
or U3161 (N_3161,N_2592,N_2619);
nor U3162 (N_3162,N_1572,N_2614);
and U3163 (N_3163,N_1985,N_2540);
and U3164 (N_3164,N_2578,N_1676);
nor U3165 (N_3165,N_1598,N_2168);
or U3166 (N_3166,N_2083,N_2799);
nand U3167 (N_3167,N_2328,N_2265);
nand U3168 (N_3168,N_2192,N_2551);
nor U3169 (N_3169,N_2980,N_2237);
nand U3170 (N_3170,N_1785,N_2295);
nor U3171 (N_3171,N_2859,N_2304);
nand U3172 (N_3172,N_2889,N_1570);
nand U3173 (N_3173,N_1784,N_2544);
nor U3174 (N_3174,N_1952,N_2966);
or U3175 (N_3175,N_1918,N_1857);
nand U3176 (N_3176,N_1804,N_1727);
xnor U3177 (N_3177,N_1519,N_2184);
nand U3178 (N_3178,N_2753,N_2041);
nor U3179 (N_3179,N_2057,N_2787);
or U3180 (N_3180,N_2142,N_1793);
nand U3181 (N_3181,N_1796,N_2342);
or U3182 (N_3182,N_1671,N_2843);
xor U3183 (N_3183,N_1645,N_2156);
nor U3184 (N_3184,N_1557,N_1559);
and U3185 (N_3185,N_2839,N_2538);
nor U3186 (N_3186,N_2632,N_1890);
nor U3187 (N_3187,N_2348,N_2448);
nor U3188 (N_3188,N_2995,N_2635);
xnor U3189 (N_3189,N_2643,N_1926);
or U3190 (N_3190,N_2351,N_2407);
nor U3191 (N_3191,N_2389,N_2483);
or U3192 (N_3192,N_2094,N_1546);
nand U3193 (N_3193,N_2827,N_2430);
nand U3194 (N_3194,N_1574,N_1743);
xor U3195 (N_3195,N_2797,N_2079);
nand U3196 (N_3196,N_2349,N_2589);
and U3197 (N_3197,N_2919,N_1799);
and U3198 (N_3198,N_2445,N_2564);
nand U3199 (N_3199,N_1975,N_2258);
nor U3200 (N_3200,N_2717,N_2982);
and U3201 (N_3201,N_1670,N_2807);
and U3202 (N_3202,N_2902,N_2586);
nand U3203 (N_3203,N_2994,N_2541);
and U3204 (N_3204,N_1887,N_1824);
xor U3205 (N_3205,N_1989,N_1635);
nor U3206 (N_3206,N_2944,N_2464);
nand U3207 (N_3207,N_1545,N_2871);
and U3208 (N_3208,N_1805,N_2515);
xnor U3209 (N_3209,N_2420,N_2465);
nor U3210 (N_3210,N_2112,N_2741);
or U3211 (N_3211,N_2432,N_1507);
xnor U3212 (N_3212,N_2996,N_1835);
xnor U3213 (N_3213,N_2818,N_2903);
xor U3214 (N_3214,N_2985,N_2408);
and U3215 (N_3215,N_2419,N_2852);
or U3216 (N_3216,N_2735,N_1921);
nand U3217 (N_3217,N_2384,N_2460);
or U3218 (N_3218,N_2499,N_2983);
and U3219 (N_3219,N_2690,N_1972);
or U3220 (N_3220,N_1912,N_2223);
or U3221 (N_3221,N_2143,N_1763);
nand U3222 (N_3222,N_1748,N_2938);
xnor U3223 (N_3223,N_1865,N_2274);
xor U3224 (N_3224,N_1755,N_1596);
xnor U3225 (N_3225,N_1767,N_2372);
and U3226 (N_3226,N_1655,N_2477);
nor U3227 (N_3227,N_2681,N_2688);
nand U3228 (N_3228,N_1558,N_2714);
and U3229 (N_3229,N_2409,N_1642);
xnor U3230 (N_3230,N_2533,N_2546);
or U3231 (N_3231,N_2744,N_1504);
and U3232 (N_3232,N_1846,N_2675);
xnor U3233 (N_3233,N_1797,N_1896);
or U3234 (N_3234,N_1965,N_2180);
nor U3235 (N_3235,N_1539,N_2934);
nand U3236 (N_3236,N_2155,N_2411);
nand U3237 (N_3237,N_2327,N_2709);
and U3238 (N_3238,N_1583,N_2971);
xnor U3239 (N_3239,N_2888,N_2922);
nand U3240 (N_3240,N_2534,N_2044);
xor U3241 (N_3241,N_2017,N_2895);
nor U3242 (N_3242,N_2671,N_1914);
nor U3243 (N_3243,N_2495,N_2117);
or U3244 (N_3244,N_1701,N_2275);
xor U3245 (N_3245,N_1874,N_2532);
nand U3246 (N_3246,N_2086,N_2647);
nor U3247 (N_3247,N_2915,N_2720);
and U3248 (N_3248,N_1885,N_2651);
and U3249 (N_3249,N_1567,N_2357);
nor U3250 (N_3250,N_2177,N_2704);
xor U3251 (N_3251,N_1600,N_2205);
or U3252 (N_3252,N_1842,N_2289);
nor U3253 (N_3253,N_1737,N_2949);
nand U3254 (N_3254,N_2116,N_1731);
nor U3255 (N_3255,N_2842,N_2722);
or U3256 (N_3256,N_2584,N_2273);
xnor U3257 (N_3257,N_2255,N_2627);
nor U3258 (N_3258,N_1923,N_1810);
nand U3259 (N_3259,N_2567,N_1963);
and U3260 (N_3260,N_1725,N_2049);
nor U3261 (N_3261,N_1682,N_2084);
nor U3262 (N_3262,N_1644,N_1729);
and U3263 (N_3263,N_2345,N_2896);
nand U3264 (N_3264,N_2174,N_2183);
and U3265 (N_3265,N_2653,N_1561);
or U3266 (N_3266,N_2779,N_2752);
or U3267 (N_3267,N_2046,N_1595);
and U3268 (N_3268,N_2513,N_1501);
or U3269 (N_3269,N_2390,N_2778);
xnor U3270 (N_3270,N_2417,N_1563);
and U3271 (N_3271,N_1747,N_2695);
and U3272 (N_3272,N_2793,N_2553);
nand U3273 (N_3273,N_1831,N_2241);
and U3274 (N_3274,N_1750,N_2637);
xnor U3275 (N_3275,N_2253,N_2563);
or U3276 (N_3276,N_2415,N_2707);
or U3277 (N_3277,N_1510,N_2519);
and U3278 (N_3278,N_2037,N_2826);
nand U3279 (N_3279,N_1786,N_1643);
and U3280 (N_3280,N_2759,N_2692);
nand U3281 (N_3281,N_2881,N_2491);
and U3282 (N_3282,N_2761,N_2625);
nor U3283 (N_3283,N_1986,N_2756);
xnor U3284 (N_3284,N_2866,N_2468);
xnor U3285 (N_3285,N_2455,N_2111);
nor U3286 (N_3286,N_1803,N_1998);
xnor U3287 (N_3287,N_2993,N_1898);
nor U3288 (N_3288,N_1788,N_2611);
xor U3289 (N_3289,N_2703,N_1537);
xnor U3290 (N_3290,N_2410,N_1970);
nand U3291 (N_3291,N_2118,N_1509);
nand U3292 (N_3292,N_2680,N_1819);
xor U3293 (N_3293,N_1776,N_2062);
nor U3294 (N_3294,N_2276,N_2438);
nand U3295 (N_3295,N_1897,N_2352);
nand U3296 (N_3296,N_1617,N_1736);
xor U3297 (N_3297,N_2970,N_2747);
nor U3298 (N_3298,N_1685,N_2321);
nand U3299 (N_3299,N_1647,N_2492);
xor U3300 (N_3300,N_2297,N_1982);
or U3301 (N_3301,N_2890,N_2356);
nand U3302 (N_3302,N_1821,N_2683);
nor U3303 (N_3303,N_2482,N_1581);
nor U3304 (N_3304,N_2502,N_1689);
xnor U3305 (N_3305,N_2421,N_1672);
nor U3306 (N_3306,N_2490,N_2951);
xor U3307 (N_3307,N_2362,N_1948);
xor U3308 (N_3308,N_1592,N_2877);
xor U3309 (N_3309,N_2375,N_2437);
nor U3310 (N_3310,N_2530,N_2060);
xor U3311 (N_3311,N_2795,N_2216);
nand U3312 (N_3312,N_1555,N_2691);
xor U3313 (N_3313,N_2260,N_1858);
and U3314 (N_3314,N_1884,N_2344);
and U3315 (N_3315,N_2066,N_2485);
or U3316 (N_3316,N_2077,N_1861);
xnor U3317 (N_3317,N_2621,N_2150);
or U3318 (N_3318,N_1849,N_2284);
xor U3319 (N_3319,N_2672,N_2382);
nor U3320 (N_3320,N_2825,N_2261);
and U3321 (N_3321,N_1902,N_1836);
nand U3322 (N_3322,N_1745,N_2721);
xnor U3323 (N_3323,N_2828,N_2130);
xor U3324 (N_3324,N_2068,N_2252);
xor U3325 (N_3325,N_2035,N_1706);
and U3326 (N_3326,N_2521,N_2686);
xnor U3327 (N_3327,N_1657,N_2815);
or U3328 (N_3328,N_1713,N_2633);
xnor U3329 (N_3329,N_2955,N_2059);
nor U3330 (N_3330,N_2609,N_2070);
and U3331 (N_3331,N_2392,N_2329);
or U3332 (N_3332,N_2291,N_2207);
xor U3333 (N_3333,N_2463,N_2098);
nor U3334 (N_3334,N_1700,N_2767);
or U3335 (N_3335,N_1855,N_2758);
or U3336 (N_3336,N_2162,N_2923);
xnor U3337 (N_3337,N_2064,N_2245);
xnor U3338 (N_3338,N_2981,N_1827);
nand U3339 (N_3339,N_2208,N_2314);
nor U3340 (N_3340,N_2333,N_1826);
or U3341 (N_3341,N_2257,N_1721);
nand U3342 (N_3342,N_2189,N_2350);
nand U3343 (N_3343,N_1844,N_2909);
nand U3344 (N_3344,N_1754,N_2542);
or U3345 (N_3345,N_2535,N_1969);
nand U3346 (N_3346,N_1869,N_1723);
nand U3347 (N_3347,N_2764,N_1847);
or U3348 (N_3348,N_2757,N_2121);
nand U3349 (N_3349,N_2835,N_1512);
nand U3350 (N_3350,N_1540,N_1549);
nor U3351 (N_3351,N_2677,N_2791);
or U3352 (N_3352,N_2528,N_2157);
and U3353 (N_3353,N_2401,N_2845);
and U3354 (N_3354,N_2036,N_2702);
and U3355 (N_3355,N_2234,N_2206);
or U3356 (N_3356,N_2361,N_2034);
xor U3357 (N_3357,N_1571,N_2812);
and U3358 (N_3358,N_1514,N_2525);
or U3359 (N_3359,N_2976,N_2918);
and U3360 (N_3360,N_2958,N_1692);
xor U3361 (N_3361,N_2608,N_2987);
nor U3362 (N_3362,N_2929,N_2685);
xor U3363 (N_3363,N_2414,N_2095);
or U3364 (N_3364,N_1553,N_2149);
xnor U3365 (N_3365,N_2148,N_1649);
nand U3366 (N_3366,N_2014,N_2857);
or U3367 (N_3367,N_2011,N_2912);
nor U3368 (N_3368,N_2371,N_2232);
nand U3369 (N_3369,N_1719,N_1881);
and U3370 (N_3370,N_2310,N_1542);
and U3371 (N_3371,N_1863,N_2577);
and U3372 (N_3372,N_1990,N_2486);
and U3373 (N_3373,N_2924,N_1845);
nor U3374 (N_3374,N_2048,N_1802);
or U3375 (N_3375,N_1552,N_2884);
nor U3376 (N_3376,N_1981,N_2235);
and U3377 (N_3377,N_2475,N_1941);
or U3378 (N_3378,N_2710,N_1705);
xor U3379 (N_3379,N_2734,N_1746);
and U3380 (N_3380,N_1954,N_2008);
nor U3381 (N_3381,N_2222,N_2078);
nor U3382 (N_3382,N_2256,N_2948);
or U3383 (N_3383,N_2474,N_1859);
and U3384 (N_3384,N_2085,N_2947);
or U3385 (N_3385,N_1653,N_1502);
or U3386 (N_3386,N_2606,N_2434);
and U3387 (N_3387,N_1800,N_2341);
xnor U3388 (N_3388,N_2454,N_1765);
and U3389 (N_3389,N_2711,N_1661);
nand U3390 (N_3390,N_2193,N_2309);
xnor U3391 (N_3391,N_1769,N_2555);
or U3392 (N_3392,N_1924,N_2399);
nand U3393 (N_3393,N_2667,N_1843);
nand U3394 (N_3394,N_1628,N_1761);
xor U3395 (N_3395,N_2840,N_2901);
and U3396 (N_3396,N_2875,N_1506);
nor U3397 (N_3397,N_1652,N_2426);
xor U3398 (N_3398,N_2642,N_2053);
or U3399 (N_3399,N_2387,N_1703);
nor U3400 (N_3400,N_1931,N_1991);
xnor U3401 (N_3401,N_2010,N_1792);
xor U3402 (N_3402,N_2347,N_1978);
nor U3403 (N_3403,N_1742,N_2898);
or U3404 (N_3404,N_1871,N_1967);
or U3405 (N_3405,N_1594,N_2940);
or U3406 (N_3406,N_1900,N_1704);
or U3407 (N_3407,N_2682,N_2279);
and U3408 (N_3408,N_1928,N_2792);
and U3409 (N_3409,N_1850,N_2395);
nor U3410 (N_3410,N_1733,N_1633);
and U3411 (N_3411,N_2199,N_2221);
nand U3412 (N_3412,N_2461,N_2713);
nor U3413 (N_3413,N_2665,N_2698);
or U3414 (N_3414,N_1911,N_2652);
and U3415 (N_3415,N_2668,N_1590);
and U3416 (N_3416,N_2003,N_2141);
xor U3417 (N_3417,N_2092,N_2801);
xor U3418 (N_3418,N_2806,N_1621);
or U3419 (N_3419,N_1735,N_2278);
nor U3420 (N_3420,N_2191,N_2634);
or U3421 (N_3421,N_2282,N_2705);
nand U3422 (N_3422,N_1772,N_1660);
nand U3423 (N_3423,N_1533,N_2883);
xnor U3424 (N_3424,N_1930,N_2914);
and U3425 (N_3425,N_2145,N_1531);
or U3426 (N_3426,N_2820,N_2600);
nand U3427 (N_3427,N_1518,N_2998);
nor U3428 (N_3428,N_2340,N_2974);
or U3429 (N_3429,N_2231,N_2088);
and U3430 (N_3430,N_1698,N_2804);
or U3431 (N_3431,N_2550,N_2559);
or U3432 (N_3432,N_1852,N_1943);
or U3433 (N_3433,N_1739,N_2963);
or U3434 (N_3434,N_1520,N_1892);
nor U3435 (N_3435,N_2654,N_2091);
and U3436 (N_3436,N_2786,N_2501);
nand U3437 (N_3437,N_2398,N_2942);
xor U3438 (N_3438,N_2190,N_1568);
and U3439 (N_3439,N_2864,N_1929);
nand U3440 (N_3440,N_1953,N_2766);
or U3441 (N_3441,N_1688,N_1886);
nor U3442 (N_3442,N_2040,N_2451);
xor U3443 (N_3443,N_1751,N_2851);
or U3444 (N_3444,N_2834,N_2109);
nand U3445 (N_3445,N_2217,N_2917);
nand U3446 (N_3446,N_1673,N_2748);
or U3447 (N_3447,N_2536,N_2450);
xnor U3448 (N_3448,N_1950,N_2569);
or U3449 (N_3449,N_2416,N_2813);
and U3450 (N_3450,N_1904,N_2841);
nor U3451 (N_3451,N_2402,N_1734);
xnor U3452 (N_3452,N_2324,N_2293);
nand U3453 (N_3453,N_2336,N_2126);
nor U3454 (N_3454,N_2370,N_2161);
and U3455 (N_3455,N_2640,N_2090);
nand U3456 (N_3456,N_2096,N_2388);
and U3457 (N_3457,N_2452,N_2441);
nor U3458 (N_3458,N_1976,N_1875);
or U3459 (N_3459,N_2369,N_2038);
or U3460 (N_3460,N_2101,N_1508);
and U3461 (N_3461,N_2277,N_2131);
or U3462 (N_3462,N_1889,N_2166);
or U3463 (N_3463,N_2099,N_2524);
nor U3464 (N_3464,N_2220,N_1958);
or U3465 (N_3465,N_1551,N_2479);
nand U3466 (N_3466,N_2715,N_2067);
nor U3467 (N_3467,N_1741,N_1758);
nand U3468 (N_3468,N_2733,N_2429);
or U3469 (N_3469,N_2823,N_2167);
nand U3470 (N_3470,N_2210,N_2047);
xnor U3471 (N_3471,N_1883,N_1956);
and U3472 (N_3472,N_1625,N_1711);
and U3473 (N_3473,N_1580,N_2972);
nor U3474 (N_3474,N_2021,N_2323);
xnor U3475 (N_3475,N_2655,N_2176);
xor U3476 (N_3476,N_2063,N_2960);
nor U3477 (N_3477,N_1837,N_2527);
nand U3478 (N_3478,N_1717,N_2473);
nor U3479 (N_3479,N_2585,N_2186);
or U3480 (N_3480,N_2716,N_2072);
nor U3481 (N_3481,N_1616,N_1683);
or U3482 (N_3482,N_2624,N_1608);
or U3483 (N_3483,N_1562,N_1740);
or U3484 (N_3484,N_2518,N_2185);
and U3485 (N_3485,N_2144,N_1664);
or U3486 (N_3486,N_2281,N_1853);
xnor U3487 (N_3487,N_2080,N_2817);
xor U3488 (N_3488,N_2316,N_2740);
nand U3489 (N_3489,N_2623,N_1694);
xnor U3490 (N_3490,N_2042,N_1936);
and U3491 (N_3491,N_2300,N_1915);
xor U3492 (N_3492,N_2202,N_2383);
and U3493 (N_3493,N_2514,N_2248);
nand U3494 (N_3494,N_1577,N_1646);
or U3495 (N_3495,N_1829,N_2058);
and U3496 (N_3496,N_2458,N_1654);
xor U3497 (N_3497,N_1648,N_2566);
and U3498 (N_3498,N_2449,N_2005);
xnor U3499 (N_3499,N_2622,N_2679);
and U3500 (N_3500,N_1543,N_2462);
xor U3501 (N_3501,N_2226,N_2119);
xor U3502 (N_3502,N_1964,N_1962);
or U3503 (N_3503,N_2650,N_2355);
nor U3504 (N_3504,N_2522,N_2952);
nand U3505 (N_3505,N_2873,N_1610);
xor U3506 (N_3506,N_2404,N_1780);
and U3507 (N_3507,N_2343,N_2381);
nor U3508 (N_3508,N_2732,N_2554);
nand U3509 (N_3509,N_2775,N_1708);
nand U3510 (N_3510,N_2872,N_2487);
nand U3511 (N_3511,N_1764,N_2082);
or U3512 (N_3512,N_1870,N_1505);
or U3513 (N_3513,N_1996,N_1532);
nand U3514 (N_3514,N_1566,N_2338);
or U3515 (N_3515,N_2894,N_2978);
and U3516 (N_3516,N_2424,N_2133);
or U3517 (N_3517,N_1781,N_2626);
nand U3518 (N_3518,N_2120,N_2224);
nand U3519 (N_3519,N_2968,N_1730);
nand U3520 (N_3520,N_2876,N_2412);
xnor U3521 (N_3521,N_1631,N_1669);
nand U3522 (N_3522,N_2882,N_2821);
xnor U3523 (N_3523,N_1820,N_1624);
or U3524 (N_3524,N_2396,N_1807);
nand U3525 (N_3525,N_2865,N_2905);
or U3526 (N_3526,N_2140,N_2648);
or U3527 (N_3527,N_2661,N_2597);
nand U3528 (N_3528,N_2358,N_2360);
and U3529 (N_3529,N_1760,N_1808);
and U3530 (N_3530,N_1867,N_2433);
nand U3531 (N_3531,N_1547,N_1838);
nor U3532 (N_3532,N_2790,N_2497);
xnor U3533 (N_3533,N_2718,N_1960);
and U3534 (N_3534,N_1801,N_2916);
nand U3535 (N_3535,N_1839,N_2102);
or U3536 (N_3536,N_2105,N_2159);
xnor U3537 (N_3537,N_2706,N_2154);
xor U3538 (N_3538,N_2754,N_2599);
nand U3539 (N_3539,N_2470,N_2367);
or U3540 (N_3540,N_1840,N_1925);
or U3541 (N_3541,N_2081,N_2956);
xnor U3542 (N_3542,N_2020,N_2669);
or U3543 (N_3543,N_2570,N_2093);
nand U3544 (N_3544,N_1517,N_1968);
or U3545 (N_3545,N_2000,N_2195);
nor U3546 (N_3546,N_1856,N_2900);
nand U3547 (N_3547,N_2480,N_2676);
nor U3548 (N_3548,N_1879,N_1905);
and U3549 (N_3549,N_2239,N_2444);
and U3550 (N_3550,N_2893,N_2181);
nor U3551 (N_3551,N_2824,N_2172);
or U3552 (N_3552,N_2055,N_2565);
nand U3553 (N_3553,N_1591,N_2574);
xor U3554 (N_3554,N_2251,N_2051);
or U3555 (N_3555,N_2097,N_1935);
or U3556 (N_3556,N_1651,N_2478);
nand U3557 (N_3557,N_2073,N_2742);
nand U3558 (N_3558,N_2613,N_2930);
xor U3559 (N_3559,N_1607,N_2418);
and U3560 (N_3560,N_2856,N_2506);
xor U3561 (N_3561,N_2287,N_1932);
or U3562 (N_3562,N_2365,N_2229);
nand U3563 (N_3563,N_2697,N_1973);
xnor U3564 (N_3564,N_2018,N_2674);
xor U3565 (N_3565,N_2110,N_1526);
or U3566 (N_3566,N_2332,N_2999);
and U3567 (N_3567,N_2805,N_1541);
or U3568 (N_3568,N_2701,N_1615);
nor U3569 (N_3569,N_2158,N_2954);
and U3570 (N_3570,N_2869,N_1550);
and U3571 (N_3571,N_2331,N_2776);
nand U3572 (N_3572,N_2493,N_1872);
xor U3573 (N_3573,N_2456,N_2488);
nor U3574 (N_3574,N_1726,N_1548);
or U3575 (N_3575,N_1641,N_2259);
nor U3576 (N_3576,N_2953,N_2313);
or U3577 (N_3577,N_1880,N_1753);
nor U3578 (N_3578,N_2466,N_2076);
and U3579 (N_3579,N_2861,N_2594);
and U3580 (N_3580,N_1994,N_2670);
nor U3581 (N_3581,N_2045,N_2965);
and U3582 (N_3582,N_2484,N_2598);
or U3583 (N_3583,N_2832,N_2727);
and U3584 (N_3584,N_2562,N_2152);
nand U3585 (N_3585,N_1916,N_2907);
nor U3586 (N_3586,N_2730,N_1834);
nand U3587 (N_3587,N_2739,N_1601);
or U3588 (N_3588,N_1693,N_1691);
nand U3589 (N_3589,N_1612,N_2368);
nand U3590 (N_3590,N_2317,N_2122);
and U3591 (N_3591,N_2403,N_2610);
nand U3592 (N_3592,N_2405,N_2394);
and U3593 (N_3593,N_2363,N_2773);
xnor U3594 (N_3594,N_2768,N_2428);
and U3595 (N_3595,N_2215,N_2628);
nand U3596 (N_3596,N_2243,N_1584);
nand U3597 (N_3597,N_2013,N_1516);
or U3598 (N_3598,N_2645,N_2558);
and U3599 (N_3599,N_2364,N_2607);
or U3600 (N_3600,N_2115,N_2457);
xor U3601 (N_3601,N_2992,N_2026);
or U3602 (N_3602,N_1920,N_2442);
nand U3603 (N_3603,N_1876,N_2374);
nand U3604 (N_3604,N_1626,N_1818);
nor U3605 (N_3605,N_2809,N_1714);
and U3606 (N_3606,N_2427,N_2811);
and U3607 (N_3607,N_2822,N_2781);
and U3608 (N_3608,N_2028,N_2123);
xor U3609 (N_3609,N_2173,N_1762);
and U3610 (N_3610,N_2615,N_1715);
nand U3611 (N_3611,N_2927,N_1848);
nor U3612 (N_3612,N_1588,N_1530);
xnor U3613 (N_3613,N_2153,N_1816);
nor U3614 (N_3614,N_2128,N_1525);
nand U3615 (N_3615,N_1961,N_2087);
nand U3616 (N_3616,N_2846,N_1585);
xor U3617 (N_3617,N_2007,N_2211);
nor U3618 (N_3618,N_2213,N_1945);
xor U3619 (N_3619,N_2784,N_1825);
and U3620 (N_3620,N_2556,N_1637);
or U3621 (N_3621,N_1513,N_2868);
nor U3622 (N_3622,N_2657,N_1718);
nand U3623 (N_3623,N_1604,N_2728);
nor U3624 (N_3624,N_1778,N_2188);
nor U3625 (N_3625,N_1696,N_1787);
and U3626 (N_3626,N_2581,N_2616);
or U3627 (N_3627,N_2312,N_1662);
and U3628 (N_3628,N_2860,N_2867);
xor U3629 (N_3629,N_1903,N_2986);
nor U3630 (N_3630,N_1891,N_1899);
xor U3631 (N_3631,N_2459,N_1951);
or U3632 (N_3632,N_2772,N_2658);
xor U3633 (N_3633,N_2796,N_2016);
nand U3634 (N_3634,N_2134,N_1854);
nand U3635 (N_3635,N_2878,N_1627);
nand U3636 (N_3636,N_2236,N_2054);
or U3637 (N_3637,N_2476,N_2182);
xnor U3638 (N_3638,N_2299,N_1681);
and U3639 (N_3639,N_1822,N_2039);
nor U3640 (N_3640,N_2200,N_2196);
nor U3641 (N_3641,N_2810,N_2294);
nor U3642 (N_3642,N_2699,N_1573);
xnor U3643 (N_3643,N_1602,N_1980);
nor U3644 (N_3644,N_1993,N_1579);
and U3645 (N_3645,N_2990,N_2214);
nor U3646 (N_3646,N_2435,N_2302);
or U3647 (N_3647,N_2175,N_2708);
or U3648 (N_3648,N_2286,N_1699);
nor U3649 (N_3649,N_2132,N_1823);
nor U3650 (N_3650,N_2656,N_2050);
xnor U3651 (N_3651,N_2002,N_2523);
nor U3652 (N_3652,N_1833,N_2891);
and U3653 (N_3653,N_1756,N_2031);
xor U3654 (N_3654,N_2573,N_2127);
and U3655 (N_3655,N_2280,N_2508);
nor U3656 (N_3656,N_1593,N_2603);
nand U3657 (N_3657,N_2962,N_1707);
nand U3658 (N_3658,N_2549,N_2520);
xnor U3659 (N_3659,N_1534,N_2552);
or U3660 (N_3660,N_2638,N_2137);
nor U3661 (N_3661,N_2004,N_2346);
nor U3662 (N_3662,N_1866,N_2926);
xor U3663 (N_3663,N_2379,N_1724);
or U3664 (N_3664,N_2831,N_1909);
or U3665 (N_3665,N_2636,N_2911);
or U3666 (N_3666,N_2298,N_1860);
xnor U3667 (N_3667,N_2673,N_2254);
or U3668 (N_3668,N_1589,N_2853);
nor U3669 (N_3669,N_1511,N_2897);
nand U3670 (N_3670,N_2510,N_1686);
xnor U3671 (N_3671,N_2246,N_1538);
or U3672 (N_3672,N_1766,N_1893);
nand U3673 (N_3673,N_2146,N_2147);
nand U3674 (N_3674,N_1806,N_2800);
and U3675 (N_3675,N_2719,N_2439);
nand U3676 (N_3676,N_2854,N_2194);
xor U3677 (N_3677,N_2373,N_1618);
or U3678 (N_3678,N_2354,N_2731);
nand U3679 (N_3679,N_2991,N_2862);
and U3680 (N_3680,N_2777,N_1894);
nand U3681 (N_3681,N_2755,N_2136);
xor U3682 (N_3682,N_2849,N_2659);
xor U3683 (N_3683,N_1927,N_1999);
or U3684 (N_3684,N_1586,N_2481);
xor U3685 (N_3685,N_2666,N_2723);
xor U3686 (N_3686,N_1768,N_2107);
and U3687 (N_3687,N_2660,N_1521);
nor U3688 (N_3688,N_2646,N_2696);
nand U3689 (N_3689,N_2694,N_2726);
or U3690 (N_3690,N_2113,N_2198);
xnor U3691 (N_3691,N_2201,N_2288);
and U3692 (N_3692,N_1523,N_2489);
and U3693 (N_3693,N_2446,N_1913);
or U3694 (N_3694,N_1684,N_2074);
and U3695 (N_3695,N_2836,N_2588);
or U3696 (N_3696,N_2391,N_1922);
xor U3697 (N_3697,N_2855,N_2366);
nor U3698 (N_3698,N_1779,N_2678);
xnor U3699 (N_3699,N_1997,N_2494);
nor U3700 (N_3700,N_2931,N_1984);
nand U3701 (N_3701,N_2847,N_2025);
nor U3702 (N_3702,N_1636,N_2100);
nand U3703 (N_3703,N_2961,N_2989);
nor U3704 (N_3704,N_2933,N_2033);
xnor U3705 (N_3705,N_2979,N_2910);
nor U3706 (N_3706,N_1659,N_2303);
xnor U3707 (N_3707,N_1675,N_2939);
and U3708 (N_3708,N_1770,N_2644);
and U3709 (N_3709,N_2590,N_2272);
or U3710 (N_3710,N_2945,N_2496);
and U3711 (N_3711,N_2568,N_1832);
or U3712 (N_3712,N_2863,N_1522);
nand U3713 (N_3713,N_2305,N_2762);
xor U3714 (N_3714,N_1940,N_2547);
nand U3715 (N_3715,N_2290,N_2263);
nor U3716 (N_3716,N_2967,N_1658);
nand U3717 (N_3717,N_2089,N_2209);
nand U3718 (N_3718,N_2103,N_2604);
or U3719 (N_3719,N_2837,N_2318);
xnor U3720 (N_3720,N_2582,N_2164);
and U3721 (N_3721,N_2769,N_2397);
nor U3722 (N_3722,N_2858,N_1524);
or U3723 (N_3723,N_1620,N_2782);
or U3724 (N_3724,N_2443,N_2531);
xor U3725 (N_3725,N_1789,N_2899);
xnor U3726 (N_3726,N_2808,N_2335);
nand U3727 (N_3727,N_2353,N_2467);
nand U3728 (N_3728,N_2250,N_2629);
nor U3729 (N_3729,N_2509,N_1667);
xor U3730 (N_3730,N_2249,N_2816);
and U3731 (N_3731,N_1995,N_2997);
nor U3732 (N_3732,N_1679,N_1609);
xor U3733 (N_3733,N_2447,N_2135);
or U3734 (N_3734,N_1946,N_1877);
nand U3735 (N_3735,N_2850,N_2204);
or U3736 (N_3736,N_2511,N_2936);
nand U3737 (N_3737,N_2662,N_1668);
and U3738 (N_3738,N_2838,N_2138);
and U3739 (N_3739,N_2029,N_1910);
nor U3740 (N_3740,N_2022,N_2061);
or U3741 (N_3741,N_2959,N_2941);
xor U3742 (N_3742,N_2244,N_1851);
or U3743 (N_3743,N_1873,N_2203);
or U3744 (N_3744,N_1619,N_2071);
or U3745 (N_3745,N_2964,N_1695);
nand U3746 (N_3746,N_2178,N_2908);
nand U3747 (N_3747,N_1503,N_2139);
xnor U3748 (N_3748,N_2306,N_2920);
nand U3749 (N_3749,N_1798,N_2617);
xor U3750 (N_3750,N_2063,N_1907);
nand U3751 (N_3751,N_2263,N_2640);
or U3752 (N_3752,N_2926,N_2440);
nor U3753 (N_3753,N_1548,N_1695);
nand U3754 (N_3754,N_1546,N_2851);
nand U3755 (N_3755,N_1953,N_2078);
and U3756 (N_3756,N_2314,N_2803);
or U3757 (N_3757,N_1684,N_2266);
nor U3758 (N_3758,N_2638,N_2513);
nand U3759 (N_3759,N_1645,N_2280);
nor U3760 (N_3760,N_2548,N_2551);
or U3761 (N_3761,N_2711,N_2845);
or U3762 (N_3762,N_1805,N_1579);
nor U3763 (N_3763,N_1966,N_2001);
nor U3764 (N_3764,N_1614,N_2461);
xnor U3765 (N_3765,N_1678,N_1851);
nand U3766 (N_3766,N_1506,N_2260);
nand U3767 (N_3767,N_2116,N_2625);
or U3768 (N_3768,N_1980,N_2039);
nand U3769 (N_3769,N_2466,N_2935);
and U3770 (N_3770,N_1717,N_2049);
and U3771 (N_3771,N_2805,N_2069);
or U3772 (N_3772,N_2961,N_2148);
or U3773 (N_3773,N_2526,N_2197);
xor U3774 (N_3774,N_1737,N_1559);
nor U3775 (N_3775,N_1603,N_2395);
nor U3776 (N_3776,N_2317,N_2183);
and U3777 (N_3777,N_1705,N_2667);
or U3778 (N_3778,N_2649,N_2127);
nand U3779 (N_3779,N_1584,N_2562);
or U3780 (N_3780,N_2008,N_2772);
xnor U3781 (N_3781,N_2695,N_2971);
and U3782 (N_3782,N_2021,N_2747);
nor U3783 (N_3783,N_2451,N_2566);
nand U3784 (N_3784,N_2025,N_2026);
and U3785 (N_3785,N_1895,N_2516);
nand U3786 (N_3786,N_2099,N_2933);
or U3787 (N_3787,N_2640,N_2335);
nor U3788 (N_3788,N_2660,N_2393);
nand U3789 (N_3789,N_1875,N_2699);
nand U3790 (N_3790,N_2137,N_2101);
and U3791 (N_3791,N_2061,N_2305);
xor U3792 (N_3792,N_2843,N_2370);
and U3793 (N_3793,N_2181,N_2574);
xnor U3794 (N_3794,N_1690,N_1800);
and U3795 (N_3795,N_2985,N_2219);
and U3796 (N_3796,N_1548,N_2194);
or U3797 (N_3797,N_2363,N_2264);
xor U3798 (N_3798,N_1900,N_1656);
or U3799 (N_3799,N_1624,N_2967);
nand U3800 (N_3800,N_2181,N_2495);
nand U3801 (N_3801,N_2425,N_1519);
xor U3802 (N_3802,N_2355,N_1627);
nand U3803 (N_3803,N_1917,N_2244);
nand U3804 (N_3804,N_2872,N_2049);
xnor U3805 (N_3805,N_2649,N_1666);
nor U3806 (N_3806,N_2872,N_1542);
and U3807 (N_3807,N_1853,N_1646);
or U3808 (N_3808,N_2702,N_2552);
nand U3809 (N_3809,N_1847,N_2701);
and U3810 (N_3810,N_2152,N_2983);
or U3811 (N_3811,N_2644,N_2746);
or U3812 (N_3812,N_2570,N_1693);
or U3813 (N_3813,N_2938,N_2449);
xor U3814 (N_3814,N_2630,N_2306);
nand U3815 (N_3815,N_2533,N_2760);
nand U3816 (N_3816,N_1756,N_2283);
or U3817 (N_3817,N_1762,N_2500);
nor U3818 (N_3818,N_2461,N_2009);
nor U3819 (N_3819,N_1874,N_1610);
or U3820 (N_3820,N_1686,N_1880);
nor U3821 (N_3821,N_1702,N_1913);
nand U3822 (N_3822,N_1806,N_2059);
nand U3823 (N_3823,N_1909,N_1680);
and U3824 (N_3824,N_2744,N_1830);
xnor U3825 (N_3825,N_2675,N_1930);
and U3826 (N_3826,N_2824,N_2056);
xor U3827 (N_3827,N_1739,N_1709);
xor U3828 (N_3828,N_2206,N_2212);
xnor U3829 (N_3829,N_2008,N_2259);
or U3830 (N_3830,N_2352,N_2230);
and U3831 (N_3831,N_2418,N_2245);
nand U3832 (N_3832,N_2967,N_2259);
xnor U3833 (N_3833,N_1933,N_1694);
or U3834 (N_3834,N_1670,N_1547);
nand U3835 (N_3835,N_1701,N_1861);
or U3836 (N_3836,N_2320,N_2932);
nor U3837 (N_3837,N_1524,N_2386);
and U3838 (N_3838,N_2013,N_1763);
nand U3839 (N_3839,N_2344,N_2737);
and U3840 (N_3840,N_2379,N_2469);
nor U3841 (N_3841,N_1921,N_1846);
xor U3842 (N_3842,N_2036,N_2965);
nor U3843 (N_3843,N_1880,N_2990);
nand U3844 (N_3844,N_1701,N_2247);
or U3845 (N_3845,N_2732,N_2961);
xor U3846 (N_3846,N_1674,N_2948);
and U3847 (N_3847,N_2422,N_1869);
nor U3848 (N_3848,N_2008,N_2050);
nor U3849 (N_3849,N_2847,N_2059);
and U3850 (N_3850,N_1751,N_2133);
xnor U3851 (N_3851,N_2820,N_1705);
and U3852 (N_3852,N_2057,N_2580);
xnor U3853 (N_3853,N_1645,N_1950);
nor U3854 (N_3854,N_2733,N_2835);
or U3855 (N_3855,N_2680,N_1685);
xor U3856 (N_3856,N_2037,N_2423);
nand U3857 (N_3857,N_2767,N_1656);
xnor U3858 (N_3858,N_1502,N_1730);
nor U3859 (N_3859,N_2072,N_2518);
xnor U3860 (N_3860,N_2641,N_1919);
xnor U3861 (N_3861,N_2713,N_2244);
nand U3862 (N_3862,N_1876,N_2594);
and U3863 (N_3863,N_2307,N_2478);
nand U3864 (N_3864,N_2509,N_2806);
xor U3865 (N_3865,N_2606,N_1669);
nand U3866 (N_3866,N_2532,N_2901);
nand U3867 (N_3867,N_2563,N_2160);
and U3868 (N_3868,N_2924,N_2899);
xor U3869 (N_3869,N_1933,N_2516);
xnor U3870 (N_3870,N_2927,N_1750);
xnor U3871 (N_3871,N_1647,N_2084);
nand U3872 (N_3872,N_2688,N_2731);
nand U3873 (N_3873,N_2813,N_1740);
nor U3874 (N_3874,N_1764,N_1900);
nand U3875 (N_3875,N_2782,N_2154);
xnor U3876 (N_3876,N_2291,N_2104);
nor U3877 (N_3877,N_1765,N_2681);
xor U3878 (N_3878,N_2208,N_1860);
nand U3879 (N_3879,N_1862,N_2433);
nor U3880 (N_3880,N_2850,N_1787);
nor U3881 (N_3881,N_2116,N_2173);
xor U3882 (N_3882,N_2985,N_1731);
nand U3883 (N_3883,N_2509,N_2482);
nor U3884 (N_3884,N_2215,N_2216);
nand U3885 (N_3885,N_2856,N_2014);
and U3886 (N_3886,N_2457,N_2110);
and U3887 (N_3887,N_2692,N_1825);
nand U3888 (N_3888,N_1592,N_2277);
nor U3889 (N_3889,N_2595,N_1756);
xnor U3890 (N_3890,N_2610,N_1614);
nor U3891 (N_3891,N_2223,N_1922);
nor U3892 (N_3892,N_2205,N_2549);
or U3893 (N_3893,N_2735,N_1528);
nand U3894 (N_3894,N_2518,N_1675);
nand U3895 (N_3895,N_1649,N_2270);
or U3896 (N_3896,N_2641,N_1679);
and U3897 (N_3897,N_1638,N_1799);
nor U3898 (N_3898,N_2912,N_2246);
nand U3899 (N_3899,N_2285,N_2839);
or U3900 (N_3900,N_2340,N_2470);
or U3901 (N_3901,N_2413,N_1819);
or U3902 (N_3902,N_2234,N_1552);
and U3903 (N_3903,N_1913,N_1673);
nand U3904 (N_3904,N_2487,N_2537);
nand U3905 (N_3905,N_2567,N_2240);
and U3906 (N_3906,N_2862,N_2617);
nor U3907 (N_3907,N_2899,N_1764);
and U3908 (N_3908,N_2182,N_2212);
or U3909 (N_3909,N_1607,N_1800);
nor U3910 (N_3910,N_2398,N_2004);
xnor U3911 (N_3911,N_2380,N_2941);
nand U3912 (N_3912,N_2310,N_2885);
and U3913 (N_3913,N_2294,N_2543);
and U3914 (N_3914,N_1505,N_1770);
xor U3915 (N_3915,N_2707,N_1627);
xnor U3916 (N_3916,N_2680,N_1743);
nor U3917 (N_3917,N_2891,N_1870);
or U3918 (N_3918,N_2771,N_2215);
and U3919 (N_3919,N_1580,N_2609);
nand U3920 (N_3920,N_2712,N_2273);
xor U3921 (N_3921,N_1750,N_2739);
and U3922 (N_3922,N_2837,N_2609);
and U3923 (N_3923,N_2870,N_1787);
or U3924 (N_3924,N_2761,N_2015);
nor U3925 (N_3925,N_2119,N_2509);
nand U3926 (N_3926,N_2263,N_2310);
and U3927 (N_3927,N_2568,N_1654);
or U3928 (N_3928,N_1849,N_1668);
nand U3929 (N_3929,N_1619,N_1943);
or U3930 (N_3930,N_2334,N_1796);
nand U3931 (N_3931,N_2220,N_1914);
xnor U3932 (N_3932,N_2035,N_1571);
xor U3933 (N_3933,N_2088,N_1677);
nor U3934 (N_3934,N_2213,N_2212);
or U3935 (N_3935,N_1802,N_2505);
nor U3936 (N_3936,N_1909,N_2749);
nor U3937 (N_3937,N_1712,N_1972);
and U3938 (N_3938,N_1535,N_2622);
and U3939 (N_3939,N_2684,N_2114);
nand U3940 (N_3940,N_2369,N_2752);
xor U3941 (N_3941,N_2911,N_2827);
or U3942 (N_3942,N_2085,N_2026);
nor U3943 (N_3943,N_2808,N_1832);
nor U3944 (N_3944,N_2149,N_2626);
nand U3945 (N_3945,N_2313,N_2148);
or U3946 (N_3946,N_2652,N_2990);
nor U3947 (N_3947,N_2901,N_2392);
and U3948 (N_3948,N_2132,N_1507);
or U3949 (N_3949,N_2007,N_2908);
and U3950 (N_3950,N_2648,N_2051);
and U3951 (N_3951,N_2117,N_2926);
and U3952 (N_3952,N_2778,N_2963);
or U3953 (N_3953,N_2316,N_2774);
nand U3954 (N_3954,N_1920,N_1519);
nand U3955 (N_3955,N_2858,N_1862);
xnor U3956 (N_3956,N_2123,N_2304);
xor U3957 (N_3957,N_2244,N_2622);
and U3958 (N_3958,N_1817,N_2335);
and U3959 (N_3959,N_2932,N_1556);
nor U3960 (N_3960,N_1679,N_1868);
xor U3961 (N_3961,N_2013,N_2839);
or U3962 (N_3962,N_2004,N_2166);
or U3963 (N_3963,N_2586,N_1649);
xor U3964 (N_3964,N_1879,N_2714);
xor U3965 (N_3965,N_2142,N_2660);
nand U3966 (N_3966,N_2677,N_2360);
nand U3967 (N_3967,N_1560,N_1866);
nor U3968 (N_3968,N_2188,N_2367);
or U3969 (N_3969,N_2782,N_1536);
xnor U3970 (N_3970,N_1825,N_2622);
and U3971 (N_3971,N_2449,N_1572);
nor U3972 (N_3972,N_1529,N_2289);
nor U3973 (N_3973,N_2263,N_1766);
nand U3974 (N_3974,N_1656,N_2718);
or U3975 (N_3975,N_2300,N_2229);
xor U3976 (N_3976,N_1806,N_2941);
or U3977 (N_3977,N_2389,N_2335);
and U3978 (N_3978,N_2017,N_2233);
nor U3979 (N_3979,N_2694,N_2250);
or U3980 (N_3980,N_2259,N_2337);
and U3981 (N_3981,N_2128,N_1859);
and U3982 (N_3982,N_1991,N_1831);
xor U3983 (N_3983,N_1524,N_2032);
or U3984 (N_3984,N_2406,N_1973);
and U3985 (N_3985,N_2914,N_2382);
nor U3986 (N_3986,N_1537,N_2287);
and U3987 (N_3987,N_1505,N_1980);
xnor U3988 (N_3988,N_2803,N_1859);
nor U3989 (N_3989,N_1799,N_1666);
or U3990 (N_3990,N_2655,N_2788);
and U3991 (N_3991,N_2296,N_2672);
or U3992 (N_3992,N_2387,N_1535);
and U3993 (N_3993,N_1517,N_2295);
and U3994 (N_3994,N_2687,N_2463);
nor U3995 (N_3995,N_2872,N_2373);
xor U3996 (N_3996,N_1694,N_2926);
and U3997 (N_3997,N_2802,N_2566);
or U3998 (N_3998,N_1637,N_1511);
nand U3999 (N_3999,N_1637,N_2093);
or U4000 (N_4000,N_2724,N_1609);
or U4001 (N_4001,N_2024,N_2917);
nor U4002 (N_4002,N_1830,N_1900);
nand U4003 (N_4003,N_2579,N_2270);
and U4004 (N_4004,N_2652,N_2274);
and U4005 (N_4005,N_1946,N_2589);
and U4006 (N_4006,N_2719,N_2622);
nand U4007 (N_4007,N_2717,N_2667);
nor U4008 (N_4008,N_2730,N_2390);
and U4009 (N_4009,N_1810,N_1626);
xor U4010 (N_4010,N_1801,N_2046);
xnor U4011 (N_4011,N_2214,N_2430);
or U4012 (N_4012,N_2324,N_2301);
and U4013 (N_4013,N_2141,N_1713);
nor U4014 (N_4014,N_2711,N_2688);
nand U4015 (N_4015,N_2755,N_2608);
nor U4016 (N_4016,N_2305,N_2854);
or U4017 (N_4017,N_1899,N_2524);
nor U4018 (N_4018,N_1910,N_2776);
nor U4019 (N_4019,N_2253,N_2043);
or U4020 (N_4020,N_2937,N_1725);
nor U4021 (N_4021,N_2842,N_1996);
xnor U4022 (N_4022,N_1902,N_2338);
nor U4023 (N_4023,N_1624,N_2642);
nor U4024 (N_4024,N_2879,N_1731);
nand U4025 (N_4025,N_1910,N_2263);
nand U4026 (N_4026,N_1856,N_2298);
or U4027 (N_4027,N_2539,N_2101);
nand U4028 (N_4028,N_2474,N_1830);
nand U4029 (N_4029,N_2056,N_1991);
or U4030 (N_4030,N_1627,N_2573);
and U4031 (N_4031,N_2556,N_2153);
and U4032 (N_4032,N_2973,N_1714);
xor U4033 (N_4033,N_2127,N_2207);
nand U4034 (N_4034,N_1973,N_1812);
nand U4035 (N_4035,N_2474,N_1647);
or U4036 (N_4036,N_2574,N_2166);
or U4037 (N_4037,N_1817,N_2519);
xor U4038 (N_4038,N_2875,N_1808);
or U4039 (N_4039,N_2899,N_2088);
and U4040 (N_4040,N_2346,N_2445);
nor U4041 (N_4041,N_2516,N_2579);
or U4042 (N_4042,N_1710,N_1959);
xor U4043 (N_4043,N_2956,N_2136);
and U4044 (N_4044,N_1746,N_2842);
nor U4045 (N_4045,N_2339,N_2674);
nand U4046 (N_4046,N_2187,N_2370);
xnor U4047 (N_4047,N_2509,N_1636);
nor U4048 (N_4048,N_2078,N_2638);
or U4049 (N_4049,N_1796,N_2944);
or U4050 (N_4050,N_2357,N_2899);
or U4051 (N_4051,N_2375,N_2866);
xnor U4052 (N_4052,N_2629,N_2255);
and U4053 (N_4053,N_2455,N_2050);
xnor U4054 (N_4054,N_2248,N_1893);
nand U4055 (N_4055,N_1708,N_2829);
nand U4056 (N_4056,N_2196,N_2359);
nand U4057 (N_4057,N_2569,N_2178);
xnor U4058 (N_4058,N_2327,N_2820);
and U4059 (N_4059,N_2928,N_2287);
nand U4060 (N_4060,N_1911,N_1727);
and U4061 (N_4061,N_1573,N_2793);
and U4062 (N_4062,N_2042,N_2891);
nand U4063 (N_4063,N_2677,N_1820);
nand U4064 (N_4064,N_1582,N_2046);
and U4065 (N_4065,N_2355,N_1898);
xor U4066 (N_4066,N_1684,N_2158);
and U4067 (N_4067,N_1905,N_1619);
nand U4068 (N_4068,N_1745,N_2514);
or U4069 (N_4069,N_2105,N_1760);
or U4070 (N_4070,N_2763,N_2398);
nor U4071 (N_4071,N_2284,N_2771);
nand U4072 (N_4072,N_2866,N_2638);
nor U4073 (N_4073,N_2115,N_2706);
or U4074 (N_4074,N_1980,N_1761);
nand U4075 (N_4075,N_2459,N_2660);
nor U4076 (N_4076,N_1830,N_1911);
xor U4077 (N_4077,N_2394,N_2833);
or U4078 (N_4078,N_2204,N_2947);
nand U4079 (N_4079,N_2677,N_1567);
nor U4080 (N_4080,N_1916,N_2310);
nand U4081 (N_4081,N_2542,N_2636);
nor U4082 (N_4082,N_2441,N_2699);
or U4083 (N_4083,N_1922,N_2362);
or U4084 (N_4084,N_2758,N_2410);
xor U4085 (N_4085,N_2396,N_2161);
nor U4086 (N_4086,N_1996,N_2855);
or U4087 (N_4087,N_2646,N_2058);
and U4088 (N_4088,N_2543,N_1979);
and U4089 (N_4089,N_2808,N_1741);
xor U4090 (N_4090,N_2437,N_2293);
or U4091 (N_4091,N_2646,N_2564);
xor U4092 (N_4092,N_2170,N_1525);
and U4093 (N_4093,N_1731,N_2268);
or U4094 (N_4094,N_2182,N_1931);
nor U4095 (N_4095,N_1982,N_2387);
nand U4096 (N_4096,N_2998,N_2273);
or U4097 (N_4097,N_2350,N_2791);
or U4098 (N_4098,N_1670,N_1815);
and U4099 (N_4099,N_1784,N_2055);
or U4100 (N_4100,N_1610,N_2938);
and U4101 (N_4101,N_2501,N_1967);
and U4102 (N_4102,N_2484,N_2644);
and U4103 (N_4103,N_2012,N_1909);
or U4104 (N_4104,N_2998,N_1713);
xnor U4105 (N_4105,N_1710,N_1674);
xor U4106 (N_4106,N_2128,N_2878);
and U4107 (N_4107,N_1876,N_1572);
nand U4108 (N_4108,N_1944,N_2661);
and U4109 (N_4109,N_2283,N_2147);
nor U4110 (N_4110,N_2757,N_2225);
nor U4111 (N_4111,N_2260,N_2197);
nand U4112 (N_4112,N_2735,N_2087);
nand U4113 (N_4113,N_2635,N_2574);
or U4114 (N_4114,N_1545,N_1912);
and U4115 (N_4115,N_2023,N_2336);
and U4116 (N_4116,N_2736,N_2151);
nand U4117 (N_4117,N_1806,N_2701);
nor U4118 (N_4118,N_2954,N_1667);
and U4119 (N_4119,N_2406,N_1868);
nor U4120 (N_4120,N_1766,N_2491);
xnor U4121 (N_4121,N_2161,N_1814);
nor U4122 (N_4122,N_2526,N_2216);
xor U4123 (N_4123,N_2194,N_2882);
nand U4124 (N_4124,N_2280,N_1821);
nand U4125 (N_4125,N_2638,N_2552);
nor U4126 (N_4126,N_1861,N_1809);
and U4127 (N_4127,N_1928,N_1972);
nand U4128 (N_4128,N_2519,N_2863);
nor U4129 (N_4129,N_2731,N_2572);
or U4130 (N_4130,N_2915,N_1506);
nor U4131 (N_4131,N_1925,N_1588);
xor U4132 (N_4132,N_1504,N_2227);
or U4133 (N_4133,N_2265,N_2193);
xnor U4134 (N_4134,N_2880,N_2461);
nand U4135 (N_4135,N_2982,N_2442);
and U4136 (N_4136,N_2894,N_2280);
xor U4137 (N_4137,N_1623,N_2358);
xnor U4138 (N_4138,N_1861,N_2110);
or U4139 (N_4139,N_2282,N_2628);
nand U4140 (N_4140,N_2714,N_2011);
xnor U4141 (N_4141,N_1869,N_1841);
nor U4142 (N_4142,N_2762,N_2556);
and U4143 (N_4143,N_2246,N_2651);
or U4144 (N_4144,N_2067,N_1803);
nand U4145 (N_4145,N_1861,N_2216);
xor U4146 (N_4146,N_2440,N_1998);
and U4147 (N_4147,N_2887,N_2569);
nand U4148 (N_4148,N_2422,N_2031);
xor U4149 (N_4149,N_1995,N_2882);
xor U4150 (N_4150,N_1608,N_1554);
nand U4151 (N_4151,N_1808,N_2714);
nor U4152 (N_4152,N_2280,N_2481);
xor U4153 (N_4153,N_2092,N_2254);
and U4154 (N_4154,N_2985,N_2703);
nand U4155 (N_4155,N_2471,N_2585);
xor U4156 (N_4156,N_1829,N_2518);
nand U4157 (N_4157,N_2497,N_2004);
nor U4158 (N_4158,N_1980,N_1702);
or U4159 (N_4159,N_2800,N_2960);
nand U4160 (N_4160,N_1587,N_1820);
xor U4161 (N_4161,N_2300,N_2122);
nor U4162 (N_4162,N_2632,N_2653);
nand U4163 (N_4163,N_2254,N_1832);
nand U4164 (N_4164,N_2123,N_1888);
and U4165 (N_4165,N_2752,N_1775);
or U4166 (N_4166,N_1755,N_2491);
xnor U4167 (N_4167,N_2583,N_1509);
nor U4168 (N_4168,N_2624,N_2336);
xor U4169 (N_4169,N_2180,N_1654);
xnor U4170 (N_4170,N_2221,N_2751);
nor U4171 (N_4171,N_1840,N_1987);
xnor U4172 (N_4172,N_2531,N_2971);
nor U4173 (N_4173,N_2389,N_2132);
or U4174 (N_4174,N_1748,N_1928);
and U4175 (N_4175,N_2706,N_2392);
nor U4176 (N_4176,N_1800,N_2752);
xor U4177 (N_4177,N_2677,N_2025);
and U4178 (N_4178,N_2536,N_2011);
and U4179 (N_4179,N_1784,N_2203);
or U4180 (N_4180,N_2673,N_2159);
and U4181 (N_4181,N_2934,N_2279);
nor U4182 (N_4182,N_2701,N_2242);
or U4183 (N_4183,N_2303,N_2581);
nand U4184 (N_4184,N_2755,N_2264);
nand U4185 (N_4185,N_1544,N_2046);
and U4186 (N_4186,N_2590,N_1818);
or U4187 (N_4187,N_2852,N_1800);
or U4188 (N_4188,N_2742,N_2754);
or U4189 (N_4189,N_1721,N_1604);
and U4190 (N_4190,N_1563,N_2093);
and U4191 (N_4191,N_1973,N_2138);
nand U4192 (N_4192,N_2940,N_2020);
nand U4193 (N_4193,N_1779,N_2685);
xnor U4194 (N_4194,N_2888,N_1881);
or U4195 (N_4195,N_1802,N_1896);
nand U4196 (N_4196,N_1900,N_1725);
nor U4197 (N_4197,N_2067,N_1610);
nor U4198 (N_4198,N_1970,N_1646);
nor U4199 (N_4199,N_1938,N_2951);
nand U4200 (N_4200,N_2308,N_2782);
nand U4201 (N_4201,N_1861,N_2009);
or U4202 (N_4202,N_2069,N_2618);
nand U4203 (N_4203,N_1682,N_2627);
nand U4204 (N_4204,N_2730,N_2534);
xnor U4205 (N_4205,N_1827,N_1550);
nor U4206 (N_4206,N_2513,N_1858);
nand U4207 (N_4207,N_1707,N_2742);
xor U4208 (N_4208,N_2786,N_2737);
and U4209 (N_4209,N_2875,N_2572);
and U4210 (N_4210,N_2746,N_2609);
xor U4211 (N_4211,N_2446,N_2822);
or U4212 (N_4212,N_2179,N_1797);
and U4213 (N_4213,N_2362,N_1850);
or U4214 (N_4214,N_2008,N_2379);
or U4215 (N_4215,N_2512,N_2029);
nor U4216 (N_4216,N_2613,N_1742);
xnor U4217 (N_4217,N_2581,N_1739);
and U4218 (N_4218,N_2022,N_2651);
and U4219 (N_4219,N_2526,N_2604);
xnor U4220 (N_4220,N_2215,N_1655);
nand U4221 (N_4221,N_1962,N_1993);
nand U4222 (N_4222,N_2376,N_2815);
or U4223 (N_4223,N_1823,N_2293);
nand U4224 (N_4224,N_2427,N_2366);
nand U4225 (N_4225,N_1877,N_2284);
nor U4226 (N_4226,N_2540,N_2614);
nand U4227 (N_4227,N_2043,N_1538);
nand U4228 (N_4228,N_1934,N_2480);
or U4229 (N_4229,N_1999,N_1787);
nor U4230 (N_4230,N_2601,N_2048);
nor U4231 (N_4231,N_2715,N_2465);
nand U4232 (N_4232,N_2229,N_1675);
and U4233 (N_4233,N_1946,N_2170);
nor U4234 (N_4234,N_2598,N_2669);
xnor U4235 (N_4235,N_2223,N_2213);
and U4236 (N_4236,N_2842,N_2759);
or U4237 (N_4237,N_2913,N_2561);
or U4238 (N_4238,N_1538,N_1880);
nor U4239 (N_4239,N_1769,N_2056);
and U4240 (N_4240,N_2007,N_2136);
xnor U4241 (N_4241,N_1807,N_2327);
or U4242 (N_4242,N_2312,N_1592);
nand U4243 (N_4243,N_2111,N_2522);
or U4244 (N_4244,N_1563,N_2621);
or U4245 (N_4245,N_1649,N_2452);
xnor U4246 (N_4246,N_1997,N_2760);
nor U4247 (N_4247,N_2694,N_2401);
xor U4248 (N_4248,N_1803,N_1760);
and U4249 (N_4249,N_2277,N_2013);
nand U4250 (N_4250,N_2899,N_2876);
and U4251 (N_4251,N_2813,N_1667);
and U4252 (N_4252,N_2274,N_2238);
nand U4253 (N_4253,N_2180,N_2988);
or U4254 (N_4254,N_2001,N_2887);
xnor U4255 (N_4255,N_1852,N_2794);
nor U4256 (N_4256,N_1737,N_2905);
and U4257 (N_4257,N_2221,N_1990);
or U4258 (N_4258,N_2267,N_2738);
xor U4259 (N_4259,N_1874,N_2590);
and U4260 (N_4260,N_1971,N_1879);
or U4261 (N_4261,N_2301,N_2933);
nor U4262 (N_4262,N_2667,N_2676);
or U4263 (N_4263,N_2506,N_1586);
nor U4264 (N_4264,N_2062,N_2317);
nor U4265 (N_4265,N_2833,N_1686);
xor U4266 (N_4266,N_2109,N_1714);
nand U4267 (N_4267,N_2226,N_1837);
nand U4268 (N_4268,N_2771,N_2191);
nand U4269 (N_4269,N_2241,N_1998);
nor U4270 (N_4270,N_1774,N_2470);
xor U4271 (N_4271,N_2967,N_2653);
nand U4272 (N_4272,N_2815,N_1724);
nand U4273 (N_4273,N_1610,N_2621);
nor U4274 (N_4274,N_1596,N_2677);
nor U4275 (N_4275,N_2764,N_2294);
nor U4276 (N_4276,N_2640,N_2028);
nand U4277 (N_4277,N_2912,N_2807);
and U4278 (N_4278,N_1505,N_1812);
nand U4279 (N_4279,N_2039,N_2263);
xor U4280 (N_4280,N_2911,N_2640);
and U4281 (N_4281,N_2342,N_2190);
nor U4282 (N_4282,N_1940,N_2870);
or U4283 (N_4283,N_2059,N_2926);
or U4284 (N_4284,N_2251,N_2360);
and U4285 (N_4285,N_2641,N_2113);
or U4286 (N_4286,N_2910,N_2614);
or U4287 (N_4287,N_2626,N_2396);
nand U4288 (N_4288,N_2892,N_1581);
or U4289 (N_4289,N_1569,N_2973);
nand U4290 (N_4290,N_2627,N_1864);
or U4291 (N_4291,N_2200,N_1918);
nand U4292 (N_4292,N_2924,N_2926);
nor U4293 (N_4293,N_1783,N_2998);
or U4294 (N_4294,N_1576,N_1601);
nor U4295 (N_4295,N_1678,N_1687);
xnor U4296 (N_4296,N_2149,N_2045);
nor U4297 (N_4297,N_1782,N_2843);
or U4298 (N_4298,N_2829,N_2675);
nor U4299 (N_4299,N_1557,N_2919);
nand U4300 (N_4300,N_1977,N_2994);
xnor U4301 (N_4301,N_2294,N_2643);
nand U4302 (N_4302,N_2826,N_2843);
nand U4303 (N_4303,N_1793,N_2440);
and U4304 (N_4304,N_2763,N_2879);
or U4305 (N_4305,N_2639,N_1839);
or U4306 (N_4306,N_2272,N_2298);
or U4307 (N_4307,N_1707,N_1837);
and U4308 (N_4308,N_2466,N_2608);
xor U4309 (N_4309,N_2434,N_2097);
and U4310 (N_4310,N_1594,N_2801);
and U4311 (N_4311,N_2619,N_2922);
nor U4312 (N_4312,N_2507,N_1709);
nor U4313 (N_4313,N_2593,N_2806);
and U4314 (N_4314,N_2689,N_1821);
and U4315 (N_4315,N_1515,N_2188);
and U4316 (N_4316,N_2550,N_1783);
xnor U4317 (N_4317,N_2192,N_2380);
xor U4318 (N_4318,N_2671,N_1603);
nor U4319 (N_4319,N_2737,N_2871);
nor U4320 (N_4320,N_2326,N_2519);
and U4321 (N_4321,N_2133,N_2860);
or U4322 (N_4322,N_2184,N_1677);
nand U4323 (N_4323,N_1973,N_2470);
and U4324 (N_4324,N_1996,N_2409);
nand U4325 (N_4325,N_2786,N_1551);
nand U4326 (N_4326,N_2667,N_2322);
nor U4327 (N_4327,N_1507,N_1592);
nand U4328 (N_4328,N_2370,N_1853);
or U4329 (N_4329,N_2033,N_2629);
nand U4330 (N_4330,N_2494,N_2115);
xor U4331 (N_4331,N_2319,N_2503);
and U4332 (N_4332,N_2738,N_1821);
nand U4333 (N_4333,N_2935,N_1964);
nor U4334 (N_4334,N_1839,N_1598);
nor U4335 (N_4335,N_2068,N_1901);
or U4336 (N_4336,N_1789,N_2166);
nand U4337 (N_4337,N_2482,N_1801);
nand U4338 (N_4338,N_1691,N_1843);
nand U4339 (N_4339,N_2091,N_1548);
and U4340 (N_4340,N_2221,N_1629);
and U4341 (N_4341,N_1797,N_1839);
nor U4342 (N_4342,N_2171,N_2874);
nor U4343 (N_4343,N_2201,N_1731);
nand U4344 (N_4344,N_2792,N_1922);
or U4345 (N_4345,N_1941,N_2075);
and U4346 (N_4346,N_2070,N_1793);
or U4347 (N_4347,N_2008,N_2667);
and U4348 (N_4348,N_2745,N_2216);
nor U4349 (N_4349,N_1743,N_2979);
and U4350 (N_4350,N_2739,N_2601);
xnor U4351 (N_4351,N_2697,N_2344);
and U4352 (N_4352,N_2925,N_2187);
xnor U4353 (N_4353,N_1984,N_1722);
nand U4354 (N_4354,N_1746,N_1884);
and U4355 (N_4355,N_2377,N_1939);
nand U4356 (N_4356,N_2061,N_1731);
nor U4357 (N_4357,N_2125,N_1853);
nand U4358 (N_4358,N_1800,N_1873);
or U4359 (N_4359,N_2165,N_1580);
xnor U4360 (N_4360,N_1533,N_2006);
and U4361 (N_4361,N_1666,N_2986);
xnor U4362 (N_4362,N_2120,N_2427);
nand U4363 (N_4363,N_2856,N_1559);
or U4364 (N_4364,N_2571,N_2093);
xnor U4365 (N_4365,N_2046,N_2975);
nand U4366 (N_4366,N_2538,N_2023);
nand U4367 (N_4367,N_2792,N_2085);
and U4368 (N_4368,N_1960,N_2566);
nor U4369 (N_4369,N_1928,N_2194);
and U4370 (N_4370,N_2907,N_2240);
and U4371 (N_4371,N_1711,N_2291);
xnor U4372 (N_4372,N_2110,N_2091);
xnor U4373 (N_4373,N_2935,N_1576);
nor U4374 (N_4374,N_2021,N_2296);
or U4375 (N_4375,N_1595,N_2498);
or U4376 (N_4376,N_2945,N_2503);
and U4377 (N_4377,N_2185,N_1624);
or U4378 (N_4378,N_2084,N_2373);
or U4379 (N_4379,N_2932,N_2891);
and U4380 (N_4380,N_1563,N_1884);
and U4381 (N_4381,N_2494,N_1795);
xor U4382 (N_4382,N_1799,N_1780);
and U4383 (N_4383,N_2010,N_2166);
and U4384 (N_4384,N_2205,N_2386);
nor U4385 (N_4385,N_2844,N_1809);
or U4386 (N_4386,N_2842,N_2979);
or U4387 (N_4387,N_2583,N_1731);
nor U4388 (N_4388,N_1558,N_1812);
xnor U4389 (N_4389,N_2965,N_1721);
or U4390 (N_4390,N_1970,N_1881);
nor U4391 (N_4391,N_2599,N_2186);
or U4392 (N_4392,N_2930,N_1550);
or U4393 (N_4393,N_2263,N_2082);
nor U4394 (N_4394,N_2544,N_1646);
and U4395 (N_4395,N_2798,N_1682);
xnor U4396 (N_4396,N_1711,N_1814);
nor U4397 (N_4397,N_2087,N_2671);
and U4398 (N_4398,N_1688,N_1529);
and U4399 (N_4399,N_2699,N_2761);
or U4400 (N_4400,N_1826,N_1798);
xor U4401 (N_4401,N_1998,N_2046);
nor U4402 (N_4402,N_1605,N_2918);
xor U4403 (N_4403,N_2169,N_2658);
or U4404 (N_4404,N_2707,N_2918);
or U4405 (N_4405,N_1896,N_1500);
nor U4406 (N_4406,N_1891,N_1648);
nor U4407 (N_4407,N_2483,N_2184);
and U4408 (N_4408,N_2560,N_1526);
nand U4409 (N_4409,N_2931,N_2928);
and U4410 (N_4410,N_2710,N_2654);
and U4411 (N_4411,N_2648,N_2759);
xor U4412 (N_4412,N_1547,N_2856);
and U4413 (N_4413,N_1587,N_2559);
and U4414 (N_4414,N_2816,N_1578);
xor U4415 (N_4415,N_2608,N_2359);
xor U4416 (N_4416,N_1904,N_1745);
nand U4417 (N_4417,N_2889,N_2289);
nand U4418 (N_4418,N_2502,N_2856);
xor U4419 (N_4419,N_1830,N_2833);
or U4420 (N_4420,N_2321,N_2086);
xnor U4421 (N_4421,N_2029,N_2193);
xnor U4422 (N_4422,N_1597,N_1914);
nand U4423 (N_4423,N_2106,N_2654);
nand U4424 (N_4424,N_2024,N_2204);
and U4425 (N_4425,N_1570,N_1709);
xor U4426 (N_4426,N_2240,N_2002);
nand U4427 (N_4427,N_2016,N_2127);
or U4428 (N_4428,N_2789,N_2037);
nor U4429 (N_4429,N_2949,N_1684);
xor U4430 (N_4430,N_2321,N_2143);
nand U4431 (N_4431,N_1708,N_2290);
xor U4432 (N_4432,N_1639,N_2005);
nor U4433 (N_4433,N_2283,N_2757);
nor U4434 (N_4434,N_2587,N_2467);
nand U4435 (N_4435,N_2445,N_2342);
or U4436 (N_4436,N_2990,N_2680);
or U4437 (N_4437,N_2052,N_2404);
xor U4438 (N_4438,N_1704,N_1849);
and U4439 (N_4439,N_2388,N_2183);
or U4440 (N_4440,N_2812,N_1814);
and U4441 (N_4441,N_2683,N_2330);
or U4442 (N_4442,N_1974,N_2129);
and U4443 (N_4443,N_1953,N_2197);
nand U4444 (N_4444,N_2671,N_2863);
xnor U4445 (N_4445,N_2045,N_2496);
nor U4446 (N_4446,N_2469,N_1843);
nand U4447 (N_4447,N_2177,N_2655);
and U4448 (N_4448,N_1693,N_2085);
nand U4449 (N_4449,N_1596,N_2337);
xnor U4450 (N_4450,N_1552,N_1557);
nand U4451 (N_4451,N_2040,N_2542);
or U4452 (N_4452,N_2229,N_1867);
or U4453 (N_4453,N_2409,N_1529);
or U4454 (N_4454,N_2437,N_1779);
xor U4455 (N_4455,N_1705,N_2587);
and U4456 (N_4456,N_2893,N_1524);
and U4457 (N_4457,N_2701,N_2355);
nand U4458 (N_4458,N_2990,N_2320);
xor U4459 (N_4459,N_2866,N_2991);
nor U4460 (N_4460,N_2811,N_2234);
nor U4461 (N_4461,N_2976,N_2372);
nand U4462 (N_4462,N_1565,N_1532);
nor U4463 (N_4463,N_2876,N_2125);
nor U4464 (N_4464,N_1754,N_1981);
nand U4465 (N_4465,N_2950,N_2077);
nor U4466 (N_4466,N_1976,N_2929);
or U4467 (N_4467,N_2893,N_1675);
nand U4468 (N_4468,N_2519,N_1541);
xor U4469 (N_4469,N_1710,N_2283);
xnor U4470 (N_4470,N_2444,N_2357);
nand U4471 (N_4471,N_2628,N_2524);
and U4472 (N_4472,N_2310,N_1831);
nor U4473 (N_4473,N_1507,N_1958);
nand U4474 (N_4474,N_2459,N_2762);
nor U4475 (N_4475,N_2989,N_2548);
xnor U4476 (N_4476,N_1741,N_2971);
or U4477 (N_4477,N_1589,N_2437);
nor U4478 (N_4478,N_1883,N_1642);
xor U4479 (N_4479,N_1570,N_2711);
xor U4480 (N_4480,N_1953,N_2125);
nand U4481 (N_4481,N_2722,N_2438);
nor U4482 (N_4482,N_1747,N_2656);
xor U4483 (N_4483,N_2104,N_1951);
nand U4484 (N_4484,N_2467,N_2619);
nor U4485 (N_4485,N_2605,N_2546);
and U4486 (N_4486,N_1529,N_2231);
and U4487 (N_4487,N_2810,N_1824);
nand U4488 (N_4488,N_1613,N_2346);
nand U4489 (N_4489,N_1748,N_2037);
nor U4490 (N_4490,N_2014,N_2751);
nand U4491 (N_4491,N_1535,N_2656);
nand U4492 (N_4492,N_2384,N_1531);
or U4493 (N_4493,N_2352,N_2588);
nand U4494 (N_4494,N_2548,N_2438);
xnor U4495 (N_4495,N_1518,N_2656);
and U4496 (N_4496,N_2252,N_2422);
xnor U4497 (N_4497,N_1842,N_2226);
and U4498 (N_4498,N_1806,N_2170);
nand U4499 (N_4499,N_2126,N_2287);
or U4500 (N_4500,N_4458,N_3657);
nand U4501 (N_4501,N_4152,N_3650);
nor U4502 (N_4502,N_3468,N_3646);
nor U4503 (N_4503,N_3005,N_3125);
xnor U4504 (N_4504,N_3945,N_4463);
xnor U4505 (N_4505,N_3420,N_3807);
xor U4506 (N_4506,N_3327,N_3557);
or U4507 (N_4507,N_4241,N_3237);
or U4508 (N_4508,N_3553,N_4027);
or U4509 (N_4509,N_3061,N_3598);
nor U4510 (N_4510,N_3530,N_4119);
nand U4511 (N_4511,N_3373,N_3589);
nor U4512 (N_4512,N_3289,N_4182);
or U4513 (N_4513,N_4403,N_3078);
and U4514 (N_4514,N_4347,N_3789);
nor U4515 (N_4515,N_3439,N_4321);
xnor U4516 (N_4516,N_3744,N_3753);
and U4517 (N_4517,N_4166,N_4485);
xor U4518 (N_4518,N_3385,N_3546);
or U4519 (N_4519,N_4419,N_3834);
xnor U4520 (N_4520,N_4102,N_4329);
xor U4521 (N_4521,N_3428,N_3678);
and U4522 (N_4522,N_3860,N_4429);
xnor U4523 (N_4523,N_4272,N_4250);
and U4524 (N_4524,N_4201,N_3474);
and U4525 (N_4525,N_3829,N_3665);
nand U4526 (N_4526,N_4083,N_3907);
nor U4527 (N_4527,N_3479,N_4376);
and U4528 (N_4528,N_3196,N_3680);
and U4529 (N_4529,N_4494,N_3785);
nor U4530 (N_4530,N_3565,N_3084);
or U4531 (N_4531,N_3914,N_3540);
or U4532 (N_4532,N_3029,N_3195);
nor U4533 (N_4533,N_4425,N_4067);
nor U4534 (N_4534,N_4495,N_4255);
or U4535 (N_4535,N_4389,N_3126);
and U4536 (N_4536,N_3316,N_4412);
and U4537 (N_4537,N_3982,N_3701);
and U4538 (N_4538,N_3086,N_3072);
or U4539 (N_4539,N_4123,N_4113);
and U4540 (N_4540,N_3963,N_3936);
xor U4541 (N_4541,N_3840,N_3525);
and U4542 (N_4542,N_4088,N_3164);
xor U4543 (N_4543,N_3376,N_3688);
xnor U4544 (N_4544,N_4072,N_4087);
and U4545 (N_4545,N_3818,N_3762);
nand U4546 (N_4546,N_3051,N_3413);
and U4547 (N_4547,N_4266,N_4396);
xor U4548 (N_4548,N_3896,N_4222);
nand U4549 (N_4549,N_3023,N_3791);
and U4550 (N_4550,N_3148,N_3802);
nor U4551 (N_4551,N_3836,N_3841);
or U4552 (N_4552,N_3358,N_4218);
nor U4553 (N_4553,N_3383,N_4183);
xnor U4554 (N_4554,N_3793,N_3177);
nor U4555 (N_4555,N_3719,N_3313);
nor U4556 (N_4556,N_3600,N_3690);
nand U4557 (N_4557,N_4033,N_4147);
nor U4558 (N_4558,N_3276,N_3891);
nor U4559 (N_4559,N_3294,N_3861);
or U4560 (N_4560,N_3070,N_3928);
nor U4561 (N_4561,N_3803,N_3496);
nor U4562 (N_4562,N_4435,N_4015);
or U4563 (N_4563,N_4338,N_4217);
nor U4564 (N_4564,N_3161,N_3894);
and U4565 (N_4565,N_4034,N_3149);
and U4566 (N_4566,N_3619,N_3140);
nor U4567 (N_4567,N_3285,N_3042);
or U4568 (N_4568,N_3938,N_3951);
xor U4569 (N_4569,N_3849,N_3142);
and U4570 (N_4570,N_3255,N_3747);
and U4571 (N_4571,N_3623,N_3563);
and U4572 (N_4572,N_3347,N_4098);
xor U4573 (N_4573,N_4068,N_3988);
or U4574 (N_4574,N_4232,N_4256);
xor U4575 (N_4575,N_4089,N_4416);
nor U4576 (N_4576,N_4176,N_4439);
nor U4577 (N_4577,N_4044,N_3918);
or U4578 (N_4578,N_4353,N_3873);
nand U4579 (N_4579,N_4137,N_4341);
and U4580 (N_4580,N_3471,N_3882);
nand U4581 (N_4581,N_3422,N_3201);
nor U4582 (N_4582,N_3721,N_3735);
nand U4583 (N_4583,N_4246,N_3733);
xnor U4584 (N_4584,N_4282,N_3737);
xnor U4585 (N_4585,N_3870,N_4368);
nor U4586 (N_4586,N_4112,N_4086);
nand U4587 (N_4587,N_3387,N_4314);
or U4588 (N_4588,N_3813,N_4358);
nand U4589 (N_4589,N_4103,N_3607);
or U4590 (N_4590,N_4342,N_4226);
nand U4591 (N_4591,N_3630,N_3390);
nor U4592 (N_4592,N_4168,N_4150);
and U4593 (N_4593,N_4165,N_3279);
xor U4594 (N_4594,N_3363,N_3094);
and U4595 (N_4595,N_3323,N_3955);
xnor U4596 (N_4596,N_3628,N_4170);
and U4597 (N_4597,N_4462,N_3476);
nand U4598 (N_4598,N_4016,N_4133);
or U4599 (N_4599,N_3238,N_3651);
nand U4600 (N_4600,N_4415,N_3093);
xor U4601 (N_4601,N_4424,N_3123);
xor U4602 (N_4602,N_3248,N_4148);
xnor U4603 (N_4603,N_3103,N_3927);
nor U4604 (N_4604,N_3585,N_4288);
or U4605 (N_4605,N_3591,N_3754);
and U4606 (N_4606,N_3906,N_4229);
and U4607 (N_4607,N_4242,N_3321);
nand U4608 (N_4608,N_3368,N_4264);
and U4609 (N_4609,N_4134,N_4049);
nand U4610 (N_4610,N_3096,N_4344);
xnor U4611 (N_4611,N_3348,N_3832);
nor U4612 (N_4612,N_3996,N_4171);
or U4613 (N_4613,N_4193,N_4230);
nand U4614 (N_4614,N_4449,N_4110);
nand U4615 (N_4615,N_4215,N_3682);
xor U4616 (N_4616,N_3709,N_4140);
nor U4617 (N_4617,N_3915,N_3118);
and U4618 (N_4618,N_3160,N_4409);
nand U4619 (N_4619,N_3231,N_3229);
xor U4620 (N_4620,N_3157,N_3887);
and U4621 (N_4621,N_3384,N_4333);
and U4622 (N_4622,N_4181,N_3169);
nor U4623 (N_4623,N_3127,N_4444);
or U4624 (N_4624,N_3819,N_3314);
xor U4625 (N_4625,N_4410,N_3909);
xor U4626 (N_4626,N_3119,N_4395);
or U4627 (N_4627,N_3505,N_4002);
nand U4628 (N_4628,N_3062,N_3147);
xor U4629 (N_4629,N_3247,N_4335);
and U4630 (N_4630,N_3026,N_4196);
nand U4631 (N_4631,N_4317,N_3179);
xor U4632 (N_4632,N_4488,N_3935);
nor U4633 (N_4633,N_3040,N_4109);
nand U4634 (N_4634,N_4418,N_3187);
and U4635 (N_4635,N_4290,N_3724);
nand U4636 (N_4636,N_3957,N_3322);
or U4637 (N_4637,N_3274,N_4178);
nor U4638 (N_4638,N_3796,N_3568);
and U4639 (N_4639,N_3240,N_4006);
or U4640 (N_4640,N_4292,N_3280);
xnor U4641 (N_4641,N_3369,N_4496);
and U4642 (N_4642,N_4008,N_3450);
or U4643 (N_4643,N_4378,N_4074);
nand U4644 (N_4644,N_3794,N_3975);
nor U4645 (N_4645,N_3020,N_3397);
xnor U4646 (N_4646,N_4304,N_3964);
xnor U4647 (N_4647,N_3635,N_3949);
xor U4648 (N_4648,N_4090,N_4271);
xnor U4649 (N_4649,N_3222,N_4312);
and U4650 (N_4650,N_3859,N_3353);
nand U4651 (N_4651,N_3720,N_3867);
nand U4652 (N_4652,N_4268,N_3488);
nor U4653 (N_4653,N_3249,N_3761);
xor U4654 (N_4654,N_3311,N_3087);
nor U4655 (N_4655,N_4153,N_4146);
nor U4656 (N_4656,N_3265,N_3204);
or U4657 (N_4657,N_3614,N_3932);
nand U4658 (N_4658,N_4190,N_3561);
xnor U4659 (N_4659,N_3245,N_3745);
nand U4660 (N_4660,N_3082,N_4469);
xnor U4661 (N_4661,N_4031,N_3017);
nor U4662 (N_4662,N_3681,N_3842);
and U4663 (N_4663,N_3624,N_4298);
and U4664 (N_4664,N_4007,N_4340);
nand U4665 (N_4665,N_3299,N_3828);
or U4666 (N_4666,N_3548,N_3770);
xnor U4667 (N_4667,N_3684,N_3729);
nor U4668 (N_4668,N_3111,N_3535);
xnor U4669 (N_4669,N_3167,N_3137);
or U4670 (N_4670,N_3267,N_3406);
and U4671 (N_4671,N_4050,N_4348);
xor U4672 (N_4672,N_3423,N_4194);
xor U4673 (N_4673,N_4057,N_3806);
nor U4674 (N_4674,N_3995,N_3604);
xnor U4675 (N_4675,N_4157,N_4004);
or U4676 (N_4676,N_4022,N_3310);
or U4677 (N_4677,N_3531,N_4077);
and U4678 (N_4678,N_4069,N_3120);
xnor U4679 (N_4679,N_3158,N_3798);
and U4680 (N_4680,N_3097,N_4399);
nand U4681 (N_4681,N_3594,N_3526);
or U4682 (N_4682,N_3966,N_3045);
nor U4683 (N_4683,N_3349,N_3226);
nor U4684 (N_4684,N_4413,N_4097);
and U4685 (N_4685,N_3595,N_3779);
xnor U4686 (N_4686,N_3482,N_3402);
nor U4687 (N_4687,N_4404,N_3025);
xor U4688 (N_4688,N_3580,N_3629);
xnor U4689 (N_4689,N_4186,N_3207);
nor U4690 (N_4690,N_3990,N_3631);
and U4691 (N_4691,N_3980,N_3795);
nor U4692 (N_4692,N_3708,N_3511);
nand U4693 (N_4693,N_3246,N_3380);
nor U4694 (N_4694,N_4203,N_4446);
nand U4695 (N_4695,N_4204,N_4056);
nor U4696 (N_4696,N_3426,N_4243);
xnor U4697 (N_4697,N_3254,N_3797);
nand U4698 (N_4698,N_4048,N_3736);
nor U4699 (N_4699,N_3883,N_4441);
nor U4700 (N_4700,N_3880,N_3277);
or U4701 (N_4701,N_3364,N_3220);
or U4702 (N_4702,N_3663,N_3816);
xor U4703 (N_4703,N_3890,N_3573);
or U4704 (N_4704,N_3083,N_4038);
or U4705 (N_4705,N_3973,N_3529);
and U4706 (N_4706,N_3054,N_4212);
nand U4707 (N_4707,N_4483,N_4065);
nor U4708 (N_4708,N_3350,N_3898);
xnor U4709 (N_4709,N_4106,N_4244);
nand U4710 (N_4710,N_4427,N_4411);
xnor U4711 (N_4711,N_3372,N_3952);
and U4712 (N_4712,N_3462,N_3637);
or U4713 (N_4713,N_3108,N_4319);
nand U4714 (N_4714,N_3773,N_3676);
nand U4715 (N_4715,N_3830,N_4258);
and U4716 (N_4716,N_3176,N_4345);
and U4717 (N_4717,N_3930,N_4346);
xnor U4718 (N_4718,N_3857,N_3702);
nor U4719 (N_4719,N_4055,N_4281);
nand U4720 (N_4720,N_4471,N_3415);
nand U4721 (N_4721,N_4421,N_3049);
nand U4722 (N_4722,N_3214,N_4401);
nand U4723 (N_4723,N_3800,N_4052);
nor U4724 (N_4724,N_3771,N_3519);
or U4725 (N_4725,N_3003,N_3257);
and U4726 (N_4726,N_3811,N_3691);
xor U4727 (N_4727,N_4267,N_3085);
xor U4728 (N_4728,N_3664,N_3694);
nor U4729 (N_4729,N_4012,N_4252);
and U4730 (N_4730,N_3200,N_4436);
or U4731 (N_4731,N_4315,N_3461);
nor U4732 (N_4732,N_4122,N_3991);
nand U4733 (N_4733,N_3292,N_3903);
nand U4734 (N_4734,N_3940,N_3617);
and U4735 (N_4735,N_3517,N_4114);
and U4736 (N_4736,N_3784,N_3258);
nor U4737 (N_4737,N_3063,N_3188);
or U4738 (N_4738,N_4035,N_3477);
or U4739 (N_4739,N_3215,N_3578);
or U4740 (N_4740,N_3414,N_4187);
or U4741 (N_4741,N_3185,N_4308);
xor U4742 (N_4742,N_3022,N_3239);
or U4743 (N_4743,N_4461,N_3850);
and U4744 (N_4744,N_3046,N_3616);
nor U4745 (N_4745,N_3053,N_3154);
and U4746 (N_4746,N_4270,N_3031);
xnor U4747 (N_4747,N_3558,N_3815);
xor U4748 (N_4748,N_3303,N_4386);
xnor U4749 (N_4749,N_3581,N_3065);
or U4750 (N_4750,N_4477,N_3560);
nor U4751 (N_4751,N_3632,N_3041);
and U4752 (N_4752,N_3218,N_3012);
xnor U4753 (N_4753,N_4082,N_3057);
xor U4754 (N_4754,N_3463,N_3067);
nor U4755 (N_4755,N_4259,N_3184);
or U4756 (N_4756,N_4286,N_3722);
and U4757 (N_4757,N_3440,N_4115);
and U4758 (N_4758,N_4111,N_3498);
nand U4759 (N_4759,N_3537,N_3693);
xnor U4760 (N_4760,N_3875,N_4126);
nand U4761 (N_4761,N_3844,N_3015);
xnor U4762 (N_4762,N_3924,N_4490);
and U4763 (N_4763,N_3804,N_4375);
nor U4764 (N_4764,N_3455,N_4239);
and U4765 (N_4765,N_3603,N_3683);
and U4766 (N_4766,N_3748,N_3534);
or U4767 (N_4767,N_3494,N_3692);
nor U4768 (N_4768,N_3432,N_3835);
and U4769 (N_4769,N_3538,N_4118);
xnor U4770 (N_4770,N_3030,N_4323);
and U4771 (N_4771,N_3933,N_3109);
xor U4772 (N_4772,N_3636,N_4400);
nor U4773 (N_4773,N_4177,N_3590);
nor U4774 (N_4774,N_4328,N_3715);
and U4775 (N_4775,N_3904,N_3901);
or U4776 (N_4776,N_3714,N_4360);
xor U4777 (N_4777,N_3344,N_3837);
nand U4778 (N_4778,N_4017,N_4433);
and U4779 (N_4779,N_4381,N_3532);
and U4780 (N_4780,N_4269,N_3317);
nor U4781 (N_4781,N_3515,N_3902);
nor U4782 (N_4782,N_3513,N_3879);
nor U4783 (N_4783,N_3886,N_3298);
and U4784 (N_4784,N_4359,N_4417);
nand U4785 (N_4785,N_4064,N_3550);
nor U4786 (N_4786,N_4382,N_3954);
or U4787 (N_4787,N_3001,N_3984);
nand U4788 (N_4788,N_4159,N_3081);
xor U4789 (N_4789,N_3472,N_4300);
nor U4790 (N_4790,N_3328,N_4213);
and U4791 (N_4791,N_3301,N_3900);
and U4792 (N_4792,N_3131,N_3679);
and U4793 (N_4793,N_4135,N_3790);
and U4794 (N_4794,N_3574,N_3166);
or U4795 (N_4795,N_3738,N_3765);
nand U4796 (N_4796,N_4330,N_3400);
nand U4797 (N_4797,N_3611,N_3981);
xnor U4798 (N_4798,N_3024,N_4060);
and U4799 (N_4799,N_4374,N_3028);
nor U4800 (N_4800,N_3270,N_4475);
and U4801 (N_4801,N_3763,N_4260);
nor U4802 (N_4802,N_4011,N_3343);
xor U4803 (N_4803,N_3809,N_3912);
xnor U4804 (N_4804,N_4265,N_4024);
xor U4805 (N_4805,N_3013,N_4043);
xnor U4806 (N_4806,N_3286,N_3689);
nor U4807 (N_4807,N_3153,N_3711);
or U4808 (N_4808,N_3506,N_3320);
nor U4809 (N_4809,N_4482,N_3055);
nand U4810 (N_4810,N_4361,N_3273);
nand U4811 (N_4811,N_3181,N_4130);
xor U4812 (N_4812,N_4388,N_3822);
nor U4813 (N_4813,N_3666,N_3817);
nor U4814 (N_4814,N_4079,N_4247);
or U4815 (N_4815,N_4339,N_3233);
nor U4816 (N_4816,N_3667,N_3340);
nor U4817 (N_4817,N_3370,N_3648);
and U4818 (N_4818,N_3307,N_3895);
and U4819 (N_4819,N_3877,N_4205);
xor U4820 (N_4820,N_3569,N_3549);
xnor U4821 (N_4821,N_3606,N_3862);
nor U4822 (N_4822,N_3979,N_3230);
or U4823 (N_4823,N_4009,N_3427);
nor U4824 (N_4824,N_3567,N_4283);
and U4825 (N_4825,N_4394,N_3002);
or U4826 (N_4826,N_3334,N_3704);
nand U4827 (N_4827,N_3244,N_3845);
nand U4828 (N_4828,N_3366,N_4357);
nor U4829 (N_4829,N_3130,N_4491);
nor U4830 (N_4830,N_3371,N_4305);
nor U4831 (N_4831,N_4116,N_3633);
nand U4832 (N_4832,N_3360,N_4192);
or U4833 (N_4833,N_4197,N_3503);
nand U4834 (N_4834,N_3252,N_3858);
nand U4835 (N_4835,N_4301,N_3814);
xor U4836 (N_4836,N_3263,N_4030);
or U4837 (N_4837,N_4443,N_3011);
or U4838 (N_4838,N_3076,N_3235);
xnor U4839 (N_4839,N_4322,N_3253);
and U4840 (N_4840,N_4263,N_3162);
nor U4841 (N_4841,N_3777,N_3009);
nand U4842 (N_4842,N_3333,N_3968);
and U4843 (N_4843,N_3958,N_3326);
and U4844 (N_4844,N_4145,N_3778);
nand U4845 (N_4845,N_3044,N_4128);
nor U4846 (N_4846,N_3592,N_3500);
nand U4847 (N_4847,N_4143,N_3706);
nand U4848 (N_4848,N_4139,N_4284);
or U4849 (N_4849,N_3998,N_4402);
or U4850 (N_4850,N_3186,N_4164);
xnor U4851 (N_4851,N_4085,N_3659);
and U4852 (N_4852,N_3319,N_3967);
nor U4853 (N_4853,N_3124,N_4296);
xnor U4854 (N_4854,N_3993,N_3473);
xnor U4855 (N_4855,N_4445,N_3740);
nor U4856 (N_4856,N_4371,N_4174);
nand U4857 (N_4857,N_4142,N_4172);
or U4858 (N_4858,N_3810,N_4450);
and U4859 (N_4859,N_3696,N_3544);
or U4860 (N_4860,N_3113,N_4051);
nand U4861 (N_4861,N_3100,N_3674);
or U4862 (N_4862,N_3172,N_3746);
nor U4863 (N_4863,N_3670,N_4005);
nor U4864 (N_4864,N_3931,N_3391);
nand U4865 (N_4865,N_3470,N_4094);
nor U4866 (N_4866,N_3758,N_3908);
or U4867 (N_4867,N_3878,N_4295);
nor U4868 (N_4868,N_3066,N_4211);
xnor U4869 (N_4869,N_3726,N_3165);
nand U4870 (N_4870,N_3377,N_3597);
or U4871 (N_4871,N_3780,N_3378);
and U4872 (N_4872,N_4431,N_3478);
xor U4873 (N_4873,N_4041,N_3487);
xnor U4874 (N_4874,N_3242,N_3512);
xor U4875 (N_4875,N_3114,N_4337);
xor U4876 (N_4876,N_3407,N_3437);
nand U4877 (N_4877,N_4362,N_3855);
or U4878 (N_4878,N_3856,N_4313);
or U4879 (N_4879,N_4216,N_3209);
nand U4880 (N_4880,N_4003,N_3232);
nor U4881 (N_4881,N_3893,N_3556);
nand U4882 (N_4882,N_3602,N_4365);
xnor U4883 (N_4883,N_3760,N_3509);
nor U4884 (N_4884,N_3059,N_3183);
xor U4885 (N_4885,N_4466,N_3922);
or U4886 (N_4886,N_3518,N_3959);
or U4887 (N_4887,N_3946,N_3944);
or U4888 (N_4888,N_3228,N_4280);
xor U4889 (N_4889,N_4163,N_4156);
xor U4890 (N_4890,N_3710,N_3545);
or U4891 (N_4891,N_3404,N_3642);
or U4892 (N_4892,N_3504,N_3189);
nand U4893 (N_4893,N_3152,N_3006);
nor U4894 (N_4894,N_3776,N_3703);
and U4895 (N_4895,N_4220,N_3934);
or U4896 (N_4896,N_4414,N_4455);
nor U4897 (N_4897,N_3480,N_4473);
or U4898 (N_4898,N_4451,N_3978);
and U4899 (N_4899,N_4294,N_3669);
and U4900 (N_4900,N_3091,N_3354);
nand U4901 (N_4901,N_4324,N_3916);
xor U4902 (N_4902,N_3582,N_3374);
or U4903 (N_4903,N_4291,N_3923);
nand U4904 (N_4904,N_3848,N_3843);
nand U4905 (N_4905,N_3889,N_4438);
and U4906 (N_4906,N_4352,N_3079);
nand U4907 (N_4907,N_3805,N_3464);
xnor U4908 (N_4908,N_3146,N_3783);
xnor U4909 (N_4909,N_4014,N_3577);
xnor U4910 (N_4910,N_4351,N_4276);
xor U4911 (N_4911,N_3297,N_3375);
nand U4912 (N_4912,N_3695,N_3520);
nand U4913 (N_4913,N_4020,N_3037);
nor U4914 (N_4914,N_3484,N_4036);
and U4915 (N_4915,N_3950,N_4096);
xor U4916 (N_4916,N_3825,N_4107);
nand U4917 (N_4917,N_4032,N_3469);
xnor U4918 (N_4918,N_3345,N_3144);
and U4919 (N_4919,N_3983,N_3994);
or U4920 (N_4920,N_3621,N_3132);
or U4921 (N_4921,N_3034,N_3444);
nor U4922 (N_4922,N_3644,N_3649);
nor U4923 (N_4923,N_3846,N_3430);
or U4924 (N_4924,N_3872,N_4208);
and U4925 (N_4925,N_3475,N_3104);
or U4926 (N_4926,N_3243,N_3361);
or U4927 (N_4927,N_4487,N_4336);
nor U4928 (N_4928,N_4149,N_3885);
or U4929 (N_4929,N_3989,N_4428);
or U4930 (N_4930,N_4363,N_3782);
nor U4931 (N_4931,N_3202,N_3128);
xnor U4932 (N_4932,N_3615,N_3864);
and U4933 (N_4933,N_4093,N_3485);
or U4934 (N_4934,N_3705,N_3921);
or U4935 (N_4935,N_3190,N_3571);
xnor U4936 (N_4936,N_3755,N_3781);
xor U4937 (N_4937,N_3775,N_3211);
or U4938 (N_4938,N_3408,N_4398);
and U4939 (N_4939,N_3174,N_3227);
nor U4940 (N_4940,N_4039,N_3730);
nand U4941 (N_4941,N_3564,N_3168);
nand U4942 (N_4942,N_4331,N_3786);
or U4943 (N_4943,N_4167,N_3388);
xor U4944 (N_4944,N_3080,N_4316);
nand U4945 (N_4945,N_4479,N_3212);
nand U4946 (N_4946,N_3351,N_4405);
or U4947 (N_4947,N_3287,N_3356);
nand U4948 (N_4948,N_3562,N_4285);
or U4949 (N_4949,N_3627,N_4155);
or U4950 (N_4950,N_3508,N_3105);
and U4951 (N_4951,N_4158,N_4202);
xnor U4952 (N_4952,N_4373,N_4081);
and U4953 (N_4953,N_3036,N_4302);
xor U4954 (N_4954,N_3295,N_3180);
and U4955 (N_4955,N_3533,N_3457);
and U4956 (N_4956,N_3260,N_3821);
and U4957 (N_4957,N_3075,N_3409);
or U4958 (N_4958,N_3839,N_4221);
nand U4959 (N_4959,N_3827,N_4499);
xnor U4960 (N_4960,N_3892,N_3974);
xor U4961 (N_4961,N_4432,N_3458);
and U4962 (N_4962,N_3357,N_4293);
or U4963 (N_4963,N_4498,N_3268);
xor U4964 (N_4964,N_4141,N_3266);
xnor U4965 (N_4965,N_3583,N_3847);
or U4966 (N_4966,N_3547,N_4198);
or U4967 (N_4967,N_3622,N_3987);
and U4968 (N_4968,N_3552,N_3739);
nand U4969 (N_4969,N_3175,N_3208);
nor U4970 (N_4970,N_4029,N_3972);
nand U4971 (N_4971,N_4227,N_4175);
xor U4972 (N_4972,N_3173,N_4231);
nand U4973 (N_4973,N_4459,N_4080);
and U4974 (N_4974,N_3435,N_3335);
xor U4975 (N_4975,N_3962,N_4073);
and U4976 (N_4976,N_3961,N_3401);
nor U4977 (N_4977,N_3223,N_3386);
xor U4978 (N_4978,N_3010,N_3121);
and U4979 (N_4979,N_3465,N_4040);
nand U4980 (N_4980,N_3008,N_4138);
nor U4981 (N_4981,N_3155,N_3102);
and U4982 (N_4982,N_4484,N_3099);
nand U4983 (N_4983,N_3416,N_4448);
and U4984 (N_4984,N_3539,N_3205);
and U4985 (N_4985,N_4406,N_4460);
and U4986 (N_4986,N_4047,N_3653);
nor U4987 (N_4987,N_3302,N_3241);
and U4988 (N_4988,N_3342,N_4307);
xnor U4989 (N_4989,N_4372,N_3454);
nor U4990 (N_4990,N_3284,N_4253);
nor U4991 (N_4991,N_3101,N_3293);
nand U4992 (N_4992,N_4179,N_4377);
or U4993 (N_4993,N_3259,N_3899);
and U4994 (N_4994,N_3884,N_4144);
xnor U4995 (N_4995,N_3399,N_3671);
nand U4996 (N_4996,N_3216,N_3074);
nand U4997 (N_4997,N_3502,N_3309);
nand U4998 (N_4998,N_4021,N_3522);
nor U4999 (N_4999,N_3283,N_3021);
and U5000 (N_5000,N_3047,N_3448);
and U5001 (N_5001,N_3584,N_3643);
and U5002 (N_5002,N_3524,N_4476);
nor U5003 (N_5003,N_3501,N_3089);
and U5004 (N_5004,N_3379,N_4430);
or U5005 (N_5005,N_3039,N_3352);
nand U5006 (N_5006,N_3403,N_3110);
nand U5007 (N_5007,N_3122,N_3660);
nand U5008 (N_5008,N_3970,N_4481);
nand U5009 (N_5009,N_3801,N_3192);
xor U5010 (N_5010,N_4129,N_3925);
or U5011 (N_5011,N_3324,N_3027);
nor U5012 (N_5012,N_4350,N_4367);
and U5013 (N_5013,N_3056,N_4369);
and U5014 (N_5014,N_3992,N_3038);
xor U5015 (N_5015,N_3141,N_3764);
or U5016 (N_5016,N_3199,N_3587);
or U5017 (N_5017,N_3262,N_3698);
nor U5018 (N_5018,N_4408,N_4364);
nand U5019 (N_5019,N_3536,N_3960);
xnor U5020 (N_5020,N_4309,N_3541);
xor U5021 (N_5021,N_3543,N_3145);
or U5022 (N_5022,N_3098,N_3171);
xor U5023 (N_5023,N_4071,N_3115);
or U5024 (N_5024,N_3442,N_3640);
and U5025 (N_5025,N_3812,N_3727);
nand U5026 (N_5026,N_4210,N_4486);
xnor U5027 (N_5027,N_4188,N_3394);
nor U5028 (N_5028,N_3939,N_3398);
and U5029 (N_5029,N_4026,N_4334);
or U5030 (N_5030,N_3217,N_4453);
or U5031 (N_5031,N_4219,N_4349);
or U5032 (N_5032,N_3528,N_3697);
and U5033 (N_5033,N_3514,N_4070);
xor U5034 (N_5034,N_3586,N_3306);
or U5035 (N_5035,N_4214,N_4180);
nor U5036 (N_5036,N_4492,N_4224);
nor U5037 (N_5037,N_4474,N_3425);
xor U5038 (N_5038,N_4061,N_4478);
nand U5039 (N_5039,N_3405,N_3919);
xnor U5040 (N_5040,N_3341,N_4391);
xnor U5041 (N_5041,N_3686,N_3107);
or U5042 (N_5042,N_3555,N_4173);
and U5043 (N_5043,N_3251,N_3143);
xor U5044 (N_5044,N_3792,N_3077);
nand U5045 (N_5045,N_3346,N_3288);
nand U5046 (N_5046,N_4160,N_4207);
nand U5047 (N_5047,N_3871,N_3820);
and U5048 (N_5048,N_4384,N_4105);
or U5049 (N_5049,N_3050,N_4018);
xor U5050 (N_5050,N_4028,N_3851);
nor U5051 (N_5051,N_3071,N_3661);
xor U5052 (N_5052,N_3300,N_3490);
nand U5053 (N_5053,N_3658,N_3510);
nor U5054 (N_5054,N_4440,N_4184);
and U5055 (N_5055,N_4189,N_3699);
or U5056 (N_5056,N_3647,N_4442);
or U5057 (N_5057,N_3677,N_3133);
and U5058 (N_5058,N_3019,N_3734);
and U5059 (N_5059,N_3138,N_4104);
xnor U5060 (N_5060,N_3355,N_3579);
or U5061 (N_5061,N_3431,N_4199);
or U5062 (N_5062,N_3865,N_3634);
nor U5063 (N_5063,N_4019,N_4370);
and U5064 (N_5064,N_3331,N_3139);
nor U5065 (N_5065,N_3163,N_3441);
and U5066 (N_5066,N_3542,N_3365);
nand U5067 (N_5067,N_3396,N_3662);
xor U5068 (N_5068,N_3225,N_4320);
xnor U5069 (N_5069,N_4489,N_3095);
nor U5070 (N_5070,N_4117,N_3905);
nand U5071 (N_5071,N_3638,N_3466);
nand U5072 (N_5072,N_4066,N_3116);
and U5073 (N_5073,N_3134,N_4426);
nand U5074 (N_5074,N_4289,N_4380);
or U5075 (N_5075,N_3605,N_3272);
or U5076 (N_5076,N_4493,N_3016);
nor U5077 (N_5077,N_3451,N_3453);
nor U5078 (N_5078,N_3868,N_3033);
or U5079 (N_5079,N_4099,N_3625);
and U5080 (N_5080,N_3459,N_4354);
and U5081 (N_5081,N_4275,N_4162);
xnor U5082 (N_5082,N_3766,N_4254);
and U5083 (N_5083,N_4434,N_4248);
and U5084 (N_5084,N_3854,N_3250);
and U5085 (N_5085,N_4326,N_4236);
and U5086 (N_5086,N_3178,N_3853);
nor U5087 (N_5087,N_3219,N_3824);
xnor U5088 (N_5088,N_4273,N_3150);
nor U5089 (N_5089,N_3718,N_3741);
or U5090 (N_5090,N_3725,N_4407);
xnor U5091 (N_5091,N_3743,N_4379);
xor U5092 (N_5092,N_3953,N_4120);
nand U5093 (N_5093,N_3645,N_3609);
nor U5094 (N_5094,N_3004,N_3808);
and U5095 (N_5095,N_3271,N_3068);
nand U5096 (N_5096,N_4076,N_3018);
nor U5097 (N_5097,N_3135,N_3948);
xnor U5098 (N_5098,N_3626,N_3194);
or U5099 (N_5099,N_3481,N_3559);
nor U5100 (N_5100,N_4311,N_4223);
or U5101 (N_5101,N_3106,N_4355);
and U5102 (N_5102,N_3863,N_4195);
and U5103 (N_5103,N_3264,N_3296);
nand U5104 (N_5104,N_3769,N_4257);
xor U5105 (N_5105,N_3869,N_4325);
and U5106 (N_5106,N_4274,N_3947);
nor U5107 (N_5107,N_4063,N_3043);
xor U5108 (N_5108,N_4423,N_4209);
xor U5109 (N_5109,N_4327,N_3088);
nand U5110 (N_5110,N_3986,N_3751);
nor U5111 (N_5111,N_3433,N_3007);
nand U5112 (N_5112,N_4127,N_4131);
nand U5113 (N_5113,N_4132,N_3064);
nor U5114 (N_5114,N_3325,N_3876);
nor U5115 (N_5115,N_3942,N_4390);
and U5116 (N_5116,N_3799,N_4437);
nor U5117 (N_5117,N_4356,N_4062);
nor U5118 (N_5118,N_3926,N_4464);
xnor U5119 (N_5119,N_3445,N_3381);
and U5120 (N_5120,N_4075,N_3956);
nand U5121 (N_5121,N_3999,N_3014);
xnor U5122 (N_5122,N_4393,N_3198);
xnor U5123 (N_5123,N_4001,N_3527);
xnor U5124 (N_5124,N_3197,N_3329);
xnor U5125 (N_5125,N_4277,N_3418);
xor U5126 (N_5126,N_4343,N_3156);
xor U5127 (N_5127,N_3234,N_4058);
or U5128 (N_5128,N_3069,N_4306);
or U5129 (N_5129,N_4310,N_4234);
xnor U5130 (N_5130,N_3593,N_3291);
xnor U5131 (N_5131,N_4228,N_4200);
xnor U5132 (N_5132,N_3460,N_4125);
and U5133 (N_5133,N_3452,N_4042);
nand U5134 (N_5134,N_3788,N_3596);
and U5135 (N_5135,N_3920,N_3447);
nor U5136 (N_5136,N_3060,N_3362);
nand U5137 (N_5137,N_4235,N_3112);
or U5138 (N_5138,N_3897,N_4121);
xnor U5139 (N_5139,N_3575,N_3256);
xor U5140 (N_5140,N_3318,N_4447);
xnor U5141 (N_5141,N_3613,N_3290);
xor U5142 (N_5142,N_3312,N_3767);
nand U5143 (N_5143,N_4472,N_3570);
nand U5144 (N_5144,N_4084,N_4101);
or U5145 (N_5145,N_3035,N_3449);
nor U5146 (N_5146,N_3888,N_3833);
nand U5147 (N_5147,N_3652,N_3997);
or U5148 (N_5148,N_3977,N_3985);
xor U5149 (N_5149,N_3768,N_3672);
nor U5150 (N_5150,N_3618,N_3337);
xnor U5151 (N_5151,N_4191,N_4245);
xor U5152 (N_5152,N_3723,N_3411);
nand U5153 (N_5153,N_3752,N_3941);
xor U5154 (N_5154,N_4206,N_4161);
nand U5155 (N_5155,N_3421,N_3608);
xor U5156 (N_5156,N_4237,N_3206);
and U5157 (N_5157,N_4287,N_3969);
or U5158 (N_5158,N_4240,N_3551);
and U5159 (N_5159,N_3483,N_3129);
xnor U5160 (N_5160,N_3117,N_3392);
and U5161 (N_5161,N_3620,N_4053);
nor U5162 (N_5162,N_3675,N_3429);
nor U5163 (N_5163,N_3151,N_3838);
and U5164 (N_5164,N_4262,N_3742);
and U5165 (N_5165,N_4251,N_4456);
and U5166 (N_5166,N_3438,N_4452);
nand U5167 (N_5167,N_3412,N_4059);
or U5168 (N_5168,N_4091,N_3913);
nor U5169 (N_5169,N_3193,N_3275);
nand U5170 (N_5170,N_4279,N_3610);
xnor U5171 (N_5171,N_3823,N_3213);
or U5172 (N_5172,N_3304,N_3685);
nor U5173 (N_5173,N_4468,N_3170);
nand U5174 (N_5174,N_3874,N_3852);
xor U5175 (N_5175,N_3491,N_3732);
xnor U5176 (N_5176,N_3424,N_3499);
and U5177 (N_5177,N_4249,N_3668);
or U5178 (N_5178,N_3599,N_3367);
xor U5179 (N_5179,N_3224,N_3092);
and U5180 (N_5180,N_3588,N_3521);
nor U5181 (N_5181,N_4046,N_3612);
and U5182 (N_5182,N_3278,N_3943);
nand U5183 (N_5183,N_3757,N_4278);
xor U5184 (N_5184,N_4154,N_3707);
nor U5185 (N_5185,N_3601,N_4095);
or U5186 (N_5186,N_4297,N_3655);
or U5187 (N_5187,N_3359,N_3700);
nand U5188 (N_5188,N_3236,N_4261);
nand U5189 (N_5189,N_4092,N_3772);
nand U5190 (N_5190,N_3516,N_3826);
or U5191 (N_5191,N_4124,N_3576);
xor U5192 (N_5192,N_3203,N_3393);
nand U5193 (N_5193,N_4470,N_3937);
or U5194 (N_5194,N_4100,N_3269);
or U5195 (N_5195,N_3673,N_3282);
and U5196 (N_5196,N_4225,N_3338);
nand U5197 (N_5197,N_3159,N_3787);
xnor U5198 (N_5198,N_4023,N_3731);
and U5199 (N_5199,N_3654,N_4332);
xnor U5200 (N_5200,N_4054,N_3210);
nor U5201 (N_5201,N_3315,N_3728);
nand U5202 (N_5202,N_3032,N_4366);
nor U5203 (N_5203,N_3507,N_3687);
xnor U5204 (N_5204,N_3486,N_3566);
nor U5205 (N_5205,N_3410,N_4010);
nor U5206 (N_5206,N_4480,N_4169);
nand U5207 (N_5207,N_3492,N_3191);
or U5208 (N_5208,N_3639,N_4185);
xnor U5209 (N_5209,N_4303,N_4037);
xor U5210 (N_5210,N_4422,N_4385);
or U5211 (N_5211,N_3831,N_3713);
or U5212 (N_5212,N_4397,N_4299);
xor U5213 (N_5213,N_3090,N_4318);
and U5214 (N_5214,N_3467,N_3182);
xor U5215 (N_5215,N_3641,N_4467);
or U5216 (N_5216,N_4465,N_3866);
or U5217 (N_5217,N_3717,N_4383);
xor U5218 (N_5218,N_4420,N_3436);
xnor U5219 (N_5219,N_3911,N_3756);
or U5220 (N_5220,N_4497,N_3712);
or U5221 (N_5221,N_3281,N_4151);
or U5222 (N_5222,N_3976,N_3749);
and U5223 (N_5223,N_4045,N_3058);
and U5224 (N_5224,N_3221,N_4454);
nand U5225 (N_5225,N_4136,N_4013);
or U5226 (N_5226,N_3446,N_3395);
and U5227 (N_5227,N_3336,N_3382);
or U5228 (N_5228,N_4238,N_3917);
nor U5229 (N_5229,N_3048,N_3332);
or U5230 (N_5230,N_3305,N_3750);
or U5231 (N_5231,N_3489,N_3073);
nor U5232 (N_5232,N_3497,N_3308);
nor U5233 (N_5233,N_3456,N_3965);
nand U5234 (N_5234,N_4025,N_3774);
xor U5235 (N_5235,N_3261,N_3656);
nand U5236 (N_5236,N_3759,N_3554);
xor U5237 (N_5237,N_4000,N_4233);
nand U5238 (N_5238,N_3417,N_4392);
nand U5239 (N_5239,N_3881,N_3523);
or U5240 (N_5240,N_3000,N_3493);
or U5241 (N_5241,N_3389,N_3330);
nand U5242 (N_5242,N_3495,N_3910);
and U5243 (N_5243,N_4108,N_4387);
nand U5244 (N_5244,N_3339,N_4457);
and U5245 (N_5245,N_3929,N_3971);
nand U5246 (N_5246,N_3443,N_3052);
and U5247 (N_5247,N_4078,N_3434);
and U5248 (N_5248,N_3716,N_3572);
nor U5249 (N_5249,N_3136,N_3419);
and U5250 (N_5250,N_3892,N_3391);
and U5251 (N_5251,N_3789,N_4262);
and U5252 (N_5252,N_3450,N_3487);
and U5253 (N_5253,N_3537,N_4377);
nor U5254 (N_5254,N_3591,N_3266);
nor U5255 (N_5255,N_3532,N_3340);
xor U5256 (N_5256,N_3309,N_3536);
nor U5257 (N_5257,N_3436,N_4024);
nand U5258 (N_5258,N_3485,N_3326);
or U5259 (N_5259,N_3343,N_3934);
or U5260 (N_5260,N_4302,N_3116);
xnor U5261 (N_5261,N_4052,N_4258);
nor U5262 (N_5262,N_3788,N_3766);
xnor U5263 (N_5263,N_3858,N_3661);
nand U5264 (N_5264,N_3591,N_4356);
nor U5265 (N_5265,N_3234,N_3643);
and U5266 (N_5266,N_3563,N_3348);
nor U5267 (N_5267,N_4463,N_3836);
or U5268 (N_5268,N_4336,N_3916);
nand U5269 (N_5269,N_3690,N_3725);
or U5270 (N_5270,N_4413,N_3406);
nor U5271 (N_5271,N_3434,N_4457);
or U5272 (N_5272,N_3750,N_3334);
or U5273 (N_5273,N_3692,N_3776);
nand U5274 (N_5274,N_3469,N_4250);
and U5275 (N_5275,N_3269,N_4164);
and U5276 (N_5276,N_4438,N_3958);
nand U5277 (N_5277,N_3350,N_3928);
and U5278 (N_5278,N_4261,N_3655);
and U5279 (N_5279,N_4069,N_4246);
and U5280 (N_5280,N_3577,N_3649);
xnor U5281 (N_5281,N_3001,N_3275);
nor U5282 (N_5282,N_4225,N_3817);
nor U5283 (N_5283,N_3564,N_4306);
or U5284 (N_5284,N_3847,N_4326);
or U5285 (N_5285,N_3925,N_3450);
nand U5286 (N_5286,N_4230,N_3512);
nor U5287 (N_5287,N_3362,N_3108);
or U5288 (N_5288,N_3723,N_3936);
or U5289 (N_5289,N_3920,N_4011);
nor U5290 (N_5290,N_3602,N_3863);
or U5291 (N_5291,N_4114,N_4110);
nand U5292 (N_5292,N_3476,N_4276);
nor U5293 (N_5293,N_3519,N_4127);
nor U5294 (N_5294,N_3469,N_3501);
nand U5295 (N_5295,N_3287,N_4364);
or U5296 (N_5296,N_4065,N_3130);
and U5297 (N_5297,N_3357,N_4260);
and U5298 (N_5298,N_4161,N_3513);
nor U5299 (N_5299,N_3768,N_4144);
and U5300 (N_5300,N_3088,N_3545);
nor U5301 (N_5301,N_4067,N_4261);
and U5302 (N_5302,N_3058,N_3191);
xor U5303 (N_5303,N_3801,N_4380);
nor U5304 (N_5304,N_4103,N_4119);
and U5305 (N_5305,N_3764,N_3664);
xnor U5306 (N_5306,N_4380,N_3954);
and U5307 (N_5307,N_3473,N_3080);
nor U5308 (N_5308,N_3229,N_3309);
and U5309 (N_5309,N_4039,N_4487);
and U5310 (N_5310,N_3889,N_3746);
or U5311 (N_5311,N_4144,N_3996);
xor U5312 (N_5312,N_3300,N_4250);
xor U5313 (N_5313,N_3745,N_3787);
or U5314 (N_5314,N_3269,N_4340);
nor U5315 (N_5315,N_3653,N_3670);
and U5316 (N_5316,N_3515,N_4446);
xor U5317 (N_5317,N_3974,N_3025);
or U5318 (N_5318,N_3195,N_3971);
xnor U5319 (N_5319,N_3107,N_3470);
nor U5320 (N_5320,N_3598,N_3324);
and U5321 (N_5321,N_3836,N_4329);
nor U5322 (N_5322,N_3384,N_3981);
nor U5323 (N_5323,N_4228,N_3956);
or U5324 (N_5324,N_3045,N_3501);
xnor U5325 (N_5325,N_4249,N_3257);
xnor U5326 (N_5326,N_4463,N_4156);
nor U5327 (N_5327,N_3341,N_4006);
and U5328 (N_5328,N_3967,N_4307);
or U5329 (N_5329,N_3387,N_3083);
nand U5330 (N_5330,N_3575,N_3227);
and U5331 (N_5331,N_3648,N_3306);
xor U5332 (N_5332,N_3075,N_3937);
nor U5333 (N_5333,N_3543,N_4053);
xnor U5334 (N_5334,N_3382,N_3209);
or U5335 (N_5335,N_3543,N_3584);
xor U5336 (N_5336,N_4246,N_3357);
or U5337 (N_5337,N_3567,N_4170);
xnor U5338 (N_5338,N_3025,N_3805);
and U5339 (N_5339,N_3323,N_3341);
nor U5340 (N_5340,N_3982,N_4310);
or U5341 (N_5341,N_3404,N_4072);
and U5342 (N_5342,N_3877,N_4065);
xnor U5343 (N_5343,N_4350,N_4457);
or U5344 (N_5344,N_3243,N_4088);
or U5345 (N_5345,N_4138,N_3659);
xor U5346 (N_5346,N_4124,N_4093);
nand U5347 (N_5347,N_4188,N_3460);
nand U5348 (N_5348,N_3868,N_4041);
nand U5349 (N_5349,N_4414,N_4410);
nand U5350 (N_5350,N_3350,N_3029);
xor U5351 (N_5351,N_3129,N_3855);
nand U5352 (N_5352,N_3041,N_4125);
nand U5353 (N_5353,N_3106,N_3318);
nand U5354 (N_5354,N_4487,N_4321);
nor U5355 (N_5355,N_3732,N_3145);
or U5356 (N_5356,N_4118,N_4344);
or U5357 (N_5357,N_3268,N_3778);
xor U5358 (N_5358,N_4199,N_4175);
nand U5359 (N_5359,N_3660,N_3686);
xor U5360 (N_5360,N_4361,N_4465);
or U5361 (N_5361,N_3073,N_3423);
xnor U5362 (N_5362,N_3257,N_3843);
or U5363 (N_5363,N_3715,N_3244);
nand U5364 (N_5364,N_3784,N_3881);
and U5365 (N_5365,N_3148,N_4249);
and U5366 (N_5366,N_3381,N_3704);
nor U5367 (N_5367,N_3724,N_3686);
and U5368 (N_5368,N_3704,N_4476);
xor U5369 (N_5369,N_3241,N_3865);
nor U5370 (N_5370,N_4113,N_3156);
xnor U5371 (N_5371,N_3783,N_3245);
or U5372 (N_5372,N_3267,N_3055);
nor U5373 (N_5373,N_4020,N_4090);
or U5374 (N_5374,N_4096,N_3544);
nand U5375 (N_5375,N_3676,N_3932);
nand U5376 (N_5376,N_3926,N_4053);
and U5377 (N_5377,N_3772,N_3606);
xnor U5378 (N_5378,N_4131,N_3820);
nor U5379 (N_5379,N_3977,N_3079);
and U5380 (N_5380,N_3354,N_3965);
nor U5381 (N_5381,N_3508,N_3849);
xor U5382 (N_5382,N_4339,N_3687);
xor U5383 (N_5383,N_3820,N_3814);
and U5384 (N_5384,N_3302,N_4074);
and U5385 (N_5385,N_3857,N_3564);
and U5386 (N_5386,N_4376,N_3187);
and U5387 (N_5387,N_3597,N_3006);
nand U5388 (N_5388,N_3086,N_4367);
xor U5389 (N_5389,N_3943,N_4320);
xnor U5390 (N_5390,N_3689,N_3679);
or U5391 (N_5391,N_3213,N_4426);
nand U5392 (N_5392,N_3892,N_4271);
or U5393 (N_5393,N_4144,N_3968);
nand U5394 (N_5394,N_3387,N_3179);
and U5395 (N_5395,N_4346,N_3801);
and U5396 (N_5396,N_3475,N_3510);
or U5397 (N_5397,N_4326,N_4377);
and U5398 (N_5398,N_3527,N_3011);
nor U5399 (N_5399,N_3212,N_3498);
and U5400 (N_5400,N_4389,N_3480);
xnor U5401 (N_5401,N_3635,N_3822);
and U5402 (N_5402,N_3598,N_4367);
nor U5403 (N_5403,N_3570,N_4355);
nand U5404 (N_5404,N_3482,N_3008);
or U5405 (N_5405,N_3439,N_3720);
nand U5406 (N_5406,N_3530,N_3098);
nor U5407 (N_5407,N_4338,N_4332);
and U5408 (N_5408,N_3197,N_3416);
xnor U5409 (N_5409,N_3347,N_3154);
and U5410 (N_5410,N_3519,N_3860);
and U5411 (N_5411,N_3299,N_3723);
nand U5412 (N_5412,N_3250,N_3282);
xnor U5413 (N_5413,N_4083,N_3116);
and U5414 (N_5414,N_3846,N_3532);
nand U5415 (N_5415,N_3493,N_3238);
xor U5416 (N_5416,N_3185,N_4099);
and U5417 (N_5417,N_4335,N_3595);
nor U5418 (N_5418,N_3672,N_4198);
or U5419 (N_5419,N_3959,N_3364);
nor U5420 (N_5420,N_4359,N_4421);
nand U5421 (N_5421,N_4248,N_3066);
nand U5422 (N_5422,N_4024,N_3869);
or U5423 (N_5423,N_4162,N_4105);
nor U5424 (N_5424,N_3884,N_3432);
and U5425 (N_5425,N_3498,N_3897);
or U5426 (N_5426,N_3355,N_3114);
nor U5427 (N_5427,N_3236,N_3621);
or U5428 (N_5428,N_3927,N_4494);
and U5429 (N_5429,N_3394,N_3423);
and U5430 (N_5430,N_3398,N_3216);
and U5431 (N_5431,N_3881,N_4051);
or U5432 (N_5432,N_4089,N_4454);
xor U5433 (N_5433,N_3411,N_4351);
or U5434 (N_5434,N_3351,N_3034);
xnor U5435 (N_5435,N_4184,N_3336);
and U5436 (N_5436,N_3750,N_3939);
and U5437 (N_5437,N_4483,N_4375);
and U5438 (N_5438,N_3893,N_4149);
xnor U5439 (N_5439,N_3113,N_3264);
nor U5440 (N_5440,N_3556,N_4314);
or U5441 (N_5441,N_4486,N_3578);
xnor U5442 (N_5442,N_3093,N_3125);
xnor U5443 (N_5443,N_4172,N_3993);
xor U5444 (N_5444,N_4308,N_3777);
nor U5445 (N_5445,N_4078,N_3744);
nand U5446 (N_5446,N_3124,N_3454);
xor U5447 (N_5447,N_4220,N_3006);
nor U5448 (N_5448,N_3304,N_3075);
nand U5449 (N_5449,N_3858,N_3202);
or U5450 (N_5450,N_4411,N_4416);
nor U5451 (N_5451,N_4455,N_3623);
xnor U5452 (N_5452,N_3158,N_4080);
or U5453 (N_5453,N_3521,N_3564);
or U5454 (N_5454,N_3136,N_3794);
and U5455 (N_5455,N_3469,N_4360);
or U5456 (N_5456,N_3929,N_3638);
or U5457 (N_5457,N_3984,N_4208);
nand U5458 (N_5458,N_4070,N_3906);
or U5459 (N_5459,N_3876,N_4401);
or U5460 (N_5460,N_4161,N_4279);
and U5461 (N_5461,N_3726,N_3095);
nand U5462 (N_5462,N_3044,N_4224);
xnor U5463 (N_5463,N_3745,N_3133);
and U5464 (N_5464,N_4153,N_4261);
or U5465 (N_5465,N_3122,N_3694);
xnor U5466 (N_5466,N_3170,N_4086);
nor U5467 (N_5467,N_4127,N_3328);
xor U5468 (N_5468,N_4495,N_3946);
nor U5469 (N_5469,N_3160,N_3702);
xnor U5470 (N_5470,N_3679,N_4266);
nand U5471 (N_5471,N_3626,N_4321);
xor U5472 (N_5472,N_4355,N_4121);
and U5473 (N_5473,N_3103,N_3226);
nor U5474 (N_5474,N_3182,N_3764);
nor U5475 (N_5475,N_3389,N_3774);
nand U5476 (N_5476,N_3628,N_4199);
nand U5477 (N_5477,N_3034,N_4219);
or U5478 (N_5478,N_4048,N_3892);
or U5479 (N_5479,N_4031,N_3052);
and U5480 (N_5480,N_3060,N_3975);
or U5481 (N_5481,N_3142,N_3148);
xor U5482 (N_5482,N_3898,N_4138);
and U5483 (N_5483,N_3083,N_4490);
xor U5484 (N_5484,N_4044,N_3444);
nor U5485 (N_5485,N_4010,N_3294);
or U5486 (N_5486,N_3306,N_3765);
xor U5487 (N_5487,N_3689,N_3307);
nand U5488 (N_5488,N_4277,N_4190);
xnor U5489 (N_5489,N_4268,N_3466);
or U5490 (N_5490,N_3526,N_3150);
xnor U5491 (N_5491,N_3748,N_3341);
nand U5492 (N_5492,N_3456,N_3413);
nor U5493 (N_5493,N_3492,N_3649);
and U5494 (N_5494,N_4368,N_3505);
nor U5495 (N_5495,N_3595,N_3089);
and U5496 (N_5496,N_3600,N_3580);
and U5497 (N_5497,N_4203,N_4295);
xnor U5498 (N_5498,N_4322,N_3786);
or U5499 (N_5499,N_4136,N_4423);
or U5500 (N_5500,N_4230,N_4403);
xnor U5501 (N_5501,N_3993,N_4038);
xor U5502 (N_5502,N_4485,N_4113);
nand U5503 (N_5503,N_3659,N_3487);
nor U5504 (N_5504,N_3153,N_4183);
xnor U5505 (N_5505,N_3205,N_4257);
nand U5506 (N_5506,N_4259,N_3148);
and U5507 (N_5507,N_4235,N_3438);
or U5508 (N_5508,N_4108,N_3670);
xor U5509 (N_5509,N_3365,N_3599);
xnor U5510 (N_5510,N_3594,N_3603);
or U5511 (N_5511,N_3055,N_3044);
xnor U5512 (N_5512,N_4148,N_3657);
or U5513 (N_5513,N_4334,N_3087);
xnor U5514 (N_5514,N_4188,N_3217);
xnor U5515 (N_5515,N_3682,N_3270);
and U5516 (N_5516,N_3098,N_4064);
xnor U5517 (N_5517,N_3792,N_4196);
nand U5518 (N_5518,N_3685,N_3261);
xnor U5519 (N_5519,N_3595,N_3038);
nand U5520 (N_5520,N_3434,N_3264);
and U5521 (N_5521,N_3033,N_4400);
nor U5522 (N_5522,N_4361,N_3365);
or U5523 (N_5523,N_3372,N_4362);
nand U5524 (N_5524,N_4181,N_3363);
xor U5525 (N_5525,N_3544,N_3353);
nand U5526 (N_5526,N_3947,N_3068);
xor U5527 (N_5527,N_4197,N_3123);
or U5528 (N_5528,N_3241,N_3144);
nand U5529 (N_5529,N_3805,N_3628);
nor U5530 (N_5530,N_4132,N_3066);
nand U5531 (N_5531,N_4057,N_4172);
or U5532 (N_5532,N_4261,N_3150);
or U5533 (N_5533,N_4196,N_3534);
nand U5534 (N_5534,N_3896,N_3660);
nor U5535 (N_5535,N_3061,N_4298);
xnor U5536 (N_5536,N_4120,N_3168);
or U5537 (N_5537,N_4212,N_3440);
nand U5538 (N_5538,N_3007,N_4473);
and U5539 (N_5539,N_3935,N_4353);
xnor U5540 (N_5540,N_3791,N_4168);
nand U5541 (N_5541,N_3127,N_3302);
and U5542 (N_5542,N_3241,N_3767);
xnor U5543 (N_5543,N_3399,N_4216);
nor U5544 (N_5544,N_3310,N_3463);
and U5545 (N_5545,N_3587,N_3741);
xor U5546 (N_5546,N_3237,N_3473);
nand U5547 (N_5547,N_4111,N_3646);
or U5548 (N_5548,N_4134,N_4259);
or U5549 (N_5549,N_4269,N_4101);
or U5550 (N_5550,N_3540,N_4075);
nor U5551 (N_5551,N_3528,N_3609);
nand U5552 (N_5552,N_3012,N_4431);
xnor U5553 (N_5553,N_3139,N_4291);
nand U5554 (N_5554,N_4197,N_3344);
xor U5555 (N_5555,N_3789,N_3363);
or U5556 (N_5556,N_3098,N_3320);
and U5557 (N_5557,N_3036,N_3873);
nand U5558 (N_5558,N_4030,N_3107);
or U5559 (N_5559,N_3393,N_4455);
nor U5560 (N_5560,N_3697,N_4072);
and U5561 (N_5561,N_4449,N_3167);
and U5562 (N_5562,N_3422,N_4269);
or U5563 (N_5563,N_4266,N_3654);
and U5564 (N_5564,N_3260,N_3876);
nor U5565 (N_5565,N_3052,N_4323);
nand U5566 (N_5566,N_4255,N_3871);
and U5567 (N_5567,N_4409,N_3386);
and U5568 (N_5568,N_3333,N_3145);
nor U5569 (N_5569,N_3965,N_4188);
xor U5570 (N_5570,N_3830,N_3597);
xnor U5571 (N_5571,N_3385,N_4433);
nand U5572 (N_5572,N_3767,N_3582);
and U5573 (N_5573,N_3929,N_3670);
or U5574 (N_5574,N_3940,N_4461);
or U5575 (N_5575,N_4016,N_4203);
xor U5576 (N_5576,N_3385,N_3178);
nand U5577 (N_5577,N_4049,N_4163);
nand U5578 (N_5578,N_3623,N_3985);
nor U5579 (N_5579,N_3070,N_3035);
xor U5580 (N_5580,N_3306,N_3515);
xor U5581 (N_5581,N_3275,N_3690);
nand U5582 (N_5582,N_3156,N_3640);
and U5583 (N_5583,N_3345,N_3023);
nor U5584 (N_5584,N_3861,N_4124);
xnor U5585 (N_5585,N_3277,N_4006);
or U5586 (N_5586,N_3401,N_3153);
xor U5587 (N_5587,N_4229,N_3057);
nand U5588 (N_5588,N_3637,N_3533);
and U5589 (N_5589,N_3849,N_4074);
or U5590 (N_5590,N_3298,N_3970);
and U5591 (N_5591,N_3682,N_3649);
nand U5592 (N_5592,N_3396,N_3308);
and U5593 (N_5593,N_4491,N_3414);
or U5594 (N_5594,N_4150,N_3627);
nor U5595 (N_5595,N_3361,N_3476);
or U5596 (N_5596,N_3623,N_3866);
nor U5597 (N_5597,N_4133,N_3326);
or U5598 (N_5598,N_3107,N_3521);
nand U5599 (N_5599,N_3829,N_4323);
nand U5600 (N_5600,N_3995,N_3427);
nor U5601 (N_5601,N_4001,N_3631);
and U5602 (N_5602,N_3957,N_4009);
nor U5603 (N_5603,N_3268,N_3066);
or U5604 (N_5604,N_3342,N_4479);
nand U5605 (N_5605,N_3168,N_3354);
or U5606 (N_5606,N_4233,N_3256);
nor U5607 (N_5607,N_4297,N_3322);
or U5608 (N_5608,N_4149,N_4235);
nand U5609 (N_5609,N_3681,N_3771);
nand U5610 (N_5610,N_4215,N_3544);
nor U5611 (N_5611,N_3186,N_3017);
and U5612 (N_5612,N_3929,N_4063);
nor U5613 (N_5613,N_3728,N_4260);
nand U5614 (N_5614,N_3612,N_4346);
xor U5615 (N_5615,N_3330,N_3258);
xor U5616 (N_5616,N_3646,N_3257);
nor U5617 (N_5617,N_3524,N_3336);
or U5618 (N_5618,N_3117,N_3851);
xnor U5619 (N_5619,N_3666,N_4356);
or U5620 (N_5620,N_3581,N_3601);
and U5621 (N_5621,N_4279,N_3208);
nor U5622 (N_5622,N_4497,N_3358);
and U5623 (N_5623,N_3654,N_4473);
and U5624 (N_5624,N_3399,N_3526);
nor U5625 (N_5625,N_3866,N_3163);
or U5626 (N_5626,N_3569,N_3817);
or U5627 (N_5627,N_4290,N_3338);
and U5628 (N_5628,N_3766,N_4091);
and U5629 (N_5629,N_3154,N_4091);
xor U5630 (N_5630,N_4466,N_3239);
nor U5631 (N_5631,N_3197,N_3315);
nand U5632 (N_5632,N_3397,N_3632);
or U5633 (N_5633,N_3916,N_4086);
and U5634 (N_5634,N_3593,N_3423);
nor U5635 (N_5635,N_3850,N_3297);
and U5636 (N_5636,N_3556,N_4188);
and U5637 (N_5637,N_3717,N_3413);
and U5638 (N_5638,N_3546,N_3312);
xnor U5639 (N_5639,N_3450,N_3472);
xor U5640 (N_5640,N_3445,N_3437);
nand U5641 (N_5641,N_3054,N_3830);
xor U5642 (N_5642,N_3122,N_4449);
and U5643 (N_5643,N_4121,N_3834);
and U5644 (N_5644,N_3684,N_3376);
nor U5645 (N_5645,N_4358,N_3474);
nor U5646 (N_5646,N_3036,N_3115);
xnor U5647 (N_5647,N_3634,N_4444);
nor U5648 (N_5648,N_3231,N_3821);
nor U5649 (N_5649,N_3437,N_4104);
nand U5650 (N_5650,N_3645,N_3581);
or U5651 (N_5651,N_4053,N_4428);
nand U5652 (N_5652,N_4112,N_3096);
nand U5653 (N_5653,N_4232,N_4329);
or U5654 (N_5654,N_4151,N_3577);
nor U5655 (N_5655,N_4425,N_4180);
and U5656 (N_5656,N_3124,N_4463);
nand U5657 (N_5657,N_4096,N_4141);
nor U5658 (N_5658,N_3509,N_4379);
nor U5659 (N_5659,N_3454,N_3058);
xor U5660 (N_5660,N_4033,N_3311);
or U5661 (N_5661,N_3124,N_3806);
nor U5662 (N_5662,N_4111,N_3462);
xor U5663 (N_5663,N_3450,N_4096);
nand U5664 (N_5664,N_3810,N_4249);
nor U5665 (N_5665,N_4299,N_3956);
xnor U5666 (N_5666,N_3626,N_3256);
xnor U5667 (N_5667,N_3189,N_4281);
xnor U5668 (N_5668,N_3149,N_3788);
and U5669 (N_5669,N_3247,N_3878);
nor U5670 (N_5670,N_3261,N_3364);
xnor U5671 (N_5671,N_3033,N_3009);
or U5672 (N_5672,N_3895,N_3673);
xor U5673 (N_5673,N_3408,N_3486);
xor U5674 (N_5674,N_3954,N_3979);
xnor U5675 (N_5675,N_4092,N_3280);
xor U5676 (N_5676,N_4413,N_3457);
and U5677 (N_5677,N_3347,N_3245);
and U5678 (N_5678,N_4038,N_3325);
nor U5679 (N_5679,N_4257,N_3077);
nor U5680 (N_5680,N_3920,N_3478);
nand U5681 (N_5681,N_4092,N_4000);
and U5682 (N_5682,N_3710,N_3514);
xor U5683 (N_5683,N_3422,N_3230);
xor U5684 (N_5684,N_4246,N_4144);
and U5685 (N_5685,N_3491,N_3044);
and U5686 (N_5686,N_3399,N_4369);
nor U5687 (N_5687,N_4371,N_3534);
nor U5688 (N_5688,N_3763,N_3344);
nor U5689 (N_5689,N_3640,N_3336);
xnor U5690 (N_5690,N_3983,N_4163);
and U5691 (N_5691,N_3128,N_3475);
or U5692 (N_5692,N_3496,N_3080);
nand U5693 (N_5693,N_3756,N_3662);
xnor U5694 (N_5694,N_3575,N_4487);
nor U5695 (N_5695,N_3143,N_4322);
nor U5696 (N_5696,N_4323,N_4267);
nor U5697 (N_5697,N_3250,N_4314);
xor U5698 (N_5698,N_3755,N_4363);
nand U5699 (N_5699,N_3601,N_3583);
xor U5700 (N_5700,N_3997,N_3829);
and U5701 (N_5701,N_4067,N_3931);
nor U5702 (N_5702,N_4380,N_3710);
nand U5703 (N_5703,N_3067,N_3150);
nand U5704 (N_5704,N_4029,N_3510);
and U5705 (N_5705,N_3781,N_3369);
xor U5706 (N_5706,N_3952,N_3054);
nand U5707 (N_5707,N_3014,N_3339);
nor U5708 (N_5708,N_3854,N_4382);
nand U5709 (N_5709,N_4028,N_4433);
or U5710 (N_5710,N_4152,N_3115);
xnor U5711 (N_5711,N_4127,N_3476);
and U5712 (N_5712,N_4497,N_3505);
or U5713 (N_5713,N_3974,N_3239);
nor U5714 (N_5714,N_3411,N_3246);
xnor U5715 (N_5715,N_4090,N_3040);
nor U5716 (N_5716,N_3264,N_4418);
or U5717 (N_5717,N_3830,N_3382);
or U5718 (N_5718,N_3678,N_3525);
nand U5719 (N_5719,N_4040,N_3964);
xnor U5720 (N_5720,N_3040,N_3301);
xnor U5721 (N_5721,N_4248,N_3656);
xor U5722 (N_5722,N_4403,N_3451);
xor U5723 (N_5723,N_3361,N_3550);
xor U5724 (N_5724,N_4301,N_3052);
and U5725 (N_5725,N_3583,N_3080);
or U5726 (N_5726,N_3201,N_3092);
and U5727 (N_5727,N_4244,N_3503);
nor U5728 (N_5728,N_4259,N_4114);
and U5729 (N_5729,N_4121,N_3552);
nor U5730 (N_5730,N_4097,N_4455);
nand U5731 (N_5731,N_3155,N_3388);
nand U5732 (N_5732,N_3566,N_3475);
xnor U5733 (N_5733,N_3560,N_3615);
nor U5734 (N_5734,N_4267,N_3516);
and U5735 (N_5735,N_3129,N_3175);
and U5736 (N_5736,N_3821,N_3042);
xor U5737 (N_5737,N_3884,N_4281);
nor U5738 (N_5738,N_4476,N_4186);
nor U5739 (N_5739,N_3479,N_3072);
nor U5740 (N_5740,N_3359,N_3155);
nand U5741 (N_5741,N_3284,N_3910);
or U5742 (N_5742,N_3593,N_3548);
nand U5743 (N_5743,N_3886,N_3792);
nand U5744 (N_5744,N_3113,N_4001);
nand U5745 (N_5745,N_4020,N_4459);
nand U5746 (N_5746,N_3143,N_4393);
nand U5747 (N_5747,N_4385,N_4380);
xor U5748 (N_5748,N_4149,N_3648);
nand U5749 (N_5749,N_4066,N_3829);
nand U5750 (N_5750,N_3177,N_3337);
nand U5751 (N_5751,N_4194,N_3500);
nor U5752 (N_5752,N_3822,N_3372);
xor U5753 (N_5753,N_3281,N_3826);
or U5754 (N_5754,N_3818,N_3403);
or U5755 (N_5755,N_3266,N_3642);
xnor U5756 (N_5756,N_4084,N_4389);
nand U5757 (N_5757,N_3340,N_4461);
xor U5758 (N_5758,N_3260,N_4179);
nor U5759 (N_5759,N_3797,N_4175);
nor U5760 (N_5760,N_4420,N_3514);
and U5761 (N_5761,N_3078,N_4231);
and U5762 (N_5762,N_4209,N_3893);
xnor U5763 (N_5763,N_3783,N_3229);
and U5764 (N_5764,N_3378,N_3697);
and U5765 (N_5765,N_4219,N_4430);
nand U5766 (N_5766,N_3420,N_3528);
xor U5767 (N_5767,N_3706,N_3318);
or U5768 (N_5768,N_3755,N_4211);
xor U5769 (N_5769,N_3576,N_4412);
xor U5770 (N_5770,N_3176,N_3913);
or U5771 (N_5771,N_3413,N_3397);
xor U5772 (N_5772,N_3237,N_3405);
and U5773 (N_5773,N_3184,N_4395);
and U5774 (N_5774,N_4315,N_3648);
nor U5775 (N_5775,N_3556,N_3281);
nor U5776 (N_5776,N_4048,N_3297);
nor U5777 (N_5777,N_3191,N_3282);
xor U5778 (N_5778,N_4001,N_3506);
nand U5779 (N_5779,N_3083,N_4428);
nand U5780 (N_5780,N_3653,N_4395);
and U5781 (N_5781,N_3559,N_3853);
xor U5782 (N_5782,N_3175,N_3891);
nor U5783 (N_5783,N_3638,N_3011);
or U5784 (N_5784,N_3573,N_3804);
nor U5785 (N_5785,N_4483,N_3241);
and U5786 (N_5786,N_4244,N_4335);
and U5787 (N_5787,N_4041,N_3644);
or U5788 (N_5788,N_4015,N_4207);
nor U5789 (N_5789,N_3472,N_3229);
nor U5790 (N_5790,N_3415,N_4426);
xnor U5791 (N_5791,N_3851,N_3020);
nor U5792 (N_5792,N_4128,N_3876);
nor U5793 (N_5793,N_4373,N_3958);
xnor U5794 (N_5794,N_4210,N_3437);
nand U5795 (N_5795,N_4181,N_4226);
and U5796 (N_5796,N_3703,N_3919);
nor U5797 (N_5797,N_3281,N_4165);
nand U5798 (N_5798,N_4395,N_3612);
nand U5799 (N_5799,N_4104,N_4148);
or U5800 (N_5800,N_3323,N_4294);
or U5801 (N_5801,N_3279,N_3798);
xnor U5802 (N_5802,N_3633,N_3054);
or U5803 (N_5803,N_3111,N_3208);
or U5804 (N_5804,N_4484,N_3201);
and U5805 (N_5805,N_3397,N_4307);
or U5806 (N_5806,N_3401,N_4145);
or U5807 (N_5807,N_4188,N_3819);
or U5808 (N_5808,N_4437,N_3131);
xor U5809 (N_5809,N_3540,N_3681);
xnor U5810 (N_5810,N_3922,N_4370);
xor U5811 (N_5811,N_4304,N_3545);
or U5812 (N_5812,N_4422,N_4386);
or U5813 (N_5813,N_3474,N_3648);
or U5814 (N_5814,N_3360,N_3985);
or U5815 (N_5815,N_3713,N_3573);
or U5816 (N_5816,N_3025,N_3109);
or U5817 (N_5817,N_3063,N_3594);
nand U5818 (N_5818,N_4384,N_3193);
or U5819 (N_5819,N_3124,N_4253);
and U5820 (N_5820,N_4452,N_3061);
or U5821 (N_5821,N_3360,N_3867);
nand U5822 (N_5822,N_3843,N_3014);
nor U5823 (N_5823,N_3312,N_3174);
nor U5824 (N_5824,N_3767,N_4400);
or U5825 (N_5825,N_3402,N_4062);
nor U5826 (N_5826,N_3139,N_3911);
nand U5827 (N_5827,N_3163,N_3501);
xnor U5828 (N_5828,N_3276,N_3851);
nand U5829 (N_5829,N_3032,N_3117);
nor U5830 (N_5830,N_3100,N_3583);
xor U5831 (N_5831,N_3297,N_3481);
and U5832 (N_5832,N_3734,N_3663);
and U5833 (N_5833,N_4389,N_4204);
nor U5834 (N_5834,N_3701,N_4340);
and U5835 (N_5835,N_3349,N_4318);
nor U5836 (N_5836,N_3547,N_3308);
nor U5837 (N_5837,N_3460,N_3662);
nand U5838 (N_5838,N_4394,N_3567);
and U5839 (N_5839,N_3902,N_3038);
or U5840 (N_5840,N_4110,N_4356);
nand U5841 (N_5841,N_4168,N_3396);
nor U5842 (N_5842,N_4465,N_4305);
and U5843 (N_5843,N_3507,N_4158);
nor U5844 (N_5844,N_3235,N_3556);
nand U5845 (N_5845,N_3823,N_3396);
or U5846 (N_5846,N_3842,N_4442);
and U5847 (N_5847,N_4025,N_3983);
nand U5848 (N_5848,N_3084,N_3818);
or U5849 (N_5849,N_3202,N_3037);
xor U5850 (N_5850,N_3482,N_3159);
and U5851 (N_5851,N_3576,N_4172);
or U5852 (N_5852,N_3725,N_3132);
nor U5853 (N_5853,N_4346,N_4483);
nand U5854 (N_5854,N_3161,N_3228);
nor U5855 (N_5855,N_3662,N_4383);
xnor U5856 (N_5856,N_3557,N_4217);
nor U5857 (N_5857,N_3766,N_3995);
and U5858 (N_5858,N_3440,N_4260);
nor U5859 (N_5859,N_3262,N_3124);
xnor U5860 (N_5860,N_3447,N_3385);
xor U5861 (N_5861,N_4075,N_3164);
or U5862 (N_5862,N_3328,N_3028);
nor U5863 (N_5863,N_4146,N_3534);
nand U5864 (N_5864,N_4327,N_3419);
or U5865 (N_5865,N_4373,N_3892);
nor U5866 (N_5866,N_3745,N_3656);
or U5867 (N_5867,N_3690,N_4255);
or U5868 (N_5868,N_3847,N_3600);
or U5869 (N_5869,N_3962,N_3300);
nor U5870 (N_5870,N_4175,N_3661);
nor U5871 (N_5871,N_4366,N_4275);
nand U5872 (N_5872,N_3160,N_3120);
and U5873 (N_5873,N_3917,N_3936);
or U5874 (N_5874,N_4252,N_3453);
and U5875 (N_5875,N_3655,N_3090);
nor U5876 (N_5876,N_4144,N_3988);
nand U5877 (N_5877,N_4418,N_4042);
or U5878 (N_5878,N_3263,N_3767);
or U5879 (N_5879,N_3535,N_4119);
or U5880 (N_5880,N_3786,N_4463);
and U5881 (N_5881,N_3020,N_3948);
xor U5882 (N_5882,N_4091,N_3652);
and U5883 (N_5883,N_3364,N_3176);
or U5884 (N_5884,N_4454,N_4285);
nand U5885 (N_5885,N_3611,N_3704);
or U5886 (N_5886,N_4142,N_4295);
nor U5887 (N_5887,N_4282,N_3670);
nand U5888 (N_5888,N_3296,N_3198);
xor U5889 (N_5889,N_3248,N_3140);
and U5890 (N_5890,N_3371,N_3722);
nor U5891 (N_5891,N_4456,N_3124);
xnor U5892 (N_5892,N_3535,N_3001);
nand U5893 (N_5893,N_3562,N_3541);
nand U5894 (N_5894,N_3234,N_4391);
nor U5895 (N_5895,N_3735,N_4471);
and U5896 (N_5896,N_3529,N_3897);
nor U5897 (N_5897,N_3197,N_3139);
or U5898 (N_5898,N_4128,N_3984);
or U5899 (N_5899,N_3265,N_3377);
xor U5900 (N_5900,N_3643,N_4421);
nand U5901 (N_5901,N_3590,N_3439);
nor U5902 (N_5902,N_3634,N_3185);
xor U5903 (N_5903,N_4262,N_3791);
xor U5904 (N_5904,N_3861,N_3080);
nor U5905 (N_5905,N_4440,N_3592);
nor U5906 (N_5906,N_4075,N_3452);
xor U5907 (N_5907,N_3011,N_4298);
nand U5908 (N_5908,N_4498,N_3639);
nand U5909 (N_5909,N_3910,N_4091);
and U5910 (N_5910,N_4392,N_4277);
nand U5911 (N_5911,N_3209,N_3072);
or U5912 (N_5912,N_4425,N_3912);
and U5913 (N_5913,N_4067,N_3816);
xnor U5914 (N_5914,N_3483,N_3494);
nor U5915 (N_5915,N_3842,N_4332);
or U5916 (N_5916,N_4131,N_3293);
nand U5917 (N_5917,N_3495,N_4098);
or U5918 (N_5918,N_4156,N_3867);
nor U5919 (N_5919,N_3591,N_4355);
and U5920 (N_5920,N_3798,N_4076);
nor U5921 (N_5921,N_3907,N_3812);
nor U5922 (N_5922,N_3020,N_3612);
and U5923 (N_5923,N_4079,N_4403);
and U5924 (N_5924,N_4490,N_4088);
or U5925 (N_5925,N_3631,N_4014);
xor U5926 (N_5926,N_4399,N_4070);
nor U5927 (N_5927,N_3375,N_4074);
nand U5928 (N_5928,N_3730,N_3572);
or U5929 (N_5929,N_3893,N_3938);
and U5930 (N_5930,N_3147,N_3138);
or U5931 (N_5931,N_4496,N_3535);
nor U5932 (N_5932,N_4367,N_4366);
xnor U5933 (N_5933,N_4341,N_3207);
nand U5934 (N_5934,N_4001,N_4077);
nand U5935 (N_5935,N_3280,N_3106);
xor U5936 (N_5936,N_3915,N_3464);
xor U5937 (N_5937,N_4263,N_4385);
nor U5938 (N_5938,N_3951,N_3182);
and U5939 (N_5939,N_3841,N_3228);
nor U5940 (N_5940,N_4024,N_4449);
xor U5941 (N_5941,N_3702,N_3867);
nand U5942 (N_5942,N_3047,N_4219);
and U5943 (N_5943,N_3583,N_4050);
xor U5944 (N_5944,N_4157,N_4427);
and U5945 (N_5945,N_4433,N_3972);
xor U5946 (N_5946,N_3625,N_4016);
or U5947 (N_5947,N_3310,N_4465);
nor U5948 (N_5948,N_3249,N_3764);
nand U5949 (N_5949,N_3719,N_3586);
nor U5950 (N_5950,N_3664,N_3431);
xnor U5951 (N_5951,N_3205,N_3902);
and U5952 (N_5952,N_3038,N_3169);
or U5953 (N_5953,N_3039,N_3295);
or U5954 (N_5954,N_3181,N_3748);
or U5955 (N_5955,N_3574,N_4262);
nor U5956 (N_5956,N_4081,N_3641);
or U5957 (N_5957,N_3624,N_3855);
xnor U5958 (N_5958,N_4377,N_3176);
xnor U5959 (N_5959,N_4195,N_3598);
nand U5960 (N_5960,N_3418,N_3109);
or U5961 (N_5961,N_4096,N_3160);
or U5962 (N_5962,N_3516,N_4174);
xnor U5963 (N_5963,N_3248,N_3699);
or U5964 (N_5964,N_4013,N_4490);
or U5965 (N_5965,N_4090,N_3143);
nand U5966 (N_5966,N_4041,N_3166);
and U5967 (N_5967,N_3754,N_3786);
nand U5968 (N_5968,N_3683,N_3738);
nand U5969 (N_5969,N_4224,N_3470);
nor U5970 (N_5970,N_3235,N_4132);
xor U5971 (N_5971,N_3995,N_3203);
or U5972 (N_5972,N_3735,N_3809);
or U5973 (N_5973,N_3402,N_3300);
and U5974 (N_5974,N_4217,N_3153);
xor U5975 (N_5975,N_3959,N_3531);
nand U5976 (N_5976,N_4127,N_3991);
or U5977 (N_5977,N_3075,N_3235);
and U5978 (N_5978,N_4428,N_3329);
nand U5979 (N_5979,N_3226,N_4308);
nand U5980 (N_5980,N_3024,N_3056);
xnor U5981 (N_5981,N_3092,N_3125);
nor U5982 (N_5982,N_3128,N_4395);
and U5983 (N_5983,N_3315,N_3564);
nor U5984 (N_5984,N_4222,N_3052);
or U5985 (N_5985,N_3861,N_4239);
nand U5986 (N_5986,N_3727,N_3040);
nor U5987 (N_5987,N_3999,N_3238);
xor U5988 (N_5988,N_4441,N_3902);
nor U5989 (N_5989,N_4286,N_4098);
or U5990 (N_5990,N_3412,N_4075);
nand U5991 (N_5991,N_4011,N_3580);
nand U5992 (N_5992,N_3063,N_3700);
or U5993 (N_5993,N_3878,N_4489);
and U5994 (N_5994,N_3780,N_3794);
and U5995 (N_5995,N_4115,N_3502);
and U5996 (N_5996,N_4019,N_3492);
nand U5997 (N_5997,N_3703,N_3299);
xor U5998 (N_5998,N_4172,N_3090);
nor U5999 (N_5999,N_4399,N_3226);
or U6000 (N_6000,N_5742,N_5264);
nand U6001 (N_6001,N_4690,N_4938);
and U6002 (N_6002,N_4726,N_5666);
nor U6003 (N_6003,N_5593,N_5265);
xor U6004 (N_6004,N_4941,N_4633);
and U6005 (N_6005,N_5288,N_5020);
nor U6006 (N_6006,N_4922,N_4934);
or U6007 (N_6007,N_5116,N_5966);
and U6008 (N_6008,N_4824,N_4780);
xor U6009 (N_6009,N_4801,N_4515);
nand U6010 (N_6010,N_4527,N_4597);
xor U6011 (N_6011,N_4870,N_5410);
xnor U6012 (N_6012,N_5325,N_5186);
nand U6013 (N_6013,N_5753,N_4644);
nand U6014 (N_6014,N_4742,N_4585);
nand U6015 (N_6015,N_4807,N_5363);
nand U6016 (N_6016,N_4538,N_5228);
or U6017 (N_6017,N_5313,N_5604);
nand U6018 (N_6018,N_5338,N_4857);
nor U6019 (N_6019,N_4884,N_5714);
and U6020 (N_6020,N_4674,N_5339);
xor U6021 (N_6021,N_5175,N_5520);
and U6022 (N_6022,N_4565,N_5305);
xor U6023 (N_6023,N_5403,N_5673);
xor U6024 (N_6024,N_4624,N_5408);
or U6025 (N_6025,N_4841,N_5668);
and U6026 (N_6026,N_4809,N_5098);
nor U6027 (N_6027,N_5999,N_4984);
nor U6028 (N_6028,N_5617,N_4792);
nor U6029 (N_6029,N_5277,N_5922);
nor U6030 (N_6030,N_5804,N_5029);
or U6031 (N_6031,N_5995,N_5214);
or U6032 (N_6032,N_5597,N_4756);
or U6033 (N_6033,N_5528,N_4897);
or U6034 (N_6034,N_5192,N_4730);
and U6035 (N_6035,N_5287,N_4510);
and U6036 (N_6036,N_5961,N_5374);
nand U6037 (N_6037,N_5881,N_4603);
and U6038 (N_6038,N_5609,N_4818);
nor U6039 (N_6039,N_5188,N_5126);
xnor U6040 (N_6040,N_5758,N_4960);
or U6041 (N_6041,N_5064,N_5868);
nor U6042 (N_6042,N_4649,N_5909);
nor U6043 (N_6043,N_4814,N_5774);
nand U6044 (N_6044,N_5902,N_5349);
nor U6045 (N_6045,N_4923,N_5889);
or U6046 (N_6046,N_5854,N_4576);
and U6047 (N_6047,N_5275,N_4868);
xor U6048 (N_6048,N_4976,N_4678);
nand U6049 (N_6049,N_5406,N_4663);
nand U6050 (N_6050,N_5424,N_5776);
nor U6051 (N_6051,N_4518,N_4547);
xor U6052 (N_6052,N_5343,N_5642);
or U6053 (N_6053,N_4973,N_5689);
xor U6054 (N_6054,N_5795,N_5835);
and U6055 (N_6055,N_5205,N_5130);
or U6056 (N_6056,N_5501,N_5887);
and U6057 (N_6057,N_5483,N_5649);
and U6058 (N_6058,N_5249,N_5346);
nand U6059 (N_6059,N_5439,N_5687);
and U6060 (N_6060,N_5762,N_4542);
or U6061 (N_6061,N_5310,N_4912);
nand U6062 (N_6062,N_4561,N_4871);
or U6063 (N_6063,N_5226,N_4901);
nor U6064 (N_6064,N_4760,N_4571);
or U6065 (N_6065,N_5820,N_4860);
and U6066 (N_6066,N_5905,N_5947);
nor U6067 (N_6067,N_5998,N_4735);
nand U6068 (N_6068,N_4757,N_5910);
and U6069 (N_6069,N_5037,N_5197);
and U6070 (N_6070,N_5153,N_5371);
nand U6071 (N_6071,N_4718,N_5353);
xor U6072 (N_6072,N_5559,N_5691);
xnor U6073 (N_6073,N_4847,N_5605);
nand U6074 (N_6074,N_4519,N_5454);
and U6075 (N_6075,N_4556,N_4570);
or U6076 (N_6076,N_5841,N_5282);
nand U6077 (N_6077,N_4671,N_4640);
and U6078 (N_6078,N_5300,N_5522);
or U6079 (N_6079,N_4721,N_5392);
nor U6080 (N_6080,N_5464,N_5179);
and U6081 (N_6081,N_5651,N_5055);
nand U6082 (N_6082,N_5561,N_5571);
or U6083 (N_6083,N_5328,N_4902);
or U6084 (N_6084,N_5811,N_4883);
xnor U6085 (N_6085,N_5019,N_5199);
and U6086 (N_6086,N_5211,N_4957);
xor U6087 (N_6087,N_5007,N_4985);
and U6088 (N_6088,N_4577,N_4851);
xor U6089 (N_6089,N_5203,N_5843);
or U6090 (N_6090,N_5735,N_5636);
xnor U6091 (N_6091,N_4692,N_4647);
xnor U6092 (N_6092,N_5252,N_5366);
nand U6093 (N_6093,N_5110,N_5629);
nor U6094 (N_6094,N_5195,N_5499);
nor U6095 (N_6095,N_5690,N_4689);
nand U6096 (N_6096,N_4521,N_4684);
and U6097 (N_6097,N_4914,N_5646);
and U6098 (N_6098,N_5564,N_4716);
or U6099 (N_6099,N_4959,N_5163);
and U6100 (N_6100,N_4790,N_4535);
xnor U6101 (N_6101,N_5993,N_5221);
nor U6102 (N_6102,N_4793,N_4995);
and U6103 (N_6103,N_5572,N_5549);
or U6104 (N_6104,N_5793,N_4778);
xor U6105 (N_6105,N_4614,N_5682);
nor U6106 (N_6106,N_5284,N_5553);
xnor U6107 (N_6107,N_5659,N_4893);
nor U6108 (N_6108,N_5273,N_5853);
and U6109 (N_6109,N_5624,N_4746);
and U6110 (N_6110,N_4864,N_5375);
and U6111 (N_6111,N_4832,N_5503);
nor U6112 (N_6112,N_5040,N_5469);
xor U6113 (N_6113,N_5451,N_5121);
nor U6114 (N_6114,N_5208,N_5162);
nor U6115 (N_6115,N_5294,N_5931);
xnor U6116 (N_6116,N_4567,N_5434);
nor U6117 (N_6117,N_5065,N_4651);
and U6118 (N_6118,N_5489,N_5465);
nor U6119 (N_6119,N_5317,N_4728);
nand U6120 (N_6120,N_5089,N_5828);
nor U6121 (N_6121,N_4619,N_5005);
nand U6122 (N_6122,N_5837,N_4963);
and U6123 (N_6123,N_4749,N_5314);
nand U6124 (N_6124,N_5747,N_5700);
nand U6125 (N_6125,N_5103,N_5036);
xor U6126 (N_6126,N_5140,N_5053);
and U6127 (N_6127,N_4930,N_5632);
and U6128 (N_6128,N_4795,N_4589);
xor U6129 (N_6129,N_4891,N_5698);
nand U6130 (N_6130,N_5918,N_4745);
and U6131 (N_6131,N_5268,N_5271);
or U6132 (N_6132,N_5033,N_5519);
or U6133 (N_6133,N_4681,N_5704);
nor U6134 (N_6134,N_4656,N_4732);
and U6135 (N_6135,N_5847,N_4849);
xnor U6136 (N_6136,N_5969,N_4541);
and U6137 (N_6137,N_5105,N_4978);
nand U6138 (N_6138,N_5091,N_5468);
nor U6139 (N_6139,N_5009,N_5183);
nor U6140 (N_6140,N_5874,N_5272);
nand U6141 (N_6141,N_4609,N_4815);
and U6142 (N_6142,N_5708,N_4805);
nand U6143 (N_6143,N_5006,N_4942);
and U6144 (N_6144,N_4968,N_5705);
and U6145 (N_6145,N_5903,N_5702);
or U6146 (N_6146,N_5027,N_4852);
nor U6147 (N_6147,N_4675,N_5832);
and U6148 (N_6148,N_5965,N_4629);
nand U6149 (N_6149,N_5808,N_4618);
or U6150 (N_6150,N_4856,N_5372);
nor U6151 (N_6151,N_5769,N_5177);
nand U6152 (N_6152,N_5633,N_5144);
or U6153 (N_6153,N_4774,N_4982);
or U6154 (N_6154,N_5679,N_5773);
nand U6155 (N_6155,N_5224,N_5759);
nor U6156 (N_6156,N_5670,N_4927);
nand U6157 (N_6157,N_5667,N_5125);
and U6158 (N_6158,N_5621,N_4586);
nand U6159 (N_6159,N_5547,N_5821);
nor U6160 (N_6160,N_4701,N_5112);
nor U6161 (N_6161,N_5723,N_5957);
and U6162 (N_6162,N_5160,N_5663);
nand U6163 (N_6163,N_5446,N_5058);
and U6164 (N_6164,N_4668,N_4940);
or U6165 (N_6165,N_4806,N_5671);
xnor U6166 (N_6166,N_4572,N_4558);
nor U6167 (N_6167,N_5817,N_5538);
or U6168 (N_6168,N_5291,N_4557);
or U6169 (N_6169,N_5100,N_4817);
nand U6170 (N_6170,N_4606,N_5435);
or U6171 (N_6171,N_5971,N_4705);
nor U6172 (N_6172,N_4588,N_4693);
nand U6173 (N_6173,N_4773,N_4990);
or U6174 (N_6174,N_5959,N_4986);
or U6175 (N_6175,N_5142,N_5643);
nor U6176 (N_6176,N_4816,N_5013);
nand U6177 (N_6177,N_5516,N_5767);
xnor U6178 (N_6178,N_5086,N_5492);
or U6179 (N_6179,N_5378,N_5757);
or U6180 (N_6180,N_4869,N_5182);
nor U6181 (N_6181,N_4833,N_5337);
and U6182 (N_6182,N_5864,N_4747);
or U6183 (N_6183,N_4639,N_5048);
nand U6184 (N_6184,N_5088,N_5109);
and U6185 (N_6185,N_5598,N_5133);
xor U6186 (N_6186,N_5258,N_4720);
or U6187 (N_6187,N_5067,N_5479);
nand U6188 (N_6188,N_5173,N_5738);
and U6189 (N_6189,N_4744,N_5049);
nor U6190 (N_6190,N_4977,N_5685);
nor U6191 (N_6191,N_4766,N_5072);
xor U6192 (N_6192,N_5229,N_4786);
nor U6193 (N_6193,N_5672,N_4611);
xor U6194 (N_6194,N_4632,N_5139);
nand U6195 (N_6195,N_4553,N_5824);
or U6196 (N_6196,N_4579,N_4712);
and U6197 (N_6197,N_5455,N_5176);
nand U6198 (N_6198,N_4789,N_4791);
nor U6199 (N_6199,N_4759,N_5584);
nand U6200 (N_6200,N_4706,N_4582);
or U6201 (N_6201,N_5567,N_4802);
nor U6202 (N_6202,N_5569,N_5216);
and U6203 (N_6203,N_5341,N_5085);
and U6204 (N_6204,N_4564,N_5780);
xnor U6205 (N_6205,N_5172,N_5122);
nand U6206 (N_6206,N_4843,N_4872);
nand U6207 (N_6207,N_5200,N_4788);
and U6208 (N_6208,N_4770,N_5857);
nor U6209 (N_6209,N_5322,N_5878);
and U6210 (N_6210,N_5482,N_4933);
and U6211 (N_6211,N_5791,N_5045);
xor U6212 (N_6212,N_4638,N_4544);
or U6213 (N_6213,N_4981,N_5478);
and U6214 (N_6214,N_5278,N_4988);
and U6215 (N_6215,N_5324,N_5494);
nor U6216 (N_6216,N_5900,N_5094);
xnor U6217 (N_6217,N_4550,N_4915);
xnor U6218 (N_6218,N_4520,N_5801);
or U6219 (N_6219,N_4636,N_5321);
nor U6220 (N_6220,N_5781,N_5137);
xor U6221 (N_6221,N_5075,N_5246);
nor U6222 (N_6222,N_5442,N_5364);
or U6223 (N_6223,N_5512,N_5823);
or U6224 (N_6224,N_5379,N_5891);
and U6225 (N_6225,N_5031,N_5296);
or U6226 (N_6226,N_5161,N_4993);
xor U6227 (N_6227,N_4669,N_5761);
nand U6228 (N_6228,N_5010,N_4787);
xnor U6229 (N_6229,N_4551,N_4729);
nor U6230 (N_6230,N_5996,N_5401);
and U6231 (N_6231,N_5985,N_5003);
xor U6232 (N_6232,N_5323,N_5008);
xnor U6233 (N_6233,N_5949,N_4574);
xor U6234 (N_6234,N_5754,N_5202);
nand U6235 (N_6235,N_5069,N_5194);
and U6236 (N_6236,N_4667,N_5231);
nor U6237 (N_6237,N_5393,N_5276);
or U6238 (N_6238,N_5653,N_5858);
nand U6239 (N_6239,N_4748,N_4830);
and U6240 (N_6240,N_5867,N_5307);
xnor U6241 (N_6241,N_5894,N_5748);
xnor U6242 (N_6242,N_5132,N_5756);
xor U6243 (N_6243,N_5213,N_5805);
nand U6244 (N_6244,N_5701,N_5413);
or U6245 (N_6245,N_5852,N_5688);
nand U6246 (N_6246,N_5627,N_4896);
xnor U6247 (N_6247,N_4661,N_5635);
xor U6248 (N_6248,N_4970,N_5071);
nand U6249 (N_6249,N_5873,N_5728);
xnor U6250 (N_6250,N_5694,N_5234);
nor U6251 (N_6251,N_5607,N_4925);
xor U6252 (N_6252,N_5380,N_5458);
or U6253 (N_6253,N_4500,N_5580);
nor U6254 (N_6254,N_5542,N_5518);
nand U6255 (N_6255,N_5746,N_4874);
nor U6256 (N_6256,N_4698,N_5897);
nor U6257 (N_6257,N_5052,N_5354);
or U6258 (N_6258,N_5243,N_5638);
nor U6259 (N_6259,N_5908,N_5493);
xor U6260 (N_6260,N_5525,N_4821);
nand U6261 (N_6261,N_5012,N_5331);
nand U6262 (N_6262,N_4514,N_5625);
or U6263 (N_6263,N_5713,N_5751);
nor U6264 (N_6264,N_5418,N_4894);
xnor U6265 (N_6265,N_5676,N_4762);
and U6266 (N_6266,N_5509,N_5540);
or U6267 (N_6267,N_5259,N_5391);
nand U6268 (N_6268,N_5718,N_5802);
or U6269 (N_6269,N_5425,N_5546);
and U6270 (N_6270,N_5241,N_5741);
xnor U6271 (N_6271,N_5506,N_5332);
or U6272 (N_6272,N_5788,N_5253);
and U6273 (N_6273,N_5395,N_4763);
nand U6274 (N_6274,N_4682,N_5591);
nand U6275 (N_6275,N_4559,N_4767);
nor U6276 (N_6276,N_4555,N_5920);
or U6277 (N_6277,N_4622,N_4879);
xor U6278 (N_6278,N_4511,N_5420);
or U6279 (N_6279,N_4642,N_4599);
or U6280 (N_6280,N_5450,N_5785);
and U6281 (N_6281,N_5002,N_4584);
or U6282 (N_6282,N_5766,N_4837);
nor U6283 (N_6283,N_5021,N_5017);
nor U6284 (N_6284,N_4994,N_5543);
nand U6285 (N_6285,N_4890,N_5462);
nand U6286 (N_6286,N_4810,N_4560);
xnor U6287 (N_6287,N_5586,N_5937);
or U6288 (N_6288,N_4964,N_5536);
or U6289 (N_6289,N_5427,N_5831);
or U6290 (N_6290,N_5926,N_5001);
nor U6291 (N_6291,N_5432,N_4835);
or U6292 (N_6292,N_4563,N_5882);
or U6293 (N_6293,N_4797,N_5476);
and U6294 (N_6294,N_4575,N_5818);
nor U6295 (N_6295,N_5846,N_5764);
xnor U6296 (N_6296,N_5712,N_5157);
xnor U6297 (N_6297,N_5026,N_4710);
nand U6298 (N_6298,N_5452,N_4549);
xor U6299 (N_6299,N_5641,N_5024);
and U6300 (N_6300,N_5825,N_5032);
nand U6301 (N_6301,N_5496,N_5815);
nand U6302 (N_6302,N_4862,N_4507);
xnor U6303 (N_6303,N_5146,N_5888);
and U6304 (N_6304,N_4943,N_4892);
or U6305 (N_6305,N_5628,N_5612);
xor U6306 (N_6306,N_4751,N_4725);
xnor U6307 (N_6307,N_5799,N_5219);
nand U6308 (N_6308,N_5958,N_5885);
nor U6309 (N_6309,N_5581,N_5204);
and U6310 (N_6310,N_5935,N_4936);
xnor U6311 (N_6311,N_4867,N_5806);
or U6312 (N_6312,N_5719,N_5365);
nor U6313 (N_6313,N_4662,N_4715);
nor U6314 (N_6314,N_5979,N_5113);
and U6315 (N_6315,N_4947,N_5099);
nand U6316 (N_6316,N_5989,N_5675);
xor U6317 (N_6317,N_4665,N_5883);
or U6318 (N_6318,N_5899,N_5967);
and U6319 (N_6319,N_5412,N_5886);
and U6320 (N_6320,N_5927,N_4889);
xnor U6321 (N_6321,N_5051,N_4630);
and U6322 (N_6322,N_5212,N_5230);
nand U6323 (N_6323,N_5645,N_4637);
nand U6324 (N_6324,N_5150,N_5149);
or U6325 (N_6325,N_5267,N_5844);
nor U6326 (N_6326,N_4741,N_5775);
or U6327 (N_6327,N_5119,N_5596);
nand U6328 (N_6328,N_5428,N_4608);
xnor U6329 (N_6329,N_5725,N_5644);
nand U6330 (N_6330,N_5640,N_5491);
or U6331 (N_6331,N_5752,N_4880);
and U6332 (N_6332,N_5715,N_5803);
nor U6333 (N_6333,N_4903,N_4910);
nor U6334 (N_6334,N_5351,N_4615);
nor U6335 (N_6335,N_4811,N_5210);
or U6336 (N_6336,N_5326,N_4881);
nand U6337 (N_6337,N_4823,N_5247);
nor U6338 (N_6338,N_4502,N_4583);
nand U6339 (N_6339,N_5181,N_5921);
nor U6340 (N_6340,N_5035,N_5991);
nand U6341 (N_6341,N_4731,N_5184);
or U6342 (N_6342,N_5656,N_4854);
nor U6343 (N_6343,N_5073,N_5426);
or U6344 (N_6344,N_5928,N_5655);
or U6345 (N_6345,N_5107,N_5980);
and U6346 (N_6346,N_4772,N_5532);
nand U6347 (N_6347,N_5892,N_5480);
xnor U6348 (N_6348,N_5855,N_4612);
nor U6349 (N_6349,N_5830,N_5616);
xor U6350 (N_6350,N_5523,N_4702);
or U6351 (N_6351,N_4782,N_4617);
nor U6352 (N_6352,N_5749,N_5608);
or U6353 (N_6353,N_5779,N_5913);
and U6354 (N_6354,N_4952,N_4524);
nor U6355 (N_6355,N_5384,N_4946);
xor U6356 (N_6356,N_5106,N_4685);
nand U6357 (N_6357,N_5526,N_5279);
nand U6358 (N_6358,N_5916,N_5626);
nand U6359 (N_6359,N_5357,N_5527);
nand U6360 (N_6360,N_5274,N_5743);
nand U6361 (N_6361,N_5495,N_5860);
nor U6362 (N_6362,N_5070,N_5535);
or U6363 (N_6363,N_4740,N_5023);
nor U6364 (N_6364,N_5034,N_5983);
xor U6365 (N_6365,N_5865,N_4935);
xor U6366 (N_6366,N_5447,N_5739);
xnor U6367 (N_6367,N_4825,N_5056);
xor U6368 (N_6368,N_5129,N_4804);
nor U6369 (N_6369,N_5409,N_5810);
and U6370 (N_6370,N_5703,N_5960);
nand U6371 (N_6371,N_4566,N_4955);
and U6372 (N_6372,N_4523,N_4727);
nor U6373 (N_6373,N_4737,N_5763);
or U6374 (N_6374,N_4664,N_5370);
and U6375 (N_6375,N_5330,N_5724);
and U6376 (N_6376,N_5449,N_5474);
xor U6377 (N_6377,N_5000,N_4808);
or U6378 (N_6378,N_5514,N_5770);
or U6379 (N_6379,N_5568,N_5639);
and U6380 (N_6380,N_4826,N_5956);
nor U6381 (N_6381,N_5551,N_5530);
and U6382 (N_6382,N_5383,N_5602);
or U6383 (N_6383,N_5360,N_5537);
and U6384 (N_6384,N_4820,N_5730);
or U6385 (N_6385,N_4828,N_5430);
and U6386 (N_6386,N_5083,N_5263);
xnor U6387 (N_6387,N_5115,N_5794);
or U6388 (N_6388,N_5912,N_5934);
nor U6389 (N_6389,N_5727,N_5101);
xor U6390 (N_6390,N_5588,N_4761);
nand U6391 (N_6391,N_5662,N_5601);
nand U6392 (N_6392,N_5373,N_4919);
xor U6393 (N_6393,N_4913,N_5510);
xor U6394 (N_6394,N_5312,N_5074);
or U6395 (N_6395,N_5185,N_5421);
nand U6396 (N_6396,N_5180,N_5444);
nor U6397 (N_6397,N_4967,N_5554);
or U6398 (N_6398,N_5654,N_5152);
or U6399 (N_6399,N_4827,N_5368);
nand U6400 (N_6400,N_4646,N_5585);
and U6401 (N_6401,N_4845,N_5982);
and U6402 (N_6402,N_4704,N_5318);
nor U6403 (N_6403,N_4873,N_4887);
and U6404 (N_6404,N_4516,N_5981);
or U6405 (N_6405,N_5481,N_4736);
nor U6406 (N_6406,N_5147,N_5484);
xor U6407 (N_6407,N_4552,N_5740);
and U6408 (N_6408,N_4711,N_5706);
nand U6409 (N_6409,N_5848,N_4595);
xor U6410 (N_6410,N_5223,N_4709);
nor U6411 (N_6411,N_4593,N_4522);
nor U6412 (N_6412,N_4954,N_5573);
nor U6413 (N_6413,N_5834,N_5164);
nor U6414 (N_6414,N_5080,N_5623);
and U6415 (N_6415,N_5377,N_5772);
and U6416 (N_6416,N_4819,N_4951);
xnor U6417 (N_6417,N_5039,N_4691);
or U6418 (N_6418,N_5155,N_4545);
and U6419 (N_6419,N_5390,N_4983);
or U6420 (N_6420,N_4532,N_5570);
nand U6421 (N_6421,N_5695,N_5787);
nand U6422 (N_6422,N_4813,N_4598);
xnor U6423 (N_6423,N_5813,N_4907);
nand U6424 (N_6424,N_5513,N_4839);
and U6425 (N_6425,N_5871,N_5678);
and U6426 (N_6426,N_5603,N_4965);
nand U6427 (N_6427,N_5304,N_5850);
or U6428 (N_6428,N_5196,N_5171);
nor U6429 (N_6429,N_5765,N_4653);
nor U6430 (N_6430,N_5260,N_4796);
nand U6431 (N_6431,N_5063,N_5558);
or U6432 (N_6432,N_5316,N_5295);
nor U6433 (N_6433,N_5952,N_5541);
nor U6434 (N_6434,N_5340,N_5220);
or U6435 (N_6435,N_5755,N_4974);
nand U6436 (N_6436,N_5309,N_5385);
xor U6437 (N_6437,N_4949,N_5433);
nand U6438 (N_6438,N_4660,N_5209);
nand U6439 (N_6439,N_4987,N_5077);
nand U6440 (N_6440,N_5497,N_4866);
and U6441 (N_6441,N_5710,N_5143);
nand U6442 (N_6442,N_5664,N_5261);
or U6443 (N_6443,N_5986,N_4714);
nor U6444 (N_6444,N_5092,N_4580);
or U6445 (N_6445,N_5108,N_5303);
and U6446 (N_6446,N_5436,N_5404);
or U6447 (N_6447,N_4505,N_5575);
or U6448 (N_6448,N_5845,N_5043);
xnor U6449 (N_6449,N_5851,N_5976);
and U6450 (N_6450,N_4855,N_5582);
and U6451 (N_6451,N_4743,N_5872);
nand U6452 (N_6452,N_5674,N_4650);
nand U6453 (N_6453,N_5217,N_4680);
nor U6454 (N_6454,N_5552,N_4548);
or U6455 (N_6455,N_5583,N_4758);
and U6456 (N_6456,N_5207,N_5944);
xnor U6457 (N_6457,N_5657,N_5789);
nand U6458 (N_6458,N_5565,N_4812);
nor U6459 (N_6459,N_4533,N_4686);
nand U6460 (N_6460,N_4623,N_4917);
and U6461 (N_6461,N_4707,N_5443);
nand U6462 (N_6462,N_5342,N_5592);
xnor U6463 (N_6463,N_5004,N_5517);
and U6464 (N_6464,N_5948,N_5336);
and U6465 (N_6465,N_5359,N_5915);
or U6466 (N_6466,N_4526,N_4937);
xor U6467 (N_6467,N_5256,N_5987);
nor U6468 (N_6468,N_5729,N_5890);
or U6469 (N_6469,N_5576,N_4604);
nand U6470 (N_6470,N_5472,N_5151);
and U6471 (N_6471,N_4590,N_5637);
xor U6472 (N_6472,N_5471,N_4752);
or U6473 (N_6473,N_5929,N_5170);
nor U6474 (N_6474,N_5327,N_4768);
xnor U6475 (N_6475,N_4676,N_4996);
nor U6476 (N_6476,N_5270,N_5650);
nor U6477 (N_6477,N_4591,N_5721);
nand U6478 (N_6478,N_5215,N_5079);
xor U6479 (N_6479,N_5333,N_5355);
nor U6480 (N_6480,N_4708,N_4562);
and U6481 (N_6481,N_5145,N_5445);
xnor U6482 (N_6482,N_4657,N_5159);
or U6483 (N_6483,N_5838,N_5135);
or U6484 (N_6484,N_5997,N_4546);
and U6485 (N_6485,N_5533,N_5136);
nand U6486 (N_6486,N_5235,N_5329);
and U6487 (N_6487,N_4648,N_5942);
nand U6488 (N_6488,N_4822,N_5093);
xnor U6489 (N_6489,N_5350,N_5233);
or U6490 (N_6490,N_5932,N_4683);
or U6491 (N_6491,N_4895,N_4635);
nand U6492 (N_6492,N_4695,N_4908);
or U6493 (N_6493,N_5500,N_5293);
or U6494 (N_6494,N_5907,N_4602);
and U6495 (N_6495,N_4528,N_4569);
and U6496 (N_6496,N_5477,N_4956);
and U6497 (N_6497,N_5941,N_5790);
or U6498 (N_6498,N_5977,N_5298);
and U6499 (N_6499,N_5485,N_5505);
and U6500 (N_6500,N_5407,N_5311);
xor U6501 (N_6501,N_4659,N_5118);
nand U6502 (N_6502,N_4932,N_4679);
nor U6503 (N_6503,N_5615,N_4775);
nor U6504 (N_6504,N_4537,N_5863);
or U6505 (N_6505,N_5978,N_5166);
or U6506 (N_6506,N_5306,N_5560);
or U6507 (N_6507,N_4800,N_5038);
xnor U6508 (N_6508,N_5722,N_4739);
nand U6509 (N_6509,N_4885,N_4850);
nand U6510 (N_6510,N_4733,N_5399);
nand U6511 (N_6511,N_5473,N_5244);
nand U6512 (N_6512,N_5281,N_4631);
nor U6513 (N_6513,N_5974,N_5193);
nand U6514 (N_6514,N_4950,N_5201);
nor U6515 (N_6515,N_5387,N_5661);
xnor U6516 (N_6516,N_5382,N_5778);
or U6517 (N_6517,N_5699,N_4876);
or U6518 (N_6518,N_4628,N_5386);
xnor U6519 (N_6519,N_4840,N_5933);
or U6520 (N_6520,N_4607,N_4643);
xnor U6521 (N_6521,N_4554,N_5614);
nand U6522 (N_6522,N_4581,N_4962);
nor U6523 (N_6523,N_5388,N_4958);
nor U6524 (N_6524,N_4997,N_4779);
nand U6525 (N_6525,N_5042,N_4610);
xnor U6526 (N_6526,N_5819,N_5796);
or U6527 (N_6527,N_5095,N_5361);
nand U6528 (N_6528,N_5812,N_5919);
xnor U6529 (N_6529,N_5784,N_5286);
nor U6530 (N_6530,N_5648,N_5745);
and U6531 (N_6531,N_4508,N_4738);
and U6532 (N_6532,N_5869,N_5356);
and U6533 (N_6533,N_5555,N_5829);
nor U6534 (N_6534,N_4525,N_5534);
nor U6535 (N_6535,N_5904,N_5285);
and U6536 (N_6536,N_5951,N_4601);
nand U6537 (N_6537,N_4717,N_4853);
nand U6538 (N_6538,N_4506,N_5248);
and U6539 (N_6539,N_4670,N_4764);
or U6540 (N_6540,N_4846,N_5315);
and U6541 (N_6541,N_5950,N_5610);
and U6542 (N_6542,N_4848,N_5893);
and U6543 (N_6543,N_4998,N_4625);
or U6544 (N_6544,N_4722,N_5429);
nor U6545 (N_6545,N_4904,N_4719);
nand U6546 (N_6546,N_4865,N_4627);
nor U6547 (N_6547,N_4765,N_4900);
xnor U6548 (N_6548,N_5453,N_5968);
and U6549 (N_6549,N_4513,N_5936);
nand U6550 (N_6550,N_5606,N_5198);
or U6551 (N_6551,N_5930,N_4621);
or U6552 (N_6552,N_5839,N_4886);
nand U6553 (N_6553,N_4605,N_4776);
and U6554 (N_6554,N_5938,N_5792);
or U6555 (N_6555,N_5044,N_5529);
nor U6556 (N_6556,N_5237,N_5964);
nand U6557 (N_6557,N_4509,N_5087);
or U6558 (N_6558,N_5084,N_5381);
and U6559 (N_6559,N_5405,N_5082);
nor U6560 (N_6560,N_5807,N_5076);
xor U6561 (N_6561,N_5797,N_4921);
or U6562 (N_6562,N_5299,N_5457);
nor U6563 (N_6563,N_5716,N_5292);
nor U6564 (N_6564,N_4530,N_4844);
and U6565 (N_6565,N_5416,N_5884);
nor U6566 (N_6566,N_4969,N_5836);
nand U6567 (N_6567,N_4803,N_5962);
or U6568 (N_6568,N_5467,N_5686);
and U6569 (N_6569,N_4699,N_5563);
nor U6570 (N_6570,N_5015,N_4931);
nand U6571 (N_6571,N_5269,N_5022);
nor U6572 (N_6572,N_4769,N_4909);
or U6573 (N_6573,N_5466,N_4972);
nor U6574 (N_6574,N_5709,N_5078);
and U6575 (N_6575,N_5397,N_5347);
nor U6576 (N_6576,N_5057,N_5511);
or U6577 (N_6577,N_4531,N_4700);
nor U6578 (N_6578,N_5396,N_4723);
and U6579 (N_6579,N_5438,N_5620);
xor U6580 (N_6580,N_5970,N_4882);
and U6581 (N_6581,N_4991,N_5448);
nor U6582 (N_6582,N_5141,N_5707);
or U6583 (N_6583,N_4842,N_5876);
and U6584 (N_6584,N_5917,N_5943);
and U6585 (N_6585,N_5826,N_5984);
or U6586 (N_6586,N_5290,N_5550);
nand U6587 (N_6587,N_4944,N_5798);
nor U6588 (N_6588,N_5441,N_4899);
nor U6589 (N_6589,N_5849,N_5548);
nand U6590 (N_6590,N_4652,N_5901);
nand U6591 (N_6591,N_4979,N_4620);
nor U6592 (N_6592,N_5068,N_4961);
or U6593 (N_6593,N_5866,N_5692);
nand U6594 (N_6594,N_5376,N_5816);
xor U6595 (N_6595,N_5302,N_4592);
nor U6596 (N_6596,N_5066,N_5218);
nor U6597 (N_6597,N_5419,N_4989);
and U6598 (N_6598,N_5711,N_5697);
and U6599 (N_6599,N_5556,N_5460);
and U6600 (N_6600,N_5524,N_5594);
and U6601 (N_6601,N_4928,N_4834);
and U6602 (N_6602,N_5744,N_5590);
xnor U6603 (N_6603,N_4953,N_5914);
nor U6604 (N_6604,N_4688,N_5250);
nor U6605 (N_6605,N_5242,N_4512);
nor U6606 (N_6606,N_5622,N_5251);
nor U6607 (N_6607,N_4703,N_4992);
nand U6608 (N_6608,N_4673,N_5880);
nand U6609 (N_6609,N_5334,N_4641);
and U6610 (N_6610,N_5061,N_5475);
and U6611 (N_6611,N_5301,N_4878);
and U6612 (N_6612,N_5400,N_5191);
xor U6613 (N_6613,N_4543,N_5158);
nand U6614 (N_6614,N_5732,N_4858);
and U6615 (N_6615,N_5600,N_5809);
nand U6616 (N_6616,N_5658,N_5939);
nor U6617 (N_6617,N_5283,N_5367);
xor U6618 (N_6618,N_4784,N_4859);
and U6619 (N_6619,N_4863,N_5280);
nand U6620 (N_6620,N_4672,N_5117);
nor U6621 (N_6621,N_5737,N_5875);
nor U6622 (N_6622,N_5955,N_5461);
nor U6623 (N_6623,N_5760,N_5239);
or U6624 (N_6624,N_4911,N_5599);
and U6625 (N_6625,N_5289,N_5059);
or U6626 (N_6626,N_5014,N_5131);
nand U6627 (N_6627,N_4654,N_5254);
xnor U6628 (N_6628,N_5030,N_5557);
nand U6629 (N_6629,N_5245,N_4697);
nand U6630 (N_6630,N_4888,N_4529);
or U6631 (N_6631,N_4539,N_5579);
and U6632 (N_6632,N_5566,N_5898);
nand U6633 (N_6633,N_4836,N_4503);
and U6634 (N_6634,N_5240,N_5440);
or U6635 (N_6635,N_5018,N_5358);
nor U6636 (N_6636,N_5507,N_5953);
nand U6637 (N_6637,N_5050,N_4877);
and U6638 (N_6638,N_4587,N_5255);
and U6639 (N_6639,N_4999,N_5502);
nand U6640 (N_6640,N_5669,N_5973);
nor U6641 (N_6641,N_5225,N_5165);
and U6642 (N_6642,N_5178,N_5206);
or U6643 (N_6643,N_5041,N_5345);
xor U6644 (N_6644,N_4504,N_4875);
xnor U6645 (N_6645,N_5777,N_4926);
nor U6646 (N_6646,N_5168,N_5634);
or U6647 (N_6647,N_5111,N_5459);
xnor U6648 (N_6648,N_5138,N_5720);
xor U6649 (N_6649,N_5946,N_4734);
or U6650 (N_6650,N_5102,N_5394);
nor U6651 (N_6651,N_5156,N_5348);
nor U6652 (N_6652,N_5028,N_4783);
nand U6653 (N_6653,N_4755,N_5362);
nor U6654 (N_6654,N_5120,N_4918);
or U6655 (N_6655,N_5266,N_5630);
or U6656 (N_6656,N_5167,N_5521);
nand U6657 (N_6657,N_4568,N_5437);
or U6658 (N_6658,N_5680,N_5487);
nand U6659 (N_6659,N_5062,N_5189);
nand U6660 (N_6660,N_5504,N_4905);
nor U6661 (N_6661,N_5677,N_5734);
and U6662 (N_6662,N_5665,N_5414);
or U6663 (N_6663,N_5940,N_5859);
nand U6664 (N_6664,N_5783,N_5988);
nand U6665 (N_6665,N_5498,N_4785);
or U6666 (N_6666,N_4798,N_4696);
and U6667 (N_6667,N_5128,N_5515);
or U6668 (N_6668,N_5589,N_4713);
xnor U6669 (N_6669,N_5490,N_4920);
nand U6670 (N_6670,N_5647,N_5148);
and U6671 (N_6671,N_5545,N_5814);
and U6672 (N_6672,N_4898,N_5423);
and U6673 (N_6673,N_4916,N_5262);
xnor U6674 (N_6674,N_5619,N_5726);
nor U6675 (N_6675,N_4831,N_5911);
and U6676 (N_6676,N_4658,N_5190);
nor U6677 (N_6677,N_5696,N_4971);
nand U6678 (N_6678,N_5431,N_4794);
and U6679 (N_6679,N_5877,N_4777);
and U6680 (N_6680,N_4929,N_5923);
and U6681 (N_6681,N_5232,N_5097);
or U6682 (N_6682,N_4694,N_5114);
or U6683 (N_6683,N_5611,N_5096);
or U6684 (N_6684,N_5011,N_5016);
nor U6685 (N_6685,N_5562,N_4594);
nand U6686 (N_6686,N_4655,N_5417);
or U6687 (N_6687,N_5963,N_5319);
xnor U6688 (N_6688,N_5369,N_5308);
or U6689 (N_6689,N_5618,N_4838);
xnor U6690 (N_6690,N_5411,N_5046);
and U6691 (N_6691,N_5297,N_5800);
or U6692 (N_6692,N_5945,N_5320);
and U6693 (N_6693,N_5771,N_4517);
xor U6694 (N_6694,N_4626,N_5236);
nand U6695 (N_6695,N_5047,N_4948);
xor U6696 (N_6696,N_5587,N_4677);
nand U6697 (N_6697,N_5994,N_4687);
or U6698 (N_6698,N_4600,N_5906);
or U6699 (N_6699,N_5238,N_5768);
and U6700 (N_6700,N_5972,N_5352);
or U6701 (N_6701,N_5415,N_5861);
xor U6702 (N_6702,N_5402,N_5896);
nand U6703 (N_6703,N_4613,N_4573);
nor U6704 (N_6704,N_5169,N_4924);
and U6705 (N_6705,N_5856,N_5127);
xnor U6706 (N_6706,N_4666,N_5104);
or U6707 (N_6707,N_5578,N_5684);
xor U6708 (N_6708,N_5123,N_5257);
and U6709 (N_6709,N_5827,N_5486);
or U6710 (N_6710,N_4945,N_5733);
and U6711 (N_6711,N_5895,N_5398);
nand U6712 (N_6712,N_5840,N_4966);
nor U6713 (N_6713,N_5786,N_4540);
nor U6714 (N_6714,N_4645,N_5736);
nor U6715 (N_6715,N_5227,N_5842);
nand U6716 (N_6716,N_5544,N_4724);
xor U6717 (N_6717,N_5683,N_5531);
or U6718 (N_6718,N_5924,N_4616);
nand U6719 (N_6719,N_5822,N_5862);
nand U6720 (N_6720,N_4534,N_4536);
and U6721 (N_6721,N_5577,N_4501);
or U6722 (N_6722,N_5463,N_5060);
nor U6723 (N_6723,N_5456,N_5595);
and U6724 (N_6724,N_5954,N_4906);
and U6725 (N_6725,N_4829,N_5025);
and U6726 (N_6726,N_5174,N_5222);
nor U6727 (N_6727,N_5660,N_5631);
nand U6728 (N_6728,N_5574,N_5975);
nand U6729 (N_6729,N_5750,N_5693);
nand U6730 (N_6730,N_4754,N_5422);
xor U6731 (N_6731,N_4980,N_4578);
nand U6732 (N_6732,N_5508,N_5134);
xnor U6733 (N_6733,N_5925,N_4596);
nand U6734 (N_6734,N_4634,N_5081);
nor U6735 (N_6735,N_5833,N_5539);
nand U6736 (N_6736,N_5870,N_4939);
or U6737 (N_6737,N_5389,N_5187);
nand U6738 (N_6738,N_5344,N_4771);
xor U6739 (N_6739,N_4753,N_5992);
nand U6740 (N_6740,N_5090,N_5335);
nand U6741 (N_6741,N_5990,N_5613);
and U6742 (N_6742,N_5879,N_5731);
xnor U6743 (N_6743,N_4799,N_4975);
and U6744 (N_6744,N_4750,N_5124);
and U6745 (N_6745,N_4781,N_5470);
and U6746 (N_6746,N_5154,N_5782);
and U6747 (N_6747,N_5054,N_5717);
or U6748 (N_6748,N_5681,N_5652);
xor U6749 (N_6749,N_4861,N_5488);
nor U6750 (N_6750,N_4581,N_4994);
and U6751 (N_6751,N_4716,N_5620);
or U6752 (N_6752,N_5631,N_5080);
and U6753 (N_6753,N_5273,N_5804);
nor U6754 (N_6754,N_4929,N_5295);
nand U6755 (N_6755,N_5050,N_5940);
nand U6756 (N_6756,N_5258,N_4535);
xnor U6757 (N_6757,N_5093,N_4981);
or U6758 (N_6758,N_5979,N_5881);
nand U6759 (N_6759,N_5788,N_5143);
nand U6760 (N_6760,N_5068,N_5617);
and U6761 (N_6761,N_4633,N_4687);
nor U6762 (N_6762,N_4889,N_4940);
nor U6763 (N_6763,N_5354,N_4807);
and U6764 (N_6764,N_5365,N_5399);
xor U6765 (N_6765,N_5820,N_4711);
nand U6766 (N_6766,N_4835,N_5968);
and U6767 (N_6767,N_5448,N_5473);
or U6768 (N_6768,N_5206,N_5803);
xnor U6769 (N_6769,N_5196,N_5299);
and U6770 (N_6770,N_4889,N_5802);
nor U6771 (N_6771,N_5827,N_5153);
or U6772 (N_6772,N_5949,N_5585);
and U6773 (N_6773,N_5698,N_4586);
nor U6774 (N_6774,N_5565,N_4864);
or U6775 (N_6775,N_5620,N_5805);
and U6776 (N_6776,N_4886,N_5983);
nand U6777 (N_6777,N_5976,N_5380);
xnor U6778 (N_6778,N_5986,N_4581);
or U6779 (N_6779,N_4903,N_5234);
and U6780 (N_6780,N_5186,N_5420);
nand U6781 (N_6781,N_5498,N_5413);
and U6782 (N_6782,N_5287,N_5925);
nand U6783 (N_6783,N_4984,N_4942);
or U6784 (N_6784,N_5741,N_5219);
nor U6785 (N_6785,N_5462,N_5018);
nand U6786 (N_6786,N_5759,N_4676);
nor U6787 (N_6787,N_4756,N_5033);
nor U6788 (N_6788,N_5993,N_4954);
or U6789 (N_6789,N_5318,N_5295);
and U6790 (N_6790,N_5386,N_5476);
nor U6791 (N_6791,N_4676,N_4912);
and U6792 (N_6792,N_5719,N_5245);
nor U6793 (N_6793,N_4953,N_5934);
or U6794 (N_6794,N_4929,N_5272);
and U6795 (N_6795,N_5266,N_4501);
or U6796 (N_6796,N_5191,N_5125);
or U6797 (N_6797,N_5062,N_5256);
nand U6798 (N_6798,N_5050,N_4948);
or U6799 (N_6799,N_4845,N_5364);
or U6800 (N_6800,N_5829,N_4830);
nand U6801 (N_6801,N_5439,N_5321);
and U6802 (N_6802,N_5996,N_4684);
and U6803 (N_6803,N_5759,N_4750);
nor U6804 (N_6804,N_5988,N_4799);
and U6805 (N_6805,N_5184,N_5952);
or U6806 (N_6806,N_5371,N_5764);
and U6807 (N_6807,N_4537,N_5966);
xor U6808 (N_6808,N_5917,N_5734);
or U6809 (N_6809,N_4967,N_5377);
nand U6810 (N_6810,N_4536,N_4605);
nand U6811 (N_6811,N_5961,N_4588);
and U6812 (N_6812,N_4575,N_5456);
and U6813 (N_6813,N_5390,N_5440);
nor U6814 (N_6814,N_5332,N_5885);
nand U6815 (N_6815,N_5414,N_4732);
xor U6816 (N_6816,N_5285,N_5506);
nand U6817 (N_6817,N_5335,N_5608);
and U6818 (N_6818,N_5987,N_5970);
or U6819 (N_6819,N_4758,N_5589);
or U6820 (N_6820,N_4944,N_4721);
nand U6821 (N_6821,N_5535,N_5360);
nor U6822 (N_6822,N_5394,N_5675);
xnor U6823 (N_6823,N_5147,N_4873);
and U6824 (N_6824,N_5806,N_5049);
xnor U6825 (N_6825,N_5839,N_5724);
and U6826 (N_6826,N_5861,N_4686);
nand U6827 (N_6827,N_5441,N_5631);
nor U6828 (N_6828,N_5214,N_5723);
and U6829 (N_6829,N_5888,N_4870);
xor U6830 (N_6830,N_4882,N_5462);
nand U6831 (N_6831,N_5156,N_5368);
nand U6832 (N_6832,N_5945,N_5442);
xnor U6833 (N_6833,N_5685,N_4790);
and U6834 (N_6834,N_5375,N_4626);
xnor U6835 (N_6835,N_4704,N_5973);
nor U6836 (N_6836,N_5756,N_4559);
xnor U6837 (N_6837,N_5218,N_5132);
xor U6838 (N_6838,N_5623,N_5885);
nand U6839 (N_6839,N_4750,N_5278);
nand U6840 (N_6840,N_4819,N_5818);
and U6841 (N_6841,N_5979,N_5264);
or U6842 (N_6842,N_5757,N_5483);
xor U6843 (N_6843,N_4608,N_4898);
xnor U6844 (N_6844,N_5015,N_5724);
nand U6845 (N_6845,N_4566,N_5201);
and U6846 (N_6846,N_5150,N_5583);
nor U6847 (N_6847,N_4789,N_5233);
xnor U6848 (N_6848,N_4930,N_5014);
or U6849 (N_6849,N_5697,N_5233);
nand U6850 (N_6850,N_5874,N_5833);
xor U6851 (N_6851,N_4623,N_4829);
xor U6852 (N_6852,N_5950,N_5618);
nor U6853 (N_6853,N_5417,N_5262);
and U6854 (N_6854,N_5415,N_5926);
nor U6855 (N_6855,N_5229,N_5119);
nor U6856 (N_6856,N_5467,N_5563);
nor U6857 (N_6857,N_4782,N_4904);
and U6858 (N_6858,N_4540,N_4616);
or U6859 (N_6859,N_5806,N_5628);
and U6860 (N_6860,N_5635,N_4727);
nor U6861 (N_6861,N_5237,N_5990);
xnor U6862 (N_6862,N_5629,N_4512);
nor U6863 (N_6863,N_4954,N_5368);
nor U6864 (N_6864,N_4542,N_5807);
and U6865 (N_6865,N_5580,N_5602);
nand U6866 (N_6866,N_5477,N_4886);
xnor U6867 (N_6867,N_5886,N_4731);
xor U6868 (N_6868,N_5165,N_5846);
nor U6869 (N_6869,N_4760,N_5782);
and U6870 (N_6870,N_5405,N_4504);
nor U6871 (N_6871,N_5110,N_5242);
or U6872 (N_6872,N_5234,N_5973);
or U6873 (N_6873,N_5821,N_5351);
and U6874 (N_6874,N_5163,N_4952);
nand U6875 (N_6875,N_5844,N_4850);
or U6876 (N_6876,N_4523,N_5188);
or U6877 (N_6877,N_5308,N_5070);
xor U6878 (N_6878,N_5462,N_5055);
or U6879 (N_6879,N_5201,N_4767);
or U6880 (N_6880,N_4922,N_5139);
nor U6881 (N_6881,N_5634,N_5862);
nand U6882 (N_6882,N_5678,N_5470);
nor U6883 (N_6883,N_5216,N_5743);
nand U6884 (N_6884,N_4695,N_4982);
xnor U6885 (N_6885,N_4958,N_4895);
or U6886 (N_6886,N_5021,N_5522);
xor U6887 (N_6887,N_4947,N_4981);
or U6888 (N_6888,N_5063,N_4904);
nand U6889 (N_6889,N_5625,N_5233);
xor U6890 (N_6890,N_4536,N_5729);
xor U6891 (N_6891,N_5473,N_5256);
and U6892 (N_6892,N_5461,N_5772);
nor U6893 (N_6893,N_5446,N_5653);
xor U6894 (N_6894,N_4580,N_5192);
nor U6895 (N_6895,N_5642,N_5375);
and U6896 (N_6896,N_5126,N_4991);
xor U6897 (N_6897,N_5223,N_4888);
xnor U6898 (N_6898,N_5351,N_5695);
and U6899 (N_6899,N_4599,N_4966);
nor U6900 (N_6900,N_5418,N_5392);
nor U6901 (N_6901,N_4798,N_5419);
xor U6902 (N_6902,N_5632,N_5433);
and U6903 (N_6903,N_4741,N_4686);
xor U6904 (N_6904,N_4704,N_5816);
nor U6905 (N_6905,N_5242,N_4955);
or U6906 (N_6906,N_5107,N_4550);
or U6907 (N_6907,N_5436,N_5844);
nand U6908 (N_6908,N_5707,N_5010);
nor U6909 (N_6909,N_5601,N_5353);
xnor U6910 (N_6910,N_5635,N_5452);
or U6911 (N_6911,N_5634,N_5543);
or U6912 (N_6912,N_5577,N_5741);
nand U6913 (N_6913,N_5622,N_4636);
nand U6914 (N_6914,N_4967,N_5445);
nor U6915 (N_6915,N_4743,N_4626);
nand U6916 (N_6916,N_4574,N_5978);
nor U6917 (N_6917,N_5485,N_5102);
nand U6918 (N_6918,N_4549,N_5828);
and U6919 (N_6919,N_4622,N_4708);
nor U6920 (N_6920,N_5302,N_4818);
xor U6921 (N_6921,N_5613,N_5237);
xor U6922 (N_6922,N_4924,N_5378);
nand U6923 (N_6923,N_5595,N_4943);
nand U6924 (N_6924,N_5549,N_4797);
and U6925 (N_6925,N_5589,N_5991);
nor U6926 (N_6926,N_5540,N_5300);
and U6927 (N_6927,N_5321,N_5652);
nor U6928 (N_6928,N_5842,N_5126);
and U6929 (N_6929,N_4540,N_5920);
nor U6930 (N_6930,N_4930,N_5764);
and U6931 (N_6931,N_4833,N_5722);
xnor U6932 (N_6932,N_5264,N_4841);
or U6933 (N_6933,N_4612,N_4847);
or U6934 (N_6934,N_5007,N_5257);
nand U6935 (N_6935,N_4829,N_4518);
nand U6936 (N_6936,N_5685,N_5370);
xnor U6937 (N_6937,N_5398,N_5280);
nand U6938 (N_6938,N_4912,N_4979);
nand U6939 (N_6939,N_5829,N_4951);
nor U6940 (N_6940,N_5598,N_5208);
nor U6941 (N_6941,N_5702,N_5019);
and U6942 (N_6942,N_5874,N_5262);
and U6943 (N_6943,N_4526,N_5125);
nor U6944 (N_6944,N_4802,N_4876);
nor U6945 (N_6945,N_4828,N_5419);
or U6946 (N_6946,N_4556,N_4660);
or U6947 (N_6947,N_5801,N_5131);
xor U6948 (N_6948,N_4859,N_4932);
nand U6949 (N_6949,N_4930,N_5960);
and U6950 (N_6950,N_5502,N_5537);
and U6951 (N_6951,N_5624,N_5999);
and U6952 (N_6952,N_5586,N_5059);
and U6953 (N_6953,N_5039,N_5668);
nand U6954 (N_6954,N_4642,N_5481);
nand U6955 (N_6955,N_5860,N_4914);
nor U6956 (N_6956,N_4917,N_4866);
or U6957 (N_6957,N_5068,N_5182);
nor U6958 (N_6958,N_5464,N_4869);
nand U6959 (N_6959,N_4635,N_5649);
xor U6960 (N_6960,N_4727,N_5188);
nor U6961 (N_6961,N_5106,N_5603);
xor U6962 (N_6962,N_4943,N_5543);
xor U6963 (N_6963,N_5267,N_4650);
and U6964 (N_6964,N_5663,N_5130);
xnor U6965 (N_6965,N_5641,N_4991);
nor U6966 (N_6966,N_5545,N_4742);
nor U6967 (N_6967,N_5782,N_5837);
xor U6968 (N_6968,N_5429,N_4890);
nand U6969 (N_6969,N_4602,N_4679);
or U6970 (N_6970,N_4715,N_5316);
nand U6971 (N_6971,N_5592,N_4803);
or U6972 (N_6972,N_5935,N_4635);
xnor U6973 (N_6973,N_5870,N_4731);
xnor U6974 (N_6974,N_5603,N_5553);
and U6975 (N_6975,N_5828,N_4773);
nand U6976 (N_6976,N_5006,N_5887);
or U6977 (N_6977,N_5975,N_5180);
and U6978 (N_6978,N_4598,N_5392);
nand U6979 (N_6979,N_5522,N_4667);
and U6980 (N_6980,N_5607,N_4535);
xnor U6981 (N_6981,N_5205,N_4520);
xnor U6982 (N_6982,N_5978,N_5211);
or U6983 (N_6983,N_4978,N_5601);
or U6984 (N_6984,N_5473,N_5161);
xnor U6985 (N_6985,N_4788,N_4554);
and U6986 (N_6986,N_5888,N_4867);
xor U6987 (N_6987,N_5571,N_4723);
and U6988 (N_6988,N_4979,N_4755);
xnor U6989 (N_6989,N_5486,N_5593);
xnor U6990 (N_6990,N_5696,N_5269);
nand U6991 (N_6991,N_4501,N_4577);
or U6992 (N_6992,N_4810,N_5350);
or U6993 (N_6993,N_5075,N_4786);
xor U6994 (N_6994,N_4509,N_5923);
and U6995 (N_6995,N_5259,N_5591);
xor U6996 (N_6996,N_4749,N_5502);
or U6997 (N_6997,N_4909,N_4799);
nand U6998 (N_6998,N_4712,N_4560);
and U6999 (N_6999,N_5429,N_5350);
and U7000 (N_7000,N_5830,N_4924);
or U7001 (N_7001,N_4572,N_5180);
xnor U7002 (N_7002,N_5336,N_4578);
nor U7003 (N_7003,N_5454,N_5614);
or U7004 (N_7004,N_5243,N_4514);
nor U7005 (N_7005,N_4546,N_5933);
nand U7006 (N_7006,N_4539,N_5387);
and U7007 (N_7007,N_5733,N_5721);
or U7008 (N_7008,N_5758,N_4603);
and U7009 (N_7009,N_5306,N_5781);
and U7010 (N_7010,N_5504,N_5410);
or U7011 (N_7011,N_4897,N_5761);
nor U7012 (N_7012,N_5574,N_5129);
nand U7013 (N_7013,N_5510,N_4590);
and U7014 (N_7014,N_5436,N_5095);
and U7015 (N_7015,N_5388,N_5040);
xnor U7016 (N_7016,N_5834,N_5368);
xnor U7017 (N_7017,N_5133,N_4948);
xor U7018 (N_7018,N_5897,N_5066);
nor U7019 (N_7019,N_5441,N_4673);
or U7020 (N_7020,N_5594,N_5848);
or U7021 (N_7021,N_5348,N_4858);
xnor U7022 (N_7022,N_5363,N_5702);
or U7023 (N_7023,N_5227,N_5772);
xnor U7024 (N_7024,N_4896,N_5004);
nor U7025 (N_7025,N_5231,N_5837);
nand U7026 (N_7026,N_5734,N_5921);
xnor U7027 (N_7027,N_5351,N_5079);
and U7028 (N_7028,N_5129,N_5193);
xor U7029 (N_7029,N_5755,N_4714);
nand U7030 (N_7030,N_5779,N_4553);
nand U7031 (N_7031,N_4663,N_4858);
or U7032 (N_7032,N_5525,N_5504);
or U7033 (N_7033,N_5572,N_5548);
xor U7034 (N_7034,N_4563,N_4948);
nor U7035 (N_7035,N_5072,N_5663);
nand U7036 (N_7036,N_5828,N_5287);
nand U7037 (N_7037,N_5641,N_5057);
and U7038 (N_7038,N_5738,N_5933);
nor U7039 (N_7039,N_5599,N_5854);
and U7040 (N_7040,N_5108,N_5116);
nor U7041 (N_7041,N_4543,N_5457);
nor U7042 (N_7042,N_5119,N_4714);
xnor U7043 (N_7043,N_5761,N_5405);
or U7044 (N_7044,N_5762,N_5491);
nor U7045 (N_7045,N_5896,N_5993);
xor U7046 (N_7046,N_4694,N_5253);
and U7047 (N_7047,N_4536,N_5350);
and U7048 (N_7048,N_4552,N_5710);
xnor U7049 (N_7049,N_5564,N_5582);
xnor U7050 (N_7050,N_5451,N_4662);
or U7051 (N_7051,N_5846,N_5213);
or U7052 (N_7052,N_4519,N_5989);
xnor U7053 (N_7053,N_5850,N_4875);
or U7054 (N_7054,N_5037,N_5935);
nand U7055 (N_7055,N_5753,N_5145);
or U7056 (N_7056,N_5294,N_4789);
nand U7057 (N_7057,N_4647,N_5460);
or U7058 (N_7058,N_5308,N_4889);
nor U7059 (N_7059,N_5708,N_4716);
and U7060 (N_7060,N_4691,N_4530);
nor U7061 (N_7061,N_5497,N_4817);
and U7062 (N_7062,N_4713,N_5089);
and U7063 (N_7063,N_4703,N_5631);
or U7064 (N_7064,N_5457,N_5812);
xnor U7065 (N_7065,N_5860,N_5313);
nor U7066 (N_7066,N_5034,N_4919);
and U7067 (N_7067,N_4638,N_4534);
xor U7068 (N_7068,N_5645,N_5734);
xor U7069 (N_7069,N_5696,N_4818);
nand U7070 (N_7070,N_5122,N_5414);
and U7071 (N_7071,N_5261,N_4595);
xnor U7072 (N_7072,N_5729,N_5378);
xnor U7073 (N_7073,N_5119,N_5240);
nor U7074 (N_7074,N_5023,N_5194);
nor U7075 (N_7075,N_5809,N_4604);
nor U7076 (N_7076,N_4612,N_4891);
nand U7077 (N_7077,N_5431,N_4606);
or U7078 (N_7078,N_4677,N_4665);
nor U7079 (N_7079,N_4729,N_4607);
and U7080 (N_7080,N_5447,N_5000);
xnor U7081 (N_7081,N_4992,N_5759);
nand U7082 (N_7082,N_5223,N_5755);
nor U7083 (N_7083,N_5175,N_4892);
or U7084 (N_7084,N_5142,N_4864);
and U7085 (N_7085,N_4759,N_5476);
nand U7086 (N_7086,N_5057,N_5753);
nand U7087 (N_7087,N_4868,N_4658);
nand U7088 (N_7088,N_5952,N_5460);
nand U7089 (N_7089,N_4913,N_5600);
xnor U7090 (N_7090,N_5988,N_5661);
nor U7091 (N_7091,N_4629,N_4510);
xor U7092 (N_7092,N_5186,N_5161);
and U7093 (N_7093,N_5383,N_4742);
nor U7094 (N_7094,N_5050,N_4658);
xnor U7095 (N_7095,N_4941,N_5479);
nor U7096 (N_7096,N_4530,N_5032);
xor U7097 (N_7097,N_4990,N_5173);
xor U7098 (N_7098,N_5879,N_5150);
xnor U7099 (N_7099,N_4707,N_5960);
nor U7100 (N_7100,N_4965,N_5481);
xor U7101 (N_7101,N_5240,N_5278);
nor U7102 (N_7102,N_5174,N_5296);
nand U7103 (N_7103,N_5480,N_5919);
nor U7104 (N_7104,N_4709,N_5650);
or U7105 (N_7105,N_5915,N_4702);
xnor U7106 (N_7106,N_4761,N_4765);
nor U7107 (N_7107,N_5564,N_4514);
or U7108 (N_7108,N_5853,N_5652);
nor U7109 (N_7109,N_5184,N_5687);
nand U7110 (N_7110,N_5604,N_4887);
xnor U7111 (N_7111,N_4944,N_5864);
or U7112 (N_7112,N_5096,N_5837);
nor U7113 (N_7113,N_4742,N_4960);
or U7114 (N_7114,N_5077,N_4858);
and U7115 (N_7115,N_4696,N_4544);
nand U7116 (N_7116,N_5115,N_5064);
nor U7117 (N_7117,N_4554,N_5809);
or U7118 (N_7118,N_5306,N_5450);
nor U7119 (N_7119,N_4952,N_4716);
nand U7120 (N_7120,N_4547,N_5845);
nand U7121 (N_7121,N_5857,N_5569);
nor U7122 (N_7122,N_5319,N_4932);
or U7123 (N_7123,N_5624,N_5348);
nor U7124 (N_7124,N_5896,N_5872);
or U7125 (N_7125,N_5810,N_4520);
and U7126 (N_7126,N_5506,N_5521);
and U7127 (N_7127,N_5176,N_5822);
or U7128 (N_7128,N_4751,N_5764);
nor U7129 (N_7129,N_5588,N_5350);
nand U7130 (N_7130,N_5738,N_5433);
or U7131 (N_7131,N_5311,N_5338);
xnor U7132 (N_7132,N_5345,N_5557);
nand U7133 (N_7133,N_5827,N_4791);
and U7134 (N_7134,N_4768,N_5287);
nand U7135 (N_7135,N_5143,N_4662);
and U7136 (N_7136,N_5797,N_5364);
nand U7137 (N_7137,N_5730,N_5018);
nand U7138 (N_7138,N_5543,N_4514);
or U7139 (N_7139,N_4999,N_4975);
and U7140 (N_7140,N_5619,N_5599);
nand U7141 (N_7141,N_5419,N_5186);
nor U7142 (N_7142,N_5738,N_4853);
xor U7143 (N_7143,N_5360,N_4569);
or U7144 (N_7144,N_4742,N_5256);
and U7145 (N_7145,N_5841,N_5733);
nand U7146 (N_7146,N_5968,N_5498);
nand U7147 (N_7147,N_4597,N_5351);
nor U7148 (N_7148,N_5160,N_5576);
nor U7149 (N_7149,N_4525,N_5848);
nor U7150 (N_7150,N_5859,N_5581);
xor U7151 (N_7151,N_4533,N_5310);
xor U7152 (N_7152,N_5867,N_4782);
xnor U7153 (N_7153,N_5860,N_5249);
nand U7154 (N_7154,N_5887,N_4669);
xor U7155 (N_7155,N_5105,N_5252);
and U7156 (N_7156,N_5581,N_5176);
xnor U7157 (N_7157,N_5202,N_4922);
xnor U7158 (N_7158,N_5517,N_5677);
nand U7159 (N_7159,N_5684,N_5222);
nand U7160 (N_7160,N_4773,N_4812);
nor U7161 (N_7161,N_5443,N_4607);
and U7162 (N_7162,N_5732,N_5059);
nand U7163 (N_7163,N_4985,N_5000);
nand U7164 (N_7164,N_5533,N_5290);
and U7165 (N_7165,N_4701,N_5884);
nor U7166 (N_7166,N_5220,N_5395);
and U7167 (N_7167,N_5081,N_5242);
or U7168 (N_7168,N_5450,N_4776);
xor U7169 (N_7169,N_5643,N_5462);
nand U7170 (N_7170,N_4733,N_5240);
and U7171 (N_7171,N_5798,N_5699);
xnor U7172 (N_7172,N_5957,N_4807);
or U7173 (N_7173,N_5200,N_5197);
nor U7174 (N_7174,N_5546,N_5417);
nor U7175 (N_7175,N_5660,N_5887);
and U7176 (N_7176,N_5061,N_5173);
nand U7177 (N_7177,N_5606,N_5136);
or U7178 (N_7178,N_5249,N_4547);
or U7179 (N_7179,N_4692,N_4501);
xnor U7180 (N_7180,N_5284,N_4836);
nor U7181 (N_7181,N_4645,N_5290);
nor U7182 (N_7182,N_5590,N_4942);
nand U7183 (N_7183,N_4578,N_5411);
nor U7184 (N_7184,N_4517,N_5746);
and U7185 (N_7185,N_5364,N_5429);
and U7186 (N_7186,N_4696,N_5573);
nor U7187 (N_7187,N_5619,N_4932);
xor U7188 (N_7188,N_4732,N_5836);
nand U7189 (N_7189,N_5612,N_5770);
nor U7190 (N_7190,N_5593,N_4662);
xor U7191 (N_7191,N_4729,N_4817);
and U7192 (N_7192,N_4607,N_4781);
xnor U7193 (N_7193,N_5359,N_5809);
and U7194 (N_7194,N_5449,N_5086);
xor U7195 (N_7195,N_5019,N_4704);
xor U7196 (N_7196,N_5683,N_5239);
or U7197 (N_7197,N_5515,N_4657);
nor U7198 (N_7198,N_5713,N_5085);
or U7199 (N_7199,N_5737,N_5162);
nor U7200 (N_7200,N_5810,N_4779);
or U7201 (N_7201,N_5526,N_5244);
nand U7202 (N_7202,N_5118,N_5012);
nor U7203 (N_7203,N_4543,N_5582);
or U7204 (N_7204,N_4660,N_4519);
nor U7205 (N_7205,N_4760,N_5832);
nor U7206 (N_7206,N_4503,N_5213);
nand U7207 (N_7207,N_5218,N_5469);
and U7208 (N_7208,N_4794,N_4618);
nor U7209 (N_7209,N_5794,N_5235);
or U7210 (N_7210,N_5390,N_4517);
nand U7211 (N_7211,N_5587,N_4568);
nand U7212 (N_7212,N_5276,N_5321);
and U7213 (N_7213,N_4532,N_5843);
nand U7214 (N_7214,N_5512,N_4650);
nor U7215 (N_7215,N_4611,N_5097);
or U7216 (N_7216,N_5344,N_5024);
nor U7217 (N_7217,N_5922,N_5694);
nand U7218 (N_7218,N_5036,N_5176);
or U7219 (N_7219,N_4963,N_4725);
xnor U7220 (N_7220,N_4892,N_4826);
and U7221 (N_7221,N_4513,N_4753);
nand U7222 (N_7222,N_4954,N_4581);
nor U7223 (N_7223,N_4890,N_4543);
nor U7224 (N_7224,N_5965,N_4768);
and U7225 (N_7225,N_5290,N_4723);
nand U7226 (N_7226,N_5889,N_5478);
nor U7227 (N_7227,N_5764,N_5688);
nand U7228 (N_7228,N_4882,N_4580);
nor U7229 (N_7229,N_5266,N_5276);
nand U7230 (N_7230,N_5859,N_4999);
and U7231 (N_7231,N_5909,N_4806);
nand U7232 (N_7232,N_5401,N_5884);
or U7233 (N_7233,N_5698,N_5529);
nand U7234 (N_7234,N_5314,N_4685);
and U7235 (N_7235,N_5805,N_4758);
or U7236 (N_7236,N_4622,N_4516);
nor U7237 (N_7237,N_4851,N_5135);
and U7238 (N_7238,N_4545,N_5198);
nor U7239 (N_7239,N_5114,N_5714);
nand U7240 (N_7240,N_4681,N_4974);
xnor U7241 (N_7241,N_4736,N_5172);
or U7242 (N_7242,N_4597,N_5762);
or U7243 (N_7243,N_5383,N_4776);
nor U7244 (N_7244,N_5947,N_5011);
nor U7245 (N_7245,N_5336,N_5225);
nand U7246 (N_7246,N_5975,N_4948);
nor U7247 (N_7247,N_5656,N_4616);
and U7248 (N_7248,N_5837,N_4841);
and U7249 (N_7249,N_5263,N_5496);
and U7250 (N_7250,N_5393,N_5338);
or U7251 (N_7251,N_4648,N_5069);
or U7252 (N_7252,N_5323,N_4893);
nand U7253 (N_7253,N_5610,N_5995);
nand U7254 (N_7254,N_4675,N_5819);
nor U7255 (N_7255,N_5511,N_4976);
xnor U7256 (N_7256,N_5604,N_5431);
xnor U7257 (N_7257,N_4569,N_5850);
nor U7258 (N_7258,N_5507,N_5267);
xor U7259 (N_7259,N_5630,N_5650);
nand U7260 (N_7260,N_4641,N_4991);
or U7261 (N_7261,N_4743,N_4671);
nor U7262 (N_7262,N_4510,N_5512);
xnor U7263 (N_7263,N_4840,N_5647);
or U7264 (N_7264,N_5896,N_5738);
xor U7265 (N_7265,N_5102,N_5337);
nand U7266 (N_7266,N_5764,N_5269);
xnor U7267 (N_7267,N_5078,N_5463);
nand U7268 (N_7268,N_5586,N_4596);
nand U7269 (N_7269,N_5486,N_4994);
and U7270 (N_7270,N_5964,N_5666);
nand U7271 (N_7271,N_5593,N_5974);
nor U7272 (N_7272,N_4918,N_5994);
xor U7273 (N_7273,N_5800,N_4638);
nor U7274 (N_7274,N_4843,N_5715);
or U7275 (N_7275,N_5651,N_5517);
or U7276 (N_7276,N_5620,N_4639);
xnor U7277 (N_7277,N_4830,N_4665);
and U7278 (N_7278,N_4835,N_4591);
nor U7279 (N_7279,N_5610,N_4653);
nor U7280 (N_7280,N_4731,N_4681);
xor U7281 (N_7281,N_5459,N_4814);
or U7282 (N_7282,N_4527,N_5895);
xor U7283 (N_7283,N_5291,N_5166);
xor U7284 (N_7284,N_5871,N_4874);
nand U7285 (N_7285,N_4506,N_4619);
or U7286 (N_7286,N_4700,N_4893);
and U7287 (N_7287,N_5907,N_4534);
nor U7288 (N_7288,N_5810,N_5505);
and U7289 (N_7289,N_5094,N_4787);
nor U7290 (N_7290,N_4750,N_4741);
xnor U7291 (N_7291,N_4957,N_5138);
or U7292 (N_7292,N_5012,N_5815);
nor U7293 (N_7293,N_5632,N_4500);
xor U7294 (N_7294,N_5630,N_4970);
nor U7295 (N_7295,N_4744,N_5671);
and U7296 (N_7296,N_5233,N_5681);
nor U7297 (N_7297,N_4931,N_5774);
and U7298 (N_7298,N_5260,N_5830);
and U7299 (N_7299,N_5272,N_5309);
or U7300 (N_7300,N_5959,N_4702);
nand U7301 (N_7301,N_5573,N_5197);
nor U7302 (N_7302,N_4525,N_4740);
nand U7303 (N_7303,N_4686,N_5474);
nand U7304 (N_7304,N_4752,N_5152);
xnor U7305 (N_7305,N_5980,N_5873);
nor U7306 (N_7306,N_5070,N_5471);
nor U7307 (N_7307,N_4689,N_5463);
xnor U7308 (N_7308,N_5262,N_5242);
and U7309 (N_7309,N_5483,N_4789);
xor U7310 (N_7310,N_4886,N_5744);
nand U7311 (N_7311,N_5766,N_5826);
or U7312 (N_7312,N_5231,N_4780);
and U7313 (N_7313,N_4723,N_4671);
or U7314 (N_7314,N_5447,N_5465);
and U7315 (N_7315,N_4681,N_5996);
and U7316 (N_7316,N_5028,N_4905);
xnor U7317 (N_7317,N_5470,N_5751);
or U7318 (N_7318,N_4639,N_5987);
or U7319 (N_7319,N_5036,N_5640);
nand U7320 (N_7320,N_4528,N_5144);
xor U7321 (N_7321,N_4574,N_5193);
xnor U7322 (N_7322,N_5752,N_5422);
or U7323 (N_7323,N_5232,N_5431);
nand U7324 (N_7324,N_4586,N_4596);
or U7325 (N_7325,N_5073,N_5790);
nand U7326 (N_7326,N_5731,N_4663);
nor U7327 (N_7327,N_4663,N_5917);
nand U7328 (N_7328,N_4568,N_4703);
nor U7329 (N_7329,N_5254,N_5828);
or U7330 (N_7330,N_5251,N_5417);
xor U7331 (N_7331,N_5993,N_4660);
nor U7332 (N_7332,N_4885,N_5488);
or U7333 (N_7333,N_4941,N_5378);
nand U7334 (N_7334,N_5951,N_5945);
nor U7335 (N_7335,N_5656,N_4993);
xnor U7336 (N_7336,N_4851,N_4848);
nor U7337 (N_7337,N_4991,N_5402);
nand U7338 (N_7338,N_5118,N_5767);
or U7339 (N_7339,N_5899,N_4957);
or U7340 (N_7340,N_5416,N_5983);
and U7341 (N_7341,N_5847,N_5129);
or U7342 (N_7342,N_5029,N_4703);
or U7343 (N_7343,N_5325,N_5692);
xor U7344 (N_7344,N_4568,N_5684);
nor U7345 (N_7345,N_5574,N_5942);
xor U7346 (N_7346,N_5604,N_5008);
xnor U7347 (N_7347,N_5679,N_5489);
nor U7348 (N_7348,N_4599,N_5932);
nand U7349 (N_7349,N_5796,N_5235);
and U7350 (N_7350,N_5382,N_4628);
nor U7351 (N_7351,N_5383,N_4561);
nor U7352 (N_7352,N_5617,N_5417);
nand U7353 (N_7353,N_5670,N_4581);
xor U7354 (N_7354,N_5943,N_5381);
xnor U7355 (N_7355,N_5158,N_5524);
nor U7356 (N_7356,N_4616,N_4951);
and U7357 (N_7357,N_4554,N_4572);
nor U7358 (N_7358,N_5531,N_4923);
xnor U7359 (N_7359,N_5467,N_5580);
nor U7360 (N_7360,N_4593,N_5172);
or U7361 (N_7361,N_5665,N_5386);
and U7362 (N_7362,N_5747,N_5932);
or U7363 (N_7363,N_5302,N_4938);
nand U7364 (N_7364,N_4729,N_5619);
xor U7365 (N_7365,N_5277,N_4881);
nand U7366 (N_7366,N_4940,N_4615);
nand U7367 (N_7367,N_5590,N_4582);
xor U7368 (N_7368,N_5864,N_4687);
xnor U7369 (N_7369,N_5068,N_5700);
or U7370 (N_7370,N_5331,N_4531);
nand U7371 (N_7371,N_5615,N_5180);
and U7372 (N_7372,N_5922,N_5364);
xnor U7373 (N_7373,N_5139,N_5639);
xnor U7374 (N_7374,N_4566,N_5669);
or U7375 (N_7375,N_4637,N_5954);
nor U7376 (N_7376,N_4765,N_4972);
xor U7377 (N_7377,N_5150,N_5012);
nand U7378 (N_7378,N_5108,N_5295);
and U7379 (N_7379,N_4717,N_5281);
nand U7380 (N_7380,N_5371,N_5626);
and U7381 (N_7381,N_5631,N_5564);
and U7382 (N_7382,N_4715,N_5546);
or U7383 (N_7383,N_5788,N_5805);
xor U7384 (N_7384,N_5279,N_5999);
and U7385 (N_7385,N_5926,N_5372);
xnor U7386 (N_7386,N_4853,N_5338);
and U7387 (N_7387,N_5391,N_5078);
nor U7388 (N_7388,N_5186,N_5731);
or U7389 (N_7389,N_5819,N_5762);
nor U7390 (N_7390,N_4902,N_5348);
xor U7391 (N_7391,N_4720,N_4736);
or U7392 (N_7392,N_4973,N_5119);
and U7393 (N_7393,N_5336,N_5759);
nand U7394 (N_7394,N_4892,N_5858);
nor U7395 (N_7395,N_5644,N_5921);
or U7396 (N_7396,N_5983,N_5614);
or U7397 (N_7397,N_4770,N_5906);
xor U7398 (N_7398,N_4704,N_4723);
or U7399 (N_7399,N_5184,N_5197);
nor U7400 (N_7400,N_4852,N_5451);
nand U7401 (N_7401,N_4999,N_4617);
and U7402 (N_7402,N_5625,N_5033);
and U7403 (N_7403,N_4672,N_4619);
nand U7404 (N_7404,N_4597,N_4962);
and U7405 (N_7405,N_4899,N_5468);
and U7406 (N_7406,N_5763,N_5040);
and U7407 (N_7407,N_5515,N_5705);
nor U7408 (N_7408,N_5927,N_5031);
nand U7409 (N_7409,N_5819,N_4663);
and U7410 (N_7410,N_5859,N_5080);
nor U7411 (N_7411,N_5783,N_5564);
or U7412 (N_7412,N_5674,N_4857);
nand U7413 (N_7413,N_5010,N_5789);
nor U7414 (N_7414,N_4516,N_5283);
nand U7415 (N_7415,N_5180,N_5133);
or U7416 (N_7416,N_5360,N_5802);
or U7417 (N_7417,N_5764,N_4805);
nor U7418 (N_7418,N_5758,N_4790);
xnor U7419 (N_7419,N_4893,N_5960);
xor U7420 (N_7420,N_4859,N_5895);
and U7421 (N_7421,N_5199,N_5971);
nor U7422 (N_7422,N_5466,N_4598);
or U7423 (N_7423,N_4899,N_4659);
and U7424 (N_7424,N_5352,N_4515);
and U7425 (N_7425,N_5457,N_4760);
nor U7426 (N_7426,N_4734,N_5128);
nand U7427 (N_7427,N_5298,N_5212);
and U7428 (N_7428,N_5150,N_5528);
xnor U7429 (N_7429,N_4728,N_5954);
nor U7430 (N_7430,N_5525,N_5329);
nor U7431 (N_7431,N_5048,N_5334);
or U7432 (N_7432,N_5128,N_5179);
and U7433 (N_7433,N_4768,N_5060);
xor U7434 (N_7434,N_5257,N_5778);
nor U7435 (N_7435,N_5162,N_4820);
nand U7436 (N_7436,N_5184,N_5051);
xnor U7437 (N_7437,N_5408,N_5983);
nor U7438 (N_7438,N_5324,N_5335);
nor U7439 (N_7439,N_4855,N_5528);
nor U7440 (N_7440,N_5449,N_4588);
nor U7441 (N_7441,N_4723,N_5199);
nand U7442 (N_7442,N_4739,N_5026);
nor U7443 (N_7443,N_5569,N_5197);
and U7444 (N_7444,N_5941,N_4840);
and U7445 (N_7445,N_5742,N_5296);
xor U7446 (N_7446,N_5369,N_4785);
and U7447 (N_7447,N_5726,N_5112);
xor U7448 (N_7448,N_5498,N_4622);
and U7449 (N_7449,N_5255,N_5968);
and U7450 (N_7450,N_5350,N_5956);
and U7451 (N_7451,N_5353,N_4635);
xor U7452 (N_7452,N_4581,N_5955);
xnor U7453 (N_7453,N_4908,N_5205);
xnor U7454 (N_7454,N_5826,N_5631);
nand U7455 (N_7455,N_4802,N_5325);
xor U7456 (N_7456,N_4508,N_5397);
or U7457 (N_7457,N_4874,N_5709);
nor U7458 (N_7458,N_5734,N_5871);
xor U7459 (N_7459,N_5670,N_4860);
xor U7460 (N_7460,N_5801,N_5182);
xor U7461 (N_7461,N_5844,N_5721);
xor U7462 (N_7462,N_5656,N_4786);
nand U7463 (N_7463,N_4743,N_5719);
nor U7464 (N_7464,N_5396,N_5377);
or U7465 (N_7465,N_5477,N_5416);
or U7466 (N_7466,N_5279,N_5520);
nand U7467 (N_7467,N_4656,N_5799);
nand U7468 (N_7468,N_5669,N_5466);
nor U7469 (N_7469,N_5480,N_4882);
nor U7470 (N_7470,N_4756,N_5375);
xnor U7471 (N_7471,N_5596,N_4908);
xor U7472 (N_7472,N_4580,N_5015);
or U7473 (N_7473,N_4632,N_4823);
or U7474 (N_7474,N_4611,N_5583);
xnor U7475 (N_7475,N_5348,N_5775);
and U7476 (N_7476,N_5663,N_5833);
xor U7477 (N_7477,N_4900,N_4513);
or U7478 (N_7478,N_4909,N_5729);
xor U7479 (N_7479,N_5820,N_5981);
nand U7480 (N_7480,N_4694,N_4667);
nor U7481 (N_7481,N_5905,N_4944);
xnor U7482 (N_7482,N_4815,N_5506);
or U7483 (N_7483,N_4595,N_4701);
or U7484 (N_7484,N_5972,N_5442);
or U7485 (N_7485,N_5252,N_5413);
or U7486 (N_7486,N_4749,N_5150);
nand U7487 (N_7487,N_5236,N_5485);
nor U7488 (N_7488,N_4587,N_5807);
nand U7489 (N_7489,N_4962,N_5967);
or U7490 (N_7490,N_5488,N_5747);
and U7491 (N_7491,N_5093,N_5847);
xor U7492 (N_7492,N_4641,N_4537);
nand U7493 (N_7493,N_4993,N_5218);
xnor U7494 (N_7494,N_5937,N_4877);
xor U7495 (N_7495,N_5642,N_4793);
nor U7496 (N_7496,N_5026,N_5315);
or U7497 (N_7497,N_5061,N_5849);
nand U7498 (N_7498,N_4857,N_5259);
xnor U7499 (N_7499,N_4960,N_5502);
and U7500 (N_7500,N_7075,N_6728);
or U7501 (N_7501,N_6814,N_6328);
or U7502 (N_7502,N_6110,N_6801);
xnor U7503 (N_7503,N_7151,N_7111);
nor U7504 (N_7504,N_6536,N_6909);
xor U7505 (N_7505,N_6989,N_7460);
nor U7506 (N_7506,N_6267,N_7192);
or U7507 (N_7507,N_6743,N_7396);
nor U7508 (N_7508,N_7057,N_6866);
nand U7509 (N_7509,N_6807,N_6407);
or U7510 (N_7510,N_7286,N_6394);
or U7511 (N_7511,N_7137,N_6222);
or U7512 (N_7512,N_6670,N_6746);
nand U7513 (N_7513,N_6220,N_7126);
or U7514 (N_7514,N_6249,N_6037);
nand U7515 (N_7515,N_6639,N_6293);
xor U7516 (N_7516,N_6868,N_6826);
nand U7517 (N_7517,N_7071,N_6829);
xor U7518 (N_7518,N_7241,N_7079);
and U7519 (N_7519,N_7437,N_6956);
xor U7520 (N_7520,N_7213,N_7227);
and U7521 (N_7521,N_6248,N_7301);
xor U7522 (N_7522,N_7013,N_6686);
and U7523 (N_7523,N_6008,N_6388);
nor U7524 (N_7524,N_6286,N_7074);
xnor U7525 (N_7525,N_6366,N_6982);
or U7526 (N_7526,N_6630,N_7365);
nor U7527 (N_7527,N_6664,N_6541);
xor U7528 (N_7528,N_7369,N_6972);
and U7529 (N_7529,N_6986,N_6393);
nor U7530 (N_7530,N_7338,N_7037);
nand U7531 (N_7531,N_6482,N_7256);
xnor U7532 (N_7532,N_6582,N_7116);
nor U7533 (N_7533,N_7159,N_6830);
nand U7534 (N_7534,N_7032,N_6887);
or U7535 (N_7535,N_6629,N_6688);
nor U7536 (N_7536,N_6895,N_7067);
nor U7537 (N_7537,N_6119,N_6931);
and U7538 (N_7538,N_6309,N_7012);
or U7539 (N_7539,N_7195,N_6631);
or U7540 (N_7540,N_6048,N_6080);
or U7541 (N_7541,N_6617,N_6127);
xor U7542 (N_7542,N_6530,N_6929);
or U7543 (N_7543,N_6789,N_6289);
and U7544 (N_7544,N_6244,N_6817);
or U7545 (N_7545,N_7284,N_6132);
nor U7546 (N_7546,N_7123,N_6567);
nand U7547 (N_7547,N_6905,N_6352);
nor U7548 (N_7548,N_6542,N_6257);
nor U7549 (N_7549,N_6644,N_6967);
nor U7550 (N_7550,N_7127,N_7435);
nor U7551 (N_7551,N_7366,N_7094);
nand U7552 (N_7552,N_7353,N_7428);
or U7553 (N_7553,N_7415,N_7334);
nor U7554 (N_7554,N_6498,N_6177);
or U7555 (N_7555,N_6233,N_7120);
or U7556 (N_7556,N_6809,N_6715);
nand U7557 (N_7557,N_7337,N_7021);
nand U7558 (N_7558,N_6418,N_6798);
and U7559 (N_7559,N_6044,N_7226);
and U7560 (N_7560,N_6572,N_7307);
and U7561 (N_7561,N_6808,N_6459);
xor U7562 (N_7562,N_7355,N_6841);
xor U7563 (N_7563,N_7097,N_7106);
xnor U7564 (N_7564,N_6063,N_7205);
nor U7565 (N_7565,N_6996,N_6270);
or U7566 (N_7566,N_6783,N_6315);
or U7567 (N_7567,N_6753,N_7038);
nand U7568 (N_7568,N_6495,N_6300);
nor U7569 (N_7569,N_6358,N_6474);
xor U7570 (N_7570,N_6872,N_6695);
nand U7571 (N_7571,N_6347,N_6974);
nand U7572 (N_7572,N_7211,N_6615);
nor U7573 (N_7573,N_7352,N_6687);
or U7574 (N_7574,N_7397,N_6272);
nand U7575 (N_7575,N_7309,N_6133);
xor U7576 (N_7576,N_6786,N_6993);
nor U7577 (N_7577,N_6638,N_7364);
or U7578 (N_7578,N_7129,N_6564);
or U7579 (N_7579,N_7197,N_7000);
xor U7580 (N_7580,N_6449,N_6741);
or U7581 (N_7581,N_6890,N_7341);
nor U7582 (N_7582,N_7168,N_7394);
and U7583 (N_7583,N_6441,N_6934);
and U7584 (N_7584,N_6634,N_6442);
and U7585 (N_7585,N_7380,N_6804);
and U7586 (N_7586,N_6384,N_6964);
nand U7587 (N_7587,N_7236,N_6475);
or U7588 (N_7588,N_7454,N_6174);
xor U7589 (N_7589,N_6955,N_6933);
nor U7590 (N_7590,N_6643,N_7183);
nand U7591 (N_7591,N_6236,N_7068);
nand U7592 (N_7592,N_6622,N_6027);
and U7593 (N_7593,N_6812,N_6253);
or U7594 (N_7594,N_6305,N_7306);
xor U7595 (N_7595,N_6528,N_6514);
xnor U7596 (N_7596,N_6576,N_7304);
or U7597 (N_7597,N_7020,N_6192);
xor U7598 (N_7598,N_6196,N_7008);
nor U7599 (N_7599,N_6769,N_6932);
nor U7600 (N_7600,N_7184,N_6780);
nor U7601 (N_7601,N_6504,N_6651);
xor U7602 (N_7602,N_7478,N_6563);
and U7603 (N_7603,N_6995,N_6428);
nand U7604 (N_7604,N_6167,N_6210);
xor U7605 (N_7605,N_7163,N_6454);
or U7606 (N_7606,N_6565,N_6460);
nand U7607 (N_7607,N_7387,N_6844);
nand U7608 (N_7608,N_7064,N_7351);
or U7609 (N_7609,N_6432,N_7017);
nor U7610 (N_7610,N_6524,N_6012);
and U7611 (N_7611,N_6710,N_6240);
nand U7612 (N_7612,N_6874,N_6461);
xnor U7613 (N_7613,N_7209,N_7110);
nor U7614 (N_7614,N_6487,N_6026);
xor U7615 (N_7615,N_7395,N_7208);
or U7616 (N_7616,N_6575,N_7407);
or U7617 (N_7617,N_6557,N_7392);
nor U7618 (N_7618,N_6232,N_6592);
nor U7619 (N_7619,N_7180,N_6509);
nand U7620 (N_7620,N_6345,N_6484);
and U7621 (N_7621,N_6537,N_6401);
nor U7622 (N_7622,N_6499,N_6785);
or U7623 (N_7623,N_7189,N_7264);
and U7624 (N_7624,N_7422,N_7065);
or U7625 (N_7625,N_6907,N_6560);
nand U7626 (N_7626,N_7354,N_6941);
nand U7627 (N_7627,N_7495,N_6251);
and U7628 (N_7628,N_6362,N_7050);
nor U7629 (N_7629,N_6417,N_6748);
and U7630 (N_7630,N_6526,N_6714);
nand U7631 (N_7631,N_6124,N_6730);
nand U7632 (N_7632,N_7091,N_6849);
or U7633 (N_7633,N_6578,N_6395);
or U7634 (N_7634,N_6344,N_6788);
or U7635 (N_7635,N_7174,N_6121);
and U7636 (N_7636,N_6260,N_6172);
or U7637 (N_7637,N_6488,N_6034);
and U7638 (N_7638,N_6370,N_6142);
or U7639 (N_7639,N_6811,N_7077);
and U7640 (N_7640,N_7031,N_6589);
xor U7641 (N_7641,N_7362,N_6773);
or U7642 (N_7642,N_7328,N_6489);
nor U7643 (N_7643,N_7316,N_6214);
nand U7644 (N_7644,N_6335,N_6953);
and U7645 (N_7645,N_7214,N_7260);
or U7646 (N_7646,N_6087,N_6337);
nor U7647 (N_7647,N_6698,N_6354);
xor U7648 (N_7648,N_6595,N_6213);
and U7649 (N_7649,N_6231,N_6060);
or U7650 (N_7650,N_7399,N_7072);
xor U7651 (N_7651,N_6556,N_7398);
xnor U7652 (N_7652,N_6111,N_7436);
xor U7653 (N_7653,N_7042,N_7432);
nor U7654 (N_7654,N_6009,N_6103);
nor U7655 (N_7655,N_6652,N_6648);
xnor U7656 (N_7656,N_7272,N_6099);
nor U7657 (N_7657,N_6481,N_7170);
xor U7658 (N_7658,N_6327,N_6666);
xnor U7659 (N_7659,N_7188,N_6294);
or U7660 (N_7660,N_6791,N_7300);
nand U7661 (N_7661,N_6371,N_7254);
xor U7662 (N_7662,N_7251,N_6752);
nor U7663 (N_7663,N_6476,N_6540);
or U7664 (N_7664,N_6448,N_6275);
nand U7665 (N_7665,N_6429,N_6502);
xor U7666 (N_7666,N_6511,N_6768);
nor U7667 (N_7667,N_6483,N_6042);
xor U7668 (N_7668,N_6451,N_7082);
and U7669 (N_7669,N_6732,N_7269);
xor U7670 (N_7670,N_7090,N_6054);
and U7671 (N_7671,N_7076,N_7470);
nor U7672 (N_7672,N_6723,N_6284);
or U7673 (N_7673,N_7348,N_7194);
xor U7674 (N_7674,N_6771,N_6558);
nor U7675 (N_7675,N_7294,N_6108);
nand U7676 (N_7676,N_6633,N_6843);
xnor U7677 (N_7677,N_6926,N_7314);
or U7678 (N_7678,N_6510,N_6884);
nor U7679 (N_7679,N_6452,N_6549);
or U7680 (N_7680,N_6479,N_6973);
xnor U7681 (N_7681,N_6170,N_6678);
nor U7682 (N_7682,N_7092,N_6225);
nor U7683 (N_7683,N_6927,N_6689);
nor U7684 (N_7684,N_6979,N_6424);
or U7685 (N_7685,N_7361,N_6923);
nor U7686 (N_7686,N_6910,N_7186);
xnor U7687 (N_7687,N_7245,N_6596);
nor U7688 (N_7688,N_6077,N_6377);
xor U7689 (N_7689,N_6107,N_7469);
xor U7690 (N_7690,N_6276,N_7280);
xnor U7691 (N_7691,N_6295,N_6935);
nor U7692 (N_7692,N_7004,N_6913);
and U7693 (N_7693,N_6543,N_6659);
nand U7694 (N_7694,N_6013,N_6039);
nand U7695 (N_7695,N_6637,N_6067);
or U7696 (N_7696,N_7144,N_6040);
and U7697 (N_7697,N_6090,N_7305);
and U7698 (N_7698,N_6379,N_6889);
xnor U7699 (N_7699,N_6463,N_7278);
and U7700 (N_7700,N_7438,N_6224);
or U7701 (N_7701,N_6400,N_6096);
or U7702 (N_7702,N_7234,N_6234);
xnor U7703 (N_7703,N_6691,N_7374);
and U7704 (N_7704,N_7499,N_6856);
or U7705 (N_7705,N_7340,N_6190);
xor U7706 (N_7706,N_7142,N_6126);
nor U7707 (N_7707,N_6477,N_6776);
nand U7708 (N_7708,N_6614,N_7325);
and U7709 (N_7709,N_6883,N_6824);
nor U7710 (N_7710,N_7448,N_7164);
nor U7711 (N_7711,N_6282,N_6645);
xor U7712 (N_7712,N_6778,N_7046);
nand U7713 (N_7713,N_7219,N_6002);
xnor U7714 (N_7714,N_6153,N_6113);
or U7715 (N_7715,N_6863,N_6492);
and U7716 (N_7716,N_6412,N_6810);
or U7717 (N_7717,N_6625,N_7084);
or U7718 (N_7718,N_6444,N_6727);
nand U7719 (N_7719,N_6827,N_7081);
and U7720 (N_7720,N_6363,N_6552);
or U7721 (N_7721,N_7440,N_7452);
xnor U7722 (N_7722,N_7393,N_6070);
nand U7723 (N_7723,N_6960,N_6600);
nand U7724 (N_7724,N_6815,N_7015);
nor U7725 (N_7725,N_6946,N_6033);
or U7726 (N_7726,N_6820,N_6961);
and U7727 (N_7727,N_7283,N_6204);
and U7728 (N_7728,N_7185,N_7177);
xnor U7729 (N_7729,N_6548,N_6274);
nor U7730 (N_7730,N_6030,N_6200);
nand U7731 (N_7731,N_6922,N_6770);
xnor U7732 (N_7732,N_7434,N_6082);
nor U7733 (N_7733,N_6246,N_6566);
xnor U7734 (N_7734,N_7212,N_7140);
or U7735 (N_7735,N_6209,N_7431);
nor U7736 (N_7736,N_6215,N_6531);
nor U7737 (N_7737,N_6265,N_6297);
xnor U7738 (N_7738,N_6292,N_7492);
nand U7739 (N_7739,N_6952,N_6500);
or U7740 (N_7740,N_7016,N_6440);
or U7741 (N_7741,N_6908,N_7166);
nor U7742 (N_7742,N_7490,N_6365);
nor U7743 (N_7743,N_6683,N_6212);
nor U7744 (N_7744,N_6386,N_7235);
nand U7745 (N_7745,N_6649,N_6657);
xnor U7746 (N_7746,N_6697,N_6045);
and U7747 (N_7747,N_6912,N_6740);
nor U7748 (N_7748,N_6273,N_7292);
and U7749 (N_7749,N_6836,N_6221);
nor U7750 (N_7750,N_6001,N_7257);
or U7751 (N_7751,N_7322,N_7481);
or U7752 (N_7752,N_7330,N_6319);
xor U7753 (N_7753,N_6436,N_6069);
xnor U7754 (N_7754,N_6782,N_7001);
xor U7755 (N_7755,N_7423,N_7139);
or U7756 (N_7756,N_7376,N_6568);
xor U7757 (N_7757,N_7253,N_7014);
nor U7758 (N_7758,N_6168,N_6779);
nor U7759 (N_7759,N_6672,N_6437);
xor U7760 (N_7760,N_6825,N_6750);
or U7761 (N_7761,N_7148,N_6179);
nor U7762 (N_7762,N_6587,N_6194);
nand U7763 (N_7763,N_6230,N_6456);
and U7764 (N_7764,N_6854,N_6144);
xor U7765 (N_7765,N_6619,N_7429);
and U7766 (N_7766,N_6405,N_6369);
nand U7767 (N_7767,N_7217,N_6373);
nand U7768 (N_7768,N_7147,N_6466);
nor U7769 (N_7769,N_6120,N_6439);
xor U7770 (N_7770,N_6660,N_6490);
nor U7771 (N_7771,N_7141,N_6711);
or U7772 (N_7772,N_7472,N_6227);
and U7773 (N_7773,N_6496,N_6161);
or U7774 (N_7774,N_6238,N_6047);
and U7775 (N_7775,N_6114,N_6925);
xor U7776 (N_7776,N_7218,N_7178);
nand U7777 (N_7777,N_6301,N_7413);
xnor U7778 (N_7778,N_7373,N_6602);
xor U7779 (N_7779,N_6937,N_6198);
and U7780 (N_7780,N_6302,N_6865);
nor U7781 (N_7781,N_6304,N_6963);
xnor U7782 (N_7782,N_7426,N_6020);
or U7783 (N_7783,N_6719,N_7158);
and U7784 (N_7784,N_7237,N_6951);
xor U7785 (N_7785,N_6433,N_7089);
xnor U7786 (N_7786,N_6739,N_7061);
or U7787 (N_7787,N_7344,N_7403);
xor U7788 (N_7788,N_7165,N_6516);
xnor U7789 (N_7789,N_6356,N_7281);
nand U7790 (N_7790,N_6193,N_7143);
nand U7791 (N_7791,N_6677,N_6331);
and U7792 (N_7792,N_7206,N_7480);
nor U7793 (N_7793,N_6413,N_6004);
nand U7794 (N_7794,N_6754,N_6202);
and U7795 (N_7795,N_7221,N_7367);
xnor U7796 (N_7796,N_7005,N_6035);
and U7797 (N_7797,N_6733,N_7486);
xor U7798 (N_7798,N_7441,N_7498);
nand U7799 (N_7799,N_7243,N_6247);
or U7800 (N_7800,N_6116,N_6936);
or U7801 (N_7801,N_7418,N_6885);
nor U7802 (N_7802,N_6078,N_6287);
nand U7803 (N_7803,N_6191,N_6692);
and U7804 (N_7804,N_6501,N_6823);
nor U7805 (N_7805,N_7493,N_7390);
and U7806 (N_7806,N_6641,N_6197);
and U7807 (N_7807,N_7066,N_6410);
and U7808 (N_7808,N_6627,N_6969);
or U7809 (N_7809,N_6999,N_6416);
nand U7810 (N_7810,N_7485,N_7190);
or U7811 (N_7811,N_6349,N_7224);
nand U7812 (N_7812,N_7095,N_7167);
nor U7813 (N_7813,N_7331,N_6053);
or U7814 (N_7814,N_7282,N_6137);
nand U7815 (N_7815,N_7115,N_7475);
nand U7816 (N_7816,N_6073,N_7179);
and U7817 (N_7817,N_6316,N_6091);
and U7818 (N_7818,N_6446,N_6832);
or U7819 (N_7819,N_7252,N_6920);
xnor U7820 (N_7820,N_7202,N_6291);
or U7821 (N_7821,N_6860,N_7319);
xnor U7822 (N_7822,N_6724,N_7276);
or U7823 (N_7823,N_6406,N_6350);
and U7824 (N_7824,N_6171,N_7047);
and U7825 (N_7825,N_7220,N_6317);
nand U7826 (N_7826,N_6296,N_6851);
xor U7827 (N_7827,N_7425,N_6195);
xor U7828 (N_7828,N_6819,N_6138);
and U7829 (N_7829,N_6129,N_7128);
nand U7830 (N_7830,N_6376,N_6593);
xnor U7831 (N_7831,N_6793,N_6403);
and U7832 (N_7832,N_7198,N_7259);
nor U7833 (N_7833,N_6330,N_6426);
and U7834 (N_7834,N_7274,N_7250);
and U7835 (N_7835,N_6324,N_6010);
xor U7836 (N_7836,N_7442,N_6464);
nand U7837 (N_7837,N_7263,N_7052);
nand U7838 (N_7838,N_6076,N_7455);
and U7839 (N_7839,N_6764,N_6065);
and U7840 (N_7840,N_6945,N_6997);
nor U7841 (N_7841,N_6792,N_7446);
xor U7842 (N_7842,N_6603,N_6427);
nand U7843 (N_7843,N_7023,N_6465);
xnor U7844 (N_7844,N_6707,N_6368);
nor U7845 (N_7845,N_7130,N_7381);
and U7846 (N_7846,N_6671,N_7296);
nand U7847 (N_7847,N_7468,N_7039);
or U7848 (N_7848,N_7402,N_7310);
xor U7849 (N_7849,N_7285,N_6383);
or U7850 (N_7850,N_6553,N_6447);
and U7851 (N_7851,N_7119,N_6506);
and U7852 (N_7852,N_6601,N_6544);
xor U7853 (N_7853,N_7203,N_6336);
nor U7854 (N_7854,N_7103,N_6462);
nor U7855 (N_7855,N_6681,N_6152);
nor U7856 (N_7856,N_7462,N_7086);
and U7857 (N_7857,N_6199,N_6699);
xnor U7858 (N_7858,N_7006,N_7474);
nor U7859 (N_7859,N_6871,N_6155);
and U7860 (N_7860,N_6712,N_6458);
xor U7861 (N_7861,N_6799,N_6092);
and U7862 (N_7862,N_6438,N_6980);
and U7863 (N_7863,N_6828,N_7336);
nor U7864 (N_7864,N_6201,N_6586);
xnor U7865 (N_7865,N_6661,N_6805);
or U7866 (N_7866,N_6313,N_6642);
nand U7867 (N_7867,N_6322,N_6188);
and U7868 (N_7868,N_7420,N_6095);
and U7869 (N_7869,N_6673,N_7419);
nor U7870 (N_7870,N_6283,N_6181);
and U7871 (N_7871,N_6850,N_6262);
nand U7872 (N_7872,N_6962,N_7410);
or U7873 (N_7873,N_6977,N_7029);
or U7874 (N_7874,N_6338,N_6408);
nor U7875 (N_7875,N_7450,N_6068);
and U7876 (N_7876,N_7121,N_7010);
nand U7877 (N_7877,N_6308,N_7223);
nor U7878 (N_7878,N_6399,N_6736);
or U7879 (N_7879,N_6512,N_6585);
xnor U7880 (N_7880,N_6051,N_7242);
nor U7881 (N_7881,N_6223,N_6071);
or U7882 (N_7882,N_7247,N_6834);
or U7883 (N_7883,N_6583,N_6421);
and U7884 (N_7884,N_6981,N_6674);
xnor U7885 (N_7885,N_7187,N_6881);
and U7886 (N_7886,N_7409,N_6747);
nand U7887 (N_7887,N_6990,N_6612);
nand U7888 (N_7888,N_6940,N_6392);
nand U7889 (N_7889,N_7293,N_6485);
xnor U7890 (N_7890,N_6915,N_6760);
or U7891 (N_7891,N_7494,N_7345);
nor U7892 (N_7892,N_7406,N_6790);
nand U7893 (N_7893,N_6577,N_6546);
nor U7894 (N_7894,N_6545,N_6140);
and U7895 (N_7895,N_6320,N_7125);
and U7896 (N_7896,N_6325,N_6493);
xnor U7897 (N_7897,N_6831,N_6391);
xnor U7898 (N_7898,N_6520,N_6017);
and U7899 (N_7899,N_6756,N_7045);
xnor U7900 (N_7900,N_6983,N_7389);
nand U7901 (N_7901,N_6314,N_6668);
nand U7902 (N_7902,N_7232,N_7018);
xnor U7903 (N_7903,N_6696,N_6876);
nor U7904 (N_7904,N_7449,N_6998);
xnor U7905 (N_7905,N_6165,N_7138);
xnor U7906 (N_7906,N_6375,N_6984);
or U7907 (N_7907,N_7153,N_7162);
or U7908 (N_7908,N_7225,N_6084);
nor U7909 (N_7909,N_7484,N_6254);
nand U7910 (N_7910,N_7258,N_6064);
xnor U7911 (N_7911,N_7482,N_7473);
and U7912 (N_7912,N_6944,N_6729);
or U7913 (N_7913,N_6947,N_7122);
xor U7914 (N_7914,N_6036,N_6404);
nand U7915 (N_7915,N_7303,N_6343);
or U7916 (N_7916,N_7324,N_6279);
xor U7917 (N_7917,N_6749,N_6611);
nor U7918 (N_7918,N_7349,N_7182);
nor U7919 (N_7919,N_6667,N_6978);
nand U7920 (N_7920,N_6074,N_7249);
and U7921 (N_7921,N_7034,N_6654);
and U7922 (N_7922,N_6310,N_7479);
xor U7923 (N_7923,N_6241,N_6538);
or U7924 (N_7924,N_6902,N_6156);
and U7925 (N_7925,N_6333,N_7372);
and U7926 (N_7926,N_6128,N_7458);
xor U7927 (N_7927,N_6919,N_6505);
or U7928 (N_7928,N_6787,N_6848);
and U7929 (N_7929,N_6985,N_7375);
xor U7930 (N_7930,N_7176,N_6473);
nor U7931 (N_7931,N_6435,N_6579);
and U7932 (N_7932,N_6148,N_6235);
nor U7933 (N_7933,N_6650,N_6574);
or U7934 (N_7934,N_6402,N_6258);
and U7935 (N_7935,N_6396,N_7114);
xor U7936 (N_7936,N_6271,N_6662);
or U7937 (N_7937,N_7048,N_6701);
or U7938 (N_7938,N_7215,N_7161);
and U7939 (N_7939,N_6838,N_7199);
nor U7940 (N_7940,N_6894,N_6864);
or U7941 (N_7941,N_6180,N_6610);
or U7942 (N_7942,N_6775,N_6043);
xor U7943 (N_7943,N_7430,N_7069);
and U7944 (N_7944,N_7457,N_6718);
and U7945 (N_7945,N_7191,N_6380);
nand U7946 (N_7946,N_7404,N_7022);
and U7947 (N_7947,N_6207,N_6855);
nor U7948 (N_7948,N_6870,N_6527);
nand U7949 (N_7949,N_7433,N_6857);
xnor U7950 (N_7950,N_6298,N_6759);
xnor U7951 (N_7951,N_6581,N_6183);
or U7952 (N_7952,N_6093,N_6959);
nor U7953 (N_7953,N_6229,N_6057);
or U7954 (N_7954,N_6519,N_7327);
xnor U7955 (N_7955,N_6332,N_6562);
xnor U7956 (N_7956,N_6050,N_6626);
nor U7957 (N_7957,N_6525,N_6079);
nand U7958 (N_7958,N_6003,N_7173);
nand U7959 (N_7959,N_6529,N_6766);
or U7960 (N_7960,N_6976,N_6216);
and U7961 (N_7961,N_6311,N_7024);
nor U7962 (N_7962,N_7136,N_6862);
nor U7963 (N_7963,N_6162,N_6359);
nand U7964 (N_7964,N_7007,N_7059);
nor U7965 (N_7965,N_6916,N_6299);
nand U7966 (N_7966,N_7093,N_6886);
and U7967 (N_7967,N_6425,N_7465);
nand U7968 (N_7968,N_6914,N_6802);
and U7969 (N_7969,N_7488,N_6751);
nor U7970 (N_7970,N_6663,N_6007);
nand U7971 (N_7971,N_6106,N_7401);
nand U7972 (N_7972,N_6117,N_7342);
and U7973 (N_7973,N_6803,N_7357);
and U7974 (N_7974,N_6713,N_6361);
nor U7975 (N_7975,N_6554,N_6182);
and U7976 (N_7976,N_6089,N_6503);
or U7977 (N_7977,N_6987,N_6762);
and U7978 (N_7978,N_7335,N_7181);
nor U7979 (N_7979,N_7002,N_6085);
nor U7980 (N_7980,N_6797,N_7255);
xor U7981 (N_7981,N_7339,N_6381);
nor U7982 (N_7982,N_7368,N_6259);
xor U7983 (N_7983,N_7098,N_6154);
nand U7984 (N_7984,N_7329,N_6684);
xor U7985 (N_7985,N_7201,N_6898);
xor U7986 (N_7986,N_7363,N_7222);
xnor U7987 (N_7987,N_7356,N_6430);
nand U7988 (N_7988,N_7231,N_6737);
or U7989 (N_7989,N_6075,N_6340);
and U7990 (N_7990,N_6621,N_6176);
or U7991 (N_7991,N_6123,N_6280);
nand U7992 (N_7992,N_7088,N_6640);
xnor U7993 (N_7993,N_6900,N_7421);
nor U7994 (N_7994,N_7467,N_6378);
xnor U7995 (N_7995,N_7053,N_6613);
xnor U7996 (N_7996,N_6968,N_7003);
or U7997 (N_7997,N_7302,N_6139);
xnor U7998 (N_7998,N_6725,N_6431);
or U7999 (N_7999,N_6219,N_6571);
nor U8000 (N_8000,N_6346,N_6341);
nor U8001 (N_8001,N_6173,N_7132);
and U8002 (N_8002,N_6590,N_7295);
nand U8003 (N_8003,N_6469,N_7371);
and U8004 (N_8004,N_7385,N_6024);
or U8005 (N_8005,N_6029,N_6398);
nor U8006 (N_8006,N_6118,N_7246);
or U8007 (N_8007,N_6561,N_6774);
nor U8008 (N_8008,N_6594,N_7175);
and U8009 (N_8009,N_6608,N_6164);
nor U8010 (N_8010,N_6605,N_6917);
nand U8011 (N_8011,N_6334,N_6877);
or U8012 (N_8012,N_7019,N_7291);
nor U8013 (N_8013,N_6970,N_7150);
nor U8014 (N_8014,N_6058,N_6387);
or U8015 (N_8015,N_7056,N_6796);
or U8016 (N_8016,N_7312,N_6821);
nand U8017 (N_8017,N_7124,N_6609);
and U8018 (N_8018,N_6653,N_6245);
nor U8019 (N_8019,N_6450,N_6205);
and U8020 (N_8020,N_7287,N_6414);
nor U8021 (N_8021,N_7377,N_6584);
nor U8022 (N_8022,N_6896,N_7228);
and U8023 (N_8023,N_6888,N_7491);
and U8024 (N_8024,N_6357,N_6604);
nand U8025 (N_8025,N_6088,N_6125);
or U8026 (N_8026,N_6928,N_6318);
nand U8027 (N_8027,N_6906,N_6535);
or U8028 (N_8028,N_7155,N_6022);
and U8029 (N_8029,N_6021,N_6597);
xnor U8030 (N_8030,N_6146,N_7487);
nand U8031 (N_8031,N_6385,N_6606);
nand U8032 (N_8032,N_6893,N_7078);
and U8033 (N_8033,N_7101,N_6072);
and U8034 (N_8034,N_6846,N_6742);
xor U8035 (N_8035,N_6323,N_6443);
and U8036 (N_8036,N_6559,N_6901);
and U8037 (N_8037,N_7320,N_6491);
nor U8038 (N_8038,N_6744,N_6497);
or U8039 (N_8039,N_6321,N_6372);
or U8040 (N_8040,N_6288,N_6134);
nor U8041 (N_8041,N_7346,N_6708);
nand U8042 (N_8042,N_6160,N_6765);
nand U8043 (N_8043,N_7035,N_6409);
or U8044 (N_8044,N_6023,N_6624);
nand U8045 (N_8045,N_7109,N_7080);
or U8046 (N_8046,N_6208,N_6264);
nor U8047 (N_8047,N_7229,N_6533);
xor U8048 (N_8048,N_6816,N_6252);
or U8049 (N_8049,N_6694,N_7131);
or U8050 (N_8050,N_7378,N_7134);
xor U8051 (N_8051,N_7049,N_6186);
nor U8052 (N_8052,N_7152,N_6389);
nand U8053 (N_8053,N_7273,N_6445);
nand U8054 (N_8054,N_7233,N_7308);
or U8055 (N_8055,N_6704,N_6680);
nor U8056 (N_8056,N_7200,N_6364);
or U8057 (N_8057,N_7154,N_6616);
or U8058 (N_8058,N_6591,N_7062);
nor U8059 (N_8059,N_6822,N_7149);
or U8060 (N_8060,N_6243,N_6097);
nand U8061 (N_8061,N_7060,N_7087);
and U8062 (N_8062,N_7315,N_6942);
nand U8063 (N_8063,N_6847,N_6066);
nor U8064 (N_8064,N_6569,N_6513);
xnor U8065 (N_8065,N_6623,N_6158);
and U8066 (N_8066,N_6706,N_7009);
xor U8067 (N_8067,N_6101,N_6360);
xor U8068 (N_8068,N_6632,N_7145);
xor U8069 (N_8069,N_6374,N_7444);
xor U8070 (N_8070,N_6859,N_7461);
nand U8071 (N_8071,N_7464,N_6948);
nand U8072 (N_8072,N_6115,N_7041);
nand U8073 (N_8073,N_6348,N_7360);
or U8074 (N_8074,N_6669,N_7196);
and U8075 (N_8075,N_6522,N_6015);
nand U8076 (N_8076,N_6539,N_7207);
xnor U8077 (N_8077,N_6206,N_7051);
nand U8078 (N_8078,N_6873,N_7096);
or U8079 (N_8079,N_6130,N_6277);
nand U8080 (N_8080,N_7026,N_6382);
xnor U8081 (N_8081,N_6758,N_6339);
xor U8082 (N_8082,N_6635,N_6028);
nor U8083 (N_8083,N_6467,N_7146);
nand U8084 (N_8084,N_6794,N_6813);
or U8085 (N_8085,N_6795,N_7299);
xnor U8086 (N_8086,N_7238,N_6656);
nor U8087 (N_8087,N_6281,N_6880);
or U8088 (N_8088,N_7288,N_6628);
xnor U8089 (N_8089,N_6508,N_6722);
nand U8090 (N_8090,N_6143,N_6109);
or U8091 (N_8091,N_7424,N_6833);
nor U8092 (N_8092,N_7117,N_6237);
or U8093 (N_8093,N_7210,N_6897);
xor U8094 (N_8094,N_6218,N_6307);
and U8095 (N_8095,N_6837,N_7477);
nand U8096 (N_8096,N_7427,N_6175);
and U8097 (N_8097,N_6965,N_6434);
xnor U8098 (N_8098,N_6005,N_6420);
or U8099 (N_8099,N_7405,N_7416);
nor U8100 (N_8100,N_6647,N_7489);
nand U8101 (N_8101,N_6938,N_6189);
xor U8102 (N_8102,N_6761,N_6781);
and U8103 (N_8103,N_7445,N_7100);
or U8104 (N_8104,N_6852,N_6468);
nand U8105 (N_8105,N_6700,N_6151);
nor U8106 (N_8106,N_7326,N_6892);
or U8107 (N_8107,N_6717,N_6924);
xnor U8108 (N_8108,N_7113,N_6971);
and U8109 (N_8109,N_7275,N_6975);
or U8110 (N_8110,N_6757,N_6157);
or U8111 (N_8111,N_6453,N_6818);
or U8112 (N_8112,N_6062,N_7157);
nor U8113 (N_8113,N_6263,N_6867);
and U8114 (N_8114,N_7343,N_7311);
nor U8115 (N_8115,N_6507,N_6994);
xnor U8116 (N_8116,N_6472,N_6958);
xnor U8117 (N_8117,N_6679,N_7483);
nor U8118 (N_8118,N_6882,N_6784);
nor U8119 (N_8119,N_6570,N_6957);
nand U8120 (N_8120,N_6184,N_7193);
nand U8121 (N_8121,N_7054,N_6256);
nor U8122 (N_8122,N_6869,N_6242);
and U8123 (N_8123,N_7104,N_7266);
xnor U8124 (N_8124,N_6891,N_6000);
nor U8125 (N_8125,N_7073,N_6228);
xnor U8126 (N_8126,N_7359,N_6105);
nand U8127 (N_8127,N_6163,N_6858);
nand U8128 (N_8128,N_6226,N_7412);
xnor U8129 (N_8129,N_7105,N_6853);
and U8130 (N_8130,N_6355,N_6515);
xnor U8131 (N_8131,N_6342,N_7028);
nand U8132 (N_8132,N_6580,N_6772);
xor U8133 (N_8133,N_6457,N_6032);
xor U8134 (N_8134,N_6018,N_6122);
or U8135 (N_8135,N_7417,N_6187);
xnor U8136 (N_8136,N_7414,N_7411);
or U8137 (N_8137,N_6285,N_6949);
or U8138 (N_8138,N_6845,N_6731);
and U8139 (N_8139,N_6081,N_7102);
nand U8140 (N_8140,N_7070,N_6094);
xor U8141 (N_8141,N_6551,N_6150);
nor U8142 (N_8142,N_7297,N_6930);
xor U8143 (N_8143,N_7451,N_6312);
xnor U8144 (N_8144,N_6056,N_6636);
xnor U8145 (N_8145,N_7271,N_6041);
and U8146 (N_8146,N_6534,N_6665);
nor U8147 (N_8147,N_6861,N_6423);
and U8148 (N_8148,N_7230,N_6598);
nor U8149 (N_8149,N_6059,N_7108);
nor U8150 (N_8150,N_7244,N_6278);
nor U8151 (N_8151,N_6086,N_7443);
nor U8152 (N_8152,N_7112,N_7408);
nand U8153 (N_8153,N_6250,N_7044);
nand U8154 (N_8154,N_6353,N_6755);
or U8155 (N_8155,N_7133,N_6777);
nor U8156 (N_8156,N_6166,N_6486);
and U8157 (N_8157,N_7248,N_6763);
and U8158 (N_8158,N_6390,N_7321);
nor U8159 (N_8159,N_6618,N_6266);
and U8160 (N_8160,N_6367,N_6878);
and U8161 (N_8161,N_6839,N_6693);
nand U8162 (N_8162,N_6083,N_6217);
or U8163 (N_8163,N_6903,N_6518);
or U8164 (N_8164,N_6709,N_6326);
nor U8165 (N_8165,N_6911,N_6658);
nand U8166 (N_8166,N_6255,N_7063);
xnor U8167 (N_8167,N_6992,N_6203);
nand U8168 (N_8168,N_6685,N_7313);
nand U8169 (N_8169,N_6178,N_7466);
nand U8170 (N_8170,N_6767,N_7171);
xnor U8171 (N_8171,N_7135,N_6676);
nor U8172 (N_8172,N_6329,N_6555);
nor U8173 (N_8173,N_6290,N_6550);
nand U8174 (N_8174,N_7370,N_6720);
nor U8175 (N_8175,N_6478,N_6840);
nand U8176 (N_8176,N_7379,N_6261);
nand U8177 (N_8177,N_6716,N_6875);
xor U8178 (N_8178,N_6031,N_7382);
or U8179 (N_8179,N_7239,N_7204);
and U8180 (N_8180,N_7456,N_7099);
and U8181 (N_8181,N_6480,N_6547);
and U8182 (N_8182,N_6159,N_6703);
nand U8183 (N_8183,N_6055,N_6011);
nand U8184 (N_8184,N_6100,N_7083);
nor U8185 (N_8185,N_6061,N_6899);
nor U8186 (N_8186,N_7160,N_6702);
nand U8187 (N_8187,N_7497,N_7459);
nor U8188 (N_8188,N_7172,N_7240);
xor U8189 (N_8189,N_6470,N_6800);
nand U8190 (N_8190,N_7496,N_6046);
and U8191 (N_8191,N_7447,N_6991);
and U8192 (N_8192,N_6131,N_6006);
or U8193 (N_8193,N_7156,N_6415);
nand U8194 (N_8194,N_7358,N_6455);
xnor U8195 (N_8195,N_7298,N_7400);
nor U8196 (N_8196,N_6735,N_7332);
and U8197 (N_8197,N_6351,N_7033);
nor U8198 (N_8198,N_6607,N_7277);
nand U8199 (N_8199,N_7388,N_7268);
or U8200 (N_8200,N_6842,N_6141);
nand U8201 (N_8201,N_7476,N_6726);
nand U8202 (N_8202,N_7216,N_6014);
or U8203 (N_8203,N_6966,N_7265);
nor U8204 (N_8204,N_7391,N_7036);
nand U8205 (N_8205,N_6835,N_6494);
and U8206 (N_8206,N_7463,N_6690);
xnor U8207 (N_8207,N_6169,N_7317);
xnor U8208 (N_8208,N_6921,N_7011);
xor U8209 (N_8209,N_7386,N_7289);
xor U8210 (N_8210,N_7169,N_6532);
xor U8211 (N_8211,N_6419,N_6620);
nand U8212 (N_8212,N_6268,N_6019);
nand U8213 (N_8213,N_6145,N_7267);
xnor U8214 (N_8214,N_6422,N_7040);
and U8215 (N_8215,N_6806,N_7453);
and U8216 (N_8216,N_6038,N_6904);
and U8217 (N_8217,N_6239,N_6136);
or U8218 (N_8218,N_7262,N_6269);
nor U8219 (N_8219,N_6397,N_7279);
nor U8220 (N_8220,N_6025,N_6016);
nand U8221 (N_8221,N_7107,N_6306);
nand U8222 (N_8222,N_6988,N_6599);
xnor U8223 (N_8223,N_6745,N_6646);
nand U8224 (N_8224,N_6211,N_6918);
or U8225 (N_8225,N_6104,N_6517);
xor U8226 (N_8226,N_7350,N_7347);
nor U8227 (N_8227,N_7471,N_6738);
xor U8228 (N_8228,N_6879,N_6149);
nor U8229 (N_8229,N_6185,N_6471);
xnor U8230 (N_8230,N_6112,N_6954);
or U8231 (N_8231,N_6523,N_6655);
or U8232 (N_8232,N_7058,N_7383);
or U8233 (N_8233,N_6675,N_6098);
or U8234 (N_8234,N_7118,N_7439);
nor U8235 (N_8235,N_6705,N_6049);
or U8236 (N_8236,N_6588,N_7055);
nand U8237 (N_8237,N_6521,N_7318);
nand U8238 (N_8238,N_6135,N_7384);
or U8239 (N_8239,N_7025,N_7323);
nor U8240 (N_8240,N_6943,N_6734);
or U8241 (N_8241,N_7333,N_7027);
nand U8242 (N_8242,N_6411,N_6573);
or U8243 (N_8243,N_6147,N_6950);
nand U8244 (N_8244,N_6939,N_7030);
and U8245 (N_8245,N_6682,N_6052);
nand U8246 (N_8246,N_6721,N_7261);
or U8247 (N_8247,N_7085,N_7290);
xor U8248 (N_8248,N_6102,N_6303);
nor U8249 (N_8249,N_7043,N_7270);
xor U8250 (N_8250,N_6593,N_6142);
and U8251 (N_8251,N_6300,N_6023);
xnor U8252 (N_8252,N_7449,N_6113);
xnor U8253 (N_8253,N_7356,N_6788);
or U8254 (N_8254,N_6601,N_6033);
xnor U8255 (N_8255,N_6213,N_6389);
nor U8256 (N_8256,N_6455,N_7297);
or U8257 (N_8257,N_7120,N_7205);
or U8258 (N_8258,N_6989,N_6509);
nor U8259 (N_8259,N_7110,N_6041);
or U8260 (N_8260,N_7494,N_6778);
or U8261 (N_8261,N_6866,N_6182);
nand U8262 (N_8262,N_6136,N_6578);
nor U8263 (N_8263,N_7322,N_6975);
nand U8264 (N_8264,N_6218,N_7320);
nand U8265 (N_8265,N_7233,N_7073);
and U8266 (N_8266,N_6786,N_6963);
or U8267 (N_8267,N_7175,N_7182);
xnor U8268 (N_8268,N_7209,N_6791);
nand U8269 (N_8269,N_6032,N_7006);
or U8270 (N_8270,N_7453,N_7014);
nor U8271 (N_8271,N_6061,N_7441);
and U8272 (N_8272,N_6134,N_6799);
or U8273 (N_8273,N_6825,N_6139);
xor U8274 (N_8274,N_6790,N_6055);
nand U8275 (N_8275,N_6785,N_7432);
xnor U8276 (N_8276,N_6681,N_6441);
nor U8277 (N_8277,N_6547,N_7143);
and U8278 (N_8278,N_6698,N_6321);
xnor U8279 (N_8279,N_6531,N_6055);
xnor U8280 (N_8280,N_7107,N_6782);
xnor U8281 (N_8281,N_6446,N_6295);
nand U8282 (N_8282,N_6824,N_6980);
or U8283 (N_8283,N_6806,N_7096);
or U8284 (N_8284,N_6053,N_7091);
and U8285 (N_8285,N_7455,N_6400);
nor U8286 (N_8286,N_7276,N_6649);
or U8287 (N_8287,N_6159,N_7459);
xnor U8288 (N_8288,N_6458,N_7368);
nand U8289 (N_8289,N_6982,N_6909);
nand U8290 (N_8290,N_7327,N_6720);
or U8291 (N_8291,N_6935,N_6289);
and U8292 (N_8292,N_6659,N_6553);
nand U8293 (N_8293,N_6914,N_6525);
nor U8294 (N_8294,N_6531,N_6394);
xnor U8295 (N_8295,N_6524,N_7017);
or U8296 (N_8296,N_7367,N_6361);
nand U8297 (N_8297,N_6271,N_6365);
and U8298 (N_8298,N_6784,N_7289);
or U8299 (N_8299,N_6156,N_6660);
and U8300 (N_8300,N_6599,N_6880);
or U8301 (N_8301,N_6802,N_7173);
nand U8302 (N_8302,N_7127,N_7104);
or U8303 (N_8303,N_6561,N_6730);
and U8304 (N_8304,N_7211,N_6212);
nor U8305 (N_8305,N_6208,N_6835);
xnor U8306 (N_8306,N_7029,N_6621);
or U8307 (N_8307,N_6380,N_6836);
xor U8308 (N_8308,N_6891,N_7155);
and U8309 (N_8309,N_7073,N_6333);
nor U8310 (N_8310,N_6943,N_6193);
or U8311 (N_8311,N_6172,N_6203);
nand U8312 (N_8312,N_6820,N_6572);
or U8313 (N_8313,N_7051,N_6158);
and U8314 (N_8314,N_6741,N_6331);
nand U8315 (N_8315,N_7244,N_7406);
and U8316 (N_8316,N_6603,N_7355);
xor U8317 (N_8317,N_6199,N_7476);
nor U8318 (N_8318,N_6689,N_6425);
or U8319 (N_8319,N_6258,N_6465);
or U8320 (N_8320,N_6716,N_6894);
nor U8321 (N_8321,N_7157,N_6032);
nand U8322 (N_8322,N_6078,N_6436);
nor U8323 (N_8323,N_6411,N_7141);
or U8324 (N_8324,N_6207,N_6249);
and U8325 (N_8325,N_6881,N_6531);
and U8326 (N_8326,N_7349,N_6616);
nor U8327 (N_8327,N_7217,N_6887);
nand U8328 (N_8328,N_6710,N_6842);
or U8329 (N_8329,N_6820,N_7492);
xnor U8330 (N_8330,N_6820,N_6273);
xnor U8331 (N_8331,N_6447,N_7211);
nor U8332 (N_8332,N_6126,N_6535);
nor U8333 (N_8333,N_7320,N_6579);
and U8334 (N_8334,N_6592,N_6058);
nand U8335 (N_8335,N_7459,N_6229);
nor U8336 (N_8336,N_6168,N_7256);
or U8337 (N_8337,N_6068,N_7438);
nand U8338 (N_8338,N_7151,N_6732);
nor U8339 (N_8339,N_6875,N_6838);
nand U8340 (N_8340,N_7058,N_6898);
nor U8341 (N_8341,N_6892,N_6251);
xor U8342 (N_8342,N_6669,N_6143);
xnor U8343 (N_8343,N_7025,N_6265);
and U8344 (N_8344,N_6190,N_7042);
xor U8345 (N_8345,N_6665,N_6381);
nor U8346 (N_8346,N_6241,N_6170);
or U8347 (N_8347,N_6228,N_6437);
and U8348 (N_8348,N_6186,N_6039);
and U8349 (N_8349,N_6404,N_6905);
xor U8350 (N_8350,N_6289,N_6938);
or U8351 (N_8351,N_7156,N_6802);
nand U8352 (N_8352,N_6730,N_6072);
xor U8353 (N_8353,N_6051,N_7353);
nand U8354 (N_8354,N_6981,N_7083);
nor U8355 (N_8355,N_6082,N_7169);
and U8356 (N_8356,N_6823,N_6965);
or U8357 (N_8357,N_6843,N_6173);
xnor U8358 (N_8358,N_6808,N_6133);
nor U8359 (N_8359,N_6931,N_6106);
xor U8360 (N_8360,N_6059,N_7356);
xnor U8361 (N_8361,N_7307,N_6928);
and U8362 (N_8362,N_6224,N_6195);
or U8363 (N_8363,N_6579,N_6870);
and U8364 (N_8364,N_7004,N_6427);
xnor U8365 (N_8365,N_7493,N_6435);
and U8366 (N_8366,N_7264,N_6479);
or U8367 (N_8367,N_6051,N_6755);
nand U8368 (N_8368,N_6241,N_7193);
or U8369 (N_8369,N_6099,N_6942);
nand U8370 (N_8370,N_7440,N_6738);
nor U8371 (N_8371,N_7157,N_6126);
nor U8372 (N_8372,N_7400,N_6615);
and U8373 (N_8373,N_6134,N_7116);
nor U8374 (N_8374,N_7385,N_6377);
xnor U8375 (N_8375,N_7152,N_6259);
and U8376 (N_8376,N_6234,N_6785);
and U8377 (N_8377,N_6781,N_6327);
or U8378 (N_8378,N_7423,N_7367);
xor U8379 (N_8379,N_7275,N_6723);
nand U8380 (N_8380,N_6119,N_6241);
nor U8381 (N_8381,N_7100,N_6157);
or U8382 (N_8382,N_6376,N_6902);
and U8383 (N_8383,N_6485,N_7436);
nor U8384 (N_8384,N_7372,N_6196);
xnor U8385 (N_8385,N_6712,N_6436);
nand U8386 (N_8386,N_6488,N_7259);
and U8387 (N_8387,N_7060,N_7449);
or U8388 (N_8388,N_6821,N_6579);
nand U8389 (N_8389,N_6256,N_6702);
xnor U8390 (N_8390,N_6715,N_6679);
xnor U8391 (N_8391,N_6100,N_6569);
nor U8392 (N_8392,N_7393,N_6624);
nor U8393 (N_8393,N_6439,N_6097);
nor U8394 (N_8394,N_7299,N_6284);
nand U8395 (N_8395,N_6874,N_6497);
nand U8396 (N_8396,N_6010,N_7203);
nor U8397 (N_8397,N_7355,N_7488);
nor U8398 (N_8398,N_6601,N_6948);
or U8399 (N_8399,N_7280,N_7376);
nand U8400 (N_8400,N_6480,N_6295);
xor U8401 (N_8401,N_6182,N_7394);
nor U8402 (N_8402,N_6285,N_6396);
nand U8403 (N_8403,N_6527,N_6057);
xnor U8404 (N_8404,N_6733,N_7029);
and U8405 (N_8405,N_7171,N_6297);
nand U8406 (N_8406,N_6297,N_6535);
nand U8407 (N_8407,N_6639,N_7406);
xor U8408 (N_8408,N_6523,N_7098);
xnor U8409 (N_8409,N_7149,N_6868);
and U8410 (N_8410,N_6914,N_6741);
nand U8411 (N_8411,N_6640,N_6391);
or U8412 (N_8412,N_6088,N_7038);
nor U8413 (N_8413,N_6517,N_6293);
nand U8414 (N_8414,N_7001,N_7307);
nand U8415 (N_8415,N_7000,N_6516);
nand U8416 (N_8416,N_6972,N_6673);
or U8417 (N_8417,N_7290,N_6891);
and U8418 (N_8418,N_6451,N_7351);
and U8419 (N_8419,N_7420,N_7205);
nand U8420 (N_8420,N_6262,N_7213);
xor U8421 (N_8421,N_6666,N_6515);
xnor U8422 (N_8422,N_6703,N_7023);
xor U8423 (N_8423,N_6898,N_6194);
nand U8424 (N_8424,N_6350,N_7179);
nand U8425 (N_8425,N_6009,N_6215);
or U8426 (N_8426,N_6061,N_6716);
nand U8427 (N_8427,N_6646,N_6055);
nor U8428 (N_8428,N_6629,N_7128);
nor U8429 (N_8429,N_6295,N_6851);
nor U8430 (N_8430,N_7173,N_6471);
and U8431 (N_8431,N_7278,N_7126);
and U8432 (N_8432,N_7175,N_6935);
nor U8433 (N_8433,N_6345,N_6126);
xor U8434 (N_8434,N_6594,N_6390);
nand U8435 (N_8435,N_6457,N_7044);
and U8436 (N_8436,N_7315,N_7405);
nand U8437 (N_8437,N_7116,N_7204);
xnor U8438 (N_8438,N_6873,N_6404);
or U8439 (N_8439,N_6703,N_6338);
nor U8440 (N_8440,N_6379,N_6398);
xnor U8441 (N_8441,N_6328,N_6112);
nor U8442 (N_8442,N_6015,N_6122);
or U8443 (N_8443,N_6249,N_6225);
xnor U8444 (N_8444,N_7213,N_6396);
nand U8445 (N_8445,N_6727,N_7197);
nor U8446 (N_8446,N_6190,N_7199);
or U8447 (N_8447,N_6574,N_7254);
xnor U8448 (N_8448,N_7357,N_6575);
or U8449 (N_8449,N_6984,N_6784);
and U8450 (N_8450,N_6144,N_7316);
nand U8451 (N_8451,N_7237,N_7077);
nand U8452 (N_8452,N_7343,N_6630);
xor U8453 (N_8453,N_7281,N_7474);
nand U8454 (N_8454,N_6323,N_7359);
and U8455 (N_8455,N_7479,N_7254);
and U8456 (N_8456,N_6387,N_6500);
or U8457 (N_8457,N_6977,N_6530);
nand U8458 (N_8458,N_7252,N_6995);
nand U8459 (N_8459,N_6800,N_7185);
nand U8460 (N_8460,N_6108,N_6395);
or U8461 (N_8461,N_6999,N_6529);
nand U8462 (N_8462,N_6878,N_6670);
and U8463 (N_8463,N_6640,N_7156);
nand U8464 (N_8464,N_7431,N_7123);
and U8465 (N_8465,N_6979,N_7098);
xnor U8466 (N_8466,N_7394,N_6148);
or U8467 (N_8467,N_6447,N_6800);
nand U8468 (N_8468,N_6345,N_6609);
xnor U8469 (N_8469,N_6478,N_6672);
nor U8470 (N_8470,N_6956,N_7193);
nand U8471 (N_8471,N_7046,N_6178);
or U8472 (N_8472,N_7385,N_6093);
nor U8473 (N_8473,N_6438,N_6637);
xor U8474 (N_8474,N_6317,N_7347);
or U8475 (N_8475,N_6116,N_6524);
or U8476 (N_8476,N_6488,N_6477);
nand U8477 (N_8477,N_6684,N_7192);
and U8478 (N_8478,N_7206,N_6052);
nor U8479 (N_8479,N_7028,N_6594);
and U8480 (N_8480,N_6916,N_6668);
and U8481 (N_8481,N_7474,N_6333);
nand U8482 (N_8482,N_6249,N_6768);
and U8483 (N_8483,N_6572,N_7028);
or U8484 (N_8484,N_7070,N_6135);
xor U8485 (N_8485,N_6253,N_6308);
nor U8486 (N_8486,N_6271,N_7007);
nor U8487 (N_8487,N_6267,N_6373);
and U8488 (N_8488,N_7125,N_6295);
and U8489 (N_8489,N_6643,N_6831);
or U8490 (N_8490,N_6166,N_7290);
and U8491 (N_8491,N_7059,N_6311);
nand U8492 (N_8492,N_6032,N_6199);
and U8493 (N_8493,N_6278,N_7030);
nor U8494 (N_8494,N_7286,N_6059);
nand U8495 (N_8495,N_7339,N_7447);
or U8496 (N_8496,N_6356,N_6658);
nand U8497 (N_8497,N_6570,N_6956);
nand U8498 (N_8498,N_7017,N_7423);
nor U8499 (N_8499,N_7136,N_6695);
xor U8500 (N_8500,N_6693,N_6935);
and U8501 (N_8501,N_7252,N_6063);
nor U8502 (N_8502,N_7027,N_7155);
nor U8503 (N_8503,N_6270,N_6051);
xor U8504 (N_8504,N_6805,N_7320);
xor U8505 (N_8505,N_6500,N_7442);
or U8506 (N_8506,N_6505,N_7353);
and U8507 (N_8507,N_7241,N_7441);
and U8508 (N_8508,N_7468,N_6318);
or U8509 (N_8509,N_7365,N_6090);
or U8510 (N_8510,N_7356,N_6776);
nor U8511 (N_8511,N_6748,N_7228);
and U8512 (N_8512,N_7274,N_6767);
nor U8513 (N_8513,N_6831,N_6240);
or U8514 (N_8514,N_6643,N_6859);
and U8515 (N_8515,N_6301,N_6773);
xnor U8516 (N_8516,N_6658,N_6196);
nand U8517 (N_8517,N_6298,N_7400);
and U8518 (N_8518,N_6907,N_6900);
nand U8519 (N_8519,N_6980,N_6163);
or U8520 (N_8520,N_7409,N_7247);
or U8521 (N_8521,N_7182,N_6302);
and U8522 (N_8522,N_6985,N_6237);
and U8523 (N_8523,N_6083,N_7399);
or U8524 (N_8524,N_6161,N_7362);
or U8525 (N_8525,N_6329,N_6138);
nor U8526 (N_8526,N_6712,N_6826);
or U8527 (N_8527,N_6876,N_6154);
and U8528 (N_8528,N_6602,N_6560);
xor U8529 (N_8529,N_6208,N_7476);
xnor U8530 (N_8530,N_7339,N_6506);
nand U8531 (N_8531,N_7351,N_7348);
nand U8532 (N_8532,N_6391,N_6723);
nor U8533 (N_8533,N_6039,N_6649);
nand U8534 (N_8534,N_6829,N_6836);
nor U8535 (N_8535,N_6451,N_6195);
nand U8536 (N_8536,N_6101,N_6657);
nand U8537 (N_8537,N_6527,N_7027);
xor U8538 (N_8538,N_7257,N_7483);
xor U8539 (N_8539,N_6116,N_6452);
or U8540 (N_8540,N_6807,N_6658);
or U8541 (N_8541,N_7110,N_7061);
xnor U8542 (N_8542,N_7213,N_6698);
xor U8543 (N_8543,N_6166,N_7367);
xor U8544 (N_8544,N_6279,N_6042);
xnor U8545 (N_8545,N_6245,N_6416);
or U8546 (N_8546,N_6919,N_6360);
or U8547 (N_8547,N_7221,N_6237);
nor U8548 (N_8548,N_6156,N_7485);
and U8549 (N_8549,N_6117,N_7481);
or U8550 (N_8550,N_6748,N_7203);
xor U8551 (N_8551,N_6948,N_6018);
xor U8552 (N_8552,N_7202,N_6877);
xor U8553 (N_8553,N_6350,N_6273);
nor U8554 (N_8554,N_6535,N_6211);
nand U8555 (N_8555,N_7339,N_7304);
nand U8556 (N_8556,N_7377,N_6688);
and U8557 (N_8557,N_6807,N_6020);
nor U8558 (N_8558,N_6063,N_6301);
nor U8559 (N_8559,N_6657,N_7362);
nor U8560 (N_8560,N_6401,N_7221);
or U8561 (N_8561,N_6533,N_6550);
xnor U8562 (N_8562,N_7411,N_6382);
xnor U8563 (N_8563,N_6855,N_7046);
xnor U8564 (N_8564,N_6502,N_7178);
nand U8565 (N_8565,N_6430,N_7488);
or U8566 (N_8566,N_6748,N_6209);
xnor U8567 (N_8567,N_7264,N_6909);
xnor U8568 (N_8568,N_6744,N_6711);
xor U8569 (N_8569,N_6537,N_7106);
xnor U8570 (N_8570,N_7126,N_6329);
and U8571 (N_8571,N_6033,N_7138);
nor U8572 (N_8572,N_7203,N_6505);
nor U8573 (N_8573,N_6632,N_6146);
and U8574 (N_8574,N_6258,N_7079);
and U8575 (N_8575,N_6238,N_6871);
nor U8576 (N_8576,N_6085,N_6389);
or U8577 (N_8577,N_6526,N_6666);
nand U8578 (N_8578,N_7373,N_6687);
nand U8579 (N_8579,N_7365,N_6281);
nor U8580 (N_8580,N_6459,N_6546);
and U8581 (N_8581,N_6038,N_7302);
and U8582 (N_8582,N_7234,N_6324);
nand U8583 (N_8583,N_7481,N_7446);
xor U8584 (N_8584,N_6205,N_6595);
nand U8585 (N_8585,N_7126,N_6151);
nor U8586 (N_8586,N_6664,N_6209);
nand U8587 (N_8587,N_6638,N_6773);
or U8588 (N_8588,N_6780,N_7214);
xnor U8589 (N_8589,N_7481,N_6990);
and U8590 (N_8590,N_6174,N_6872);
nor U8591 (N_8591,N_7056,N_7114);
and U8592 (N_8592,N_7455,N_7214);
or U8593 (N_8593,N_6631,N_6670);
nand U8594 (N_8594,N_7294,N_6478);
nor U8595 (N_8595,N_6372,N_7362);
nor U8596 (N_8596,N_6765,N_6659);
nand U8597 (N_8597,N_6347,N_6209);
xor U8598 (N_8598,N_6390,N_6849);
nor U8599 (N_8599,N_6145,N_7363);
nand U8600 (N_8600,N_6992,N_7201);
xnor U8601 (N_8601,N_7107,N_6506);
or U8602 (N_8602,N_7160,N_6694);
xnor U8603 (N_8603,N_7062,N_6132);
nand U8604 (N_8604,N_6261,N_6697);
nand U8605 (N_8605,N_6941,N_7172);
and U8606 (N_8606,N_6943,N_6114);
xor U8607 (N_8607,N_6442,N_6201);
xnor U8608 (N_8608,N_7050,N_6223);
or U8609 (N_8609,N_6671,N_6498);
nand U8610 (N_8610,N_6592,N_6122);
xor U8611 (N_8611,N_7286,N_7009);
nand U8612 (N_8612,N_6329,N_7226);
or U8613 (N_8613,N_7414,N_6658);
nor U8614 (N_8614,N_7371,N_6919);
nand U8615 (N_8615,N_7211,N_7447);
nor U8616 (N_8616,N_6578,N_6117);
nand U8617 (N_8617,N_7219,N_6529);
nor U8618 (N_8618,N_7267,N_7473);
and U8619 (N_8619,N_7284,N_7312);
xnor U8620 (N_8620,N_7141,N_6149);
nand U8621 (N_8621,N_6804,N_7163);
nor U8622 (N_8622,N_6000,N_7498);
xnor U8623 (N_8623,N_6393,N_7128);
or U8624 (N_8624,N_6504,N_6468);
xnor U8625 (N_8625,N_6444,N_6296);
and U8626 (N_8626,N_7324,N_7497);
xnor U8627 (N_8627,N_6207,N_6427);
nor U8628 (N_8628,N_7411,N_7086);
nand U8629 (N_8629,N_6660,N_6476);
or U8630 (N_8630,N_6391,N_7285);
or U8631 (N_8631,N_7015,N_6044);
nand U8632 (N_8632,N_6273,N_6591);
nand U8633 (N_8633,N_7085,N_6319);
nor U8634 (N_8634,N_6489,N_6095);
nor U8635 (N_8635,N_6362,N_6638);
or U8636 (N_8636,N_6368,N_7044);
nor U8637 (N_8637,N_6610,N_6375);
or U8638 (N_8638,N_6783,N_7129);
nand U8639 (N_8639,N_6388,N_6177);
or U8640 (N_8640,N_6113,N_6540);
and U8641 (N_8641,N_7098,N_6493);
nand U8642 (N_8642,N_6851,N_6404);
xnor U8643 (N_8643,N_6149,N_6450);
and U8644 (N_8644,N_6810,N_6613);
xnor U8645 (N_8645,N_6414,N_7266);
xor U8646 (N_8646,N_6701,N_6370);
or U8647 (N_8647,N_7465,N_6542);
xnor U8648 (N_8648,N_6015,N_6405);
and U8649 (N_8649,N_6208,N_6350);
xor U8650 (N_8650,N_6438,N_7075);
xnor U8651 (N_8651,N_6088,N_6337);
xor U8652 (N_8652,N_6064,N_7076);
nor U8653 (N_8653,N_6253,N_7039);
nor U8654 (N_8654,N_7066,N_6468);
nand U8655 (N_8655,N_6169,N_6936);
or U8656 (N_8656,N_6291,N_7362);
or U8657 (N_8657,N_6166,N_6687);
or U8658 (N_8658,N_7301,N_6332);
nor U8659 (N_8659,N_6794,N_7090);
and U8660 (N_8660,N_6911,N_7002);
or U8661 (N_8661,N_7491,N_7263);
and U8662 (N_8662,N_6546,N_6045);
and U8663 (N_8663,N_6336,N_7060);
xnor U8664 (N_8664,N_6590,N_7294);
nand U8665 (N_8665,N_7400,N_7305);
nor U8666 (N_8666,N_6276,N_6260);
xor U8667 (N_8667,N_6142,N_7164);
or U8668 (N_8668,N_6672,N_7092);
nand U8669 (N_8669,N_7312,N_6083);
or U8670 (N_8670,N_6356,N_6099);
nor U8671 (N_8671,N_6882,N_6432);
xor U8672 (N_8672,N_6961,N_7242);
nor U8673 (N_8673,N_6275,N_7413);
xor U8674 (N_8674,N_6054,N_6261);
nor U8675 (N_8675,N_7117,N_6272);
and U8676 (N_8676,N_6508,N_6180);
nor U8677 (N_8677,N_6549,N_7259);
nor U8678 (N_8678,N_6439,N_6672);
or U8679 (N_8679,N_6150,N_6939);
or U8680 (N_8680,N_7120,N_6866);
or U8681 (N_8681,N_6190,N_6648);
and U8682 (N_8682,N_6290,N_7133);
and U8683 (N_8683,N_6902,N_6899);
and U8684 (N_8684,N_6259,N_7024);
or U8685 (N_8685,N_7404,N_6302);
nor U8686 (N_8686,N_6946,N_7179);
and U8687 (N_8687,N_6231,N_6808);
and U8688 (N_8688,N_6226,N_7424);
xnor U8689 (N_8689,N_6794,N_7345);
nor U8690 (N_8690,N_7035,N_6086);
and U8691 (N_8691,N_7477,N_6654);
nor U8692 (N_8692,N_7113,N_6768);
and U8693 (N_8693,N_6252,N_7332);
xor U8694 (N_8694,N_6563,N_6919);
nand U8695 (N_8695,N_7022,N_6600);
xnor U8696 (N_8696,N_7131,N_7035);
xor U8697 (N_8697,N_6725,N_7425);
xnor U8698 (N_8698,N_6740,N_7116);
xor U8699 (N_8699,N_6076,N_6724);
and U8700 (N_8700,N_6820,N_6319);
nand U8701 (N_8701,N_6226,N_7487);
or U8702 (N_8702,N_6955,N_7003);
and U8703 (N_8703,N_7228,N_6781);
and U8704 (N_8704,N_6997,N_6378);
and U8705 (N_8705,N_6022,N_6637);
nor U8706 (N_8706,N_6422,N_6576);
nor U8707 (N_8707,N_6778,N_6733);
xor U8708 (N_8708,N_6712,N_6718);
or U8709 (N_8709,N_6199,N_6142);
nand U8710 (N_8710,N_7065,N_7164);
and U8711 (N_8711,N_7081,N_6669);
or U8712 (N_8712,N_7151,N_6433);
nand U8713 (N_8713,N_6681,N_7319);
nand U8714 (N_8714,N_7054,N_6639);
nor U8715 (N_8715,N_7231,N_7191);
and U8716 (N_8716,N_6296,N_7388);
xnor U8717 (N_8717,N_6676,N_6011);
xor U8718 (N_8718,N_7388,N_6791);
nand U8719 (N_8719,N_7013,N_6048);
xnor U8720 (N_8720,N_6250,N_6692);
nand U8721 (N_8721,N_7355,N_6979);
or U8722 (N_8722,N_6770,N_6472);
nand U8723 (N_8723,N_6346,N_6177);
xnor U8724 (N_8724,N_7164,N_6220);
nand U8725 (N_8725,N_6544,N_6288);
or U8726 (N_8726,N_7030,N_6813);
xnor U8727 (N_8727,N_6618,N_7188);
nor U8728 (N_8728,N_7478,N_6151);
or U8729 (N_8729,N_6654,N_6447);
nand U8730 (N_8730,N_6714,N_6783);
nand U8731 (N_8731,N_7405,N_6510);
nand U8732 (N_8732,N_6207,N_7293);
nand U8733 (N_8733,N_7308,N_6526);
xor U8734 (N_8734,N_6743,N_6491);
xor U8735 (N_8735,N_7281,N_7362);
nor U8736 (N_8736,N_7223,N_6581);
or U8737 (N_8737,N_7166,N_7448);
xor U8738 (N_8738,N_6834,N_6156);
or U8739 (N_8739,N_6969,N_6938);
nor U8740 (N_8740,N_6098,N_6787);
nor U8741 (N_8741,N_6186,N_7059);
nor U8742 (N_8742,N_6720,N_6117);
and U8743 (N_8743,N_7375,N_6368);
or U8744 (N_8744,N_6846,N_6144);
nand U8745 (N_8745,N_7268,N_7243);
or U8746 (N_8746,N_7372,N_6826);
nand U8747 (N_8747,N_6072,N_6368);
nor U8748 (N_8748,N_6367,N_6235);
xnor U8749 (N_8749,N_6373,N_6646);
nand U8750 (N_8750,N_6310,N_6776);
and U8751 (N_8751,N_6836,N_6312);
or U8752 (N_8752,N_7024,N_6681);
nor U8753 (N_8753,N_6016,N_6801);
nand U8754 (N_8754,N_7464,N_6057);
nor U8755 (N_8755,N_6327,N_7404);
nor U8756 (N_8756,N_6519,N_6358);
nor U8757 (N_8757,N_6494,N_7364);
xnor U8758 (N_8758,N_6598,N_6682);
xnor U8759 (N_8759,N_7215,N_6132);
nand U8760 (N_8760,N_7104,N_7331);
xnor U8761 (N_8761,N_6851,N_6833);
xnor U8762 (N_8762,N_6629,N_6491);
or U8763 (N_8763,N_6463,N_6192);
or U8764 (N_8764,N_6045,N_6541);
or U8765 (N_8765,N_6268,N_7281);
xnor U8766 (N_8766,N_6642,N_6447);
nor U8767 (N_8767,N_6552,N_6498);
nand U8768 (N_8768,N_7019,N_7214);
nor U8769 (N_8769,N_6382,N_6624);
xnor U8770 (N_8770,N_6747,N_7140);
and U8771 (N_8771,N_6981,N_7235);
nor U8772 (N_8772,N_7076,N_6094);
and U8773 (N_8773,N_7415,N_6674);
xnor U8774 (N_8774,N_6129,N_6452);
or U8775 (N_8775,N_6186,N_6033);
nand U8776 (N_8776,N_6444,N_6274);
nor U8777 (N_8777,N_6405,N_6246);
or U8778 (N_8778,N_7023,N_6682);
or U8779 (N_8779,N_7046,N_6081);
and U8780 (N_8780,N_6187,N_7219);
or U8781 (N_8781,N_6800,N_6945);
nor U8782 (N_8782,N_6268,N_7250);
or U8783 (N_8783,N_6821,N_6946);
nand U8784 (N_8784,N_6980,N_6346);
nand U8785 (N_8785,N_6477,N_6539);
nor U8786 (N_8786,N_6635,N_6716);
nor U8787 (N_8787,N_6775,N_6236);
or U8788 (N_8788,N_6143,N_7290);
nor U8789 (N_8789,N_6899,N_6421);
nor U8790 (N_8790,N_7400,N_6716);
nand U8791 (N_8791,N_6354,N_6821);
xnor U8792 (N_8792,N_6009,N_6666);
or U8793 (N_8793,N_6499,N_7208);
and U8794 (N_8794,N_6606,N_7148);
nor U8795 (N_8795,N_7285,N_6916);
xnor U8796 (N_8796,N_6605,N_6579);
and U8797 (N_8797,N_6439,N_6667);
xnor U8798 (N_8798,N_7473,N_6060);
and U8799 (N_8799,N_6849,N_6326);
nor U8800 (N_8800,N_7437,N_6718);
or U8801 (N_8801,N_7234,N_6905);
or U8802 (N_8802,N_6048,N_7411);
or U8803 (N_8803,N_7369,N_6406);
or U8804 (N_8804,N_6335,N_6878);
xor U8805 (N_8805,N_6324,N_6570);
nor U8806 (N_8806,N_6636,N_6998);
xnor U8807 (N_8807,N_6847,N_6712);
nor U8808 (N_8808,N_6110,N_6347);
and U8809 (N_8809,N_6860,N_6077);
and U8810 (N_8810,N_6579,N_7143);
or U8811 (N_8811,N_7382,N_6572);
and U8812 (N_8812,N_6773,N_7248);
xnor U8813 (N_8813,N_6076,N_7132);
or U8814 (N_8814,N_6271,N_6044);
or U8815 (N_8815,N_6215,N_7382);
or U8816 (N_8816,N_6627,N_6657);
or U8817 (N_8817,N_6021,N_7346);
nand U8818 (N_8818,N_6278,N_6929);
nand U8819 (N_8819,N_7411,N_6872);
nor U8820 (N_8820,N_7134,N_6661);
and U8821 (N_8821,N_7355,N_6154);
or U8822 (N_8822,N_7258,N_6676);
nor U8823 (N_8823,N_6678,N_7216);
or U8824 (N_8824,N_7324,N_7090);
nor U8825 (N_8825,N_6120,N_7417);
and U8826 (N_8826,N_6551,N_7259);
or U8827 (N_8827,N_6659,N_6403);
or U8828 (N_8828,N_6250,N_7405);
or U8829 (N_8829,N_6209,N_7432);
and U8830 (N_8830,N_6193,N_6484);
or U8831 (N_8831,N_7111,N_6084);
xor U8832 (N_8832,N_6903,N_6801);
nand U8833 (N_8833,N_6882,N_6512);
xor U8834 (N_8834,N_6191,N_7338);
nand U8835 (N_8835,N_7087,N_7371);
nand U8836 (N_8836,N_6524,N_6715);
or U8837 (N_8837,N_6058,N_6280);
nor U8838 (N_8838,N_6168,N_6206);
nor U8839 (N_8839,N_7475,N_6260);
and U8840 (N_8840,N_7259,N_6739);
and U8841 (N_8841,N_7211,N_6779);
nor U8842 (N_8842,N_6268,N_6696);
nor U8843 (N_8843,N_7018,N_6423);
nand U8844 (N_8844,N_7323,N_6766);
or U8845 (N_8845,N_7027,N_6076);
xor U8846 (N_8846,N_6814,N_6513);
nand U8847 (N_8847,N_6298,N_7256);
or U8848 (N_8848,N_7139,N_7424);
nand U8849 (N_8849,N_7454,N_6286);
or U8850 (N_8850,N_6385,N_7116);
nor U8851 (N_8851,N_6246,N_6944);
and U8852 (N_8852,N_6749,N_7111);
nor U8853 (N_8853,N_7387,N_6846);
nand U8854 (N_8854,N_6786,N_6331);
xnor U8855 (N_8855,N_7443,N_6383);
xor U8856 (N_8856,N_6312,N_7167);
nor U8857 (N_8857,N_6069,N_6481);
or U8858 (N_8858,N_7211,N_6508);
or U8859 (N_8859,N_6335,N_7120);
xor U8860 (N_8860,N_7393,N_6366);
xor U8861 (N_8861,N_6332,N_6627);
or U8862 (N_8862,N_7254,N_6620);
or U8863 (N_8863,N_6641,N_6168);
xnor U8864 (N_8864,N_6805,N_6330);
xor U8865 (N_8865,N_6565,N_6570);
nor U8866 (N_8866,N_6960,N_6139);
and U8867 (N_8867,N_7043,N_6612);
nand U8868 (N_8868,N_6141,N_6136);
nor U8869 (N_8869,N_6882,N_6966);
and U8870 (N_8870,N_6855,N_6819);
or U8871 (N_8871,N_6004,N_6266);
nor U8872 (N_8872,N_6572,N_6239);
nor U8873 (N_8873,N_6089,N_6751);
nor U8874 (N_8874,N_6421,N_6563);
or U8875 (N_8875,N_6114,N_6020);
and U8876 (N_8876,N_6347,N_7167);
nand U8877 (N_8877,N_6479,N_6864);
or U8878 (N_8878,N_7035,N_7493);
xor U8879 (N_8879,N_6929,N_6100);
nand U8880 (N_8880,N_6594,N_6050);
nor U8881 (N_8881,N_6085,N_7196);
nand U8882 (N_8882,N_7273,N_7324);
nor U8883 (N_8883,N_7226,N_6522);
or U8884 (N_8884,N_6104,N_7426);
or U8885 (N_8885,N_7312,N_6151);
nand U8886 (N_8886,N_6876,N_6639);
nor U8887 (N_8887,N_7241,N_6570);
and U8888 (N_8888,N_6036,N_6511);
nand U8889 (N_8889,N_6020,N_6586);
nand U8890 (N_8890,N_7231,N_7175);
or U8891 (N_8891,N_7349,N_6583);
nor U8892 (N_8892,N_6495,N_7370);
xor U8893 (N_8893,N_7152,N_6491);
nor U8894 (N_8894,N_7155,N_6939);
xor U8895 (N_8895,N_6054,N_6262);
xor U8896 (N_8896,N_6802,N_6939);
or U8897 (N_8897,N_6429,N_7428);
nor U8898 (N_8898,N_6715,N_6263);
nor U8899 (N_8899,N_6491,N_7039);
nand U8900 (N_8900,N_6341,N_6890);
xnor U8901 (N_8901,N_6037,N_6069);
or U8902 (N_8902,N_7232,N_7053);
nand U8903 (N_8903,N_6168,N_6594);
or U8904 (N_8904,N_6110,N_6499);
and U8905 (N_8905,N_6372,N_6109);
or U8906 (N_8906,N_6524,N_6477);
or U8907 (N_8907,N_7376,N_6024);
and U8908 (N_8908,N_7192,N_6135);
and U8909 (N_8909,N_6876,N_7488);
and U8910 (N_8910,N_6501,N_7146);
nand U8911 (N_8911,N_7461,N_7128);
and U8912 (N_8912,N_7137,N_6287);
or U8913 (N_8913,N_6188,N_6024);
and U8914 (N_8914,N_7161,N_6508);
and U8915 (N_8915,N_7200,N_6223);
and U8916 (N_8916,N_6618,N_7071);
xnor U8917 (N_8917,N_6435,N_6035);
nand U8918 (N_8918,N_6838,N_6668);
xor U8919 (N_8919,N_6046,N_6594);
or U8920 (N_8920,N_6667,N_6102);
and U8921 (N_8921,N_6901,N_6336);
and U8922 (N_8922,N_6123,N_6698);
nor U8923 (N_8923,N_6302,N_6361);
nand U8924 (N_8924,N_7383,N_7219);
nand U8925 (N_8925,N_7498,N_7281);
nor U8926 (N_8926,N_6871,N_6990);
and U8927 (N_8927,N_6033,N_6154);
xnor U8928 (N_8928,N_6906,N_7394);
or U8929 (N_8929,N_6542,N_6845);
nand U8930 (N_8930,N_6883,N_7269);
and U8931 (N_8931,N_6323,N_6249);
or U8932 (N_8932,N_6533,N_6556);
xor U8933 (N_8933,N_6544,N_7264);
nor U8934 (N_8934,N_7268,N_6501);
nand U8935 (N_8935,N_6553,N_6424);
or U8936 (N_8936,N_6908,N_6120);
nand U8937 (N_8937,N_6248,N_7260);
xnor U8938 (N_8938,N_6019,N_6271);
nand U8939 (N_8939,N_6000,N_7296);
nor U8940 (N_8940,N_6768,N_7287);
and U8941 (N_8941,N_6114,N_6430);
nand U8942 (N_8942,N_6112,N_7340);
nand U8943 (N_8943,N_6855,N_7253);
xor U8944 (N_8944,N_7438,N_6335);
xor U8945 (N_8945,N_6847,N_7160);
or U8946 (N_8946,N_6932,N_6589);
and U8947 (N_8947,N_6841,N_6175);
xnor U8948 (N_8948,N_6997,N_7402);
and U8949 (N_8949,N_7013,N_6201);
and U8950 (N_8950,N_7187,N_6044);
and U8951 (N_8951,N_6799,N_7206);
xnor U8952 (N_8952,N_7320,N_6871);
nand U8953 (N_8953,N_6977,N_6678);
and U8954 (N_8954,N_6183,N_7485);
nor U8955 (N_8955,N_6224,N_6436);
nand U8956 (N_8956,N_6201,N_6752);
nand U8957 (N_8957,N_6985,N_7103);
nand U8958 (N_8958,N_6386,N_6413);
xor U8959 (N_8959,N_6154,N_7171);
nor U8960 (N_8960,N_7284,N_6693);
and U8961 (N_8961,N_7010,N_6621);
or U8962 (N_8962,N_6100,N_7193);
nor U8963 (N_8963,N_7398,N_6333);
or U8964 (N_8964,N_6201,N_7124);
xnor U8965 (N_8965,N_7047,N_6403);
or U8966 (N_8966,N_7430,N_6857);
nor U8967 (N_8967,N_6390,N_7171);
nor U8968 (N_8968,N_6954,N_6104);
or U8969 (N_8969,N_6251,N_7259);
nor U8970 (N_8970,N_6878,N_6552);
and U8971 (N_8971,N_6490,N_6565);
nor U8972 (N_8972,N_6586,N_6478);
or U8973 (N_8973,N_6733,N_6528);
or U8974 (N_8974,N_7408,N_6332);
xor U8975 (N_8975,N_6733,N_6357);
and U8976 (N_8976,N_6339,N_6141);
nor U8977 (N_8977,N_6289,N_6841);
nand U8978 (N_8978,N_6747,N_6899);
nor U8979 (N_8979,N_6894,N_7310);
xnor U8980 (N_8980,N_6287,N_7291);
and U8981 (N_8981,N_6548,N_6938);
nor U8982 (N_8982,N_6180,N_7207);
and U8983 (N_8983,N_6904,N_6694);
nand U8984 (N_8984,N_7378,N_6416);
and U8985 (N_8985,N_7358,N_6110);
nor U8986 (N_8986,N_7396,N_6892);
nor U8987 (N_8987,N_7431,N_7189);
nor U8988 (N_8988,N_6479,N_7386);
xnor U8989 (N_8989,N_7353,N_6464);
xor U8990 (N_8990,N_6746,N_6078);
nand U8991 (N_8991,N_6060,N_7381);
or U8992 (N_8992,N_7064,N_6927);
nor U8993 (N_8993,N_6942,N_6032);
nand U8994 (N_8994,N_7071,N_7443);
nand U8995 (N_8995,N_6809,N_7429);
and U8996 (N_8996,N_6172,N_6282);
nand U8997 (N_8997,N_6842,N_7438);
xor U8998 (N_8998,N_7441,N_6465);
and U8999 (N_8999,N_6360,N_7205);
and U9000 (N_9000,N_7526,N_7722);
or U9001 (N_9001,N_8843,N_8543);
nor U9002 (N_9002,N_8077,N_8133);
or U9003 (N_9003,N_8373,N_8545);
nor U9004 (N_9004,N_8464,N_8780);
xnor U9005 (N_9005,N_8598,N_7568);
xor U9006 (N_9006,N_8054,N_8492);
and U9007 (N_9007,N_8755,N_8297);
and U9008 (N_9008,N_7583,N_8443);
and U9009 (N_9009,N_7696,N_7978);
nand U9010 (N_9010,N_8904,N_7604);
nand U9011 (N_9011,N_8895,N_7532);
and U9012 (N_9012,N_8717,N_8105);
nor U9013 (N_9013,N_8031,N_8789);
xor U9014 (N_9014,N_8651,N_8983);
nand U9015 (N_9015,N_8971,N_8461);
nor U9016 (N_9016,N_8158,N_8231);
nor U9017 (N_9017,N_7525,N_7634);
nor U9018 (N_9018,N_7614,N_7761);
nand U9019 (N_9019,N_7742,N_7562);
and U9020 (N_9020,N_7951,N_8756);
and U9021 (N_9021,N_8529,N_7654);
xnor U9022 (N_9022,N_8386,N_7503);
and U9023 (N_9023,N_7546,N_8124);
or U9024 (N_9024,N_8264,N_8699);
nand U9025 (N_9025,N_8757,N_7536);
and U9026 (N_9026,N_8086,N_8076);
xnor U9027 (N_9027,N_7796,N_8608);
and U9028 (N_9028,N_8592,N_8857);
or U9029 (N_9029,N_8030,N_8644);
nand U9030 (N_9030,N_8062,N_7926);
and U9031 (N_9031,N_7640,N_8694);
xnor U9032 (N_9032,N_8115,N_8779);
and U9033 (N_9033,N_7585,N_8819);
and U9034 (N_9034,N_7533,N_8700);
or U9035 (N_9035,N_7650,N_8063);
nor U9036 (N_9036,N_8791,N_8449);
nor U9037 (N_9037,N_8527,N_8265);
nand U9038 (N_9038,N_8419,N_8479);
nand U9039 (N_9039,N_8456,N_8038);
nor U9040 (N_9040,N_8961,N_8211);
or U9041 (N_9041,N_7707,N_8932);
nor U9042 (N_9042,N_7857,N_8248);
and U9043 (N_9043,N_8067,N_8007);
nand U9044 (N_9044,N_7944,N_7671);
xnor U9045 (N_9045,N_7972,N_8320);
nor U9046 (N_9046,N_8128,N_8168);
and U9047 (N_9047,N_8226,N_8083);
and U9048 (N_9048,N_8438,N_7805);
and U9049 (N_9049,N_8247,N_8179);
xor U9050 (N_9050,N_8869,N_8368);
nand U9051 (N_9051,N_8627,N_8950);
nor U9052 (N_9052,N_8222,N_8065);
and U9053 (N_9053,N_8984,N_8890);
or U9054 (N_9054,N_8974,N_7779);
nor U9055 (N_9055,N_7517,N_7806);
and U9056 (N_9056,N_8671,N_8965);
nor U9057 (N_9057,N_7811,N_7991);
nand U9058 (N_9058,N_8737,N_8333);
nor U9059 (N_9059,N_8859,N_8421);
xnor U9060 (N_9060,N_7687,N_7595);
xor U9061 (N_9061,N_8880,N_8860);
nand U9062 (N_9062,N_8216,N_8398);
or U9063 (N_9063,N_8794,N_7860);
nand U9064 (N_9064,N_7572,N_8374);
nand U9065 (N_9065,N_8992,N_8662);
xor U9066 (N_9066,N_8707,N_8462);
nor U9067 (N_9067,N_8810,N_8519);
nor U9068 (N_9068,N_7947,N_7581);
xor U9069 (N_9069,N_7518,N_8500);
nand U9070 (N_9070,N_8738,N_8162);
nor U9071 (N_9071,N_7768,N_7727);
nand U9072 (N_9072,N_7635,N_8146);
and U9073 (N_9073,N_7890,N_7868);
nor U9074 (N_9074,N_8595,N_8301);
nor U9075 (N_9075,N_8748,N_8256);
and U9076 (N_9076,N_8724,N_7704);
xnor U9077 (N_9077,N_8006,N_8808);
xor U9078 (N_9078,N_8477,N_8329);
or U9079 (N_9079,N_8742,N_7826);
xnor U9080 (N_9080,N_7793,N_7919);
nor U9081 (N_9081,N_8713,N_8305);
or U9082 (N_9082,N_8420,N_8385);
xnor U9083 (N_9083,N_7829,N_8568);
and U9084 (N_9084,N_8437,N_7611);
nand U9085 (N_9085,N_7542,N_7885);
xnor U9086 (N_9086,N_8383,N_7981);
or U9087 (N_9087,N_8528,N_8560);
xnor U9088 (N_9088,N_8704,N_8966);
or U9089 (N_9089,N_7932,N_8440);
nor U9090 (N_9090,N_7644,N_8572);
xnor U9091 (N_9091,N_7748,N_8986);
nand U9092 (N_9092,N_8463,N_7553);
nand U9093 (N_9093,N_8823,N_7565);
or U9094 (N_9094,N_8814,N_7739);
xnor U9095 (N_9095,N_7965,N_7788);
and U9096 (N_9096,N_8559,N_8195);
nor U9097 (N_9097,N_7942,N_7712);
or U9098 (N_9098,N_8523,N_7612);
xor U9099 (N_9099,N_8059,N_7856);
or U9100 (N_9100,N_7916,N_8027);
and U9101 (N_9101,N_8299,N_7523);
or U9102 (N_9102,N_7818,N_8563);
or U9103 (N_9103,N_7744,N_8404);
and U9104 (N_9104,N_8000,N_7705);
and U9105 (N_9105,N_8130,N_8982);
and U9106 (N_9106,N_8744,N_8617);
nor U9107 (N_9107,N_8073,N_8611);
xor U9108 (N_9108,N_8505,N_8589);
and U9109 (N_9109,N_8706,N_7809);
xnor U9110 (N_9110,N_8858,N_7958);
nand U9111 (N_9111,N_8106,N_7545);
or U9112 (N_9112,N_8176,N_8257);
and U9113 (N_9113,N_8005,N_8618);
or U9114 (N_9114,N_8612,N_7871);
or U9115 (N_9115,N_8402,N_7694);
xnor U9116 (N_9116,N_7680,N_8583);
nor U9117 (N_9117,N_8674,N_8802);
nand U9118 (N_9118,N_8021,N_7887);
nand U9119 (N_9119,N_8003,N_7827);
xnor U9120 (N_9120,N_7957,N_8512);
nor U9121 (N_9121,N_7921,N_7560);
nand U9122 (N_9122,N_8164,N_7952);
nor U9123 (N_9123,N_8837,N_7756);
and U9124 (N_9124,N_8854,N_8769);
nand U9125 (N_9125,N_7683,N_8131);
nand U9126 (N_9126,N_8225,N_7927);
nand U9127 (N_9127,N_7681,N_8958);
xor U9128 (N_9128,N_8422,N_8088);
xor U9129 (N_9129,N_8535,N_7516);
nor U9130 (N_9130,N_8927,N_8378);
xor U9131 (N_9131,N_8401,N_8145);
nand U9132 (N_9132,N_7902,N_8676);
nor U9133 (N_9133,N_8471,N_8278);
and U9134 (N_9134,N_7808,N_8571);
and U9135 (N_9135,N_8580,N_7636);
nor U9136 (N_9136,N_8331,N_8046);
nand U9137 (N_9137,N_8531,N_8008);
and U9138 (N_9138,N_8254,N_8291);
nor U9139 (N_9139,N_7875,N_8630);
xor U9140 (N_9140,N_8116,N_8460);
nand U9141 (N_9141,N_8185,N_8240);
nor U9142 (N_9142,N_7743,N_7616);
nor U9143 (N_9143,N_7955,N_7997);
and U9144 (N_9144,N_7782,N_8962);
or U9145 (N_9145,N_8605,N_8922);
xnor U9146 (N_9146,N_7734,N_8221);
or U9147 (N_9147,N_7894,N_8103);
nand U9148 (N_9148,N_8619,N_8872);
xor U9149 (N_9149,N_8661,N_8767);
or U9150 (N_9150,N_8784,N_8358);
and U9151 (N_9151,N_8107,N_8715);
or U9152 (N_9152,N_7508,N_8082);
or U9153 (N_9153,N_8308,N_7945);
or U9154 (N_9154,N_7822,N_8613);
and U9155 (N_9155,N_7594,N_7755);
nor U9156 (N_9156,N_7765,N_8285);
xnor U9157 (N_9157,N_7661,N_8926);
and U9158 (N_9158,N_8815,N_8692);
xor U9159 (N_9159,N_8089,N_7576);
or U9160 (N_9160,N_8346,N_8154);
nand U9161 (N_9161,N_8733,N_8963);
nor U9162 (N_9162,N_8553,N_8988);
and U9163 (N_9163,N_8208,N_8518);
nand U9164 (N_9164,N_7941,N_8311);
and U9165 (N_9165,N_8242,N_8336);
nand U9166 (N_9166,N_7590,N_8989);
and U9167 (N_9167,N_7676,N_7600);
nand U9168 (N_9168,N_8213,N_8524);
nand U9169 (N_9169,N_8180,N_8656);
or U9170 (N_9170,N_7895,N_8809);
or U9171 (N_9171,N_8499,N_7881);
xnor U9172 (N_9172,N_8501,N_8881);
or U9173 (N_9173,N_8975,N_7917);
or U9174 (N_9174,N_8831,N_8098);
or U9175 (N_9175,N_8224,N_7720);
or U9176 (N_9176,N_7552,N_8749);
and U9177 (N_9177,N_8842,N_7989);
xor U9178 (N_9178,N_8604,N_8788);
or U9179 (N_9179,N_8032,N_8636);
or U9180 (N_9180,N_8365,N_8758);
or U9181 (N_9181,N_8396,N_8973);
and U9182 (N_9182,N_8428,N_7961);
and U9183 (N_9183,N_8773,N_8472);
or U9184 (N_9184,N_8141,N_7638);
nand U9185 (N_9185,N_8425,N_8610);
xor U9186 (N_9186,N_7897,N_7848);
or U9187 (N_9187,N_7964,N_8313);
or U9188 (N_9188,N_8522,N_8393);
or U9189 (N_9189,N_8108,N_8478);
nand U9190 (N_9190,N_8623,N_8771);
nor U9191 (N_9191,N_7799,N_8670);
nand U9192 (N_9192,N_8684,N_8805);
and U9193 (N_9193,N_8969,N_8068);
or U9194 (N_9194,N_8639,N_8266);
xor U9195 (N_9195,N_7719,N_8693);
nand U9196 (N_9196,N_7915,N_7586);
nor U9197 (N_9197,N_7535,N_8300);
nand U9198 (N_9198,N_7759,N_7506);
xor U9199 (N_9199,N_8734,N_8918);
or U9200 (N_9200,N_8360,N_8936);
xor U9201 (N_9201,N_8244,N_7729);
and U9202 (N_9202,N_8600,N_8468);
nor U9203 (N_9203,N_8847,N_7675);
or U9204 (N_9204,N_7976,N_7962);
and U9205 (N_9205,N_8296,N_7994);
and U9206 (N_9206,N_8286,N_8095);
nor U9207 (N_9207,N_8439,N_8429);
or U9208 (N_9208,N_8978,N_8538);
nor U9209 (N_9209,N_7835,N_8444);
xnor U9210 (N_9210,N_8453,N_8807);
nor U9211 (N_9211,N_7664,N_8747);
and U9212 (N_9212,N_8570,N_7556);
xor U9213 (N_9213,N_7670,N_7567);
nor U9214 (N_9214,N_7723,N_7602);
and U9215 (N_9215,N_8775,N_8084);
nand U9216 (N_9216,N_7524,N_7544);
and U9217 (N_9217,N_8503,N_7781);
and U9218 (N_9218,N_8061,N_7682);
and U9219 (N_9219,N_8811,N_7702);
and U9220 (N_9220,N_8996,N_8935);
nand U9221 (N_9221,N_7933,N_8793);
and U9222 (N_9222,N_7867,N_8885);
and U9223 (N_9223,N_8252,N_7775);
or U9224 (N_9224,N_8347,N_8283);
nor U9225 (N_9225,N_8657,N_7833);
or U9226 (N_9226,N_8215,N_7543);
or U9227 (N_9227,N_7691,N_7579);
or U9228 (N_9228,N_8551,N_8343);
nand U9229 (N_9229,N_7814,N_7813);
xnor U9230 (N_9230,N_8884,N_8362);
or U9231 (N_9231,N_8376,N_7564);
and U9232 (N_9232,N_8999,N_7569);
or U9233 (N_9233,N_7943,N_7732);
nand U9234 (N_9234,N_8205,N_8060);
and U9235 (N_9235,N_7738,N_7975);
xor U9236 (N_9236,N_8435,N_7577);
and U9237 (N_9237,N_8199,N_7555);
or U9238 (N_9238,N_8016,N_8044);
or U9239 (N_9239,N_8410,N_8530);
nor U9240 (N_9240,N_8658,N_8483);
or U9241 (N_9241,N_8117,N_7832);
nand U9242 (N_9242,N_8263,N_8997);
or U9243 (N_9243,N_8189,N_8272);
or U9244 (N_9244,N_8725,N_7721);
nor U9245 (N_9245,N_7618,N_8678);
nor U9246 (N_9246,N_8774,N_8157);
xor U9247 (N_9247,N_8597,N_7686);
or U9248 (N_9248,N_7783,N_8465);
and U9249 (N_9249,N_7766,N_7772);
nor U9250 (N_9250,N_8609,N_8907);
nor U9251 (N_9251,N_8941,N_7821);
xnor U9252 (N_9252,N_7728,N_8798);
xor U9253 (N_9253,N_8191,N_7900);
or U9254 (N_9254,N_8281,N_7643);
or U9255 (N_9255,N_7846,N_8790);
and U9256 (N_9256,N_8484,N_8536);
nor U9257 (N_9257,N_7665,N_8140);
or U9258 (N_9258,N_8898,N_7531);
or U9259 (N_9259,N_7763,N_8387);
or U9260 (N_9260,N_8127,N_8905);
or U9261 (N_9261,N_8085,N_8901);
and U9262 (N_9262,N_7841,N_8136);
nor U9263 (N_9263,N_7538,N_7653);
or U9264 (N_9264,N_7886,N_7971);
nor U9265 (N_9265,N_8840,N_8893);
or U9266 (N_9266,N_7801,N_8186);
or U9267 (N_9267,N_8718,N_7777);
xor U9268 (N_9268,N_8233,N_8532);
and U9269 (N_9269,N_8667,N_7790);
and U9270 (N_9270,N_7948,N_7685);
or U9271 (N_9271,N_7791,N_8304);
xnor U9272 (N_9272,N_8721,N_7896);
nand U9273 (N_9273,N_8269,N_8327);
and U9274 (N_9274,N_8293,N_7865);
nand U9275 (N_9275,N_7879,N_7780);
xor U9276 (N_9276,N_7774,N_8175);
or U9277 (N_9277,N_8506,N_8002);
nand U9278 (N_9278,N_8614,N_8167);
nand U9279 (N_9279,N_8070,N_8516);
nor U9280 (N_9280,N_8835,N_7819);
and U9281 (N_9281,N_7699,N_7607);
nand U9282 (N_9282,N_8397,N_8372);
xor U9283 (N_9283,N_7645,N_8920);
xnor U9284 (N_9284,N_8566,N_7642);
xnor U9285 (N_9285,N_8625,N_7629);
xnor U9286 (N_9286,N_7619,N_7700);
xor U9287 (N_9287,N_8114,N_8672);
nor U9288 (N_9288,N_8933,N_7776);
nand U9289 (N_9289,N_8727,N_8900);
xnor U9290 (N_9290,N_8228,N_8491);
and U9291 (N_9291,N_8206,N_8212);
xnor U9292 (N_9292,N_8648,N_8925);
or U9293 (N_9293,N_8943,N_8868);
nand U9294 (N_9294,N_7563,N_7733);
or U9295 (N_9295,N_8877,N_8822);
nand U9296 (N_9296,N_8637,N_8232);
nor U9297 (N_9297,N_7514,N_8151);
and U9298 (N_9298,N_8391,N_8147);
nand U9299 (N_9299,N_7903,N_7548);
xor U9300 (N_9300,N_8663,N_7834);
or U9301 (N_9301,N_8357,N_8812);
and U9302 (N_9302,N_8569,N_8328);
nand U9303 (N_9303,N_8203,N_7864);
xor U9304 (N_9304,N_7824,N_8352);
or U9305 (N_9305,N_8403,N_7693);
nor U9306 (N_9306,N_8087,N_8409);
nor U9307 (N_9307,N_8366,N_7937);
xor U9308 (N_9308,N_8041,N_8253);
or U9309 (N_9309,N_8298,N_8099);
nand U9310 (N_9310,N_8856,N_8894);
xnor U9311 (N_9311,N_8497,N_8855);
and U9312 (N_9312,N_7689,N_8792);
or U9313 (N_9313,N_8778,N_8934);
nand U9314 (N_9314,N_8200,N_7850);
nand U9315 (N_9315,N_7551,N_7575);
nor U9316 (N_9316,N_7914,N_8581);
xor U9317 (N_9317,N_7519,N_7547);
and U9318 (N_9318,N_7566,N_7767);
and U9319 (N_9319,N_8955,N_8056);
and U9320 (N_9320,N_8332,N_8964);
nor U9321 (N_9321,N_8817,N_8028);
and U9322 (N_9322,N_7984,N_8818);
nor U9323 (N_9323,N_8797,N_8590);
and U9324 (N_9324,N_8921,N_8621);
nand U9325 (N_9325,N_8534,N_8183);
nor U9326 (N_9326,N_8122,N_8687);
and U9327 (N_9327,N_8017,N_8284);
nand U9328 (N_9328,N_8555,N_8093);
or U9329 (N_9329,N_8258,N_8586);
xor U9330 (N_9330,N_7678,N_8628);
nor U9331 (N_9331,N_8040,N_8760);
nand U9332 (N_9332,N_7561,N_8564);
and U9333 (N_9333,N_8526,N_8190);
nor U9334 (N_9334,N_7537,N_8159);
xnor U9335 (N_9335,N_8335,N_8649);
and U9336 (N_9336,N_7620,N_7549);
nor U9337 (N_9337,N_8763,N_8413);
xor U9338 (N_9338,N_8697,N_7847);
or U9339 (N_9339,N_8367,N_8406);
nor U9340 (N_9340,N_8118,N_7880);
nor U9341 (N_9341,N_7628,N_8556);
xor U9342 (N_9342,N_8187,N_8681);
and U9343 (N_9343,N_7854,N_7501);
nor U9344 (N_9344,N_7690,N_8677);
nand U9345 (N_9345,N_8507,N_8533);
nor U9346 (N_9346,N_7657,N_8037);
xor U9347 (N_9347,N_8902,N_8875);
and U9348 (N_9348,N_8223,N_8695);
nand U9349 (N_9349,N_8431,N_8680);
xor U9350 (N_9350,N_7922,N_7934);
or U9351 (N_9351,N_8754,N_8149);
or U9352 (N_9352,N_8342,N_8457);
and U9353 (N_9353,N_7874,N_7803);
nor U9354 (N_9354,N_8390,N_7709);
nand U9355 (N_9355,N_8081,N_8137);
nor U9356 (N_9356,N_7999,N_8730);
and U9357 (N_9357,N_7633,N_7534);
and U9358 (N_9358,N_8091,N_8701);
nand U9359 (N_9359,N_7882,N_8683);
nor U9360 (N_9360,N_8547,N_8451);
nand U9361 (N_9361,N_7603,N_8169);
nor U9362 (N_9362,N_8234,N_7816);
nand U9363 (N_9363,N_7504,N_8192);
xor U9364 (N_9364,N_8277,N_8979);
nor U9365 (N_9365,N_7672,N_7870);
nand U9366 (N_9366,N_7507,N_8455);
nor U9367 (N_9367,N_7988,N_7977);
nand U9368 (N_9368,N_8772,N_8510);
nand U9369 (N_9369,N_7509,N_8178);
nand U9370 (N_9370,N_7598,N_8753);
nor U9371 (N_9371,N_7936,N_7527);
nand U9372 (N_9372,N_8567,N_8156);
nor U9373 (N_9373,N_8267,N_8655);
nand U9374 (N_9374,N_8541,N_8018);
nor U9375 (N_9375,N_8426,N_8274);
and U9376 (N_9376,N_7979,N_7584);
and U9377 (N_9377,N_7858,N_8696);
or U9378 (N_9378,N_7674,N_8584);
nand U9379 (N_9379,N_8645,N_8953);
and U9380 (N_9380,N_8740,N_7753);
xor U9381 (N_9381,N_8043,N_7695);
xor U9382 (N_9382,N_7578,N_7502);
nand U9383 (N_9383,N_8494,N_8762);
nor U9384 (N_9384,N_8827,N_7684);
xor U9385 (N_9385,N_8712,N_8624);
xnor U9386 (N_9386,N_8289,N_8412);
nor U9387 (N_9387,N_7980,N_8923);
nand U9388 (N_9388,N_8972,N_8602);
nand U9389 (N_9389,N_7648,N_8090);
and U9390 (N_9390,N_8042,N_8408);
or U9391 (N_9391,N_7574,N_8876);
or U9392 (N_9392,N_8682,N_8321);
nand U9393 (N_9393,N_7520,N_8488);
nor U9394 (N_9394,N_8853,N_8652);
nand U9395 (N_9395,N_8476,N_8865);
and U9396 (N_9396,N_7815,N_8669);
or U9397 (N_9397,N_8182,N_8585);
nand U9398 (N_9398,N_8825,N_8970);
or U9399 (N_9399,N_8646,N_8375);
nand U9400 (N_9400,N_8270,N_8152);
or U9401 (N_9401,N_8887,N_8036);
nor U9402 (N_9402,N_8739,N_8325);
and U9403 (N_9403,N_7953,N_8150);
nor U9404 (N_9404,N_7913,N_7697);
and U9405 (N_9405,N_8261,N_8641);
or U9406 (N_9406,N_8642,N_7986);
xnor U9407 (N_9407,N_8729,N_8448);
nor U9408 (N_9408,N_8801,N_8917);
and U9409 (N_9409,N_8851,N_8132);
xor U9410 (N_9410,N_7737,N_8048);
nand U9411 (N_9411,N_8142,N_8698);
or U9412 (N_9412,N_8606,N_8356);
nand U9413 (N_9413,N_8026,N_8879);
and U9414 (N_9414,N_8348,N_7830);
xnor U9415 (N_9415,N_8948,N_7500);
and U9416 (N_9416,N_8591,N_8783);
or U9417 (N_9417,N_7795,N_8470);
and U9418 (N_9418,N_7995,N_7610);
nor U9419 (N_9419,N_8450,N_8496);
xor U9420 (N_9420,N_8867,N_8521);
nand U9421 (N_9421,N_7667,N_7923);
nand U9422 (N_9422,N_8295,N_7609);
xnor U9423 (N_9423,N_8650,N_7863);
nand U9424 (N_9424,N_7859,N_7898);
nor U9425 (N_9425,N_8990,N_8275);
nor U9426 (N_9426,N_7853,N_7513);
nand U9427 (N_9427,N_8125,N_8307);
and U9428 (N_9428,N_8746,N_8075);
and U9429 (N_9429,N_8806,N_7877);
or U9430 (N_9430,N_7908,N_8334);
and U9431 (N_9431,N_7646,N_8259);
nor U9432 (N_9432,N_8554,N_8345);
xnor U9433 (N_9433,N_8863,N_7884);
or U9434 (N_9434,N_8726,N_8719);
and U9435 (N_9435,N_7855,N_7869);
or U9436 (N_9436,N_8849,N_8838);
nor U9437 (N_9437,N_7929,N_8765);
nand U9438 (N_9438,N_8350,N_8024);
nand U9439 (N_9439,N_8094,N_8852);
nor U9440 (N_9440,N_8013,N_8097);
nor U9441 (N_9441,N_7652,N_8012);
nor U9442 (N_9442,N_8751,N_8947);
and U9443 (N_9443,N_8382,N_7828);
and U9444 (N_9444,N_7852,N_8931);
nand U9445 (N_9445,N_7637,N_7956);
nor U9446 (N_9446,N_8689,N_8513);
and U9447 (N_9447,N_8020,N_8803);
xnor U9448 (N_9448,N_8573,N_7679);
nor U9449 (N_9449,N_8782,N_7925);
nand U9450 (N_9450,N_7836,N_8777);
or U9451 (N_9451,N_7541,N_8493);
and U9452 (N_9452,N_7905,N_7985);
xnor U9453 (N_9453,N_7639,N_8883);
and U9454 (N_9454,N_8959,N_8930);
xor U9455 (N_9455,N_8903,N_8045);
or U9456 (N_9456,N_8010,N_8705);
xor U9457 (N_9457,N_8498,N_8317);
xnor U9458 (N_9458,N_8702,N_8720);
nand U9459 (N_9459,N_8640,N_8906);
or U9460 (N_9460,N_8781,N_8339);
nor U9461 (N_9461,N_7591,N_7792);
or U9462 (N_9462,N_8025,N_8578);
or U9463 (N_9463,N_8514,N_7539);
and U9464 (N_9464,N_8861,N_8138);
nand U9465 (N_9465,N_8341,N_8834);
nor U9466 (N_9466,N_8210,N_7655);
and U9467 (N_9467,N_8685,N_8550);
or U9468 (N_9468,N_8520,N_8480);
or U9469 (N_9469,N_8482,N_7521);
nor U9470 (N_9470,N_7842,N_7771);
or U9471 (N_9471,N_8029,N_7571);
and U9472 (N_9472,N_8079,N_8135);
xor U9473 (N_9473,N_7787,N_8710);
or U9474 (N_9474,N_8184,N_7641);
or U9475 (N_9475,N_7838,N_7724);
nor U9476 (N_9476,N_8324,N_8458);
and U9477 (N_9477,N_8220,N_7715);
or U9478 (N_9478,N_8490,N_7663);
nor U9479 (N_9479,N_8246,N_8473);
or U9480 (N_9480,N_7613,N_7725);
or U9481 (N_9481,N_8968,N_7998);
nor U9482 (N_9482,N_8229,N_8634);
and U9483 (N_9483,N_8459,N_8829);
and U9484 (N_9484,N_7741,N_8442);
xor U9485 (N_9485,N_8911,N_8326);
nand U9486 (N_9486,N_8243,N_8928);
and U9487 (N_9487,N_7752,N_8282);
nand U9488 (N_9488,N_8123,N_7615);
nor U9489 (N_9489,N_8537,N_7892);
or U9490 (N_9490,N_7878,N_8743);
nor U9491 (N_9491,N_8828,N_7557);
and U9492 (N_9492,N_8236,N_8113);
xor U9493 (N_9493,N_8174,N_8280);
or U9494 (N_9494,N_8908,N_8632);
xnor U9495 (N_9495,N_8287,N_8576);
nor U9496 (N_9496,N_7960,N_8249);
nand U9497 (N_9497,N_8489,N_7747);
nor U9498 (N_9498,N_7992,N_7889);
xor U9499 (N_9499,N_8635,N_7589);
nand U9500 (N_9500,N_8804,N_7625);
nand U9501 (N_9501,N_8069,N_7966);
or U9502 (N_9502,N_8631,N_8262);
nand U9503 (N_9503,N_7930,N_8194);
nor U9504 (N_9504,N_8209,N_7528);
and U9505 (N_9505,N_8951,N_8795);
nand U9506 (N_9506,N_8330,N_8690);
and U9507 (N_9507,N_8485,N_7730);
nor U9508 (N_9508,N_8776,N_7658);
nor U9509 (N_9509,N_8714,N_7716);
or U9510 (N_9510,N_7599,N_8957);
nand U9511 (N_9511,N_8502,N_8467);
nor U9512 (N_9512,N_7907,N_7866);
and U9513 (N_9513,N_7911,N_7820);
nor U9514 (N_9514,N_7800,N_7605);
or U9515 (N_9515,N_8049,N_8873);
and U9516 (N_9516,N_7659,N_7924);
nand U9517 (N_9517,N_8882,N_8668);
nor U9518 (N_9518,N_8316,N_8616);
or U9519 (N_9519,N_8991,N_8064);
and U9520 (N_9520,N_7668,N_8389);
nor U9521 (N_9521,N_7950,N_7649);
nand U9522 (N_9522,N_8956,N_8197);
nor U9523 (N_9523,N_7983,N_8237);
nor U9524 (N_9524,N_8441,N_7910);
nand U9525 (N_9525,N_8596,N_8799);
nand U9526 (N_9526,N_7918,N_7530);
or U9527 (N_9527,N_7851,N_8736);
xnor U9528 (N_9528,N_8411,N_7651);
nand U9529 (N_9529,N_8314,N_8377);
nor U9530 (N_9530,N_7617,N_8121);
xor U9531 (N_9531,N_7726,N_8312);
nor U9532 (N_9532,N_8525,N_8349);
and U9533 (N_9533,N_8445,N_8659);
xor U9534 (N_9534,N_8309,N_7624);
xnor U9535 (N_9535,N_8100,N_8434);
and U9536 (N_9536,N_8509,N_7701);
nand U9537 (N_9537,N_8770,N_7789);
nand U9538 (N_9538,N_8134,N_7606);
and U9539 (N_9539,N_8557,N_8998);
and U9540 (N_9540,N_8430,N_8322);
nor U9541 (N_9541,N_8227,N_8980);
and U9542 (N_9542,N_8848,N_8104);
nor U9543 (N_9543,N_8171,N_8954);
nor U9544 (N_9544,N_8014,N_7626);
xor U9545 (N_9545,N_8976,N_7901);
nand U9546 (N_9546,N_8166,N_7698);
xnor U9547 (N_9547,N_8379,N_8504);
xor U9548 (N_9548,N_8279,N_7845);
or U9549 (N_9549,N_8864,N_7825);
or U9550 (N_9550,N_8004,N_7601);
nor U9551 (N_9551,N_8474,N_7770);
and U9552 (N_9552,N_8723,N_8665);
nor U9553 (N_9553,N_8447,N_7596);
nand U9554 (N_9554,N_8845,N_8866);
nand U9555 (N_9555,N_8102,N_7677);
and U9556 (N_9556,N_8071,N_8653);
and U9557 (N_9557,N_8238,N_8977);
or U9558 (N_9558,N_7893,N_8546);
or U9559 (N_9559,N_8985,N_7673);
xor U9560 (N_9560,N_8562,N_8288);
nor U9561 (N_9561,N_7891,N_8198);
xnor U9562 (N_9562,N_8074,N_8841);
and U9563 (N_9563,N_8732,N_8338);
and U9564 (N_9564,N_8561,N_7876);
nor U9565 (N_9565,N_8673,N_7843);
xnor U9566 (N_9566,N_8009,N_8735);
nand U9567 (N_9567,N_8622,N_8416);
nor U9568 (N_9568,N_8599,N_7840);
or U9569 (N_9569,N_7839,N_8160);
and U9570 (N_9570,N_7735,N_8015);
xor U9571 (N_9571,N_7872,N_8643);
nor U9572 (N_9572,N_7703,N_7762);
nor U9573 (N_9573,N_8981,N_8188);
nand U9574 (N_9574,N_8741,N_8432);
and U9575 (N_9575,N_8548,N_8235);
nand U9576 (N_9576,N_7883,N_8914);
nand U9577 (N_9577,N_8638,N_8315);
xnor U9578 (N_9578,N_8033,N_7597);
nand U9579 (N_9579,N_7587,N_8139);
and U9580 (N_9580,N_8620,N_7529);
nor U9581 (N_9581,N_8303,N_7623);
or U9582 (N_9582,N_8539,N_8414);
or U9583 (N_9583,N_7906,N_8542);
nor U9584 (N_9584,N_8423,N_8392);
nand U9585 (N_9585,N_7794,N_7582);
nand U9586 (N_9586,N_8201,N_8844);
nand U9587 (N_9587,N_8626,N_7550);
or U9588 (N_9588,N_8761,N_7931);
nor U9589 (N_9589,N_7692,N_8218);
nand U9590 (N_9590,N_8369,N_7573);
nand U9591 (N_9591,N_8294,N_8886);
xnor U9592 (N_9592,N_8370,N_8675);
nor U9593 (N_9593,N_8945,N_7804);
nand U9594 (N_9594,N_7993,N_8424);
nand U9595 (N_9595,N_7662,N_8023);
nor U9596 (N_9596,N_8053,N_7939);
nor U9597 (N_9597,N_7982,N_8558);
xnor U9598 (N_9598,N_8745,N_8394);
nor U9599 (N_9599,N_8306,N_7647);
nand U9600 (N_9600,N_8155,N_7688);
nor U9601 (N_9601,N_8072,N_7522);
or U9602 (N_9602,N_8380,N_7823);
nand U9603 (N_9603,N_8666,N_8481);
and U9604 (N_9604,N_8870,N_7904);
or U9605 (N_9605,N_8078,N_8629);
nor U9606 (N_9606,N_8691,N_8994);
nand U9607 (N_9607,N_8833,N_7810);
or U9608 (N_9608,N_8711,N_7954);
xor U9609 (N_9609,N_7656,N_7622);
nand U9610 (N_9610,N_8318,N_8601);
or U9611 (N_9611,N_8709,N_7949);
xor U9612 (N_9612,N_8892,N_7802);
xor U9613 (N_9613,N_8593,N_7967);
nand U9614 (N_9614,N_8785,N_7969);
or U9615 (N_9615,N_8177,N_7807);
and U9616 (N_9616,N_7990,N_7750);
and U9617 (N_9617,N_7912,N_7554);
and U9618 (N_9618,N_8110,N_8371);
and U9619 (N_9619,N_8310,N_8766);
nor U9620 (N_9620,N_7632,N_8816);
nor U9621 (N_9621,N_8633,N_8508);
or U9622 (N_9622,N_7757,N_7769);
xnor U9623 (N_9623,N_8929,N_8575);
nand U9624 (N_9624,N_8850,N_8418);
nand U9625 (N_9625,N_7731,N_7608);
and U9626 (N_9626,N_8910,N_8011);
nand U9627 (N_9627,N_8241,N_7758);
nor U9628 (N_9628,N_8796,N_8664);
nor U9629 (N_9629,N_8111,N_7996);
nand U9630 (N_9630,N_8096,N_7946);
nand U9631 (N_9631,N_8731,N_8255);
xor U9632 (N_9632,N_7588,N_8615);
nand U9633 (N_9633,N_8276,N_8603);
and U9634 (N_9634,N_8153,N_7849);
nor U9635 (N_9635,N_8066,N_8515);
nand U9636 (N_9636,N_8381,N_7754);
and U9637 (N_9637,N_8057,N_8939);
or U9638 (N_9638,N_8937,N_8207);
nor U9639 (N_9639,N_8001,N_8899);
nand U9640 (N_9640,N_8436,N_8768);
nor U9641 (N_9641,N_8268,N_8407);
or U9642 (N_9642,N_7713,N_7512);
and U9643 (N_9643,N_8469,N_7505);
or U9644 (N_9644,N_8022,N_7938);
nand U9645 (N_9645,N_8058,N_8219);
and U9646 (N_9646,N_7630,N_8949);
nand U9647 (N_9647,N_7627,N_8196);
or U9648 (N_9648,N_8688,N_7963);
xor U9649 (N_9649,N_8319,N_7831);
xor U9650 (N_9650,N_8170,N_8952);
and U9651 (N_9651,N_8896,N_7773);
nand U9652 (N_9652,N_8172,N_8399);
xnor U9653 (N_9653,N_8214,N_8245);
nor U9654 (N_9654,N_8647,N_8144);
or U9655 (N_9655,N_8120,N_8052);
or U9656 (N_9656,N_8813,N_7778);
nand U9657 (N_9657,N_8888,N_8454);
xnor U9658 (N_9658,N_7740,N_8946);
and U9659 (N_9659,N_8588,N_8679);
or U9660 (N_9660,N_8607,N_8995);
xnor U9661 (N_9661,N_8395,N_8035);
nor U9662 (N_9662,N_8871,N_7987);
xnor U9663 (N_9663,N_7784,N_8820);
or U9664 (N_9664,N_7714,N_8034);
xor U9665 (N_9665,N_7974,N_7631);
nand U9666 (N_9666,N_8351,N_8750);
and U9667 (N_9667,N_8878,N_7710);
or U9668 (N_9668,N_7515,N_7760);
and U9669 (N_9669,N_8204,N_8260);
xnor U9670 (N_9670,N_7593,N_7970);
and U9671 (N_9671,N_8486,N_8912);
xor U9672 (N_9672,N_8039,N_7873);
nand U9673 (N_9673,N_8361,N_8302);
nor U9674 (N_9674,N_8292,N_8967);
nand U9675 (N_9675,N_7559,N_8582);
nor U9676 (N_9676,N_7928,N_8047);
nor U9677 (N_9677,N_8271,N_8250);
or U9678 (N_9678,N_8019,N_8129);
nand U9679 (N_9679,N_8239,N_8654);
nand U9680 (N_9680,N_7540,N_8800);
xor U9681 (N_9681,N_7935,N_8092);
xor U9682 (N_9682,N_8400,N_8786);
and U9683 (N_9683,N_8051,N_8517);
and U9684 (N_9684,N_8759,N_8143);
or U9685 (N_9685,N_8101,N_8354);
or U9686 (N_9686,N_8202,N_8940);
xnor U9687 (N_9687,N_8405,N_7736);
nand U9688 (N_9688,N_8388,N_8832);
and U9689 (N_9689,N_8161,N_8417);
or U9690 (N_9690,N_8728,N_8897);
or U9691 (N_9691,N_8165,N_7844);
and U9692 (N_9692,N_7745,N_7968);
nor U9693 (N_9693,N_8993,N_8787);
or U9694 (N_9694,N_8126,N_8273);
and U9695 (N_9695,N_7862,N_8889);
or U9696 (N_9696,N_8323,N_8355);
nand U9697 (N_9697,N_8433,N_7570);
xnor U9698 (N_9698,N_8359,N_7812);
or U9699 (N_9699,N_8874,N_7669);
and U9700 (N_9700,N_8217,N_8826);
nand U9701 (N_9701,N_8080,N_7708);
and U9702 (N_9702,N_8909,N_7940);
xor U9703 (N_9703,N_8579,N_8824);
or U9704 (N_9704,N_7706,N_8594);
or U9705 (N_9705,N_8363,N_8109);
or U9706 (N_9706,N_7764,N_8565);
nand U9707 (N_9707,N_8415,N_8119);
and U9708 (N_9708,N_8230,N_8924);
nor U9709 (N_9709,N_8916,N_8340);
and U9710 (N_9710,N_7592,N_8364);
or U9711 (N_9711,N_7511,N_8821);
and U9712 (N_9712,N_8487,N_8839);
nand U9713 (N_9713,N_8384,N_8112);
nand U9714 (N_9714,N_8913,N_8495);
or U9715 (N_9715,N_8846,N_7837);
nand U9716 (N_9716,N_7558,N_8050);
and U9717 (N_9717,N_7785,N_7797);
nand U9718 (N_9718,N_7973,N_8574);
nor U9719 (N_9719,N_8891,N_8938);
xor U9720 (N_9720,N_8544,N_7666);
xor U9721 (N_9721,N_8344,N_8942);
nor U9722 (N_9722,N_7711,N_7751);
and U9723 (N_9723,N_8181,N_8752);
xor U9724 (N_9724,N_8703,N_8587);
xor U9725 (N_9725,N_8193,N_8163);
nor U9726 (N_9726,N_7718,N_7899);
xnor U9727 (N_9727,N_8830,N_8251);
xnor U9728 (N_9728,N_7749,N_7660);
or U9729 (N_9729,N_7959,N_8686);
nor U9730 (N_9730,N_8446,N_8540);
and U9731 (N_9731,N_8511,N_8764);
nor U9732 (N_9732,N_7717,N_7861);
xor U9733 (N_9733,N_8862,N_8708);
nor U9734 (N_9734,N_8549,N_8173);
xnor U9735 (N_9735,N_7920,N_8577);
nand U9736 (N_9736,N_8466,N_8290);
and U9737 (N_9737,N_7580,N_8944);
nor U9738 (N_9738,N_8452,N_7621);
nand U9739 (N_9739,N_7798,N_8960);
or U9740 (N_9740,N_8337,N_7510);
nor U9741 (N_9741,N_8353,N_8919);
or U9742 (N_9742,N_8915,N_7909);
nor U9743 (N_9743,N_8475,N_7786);
xor U9744 (N_9744,N_8836,N_8987);
xnor U9745 (N_9745,N_8055,N_8148);
nor U9746 (N_9746,N_8552,N_8660);
or U9747 (N_9747,N_7817,N_7746);
nand U9748 (N_9748,N_8716,N_8427);
and U9749 (N_9749,N_8722,N_7888);
or U9750 (N_9750,N_8636,N_8059);
nand U9751 (N_9751,N_7877,N_7624);
nor U9752 (N_9752,N_8959,N_8728);
and U9753 (N_9753,N_7873,N_8282);
and U9754 (N_9754,N_7878,N_7807);
and U9755 (N_9755,N_8852,N_8030);
or U9756 (N_9756,N_8781,N_8218);
or U9757 (N_9757,N_7505,N_8249);
nor U9758 (N_9758,N_7666,N_7512);
and U9759 (N_9759,N_8268,N_8526);
xnor U9760 (N_9760,N_8382,N_7760);
and U9761 (N_9761,N_8164,N_8671);
xnor U9762 (N_9762,N_8674,N_7939);
nor U9763 (N_9763,N_8969,N_8255);
or U9764 (N_9764,N_8276,N_8604);
nor U9765 (N_9765,N_8071,N_8126);
nand U9766 (N_9766,N_8895,N_7541);
and U9767 (N_9767,N_8299,N_7676);
nand U9768 (N_9768,N_7623,N_8717);
nor U9769 (N_9769,N_8758,N_8569);
nand U9770 (N_9770,N_8614,N_8994);
or U9771 (N_9771,N_8762,N_8591);
or U9772 (N_9772,N_8234,N_8934);
xor U9773 (N_9773,N_8576,N_8388);
nor U9774 (N_9774,N_7950,N_8255);
or U9775 (N_9775,N_8493,N_7947);
xor U9776 (N_9776,N_7760,N_8334);
xnor U9777 (N_9777,N_8365,N_8419);
or U9778 (N_9778,N_8664,N_8625);
nand U9779 (N_9779,N_8173,N_8032);
xor U9780 (N_9780,N_8679,N_7558);
or U9781 (N_9781,N_8330,N_8779);
or U9782 (N_9782,N_8484,N_7508);
xnor U9783 (N_9783,N_7861,N_8739);
nor U9784 (N_9784,N_8067,N_8615);
or U9785 (N_9785,N_8308,N_8212);
nand U9786 (N_9786,N_8808,N_7643);
nand U9787 (N_9787,N_8925,N_7899);
nand U9788 (N_9788,N_8833,N_8836);
or U9789 (N_9789,N_8971,N_8804);
nor U9790 (N_9790,N_8784,N_7613);
nand U9791 (N_9791,N_8582,N_7671);
and U9792 (N_9792,N_7700,N_8955);
nand U9793 (N_9793,N_8682,N_8884);
or U9794 (N_9794,N_7590,N_8478);
or U9795 (N_9795,N_7622,N_8387);
or U9796 (N_9796,N_8499,N_8745);
and U9797 (N_9797,N_7578,N_8133);
nor U9798 (N_9798,N_8619,N_8089);
and U9799 (N_9799,N_8831,N_8102);
nor U9800 (N_9800,N_7969,N_8791);
nor U9801 (N_9801,N_8312,N_8996);
nor U9802 (N_9802,N_8303,N_8595);
xnor U9803 (N_9803,N_7950,N_8443);
xnor U9804 (N_9804,N_7972,N_8197);
nand U9805 (N_9805,N_8548,N_8273);
nor U9806 (N_9806,N_7770,N_8581);
xor U9807 (N_9807,N_8978,N_7671);
or U9808 (N_9808,N_8296,N_8535);
nand U9809 (N_9809,N_8077,N_8061);
or U9810 (N_9810,N_7553,N_8064);
nand U9811 (N_9811,N_8021,N_7995);
xnor U9812 (N_9812,N_8618,N_7782);
xor U9813 (N_9813,N_8192,N_7760);
nand U9814 (N_9814,N_8968,N_7942);
nand U9815 (N_9815,N_7731,N_8215);
or U9816 (N_9816,N_8786,N_8762);
or U9817 (N_9817,N_8329,N_8875);
or U9818 (N_9818,N_8846,N_8476);
nor U9819 (N_9819,N_7867,N_8662);
xor U9820 (N_9820,N_8348,N_7801);
and U9821 (N_9821,N_8570,N_8508);
xor U9822 (N_9822,N_8761,N_7930);
and U9823 (N_9823,N_8692,N_8241);
and U9824 (N_9824,N_8899,N_7513);
and U9825 (N_9825,N_7593,N_7756);
or U9826 (N_9826,N_8356,N_8650);
nor U9827 (N_9827,N_7984,N_8091);
or U9828 (N_9828,N_8386,N_8223);
and U9829 (N_9829,N_8701,N_7599);
xnor U9830 (N_9830,N_8203,N_7994);
xnor U9831 (N_9831,N_7902,N_7717);
nand U9832 (N_9832,N_8207,N_7853);
nand U9833 (N_9833,N_8964,N_7795);
or U9834 (N_9834,N_7685,N_7609);
nand U9835 (N_9835,N_8197,N_7887);
or U9836 (N_9836,N_7859,N_7940);
and U9837 (N_9837,N_8733,N_8091);
nand U9838 (N_9838,N_8104,N_8051);
or U9839 (N_9839,N_7549,N_7681);
xor U9840 (N_9840,N_8026,N_8204);
or U9841 (N_9841,N_7838,N_8327);
nor U9842 (N_9842,N_7502,N_7671);
nand U9843 (N_9843,N_7531,N_8201);
or U9844 (N_9844,N_8722,N_8940);
nand U9845 (N_9845,N_8059,N_8776);
nand U9846 (N_9846,N_8774,N_8561);
or U9847 (N_9847,N_8413,N_8907);
nand U9848 (N_9848,N_7740,N_7877);
nor U9849 (N_9849,N_7638,N_8931);
and U9850 (N_9850,N_7568,N_7856);
nor U9851 (N_9851,N_8098,N_7673);
xnor U9852 (N_9852,N_8406,N_8660);
nand U9853 (N_9853,N_8804,N_8826);
nor U9854 (N_9854,N_8014,N_8512);
nor U9855 (N_9855,N_8603,N_8279);
and U9856 (N_9856,N_8827,N_8987);
xor U9857 (N_9857,N_8921,N_8978);
nand U9858 (N_9858,N_7749,N_8526);
nor U9859 (N_9859,N_8694,N_7806);
xor U9860 (N_9860,N_8462,N_8203);
and U9861 (N_9861,N_7770,N_8288);
nand U9862 (N_9862,N_7951,N_8157);
xor U9863 (N_9863,N_7748,N_7899);
or U9864 (N_9864,N_7787,N_7979);
nand U9865 (N_9865,N_7948,N_8713);
xnor U9866 (N_9866,N_7920,N_8490);
nand U9867 (N_9867,N_7839,N_7821);
or U9868 (N_9868,N_8559,N_8767);
nand U9869 (N_9869,N_8820,N_7815);
and U9870 (N_9870,N_8707,N_7780);
and U9871 (N_9871,N_8716,N_7852);
xnor U9872 (N_9872,N_8953,N_8598);
and U9873 (N_9873,N_8765,N_7653);
and U9874 (N_9874,N_8056,N_8514);
nand U9875 (N_9875,N_8895,N_7735);
nor U9876 (N_9876,N_7541,N_8317);
or U9877 (N_9877,N_8385,N_7522);
nor U9878 (N_9878,N_8769,N_8849);
and U9879 (N_9879,N_8449,N_8660);
nor U9880 (N_9880,N_8729,N_8677);
nor U9881 (N_9881,N_8613,N_8522);
nand U9882 (N_9882,N_7564,N_8242);
nand U9883 (N_9883,N_7787,N_7701);
xor U9884 (N_9884,N_8718,N_8490);
or U9885 (N_9885,N_7630,N_8300);
nand U9886 (N_9886,N_8997,N_8011);
nor U9887 (N_9887,N_7922,N_8978);
nor U9888 (N_9888,N_7769,N_8484);
nand U9889 (N_9889,N_7729,N_8526);
and U9890 (N_9890,N_8932,N_7879);
nor U9891 (N_9891,N_8785,N_7884);
or U9892 (N_9892,N_8047,N_7835);
and U9893 (N_9893,N_8091,N_7658);
and U9894 (N_9894,N_8258,N_8007);
or U9895 (N_9895,N_8272,N_8727);
and U9896 (N_9896,N_8339,N_8395);
and U9897 (N_9897,N_8806,N_8484);
nand U9898 (N_9898,N_7967,N_8897);
nor U9899 (N_9899,N_8452,N_7911);
or U9900 (N_9900,N_7939,N_8784);
and U9901 (N_9901,N_8897,N_7634);
and U9902 (N_9902,N_7626,N_8851);
nor U9903 (N_9903,N_7830,N_8390);
nor U9904 (N_9904,N_8838,N_7982);
or U9905 (N_9905,N_8558,N_8060);
xor U9906 (N_9906,N_7540,N_7723);
xor U9907 (N_9907,N_8595,N_8837);
xor U9908 (N_9908,N_7913,N_8384);
and U9909 (N_9909,N_8062,N_8607);
or U9910 (N_9910,N_7754,N_8227);
nor U9911 (N_9911,N_8367,N_8130);
or U9912 (N_9912,N_8621,N_8804);
or U9913 (N_9913,N_8986,N_7740);
nand U9914 (N_9914,N_7707,N_8539);
nor U9915 (N_9915,N_7582,N_8969);
xnor U9916 (N_9916,N_8766,N_8980);
xnor U9917 (N_9917,N_8236,N_7663);
and U9918 (N_9918,N_8372,N_8545);
or U9919 (N_9919,N_7831,N_7795);
xor U9920 (N_9920,N_7979,N_7801);
and U9921 (N_9921,N_8389,N_7872);
or U9922 (N_9922,N_7626,N_8882);
xnor U9923 (N_9923,N_8233,N_7820);
nor U9924 (N_9924,N_8646,N_8588);
and U9925 (N_9925,N_8869,N_8591);
nand U9926 (N_9926,N_8449,N_8718);
and U9927 (N_9927,N_8464,N_7902);
nor U9928 (N_9928,N_8467,N_8774);
or U9929 (N_9929,N_7928,N_7692);
and U9930 (N_9930,N_7676,N_8305);
or U9931 (N_9931,N_8264,N_8539);
xnor U9932 (N_9932,N_8335,N_7818);
and U9933 (N_9933,N_7740,N_7501);
or U9934 (N_9934,N_7616,N_8879);
xnor U9935 (N_9935,N_8635,N_7882);
nor U9936 (N_9936,N_7949,N_8369);
and U9937 (N_9937,N_7835,N_7970);
xnor U9938 (N_9938,N_8676,N_7660);
nor U9939 (N_9939,N_8338,N_8358);
nand U9940 (N_9940,N_7682,N_7976);
and U9941 (N_9941,N_8263,N_8063);
xnor U9942 (N_9942,N_8733,N_7996);
and U9943 (N_9943,N_8902,N_8841);
or U9944 (N_9944,N_7742,N_7659);
and U9945 (N_9945,N_8116,N_7669);
and U9946 (N_9946,N_8582,N_7831);
xor U9947 (N_9947,N_8499,N_8477);
or U9948 (N_9948,N_8194,N_8207);
and U9949 (N_9949,N_7572,N_7729);
or U9950 (N_9950,N_8784,N_8070);
xor U9951 (N_9951,N_8173,N_7669);
or U9952 (N_9952,N_7507,N_8302);
or U9953 (N_9953,N_8160,N_8168);
nor U9954 (N_9954,N_8742,N_8122);
nand U9955 (N_9955,N_8479,N_8624);
or U9956 (N_9956,N_7998,N_8610);
nand U9957 (N_9957,N_8503,N_8565);
or U9958 (N_9958,N_7972,N_7763);
xor U9959 (N_9959,N_7598,N_8203);
and U9960 (N_9960,N_8252,N_8144);
nand U9961 (N_9961,N_7710,N_8748);
nor U9962 (N_9962,N_8876,N_8988);
and U9963 (N_9963,N_7573,N_8466);
nor U9964 (N_9964,N_8422,N_8291);
or U9965 (N_9965,N_8237,N_8456);
nand U9966 (N_9966,N_8455,N_7795);
nor U9967 (N_9967,N_8969,N_8069);
nand U9968 (N_9968,N_8316,N_8939);
nor U9969 (N_9969,N_7879,N_8362);
or U9970 (N_9970,N_8324,N_8785);
xor U9971 (N_9971,N_7522,N_8915);
and U9972 (N_9972,N_8056,N_8345);
or U9973 (N_9973,N_8348,N_7641);
nand U9974 (N_9974,N_8846,N_8857);
and U9975 (N_9975,N_7681,N_8284);
xor U9976 (N_9976,N_8398,N_8325);
nor U9977 (N_9977,N_7953,N_8807);
nand U9978 (N_9978,N_8854,N_7741);
nand U9979 (N_9979,N_8099,N_7692);
nand U9980 (N_9980,N_8224,N_8899);
xor U9981 (N_9981,N_7515,N_8330);
or U9982 (N_9982,N_8473,N_7684);
nand U9983 (N_9983,N_8676,N_8295);
nand U9984 (N_9984,N_8805,N_7648);
nand U9985 (N_9985,N_8803,N_8437);
or U9986 (N_9986,N_7949,N_7943);
nand U9987 (N_9987,N_7584,N_8726);
nand U9988 (N_9988,N_8463,N_8569);
and U9989 (N_9989,N_7624,N_8932);
or U9990 (N_9990,N_7583,N_7679);
nor U9991 (N_9991,N_8748,N_7896);
xnor U9992 (N_9992,N_8063,N_7684);
xor U9993 (N_9993,N_7781,N_8157);
nand U9994 (N_9994,N_7539,N_8624);
xnor U9995 (N_9995,N_7782,N_7902);
xnor U9996 (N_9996,N_7575,N_8001);
nor U9997 (N_9997,N_8378,N_8357);
nand U9998 (N_9998,N_7785,N_7692);
nand U9999 (N_9999,N_8827,N_7942);
or U10000 (N_10000,N_8103,N_8096);
and U10001 (N_10001,N_8485,N_8365);
or U10002 (N_10002,N_8675,N_8575);
nor U10003 (N_10003,N_8427,N_8816);
or U10004 (N_10004,N_8194,N_8133);
or U10005 (N_10005,N_7584,N_8283);
nand U10006 (N_10006,N_7828,N_7731);
nand U10007 (N_10007,N_7597,N_8770);
xor U10008 (N_10008,N_8982,N_8270);
xnor U10009 (N_10009,N_8338,N_7734);
or U10010 (N_10010,N_8738,N_8132);
or U10011 (N_10011,N_8319,N_8847);
or U10012 (N_10012,N_7955,N_7500);
nor U10013 (N_10013,N_8633,N_8515);
xor U10014 (N_10014,N_7959,N_8100);
and U10015 (N_10015,N_7732,N_8986);
nor U10016 (N_10016,N_8273,N_8681);
and U10017 (N_10017,N_8373,N_8154);
nor U10018 (N_10018,N_8885,N_8471);
or U10019 (N_10019,N_8314,N_7995);
xnor U10020 (N_10020,N_7709,N_7740);
nor U10021 (N_10021,N_7522,N_8898);
nand U10022 (N_10022,N_8605,N_7807);
nor U10023 (N_10023,N_8000,N_8694);
or U10024 (N_10024,N_8292,N_7792);
or U10025 (N_10025,N_8994,N_8492);
xnor U10026 (N_10026,N_7666,N_7587);
nor U10027 (N_10027,N_8893,N_8366);
xnor U10028 (N_10028,N_8711,N_8061);
nor U10029 (N_10029,N_7581,N_7667);
nor U10030 (N_10030,N_7546,N_7541);
or U10031 (N_10031,N_7867,N_7558);
or U10032 (N_10032,N_8573,N_7693);
nand U10033 (N_10033,N_8722,N_8647);
or U10034 (N_10034,N_7999,N_8804);
xnor U10035 (N_10035,N_8849,N_8273);
or U10036 (N_10036,N_7564,N_7904);
nor U10037 (N_10037,N_8685,N_8974);
nand U10038 (N_10038,N_7540,N_7794);
nand U10039 (N_10039,N_7712,N_8075);
and U10040 (N_10040,N_8773,N_8846);
nand U10041 (N_10041,N_8587,N_8129);
and U10042 (N_10042,N_7734,N_7543);
xor U10043 (N_10043,N_8743,N_8572);
or U10044 (N_10044,N_8518,N_7605);
or U10045 (N_10045,N_8629,N_8374);
nor U10046 (N_10046,N_8913,N_8674);
xnor U10047 (N_10047,N_8502,N_8695);
xnor U10048 (N_10048,N_8556,N_8482);
and U10049 (N_10049,N_8619,N_8122);
and U10050 (N_10050,N_7654,N_8002);
xnor U10051 (N_10051,N_8112,N_7881);
xor U10052 (N_10052,N_7546,N_8772);
nand U10053 (N_10053,N_8404,N_7581);
xnor U10054 (N_10054,N_7612,N_8227);
nor U10055 (N_10055,N_8295,N_7751);
or U10056 (N_10056,N_8857,N_8690);
nor U10057 (N_10057,N_8832,N_7795);
and U10058 (N_10058,N_7518,N_8587);
and U10059 (N_10059,N_7851,N_8998);
nor U10060 (N_10060,N_8673,N_8334);
xor U10061 (N_10061,N_7699,N_8410);
and U10062 (N_10062,N_7874,N_7569);
or U10063 (N_10063,N_8942,N_7595);
nor U10064 (N_10064,N_8083,N_8500);
nand U10065 (N_10065,N_7772,N_8953);
and U10066 (N_10066,N_7544,N_7981);
xnor U10067 (N_10067,N_8109,N_7548);
nor U10068 (N_10068,N_8907,N_8025);
xnor U10069 (N_10069,N_7655,N_8209);
and U10070 (N_10070,N_7793,N_7843);
nand U10071 (N_10071,N_7631,N_7756);
nor U10072 (N_10072,N_8386,N_7570);
nand U10073 (N_10073,N_8092,N_7862);
xor U10074 (N_10074,N_8994,N_8211);
nand U10075 (N_10075,N_7907,N_8685);
or U10076 (N_10076,N_8250,N_7891);
nand U10077 (N_10077,N_8834,N_8405);
and U10078 (N_10078,N_7620,N_8145);
nor U10079 (N_10079,N_7882,N_7742);
nand U10080 (N_10080,N_8088,N_7827);
nor U10081 (N_10081,N_7887,N_8765);
and U10082 (N_10082,N_8531,N_7817);
nor U10083 (N_10083,N_7632,N_8453);
xor U10084 (N_10084,N_8376,N_8698);
nand U10085 (N_10085,N_8413,N_8924);
xnor U10086 (N_10086,N_7603,N_8177);
nor U10087 (N_10087,N_8257,N_8478);
xor U10088 (N_10088,N_8875,N_8191);
nand U10089 (N_10089,N_8322,N_8871);
xor U10090 (N_10090,N_8723,N_7933);
nand U10091 (N_10091,N_7879,N_7773);
nor U10092 (N_10092,N_7557,N_7534);
xnor U10093 (N_10093,N_8896,N_8565);
nor U10094 (N_10094,N_8137,N_8559);
nor U10095 (N_10095,N_7530,N_8131);
nand U10096 (N_10096,N_7545,N_7767);
xnor U10097 (N_10097,N_8746,N_8700);
nand U10098 (N_10098,N_8394,N_7923);
and U10099 (N_10099,N_8568,N_7503);
and U10100 (N_10100,N_8208,N_8856);
nand U10101 (N_10101,N_8188,N_8529);
nor U10102 (N_10102,N_8425,N_7720);
and U10103 (N_10103,N_7619,N_8979);
nand U10104 (N_10104,N_7677,N_8040);
or U10105 (N_10105,N_7630,N_7762);
and U10106 (N_10106,N_8133,N_8303);
or U10107 (N_10107,N_7786,N_7920);
nand U10108 (N_10108,N_8522,N_8309);
nor U10109 (N_10109,N_8768,N_7699);
nor U10110 (N_10110,N_7805,N_7581);
and U10111 (N_10111,N_7637,N_7824);
xnor U10112 (N_10112,N_8895,N_8268);
or U10113 (N_10113,N_7786,N_8865);
xor U10114 (N_10114,N_7840,N_8133);
and U10115 (N_10115,N_8864,N_8268);
nand U10116 (N_10116,N_8485,N_8507);
nor U10117 (N_10117,N_7964,N_8520);
or U10118 (N_10118,N_8572,N_8477);
nor U10119 (N_10119,N_7894,N_8876);
or U10120 (N_10120,N_8859,N_8755);
xor U10121 (N_10121,N_8001,N_7556);
and U10122 (N_10122,N_7997,N_8543);
nor U10123 (N_10123,N_7807,N_8321);
nand U10124 (N_10124,N_8742,N_8126);
xnor U10125 (N_10125,N_8697,N_8823);
xnor U10126 (N_10126,N_8268,N_8393);
and U10127 (N_10127,N_8482,N_8731);
nand U10128 (N_10128,N_7554,N_8505);
xnor U10129 (N_10129,N_7590,N_7724);
nand U10130 (N_10130,N_8611,N_7663);
nand U10131 (N_10131,N_7528,N_8392);
or U10132 (N_10132,N_8908,N_8096);
or U10133 (N_10133,N_7679,N_8958);
and U10134 (N_10134,N_8333,N_8498);
nand U10135 (N_10135,N_7594,N_7525);
xnor U10136 (N_10136,N_7658,N_8204);
nor U10137 (N_10137,N_8927,N_8728);
nor U10138 (N_10138,N_7963,N_8397);
xnor U10139 (N_10139,N_7634,N_7647);
nor U10140 (N_10140,N_8801,N_7780);
or U10141 (N_10141,N_7773,N_8002);
nand U10142 (N_10142,N_7877,N_8271);
and U10143 (N_10143,N_7930,N_8722);
xnor U10144 (N_10144,N_8570,N_8176);
nor U10145 (N_10145,N_8760,N_7607);
or U10146 (N_10146,N_8172,N_8046);
or U10147 (N_10147,N_7719,N_7606);
xor U10148 (N_10148,N_8876,N_8539);
nor U10149 (N_10149,N_7941,N_8779);
and U10150 (N_10150,N_8337,N_8935);
and U10151 (N_10151,N_7984,N_8877);
or U10152 (N_10152,N_7744,N_7699);
and U10153 (N_10153,N_7853,N_8927);
nor U10154 (N_10154,N_7608,N_7510);
and U10155 (N_10155,N_7943,N_7805);
xor U10156 (N_10156,N_7556,N_8019);
or U10157 (N_10157,N_8793,N_8145);
xor U10158 (N_10158,N_8751,N_8566);
nor U10159 (N_10159,N_8764,N_8123);
xor U10160 (N_10160,N_7862,N_8308);
xor U10161 (N_10161,N_8665,N_7878);
xor U10162 (N_10162,N_7984,N_8488);
nor U10163 (N_10163,N_7792,N_8983);
nand U10164 (N_10164,N_8764,N_8021);
xor U10165 (N_10165,N_7526,N_7980);
nor U10166 (N_10166,N_7672,N_8128);
xor U10167 (N_10167,N_7551,N_8902);
xnor U10168 (N_10168,N_8346,N_8769);
xnor U10169 (N_10169,N_8339,N_8216);
or U10170 (N_10170,N_7699,N_7929);
nand U10171 (N_10171,N_8772,N_8320);
and U10172 (N_10172,N_8431,N_7605);
xnor U10173 (N_10173,N_7905,N_8777);
nand U10174 (N_10174,N_7670,N_7625);
xor U10175 (N_10175,N_7864,N_7939);
or U10176 (N_10176,N_7515,N_8056);
and U10177 (N_10177,N_7876,N_8993);
nor U10178 (N_10178,N_7527,N_8021);
nor U10179 (N_10179,N_8196,N_8211);
nand U10180 (N_10180,N_8611,N_8686);
xnor U10181 (N_10181,N_7766,N_8019);
nand U10182 (N_10182,N_8819,N_8667);
or U10183 (N_10183,N_8052,N_7738);
or U10184 (N_10184,N_7818,N_7616);
nand U10185 (N_10185,N_8550,N_8318);
or U10186 (N_10186,N_8372,N_7913);
xnor U10187 (N_10187,N_8798,N_8175);
or U10188 (N_10188,N_8890,N_8739);
xor U10189 (N_10189,N_7997,N_8503);
xor U10190 (N_10190,N_8644,N_8181);
nand U10191 (N_10191,N_8180,N_8784);
nor U10192 (N_10192,N_7903,N_8754);
and U10193 (N_10193,N_8059,N_8632);
nand U10194 (N_10194,N_8843,N_8453);
or U10195 (N_10195,N_8662,N_8108);
nand U10196 (N_10196,N_8881,N_7526);
or U10197 (N_10197,N_7782,N_8070);
nor U10198 (N_10198,N_7533,N_8423);
and U10199 (N_10199,N_7780,N_7544);
xnor U10200 (N_10200,N_8327,N_8151);
xor U10201 (N_10201,N_8945,N_8104);
xor U10202 (N_10202,N_7665,N_8391);
or U10203 (N_10203,N_7812,N_7793);
xor U10204 (N_10204,N_8327,N_7752);
nand U10205 (N_10205,N_8771,N_7957);
nand U10206 (N_10206,N_8397,N_8698);
and U10207 (N_10207,N_8619,N_8016);
or U10208 (N_10208,N_8619,N_8686);
nand U10209 (N_10209,N_8525,N_7999);
xnor U10210 (N_10210,N_7912,N_8434);
and U10211 (N_10211,N_8878,N_8900);
and U10212 (N_10212,N_8306,N_8779);
xnor U10213 (N_10213,N_7541,N_7689);
and U10214 (N_10214,N_8160,N_8827);
xor U10215 (N_10215,N_8616,N_8796);
xnor U10216 (N_10216,N_8889,N_8437);
and U10217 (N_10217,N_8414,N_8088);
nand U10218 (N_10218,N_8184,N_8066);
or U10219 (N_10219,N_7835,N_8516);
xor U10220 (N_10220,N_7677,N_7908);
xnor U10221 (N_10221,N_8372,N_8176);
nand U10222 (N_10222,N_8878,N_8604);
nor U10223 (N_10223,N_8908,N_8036);
nor U10224 (N_10224,N_8745,N_8041);
xor U10225 (N_10225,N_7657,N_8488);
xnor U10226 (N_10226,N_8396,N_7501);
nand U10227 (N_10227,N_7870,N_8784);
and U10228 (N_10228,N_8452,N_8172);
nand U10229 (N_10229,N_8959,N_8422);
nor U10230 (N_10230,N_8395,N_7773);
or U10231 (N_10231,N_8946,N_7523);
nand U10232 (N_10232,N_8430,N_8542);
and U10233 (N_10233,N_8226,N_8445);
and U10234 (N_10234,N_7518,N_8584);
nand U10235 (N_10235,N_8577,N_8482);
or U10236 (N_10236,N_7726,N_7876);
nand U10237 (N_10237,N_8663,N_7509);
or U10238 (N_10238,N_8952,N_8846);
nand U10239 (N_10239,N_8208,N_8620);
and U10240 (N_10240,N_7936,N_7560);
xor U10241 (N_10241,N_8725,N_8794);
xor U10242 (N_10242,N_7904,N_8143);
and U10243 (N_10243,N_7679,N_8988);
or U10244 (N_10244,N_7515,N_7832);
nor U10245 (N_10245,N_7590,N_8891);
and U10246 (N_10246,N_8922,N_7503);
or U10247 (N_10247,N_7905,N_8086);
xnor U10248 (N_10248,N_7854,N_8946);
xor U10249 (N_10249,N_7583,N_8633);
xnor U10250 (N_10250,N_7977,N_7840);
and U10251 (N_10251,N_7877,N_7656);
or U10252 (N_10252,N_8552,N_7570);
and U10253 (N_10253,N_8008,N_8617);
xor U10254 (N_10254,N_8720,N_8801);
nand U10255 (N_10255,N_7636,N_8184);
and U10256 (N_10256,N_7917,N_7522);
or U10257 (N_10257,N_8328,N_8782);
nor U10258 (N_10258,N_8266,N_8127);
and U10259 (N_10259,N_8093,N_8316);
nand U10260 (N_10260,N_7727,N_7686);
xnor U10261 (N_10261,N_8384,N_7611);
xnor U10262 (N_10262,N_7758,N_8695);
or U10263 (N_10263,N_8299,N_7513);
nor U10264 (N_10264,N_8779,N_8556);
nor U10265 (N_10265,N_8486,N_8938);
nor U10266 (N_10266,N_8309,N_8471);
or U10267 (N_10267,N_7611,N_7823);
xor U10268 (N_10268,N_8116,N_7704);
or U10269 (N_10269,N_8832,N_8024);
xor U10270 (N_10270,N_8007,N_8748);
and U10271 (N_10271,N_7708,N_8194);
or U10272 (N_10272,N_8120,N_8197);
and U10273 (N_10273,N_7625,N_8698);
xor U10274 (N_10274,N_8594,N_7872);
nand U10275 (N_10275,N_8173,N_8246);
or U10276 (N_10276,N_8028,N_8385);
xor U10277 (N_10277,N_8608,N_8331);
nor U10278 (N_10278,N_8889,N_8285);
nor U10279 (N_10279,N_8598,N_8778);
nor U10280 (N_10280,N_7534,N_8175);
nor U10281 (N_10281,N_7917,N_7571);
and U10282 (N_10282,N_8648,N_8711);
xnor U10283 (N_10283,N_7574,N_8310);
and U10284 (N_10284,N_8928,N_8291);
and U10285 (N_10285,N_7627,N_8025);
and U10286 (N_10286,N_8064,N_7652);
nand U10287 (N_10287,N_8257,N_8743);
xor U10288 (N_10288,N_7576,N_8669);
and U10289 (N_10289,N_8274,N_7508);
or U10290 (N_10290,N_7648,N_8562);
nor U10291 (N_10291,N_7939,N_8459);
xnor U10292 (N_10292,N_7755,N_8711);
nand U10293 (N_10293,N_8869,N_7525);
xor U10294 (N_10294,N_8605,N_7764);
nand U10295 (N_10295,N_8013,N_7782);
xor U10296 (N_10296,N_7591,N_8359);
nand U10297 (N_10297,N_8835,N_8929);
or U10298 (N_10298,N_8066,N_7524);
nand U10299 (N_10299,N_8823,N_8598);
or U10300 (N_10300,N_7963,N_8098);
nor U10301 (N_10301,N_8347,N_8035);
xor U10302 (N_10302,N_7569,N_7713);
nand U10303 (N_10303,N_8891,N_7578);
or U10304 (N_10304,N_8265,N_8734);
xor U10305 (N_10305,N_7873,N_8128);
xor U10306 (N_10306,N_7962,N_7883);
nor U10307 (N_10307,N_7536,N_8098);
or U10308 (N_10308,N_7975,N_8707);
or U10309 (N_10309,N_8934,N_8750);
nand U10310 (N_10310,N_8309,N_8489);
and U10311 (N_10311,N_8505,N_8973);
nand U10312 (N_10312,N_8465,N_7684);
nand U10313 (N_10313,N_8744,N_8425);
or U10314 (N_10314,N_7737,N_8854);
nor U10315 (N_10315,N_8249,N_8078);
nand U10316 (N_10316,N_8221,N_8406);
nor U10317 (N_10317,N_7740,N_7959);
nor U10318 (N_10318,N_8573,N_7947);
nor U10319 (N_10319,N_8641,N_8735);
or U10320 (N_10320,N_8290,N_8552);
xor U10321 (N_10321,N_7555,N_8566);
or U10322 (N_10322,N_8204,N_8550);
nor U10323 (N_10323,N_7542,N_7528);
xnor U10324 (N_10324,N_8744,N_8702);
nand U10325 (N_10325,N_7614,N_7690);
or U10326 (N_10326,N_7684,N_8742);
nand U10327 (N_10327,N_8278,N_8828);
or U10328 (N_10328,N_8971,N_8459);
xnor U10329 (N_10329,N_7620,N_8766);
and U10330 (N_10330,N_8813,N_8270);
and U10331 (N_10331,N_8239,N_8051);
and U10332 (N_10332,N_8373,N_7901);
and U10333 (N_10333,N_8376,N_8783);
or U10334 (N_10334,N_8828,N_7789);
and U10335 (N_10335,N_8291,N_8344);
xnor U10336 (N_10336,N_8330,N_8160);
or U10337 (N_10337,N_8350,N_8727);
nand U10338 (N_10338,N_8612,N_8327);
nand U10339 (N_10339,N_8142,N_7876);
or U10340 (N_10340,N_7950,N_7796);
xor U10341 (N_10341,N_7756,N_8525);
nand U10342 (N_10342,N_8474,N_8850);
nor U10343 (N_10343,N_8904,N_7665);
and U10344 (N_10344,N_8237,N_8024);
nand U10345 (N_10345,N_8749,N_7866);
xnor U10346 (N_10346,N_7970,N_7752);
nor U10347 (N_10347,N_7825,N_8650);
nand U10348 (N_10348,N_7518,N_7546);
and U10349 (N_10349,N_8570,N_7891);
xor U10350 (N_10350,N_7852,N_8797);
and U10351 (N_10351,N_8547,N_8686);
and U10352 (N_10352,N_8586,N_8545);
and U10353 (N_10353,N_8674,N_8836);
or U10354 (N_10354,N_7842,N_8288);
nor U10355 (N_10355,N_8290,N_8541);
xor U10356 (N_10356,N_8211,N_8453);
xor U10357 (N_10357,N_8409,N_8249);
xnor U10358 (N_10358,N_8289,N_7666);
nand U10359 (N_10359,N_7738,N_7521);
or U10360 (N_10360,N_7758,N_8736);
nor U10361 (N_10361,N_7859,N_8715);
nand U10362 (N_10362,N_8011,N_8666);
nand U10363 (N_10363,N_7982,N_8195);
or U10364 (N_10364,N_8342,N_8160);
xnor U10365 (N_10365,N_8350,N_8604);
nand U10366 (N_10366,N_8400,N_7550);
nor U10367 (N_10367,N_8173,N_8383);
nor U10368 (N_10368,N_8994,N_8831);
or U10369 (N_10369,N_7930,N_8401);
xor U10370 (N_10370,N_8184,N_8693);
and U10371 (N_10371,N_8488,N_8762);
nor U10372 (N_10372,N_8545,N_8734);
nand U10373 (N_10373,N_8777,N_7704);
nor U10374 (N_10374,N_7948,N_7621);
nand U10375 (N_10375,N_8193,N_8322);
xor U10376 (N_10376,N_8837,N_7649);
nor U10377 (N_10377,N_8515,N_8808);
nor U10378 (N_10378,N_7736,N_8519);
nand U10379 (N_10379,N_8642,N_8735);
or U10380 (N_10380,N_8955,N_8725);
or U10381 (N_10381,N_8276,N_8262);
nand U10382 (N_10382,N_8607,N_8293);
xnor U10383 (N_10383,N_7753,N_7756);
and U10384 (N_10384,N_7861,N_8328);
and U10385 (N_10385,N_7798,N_7662);
nand U10386 (N_10386,N_8896,N_8062);
xor U10387 (N_10387,N_8365,N_8303);
and U10388 (N_10388,N_7717,N_8467);
nand U10389 (N_10389,N_7610,N_8903);
xnor U10390 (N_10390,N_8471,N_8092);
or U10391 (N_10391,N_7629,N_7972);
and U10392 (N_10392,N_7895,N_7638);
nand U10393 (N_10393,N_8718,N_7557);
nor U10394 (N_10394,N_7611,N_8993);
xor U10395 (N_10395,N_8028,N_7880);
or U10396 (N_10396,N_8661,N_8157);
xor U10397 (N_10397,N_8321,N_8884);
nor U10398 (N_10398,N_8884,N_8595);
nor U10399 (N_10399,N_8891,N_8342);
and U10400 (N_10400,N_7635,N_7538);
and U10401 (N_10401,N_8625,N_8698);
nand U10402 (N_10402,N_8316,N_7943);
nand U10403 (N_10403,N_7846,N_8672);
and U10404 (N_10404,N_7881,N_8880);
or U10405 (N_10405,N_7695,N_8406);
nand U10406 (N_10406,N_7905,N_8120);
xnor U10407 (N_10407,N_8576,N_7567);
nand U10408 (N_10408,N_8844,N_8033);
xor U10409 (N_10409,N_7602,N_8390);
xnor U10410 (N_10410,N_8145,N_8695);
xor U10411 (N_10411,N_7586,N_7767);
and U10412 (N_10412,N_8931,N_7858);
xnor U10413 (N_10413,N_8855,N_8607);
xnor U10414 (N_10414,N_8750,N_8860);
xor U10415 (N_10415,N_7531,N_8411);
or U10416 (N_10416,N_7538,N_8704);
or U10417 (N_10417,N_8345,N_8298);
or U10418 (N_10418,N_8245,N_7850);
nand U10419 (N_10419,N_7857,N_8020);
xnor U10420 (N_10420,N_8373,N_8094);
xnor U10421 (N_10421,N_7980,N_8451);
or U10422 (N_10422,N_8132,N_8923);
or U10423 (N_10423,N_7833,N_8772);
xnor U10424 (N_10424,N_8647,N_8616);
nor U10425 (N_10425,N_8828,N_8294);
nor U10426 (N_10426,N_8241,N_7700);
xnor U10427 (N_10427,N_8640,N_7690);
nor U10428 (N_10428,N_7939,N_8500);
or U10429 (N_10429,N_7773,N_8461);
and U10430 (N_10430,N_8281,N_8896);
and U10431 (N_10431,N_7737,N_8317);
xnor U10432 (N_10432,N_8500,N_8336);
or U10433 (N_10433,N_8475,N_8328);
or U10434 (N_10434,N_8117,N_8232);
and U10435 (N_10435,N_8069,N_7509);
or U10436 (N_10436,N_8437,N_7645);
or U10437 (N_10437,N_7640,N_8022);
or U10438 (N_10438,N_7822,N_8855);
nand U10439 (N_10439,N_7683,N_8104);
and U10440 (N_10440,N_7977,N_7782);
and U10441 (N_10441,N_7574,N_8524);
nand U10442 (N_10442,N_8333,N_8393);
nand U10443 (N_10443,N_8549,N_8432);
or U10444 (N_10444,N_7842,N_7568);
nor U10445 (N_10445,N_8252,N_7971);
or U10446 (N_10446,N_8861,N_7606);
nor U10447 (N_10447,N_7963,N_8987);
nand U10448 (N_10448,N_8211,N_8894);
or U10449 (N_10449,N_8698,N_8350);
or U10450 (N_10450,N_8324,N_8612);
nand U10451 (N_10451,N_8627,N_7766);
xor U10452 (N_10452,N_8478,N_7678);
or U10453 (N_10453,N_7708,N_8095);
and U10454 (N_10454,N_8879,N_8887);
or U10455 (N_10455,N_8646,N_8986);
nor U10456 (N_10456,N_7968,N_8869);
xnor U10457 (N_10457,N_8981,N_7548);
or U10458 (N_10458,N_8672,N_7665);
nor U10459 (N_10459,N_7554,N_8981);
or U10460 (N_10460,N_8753,N_8807);
xor U10461 (N_10461,N_8384,N_7795);
or U10462 (N_10462,N_8509,N_8673);
nand U10463 (N_10463,N_7623,N_7834);
xnor U10464 (N_10464,N_8320,N_7695);
and U10465 (N_10465,N_8510,N_7680);
or U10466 (N_10466,N_7929,N_8149);
or U10467 (N_10467,N_8320,N_7631);
nand U10468 (N_10468,N_8335,N_8944);
nor U10469 (N_10469,N_8684,N_8252);
nand U10470 (N_10470,N_7635,N_7599);
nand U10471 (N_10471,N_7789,N_8862);
nor U10472 (N_10472,N_7843,N_7673);
or U10473 (N_10473,N_8225,N_7926);
nand U10474 (N_10474,N_8761,N_8709);
xor U10475 (N_10475,N_8267,N_8297);
and U10476 (N_10476,N_7700,N_7519);
nand U10477 (N_10477,N_8864,N_8215);
or U10478 (N_10478,N_8087,N_7608);
xnor U10479 (N_10479,N_8755,N_7829);
nand U10480 (N_10480,N_7545,N_7937);
and U10481 (N_10481,N_8533,N_8412);
or U10482 (N_10482,N_7970,N_7637);
nor U10483 (N_10483,N_8474,N_8371);
nor U10484 (N_10484,N_7810,N_8750);
xor U10485 (N_10485,N_8263,N_7936);
xor U10486 (N_10486,N_8110,N_8672);
or U10487 (N_10487,N_8750,N_8444);
nand U10488 (N_10488,N_8395,N_8982);
nand U10489 (N_10489,N_8200,N_7886);
nand U10490 (N_10490,N_7809,N_7928);
or U10491 (N_10491,N_7738,N_8594);
nand U10492 (N_10492,N_8959,N_7878);
and U10493 (N_10493,N_8514,N_7959);
xnor U10494 (N_10494,N_8317,N_8183);
nor U10495 (N_10495,N_8928,N_8123);
nand U10496 (N_10496,N_7751,N_7652);
nand U10497 (N_10497,N_7549,N_8326);
xnor U10498 (N_10498,N_8195,N_8060);
and U10499 (N_10499,N_8252,N_8912);
nand U10500 (N_10500,N_9618,N_9507);
or U10501 (N_10501,N_9905,N_9551);
nor U10502 (N_10502,N_9265,N_10444);
xor U10503 (N_10503,N_9407,N_9620);
nor U10504 (N_10504,N_9302,N_10274);
xnor U10505 (N_10505,N_9818,N_10424);
and U10506 (N_10506,N_10165,N_9579);
and U10507 (N_10507,N_9002,N_9346);
and U10508 (N_10508,N_9648,N_9247);
nand U10509 (N_10509,N_9562,N_9695);
nor U10510 (N_10510,N_10351,N_10314);
nor U10511 (N_10511,N_10028,N_9372);
nor U10512 (N_10512,N_9864,N_9472);
nor U10513 (N_10513,N_9787,N_9667);
nand U10514 (N_10514,N_9324,N_9671);
nor U10515 (N_10515,N_9487,N_9808);
or U10516 (N_10516,N_9763,N_9884);
xnor U10517 (N_10517,N_9894,N_9570);
xor U10518 (N_10518,N_10061,N_9046);
xnor U10519 (N_10519,N_10139,N_10159);
nor U10520 (N_10520,N_10377,N_10022);
xor U10521 (N_10521,N_9747,N_9429);
nor U10522 (N_10522,N_9073,N_9779);
nand U10523 (N_10523,N_9781,N_9212);
and U10524 (N_10524,N_9499,N_9772);
and U10525 (N_10525,N_10386,N_9746);
or U10526 (N_10526,N_9843,N_9557);
or U10527 (N_10527,N_9035,N_10492);
nor U10528 (N_10528,N_9568,N_9368);
and U10529 (N_10529,N_10033,N_9099);
xor U10530 (N_10530,N_9660,N_9513);
nand U10531 (N_10531,N_10345,N_10258);
and U10532 (N_10532,N_9474,N_9928);
nor U10533 (N_10533,N_10035,N_9445);
nand U10534 (N_10534,N_10065,N_9872);
xor U10535 (N_10535,N_10462,N_9113);
nand U10536 (N_10536,N_10146,N_9389);
nand U10537 (N_10537,N_9801,N_9185);
nand U10538 (N_10538,N_10103,N_10114);
nor U10539 (N_10539,N_9900,N_9606);
nand U10540 (N_10540,N_10463,N_10242);
or U10541 (N_10541,N_10023,N_9912);
nand U10542 (N_10542,N_9491,N_9564);
nor U10543 (N_10543,N_9208,N_10153);
nand U10544 (N_10544,N_10355,N_9910);
nor U10545 (N_10545,N_9154,N_9956);
nor U10546 (N_10546,N_9799,N_10266);
xnor U10547 (N_10547,N_9626,N_9714);
nand U10548 (N_10548,N_10180,N_10064);
nor U10549 (N_10549,N_9304,N_9183);
or U10550 (N_10550,N_9005,N_9221);
nor U10551 (N_10551,N_9362,N_9042);
and U10552 (N_10552,N_9679,N_9641);
or U10553 (N_10553,N_9147,N_9462);
xor U10554 (N_10554,N_10095,N_9759);
and U10555 (N_10555,N_9531,N_10495);
nand U10556 (N_10556,N_10066,N_10145);
nor U10557 (N_10557,N_9446,N_9773);
nand U10558 (N_10558,N_9321,N_10332);
nor U10559 (N_10559,N_9088,N_9934);
xor U10560 (N_10560,N_9401,N_9502);
and U10561 (N_10561,N_9039,N_9837);
or U10562 (N_10562,N_10264,N_9343);
nand U10563 (N_10563,N_9254,N_9998);
xor U10564 (N_10564,N_10002,N_9397);
or U10565 (N_10565,N_9784,N_10447);
and U10566 (N_10566,N_10098,N_9237);
nand U10567 (N_10567,N_10236,N_9596);
and U10568 (N_10568,N_9096,N_10148);
and U10569 (N_10569,N_10372,N_9335);
nand U10570 (N_10570,N_9024,N_9790);
and U10571 (N_10571,N_9599,N_10392);
nor U10572 (N_10572,N_9358,N_10091);
or U10573 (N_10573,N_10164,N_9810);
nor U10574 (N_10574,N_9242,N_10073);
xor U10575 (N_10575,N_10341,N_10457);
or U10576 (N_10576,N_9535,N_9833);
nor U10577 (N_10577,N_9105,N_9316);
or U10578 (N_10578,N_9049,N_9654);
and U10579 (N_10579,N_10018,N_9421);
and U10580 (N_10580,N_10193,N_10298);
nor U10581 (N_10581,N_9844,N_10453);
and U10582 (N_10582,N_9268,N_9451);
xor U10583 (N_10583,N_9238,N_9216);
or U10584 (N_10584,N_10250,N_9394);
xnor U10585 (N_10585,N_9942,N_10320);
or U10586 (N_10586,N_9682,N_10483);
nand U10587 (N_10587,N_9293,N_9341);
xor U10588 (N_10588,N_9322,N_10081);
and U10589 (N_10589,N_9792,N_9812);
xnor U10590 (N_10590,N_9351,N_9732);
nand U10591 (N_10591,N_10059,N_9288);
or U10592 (N_10592,N_10203,N_9926);
nor U10593 (N_10593,N_9738,N_10204);
or U10594 (N_10594,N_9526,N_10257);
xnor U10595 (N_10595,N_9659,N_9997);
nor U10596 (N_10596,N_9767,N_9138);
xnor U10597 (N_10597,N_10256,N_9093);
nand U10598 (N_10598,N_9820,N_9774);
xnor U10599 (N_10599,N_9179,N_9940);
and U10600 (N_10600,N_9938,N_9198);
nand U10601 (N_10601,N_10043,N_9553);
nand U10602 (N_10602,N_10381,N_9455);
nor U10603 (N_10603,N_9701,N_9226);
xnor U10604 (N_10604,N_9328,N_9357);
nand U10605 (N_10605,N_9033,N_9215);
nand U10606 (N_10606,N_9388,N_10049);
nand U10607 (N_10607,N_9704,N_10390);
nand U10608 (N_10608,N_10356,N_9995);
nand U10609 (N_10609,N_10078,N_9018);
and U10610 (N_10610,N_9257,N_9101);
nor U10611 (N_10611,N_9067,N_9271);
nor U10612 (N_10612,N_9887,N_9827);
nor U10613 (N_10613,N_9727,N_10003);
or U10614 (N_10614,N_9760,N_10294);
or U10615 (N_10615,N_10430,N_9139);
xnor U10616 (N_10616,N_10089,N_9611);
and U10617 (N_10617,N_9510,N_9993);
nand U10618 (N_10618,N_9987,N_9415);
xnor U10619 (N_10619,N_9501,N_10221);
nor U10620 (N_10620,N_9209,N_9286);
nor U10621 (N_10621,N_9466,N_9306);
or U10622 (N_10622,N_10046,N_9831);
or U10623 (N_10623,N_10413,N_10053);
and U10624 (N_10624,N_10346,N_9115);
xor U10625 (N_10625,N_9793,N_10223);
nor U10626 (N_10626,N_9556,N_10283);
xnor U10627 (N_10627,N_9635,N_9698);
and U10628 (N_10628,N_10321,N_10036);
and U10629 (N_10629,N_9206,N_9913);
xor U10630 (N_10630,N_9180,N_9225);
nand U10631 (N_10631,N_9334,N_9608);
and U10632 (N_10632,N_9525,N_9640);
or U10633 (N_10633,N_10263,N_10175);
nor U10634 (N_10634,N_9986,N_10358);
nand U10635 (N_10635,N_9140,N_9952);
and U10636 (N_10636,N_9460,N_9669);
nand U10637 (N_10637,N_9036,N_9674);
and U10638 (N_10638,N_10048,N_10420);
or U10639 (N_10639,N_9026,N_10253);
nand U10640 (N_10640,N_10251,N_9643);
nor U10641 (N_10641,N_10135,N_9051);
xor U10642 (N_10642,N_10201,N_9908);
nor U10643 (N_10643,N_9824,N_9518);
and U10644 (N_10644,N_10155,N_9381);
or U10645 (N_10645,N_9645,N_10209);
or U10646 (N_10646,N_9676,N_10388);
xor U10647 (N_10647,N_9292,N_10076);
xnor U10648 (N_10648,N_9156,N_10016);
or U10649 (N_10649,N_9861,N_9365);
or U10650 (N_10650,N_9418,N_9151);
and U10651 (N_10651,N_9892,N_9916);
nand U10652 (N_10652,N_9001,N_10099);
or U10653 (N_10653,N_10366,N_9735);
and U10654 (N_10654,N_9166,N_9106);
xor U10655 (N_10655,N_9404,N_9971);
and U10656 (N_10656,N_9329,N_10436);
nor U10657 (N_10657,N_9379,N_10437);
or U10658 (N_10658,N_9269,N_9743);
or U10659 (N_10659,N_10246,N_9741);
or U10660 (N_10660,N_9985,N_10205);
nand U10661 (N_10661,N_10234,N_10063);
nor U10662 (N_10662,N_9481,N_9829);
or U10663 (N_10663,N_9373,N_9276);
xnor U10664 (N_10664,N_10401,N_10183);
xor U10665 (N_10665,N_10130,N_10229);
or U10666 (N_10666,N_9435,N_10170);
nor U10667 (N_10667,N_9108,N_9473);
xor U10668 (N_10668,N_9673,N_9390);
xnor U10669 (N_10669,N_9691,N_10333);
xnor U10670 (N_10670,N_10306,N_9142);
and U10671 (N_10671,N_9434,N_9874);
nor U10672 (N_10672,N_10113,N_9975);
nor U10673 (N_10673,N_9653,N_9210);
nand U10674 (N_10674,N_9898,N_9326);
or U10675 (N_10675,N_10295,N_9342);
and U10676 (N_10676,N_9871,N_10231);
or U10677 (N_10677,N_9246,N_10104);
and U10678 (N_10678,N_10019,N_10443);
nor U10679 (N_10679,N_9402,N_10010);
and U10680 (N_10680,N_9528,N_9300);
and U10681 (N_10681,N_9174,N_9838);
and U10682 (N_10682,N_9440,N_9696);
nand U10683 (N_10683,N_9011,N_9954);
nand U10684 (N_10684,N_10265,N_10387);
xnor U10685 (N_10685,N_9605,N_9345);
nand U10686 (N_10686,N_9173,N_9413);
or U10687 (N_10687,N_9515,N_9762);
nand U10688 (N_10688,N_9157,N_10403);
nor U10689 (N_10689,N_9214,N_9572);
or U10690 (N_10690,N_9802,N_9554);
nand U10691 (N_10691,N_10292,N_10186);
xor U10692 (N_10692,N_10293,N_9955);
nand U10693 (N_10693,N_9619,N_9523);
nand U10694 (N_10694,N_9646,N_9273);
and U10695 (N_10695,N_9542,N_10326);
and U10696 (N_10696,N_9739,N_9835);
or U10697 (N_10697,N_9124,N_9860);
nand U10698 (N_10698,N_9665,N_10433);
nor U10699 (N_10699,N_9930,N_9178);
nor U10700 (N_10700,N_9896,N_9612);
and U10701 (N_10701,N_9081,N_9162);
or U10702 (N_10702,N_9496,N_9432);
nand U10703 (N_10703,N_10196,N_9724);
or U10704 (N_10704,N_9720,N_9331);
nand U10705 (N_10705,N_10005,N_9711);
xor U10706 (N_10706,N_9539,N_10026);
or U10707 (N_10707,N_9052,N_9764);
nand U10708 (N_10708,N_9017,N_9374);
or U10709 (N_10709,N_9274,N_10021);
nand U10710 (N_10710,N_10328,N_10473);
and U10711 (N_10711,N_9047,N_9436);
xor U10712 (N_10712,N_9332,N_9171);
xnor U10713 (N_10713,N_9443,N_10300);
xnor U10714 (N_10714,N_9217,N_9256);
xnor U10715 (N_10715,N_9685,N_10038);
or U10716 (N_10716,N_9703,N_9649);
and U10717 (N_10717,N_9642,N_10045);
or U10718 (N_10718,N_10161,N_9119);
and U10719 (N_10719,N_9480,N_9914);
and U10720 (N_10720,N_9158,N_9947);
or U10721 (N_10721,N_9153,N_10208);
nor U10722 (N_10722,N_9264,N_9449);
xor U10723 (N_10723,N_9868,N_10254);
or U10724 (N_10724,N_9236,N_9690);
and U10725 (N_10725,N_9133,N_9089);
xor U10726 (N_10726,N_9869,N_10270);
nor U10727 (N_10727,N_9177,N_10286);
nor U10728 (N_10728,N_10389,N_9412);
nand U10729 (N_10729,N_10004,N_9856);
nor U10730 (N_10730,N_9193,N_9100);
or U10731 (N_10731,N_9909,N_9736);
nand U10732 (N_10732,N_9055,N_9516);
nor U10733 (N_10733,N_10405,N_9310);
and U10734 (N_10734,N_9983,N_10122);
nor U10735 (N_10735,N_9577,N_9768);
nand U10736 (N_10736,N_9354,N_9146);
and U10737 (N_10737,N_10216,N_10219);
or U10738 (N_10738,N_9881,N_9311);
xnor U10739 (N_10739,N_10160,N_9060);
nor U10740 (N_10740,N_9469,N_9369);
and U10741 (N_10741,N_9822,N_10281);
or U10742 (N_10742,N_9875,N_9485);
or U10743 (N_10743,N_9907,N_10125);
nand U10744 (N_10744,N_9229,N_9728);
or U10745 (N_10745,N_9076,N_9399);
and U10746 (N_10746,N_9651,N_10365);
and U10747 (N_10747,N_9550,N_9621);
or U10748 (N_10748,N_9598,N_10435);
and U10749 (N_10749,N_10307,N_10044);
and U10750 (N_10750,N_9475,N_9733);
nand U10751 (N_10751,N_9823,N_9087);
and U10752 (N_10752,N_10001,N_9776);
or U10753 (N_10753,N_10154,N_10400);
and U10754 (N_10754,N_9423,N_10417);
or U10755 (N_10755,N_9842,N_9616);
and U10756 (N_10756,N_10419,N_10481);
or U10757 (N_10757,N_9202,N_9069);
xnor U10758 (N_10758,N_9280,N_9454);
nand U10759 (N_10759,N_9984,N_9251);
or U10760 (N_10760,N_9624,N_9585);
xor U10761 (N_10761,N_9593,N_10340);
nand U10762 (N_10762,N_10376,N_10451);
xor U10763 (N_10763,N_10499,N_9731);
nand U10764 (N_10764,N_10244,N_9689);
nand U10765 (N_10765,N_9841,N_9309);
or U10766 (N_10766,N_9963,N_9786);
nor U10767 (N_10767,N_9663,N_10312);
nor U10768 (N_10768,N_9623,N_9677);
or U10769 (N_10769,N_9748,N_9941);
nand U10770 (N_10770,N_9493,N_9662);
xnor U10771 (N_10771,N_9131,N_9639);
nor U10772 (N_10772,N_9761,N_9197);
nor U10773 (N_10773,N_10117,N_9128);
nor U10774 (N_10774,N_9709,N_9949);
and U10775 (N_10775,N_9960,N_9540);
or U10776 (N_10776,N_9541,N_10230);
and U10777 (N_10777,N_9029,N_9610);
or U10778 (N_10778,N_10067,N_10344);
or U10779 (N_10779,N_10020,N_9770);
nand U10780 (N_10780,N_10411,N_9315);
and U10781 (N_10781,N_10334,N_9805);
nand U10782 (N_10782,N_10238,N_9816);
xor U10783 (N_10783,N_9467,N_9092);
and U10784 (N_10784,N_10385,N_9559);
and U10785 (N_10785,N_10108,N_9924);
nor U10786 (N_10786,N_9803,N_10329);
or U10787 (N_10787,N_9370,N_9453);
nor U10788 (N_10788,N_10308,N_9584);
xnor U10789 (N_10789,N_10452,N_9967);
or U10790 (N_10790,N_9203,N_9048);
or U10791 (N_10791,N_10282,N_10197);
xor U10792 (N_10792,N_10166,N_9050);
nand U10793 (N_10793,N_9118,N_10042);
and U10794 (N_10794,N_9301,N_9098);
nor U10795 (N_10795,N_9160,N_9058);
nand U10796 (N_10796,N_9014,N_9769);
or U10797 (N_10797,N_9305,N_10396);
nor U10798 (N_10798,N_10468,N_9488);
or U10799 (N_10799,N_9495,N_10335);
and U10800 (N_10800,N_9490,N_9514);
or U10801 (N_10801,N_9836,N_9604);
and U10802 (N_10802,N_9758,N_9527);
nor U10803 (N_10803,N_9114,N_10271);
xor U10804 (N_10804,N_9990,N_10202);
nand U10805 (N_10805,N_9313,N_10434);
xor U10806 (N_10806,N_10297,N_9330);
xor U10807 (N_10807,N_10379,N_9870);
xor U10808 (N_10808,N_9922,N_9410);
xor U10809 (N_10809,N_9112,N_9396);
and U10810 (N_10810,N_9688,N_10169);
or U10811 (N_10811,N_9107,N_9684);
nor U10812 (N_10812,N_9103,N_9385);
xor U10813 (N_10813,N_10136,N_9259);
nand U10814 (N_10814,N_9136,N_10259);
and U10815 (N_10815,N_9590,N_9532);
and U10816 (N_10816,N_10047,N_10375);
xnor U10817 (N_10817,N_10267,N_9095);
nor U10818 (N_10818,N_9849,N_9613);
xor U10819 (N_10819,N_9615,N_9211);
nor U10820 (N_10820,N_9726,N_10382);
or U10821 (N_10821,N_9348,N_9129);
or U10822 (N_10822,N_10171,N_10336);
nand U10823 (N_10823,N_9375,N_10367);
xnor U10824 (N_10824,N_10418,N_9522);
or U10825 (N_10825,N_9814,N_10440);
and U10826 (N_10826,N_10415,N_9622);
or U10827 (N_10827,N_10093,N_9583);
or U10828 (N_10828,N_9289,N_10338);
or U10829 (N_10829,N_10068,N_10150);
and U10830 (N_10830,N_9798,N_9509);
nand U10831 (N_10831,N_9478,N_9470);
and U10832 (N_10832,N_10316,N_9419);
nor U10833 (N_10833,N_10174,N_10207);
and U10834 (N_10834,N_10474,N_10194);
or U10835 (N_10835,N_9380,N_9320);
nor U10836 (N_10836,N_10486,N_10353);
and U10837 (N_10837,N_9270,N_10406);
or U10838 (N_10838,N_9923,N_9666);
and U10839 (N_10839,N_9122,N_10052);
or U10840 (N_10840,N_9890,N_9184);
nand U10841 (N_10841,N_10348,N_10252);
nor U10842 (N_10842,N_10027,N_9297);
nor U10843 (N_10843,N_9601,N_10152);
nor U10844 (N_10844,N_10009,N_9692);
and U10845 (N_10845,N_10427,N_9777);
xor U10846 (N_10846,N_10352,N_9045);
nor U10847 (N_10847,N_9863,N_10115);
nor U10848 (N_10848,N_10079,N_9497);
nand U10849 (N_10849,N_10373,N_9977);
or U10850 (N_10850,N_10008,N_9629);
or U10851 (N_10851,N_9285,N_10260);
or U10852 (N_10852,N_10277,N_9745);
and U10853 (N_10853,N_9806,N_10157);
or U10854 (N_10854,N_9529,N_9006);
and U10855 (N_10855,N_10015,N_10359);
or U10856 (N_10856,N_10239,N_10012);
nand U10857 (N_10857,N_9575,N_10031);
or U10858 (N_10858,N_10206,N_9706);
nand U10859 (N_10859,N_10121,N_9638);
or U10860 (N_10860,N_10339,N_9181);
nor U10861 (N_10861,N_9927,N_9700);
nor U10862 (N_10862,N_10062,N_10144);
and U10863 (N_10863,N_9350,N_10102);
nor U10864 (N_10864,N_9899,N_10195);
and U10865 (N_10865,N_9291,N_9000);
and U10866 (N_10866,N_10217,N_10496);
or U10867 (N_10867,N_10111,N_9504);
or U10868 (N_10868,N_9457,N_9471);
nor U10869 (N_10869,N_10383,N_10191);
nor U10870 (N_10870,N_9888,N_9637);
and U10871 (N_10871,N_9068,N_10212);
and U10872 (N_10872,N_10187,N_9788);
xnor U10873 (N_10873,N_9126,N_10245);
nor U10874 (N_10874,N_10077,N_9169);
nor U10875 (N_10875,N_9143,N_9715);
xnor U10876 (N_10876,N_9059,N_10030);
nand U10877 (N_10877,N_9614,N_9258);
nor U10878 (N_10878,N_9809,N_10133);
nand U10879 (N_10879,N_9015,N_10100);
nand U10880 (N_10880,N_10000,N_9376);
and U10881 (N_10881,N_9519,N_10181);
nor U10882 (N_10882,N_10007,N_9897);
xnor U10883 (N_10883,N_9589,N_10014);
nand U10884 (N_10884,N_10399,N_10147);
xor U10885 (N_10885,N_10051,N_9972);
and U10886 (N_10886,N_9111,N_9549);
xnor U10887 (N_10887,N_9420,N_9022);
or U10888 (N_10888,N_9876,N_9749);
nand U10889 (N_10889,N_9573,N_10075);
xnor U10890 (N_10890,N_9308,N_9458);
and U10891 (N_10891,N_9530,N_10060);
and U10892 (N_10892,N_9969,N_9680);
and U10893 (N_10893,N_9392,N_10414);
nor U10894 (N_10894,N_10485,N_9965);
and U10895 (N_10895,N_10302,N_9065);
or U10896 (N_10896,N_9866,N_9431);
nor U10897 (N_10897,N_9057,N_9083);
xor U10898 (N_10898,N_10096,N_9425);
or U10899 (N_10899,N_10087,N_10222);
and U10900 (N_10900,N_9791,N_9327);
or U10901 (N_10901,N_9150,N_9982);
nor U10902 (N_10902,N_9323,N_9278);
nand U10903 (N_10903,N_9817,N_10454);
nand U10904 (N_10904,N_9465,N_9734);
or U10905 (N_10905,N_9839,N_9428);
or U10906 (N_10906,N_9789,N_10172);
nor U10907 (N_10907,N_9880,N_9891);
xor U10908 (N_10908,N_9172,N_9452);
nor U10909 (N_10909,N_10445,N_9020);
and U10910 (N_10910,N_10290,N_9533);
nand U10911 (N_10911,N_9929,N_10041);
nor U10912 (N_10912,N_9580,N_9163);
or U10913 (N_10913,N_9248,N_9031);
and U10914 (N_10914,N_9352,N_9430);
nand U10915 (N_10915,N_9565,N_10092);
or U10916 (N_10916,N_9921,N_9534);
nor U10917 (N_10917,N_10378,N_10458);
xnor U10918 (N_10918,N_10235,N_9946);
nor U10919 (N_10919,N_9834,N_9041);
xor U10920 (N_10920,N_9168,N_9008);
or U10921 (N_10921,N_9344,N_10369);
xnor U10922 (N_10922,N_9958,N_10416);
xnor U10923 (N_10923,N_9340,N_10397);
or U10924 (N_10924,N_10354,N_9398);
or U10925 (N_10925,N_9377,N_9070);
xor U10926 (N_10926,N_10006,N_9647);
nor U10927 (N_10927,N_9170,N_10469);
nand U10928 (N_10928,N_9708,N_9832);
and U10929 (N_10929,N_9576,N_9450);
and U10930 (N_10930,N_9634,N_9207);
xor U10931 (N_10931,N_9775,N_9367);
nand U10932 (N_10932,N_10425,N_10137);
nand U10933 (N_10933,N_9851,N_9296);
xnor U10934 (N_10934,N_9994,N_9950);
or U10935 (N_10935,N_9232,N_10177);
and U10936 (N_10936,N_9164,N_9721);
or U10937 (N_10937,N_10317,N_9600);
and U10938 (N_10938,N_9686,N_9494);
nor U10939 (N_10939,N_9931,N_10029);
xor U10940 (N_10940,N_10192,N_9391);
nand U10941 (N_10941,N_9574,N_9338);
xnor U10942 (N_10942,N_10248,N_9710);
xnor U10943 (N_10943,N_9027,N_10479);
or U10944 (N_10944,N_9094,N_10269);
nor U10945 (N_10945,N_9627,N_9882);
nor U10946 (N_10946,N_9267,N_10467);
nor U10947 (N_10947,N_10459,N_10476);
nand U10948 (N_10948,N_9578,N_10188);
nor U10949 (N_10949,N_9591,N_9190);
and U10950 (N_10950,N_10132,N_9719);
nor U10951 (N_10951,N_9079,N_9080);
nor U10952 (N_10952,N_9636,N_9979);
nor U10953 (N_10953,N_9347,N_9299);
nor U10954 (N_10954,N_9609,N_10466);
or U10955 (N_10955,N_9123,N_9424);
xnor U10956 (N_10956,N_9672,N_9937);
or U10957 (N_10957,N_10487,N_10291);
nor U10958 (N_10958,N_9295,N_9795);
or U10959 (N_10959,N_10129,N_9702);
and U10960 (N_10960,N_10057,N_9902);
nor U10961 (N_10961,N_9078,N_9904);
or U10962 (N_10962,N_9723,N_9130);
xor U10963 (N_10963,N_9846,N_10289);
and U10964 (N_10964,N_9545,N_9678);
xnor U10965 (N_10965,N_9730,N_9906);
and U10966 (N_10966,N_9765,N_9109);
xor U10967 (N_10967,N_10039,N_9631);
nand U10968 (N_10968,N_10119,N_9149);
nor U10969 (N_10969,N_9976,N_9165);
xnor U10970 (N_10970,N_10284,N_9104);
nor U10971 (N_10971,N_9228,N_9594);
nor U10972 (N_10972,N_10124,N_10325);
nand U10973 (N_10973,N_9038,N_9075);
nand U10974 (N_10974,N_9152,N_9243);
or U10975 (N_10975,N_10368,N_9234);
nand U10976 (N_10976,N_9943,N_9134);
xor U10977 (N_10977,N_9132,N_9988);
and U10978 (N_10978,N_9378,N_10363);
or U10979 (N_10979,N_9819,N_9740);
nor U10980 (N_10980,N_9505,N_10189);
nor U10981 (N_10981,N_10391,N_9668);
nand U10982 (N_10982,N_9249,N_9694);
xor U10983 (N_10983,N_10490,N_9116);
xnor U10984 (N_10984,N_9056,N_10083);
and U10985 (N_10985,N_10120,N_9959);
xnor U10986 (N_10986,N_9371,N_9850);
or U10987 (N_10987,N_10240,N_9705);
nor U10988 (N_10988,N_10327,N_9925);
nor U10989 (N_10989,N_9220,N_10331);
xnor U10990 (N_10990,N_10198,N_9644);
nor U10991 (N_10991,N_9414,N_9957);
or U10992 (N_10992,N_10261,N_9186);
and U10993 (N_10993,N_9482,N_9915);
nand U10994 (N_10994,N_9427,N_9981);
xor U10995 (N_10995,N_9566,N_10156);
and U10996 (N_10996,N_9961,N_9061);
nand U10997 (N_10997,N_10477,N_10032);
or U10998 (N_10998,N_9298,N_9655);
or U10999 (N_10999,N_9486,N_9537);
or U11000 (N_11000,N_10410,N_9586);
xor U11001 (N_11001,N_10268,N_10384);
and U11002 (N_11002,N_9175,N_9847);
xnor U11003 (N_11003,N_10360,N_9227);
nor U11004 (N_11004,N_10278,N_10315);
or U11005 (N_11005,N_9607,N_9034);
nor U11006 (N_11006,N_9737,N_9287);
xnor U11007 (N_11007,N_9387,N_9563);
nor U11008 (N_11008,N_9077,N_10262);
nand U11009 (N_11009,N_10301,N_9617);
nor U11010 (N_11010,N_10128,N_9895);
nor U11011 (N_11011,N_9205,N_9999);
or U11012 (N_11012,N_9800,N_9858);
and U11013 (N_11013,N_9944,N_9196);
nor U11014 (N_11014,N_9363,N_9520);
or U11015 (N_11015,N_10241,N_9582);
and U11016 (N_11016,N_10088,N_9713);
xor U11017 (N_11017,N_9828,N_9120);
and U11018 (N_11018,N_9461,N_10176);
nor U11019 (N_11019,N_9722,N_9893);
or U11020 (N_11020,N_9383,N_10398);
xnor U11021 (N_11021,N_9110,N_10404);
nand U11022 (N_11022,N_10460,N_9364);
nor U11023 (N_11023,N_9811,N_9751);
xnor U11024 (N_11024,N_9062,N_10448);
nand U11025 (N_11025,N_9857,N_9195);
nor U11026 (N_11026,N_9386,N_10105);
and U11027 (N_11027,N_10370,N_9409);
or U11028 (N_11028,N_10428,N_10442);
xor U11029 (N_11029,N_9650,N_10347);
nand U11030 (N_11030,N_9948,N_10140);
xnor U11031 (N_11031,N_10101,N_9444);
or U11032 (N_11032,N_10371,N_9084);
nor U11033 (N_11033,N_9602,N_10071);
and U11034 (N_11034,N_10275,N_10178);
nand U11035 (N_11035,N_9813,N_9503);
nor U11036 (N_11036,N_9920,N_9422);
xor U11037 (N_11037,N_9155,N_10319);
nand U11038 (N_11038,N_10055,N_9233);
and U11039 (N_11039,N_9511,N_10109);
xor U11040 (N_11040,N_9144,N_9013);
xor U11041 (N_11041,N_9125,N_10493);
xnor U11042 (N_11042,N_9918,N_10322);
nor U11043 (N_11043,N_9400,N_9889);
xnor U11044 (N_11044,N_10475,N_10303);
and U11045 (N_11045,N_9825,N_9010);
or U11046 (N_11046,N_9561,N_9489);
or U11047 (N_11047,N_9201,N_10163);
and U11048 (N_11048,N_9044,N_9498);
and U11049 (N_11049,N_10141,N_9592);
or U11050 (N_11050,N_9855,N_9353);
or U11051 (N_11051,N_10072,N_10408);
and U11052 (N_11052,N_10090,N_10489);
nand U11053 (N_11053,N_10407,N_10158);
and U11054 (N_11054,N_10082,N_10380);
and U11055 (N_11055,N_9980,N_9917);
xor U11056 (N_11056,N_9272,N_9030);
xor U11057 (N_11057,N_10112,N_9712);
nor U11058 (N_11058,N_9867,N_9729);
or U11059 (N_11059,N_9945,N_9337);
xnor U11060 (N_11060,N_10127,N_9796);
or U11061 (N_11061,N_9063,N_9349);
nor U11062 (N_11062,N_10094,N_9426);
xnor U11063 (N_11063,N_10213,N_9707);
and U11064 (N_11064,N_9974,N_9794);
or U11065 (N_11065,N_9137,N_9699);
nand U11066 (N_11066,N_10276,N_9661);
nand U11067 (N_11067,N_9040,N_9360);
nor U11068 (N_11068,N_9782,N_9536);
nand U11069 (N_11069,N_9245,N_9632);
nor U11070 (N_11070,N_9755,N_10441);
and U11071 (N_11071,N_10304,N_9883);
xor U11072 (N_11072,N_10226,N_9718);
nand U11073 (N_11073,N_9148,N_9263);
nor U11074 (N_11074,N_9382,N_9303);
xnor U11075 (N_11075,N_9355,N_9255);
nor U11076 (N_11076,N_9417,N_9966);
or U11077 (N_11077,N_10402,N_9657);
and U11078 (N_11078,N_9007,N_9815);
nor U11079 (N_11079,N_9989,N_10431);
nand U11080 (N_11080,N_9403,N_9053);
and U11081 (N_11081,N_10107,N_10438);
nand U11082 (N_11082,N_10097,N_9199);
nand U11083 (N_11083,N_10350,N_10310);
or U11084 (N_11084,N_10126,N_9071);
or U11085 (N_11085,N_9821,N_9009);
xnor U11086 (N_11086,N_10131,N_9135);
xnor U11087 (N_11087,N_9517,N_10106);
xor U11088 (N_11088,N_9240,N_10461);
and U11089 (N_11089,N_9393,N_10482);
xor U11090 (N_11090,N_10162,N_10143);
nor U11091 (N_11091,N_9973,N_10472);
and U11092 (N_11092,N_9603,N_10323);
xnor U11093 (N_11093,N_9521,N_9102);
xor U11094 (N_11094,N_10446,N_9970);
xnor U11095 (N_11095,N_10025,N_9548);
nor U11096 (N_11096,N_9964,N_9191);
xor U11097 (N_11097,N_10054,N_10237);
or U11098 (N_11098,N_9807,N_9312);
and U11099 (N_11099,N_9756,N_10149);
nand U11100 (N_11100,N_9744,N_10279);
and U11101 (N_11101,N_10285,N_9656);
xnor U11102 (N_11102,N_10084,N_9476);
and U11103 (N_11103,N_9859,N_10040);
or U11104 (N_11104,N_9072,N_9992);
and U11105 (N_11105,N_9012,N_9512);
xor U11106 (N_11106,N_9325,N_9253);
and U11107 (N_11107,N_9442,N_10211);
and U11108 (N_11108,N_10478,N_9919);
nor U11109 (N_11109,N_9932,N_9456);
xor U11110 (N_11110,N_10069,N_10449);
and U11111 (N_11111,N_9188,N_10110);
nor U11112 (N_11112,N_9082,N_9281);
xnor U11113 (N_11113,N_9848,N_9194);
nand U11114 (N_11114,N_9239,N_9683);
xor U11115 (N_11115,N_10288,N_9066);
nand U11116 (N_11116,N_9546,N_10361);
nor U11117 (N_11117,N_9853,N_10086);
xnor U11118 (N_11118,N_9752,N_9361);
nor U11119 (N_11119,N_9625,N_9935);
nor U11120 (N_11120,N_9241,N_10173);
xor U11121 (N_11121,N_9235,N_9252);
nand U11122 (N_11122,N_9569,N_10498);
xnor U11123 (N_11123,N_9885,N_9753);
nand U11124 (N_11124,N_10074,N_9159);
xnor U11125 (N_11125,N_10421,N_9192);
xnor U11126 (N_11126,N_10455,N_9437);
and U11127 (N_11127,N_9037,N_9200);
nor U11128 (N_11128,N_9939,N_10034);
nor U11129 (N_11129,N_9405,N_10299);
or U11130 (N_11130,N_9411,N_10247);
and U11131 (N_11131,N_9597,N_10118);
nand U11132 (N_11132,N_9333,N_9438);
nand U11133 (N_11133,N_9230,N_10470);
nor U11134 (N_11134,N_9016,N_10224);
nor U11135 (N_11135,N_9500,N_9176);
or U11136 (N_11136,N_10228,N_10494);
nor U11137 (N_11137,N_10200,N_9778);
nand U11138 (N_11138,N_10412,N_9571);
xor U11139 (N_11139,N_9477,N_9681);
and U11140 (N_11140,N_9319,N_9439);
xnor U11141 (N_11141,N_10296,N_9356);
and U11142 (N_11142,N_9359,N_9117);
and U11143 (N_11143,N_9261,N_9127);
and U11144 (N_11144,N_10422,N_10480);
or U11145 (N_11145,N_10227,N_9003);
or U11146 (N_11146,N_9479,N_9187);
and U11147 (N_11147,N_9384,N_10311);
nor U11148 (N_11148,N_9886,N_9587);
or U11149 (N_11149,N_9307,N_10184);
and U11150 (N_11150,N_9366,N_10225);
or U11151 (N_11151,N_9804,N_9780);
or U11152 (N_11152,N_10070,N_10168);
xnor U11153 (N_11153,N_10484,N_10255);
and U11154 (N_11154,N_10134,N_9182);
and U11155 (N_11155,N_10374,N_10050);
nor U11156 (N_11156,N_10085,N_10214);
or U11157 (N_11157,N_10080,N_9951);
xor U11158 (N_11158,N_10199,N_10395);
nor U11159 (N_11159,N_10220,N_9852);
xnor U11160 (N_11160,N_10349,N_10167);
and U11161 (N_11161,N_9783,N_9716);
xor U11162 (N_11162,N_10058,N_9464);
and U11163 (N_11163,N_10123,N_10273);
xnor U11164 (N_11164,N_10464,N_9433);
nor U11165 (N_11165,N_9218,N_10249);
xor U11166 (N_11166,N_9968,N_9742);
nand U11167 (N_11167,N_9262,N_10305);
nand U11168 (N_11168,N_9317,N_9223);
nor U11169 (N_11169,N_10037,N_10011);
and U11170 (N_11170,N_9250,N_9204);
and U11171 (N_11171,N_9544,N_10324);
nor U11172 (N_11172,N_9441,N_9406);
nand U11173 (N_11173,N_9826,N_9408);
nor U11174 (N_11174,N_9543,N_9028);
and U11175 (N_11175,N_9021,N_9282);
and U11176 (N_11176,N_9750,N_9879);
or U11177 (N_11177,N_9658,N_9581);
nor U11178 (N_11178,N_10471,N_10426);
nor U11179 (N_11179,N_9244,N_10318);
xor U11180 (N_11180,N_9996,N_9275);
xnor U11181 (N_11181,N_9552,N_10313);
nor U11182 (N_11182,N_9797,N_10342);
nand U11183 (N_11183,N_9962,N_9025);
nor U11184 (N_11184,N_9290,N_9725);
or U11185 (N_11185,N_9911,N_10450);
nor U11186 (N_11186,N_10243,N_10439);
nor U11187 (N_11187,N_9555,N_9416);
or U11188 (N_11188,N_9628,N_9284);
nand U11189 (N_11189,N_10429,N_9670);
nor U11190 (N_11190,N_10142,N_9991);
nand U11191 (N_11191,N_10330,N_9086);
and U11192 (N_11192,N_9717,N_10456);
and U11193 (N_11193,N_9231,N_9064);
and U11194 (N_11194,N_9978,N_9004);
nand U11195 (N_11195,N_9314,N_9693);
xnor U11196 (N_11196,N_9877,N_10287);
or U11197 (N_11197,N_9664,N_9091);
nor U11198 (N_11198,N_9697,N_9845);
xor U11199 (N_11199,N_10272,N_9447);
xnor U11200 (N_11200,N_9508,N_9558);
nor U11201 (N_11201,N_10497,N_9953);
or U11202 (N_11202,N_10309,N_9687);
xor U11203 (N_11203,N_9448,N_10491);
and U11204 (N_11204,N_9854,N_9224);
xor U11205 (N_11205,N_9771,N_9074);
xnor U11206 (N_11206,N_9873,N_9862);
nand U11207 (N_11207,N_10364,N_10233);
nor U11208 (N_11208,N_10024,N_9043);
nand U11209 (N_11209,N_9933,N_9567);
nor U11210 (N_11210,N_9283,N_9506);
nor U11211 (N_11211,N_9019,N_10179);
nand U11212 (N_11212,N_9547,N_9785);
nand U11213 (N_11213,N_9903,N_10337);
nand U11214 (N_11214,N_9266,N_9757);
xnor U11215 (N_11215,N_9588,N_9032);
xor U11216 (N_11216,N_10017,N_10409);
and U11217 (N_11217,N_9023,N_9085);
or U11218 (N_11218,N_10182,N_10138);
or U11219 (N_11219,N_9630,N_9468);
and U11220 (N_11220,N_9538,N_9161);
xnor U11221 (N_11221,N_10343,N_9766);
xnor U11222 (N_11222,N_10190,N_10423);
xor U11223 (N_11223,N_9560,N_9459);
nand U11224 (N_11224,N_9524,N_10232);
nand U11225 (N_11225,N_9260,N_9279);
and U11226 (N_11226,N_9222,N_10215);
and U11227 (N_11227,N_9121,N_9675);
and U11228 (N_11228,N_9652,N_10432);
xnor U11229 (N_11229,N_10362,N_9463);
nand U11230 (N_11230,N_9294,N_9936);
or U11231 (N_11231,N_9167,N_9840);
and U11232 (N_11232,N_9492,N_10185);
and U11233 (N_11233,N_9336,N_9141);
nor U11234 (N_11234,N_9189,N_9633);
or U11235 (N_11235,N_9595,N_10488);
or U11236 (N_11236,N_9901,N_9090);
and U11237 (N_11237,N_9054,N_10210);
or U11238 (N_11238,N_10056,N_9339);
and U11239 (N_11239,N_9277,N_10218);
and U11240 (N_11240,N_9830,N_10357);
nor U11241 (N_11241,N_9213,N_9145);
nor U11242 (N_11242,N_9878,N_10393);
and U11243 (N_11243,N_10280,N_9395);
or U11244 (N_11244,N_10151,N_10394);
and U11245 (N_11245,N_9097,N_9754);
nand U11246 (N_11246,N_10013,N_9484);
nand U11247 (N_11247,N_9865,N_10465);
nor U11248 (N_11248,N_9318,N_9219);
and U11249 (N_11249,N_9483,N_10116);
nor U11250 (N_11250,N_9560,N_10110);
xor U11251 (N_11251,N_9712,N_9271);
or U11252 (N_11252,N_9202,N_10275);
nand U11253 (N_11253,N_9284,N_9155);
or U11254 (N_11254,N_10381,N_9734);
or U11255 (N_11255,N_9480,N_10279);
and U11256 (N_11256,N_9518,N_10117);
xor U11257 (N_11257,N_10144,N_9336);
nand U11258 (N_11258,N_9515,N_9211);
nor U11259 (N_11259,N_10457,N_10385);
and U11260 (N_11260,N_10111,N_10481);
xnor U11261 (N_11261,N_10162,N_10125);
xnor U11262 (N_11262,N_9620,N_9819);
nor U11263 (N_11263,N_9257,N_9567);
nand U11264 (N_11264,N_10093,N_9350);
nor U11265 (N_11265,N_9081,N_10218);
and U11266 (N_11266,N_10106,N_9938);
or U11267 (N_11267,N_9913,N_9364);
or U11268 (N_11268,N_9927,N_9170);
and U11269 (N_11269,N_9721,N_9259);
nand U11270 (N_11270,N_9746,N_9165);
nand U11271 (N_11271,N_9715,N_10049);
xnor U11272 (N_11272,N_9998,N_9652);
nor U11273 (N_11273,N_9705,N_9879);
and U11274 (N_11274,N_10475,N_10334);
nand U11275 (N_11275,N_9273,N_9390);
xnor U11276 (N_11276,N_9360,N_9517);
or U11277 (N_11277,N_9997,N_9833);
or U11278 (N_11278,N_9544,N_9000);
xor U11279 (N_11279,N_9992,N_9143);
xor U11280 (N_11280,N_9915,N_10215);
or U11281 (N_11281,N_9933,N_9357);
and U11282 (N_11282,N_10231,N_9816);
or U11283 (N_11283,N_9518,N_10450);
and U11284 (N_11284,N_9945,N_9269);
xnor U11285 (N_11285,N_9136,N_9956);
nor U11286 (N_11286,N_9477,N_10119);
and U11287 (N_11287,N_9371,N_9708);
nand U11288 (N_11288,N_9355,N_9893);
or U11289 (N_11289,N_9670,N_10250);
and U11290 (N_11290,N_10462,N_10390);
xnor U11291 (N_11291,N_9657,N_10398);
nor U11292 (N_11292,N_9569,N_10137);
nand U11293 (N_11293,N_9804,N_9670);
nand U11294 (N_11294,N_9531,N_9880);
or U11295 (N_11295,N_9395,N_9405);
and U11296 (N_11296,N_9213,N_9093);
xnor U11297 (N_11297,N_10137,N_10212);
and U11298 (N_11298,N_9480,N_9115);
or U11299 (N_11299,N_10130,N_9673);
xnor U11300 (N_11300,N_9466,N_9313);
xor U11301 (N_11301,N_10353,N_10035);
and U11302 (N_11302,N_9963,N_9185);
xor U11303 (N_11303,N_9777,N_9546);
xor U11304 (N_11304,N_9502,N_9267);
or U11305 (N_11305,N_10048,N_10207);
xor U11306 (N_11306,N_9140,N_9731);
xor U11307 (N_11307,N_10291,N_9620);
xnor U11308 (N_11308,N_9731,N_9723);
nand U11309 (N_11309,N_9135,N_9595);
xor U11310 (N_11310,N_10389,N_10339);
nand U11311 (N_11311,N_9214,N_9525);
nor U11312 (N_11312,N_9298,N_10233);
xor U11313 (N_11313,N_10029,N_9414);
or U11314 (N_11314,N_9514,N_9113);
or U11315 (N_11315,N_10407,N_10002);
and U11316 (N_11316,N_10070,N_10228);
and U11317 (N_11317,N_9674,N_9627);
nand U11318 (N_11318,N_9081,N_9240);
nand U11319 (N_11319,N_10247,N_10027);
nor U11320 (N_11320,N_10137,N_9839);
or U11321 (N_11321,N_10053,N_9445);
nand U11322 (N_11322,N_10437,N_9633);
xor U11323 (N_11323,N_9717,N_10076);
and U11324 (N_11324,N_9827,N_10075);
or U11325 (N_11325,N_9245,N_9208);
xor U11326 (N_11326,N_10081,N_9633);
or U11327 (N_11327,N_10439,N_10434);
nand U11328 (N_11328,N_10242,N_10016);
or U11329 (N_11329,N_9523,N_9787);
nand U11330 (N_11330,N_9550,N_10245);
xor U11331 (N_11331,N_9229,N_9816);
nand U11332 (N_11332,N_9384,N_9390);
nand U11333 (N_11333,N_9432,N_10020);
xnor U11334 (N_11334,N_10237,N_9485);
and U11335 (N_11335,N_9906,N_9426);
or U11336 (N_11336,N_10374,N_9399);
xnor U11337 (N_11337,N_9206,N_9334);
nor U11338 (N_11338,N_10261,N_9064);
or U11339 (N_11339,N_9292,N_9183);
or U11340 (N_11340,N_9889,N_9132);
nand U11341 (N_11341,N_9959,N_9382);
xnor U11342 (N_11342,N_9826,N_10014);
nand U11343 (N_11343,N_10306,N_10253);
and U11344 (N_11344,N_9372,N_9357);
and U11345 (N_11345,N_10314,N_9413);
or U11346 (N_11346,N_9741,N_10164);
xnor U11347 (N_11347,N_9181,N_9160);
and U11348 (N_11348,N_10476,N_9470);
xnor U11349 (N_11349,N_10382,N_9593);
and U11350 (N_11350,N_9680,N_9629);
or U11351 (N_11351,N_9103,N_10302);
or U11352 (N_11352,N_9282,N_9307);
nor U11353 (N_11353,N_9185,N_9687);
nor U11354 (N_11354,N_9830,N_9047);
nand U11355 (N_11355,N_9069,N_9895);
nor U11356 (N_11356,N_9186,N_9375);
and U11357 (N_11357,N_9144,N_9531);
and U11358 (N_11358,N_9530,N_9330);
or U11359 (N_11359,N_10119,N_9938);
nand U11360 (N_11360,N_10380,N_9822);
nand U11361 (N_11361,N_9440,N_10118);
nor U11362 (N_11362,N_9964,N_10070);
xor U11363 (N_11363,N_10369,N_9110);
nand U11364 (N_11364,N_9341,N_10152);
and U11365 (N_11365,N_10160,N_9427);
and U11366 (N_11366,N_10353,N_10275);
nand U11367 (N_11367,N_10217,N_10132);
and U11368 (N_11368,N_10260,N_9321);
or U11369 (N_11369,N_9710,N_9197);
or U11370 (N_11370,N_10221,N_9828);
nor U11371 (N_11371,N_10126,N_9081);
nor U11372 (N_11372,N_10086,N_10339);
nand U11373 (N_11373,N_9654,N_9280);
nand U11374 (N_11374,N_10102,N_9089);
nand U11375 (N_11375,N_10197,N_9850);
xnor U11376 (N_11376,N_10285,N_10327);
nor U11377 (N_11377,N_10462,N_9215);
or U11378 (N_11378,N_9747,N_9578);
and U11379 (N_11379,N_10045,N_9051);
nor U11380 (N_11380,N_9662,N_10063);
xnor U11381 (N_11381,N_10248,N_9661);
nor U11382 (N_11382,N_9366,N_10465);
and U11383 (N_11383,N_9499,N_9090);
nor U11384 (N_11384,N_9824,N_10499);
and U11385 (N_11385,N_9857,N_9133);
nand U11386 (N_11386,N_9371,N_10396);
xor U11387 (N_11387,N_10317,N_10256);
nand U11388 (N_11388,N_9248,N_10190);
nand U11389 (N_11389,N_10407,N_9758);
nor U11390 (N_11390,N_10038,N_9411);
nand U11391 (N_11391,N_9200,N_9506);
xor U11392 (N_11392,N_9522,N_9760);
and U11393 (N_11393,N_10098,N_9783);
nor U11394 (N_11394,N_9894,N_9026);
nand U11395 (N_11395,N_9518,N_9913);
nor U11396 (N_11396,N_9396,N_9417);
and U11397 (N_11397,N_9405,N_9922);
nor U11398 (N_11398,N_9831,N_9880);
or U11399 (N_11399,N_9217,N_10480);
nand U11400 (N_11400,N_10037,N_10210);
or U11401 (N_11401,N_10324,N_10010);
xor U11402 (N_11402,N_9939,N_9364);
and U11403 (N_11403,N_10015,N_9014);
nor U11404 (N_11404,N_10385,N_9082);
xor U11405 (N_11405,N_9453,N_10075);
xor U11406 (N_11406,N_10221,N_9992);
xor U11407 (N_11407,N_10039,N_9208);
xor U11408 (N_11408,N_9968,N_9699);
xor U11409 (N_11409,N_9680,N_9188);
nand U11410 (N_11410,N_9423,N_9297);
or U11411 (N_11411,N_10426,N_9277);
and U11412 (N_11412,N_9899,N_9627);
nor U11413 (N_11413,N_9746,N_10339);
nor U11414 (N_11414,N_10262,N_10057);
nor U11415 (N_11415,N_9774,N_9201);
nor U11416 (N_11416,N_9189,N_9969);
xor U11417 (N_11417,N_9799,N_9278);
xnor U11418 (N_11418,N_9578,N_9739);
or U11419 (N_11419,N_9704,N_9178);
or U11420 (N_11420,N_9676,N_9573);
xor U11421 (N_11421,N_9104,N_9877);
xnor U11422 (N_11422,N_10215,N_9572);
and U11423 (N_11423,N_9507,N_9701);
and U11424 (N_11424,N_9958,N_10190);
nand U11425 (N_11425,N_9683,N_9543);
or U11426 (N_11426,N_10493,N_9854);
xnor U11427 (N_11427,N_9961,N_9913);
and U11428 (N_11428,N_9620,N_10147);
and U11429 (N_11429,N_9469,N_9211);
and U11430 (N_11430,N_9354,N_9975);
or U11431 (N_11431,N_9017,N_9964);
nand U11432 (N_11432,N_9962,N_9080);
or U11433 (N_11433,N_9766,N_9828);
xnor U11434 (N_11434,N_10168,N_9296);
nor U11435 (N_11435,N_9697,N_9541);
nand U11436 (N_11436,N_9345,N_9673);
xor U11437 (N_11437,N_9814,N_9238);
nand U11438 (N_11438,N_9924,N_10418);
nor U11439 (N_11439,N_10390,N_9189);
and U11440 (N_11440,N_9709,N_10128);
nand U11441 (N_11441,N_10357,N_9422);
nand U11442 (N_11442,N_9040,N_9686);
or U11443 (N_11443,N_9537,N_9358);
xnor U11444 (N_11444,N_9653,N_9478);
nor U11445 (N_11445,N_9432,N_9772);
or U11446 (N_11446,N_9853,N_9071);
and U11447 (N_11447,N_9058,N_9877);
nand U11448 (N_11448,N_10112,N_9016);
nand U11449 (N_11449,N_10361,N_9512);
nor U11450 (N_11450,N_10363,N_9998);
nand U11451 (N_11451,N_9693,N_10236);
nand U11452 (N_11452,N_10184,N_10229);
nand U11453 (N_11453,N_9577,N_9476);
or U11454 (N_11454,N_9459,N_10054);
or U11455 (N_11455,N_10203,N_10237);
or U11456 (N_11456,N_9796,N_9964);
nand U11457 (N_11457,N_10021,N_9492);
xor U11458 (N_11458,N_9212,N_9571);
nand U11459 (N_11459,N_9156,N_9325);
or U11460 (N_11460,N_9678,N_9497);
nor U11461 (N_11461,N_10014,N_9495);
xor U11462 (N_11462,N_9308,N_9926);
nor U11463 (N_11463,N_9592,N_10441);
nand U11464 (N_11464,N_9040,N_9486);
nand U11465 (N_11465,N_9838,N_10194);
nand U11466 (N_11466,N_9043,N_9076);
nand U11467 (N_11467,N_9167,N_9325);
nor U11468 (N_11468,N_9587,N_9574);
nor U11469 (N_11469,N_9605,N_10039);
and U11470 (N_11470,N_9388,N_9550);
and U11471 (N_11471,N_10382,N_9098);
xnor U11472 (N_11472,N_9878,N_10006);
and U11473 (N_11473,N_9487,N_9047);
or U11474 (N_11474,N_9312,N_9183);
nor U11475 (N_11475,N_9355,N_9581);
and U11476 (N_11476,N_9239,N_9271);
nor U11477 (N_11477,N_9413,N_10117);
nor U11478 (N_11478,N_9989,N_10437);
xnor U11479 (N_11479,N_9113,N_10039);
or U11480 (N_11480,N_10432,N_9191);
or U11481 (N_11481,N_10448,N_10089);
and U11482 (N_11482,N_9195,N_10206);
and U11483 (N_11483,N_9992,N_10026);
or U11484 (N_11484,N_9883,N_9446);
xor U11485 (N_11485,N_10017,N_9200);
nor U11486 (N_11486,N_10259,N_9989);
nand U11487 (N_11487,N_9210,N_9497);
or U11488 (N_11488,N_10257,N_10165);
and U11489 (N_11489,N_9821,N_10307);
and U11490 (N_11490,N_10161,N_9123);
nor U11491 (N_11491,N_9819,N_9890);
nor U11492 (N_11492,N_9428,N_9735);
xnor U11493 (N_11493,N_9955,N_10363);
or U11494 (N_11494,N_9982,N_9823);
and U11495 (N_11495,N_9039,N_10008);
xnor U11496 (N_11496,N_10219,N_9839);
or U11497 (N_11497,N_9821,N_9177);
xnor U11498 (N_11498,N_9603,N_10014);
and U11499 (N_11499,N_10078,N_9341);
nand U11500 (N_11500,N_9826,N_9263);
or U11501 (N_11501,N_9887,N_10236);
xor U11502 (N_11502,N_9174,N_9666);
and U11503 (N_11503,N_9316,N_9423);
and U11504 (N_11504,N_9848,N_9767);
xor U11505 (N_11505,N_9257,N_9321);
nand U11506 (N_11506,N_9430,N_9229);
nand U11507 (N_11507,N_9519,N_9509);
nand U11508 (N_11508,N_9904,N_9136);
nand U11509 (N_11509,N_9024,N_10131);
nand U11510 (N_11510,N_10093,N_10006);
and U11511 (N_11511,N_10103,N_9600);
xor U11512 (N_11512,N_10055,N_9251);
and U11513 (N_11513,N_9201,N_9098);
and U11514 (N_11514,N_10243,N_10053);
and U11515 (N_11515,N_9112,N_10163);
and U11516 (N_11516,N_9129,N_9917);
or U11517 (N_11517,N_10287,N_10398);
nor U11518 (N_11518,N_9281,N_10265);
nor U11519 (N_11519,N_10281,N_10414);
nand U11520 (N_11520,N_9024,N_9665);
nor U11521 (N_11521,N_9102,N_9922);
nand U11522 (N_11522,N_9752,N_10079);
and U11523 (N_11523,N_10285,N_9296);
nand U11524 (N_11524,N_9954,N_9878);
xor U11525 (N_11525,N_9615,N_9085);
and U11526 (N_11526,N_9607,N_10208);
xnor U11527 (N_11527,N_9390,N_9383);
or U11528 (N_11528,N_9236,N_9864);
nand U11529 (N_11529,N_10433,N_10280);
or U11530 (N_11530,N_10173,N_9934);
or U11531 (N_11531,N_10388,N_9113);
nor U11532 (N_11532,N_9349,N_9472);
nand U11533 (N_11533,N_10072,N_9198);
nor U11534 (N_11534,N_9960,N_9351);
xor U11535 (N_11535,N_9873,N_9211);
xnor U11536 (N_11536,N_9830,N_9219);
or U11537 (N_11537,N_10060,N_9426);
nand U11538 (N_11538,N_9116,N_9817);
nor U11539 (N_11539,N_10114,N_9768);
and U11540 (N_11540,N_9282,N_10422);
or U11541 (N_11541,N_10086,N_10238);
nand U11542 (N_11542,N_9327,N_9440);
and U11543 (N_11543,N_9249,N_9458);
or U11544 (N_11544,N_9477,N_9442);
and U11545 (N_11545,N_10390,N_10009);
or U11546 (N_11546,N_9123,N_9221);
or U11547 (N_11547,N_9315,N_9502);
xor U11548 (N_11548,N_9305,N_9182);
and U11549 (N_11549,N_9139,N_9381);
xnor U11550 (N_11550,N_10338,N_9746);
or U11551 (N_11551,N_9782,N_9700);
nand U11552 (N_11552,N_10131,N_10312);
or U11553 (N_11553,N_9947,N_9560);
nor U11554 (N_11554,N_9194,N_9902);
nand U11555 (N_11555,N_10442,N_10235);
nor U11556 (N_11556,N_10012,N_9000);
or U11557 (N_11557,N_10126,N_10430);
nor U11558 (N_11558,N_10007,N_9530);
and U11559 (N_11559,N_9422,N_9056);
xor U11560 (N_11560,N_10179,N_9393);
or U11561 (N_11561,N_9244,N_10023);
nor U11562 (N_11562,N_9289,N_9225);
or U11563 (N_11563,N_9859,N_9113);
and U11564 (N_11564,N_9943,N_10212);
xnor U11565 (N_11565,N_9209,N_9321);
and U11566 (N_11566,N_10033,N_10483);
nor U11567 (N_11567,N_9432,N_9029);
nor U11568 (N_11568,N_9018,N_9289);
or U11569 (N_11569,N_9475,N_10280);
xnor U11570 (N_11570,N_9551,N_9377);
xor U11571 (N_11571,N_9424,N_9091);
or U11572 (N_11572,N_10409,N_10287);
xor U11573 (N_11573,N_10195,N_10348);
or U11574 (N_11574,N_9638,N_9508);
xnor U11575 (N_11575,N_10335,N_10464);
and U11576 (N_11576,N_9357,N_9813);
nor U11577 (N_11577,N_10140,N_9076);
nor U11578 (N_11578,N_10231,N_9298);
nor U11579 (N_11579,N_9155,N_10304);
nor U11580 (N_11580,N_10313,N_9484);
xnor U11581 (N_11581,N_9434,N_9822);
or U11582 (N_11582,N_9936,N_10238);
nor U11583 (N_11583,N_9388,N_9575);
xor U11584 (N_11584,N_10075,N_9638);
nand U11585 (N_11585,N_10246,N_9399);
and U11586 (N_11586,N_10311,N_9371);
and U11587 (N_11587,N_9203,N_9289);
or U11588 (N_11588,N_10063,N_10296);
nand U11589 (N_11589,N_10307,N_9242);
nand U11590 (N_11590,N_9001,N_10213);
nand U11591 (N_11591,N_9980,N_9214);
and U11592 (N_11592,N_9666,N_9403);
xor U11593 (N_11593,N_10226,N_9002);
or U11594 (N_11594,N_9009,N_9596);
nand U11595 (N_11595,N_10393,N_9071);
nor U11596 (N_11596,N_9904,N_9514);
and U11597 (N_11597,N_10081,N_9582);
or U11598 (N_11598,N_9308,N_9812);
nand U11599 (N_11599,N_9391,N_9148);
nand U11600 (N_11600,N_9864,N_9831);
nor U11601 (N_11601,N_10095,N_9497);
and U11602 (N_11602,N_10446,N_9383);
or U11603 (N_11603,N_10274,N_10070);
and U11604 (N_11604,N_10349,N_9250);
or U11605 (N_11605,N_10329,N_9933);
and U11606 (N_11606,N_10121,N_10473);
and U11607 (N_11607,N_10470,N_9175);
xnor U11608 (N_11608,N_10162,N_9657);
nor U11609 (N_11609,N_10096,N_9697);
xor U11610 (N_11610,N_10179,N_9619);
nor U11611 (N_11611,N_10163,N_10246);
or U11612 (N_11612,N_9824,N_9531);
nand U11613 (N_11613,N_9453,N_9886);
xor U11614 (N_11614,N_10361,N_9048);
nand U11615 (N_11615,N_9894,N_9376);
nand U11616 (N_11616,N_10267,N_9556);
or U11617 (N_11617,N_9468,N_10444);
or U11618 (N_11618,N_10212,N_9220);
or U11619 (N_11619,N_9297,N_9147);
nand U11620 (N_11620,N_10499,N_10290);
or U11621 (N_11621,N_10203,N_9152);
nor U11622 (N_11622,N_9657,N_9361);
nand U11623 (N_11623,N_9030,N_9048);
or U11624 (N_11624,N_9914,N_9625);
or U11625 (N_11625,N_9577,N_9509);
nand U11626 (N_11626,N_10346,N_10084);
nand U11627 (N_11627,N_9128,N_9163);
and U11628 (N_11628,N_10226,N_10242);
or U11629 (N_11629,N_9641,N_10322);
xnor U11630 (N_11630,N_10371,N_9607);
or U11631 (N_11631,N_9230,N_10468);
or U11632 (N_11632,N_10332,N_9955);
and U11633 (N_11633,N_10403,N_9475);
xor U11634 (N_11634,N_9952,N_9017);
nand U11635 (N_11635,N_10042,N_9449);
or U11636 (N_11636,N_10260,N_9793);
nand U11637 (N_11637,N_9578,N_9648);
nor U11638 (N_11638,N_9650,N_9540);
nor U11639 (N_11639,N_9964,N_9374);
xnor U11640 (N_11640,N_9076,N_9878);
nand U11641 (N_11641,N_9457,N_9705);
or U11642 (N_11642,N_9386,N_9193);
or U11643 (N_11643,N_9869,N_9271);
nand U11644 (N_11644,N_9713,N_9794);
and U11645 (N_11645,N_10068,N_9469);
nor U11646 (N_11646,N_9998,N_10486);
nand U11647 (N_11647,N_10222,N_10272);
nand U11648 (N_11648,N_9101,N_9146);
xnor U11649 (N_11649,N_9570,N_10364);
nor U11650 (N_11650,N_9258,N_9340);
nand U11651 (N_11651,N_10166,N_10234);
nand U11652 (N_11652,N_9732,N_9706);
or U11653 (N_11653,N_10004,N_10268);
xnor U11654 (N_11654,N_10316,N_10471);
and U11655 (N_11655,N_9610,N_9037);
nand U11656 (N_11656,N_10247,N_10371);
nor U11657 (N_11657,N_9116,N_10458);
and U11658 (N_11658,N_10047,N_10291);
nor U11659 (N_11659,N_10380,N_9345);
xnor U11660 (N_11660,N_10296,N_9486);
nor U11661 (N_11661,N_9139,N_9062);
or U11662 (N_11662,N_9923,N_10314);
nand U11663 (N_11663,N_10271,N_10132);
or U11664 (N_11664,N_9044,N_10071);
nor U11665 (N_11665,N_9401,N_9254);
xnor U11666 (N_11666,N_10216,N_9590);
or U11667 (N_11667,N_9427,N_10042);
nand U11668 (N_11668,N_9590,N_10061);
xor U11669 (N_11669,N_9204,N_9271);
or U11670 (N_11670,N_9058,N_10027);
and U11671 (N_11671,N_9256,N_10335);
nor U11672 (N_11672,N_9890,N_9603);
or U11673 (N_11673,N_9365,N_9711);
nand U11674 (N_11674,N_9037,N_10361);
nor U11675 (N_11675,N_10163,N_9740);
nand U11676 (N_11676,N_9998,N_9480);
xnor U11677 (N_11677,N_9167,N_9049);
nand U11678 (N_11678,N_9359,N_9955);
nand U11679 (N_11679,N_10122,N_9163);
nor U11680 (N_11680,N_9960,N_9068);
xor U11681 (N_11681,N_10187,N_9362);
or U11682 (N_11682,N_9942,N_10263);
nor U11683 (N_11683,N_9364,N_9780);
or U11684 (N_11684,N_9465,N_9127);
and U11685 (N_11685,N_9932,N_9333);
and U11686 (N_11686,N_10292,N_10263);
or U11687 (N_11687,N_10085,N_10462);
nor U11688 (N_11688,N_9080,N_9248);
nor U11689 (N_11689,N_9744,N_9411);
and U11690 (N_11690,N_9690,N_9480);
and U11691 (N_11691,N_10400,N_10060);
nor U11692 (N_11692,N_9318,N_9016);
xor U11693 (N_11693,N_10450,N_9111);
nor U11694 (N_11694,N_10085,N_9142);
or U11695 (N_11695,N_9145,N_10360);
nand U11696 (N_11696,N_9177,N_10447);
xor U11697 (N_11697,N_9618,N_9466);
nor U11698 (N_11698,N_9584,N_9652);
xor U11699 (N_11699,N_9446,N_9894);
and U11700 (N_11700,N_9625,N_9093);
and U11701 (N_11701,N_9216,N_10015);
nand U11702 (N_11702,N_9962,N_9287);
nand U11703 (N_11703,N_9707,N_9029);
nor U11704 (N_11704,N_10486,N_9810);
nand U11705 (N_11705,N_9968,N_9191);
xnor U11706 (N_11706,N_9391,N_10480);
and U11707 (N_11707,N_9201,N_9912);
xor U11708 (N_11708,N_9290,N_9775);
xor U11709 (N_11709,N_9146,N_9752);
nand U11710 (N_11710,N_10255,N_9281);
xor U11711 (N_11711,N_9178,N_10210);
xor U11712 (N_11712,N_9682,N_10475);
nor U11713 (N_11713,N_9063,N_9229);
and U11714 (N_11714,N_9759,N_9217);
xnor U11715 (N_11715,N_9365,N_9034);
nor U11716 (N_11716,N_9493,N_9694);
xnor U11717 (N_11717,N_10069,N_9668);
xnor U11718 (N_11718,N_10099,N_9428);
and U11719 (N_11719,N_9465,N_9806);
or U11720 (N_11720,N_9526,N_9458);
nand U11721 (N_11721,N_10209,N_9390);
nor U11722 (N_11722,N_10361,N_9349);
xnor U11723 (N_11723,N_9701,N_10431);
or U11724 (N_11724,N_9741,N_9229);
xor U11725 (N_11725,N_10231,N_9400);
or U11726 (N_11726,N_9214,N_10434);
and U11727 (N_11727,N_9853,N_10222);
nand U11728 (N_11728,N_9988,N_10234);
nand U11729 (N_11729,N_9904,N_9433);
nand U11730 (N_11730,N_9937,N_9105);
or U11731 (N_11731,N_10439,N_10056);
nor U11732 (N_11732,N_10171,N_9388);
xnor U11733 (N_11733,N_10285,N_9070);
xor U11734 (N_11734,N_9731,N_10219);
nor U11735 (N_11735,N_10059,N_10411);
xnor U11736 (N_11736,N_9281,N_10359);
and U11737 (N_11737,N_10262,N_9867);
xnor U11738 (N_11738,N_9709,N_10049);
xnor U11739 (N_11739,N_9700,N_10483);
nor U11740 (N_11740,N_9468,N_10338);
nor U11741 (N_11741,N_10229,N_9026);
and U11742 (N_11742,N_10017,N_10175);
nand U11743 (N_11743,N_9118,N_9919);
nand U11744 (N_11744,N_10169,N_9658);
and U11745 (N_11745,N_9858,N_9979);
nand U11746 (N_11746,N_10189,N_10230);
xor U11747 (N_11747,N_10445,N_9476);
xnor U11748 (N_11748,N_9337,N_10132);
nand U11749 (N_11749,N_9321,N_9174);
nor U11750 (N_11750,N_9794,N_10070);
nand U11751 (N_11751,N_9166,N_9889);
xor U11752 (N_11752,N_9924,N_9099);
xnor U11753 (N_11753,N_10446,N_9216);
nand U11754 (N_11754,N_9644,N_9477);
or U11755 (N_11755,N_9936,N_9869);
nand U11756 (N_11756,N_9591,N_9121);
xnor U11757 (N_11757,N_9909,N_9332);
or U11758 (N_11758,N_10289,N_9956);
or U11759 (N_11759,N_9972,N_9189);
or U11760 (N_11760,N_9488,N_9127);
nand U11761 (N_11761,N_9116,N_9944);
xor U11762 (N_11762,N_9745,N_9005);
and U11763 (N_11763,N_10450,N_9020);
or U11764 (N_11764,N_9901,N_9865);
or U11765 (N_11765,N_9188,N_9580);
nor U11766 (N_11766,N_9352,N_9983);
or U11767 (N_11767,N_9291,N_10150);
and U11768 (N_11768,N_9968,N_9058);
xor U11769 (N_11769,N_10292,N_10403);
nor U11770 (N_11770,N_9312,N_9435);
or U11771 (N_11771,N_9546,N_9955);
nand U11772 (N_11772,N_10195,N_9446);
nor U11773 (N_11773,N_9457,N_9644);
nand U11774 (N_11774,N_10190,N_9581);
xnor U11775 (N_11775,N_9389,N_9363);
or U11776 (N_11776,N_9793,N_9101);
nor U11777 (N_11777,N_10275,N_9286);
nor U11778 (N_11778,N_9102,N_9736);
nor U11779 (N_11779,N_10284,N_9561);
nor U11780 (N_11780,N_10422,N_9023);
nand U11781 (N_11781,N_9363,N_9745);
xnor U11782 (N_11782,N_9552,N_9015);
nor U11783 (N_11783,N_9032,N_9372);
nand U11784 (N_11784,N_10292,N_9170);
nor U11785 (N_11785,N_10393,N_9327);
xor U11786 (N_11786,N_9804,N_10050);
xor U11787 (N_11787,N_9987,N_10072);
and U11788 (N_11788,N_10174,N_9255);
nand U11789 (N_11789,N_10340,N_9421);
and U11790 (N_11790,N_10434,N_9501);
xor U11791 (N_11791,N_9566,N_9139);
nor U11792 (N_11792,N_9365,N_9839);
or U11793 (N_11793,N_10170,N_10361);
and U11794 (N_11794,N_10190,N_10030);
or U11795 (N_11795,N_10030,N_9002);
nor U11796 (N_11796,N_9001,N_9415);
nor U11797 (N_11797,N_9045,N_10237);
nor U11798 (N_11798,N_10362,N_10423);
xor U11799 (N_11799,N_10357,N_9506);
or U11800 (N_11800,N_9428,N_9380);
nand U11801 (N_11801,N_10143,N_10433);
or U11802 (N_11802,N_9838,N_10467);
or U11803 (N_11803,N_9763,N_9965);
and U11804 (N_11804,N_9970,N_9502);
nand U11805 (N_11805,N_9485,N_10068);
xnor U11806 (N_11806,N_9552,N_10139);
and U11807 (N_11807,N_9248,N_9734);
and U11808 (N_11808,N_10442,N_9386);
nand U11809 (N_11809,N_9347,N_9296);
nor U11810 (N_11810,N_10277,N_10439);
and U11811 (N_11811,N_9703,N_10427);
nor U11812 (N_11812,N_9004,N_9761);
nand U11813 (N_11813,N_9374,N_9415);
nor U11814 (N_11814,N_9267,N_10031);
nor U11815 (N_11815,N_10206,N_9142);
nor U11816 (N_11816,N_9861,N_9922);
xor U11817 (N_11817,N_9379,N_10316);
and U11818 (N_11818,N_10370,N_9894);
and U11819 (N_11819,N_10482,N_9583);
or U11820 (N_11820,N_9116,N_10181);
or U11821 (N_11821,N_9886,N_9455);
nand U11822 (N_11822,N_9748,N_10225);
nand U11823 (N_11823,N_9819,N_9157);
nor U11824 (N_11824,N_9275,N_9119);
nor U11825 (N_11825,N_10057,N_9925);
xnor U11826 (N_11826,N_9947,N_10050);
nand U11827 (N_11827,N_9982,N_10277);
and U11828 (N_11828,N_10431,N_10114);
nor U11829 (N_11829,N_10058,N_9754);
or U11830 (N_11830,N_10211,N_9954);
xor U11831 (N_11831,N_9043,N_10405);
nand U11832 (N_11832,N_9284,N_9433);
nand U11833 (N_11833,N_9842,N_10136);
nor U11834 (N_11834,N_9890,N_9439);
and U11835 (N_11835,N_10377,N_9171);
nor U11836 (N_11836,N_10387,N_9563);
or U11837 (N_11837,N_9483,N_9148);
nand U11838 (N_11838,N_10255,N_10155);
or U11839 (N_11839,N_10458,N_9227);
nand U11840 (N_11840,N_9627,N_9239);
nand U11841 (N_11841,N_9764,N_9602);
nand U11842 (N_11842,N_9928,N_9329);
or U11843 (N_11843,N_10446,N_9788);
xor U11844 (N_11844,N_10080,N_10421);
and U11845 (N_11845,N_9402,N_9307);
nand U11846 (N_11846,N_10406,N_9552);
nor U11847 (N_11847,N_9241,N_9844);
nand U11848 (N_11848,N_10068,N_9217);
xnor U11849 (N_11849,N_9738,N_10155);
nor U11850 (N_11850,N_9832,N_9931);
and U11851 (N_11851,N_10408,N_10463);
xnor U11852 (N_11852,N_9894,N_9229);
nand U11853 (N_11853,N_9635,N_9566);
xnor U11854 (N_11854,N_10109,N_10431);
and U11855 (N_11855,N_9379,N_9624);
and U11856 (N_11856,N_9971,N_9282);
xnor U11857 (N_11857,N_9796,N_9812);
nor U11858 (N_11858,N_9876,N_9365);
and U11859 (N_11859,N_9519,N_9073);
xor U11860 (N_11860,N_9995,N_10371);
and U11861 (N_11861,N_10216,N_9725);
nand U11862 (N_11862,N_9990,N_9735);
nor U11863 (N_11863,N_9731,N_10393);
or U11864 (N_11864,N_10091,N_9136);
xor U11865 (N_11865,N_9401,N_9061);
nor U11866 (N_11866,N_10055,N_10218);
nand U11867 (N_11867,N_10376,N_9573);
and U11868 (N_11868,N_10375,N_10301);
or U11869 (N_11869,N_9298,N_9613);
xnor U11870 (N_11870,N_9929,N_9640);
and U11871 (N_11871,N_10449,N_10458);
nand U11872 (N_11872,N_10023,N_9660);
nor U11873 (N_11873,N_10103,N_10139);
nand U11874 (N_11874,N_10214,N_10320);
nand U11875 (N_11875,N_9289,N_9087);
xor U11876 (N_11876,N_9883,N_9060);
or U11877 (N_11877,N_9414,N_9089);
xnor U11878 (N_11878,N_10451,N_9036);
or U11879 (N_11879,N_10254,N_9333);
and U11880 (N_11880,N_9272,N_9460);
nand U11881 (N_11881,N_9641,N_9533);
or U11882 (N_11882,N_9456,N_9346);
and U11883 (N_11883,N_9941,N_9692);
nand U11884 (N_11884,N_10087,N_9882);
nor U11885 (N_11885,N_10160,N_9817);
nor U11886 (N_11886,N_9701,N_9248);
and U11887 (N_11887,N_9275,N_10025);
nand U11888 (N_11888,N_9237,N_9284);
nor U11889 (N_11889,N_9999,N_9640);
or U11890 (N_11890,N_10056,N_9265);
xor U11891 (N_11891,N_9826,N_9588);
nand U11892 (N_11892,N_9749,N_9018);
nor U11893 (N_11893,N_10043,N_10194);
or U11894 (N_11894,N_10453,N_9795);
xnor U11895 (N_11895,N_10372,N_10363);
and U11896 (N_11896,N_9250,N_9572);
nor U11897 (N_11897,N_9704,N_9853);
nor U11898 (N_11898,N_9108,N_9120);
nand U11899 (N_11899,N_9347,N_10240);
or U11900 (N_11900,N_9771,N_9835);
or U11901 (N_11901,N_9983,N_9458);
and U11902 (N_11902,N_10111,N_9624);
xnor U11903 (N_11903,N_9266,N_9064);
or U11904 (N_11904,N_9623,N_10263);
and U11905 (N_11905,N_9645,N_10470);
nor U11906 (N_11906,N_9073,N_10205);
and U11907 (N_11907,N_10102,N_10131);
nand U11908 (N_11908,N_9242,N_9858);
xnor U11909 (N_11909,N_9515,N_9729);
nor U11910 (N_11910,N_9977,N_10060);
xnor U11911 (N_11911,N_10227,N_10175);
and U11912 (N_11912,N_9619,N_9388);
or U11913 (N_11913,N_10272,N_10466);
or U11914 (N_11914,N_9657,N_10424);
xor U11915 (N_11915,N_10273,N_9305);
xor U11916 (N_11916,N_9612,N_9821);
and U11917 (N_11917,N_10003,N_9213);
xor U11918 (N_11918,N_9604,N_9255);
or U11919 (N_11919,N_10080,N_9092);
nor U11920 (N_11920,N_10010,N_10058);
or U11921 (N_11921,N_9767,N_10036);
or U11922 (N_11922,N_10020,N_10286);
xnor U11923 (N_11923,N_9779,N_9576);
xnor U11924 (N_11924,N_9795,N_9811);
and U11925 (N_11925,N_10237,N_10338);
xor U11926 (N_11926,N_9599,N_9802);
nand U11927 (N_11927,N_9631,N_9176);
nor U11928 (N_11928,N_10377,N_10490);
xor U11929 (N_11929,N_9393,N_9717);
nor U11930 (N_11930,N_10399,N_10368);
nor U11931 (N_11931,N_9369,N_9291);
xor U11932 (N_11932,N_9718,N_9957);
and U11933 (N_11933,N_10128,N_9251);
or U11934 (N_11934,N_9337,N_9458);
nand U11935 (N_11935,N_10090,N_9770);
and U11936 (N_11936,N_9423,N_9165);
nand U11937 (N_11937,N_9520,N_9330);
and U11938 (N_11938,N_9347,N_9481);
nand U11939 (N_11939,N_9287,N_9686);
xor U11940 (N_11940,N_10101,N_9504);
or U11941 (N_11941,N_10040,N_9343);
nor U11942 (N_11942,N_9836,N_9222);
or U11943 (N_11943,N_10197,N_10126);
xor U11944 (N_11944,N_9622,N_9956);
or U11945 (N_11945,N_10333,N_10382);
xor U11946 (N_11946,N_9998,N_10476);
xor U11947 (N_11947,N_10130,N_9422);
xnor U11948 (N_11948,N_9543,N_10077);
nand U11949 (N_11949,N_10140,N_10332);
xnor U11950 (N_11950,N_9277,N_9000);
and U11951 (N_11951,N_9174,N_10321);
xor U11952 (N_11952,N_9002,N_10060);
or U11953 (N_11953,N_9422,N_10097);
xor U11954 (N_11954,N_9473,N_10114);
nor U11955 (N_11955,N_10262,N_9642);
nand U11956 (N_11956,N_9997,N_10108);
or U11957 (N_11957,N_9466,N_9006);
xor U11958 (N_11958,N_9050,N_9423);
or U11959 (N_11959,N_9487,N_10322);
nor U11960 (N_11960,N_10003,N_9770);
xor U11961 (N_11961,N_10074,N_9721);
or U11962 (N_11962,N_9000,N_10089);
or U11963 (N_11963,N_10445,N_9496);
and U11964 (N_11964,N_9304,N_9864);
xnor U11965 (N_11965,N_9763,N_10285);
xnor U11966 (N_11966,N_9151,N_9467);
or U11967 (N_11967,N_9834,N_10155);
nand U11968 (N_11968,N_9709,N_9889);
nand U11969 (N_11969,N_10225,N_9525);
nand U11970 (N_11970,N_10365,N_9835);
nor U11971 (N_11971,N_9808,N_10338);
or U11972 (N_11972,N_10266,N_9156);
and U11973 (N_11973,N_9718,N_9412);
and U11974 (N_11974,N_10032,N_9102);
nor U11975 (N_11975,N_9485,N_9745);
or U11976 (N_11976,N_9722,N_9977);
nor U11977 (N_11977,N_10222,N_9286);
and U11978 (N_11978,N_10403,N_9881);
nand U11979 (N_11979,N_9801,N_10319);
or U11980 (N_11980,N_10004,N_9055);
nand U11981 (N_11981,N_9608,N_10091);
nand U11982 (N_11982,N_9529,N_10408);
nor U11983 (N_11983,N_10217,N_9625);
or U11984 (N_11984,N_9451,N_9929);
or U11985 (N_11985,N_9204,N_9466);
and U11986 (N_11986,N_9710,N_9489);
or U11987 (N_11987,N_9519,N_10437);
nand U11988 (N_11988,N_9645,N_9237);
or U11989 (N_11989,N_9307,N_10345);
nor U11990 (N_11990,N_10051,N_9004);
nor U11991 (N_11991,N_9546,N_9427);
or U11992 (N_11992,N_9058,N_10065);
nand U11993 (N_11993,N_9073,N_9969);
and U11994 (N_11994,N_9962,N_10204);
xor U11995 (N_11995,N_10453,N_10403);
xor U11996 (N_11996,N_9665,N_9232);
nand U11997 (N_11997,N_9572,N_9517);
nor U11998 (N_11998,N_9953,N_9382);
nor U11999 (N_11999,N_10458,N_9339);
xor U12000 (N_12000,N_11335,N_11338);
or U12001 (N_12001,N_10518,N_11392);
and U12002 (N_12002,N_11267,N_11479);
nor U12003 (N_12003,N_10760,N_11975);
nand U12004 (N_12004,N_11353,N_11913);
xor U12005 (N_12005,N_10539,N_11684);
nand U12006 (N_12006,N_11596,N_11163);
xnor U12007 (N_12007,N_11258,N_11145);
and U12008 (N_12008,N_10975,N_10746);
xnor U12009 (N_12009,N_10784,N_10998);
and U12010 (N_12010,N_11079,N_11412);
or U12011 (N_12011,N_10946,N_11370);
xnor U12012 (N_12012,N_10620,N_11047);
or U12013 (N_12013,N_10502,N_10675);
or U12014 (N_12014,N_11589,N_10773);
xnor U12015 (N_12015,N_11577,N_10642);
and U12016 (N_12016,N_11890,N_11033);
and U12017 (N_12017,N_11942,N_11151);
xnor U12018 (N_12018,N_11808,N_11509);
and U12019 (N_12019,N_11055,N_11778);
and U12020 (N_12020,N_11834,N_10990);
or U12021 (N_12021,N_10657,N_10622);
nand U12022 (N_12022,N_11679,N_11631);
nor U12023 (N_12023,N_11235,N_11226);
xnor U12024 (N_12024,N_11248,N_11739);
or U12025 (N_12025,N_11358,N_11899);
nand U12026 (N_12026,N_10526,N_11460);
xnor U12027 (N_12027,N_10651,N_11557);
nand U12028 (N_12028,N_11422,N_11617);
nor U12029 (N_12029,N_10611,N_11597);
nor U12030 (N_12030,N_10879,N_11581);
xor U12031 (N_12031,N_11371,N_11906);
or U12032 (N_12032,N_11575,N_11578);
or U12033 (N_12033,N_11819,N_10796);
and U12034 (N_12034,N_11315,N_10633);
nor U12035 (N_12035,N_11729,N_10818);
nand U12036 (N_12036,N_10677,N_11757);
nand U12037 (N_12037,N_11065,N_11489);
nor U12038 (N_12038,N_10598,N_11918);
or U12039 (N_12039,N_11718,N_11636);
xor U12040 (N_12040,N_10788,N_10789);
nor U12041 (N_12041,N_11020,N_11482);
and U12042 (N_12042,N_10577,N_11302);
nand U12043 (N_12043,N_11749,N_11635);
xor U12044 (N_12044,N_10954,N_11524);
and U12045 (N_12045,N_11949,N_11139);
nor U12046 (N_12046,N_11814,N_10972);
or U12047 (N_12047,N_10889,N_11579);
nand U12048 (N_12048,N_10810,N_11584);
or U12049 (N_12049,N_11947,N_10585);
or U12050 (N_12050,N_11205,N_11376);
xnor U12051 (N_12051,N_10872,N_10700);
nand U12052 (N_12052,N_11735,N_11936);
nor U12053 (N_12053,N_11399,N_11468);
xnor U12054 (N_12054,N_11332,N_11326);
nor U12055 (N_12055,N_11884,N_10586);
nor U12056 (N_12056,N_11062,N_11471);
nor U12057 (N_12057,N_11415,N_11212);
nand U12058 (N_12058,N_10776,N_11637);
or U12059 (N_12059,N_10676,N_11278);
or U12060 (N_12060,N_11916,N_10926);
nand U12061 (N_12061,N_10531,N_11229);
or U12062 (N_12062,N_11880,N_10716);
nand U12063 (N_12063,N_11061,N_11621);
xor U12064 (N_12064,N_11955,N_10942);
xor U12065 (N_12065,N_11765,N_11303);
nor U12066 (N_12066,N_11238,N_11296);
nand U12067 (N_12067,N_11200,N_10823);
xnor U12068 (N_12068,N_11064,N_10659);
nor U12069 (N_12069,N_11364,N_10909);
xor U12070 (N_12070,N_11943,N_11649);
nand U12071 (N_12071,N_11246,N_11701);
and U12072 (N_12072,N_11395,N_11845);
nor U12073 (N_12073,N_11381,N_10956);
nand U12074 (N_12074,N_11904,N_11158);
xnor U12075 (N_12075,N_10519,N_11807);
nor U12076 (N_12076,N_11506,N_11515);
and U12077 (N_12077,N_10530,N_10532);
and U12078 (N_12078,N_10898,N_10547);
and U12079 (N_12079,N_10664,N_10825);
xor U12080 (N_12080,N_11223,N_11888);
and U12081 (N_12081,N_11723,N_11003);
or U12082 (N_12082,N_11365,N_10793);
and U12083 (N_12083,N_11241,N_11012);
xor U12084 (N_12084,N_10635,N_10573);
and U12085 (N_12085,N_11944,N_11245);
nand U12086 (N_12086,N_11754,N_11776);
xor U12087 (N_12087,N_11492,N_10875);
or U12088 (N_12088,N_11292,N_11962);
or U12089 (N_12089,N_10874,N_11623);
nor U12090 (N_12090,N_11646,N_11774);
nor U12091 (N_12091,N_10999,N_11091);
nor U12092 (N_12092,N_11184,N_11606);
nand U12093 (N_12093,N_10609,N_10572);
xnor U12094 (N_12094,N_11678,N_11447);
and U12095 (N_12095,N_11901,N_10738);
and U12096 (N_12096,N_10978,N_11772);
nor U12097 (N_12097,N_11634,N_10636);
xor U12098 (N_12098,N_11831,N_11115);
or U12099 (N_12099,N_11762,N_11505);
and U12100 (N_12100,N_11112,N_10578);
nand U12101 (N_12101,N_11101,N_10625);
and U12102 (N_12102,N_10890,N_11963);
nand U12103 (N_12103,N_11743,N_11816);
nor U12104 (N_12104,N_11499,N_10994);
and U12105 (N_12105,N_11144,N_11086);
or U12106 (N_12106,N_11340,N_10720);
nand U12107 (N_12107,N_10691,N_10543);
nor U12108 (N_12108,N_11030,N_11025);
nor U12109 (N_12109,N_10535,N_10771);
and U12110 (N_12110,N_11465,N_10802);
nand U12111 (N_12111,N_10882,N_11582);
or U12112 (N_12112,N_10589,N_11361);
xor U12113 (N_12113,N_11952,N_11941);
or U12114 (N_12114,N_11263,N_11806);
and U12115 (N_12115,N_11549,N_11734);
or U12116 (N_12116,N_10919,N_11789);
nor U12117 (N_12117,N_11357,N_11601);
or U12118 (N_12118,N_11454,N_11847);
nand U12119 (N_12119,N_11491,N_11408);
nand U12120 (N_12120,N_10571,N_11493);
and U12121 (N_12121,N_11536,N_10637);
xnor U12122 (N_12122,N_10912,N_11313);
or U12123 (N_12123,N_10721,N_11985);
and U12124 (N_12124,N_11174,N_11182);
and U12125 (N_12125,N_11935,N_11045);
or U12126 (N_12126,N_10991,N_11771);
nand U12127 (N_12127,N_11930,N_11574);
nor U12128 (N_12128,N_10932,N_11783);
and U12129 (N_12129,N_11374,N_11852);
nand U12130 (N_12130,N_11910,N_11194);
or U12131 (N_12131,N_11630,N_11432);
nand U12132 (N_12132,N_11879,N_11948);
nand U12133 (N_12133,N_11472,N_11450);
or U12134 (N_12134,N_10517,N_11481);
nand U12135 (N_12135,N_10834,N_10768);
or U12136 (N_12136,N_10566,N_10618);
or U12137 (N_12137,N_11274,N_10648);
nor U12138 (N_12138,N_10910,N_11236);
nand U12139 (N_12139,N_11198,N_11530);
or U12140 (N_12140,N_11002,N_10590);
or U12141 (N_12141,N_11976,N_10613);
and U12142 (N_12142,N_10682,N_11680);
or U12143 (N_12143,N_11440,N_10866);
or U12144 (N_12144,N_11853,N_10701);
nand U12145 (N_12145,N_11893,N_11484);
xor U12146 (N_12146,N_10629,N_11475);
and U12147 (N_12147,N_11915,N_11925);
nand U12148 (N_12148,N_10923,N_11339);
nand U12149 (N_12149,N_11034,N_11953);
nor U12150 (N_12150,N_11529,N_10544);
nor U12151 (N_12151,N_11160,N_11697);
or U12152 (N_12152,N_11728,N_11560);
and U12153 (N_12153,N_11161,N_11257);
nor U12154 (N_12154,N_10827,N_10928);
and U12155 (N_12155,N_10698,N_11812);
or U12156 (N_12156,N_11827,N_10982);
nand U12157 (N_12157,N_10709,N_10714);
nor U12158 (N_12158,N_11037,N_10971);
nand U12159 (N_12159,N_10908,N_11396);
xor U12160 (N_12160,N_11090,N_10934);
and U12161 (N_12161,N_11222,N_11561);
nor U12162 (N_12162,N_11881,N_11685);
nand U12163 (N_12163,N_11978,N_10688);
and U12164 (N_12164,N_11638,N_10754);
and U12165 (N_12165,N_11049,N_10557);
nand U12166 (N_12166,N_10901,N_10729);
xnor U12167 (N_12167,N_10570,N_10948);
nand U12168 (N_12168,N_11923,N_10937);
nand U12169 (N_12169,N_10758,N_11767);
and U12170 (N_12170,N_11240,N_10766);
or U12171 (N_12171,N_11874,N_10945);
nand U12172 (N_12172,N_11427,N_11883);
nand U12173 (N_12173,N_10608,N_11871);
or U12174 (N_12174,N_11297,N_11074);
and U12175 (N_12175,N_10761,N_11331);
and U12176 (N_12176,N_11995,N_10895);
nand U12177 (N_12177,N_10512,N_10896);
xnor U12178 (N_12178,N_10681,N_11780);
nand U12179 (N_12179,N_11805,N_11689);
xnor U12180 (N_12180,N_10851,N_11096);
nor U12181 (N_12181,N_11615,N_11155);
xor U12182 (N_12182,N_11394,N_10616);
or U12183 (N_12183,N_11398,N_11262);
xor U12184 (N_12184,N_11154,N_10941);
xor U12185 (N_12185,N_11945,N_11193);
or U12186 (N_12186,N_11775,N_10985);
xor U12187 (N_12187,N_11233,N_11627);
nor U12188 (N_12188,N_11732,N_11616);
xnor U12189 (N_12189,N_11736,N_10816);
nand U12190 (N_12190,N_11900,N_11875);
nor U12191 (N_12191,N_11157,N_11379);
nand U12192 (N_12192,N_10638,N_10778);
xnor U12193 (N_12193,N_11803,N_10787);
and U12194 (N_12194,N_10737,N_10567);
nand U12195 (N_12195,N_11021,N_11826);
nor U12196 (N_12196,N_11169,N_10696);
or U12197 (N_12197,N_11330,N_10838);
xor U12198 (N_12198,N_11537,N_10870);
xor U12199 (N_12199,N_11197,N_11362);
nor U12200 (N_12200,N_11372,N_10809);
nand U12201 (N_12201,N_10563,N_10974);
or U12202 (N_12202,N_11368,N_11603);
or U12203 (N_12203,N_11420,N_11019);
nor U12204 (N_12204,N_11657,N_11230);
nor U12205 (N_12205,N_11719,N_11971);
and U12206 (N_12206,N_10580,N_11063);
or U12207 (N_12207,N_11797,N_11703);
nand U12208 (N_12208,N_11406,N_11609);
or U12209 (N_12209,N_11266,N_11428);
nand U12210 (N_12210,N_10894,N_10981);
or U12211 (N_12211,N_11760,N_10905);
or U12212 (N_12212,N_10992,N_11221);
and U12213 (N_12213,N_10538,N_11443);
and U12214 (N_12214,N_10917,N_10646);
and U12215 (N_12215,N_11289,N_11958);
or U12216 (N_12216,N_11629,N_11706);
and U12217 (N_12217,N_10943,N_11419);
xnor U12218 (N_12218,N_11401,N_11591);
and U12219 (N_12219,N_10630,N_10808);
nor U12220 (N_12220,N_11547,N_11452);
nor U12221 (N_12221,N_11625,N_10755);
nor U12222 (N_12222,N_11043,N_10631);
or U12223 (N_12223,N_10846,N_10840);
or U12224 (N_12224,N_10939,N_11269);
and U12225 (N_12225,N_11015,N_11494);
or U12226 (N_12226,N_11572,N_10730);
and U12227 (N_12227,N_10645,N_11698);
or U12228 (N_12228,N_11983,N_11177);
nor U12229 (N_12229,N_11640,N_11960);
or U12230 (N_12230,N_11093,N_10607);
nor U12231 (N_12231,N_11252,N_10509);
xnor U12232 (N_12232,N_11299,N_11510);
nand U12233 (N_12233,N_10899,N_11533);
xor U12234 (N_12234,N_11288,N_11334);
and U12235 (N_12235,N_10938,N_11987);
nand U12236 (N_12236,N_11310,N_10892);
or U12237 (N_12237,N_11018,N_10710);
xnor U12238 (N_12238,N_11521,N_11458);
nand U12239 (N_12239,N_11275,N_11946);
and U12240 (N_12240,N_11084,N_11868);
or U12241 (N_12241,N_11416,N_11414);
xnor U12242 (N_12242,N_11192,N_11683);
nor U12243 (N_12243,N_10891,N_10548);
xnor U12244 (N_12244,N_10833,N_10627);
nor U12245 (N_12245,N_11988,N_10961);
and U12246 (N_12246,N_11191,N_10516);
nand U12247 (N_12247,N_10952,N_10558);
xnor U12248 (N_12248,N_11742,N_10826);
nor U12249 (N_12249,N_11350,N_11932);
and U12250 (N_12250,N_11470,N_10705);
xor U12251 (N_12251,N_11598,N_10759);
xnor U12252 (N_12252,N_10718,N_10575);
nand U12253 (N_12253,N_11451,N_10782);
and U12254 (N_12254,N_11761,N_11060);
nand U12255 (N_12255,N_11804,N_11309);
nand U12256 (N_12256,N_11463,N_10503);
nor U12257 (N_12257,N_11608,N_10545);
nand U12258 (N_12258,N_11066,N_11426);
nor U12259 (N_12259,N_11840,N_11039);
and U12260 (N_12260,N_10853,N_11186);
or U12261 (N_12261,N_11858,N_11284);
xor U12262 (N_12262,N_11725,N_11125);
nor U12263 (N_12263,N_11702,N_11800);
and U12264 (N_12264,N_10756,N_11010);
and U12265 (N_12265,N_11891,N_11004);
nor U12266 (N_12266,N_11956,N_10753);
nor U12267 (N_12267,N_11367,N_11788);
xor U12268 (N_12268,N_11565,N_11854);
nor U12269 (N_12269,N_10960,N_11818);
nand U12270 (N_12270,N_10900,N_11820);
and U12271 (N_12271,N_11052,N_10614);
xnor U12272 (N_12272,N_11410,N_10731);
nor U12273 (N_12273,N_11176,N_11977);
nand U12274 (N_12274,N_11234,N_10967);
nand U12275 (N_12275,N_11795,N_11828);
or U12276 (N_12276,N_10528,N_11078);
and U12277 (N_12277,N_10769,N_11153);
nand U12278 (N_12278,N_10862,N_11905);
nand U12279 (N_12279,N_11518,N_11279);
nand U12280 (N_12280,N_11994,N_11724);
xor U12281 (N_12281,N_11285,N_10565);
nor U12282 (N_12282,N_11516,N_11571);
xnor U12283 (N_12283,N_10977,N_11504);
nor U12284 (N_12284,N_11552,N_10887);
nand U12285 (N_12285,N_10918,N_11425);
and U12286 (N_12286,N_11914,N_11405);
or U12287 (N_12287,N_11855,N_10593);
and U12288 (N_12288,N_11005,N_11710);
xor U12289 (N_12289,N_11317,N_11423);
or U12290 (N_12290,N_11662,N_11912);
xnor U12291 (N_12291,N_11903,N_11573);
and U12292 (N_12292,N_10727,N_10581);
and U12293 (N_12293,N_11986,N_11534);
nand U12294 (N_12294,N_11369,N_10876);
nand U12295 (N_12295,N_10711,N_11342);
nand U12296 (N_12296,N_10678,N_11261);
or U12297 (N_12297,N_10806,N_10799);
xnor U12298 (N_12298,N_11967,N_11558);
and U12299 (N_12299,N_11437,N_10924);
nor U12300 (N_12300,N_10829,N_10790);
nor U12301 (N_12301,N_10674,N_10973);
nor U12302 (N_12302,N_11907,N_10549);
nand U12303 (N_12303,N_11250,N_10881);
nor U12304 (N_12304,N_11276,N_10821);
and U12305 (N_12305,N_11188,N_11894);
nor U12306 (N_12306,N_10725,N_10582);
xnor U12307 (N_12307,N_11103,N_11794);
nor U12308 (N_12308,N_11919,N_11528);
and U12309 (N_12309,N_10656,N_11270);
or U12310 (N_12310,N_11273,N_11337);
nor U12311 (N_12311,N_10594,N_11383);
nand U12312 (N_12312,N_11098,N_10508);
nor U12313 (N_12313,N_11487,N_11641);
or U12314 (N_12314,N_11300,N_11210);
and U12315 (N_12315,N_11730,N_10968);
nor U12316 (N_12316,N_10736,N_11654);
or U12317 (N_12317,N_11700,N_10949);
and U12318 (N_12318,N_11889,N_11922);
nand U12319 (N_12319,N_10830,N_10979);
or U12320 (N_12320,N_11622,N_11802);
and U12321 (N_12321,N_10950,N_10868);
nor U12322 (N_12322,N_11308,N_11787);
nand U12323 (N_12323,N_11291,N_11108);
or U12324 (N_12324,N_11072,N_11319);
or U12325 (N_12325,N_11691,N_11109);
xnor U12326 (N_12326,N_10715,N_10860);
or U12327 (N_12327,N_11931,N_11860);
or U12328 (N_12328,N_11295,N_11570);
nor U12329 (N_12329,N_10723,N_11307);
xnor U12330 (N_12330,N_11146,N_11653);
and U12331 (N_12331,N_10770,N_10963);
nand U12332 (N_12332,N_10525,N_11954);
xor U12333 (N_12333,N_11864,N_11551);
nand U12334 (N_12334,N_11469,N_11642);
or U12335 (N_12335,N_11522,N_11605);
xnor U12336 (N_12336,N_11567,N_10842);
or U12337 (N_12337,N_11007,N_10728);
or U12338 (N_12338,N_11793,N_11445);
and U12339 (N_12339,N_10597,N_11073);
nand U12340 (N_12340,N_11542,N_11283);
nand U12341 (N_12341,N_11546,N_10740);
xnor U12342 (N_12342,N_10683,N_11850);
nand U12343 (N_12343,N_11027,N_11607);
and U12344 (N_12344,N_10667,N_11999);
or U12345 (N_12345,N_11206,N_11321);
or U12346 (N_12346,N_11175,N_10831);
xnor U12347 (N_12347,N_11569,N_11838);
nand U12348 (N_12348,N_11696,N_10820);
xnor U12349 (N_12349,N_11782,N_10680);
or U12350 (N_12350,N_11990,N_11260);
and U12351 (N_12351,N_10692,N_10837);
xor U12352 (N_12352,N_11247,N_11859);
or U12353 (N_12353,N_11937,N_11934);
xnor U12354 (N_12354,N_10739,N_11333);
or U12355 (N_12355,N_11989,N_10743);
xor U12356 (N_12356,N_11791,N_10704);
and U12357 (N_12357,N_11254,N_10596);
xor U12358 (N_12358,N_11122,N_11737);
or U12359 (N_12359,N_11069,N_10907);
and U12360 (N_12360,N_11950,N_11179);
or U12361 (N_12361,N_11213,N_11189);
nand U12362 (N_12362,N_10653,N_11298);
nand U12363 (N_12363,N_11556,N_11766);
xor U12364 (N_12364,N_11924,N_11346);
nor U12365 (N_12365,N_11202,N_11111);
nor U12366 (N_12366,N_11592,N_10673);
xnor U12367 (N_12367,N_11526,N_10933);
xnor U12368 (N_12368,N_10989,N_11017);
xnor U12369 (N_12369,N_11866,N_10987);
or U12370 (N_12370,N_11253,N_11835);
xnor U12371 (N_12371,N_11271,N_10764);
or U12372 (N_12372,N_11436,N_10897);
xor U12373 (N_12373,N_10884,N_11391);
or U12374 (N_12374,N_11418,N_11779);
nor U12375 (N_12375,N_11323,N_11159);
nand U12376 (N_12376,N_11360,N_10588);
and U12377 (N_12377,N_11409,N_10970);
nand U12378 (N_12378,N_11809,N_11190);
xor U12379 (N_12379,N_10551,N_11466);
xor U12380 (N_12380,N_11135,N_10561);
nand U12381 (N_12381,N_11659,N_11585);
and U12382 (N_12382,N_11377,N_11704);
or U12383 (N_12383,N_11844,N_11555);
xnor U12384 (N_12384,N_10822,N_11455);
or U12385 (N_12385,N_10914,N_10592);
and U12386 (N_12386,N_10867,N_11686);
xnor U12387 (N_12387,N_11476,N_11563);
or U12388 (N_12388,N_11215,N_11882);
nand U12389 (N_12389,N_11224,N_11676);
nand U12390 (N_12390,N_11513,N_10813);
xor U12391 (N_12391,N_11650,N_11119);
nand U12392 (N_12392,N_10552,N_10958);
nand U12393 (N_12393,N_10812,N_11023);
nor U12394 (N_12394,N_10925,N_11277);
xnor U12395 (N_12395,N_11041,N_10886);
or U12396 (N_12396,N_11752,N_11525);
xnor U12397 (N_12397,N_10523,N_11969);
nor U12398 (N_12398,N_11645,N_10836);
xnor U12399 (N_12399,N_11687,N_11682);
xor U12400 (N_12400,N_11344,N_10878);
or U12401 (N_12401,N_11926,N_11327);
nand U12402 (N_12402,N_10719,N_11712);
nand U12403 (N_12403,N_11128,N_11441);
nor U12404 (N_12404,N_11624,N_11424);
xnor U12405 (N_12405,N_11272,N_10670);
or U12406 (N_12406,N_11902,N_11070);
and U12407 (N_12407,N_11094,N_10540);
nor U12408 (N_12408,N_11130,N_10861);
xor U12409 (N_12409,N_11322,N_10672);
nand U12410 (N_12410,N_11026,N_10612);
xor U12411 (N_12411,N_11957,N_10717);
nor U12412 (N_12412,N_11731,N_11439);
xor U12413 (N_12413,N_10640,N_11548);
nand U12414 (N_12414,N_11660,N_11527);
nand U12415 (N_12415,N_11137,N_11965);
nand U12416 (N_12416,N_11051,N_11628);
xnor U12417 (N_12417,N_11610,N_10668);
and U12418 (N_12418,N_11036,N_10584);
xnor U12419 (N_12419,N_11755,N_11927);
nor U12420 (N_12420,N_10835,N_10639);
and U12421 (N_12421,N_11397,N_11196);
and U12422 (N_12422,N_10841,N_11456);
xor U12423 (N_12423,N_10983,N_11973);
nor U12424 (N_12424,N_11974,N_10996);
nand U12425 (N_12425,N_10805,N_11359);
and U12426 (N_12426,N_10559,N_10795);
nand U12427 (N_12427,N_10751,N_11669);
xnor U12428 (N_12428,N_11448,N_11824);
or U12429 (N_12429,N_11336,N_10767);
nand U12430 (N_12430,N_11403,N_11014);
nor U12431 (N_12431,N_10888,N_10986);
and U12432 (N_12432,N_11633,N_10786);
xor U12433 (N_12433,N_11486,N_11038);
nor U12434 (N_12434,N_11329,N_11770);
nor U12435 (N_12435,N_11393,N_11172);
nor U12436 (N_12436,N_11741,N_11328);
nor U12437 (N_12437,N_11693,N_11588);
nor U12438 (N_12438,N_11217,N_10576);
nand U12439 (N_12439,N_10747,N_11675);
nand U12440 (N_12440,N_10930,N_11016);
and U12441 (N_12441,N_11520,N_11162);
or U12442 (N_12442,N_11228,N_11758);
xnor U12443 (N_12443,N_10520,N_11166);
xnor U12444 (N_12444,N_11707,N_11892);
and U12445 (N_12445,N_11259,N_11594);
nand U12446 (N_12446,N_11059,N_11022);
nor U12447 (N_12447,N_11180,N_11001);
or U12448 (N_12448,N_10783,N_11738);
nor U12449 (N_12449,N_10703,N_10797);
nand U12450 (N_12450,N_11239,N_10828);
xor U12451 (N_12451,N_11717,N_11165);
or U12452 (N_12452,N_11237,N_10944);
nand U12453 (N_12453,N_11961,N_11639);
or U12454 (N_12454,N_11540,N_11201);
or U12455 (N_12455,N_11343,N_10864);
or U12456 (N_12456,N_11535,N_10906);
xnor U12457 (N_12457,N_11863,N_11048);
nor U12458 (N_12458,N_10921,N_11709);
nor U12459 (N_12459,N_10643,N_11265);
nor U12460 (N_12460,N_11773,N_11281);
nand U12461 (N_12461,N_11611,N_10904);
nor U12462 (N_12462,N_11187,N_10858);
nor U12463 (N_12463,N_11595,N_11673);
or U12464 (N_12464,N_11242,N_10601);
xnor U12465 (N_12465,N_11825,N_11671);
nand U12466 (N_12466,N_10685,N_10615);
or U12467 (N_12467,N_11227,N_11543);
or U12468 (N_12468,N_11681,N_10560);
nor U12469 (N_12469,N_11387,N_11668);
and U12470 (N_12470,N_11304,N_10936);
nor U12471 (N_12471,N_10505,N_10969);
and U12472 (N_12472,N_11388,N_11796);
nor U12473 (N_12473,N_10724,N_10521);
nor U12474 (N_12474,N_10619,N_11028);
or U12475 (N_12475,N_11148,N_11363);
nor U12476 (N_12476,N_11088,N_11356);
nor U12477 (N_12477,N_10605,N_11720);
or U12478 (N_12478,N_11841,N_10628);
xnor U12479 (N_12479,N_11559,N_11851);
nand U12480 (N_12480,N_10697,N_11209);
nand U12481 (N_12481,N_11823,N_11785);
or U12482 (N_12482,N_11068,N_10569);
nand U12483 (N_12483,N_10712,N_10626);
xor U12484 (N_12484,N_11694,N_10562);
xor U12485 (N_12485,N_10621,N_11740);
nand U12486 (N_12486,N_10966,N_11120);
and U12487 (N_12487,N_11982,N_10686);
nand U12488 (N_12488,N_10763,N_10785);
xor U12489 (N_12489,N_10995,N_11656);
and U12490 (N_12490,N_11386,N_11769);
xnor U12491 (N_12491,N_11077,N_11920);
nor U12492 (N_12492,N_11620,N_11433);
nand U12493 (N_12493,N_11488,N_11677);
or U12494 (N_12494,N_11220,N_11964);
nor U12495 (N_12495,N_10857,N_10568);
or U12496 (N_12496,N_11507,N_11121);
or U12497 (N_12497,N_11100,N_11618);
or U12498 (N_12498,N_11008,N_11517);
xnor U12499 (N_12499,N_11286,N_10684);
xnor U12500 (N_12500,N_11117,N_11856);
nor U12501 (N_12501,N_11873,N_10903);
nand U12502 (N_12502,N_11544,N_10687);
nor U12503 (N_12503,N_11294,N_11417);
or U12504 (N_12504,N_11462,N_11290);
nor U12505 (N_12505,N_11389,N_11080);
nor U12506 (N_12506,N_11786,N_10722);
nand U12507 (N_12507,N_11106,N_11981);
nor U12508 (N_12508,N_11496,N_11566);
xor U12509 (N_12509,N_10980,N_11614);
and U12510 (N_12510,N_10955,N_11050);
nand U12511 (N_12511,N_11870,N_11503);
or U12512 (N_12512,N_11590,N_11404);
and U12513 (N_12513,N_11243,N_11695);
xnor U12514 (N_12514,N_11539,N_10541);
xor U12515 (N_12515,N_11046,N_11626);
and U12516 (N_12516,N_11508,N_11171);
and U12517 (N_12517,N_11349,N_11057);
nor U12518 (N_12518,N_11256,N_11421);
xor U12519 (N_12519,N_11532,N_10515);
and U12520 (N_12520,N_10735,N_11013);
or U12521 (N_12521,N_11714,N_11756);
and U12522 (N_12522,N_11593,N_11341);
nor U12523 (N_12523,N_11619,N_11127);
nor U12524 (N_12524,N_11612,N_10811);
nor U12525 (N_12525,N_11876,N_11413);
nor U12526 (N_12526,N_10777,N_10775);
nor U12527 (N_12527,N_10603,N_10665);
nand U12528 (N_12528,N_11054,N_11836);
xnor U12529 (N_12529,N_11861,N_10533);
or U12530 (N_12530,N_11087,N_11843);
nor U12531 (N_12531,N_10997,N_11390);
xnor U12532 (N_12532,N_10550,N_10644);
or U12533 (N_12533,N_11991,N_10732);
xnor U12534 (N_12534,N_10847,N_11867);
or U12535 (N_12535,N_10663,N_11658);
and U12536 (N_12536,N_11970,N_11464);
xor U12537 (N_12537,N_10623,N_11129);
xor U12538 (N_12538,N_10965,N_11402);
nand U12539 (N_12539,N_11538,N_11777);
xor U12540 (N_12540,N_10880,N_11784);
nor U12541 (N_12541,N_10655,N_11147);
nand U12542 (N_12542,N_11280,N_11104);
and U12543 (N_12543,N_11181,N_11705);
nand U12544 (N_12544,N_10750,N_11293);
nor U12545 (N_12545,N_11502,N_10885);
xnor U12546 (N_12546,N_11480,N_11651);
and U12547 (N_12547,N_11798,N_10781);
xnor U12548 (N_12548,N_11282,N_10591);
xor U12549 (N_12549,N_11959,N_11810);
xnor U12550 (N_12550,N_11301,N_10742);
xor U12551 (N_12551,N_11156,N_11311);
nor U12552 (N_12552,N_11211,N_10817);
nand U12553 (N_12553,N_10902,N_10602);
xnor U12554 (N_12554,N_10947,N_10511);
xnor U12555 (N_12555,N_11219,N_11721);
and U12556 (N_12556,N_11848,N_10844);
or U12557 (N_12557,N_11750,N_11126);
or U12558 (N_12558,N_10957,N_11746);
or U12559 (N_12559,N_11268,N_10660);
or U12560 (N_12560,N_10632,N_11670);
or U12561 (N_12561,N_11152,N_11692);
nand U12562 (N_12562,N_10600,N_11664);
and U12563 (N_12563,N_11216,N_10929);
xnor U12564 (N_12564,N_10706,N_11136);
nand U12565 (N_12565,N_11652,N_11715);
xnor U12566 (N_12566,N_11461,N_11887);
nand U12567 (N_12567,N_10815,N_11583);
or U12568 (N_12568,N_10606,N_11457);
and U12569 (N_12569,N_10839,N_10658);
xnor U12570 (N_12570,N_11966,N_11324);
xor U12571 (N_12571,N_11314,N_11497);
nor U12572 (N_12572,N_10679,N_11763);
nand U12573 (N_12573,N_11495,N_10931);
xor U12574 (N_12574,N_11655,N_11431);
and U12575 (N_12575,N_10599,N_11477);
nor U12576 (N_12576,N_10537,N_11208);
xor U12577 (N_12577,N_11554,N_10666);
and U12578 (N_12578,N_11821,N_10734);
and U12579 (N_12579,N_11075,N_10953);
and U12580 (N_12580,N_11107,N_11105);
nand U12581 (N_12581,N_11602,N_11058);
nand U12582 (N_12582,N_10506,N_11799);
xnor U12583 (N_12583,N_11790,N_11511);
or U12584 (N_12584,N_11997,N_11114);
or U12585 (N_12585,N_10848,N_11131);
nand U12586 (N_12586,N_11951,N_11917);
xnor U12587 (N_12587,N_10819,N_11143);
xor U12588 (N_12588,N_11781,N_11095);
nor U12589 (N_12589,N_10927,N_11822);
or U12590 (N_12590,N_11811,N_11564);
xnor U12591 (N_12591,N_10852,N_11124);
xnor U12592 (N_12592,N_11312,N_10873);
nand U12593 (N_12593,N_11035,N_11024);
and U12594 (N_12594,N_11325,N_11613);
nand U12595 (N_12595,N_11897,N_11523);
nand U12596 (N_12596,N_10792,N_11708);
xor U12597 (N_12597,N_10748,N_10555);
and U12598 (N_12598,N_11133,N_10513);
and U12599 (N_12599,N_11672,N_11138);
nand U12600 (N_12600,N_11199,N_11815);
nand U12601 (N_12601,N_10801,N_11663);
nor U12602 (N_12602,N_11751,N_10922);
nand U12603 (N_12603,N_11753,N_10757);
xnor U12604 (N_12604,N_11722,N_10534);
nand U12605 (N_12605,N_11429,N_11674);
and U12606 (N_12606,N_11102,N_10869);
nor U12607 (N_12607,N_10574,N_10850);
xor U12608 (N_12608,N_11378,N_11099);
xnor U12609 (N_12609,N_10661,N_11142);
xnor U12610 (N_12610,N_11562,N_10845);
or U12611 (N_12611,N_10617,N_11647);
nor U12612 (N_12612,N_10610,N_11085);
nand U12613 (N_12613,N_10604,N_11580);
xnor U12614 (N_12614,N_10504,N_10522);
or U12615 (N_12615,N_10553,N_11711);
or U12616 (N_12616,N_11839,N_11661);
xor U12617 (N_12617,N_10690,N_10807);
or U12618 (N_12618,N_10652,N_10527);
xnor U12619 (N_12619,N_10595,N_10556);
or U12620 (N_12620,N_10699,N_10749);
or U12621 (N_12621,N_11909,N_11195);
nor U12622 (N_12622,N_11173,N_11716);
nor U12623 (N_12623,N_11204,N_11167);
or U12624 (N_12624,N_10859,N_11053);
or U12625 (N_12625,N_10976,N_10649);
nor U12626 (N_12626,N_11744,N_11643);
or U12627 (N_12627,N_10579,N_10984);
and U12628 (N_12628,N_11031,N_11632);
xnor U12629 (N_12629,N_10865,N_11885);
nand U12630 (N_12630,N_10536,N_11832);
and U12631 (N_12631,N_11097,N_11170);
xnor U12632 (N_12632,N_11928,N_10694);
and U12633 (N_12633,N_11898,N_11972);
or U12634 (N_12634,N_11110,N_11490);
and U12635 (N_12635,N_10744,N_10951);
nand U12636 (N_12636,N_11768,N_10702);
nand U12637 (N_12637,N_10689,N_11287);
xor U12638 (N_12638,N_10871,N_11857);
and U12639 (N_12639,N_11519,N_11141);
and U12640 (N_12640,N_11713,N_11531);
xor U12641 (N_12641,N_11225,N_11667);
nand U12642 (N_12642,N_11232,N_10856);
nor U12643 (N_12643,N_11541,N_10708);
and U12644 (N_12644,N_11599,N_11373);
nor U12645 (N_12645,N_11348,N_11459);
and U12646 (N_12646,N_10507,N_11029);
nand U12647 (N_12647,N_11116,N_10843);
nor U12648 (N_12648,N_10824,N_11185);
nand U12649 (N_12649,N_11747,N_10920);
nor U12650 (N_12650,N_11553,N_10916);
or U12651 (N_12651,N_10940,N_10741);
and U12652 (N_12652,N_11407,N_10962);
nor U12653 (N_12653,N_11690,N_11846);
nor U12654 (N_12654,N_10794,N_10500);
and U12655 (N_12655,N_11183,N_10762);
nand U12656 (N_12656,N_11214,N_11355);
and U12657 (N_12657,N_11305,N_11231);
and U12658 (N_12658,N_11911,N_10647);
xnor U12659 (N_12659,N_11968,N_11076);
nor U12660 (N_12660,N_10911,N_11586);
xor U12661 (N_12661,N_11453,N_11501);
xnor U12662 (N_12662,N_11438,N_11842);
or U12663 (N_12663,N_10913,N_11092);
xnor U12664 (N_12664,N_11837,N_11938);
or U12665 (N_12665,N_11665,N_11032);
nand U12666 (N_12666,N_11044,N_11000);
nor U12667 (N_12667,N_11089,N_11320);
xor U12668 (N_12668,N_11474,N_11168);
xor U12669 (N_12669,N_11498,N_11984);
xor U12670 (N_12670,N_10669,N_10671);
or U12671 (N_12671,N_11568,N_11666);
nand U12672 (N_12672,N_11829,N_10514);
or U12673 (N_12673,N_11587,N_11434);
or U12674 (N_12674,N_11869,N_11132);
xor U12675 (N_12675,N_10814,N_10524);
xnor U12676 (N_12676,N_11813,N_10624);
xnor U12677 (N_12677,N_10893,N_11056);
xnor U12678 (N_12678,N_11347,N_11366);
and U12679 (N_12679,N_11733,N_10765);
or U12680 (N_12680,N_11446,N_11249);
nor U12681 (N_12681,N_11382,N_10772);
xor U12682 (N_12682,N_10542,N_11545);
nand U12683 (N_12683,N_10752,N_11400);
or U12684 (N_12684,N_10855,N_10662);
or U12685 (N_12685,N_11473,N_10713);
or U12686 (N_12686,N_11726,N_11082);
nand U12687 (N_12687,N_11878,N_11745);
and U12688 (N_12688,N_11896,N_10959);
xnor U12689 (N_12689,N_11040,N_11998);
or U12690 (N_12690,N_11550,N_11251);
xor U12691 (N_12691,N_10745,N_10695);
or U12692 (N_12692,N_11699,N_11067);
or U12693 (N_12693,N_11354,N_10935);
and U12694 (N_12694,N_10650,N_10915);
and U12695 (N_12695,N_11764,N_10587);
or U12696 (N_12696,N_11877,N_11375);
or U12697 (N_12697,N_11071,N_11600);
or U12698 (N_12698,N_11644,N_11921);
and U12699 (N_12699,N_11123,N_11442);
and U12700 (N_12700,N_11042,N_11939);
xor U12701 (N_12701,N_11908,N_11318);
nand U12702 (N_12702,N_11979,N_10501);
xnor U12703 (N_12703,N_11385,N_11255);
nor U12704 (N_12704,N_10849,N_10564);
xnor U12705 (N_12705,N_11164,N_11980);
or U12706 (N_12706,N_10832,N_11009);
nand U12707 (N_12707,N_10654,N_11748);
and U12708 (N_12708,N_10554,N_10791);
nor U12709 (N_12709,N_10883,N_11512);
xnor U12710 (N_12710,N_11244,N_11817);
xor U12711 (N_12711,N_11011,N_11895);
or U12712 (N_12712,N_11849,N_10693);
xnor U12713 (N_12713,N_11478,N_10733);
and U12714 (N_12714,N_11865,N_11306);
nor U12715 (N_12715,N_10583,N_11345);
xnor U12716 (N_12716,N_11203,N_11485);
nor U12717 (N_12717,N_11576,N_10529);
or U12718 (N_12718,N_11648,N_10877);
or U12719 (N_12719,N_11149,N_10774);
xnor U12720 (N_12720,N_11872,N_10804);
nand U12721 (N_12721,N_11933,N_10798);
and U12722 (N_12722,N_11449,N_11688);
nand U12723 (N_12723,N_11113,N_11083);
or U12724 (N_12724,N_11929,N_11801);
and U12725 (N_12725,N_11430,N_11444);
or U12726 (N_12726,N_10988,N_11264);
or U12727 (N_12727,N_11940,N_11380);
nand U12728 (N_12728,N_10779,N_11604);
xnor U12729 (N_12729,N_11886,N_11514);
xnor U12730 (N_12730,N_11140,N_10707);
nor U12731 (N_12731,N_11150,N_11316);
nor U12732 (N_12732,N_11351,N_10510);
nand U12733 (N_12733,N_10546,N_11006);
nor U12734 (N_12734,N_11134,N_11500);
nand U12735 (N_12735,N_11996,N_11830);
and U12736 (N_12736,N_11178,N_10800);
or U12737 (N_12737,N_11727,N_10993);
or U12738 (N_12738,N_10854,N_11862);
xor U12739 (N_12739,N_11384,N_11207);
and U12740 (N_12740,N_11792,N_11411);
nor U12741 (N_12741,N_11759,N_11833);
xnor U12742 (N_12742,N_11118,N_11992);
nand U12743 (N_12743,N_11483,N_11081);
xnor U12744 (N_12744,N_10641,N_11467);
xor U12745 (N_12745,N_11218,N_11352);
nand U12746 (N_12746,N_10634,N_10726);
and U12747 (N_12747,N_10964,N_11993);
or U12748 (N_12748,N_10803,N_10863);
or U12749 (N_12749,N_11435,N_10780);
nand U12750 (N_12750,N_11330,N_10654);
xor U12751 (N_12751,N_11559,N_10817);
nand U12752 (N_12752,N_11011,N_10994);
nand U12753 (N_12753,N_11544,N_10825);
nand U12754 (N_12754,N_11271,N_11073);
xor U12755 (N_12755,N_10706,N_11873);
xor U12756 (N_12756,N_11952,N_10600);
nand U12757 (N_12757,N_11763,N_10973);
nand U12758 (N_12758,N_11570,N_11666);
nand U12759 (N_12759,N_11282,N_11885);
xnor U12760 (N_12760,N_10673,N_11914);
xor U12761 (N_12761,N_11725,N_11854);
and U12762 (N_12762,N_11745,N_11545);
xnor U12763 (N_12763,N_10902,N_11333);
nor U12764 (N_12764,N_11774,N_11508);
and U12765 (N_12765,N_11440,N_11672);
xnor U12766 (N_12766,N_11745,N_11974);
nand U12767 (N_12767,N_11685,N_10870);
and U12768 (N_12768,N_10595,N_11859);
nor U12769 (N_12769,N_11207,N_11792);
nor U12770 (N_12770,N_11098,N_11653);
nand U12771 (N_12771,N_10768,N_11679);
and U12772 (N_12772,N_10729,N_11287);
nand U12773 (N_12773,N_10740,N_11494);
or U12774 (N_12774,N_10961,N_11370);
or U12775 (N_12775,N_11485,N_10509);
nand U12776 (N_12776,N_11192,N_10941);
or U12777 (N_12777,N_11305,N_11218);
and U12778 (N_12778,N_11897,N_11878);
or U12779 (N_12779,N_11097,N_11678);
or U12780 (N_12780,N_11379,N_11847);
nor U12781 (N_12781,N_11316,N_10729);
or U12782 (N_12782,N_11691,N_11318);
and U12783 (N_12783,N_10902,N_10884);
nor U12784 (N_12784,N_11938,N_10881);
nand U12785 (N_12785,N_11629,N_10583);
and U12786 (N_12786,N_11049,N_11879);
and U12787 (N_12787,N_11617,N_11759);
and U12788 (N_12788,N_11721,N_11173);
nor U12789 (N_12789,N_11774,N_11316);
nand U12790 (N_12790,N_10926,N_10594);
xnor U12791 (N_12791,N_11320,N_11560);
or U12792 (N_12792,N_11249,N_11602);
nor U12793 (N_12793,N_10924,N_11932);
nor U12794 (N_12794,N_11428,N_10677);
or U12795 (N_12795,N_11825,N_10540);
or U12796 (N_12796,N_10932,N_10536);
nand U12797 (N_12797,N_11003,N_11071);
nor U12798 (N_12798,N_11423,N_10741);
and U12799 (N_12799,N_11435,N_11467);
xor U12800 (N_12800,N_11217,N_11543);
xor U12801 (N_12801,N_11455,N_10885);
nor U12802 (N_12802,N_11717,N_11381);
nand U12803 (N_12803,N_10521,N_10506);
nand U12804 (N_12804,N_11860,N_11617);
or U12805 (N_12805,N_11609,N_11118);
or U12806 (N_12806,N_10618,N_11737);
nor U12807 (N_12807,N_11598,N_11701);
nand U12808 (N_12808,N_11443,N_11332);
nand U12809 (N_12809,N_11958,N_11545);
nor U12810 (N_12810,N_11227,N_11008);
nor U12811 (N_12811,N_11693,N_11050);
nand U12812 (N_12812,N_10538,N_11863);
or U12813 (N_12813,N_10779,N_11329);
nand U12814 (N_12814,N_11718,N_11885);
or U12815 (N_12815,N_10711,N_11600);
nand U12816 (N_12816,N_11129,N_10663);
or U12817 (N_12817,N_10754,N_11965);
xor U12818 (N_12818,N_11695,N_10681);
nor U12819 (N_12819,N_10860,N_10725);
or U12820 (N_12820,N_11287,N_11788);
nand U12821 (N_12821,N_10859,N_11962);
nand U12822 (N_12822,N_10661,N_10537);
or U12823 (N_12823,N_10507,N_11373);
or U12824 (N_12824,N_11117,N_11597);
xor U12825 (N_12825,N_11567,N_11676);
nor U12826 (N_12826,N_10861,N_11162);
or U12827 (N_12827,N_11510,N_11440);
and U12828 (N_12828,N_10610,N_11241);
and U12829 (N_12829,N_10883,N_11886);
nand U12830 (N_12830,N_10734,N_10872);
or U12831 (N_12831,N_11565,N_11770);
xor U12832 (N_12832,N_10784,N_10854);
nand U12833 (N_12833,N_11020,N_11708);
nand U12834 (N_12834,N_11729,N_11105);
nand U12835 (N_12835,N_11422,N_11639);
nor U12836 (N_12836,N_11631,N_11798);
xnor U12837 (N_12837,N_11557,N_10532);
nand U12838 (N_12838,N_11229,N_10696);
or U12839 (N_12839,N_11812,N_10665);
xor U12840 (N_12840,N_11364,N_11243);
xor U12841 (N_12841,N_11929,N_11285);
and U12842 (N_12842,N_11820,N_11575);
nand U12843 (N_12843,N_10720,N_11006);
nor U12844 (N_12844,N_10851,N_10784);
xnor U12845 (N_12845,N_11370,N_11832);
and U12846 (N_12846,N_11990,N_11636);
nor U12847 (N_12847,N_11903,N_10787);
and U12848 (N_12848,N_11328,N_11591);
nand U12849 (N_12849,N_11233,N_11516);
xor U12850 (N_12850,N_10996,N_11898);
and U12851 (N_12851,N_10705,N_11798);
and U12852 (N_12852,N_11455,N_11770);
nor U12853 (N_12853,N_10826,N_11953);
nor U12854 (N_12854,N_10540,N_11415);
or U12855 (N_12855,N_11479,N_10983);
nor U12856 (N_12856,N_11374,N_10613);
nand U12857 (N_12857,N_11255,N_11022);
nand U12858 (N_12858,N_10642,N_10940);
nor U12859 (N_12859,N_11651,N_11174);
nand U12860 (N_12860,N_10662,N_11468);
nand U12861 (N_12861,N_11851,N_11748);
and U12862 (N_12862,N_11274,N_10663);
nand U12863 (N_12863,N_11344,N_11405);
and U12864 (N_12864,N_11759,N_10918);
and U12865 (N_12865,N_10716,N_11982);
nor U12866 (N_12866,N_11720,N_10583);
and U12867 (N_12867,N_11780,N_10731);
and U12868 (N_12868,N_11169,N_11210);
nor U12869 (N_12869,N_10680,N_11655);
xnor U12870 (N_12870,N_11814,N_11012);
nand U12871 (N_12871,N_11027,N_11805);
and U12872 (N_12872,N_10960,N_11246);
xnor U12873 (N_12873,N_10766,N_11719);
or U12874 (N_12874,N_11254,N_11125);
xnor U12875 (N_12875,N_10848,N_10816);
nor U12876 (N_12876,N_11950,N_11523);
xor U12877 (N_12877,N_10743,N_11187);
and U12878 (N_12878,N_10553,N_10876);
nor U12879 (N_12879,N_11730,N_11318);
or U12880 (N_12880,N_11822,N_11863);
or U12881 (N_12881,N_11766,N_11480);
and U12882 (N_12882,N_10782,N_11791);
nand U12883 (N_12883,N_11464,N_11002);
and U12884 (N_12884,N_10949,N_11548);
nand U12885 (N_12885,N_11633,N_10819);
nor U12886 (N_12886,N_11155,N_10769);
or U12887 (N_12887,N_11186,N_10722);
xnor U12888 (N_12888,N_11396,N_11808);
nor U12889 (N_12889,N_10524,N_11530);
nand U12890 (N_12890,N_10817,N_11405);
or U12891 (N_12891,N_10917,N_11481);
nor U12892 (N_12892,N_10887,N_10912);
xnor U12893 (N_12893,N_11449,N_11680);
xnor U12894 (N_12894,N_11796,N_11899);
xor U12895 (N_12895,N_11538,N_10777);
nand U12896 (N_12896,N_11857,N_10825);
xnor U12897 (N_12897,N_11602,N_11828);
nand U12898 (N_12898,N_11127,N_11494);
nor U12899 (N_12899,N_11174,N_11605);
and U12900 (N_12900,N_11811,N_11068);
xnor U12901 (N_12901,N_10864,N_11680);
nand U12902 (N_12902,N_10896,N_11016);
nor U12903 (N_12903,N_10503,N_11114);
nand U12904 (N_12904,N_10767,N_11748);
xor U12905 (N_12905,N_11455,N_11939);
nor U12906 (N_12906,N_11567,N_10511);
nand U12907 (N_12907,N_11529,N_11403);
nand U12908 (N_12908,N_11062,N_10726);
nand U12909 (N_12909,N_11754,N_11625);
or U12910 (N_12910,N_10986,N_10597);
nor U12911 (N_12911,N_11726,N_11292);
nand U12912 (N_12912,N_11277,N_10745);
or U12913 (N_12913,N_11810,N_11478);
nand U12914 (N_12914,N_11901,N_10739);
nor U12915 (N_12915,N_11675,N_11999);
and U12916 (N_12916,N_11289,N_11296);
xnor U12917 (N_12917,N_11170,N_10664);
nand U12918 (N_12918,N_11052,N_10720);
or U12919 (N_12919,N_10984,N_10560);
xor U12920 (N_12920,N_11045,N_10744);
or U12921 (N_12921,N_10697,N_11182);
nand U12922 (N_12922,N_11346,N_11842);
nand U12923 (N_12923,N_11135,N_11854);
or U12924 (N_12924,N_11664,N_11098);
nor U12925 (N_12925,N_11319,N_10989);
nand U12926 (N_12926,N_11992,N_11624);
nand U12927 (N_12927,N_11367,N_11674);
nor U12928 (N_12928,N_11470,N_11184);
xor U12929 (N_12929,N_11145,N_10891);
nor U12930 (N_12930,N_10885,N_11513);
and U12931 (N_12931,N_10893,N_11201);
and U12932 (N_12932,N_11242,N_11624);
and U12933 (N_12933,N_11656,N_11434);
nand U12934 (N_12934,N_11241,N_10547);
or U12935 (N_12935,N_11968,N_11414);
nand U12936 (N_12936,N_11236,N_11374);
xnor U12937 (N_12937,N_11387,N_10876);
or U12938 (N_12938,N_10673,N_10990);
nor U12939 (N_12939,N_11861,N_11087);
xnor U12940 (N_12940,N_11406,N_11500);
nor U12941 (N_12941,N_11199,N_11824);
nor U12942 (N_12942,N_10979,N_10599);
nand U12943 (N_12943,N_11313,N_11705);
and U12944 (N_12944,N_11844,N_11820);
xor U12945 (N_12945,N_11114,N_10730);
nor U12946 (N_12946,N_11709,N_11721);
nor U12947 (N_12947,N_10682,N_11185);
nor U12948 (N_12948,N_11790,N_10607);
and U12949 (N_12949,N_10828,N_11419);
and U12950 (N_12950,N_10920,N_11301);
nor U12951 (N_12951,N_10813,N_11148);
or U12952 (N_12952,N_11301,N_11053);
xnor U12953 (N_12953,N_11651,N_11629);
or U12954 (N_12954,N_10738,N_11052);
and U12955 (N_12955,N_11724,N_11530);
xnor U12956 (N_12956,N_11380,N_10510);
nor U12957 (N_12957,N_11887,N_11486);
xnor U12958 (N_12958,N_11013,N_11680);
and U12959 (N_12959,N_10791,N_11150);
xnor U12960 (N_12960,N_11222,N_11300);
xor U12961 (N_12961,N_10984,N_11435);
and U12962 (N_12962,N_11483,N_11813);
xnor U12963 (N_12963,N_11293,N_10594);
nand U12964 (N_12964,N_11490,N_10886);
xor U12965 (N_12965,N_10566,N_10766);
xnor U12966 (N_12966,N_11168,N_10804);
or U12967 (N_12967,N_11979,N_10745);
nor U12968 (N_12968,N_11599,N_10803);
nand U12969 (N_12969,N_11205,N_11984);
or U12970 (N_12970,N_11159,N_11497);
or U12971 (N_12971,N_11056,N_10855);
or U12972 (N_12972,N_11894,N_11921);
nand U12973 (N_12973,N_11380,N_11472);
and U12974 (N_12974,N_11597,N_11263);
nand U12975 (N_12975,N_11970,N_11607);
nor U12976 (N_12976,N_11313,N_11509);
or U12977 (N_12977,N_11219,N_11168);
nor U12978 (N_12978,N_11128,N_10904);
or U12979 (N_12979,N_10902,N_10898);
nand U12980 (N_12980,N_11538,N_11267);
and U12981 (N_12981,N_11483,N_11166);
and U12982 (N_12982,N_10757,N_11845);
nor U12983 (N_12983,N_11553,N_10962);
and U12984 (N_12984,N_10828,N_11317);
nor U12985 (N_12985,N_11967,N_11638);
nor U12986 (N_12986,N_10774,N_11028);
or U12987 (N_12987,N_10610,N_11508);
xnor U12988 (N_12988,N_11440,N_11638);
and U12989 (N_12989,N_11339,N_11545);
nor U12990 (N_12990,N_10581,N_10568);
nor U12991 (N_12991,N_10955,N_11153);
nor U12992 (N_12992,N_10818,N_10846);
xor U12993 (N_12993,N_11030,N_11834);
and U12994 (N_12994,N_11583,N_11588);
nor U12995 (N_12995,N_10546,N_11268);
nor U12996 (N_12996,N_11905,N_10658);
nor U12997 (N_12997,N_11870,N_10956);
nand U12998 (N_12998,N_10959,N_11569);
xor U12999 (N_12999,N_10928,N_10667);
and U13000 (N_13000,N_10792,N_11710);
and U13001 (N_13001,N_11113,N_11106);
xnor U13002 (N_13002,N_11550,N_11735);
or U13003 (N_13003,N_10957,N_11825);
or U13004 (N_13004,N_10502,N_10539);
or U13005 (N_13005,N_11441,N_11636);
and U13006 (N_13006,N_11118,N_10599);
xnor U13007 (N_13007,N_11163,N_11500);
nand U13008 (N_13008,N_11970,N_11197);
and U13009 (N_13009,N_11363,N_10748);
nand U13010 (N_13010,N_11200,N_11584);
and U13011 (N_13011,N_10516,N_10563);
and U13012 (N_13012,N_10918,N_10644);
xnor U13013 (N_13013,N_11304,N_10966);
and U13014 (N_13014,N_11006,N_11641);
or U13015 (N_13015,N_11911,N_11731);
or U13016 (N_13016,N_10788,N_10747);
and U13017 (N_13017,N_10806,N_11092);
or U13018 (N_13018,N_10572,N_11136);
nand U13019 (N_13019,N_10821,N_11037);
nor U13020 (N_13020,N_11834,N_11605);
or U13021 (N_13021,N_11712,N_10509);
nand U13022 (N_13022,N_10685,N_11066);
and U13023 (N_13023,N_11311,N_10904);
or U13024 (N_13024,N_11394,N_11771);
and U13025 (N_13025,N_11403,N_11001);
nor U13026 (N_13026,N_10811,N_11676);
xor U13027 (N_13027,N_11130,N_11140);
xnor U13028 (N_13028,N_11641,N_11501);
and U13029 (N_13029,N_10845,N_10616);
nand U13030 (N_13030,N_11805,N_10962);
nand U13031 (N_13031,N_11770,N_10929);
xor U13032 (N_13032,N_11507,N_11188);
nor U13033 (N_13033,N_11679,N_10535);
nand U13034 (N_13034,N_11509,N_10712);
xor U13035 (N_13035,N_10768,N_11970);
or U13036 (N_13036,N_11187,N_11148);
and U13037 (N_13037,N_11772,N_11333);
nor U13038 (N_13038,N_10608,N_10672);
nor U13039 (N_13039,N_11930,N_10658);
and U13040 (N_13040,N_11981,N_10685);
nand U13041 (N_13041,N_10500,N_11277);
xor U13042 (N_13042,N_11877,N_10813);
xor U13043 (N_13043,N_11054,N_11587);
nor U13044 (N_13044,N_10911,N_11740);
and U13045 (N_13045,N_11079,N_10928);
and U13046 (N_13046,N_11988,N_11098);
xor U13047 (N_13047,N_11057,N_11034);
xnor U13048 (N_13048,N_11516,N_10944);
xor U13049 (N_13049,N_11038,N_11099);
nor U13050 (N_13050,N_10849,N_11207);
nor U13051 (N_13051,N_11856,N_11078);
nor U13052 (N_13052,N_11231,N_11778);
or U13053 (N_13053,N_10542,N_11843);
and U13054 (N_13054,N_11325,N_11973);
and U13055 (N_13055,N_10732,N_10797);
and U13056 (N_13056,N_10779,N_10901);
nand U13057 (N_13057,N_11582,N_11327);
nor U13058 (N_13058,N_11296,N_11905);
nor U13059 (N_13059,N_11641,N_10706);
xnor U13060 (N_13060,N_11949,N_10611);
nand U13061 (N_13061,N_10972,N_11169);
and U13062 (N_13062,N_11778,N_10973);
and U13063 (N_13063,N_10992,N_11700);
xnor U13064 (N_13064,N_11155,N_10727);
and U13065 (N_13065,N_10630,N_11934);
nand U13066 (N_13066,N_11617,N_10628);
or U13067 (N_13067,N_11894,N_11609);
and U13068 (N_13068,N_11917,N_11255);
or U13069 (N_13069,N_11489,N_11067);
or U13070 (N_13070,N_11982,N_11540);
nor U13071 (N_13071,N_11408,N_10762);
nand U13072 (N_13072,N_11318,N_10506);
nor U13073 (N_13073,N_11693,N_10815);
and U13074 (N_13074,N_11853,N_10584);
xnor U13075 (N_13075,N_11772,N_11209);
xor U13076 (N_13076,N_11451,N_11320);
nor U13077 (N_13077,N_11426,N_11971);
nor U13078 (N_13078,N_11282,N_10967);
nand U13079 (N_13079,N_11033,N_10781);
nand U13080 (N_13080,N_11020,N_11539);
nand U13081 (N_13081,N_10989,N_11925);
nand U13082 (N_13082,N_10686,N_11698);
nand U13083 (N_13083,N_11707,N_11049);
nand U13084 (N_13084,N_11098,N_11579);
xnor U13085 (N_13085,N_10602,N_11341);
xnor U13086 (N_13086,N_11056,N_11809);
or U13087 (N_13087,N_11191,N_11038);
and U13088 (N_13088,N_11144,N_10533);
nor U13089 (N_13089,N_10633,N_11976);
and U13090 (N_13090,N_10897,N_11424);
xor U13091 (N_13091,N_11234,N_11980);
xor U13092 (N_13092,N_10704,N_11444);
nor U13093 (N_13093,N_10634,N_10794);
nor U13094 (N_13094,N_11057,N_10520);
or U13095 (N_13095,N_11299,N_10869);
nor U13096 (N_13096,N_10939,N_10839);
xor U13097 (N_13097,N_11175,N_11796);
and U13098 (N_13098,N_11135,N_10953);
or U13099 (N_13099,N_10936,N_10960);
and U13100 (N_13100,N_11042,N_11385);
nand U13101 (N_13101,N_10890,N_11689);
or U13102 (N_13102,N_11803,N_11359);
nor U13103 (N_13103,N_10635,N_11094);
nor U13104 (N_13104,N_11285,N_10620);
or U13105 (N_13105,N_11428,N_11002);
or U13106 (N_13106,N_10539,N_10547);
or U13107 (N_13107,N_11284,N_10705);
nand U13108 (N_13108,N_11350,N_11204);
and U13109 (N_13109,N_10528,N_11373);
and U13110 (N_13110,N_11710,N_11640);
and U13111 (N_13111,N_10812,N_11318);
nor U13112 (N_13112,N_10814,N_11955);
and U13113 (N_13113,N_11579,N_10663);
xor U13114 (N_13114,N_11518,N_11551);
xnor U13115 (N_13115,N_11682,N_10724);
nor U13116 (N_13116,N_10864,N_11198);
or U13117 (N_13117,N_11678,N_11144);
and U13118 (N_13118,N_10910,N_11100);
nand U13119 (N_13119,N_11824,N_11416);
nand U13120 (N_13120,N_10811,N_11606);
xnor U13121 (N_13121,N_10844,N_10948);
nor U13122 (N_13122,N_10782,N_11742);
nor U13123 (N_13123,N_11865,N_11353);
nand U13124 (N_13124,N_11600,N_10965);
nor U13125 (N_13125,N_10566,N_11345);
and U13126 (N_13126,N_11728,N_11301);
nor U13127 (N_13127,N_11244,N_11946);
and U13128 (N_13128,N_11266,N_11882);
nor U13129 (N_13129,N_10943,N_11134);
xnor U13130 (N_13130,N_11352,N_11423);
xor U13131 (N_13131,N_11762,N_10644);
nor U13132 (N_13132,N_11879,N_11064);
xnor U13133 (N_13133,N_10989,N_11636);
xor U13134 (N_13134,N_10507,N_11136);
nor U13135 (N_13135,N_10844,N_10764);
nand U13136 (N_13136,N_11828,N_10662);
and U13137 (N_13137,N_11956,N_10763);
or U13138 (N_13138,N_11996,N_10899);
and U13139 (N_13139,N_10888,N_11193);
and U13140 (N_13140,N_11740,N_10772);
nor U13141 (N_13141,N_10874,N_11885);
or U13142 (N_13142,N_11912,N_11404);
and U13143 (N_13143,N_11713,N_11101);
nand U13144 (N_13144,N_10749,N_11931);
xnor U13145 (N_13145,N_11469,N_10992);
or U13146 (N_13146,N_11022,N_11072);
nor U13147 (N_13147,N_11785,N_10598);
xnor U13148 (N_13148,N_10567,N_11569);
nand U13149 (N_13149,N_11456,N_11100);
nor U13150 (N_13150,N_11081,N_10807);
nor U13151 (N_13151,N_10668,N_11343);
and U13152 (N_13152,N_11284,N_11970);
and U13153 (N_13153,N_11514,N_10647);
xnor U13154 (N_13154,N_11964,N_11253);
or U13155 (N_13155,N_11061,N_10772);
xor U13156 (N_13156,N_10590,N_11129);
or U13157 (N_13157,N_11685,N_11181);
nand U13158 (N_13158,N_11456,N_11076);
xor U13159 (N_13159,N_11144,N_11930);
xor U13160 (N_13160,N_10529,N_11591);
and U13161 (N_13161,N_10600,N_10791);
or U13162 (N_13162,N_10779,N_10578);
or U13163 (N_13163,N_11353,N_10644);
and U13164 (N_13164,N_11147,N_11154);
or U13165 (N_13165,N_11814,N_11163);
xor U13166 (N_13166,N_10805,N_11952);
nor U13167 (N_13167,N_11651,N_11949);
nand U13168 (N_13168,N_10676,N_11786);
nor U13169 (N_13169,N_11808,N_10546);
or U13170 (N_13170,N_10905,N_11534);
nor U13171 (N_13171,N_11584,N_11831);
xor U13172 (N_13172,N_10521,N_11506);
nand U13173 (N_13173,N_11742,N_10893);
and U13174 (N_13174,N_10705,N_11545);
and U13175 (N_13175,N_11837,N_11462);
nand U13176 (N_13176,N_10832,N_11664);
or U13177 (N_13177,N_11473,N_11491);
xor U13178 (N_13178,N_11532,N_11413);
and U13179 (N_13179,N_11850,N_11426);
or U13180 (N_13180,N_10889,N_10931);
nand U13181 (N_13181,N_11212,N_10547);
nor U13182 (N_13182,N_11420,N_11073);
and U13183 (N_13183,N_10790,N_11400);
xor U13184 (N_13184,N_11705,N_11371);
and U13185 (N_13185,N_10923,N_10617);
and U13186 (N_13186,N_11601,N_11714);
and U13187 (N_13187,N_11290,N_11386);
or U13188 (N_13188,N_10938,N_11223);
and U13189 (N_13189,N_10576,N_10584);
and U13190 (N_13190,N_11043,N_10567);
and U13191 (N_13191,N_11507,N_11162);
and U13192 (N_13192,N_11651,N_11451);
nand U13193 (N_13193,N_10527,N_11568);
nand U13194 (N_13194,N_11053,N_11956);
or U13195 (N_13195,N_11905,N_11825);
and U13196 (N_13196,N_11826,N_11314);
or U13197 (N_13197,N_10736,N_11805);
nand U13198 (N_13198,N_11575,N_11227);
nor U13199 (N_13199,N_10978,N_11419);
nand U13200 (N_13200,N_10717,N_11646);
xnor U13201 (N_13201,N_11809,N_11099);
and U13202 (N_13202,N_11193,N_11697);
nand U13203 (N_13203,N_11561,N_11866);
or U13204 (N_13204,N_10624,N_10731);
or U13205 (N_13205,N_11885,N_11771);
or U13206 (N_13206,N_10849,N_10522);
nand U13207 (N_13207,N_11487,N_11958);
nand U13208 (N_13208,N_11937,N_11919);
nor U13209 (N_13209,N_11131,N_11278);
and U13210 (N_13210,N_11256,N_10584);
nand U13211 (N_13211,N_11418,N_10761);
and U13212 (N_13212,N_11762,N_10600);
nor U13213 (N_13213,N_11259,N_11514);
and U13214 (N_13214,N_10787,N_11653);
nor U13215 (N_13215,N_11851,N_11737);
or U13216 (N_13216,N_11583,N_10812);
nor U13217 (N_13217,N_11806,N_11310);
or U13218 (N_13218,N_11123,N_11350);
or U13219 (N_13219,N_11024,N_11280);
and U13220 (N_13220,N_10693,N_11215);
nand U13221 (N_13221,N_11983,N_11183);
xnor U13222 (N_13222,N_10648,N_10890);
or U13223 (N_13223,N_11092,N_11716);
or U13224 (N_13224,N_10925,N_10889);
xnor U13225 (N_13225,N_11722,N_10529);
nand U13226 (N_13226,N_11633,N_11454);
or U13227 (N_13227,N_10671,N_10753);
nand U13228 (N_13228,N_11573,N_11316);
nand U13229 (N_13229,N_11248,N_11229);
xnor U13230 (N_13230,N_11634,N_11983);
nor U13231 (N_13231,N_11264,N_11394);
xnor U13232 (N_13232,N_10849,N_11464);
nand U13233 (N_13233,N_11630,N_11830);
xor U13234 (N_13234,N_11041,N_11148);
xor U13235 (N_13235,N_11372,N_11494);
and U13236 (N_13236,N_11673,N_11250);
xnor U13237 (N_13237,N_11219,N_10517);
or U13238 (N_13238,N_11993,N_11465);
xor U13239 (N_13239,N_10827,N_11544);
and U13240 (N_13240,N_11881,N_11302);
or U13241 (N_13241,N_10608,N_10801);
and U13242 (N_13242,N_10504,N_11731);
nand U13243 (N_13243,N_11360,N_11803);
or U13244 (N_13244,N_10759,N_11512);
xnor U13245 (N_13245,N_11005,N_10531);
and U13246 (N_13246,N_11564,N_10737);
nand U13247 (N_13247,N_11558,N_11465);
nand U13248 (N_13248,N_10997,N_11167);
and U13249 (N_13249,N_11097,N_10526);
or U13250 (N_13250,N_10685,N_11385);
nor U13251 (N_13251,N_11532,N_10991);
xor U13252 (N_13252,N_11195,N_11777);
xor U13253 (N_13253,N_11081,N_11080);
or U13254 (N_13254,N_11334,N_11107);
or U13255 (N_13255,N_11919,N_10576);
and U13256 (N_13256,N_10900,N_11162);
xor U13257 (N_13257,N_10886,N_11825);
and U13258 (N_13258,N_11251,N_10561);
xor U13259 (N_13259,N_11412,N_11815);
xnor U13260 (N_13260,N_10821,N_11142);
nand U13261 (N_13261,N_11397,N_11702);
nand U13262 (N_13262,N_10528,N_11499);
nor U13263 (N_13263,N_11772,N_11700);
or U13264 (N_13264,N_10600,N_10665);
nand U13265 (N_13265,N_11604,N_11286);
or U13266 (N_13266,N_11402,N_11517);
nor U13267 (N_13267,N_11806,N_10776);
nand U13268 (N_13268,N_10592,N_10544);
xor U13269 (N_13269,N_11826,N_10513);
nor U13270 (N_13270,N_11686,N_11415);
and U13271 (N_13271,N_11919,N_10869);
or U13272 (N_13272,N_10740,N_11092);
nand U13273 (N_13273,N_10728,N_11625);
or U13274 (N_13274,N_11778,N_11096);
and U13275 (N_13275,N_11886,N_11016);
or U13276 (N_13276,N_11784,N_10859);
and U13277 (N_13277,N_10633,N_11380);
or U13278 (N_13278,N_11264,N_11541);
or U13279 (N_13279,N_11209,N_11883);
and U13280 (N_13280,N_11991,N_10908);
nor U13281 (N_13281,N_11907,N_11179);
or U13282 (N_13282,N_10952,N_11476);
nor U13283 (N_13283,N_11299,N_11467);
nand U13284 (N_13284,N_11356,N_10862);
or U13285 (N_13285,N_11839,N_10519);
xor U13286 (N_13286,N_10804,N_10559);
nand U13287 (N_13287,N_10658,N_11590);
and U13288 (N_13288,N_10952,N_11410);
or U13289 (N_13289,N_11380,N_10883);
or U13290 (N_13290,N_11962,N_10680);
or U13291 (N_13291,N_10766,N_10757);
or U13292 (N_13292,N_11984,N_10785);
nor U13293 (N_13293,N_11111,N_11953);
and U13294 (N_13294,N_10860,N_11734);
nor U13295 (N_13295,N_10862,N_11545);
xor U13296 (N_13296,N_11184,N_10514);
nor U13297 (N_13297,N_11263,N_11342);
nand U13298 (N_13298,N_10577,N_11496);
xor U13299 (N_13299,N_11859,N_11492);
xnor U13300 (N_13300,N_11454,N_11038);
and U13301 (N_13301,N_11373,N_10789);
or U13302 (N_13302,N_10858,N_11208);
and U13303 (N_13303,N_11798,N_10793);
xnor U13304 (N_13304,N_11774,N_11038);
or U13305 (N_13305,N_10740,N_10506);
nand U13306 (N_13306,N_10644,N_11988);
nor U13307 (N_13307,N_11065,N_11174);
and U13308 (N_13308,N_10742,N_11008);
and U13309 (N_13309,N_10733,N_10607);
nor U13310 (N_13310,N_10866,N_11217);
nand U13311 (N_13311,N_10587,N_10979);
nor U13312 (N_13312,N_10530,N_11710);
and U13313 (N_13313,N_11600,N_11962);
and U13314 (N_13314,N_11228,N_10621);
nor U13315 (N_13315,N_11710,N_11201);
xor U13316 (N_13316,N_10705,N_11056);
nor U13317 (N_13317,N_10835,N_10852);
xor U13318 (N_13318,N_11831,N_11109);
nand U13319 (N_13319,N_10834,N_11003);
nor U13320 (N_13320,N_11296,N_11430);
nor U13321 (N_13321,N_11586,N_11286);
xor U13322 (N_13322,N_11300,N_10510);
xor U13323 (N_13323,N_10729,N_11238);
xnor U13324 (N_13324,N_11937,N_11731);
and U13325 (N_13325,N_10715,N_11868);
xor U13326 (N_13326,N_11393,N_11718);
xnor U13327 (N_13327,N_11878,N_11587);
nor U13328 (N_13328,N_10595,N_11459);
and U13329 (N_13329,N_10640,N_10722);
xor U13330 (N_13330,N_11286,N_11162);
or U13331 (N_13331,N_11773,N_11526);
xnor U13332 (N_13332,N_10893,N_10932);
nor U13333 (N_13333,N_10828,N_11104);
or U13334 (N_13334,N_10997,N_11458);
nand U13335 (N_13335,N_11098,N_11533);
nor U13336 (N_13336,N_11262,N_10647);
nand U13337 (N_13337,N_10654,N_11526);
or U13338 (N_13338,N_11025,N_11394);
or U13339 (N_13339,N_11217,N_11727);
nor U13340 (N_13340,N_11680,N_11872);
nor U13341 (N_13341,N_11383,N_11586);
nand U13342 (N_13342,N_11109,N_11531);
and U13343 (N_13343,N_10846,N_10851);
nor U13344 (N_13344,N_10819,N_11812);
nor U13345 (N_13345,N_10705,N_11898);
and U13346 (N_13346,N_11491,N_11777);
or U13347 (N_13347,N_11101,N_10535);
nor U13348 (N_13348,N_11010,N_10515);
and U13349 (N_13349,N_11896,N_11439);
xor U13350 (N_13350,N_11426,N_10887);
nand U13351 (N_13351,N_11608,N_11616);
and U13352 (N_13352,N_11359,N_11724);
and U13353 (N_13353,N_11348,N_11722);
or U13354 (N_13354,N_10835,N_11114);
and U13355 (N_13355,N_11277,N_11390);
nand U13356 (N_13356,N_10523,N_10816);
or U13357 (N_13357,N_11680,N_10662);
nor U13358 (N_13358,N_10766,N_10562);
and U13359 (N_13359,N_10837,N_10981);
and U13360 (N_13360,N_11849,N_10825);
or U13361 (N_13361,N_10908,N_11760);
or U13362 (N_13362,N_11521,N_11219);
nor U13363 (N_13363,N_11762,N_11310);
xnor U13364 (N_13364,N_11536,N_10925);
and U13365 (N_13365,N_10949,N_11931);
nor U13366 (N_13366,N_11298,N_11947);
xor U13367 (N_13367,N_11217,N_11084);
or U13368 (N_13368,N_11906,N_11494);
and U13369 (N_13369,N_11109,N_11773);
xnor U13370 (N_13370,N_11711,N_11609);
or U13371 (N_13371,N_10933,N_11854);
nor U13372 (N_13372,N_10575,N_11909);
or U13373 (N_13373,N_11128,N_11592);
nand U13374 (N_13374,N_11787,N_11126);
and U13375 (N_13375,N_11883,N_11405);
xor U13376 (N_13376,N_11096,N_11240);
nor U13377 (N_13377,N_11971,N_11464);
nand U13378 (N_13378,N_11338,N_11141);
xor U13379 (N_13379,N_10871,N_10526);
or U13380 (N_13380,N_11648,N_11972);
nand U13381 (N_13381,N_11191,N_10870);
nand U13382 (N_13382,N_10514,N_10936);
xor U13383 (N_13383,N_10556,N_11263);
xnor U13384 (N_13384,N_11951,N_10553);
and U13385 (N_13385,N_11701,N_11509);
nand U13386 (N_13386,N_11002,N_11265);
nor U13387 (N_13387,N_11784,N_10937);
or U13388 (N_13388,N_10992,N_10950);
nand U13389 (N_13389,N_10564,N_11465);
or U13390 (N_13390,N_10505,N_10589);
nor U13391 (N_13391,N_11797,N_10971);
xnor U13392 (N_13392,N_11165,N_11101);
nand U13393 (N_13393,N_11309,N_11811);
xnor U13394 (N_13394,N_11787,N_11906);
or U13395 (N_13395,N_11225,N_11186);
nor U13396 (N_13396,N_11757,N_11943);
or U13397 (N_13397,N_11887,N_11226);
and U13398 (N_13398,N_10867,N_10715);
nor U13399 (N_13399,N_11978,N_11857);
nor U13400 (N_13400,N_11915,N_11199);
xor U13401 (N_13401,N_11345,N_11805);
nor U13402 (N_13402,N_11532,N_10850);
xnor U13403 (N_13403,N_11990,N_11499);
or U13404 (N_13404,N_11388,N_11820);
nor U13405 (N_13405,N_11761,N_11823);
nor U13406 (N_13406,N_10889,N_11970);
nor U13407 (N_13407,N_11652,N_10709);
nand U13408 (N_13408,N_10538,N_10990);
or U13409 (N_13409,N_10621,N_11422);
xor U13410 (N_13410,N_11018,N_10639);
nand U13411 (N_13411,N_11823,N_11669);
and U13412 (N_13412,N_11619,N_11885);
nand U13413 (N_13413,N_11244,N_11038);
nor U13414 (N_13414,N_11693,N_10570);
nor U13415 (N_13415,N_11667,N_11513);
nor U13416 (N_13416,N_11050,N_11194);
xnor U13417 (N_13417,N_11017,N_10626);
nor U13418 (N_13418,N_10831,N_10632);
and U13419 (N_13419,N_10866,N_10618);
xor U13420 (N_13420,N_11786,N_11323);
nand U13421 (N_13421,N_11156,N_10528);
xor U13422 (N_13422,N_10549,N_11879);
xor U13423 (N_13423,N_11193,N_10897);
and U13424 (N_13424,N_11011,N_10892);
nor U13425 (N_13425,N_11443,N_11625);
nand U13426 (N_13426,N_11971,N_11474);
nand U13427 (N_13427,N_10721,N_10513);
xnor U13428 (N_13428,N_11746,N_11884);
nor U13429 (N_13429,N_10544,N_11457);
nand U13430 (N_13430,N_11319,N_11206);
and U13431 (N_13431,N_11228,N_11514);
xnor U13432 (N_13432,N_10805,N_10706);
or U13433 (N_13433,N_10668,N_11265);
nand U13434 (N_13434,N_11829,N_10588);
nor U13435 (N_13435,N_10544,N_11186);
nand U13436 (N_13436,N_11587,N_11102);
xor U13437 (N_13437,N_11794,N_11378);
or U13438 (N_13438,N_10733,N_11146);
and U13439 (N_13439,N_11623,N_10547);
or U13440 (N_13440,N_11876,N_10872);
or U13441 (N_13441,N_11502,N_11128);
and U13442 (N_13442,N_10551,N_10660);
and U13443 (N_13443,N_10715,N_11246);
or U13444 (N_13444,N_10640,N_10763);
xnor U13445 (N_13445,N_11741,N_11306);
nand U13446 (N_13446,N_10917,N_10767);
or U13447 (N_13447,N_11904,N_11500);
or U13448 (N_13448,N_10752,N_10936);
or U13449 (N_13449,N_10769,N_10525);
and U13450 (N_13450,N_11359,N_10921);
or U13451 (N_13451,N_11532,N_10613);
or U13452 (N_13452,N_11295,N_11263);
and U13453 (N_13453,N_10560,N_11809);
xnor U13454 (N_13454,N_11261,N_11752);
nor U13455 (N_13455,N_10849,N_11217);
xor U13456 (N_13456,N_10904,N_11063);
and U13457 (N_13457,N_11509,N_10778);
xnor U13458 (N_13458,N_11754,N_11099);
and U13459 (N_13459,N_11849,N_11545);
xnor U13460 (N_13460,N_10954,N_11901);
nor U13461 (N_13461,N_10588,N_11760);
and U13462 (N_13462,N_10907,N_10682);
or U13463 (N_13463,N_10786,N_11991);
xor U13464 (N_13464,N_11226,N_11868);
and U13465 (N_13465,N_10872,N_10790);
nor U13466 (N_13466,N_11487,N_11205);
and U13467 (N_13467,N_11045,N_11462);
or U13468 (N_13468,N_11851,N_11235);
and U13469 (N_13469,N_11491,N_11655);
nor U13470 (N_13470,N_10704,N_11765);
nand U13471 (N_13471,N_11622,N_11957);
xor U13472 (N_13472,N_11709,N_11150);
and U13473 (N_13473,N_10851,N_11194);
nand U13474 (N_13474,N_11428,N_11210);
xor U13475 (N_13475,N_11129,N_10963);
nor U13476 (N_13476,N_10723,N_11510);
nand U13477 (N_13477,N_11221,N_11974);
nand U13478 (N_13478,N_11099,N_10586);
and U13479 (N_13479,N_11125,N_10599);
or U13480 (N_13480,N_11800,N_11076);
and U13481 (N_13481,N_11132,N_11552);
nor U13482 (N_13482,N_11150,N_11474);
or U13483 (N_13483,N_11401,N_11353);
or U13484 (N_13484,N_10723,N_10892);
nor U13485 (N_13485,N_11498,N_10674);
and U13486 (N_13486,N_11042,N_11154);
nand U13487 (N_13487,N_11912,N_11477);
xnor U13488 (N_13488,N_11237,N_11424);
nor U13489 (N_13489,N_11695,N_11326);
xor U13490 (N_13490,N_10825,N_10901);
nand U13491 (N_13491,N_11254,N_10675);
and U13492 (N_13492,N_10580,N_10837);
and U13493 (N_13493,N_10602,N_11847);
xnor U13494 (N_13494,N_11819,N_11116);
nor U13495 (N_13495,N_10765,N_11322);
nand U13496 (N_13496,N_11462,N_11507);
or U13497 (N_13497,N_11408,N_11190);
or U13498 (N_13498,N_11794,N_10866);
nand U13499 (N_13499,N_10946,N_11724);
and U13500 (N_13500,N_12020,N_12027);
and U13501 (N_13501,N_12989,N_12024);
and U13502 (N_13502,N_13447,N_12844);
or U13503 (N_13503,N_12992,N_12053);
nand U13504 (N_13504,N_12002,N_12095);
nand U13505 (N_13505,N_12284,N_12650);
nor U13506 (N_13506,N_12398,N_12167);
nor U13507 (N_13507,N_12474,N_12191);
nand U13508 (N_13508,N_12213,N_12573);
xor U13509 (N_13509,N_12156,N_12585);
xnor U13510 (N_13510,N_12238,N_13190);
nor U13511 (N_13511,N_12139,N_12807);
nand U13512 (N_13512,N_13259,N_12455);
and U13513 (N_13513,N_12374,N_13392);
or U13514 (N_13514,N_13154,N_12879);
xor U13515 (N_13515,N_12184,N_13384);
or U13516 (N_13516,N_13039,N_12819);
or U13517 (N_13517,N_13306,N_12884);
or U13518 (N_13518,N_12193,N_12952);
nor U13519 (N_13519,N_12604,N_12809);
nand U13520 (N_13520,N_12037,N_12522);
and U13521 (N_13521,N_12559,N_13243);
nand U13522 (N_13522,N_12436,N_12306);
or U13523 (N_13523,N_12896,N_12640);
xnor U13524 (N_13524,N_12043,N_12251);
nand U13525 (N_13525,N_13491,N_12851);
nor U13526 (N_13526,N_13409,N_13041);
and U13527 (N_13527,N_12719,N_12003);
nand U13528 (N_13528,N_12776,N_13371);
nor U13529 (N_13529,N_13000,N_12326);
or U13530 (N_13530,N_12483,N_12810);
nand U13531 (N_13531,N_12300,N_12386);
or U13532 (N_13532,N_12318,N_12293);
xor U13533 (N_13533,N_12970,N_12246);
xor U13534 (N_13534,N_12791,N_13167);
nor U13535 (N_13535,N_12537,N_12951);
nand U13536 (N_13536,N_13382,N_13493);
nor U13537 (N_13537,N_13426,N_13304);
nor U13538 (N_13538,N_12907,N_12968);
nand U13539 (N_13539,N_13239,N_12305);
xnor U13540 (N_13540,N_12571,N_12128);
and U13541 (N_13541,N_12085,N_12860);
nor U13542 (N_13542,N_12721,N_12836);
nor U13543 (N_13543,N_12515,N_12667);
nor U13544 (N_13544,N_12308,N_12096);
and U13545 (N_13545,N_12545,N_13488);
or U13546 (N_13546,N_13494,N_12120);
xnor U13547 (N_13547,N_13347,N_13081);
or U13548 (N_13548,N_12174,N_12507);
nand U13549 (N_13549,N_13354,N_12105);
or U13550 (N_13550,N_13127,N_12966);
xor U13551 (N_13551,N_13102,N_13018);
nor U13552 (N_13552,N_13029,N_13476);
nand U13553 (N_13553,N_12116,N_13153);
nand U13554 (N_13554,N_12596,N_13189);
or U13555 (N_13555,N_12449,N_13214);
nor U13556 (N_13556,N_13182,N_12677);
and U13557 (N_13557,N_13463,N_12025);
nor U13558 (N_13558,N_12710,N_12083);
xnor U13559 (N_13559,N_12565,N_12220);
xor U13560 (N_13560,N_13397,N_12421);
and U13561 (N_13561,N_12379,N_13183);
xnor U13562 (N_13562,N_12853,N_13475);
or U13563 (N_13563,N_12689,N_12115);
xnor U13564 (N_13564,N_13341,N_12550);
nand U13565 (N_13565,N_12804,N_12378);
nand U13566 (N_13566,N_12649,N_12781);
nor U13567 (N_13567,N_12646,N_13107);
nand U13568 (N_13568,N_12605,N_13236);
or U13569 (N_13569,N_13356,N_12200);
nor U13570 (N_13570,N_13066,N_13418);
nor U13571 (N_13571,N_13301,N_13380);
nor U13572 (N_13572,N_12471,N_13440);
nor U13573 (N_13573,N_12936,N_12501);
nor U13574 (N_13574,N_12314,N_12068);
nand U13575 (N_13575,N_12316,N_12842);
nor U13576 (N_13576,N_13288,N_12877);
nand U13577 (N_13577,N_12761,N_12848);
nand U13578 (N_13578,N_12948,N_12103);
xor U13579 (N_13579,N_13485,N_13372);
nor U13580 (N_13580,N_12814,N_12023);
xnor U13581 (N_13581,N_12445,N_12777);
or U13582 (N_13582,N_12558,N_13135);
nor U13583 (N_13583,N_13121,N_13109);
nor U13584 (N_13584,N_12711,N_12614);
and U13585 (N_13585,N_13100,N_12375);
nor U13586 (N_13586,N_13191,N_13360);
nand U13587 (N_13587,N_12199,N_12000);
and U13588 (N_13588,N_12756,N_12938);
xor U13589 (N_13589,N_12214,N_12429);
xnor U13590 (N_13590,N_12805,N_13162);
or U13591 (N_13591,N_13312,N_12882);
nand U13592 (N_13592,N_13231,N_13052);
xor U13593 (N_13593,N_12399,N_12979);
and U13594 (N_13594,N_13076,N_12747);
or U13595 (N_13595,N_12051,N_12491);
or U13596 (N_13596,N_13155,N_12690);
and U13597 (N_13597,N_13496,N_12612);
nand U13598 (N_13598,N_13298,N_12930);
nor U13599 (N_13599,N_12385,N_12289);
nand U13600 (N_13600,N_13205,N_12917);
nand U13601 (N_13601,N_13224,N_12475);
nor U13602 (N_13602,N_12658,N_12058);
and U13603 (N_13603,N_13391,N_13203);
and U13604 (N_13604,N_13229,N_12755);
and U13605 (N_13605,N_12588,N_12465);
xnor U13606 (N_13606,N_12204,N_12880);
and U13607 (N_13607,N_13201,N_13471);
or U13608 (N_13608,N_12619,N_13207);
nand U13609 (N_13609,N_13209,N_12766);
or U13610 (N_13610,N_12933,N_12716);
and U13611 (N_13611,N_12392,N_13446);
or U13612 (N_13612,N_12134,N_12090);
or U13613 (N_13613,N_12878,N_12542);
and U13614 (N_13614,N_13035,N_13221);
and U13615 (N_13615,N_12922,N_12180);
nor U13616 (N_13616,N_13065,N_12787);
and U13617 (N_13617,N_13443,N_12151);
and U13618 (N_13618,N_12744,N_12950);
nor U13619 (N_13619,N_13200,N_12135);
xor U13620 (N_13620,N_12118,N_12645);
and U13621 (N_13621,N_13194,N_12126);
nor U13622 (N_13622,N_12488,N_12476);
and U13623 (N_13623,N_13262,N_12397);
or U13624 (N_13624,N_13444,N_13110);
nand U13625 (N_13625,N_12955,N_13142);
nor U13626 (N_13626,N_12531,N_12357);
and U13627 (N_13627,N_13406,N_13385);
and U13628 (N_13628,N_12282,N_12256);
and U13629 (N_13629,N_12201,N_13405);
or U13630 (N_13630,N_12643,N_13428);
nand U13631 (N_13631,N_12462,N_13365);
and U13632 (N_13632,N_13055,N_12901);
nand U13633 (N_13633,N_12629,N_12358);
xnor U13634 (N_13634,N_12954,N_13098);
nand U13635 (N_13635,N_12353,N_12048);
and U13636 (N_13636,N_12500,N_12235);
and U13637 (N_13637,N_12827,N_12290);
or U13638 (N_13638,N_12811,N_12511);
nand U13639 (N_13639,N_12541,N_12032);
nand U13640 (N_13640,N_12258,N_12112);
and U13641 (N_13641,N_12188,N_13343);
and U13642 (N_13642,N_13139,N_12798);
or U13643 (N_13643,N_13060,N_12826);
or U13644 (N_13644,N_12816,N_12957);
or U13645 (N_13645,N_12803,N_12919);
xnor U13646 (N_13646,N_12533,N_13241);
nand U13647 (N_13647,N_12363,N_12109);
xnor U13648 (N_13648,N_12539,N_12015);
xor U13649 (N_13649,N_12228,N_13078);
and U13650 (N_13650,N_12005,N_12270);
nand U13651 (N_13651,N_12010,N_13174);
xor U13652 (N_13652,N_12050,N_12143);
nor U13653 (N_13653,N_12381,N_12028);
nor U13654 (N_13654,N_12762,N_12327);
or U13655 (N_13655,N_12124,N_12872);
xnor U13656 (N_13656,N_13086,N_12260);
nand U13657 (N_13657,N_12724,N_12442);
xnor U13658 (N_13658,N_13411,N_12976);
nor U13659 (N_13659,N_12609,N_12944);
nand U13660 (N_13660,N_12606,N_12031);
nand U13661 (N_13661,N_12924,N_12457);
nor U13662 (N_13662,N_13091,N_12998);
nor U13663 (N_13663,N_12740,N_12712);
and U13664 (N_13664,N_12017,N_12163);
or U13665 (N_13665,N_13416,N_12512);
and U13666 (N_13666,N_13219,N_12245);
or U13667 (N_13667,N_12767,N_12893);
nor U13668 (N_13668,N_13001,N_12407);
and U13669 (N_13669,N_13332,N_12106);
nor U13670 (N_13670,N_13187,N_12557);
nor U13671 (N_13671,N_12775,N_12732);
nor U13672 (N_13672,N_12613,N_12611);
nand U13673 (N_13673,N_12789,N_12838);
or U13674 (N_13674,N_12699,N_13019);
nand U13675 (N_13675,N_12945,N_12946);
nor U13676 (N_13676,N_12348,N_13075);
and U13677 (N_13677,N_13467,N_12082);
or U13678 (N_13678,N_12279,N_13253);
and U13679 (N_13679,N_13160,N_13492);
nor U13680 (N_13680,N_13090,N_12865);
nor U13681 (N_13681,N_12013,N_13292);
nor U13682 (N_13682,N_12864,N_12543);
nor U13683 (N_13683,N_12499,N_12519);
or U13684 (N_13684,N_12546,N_12837);
nand U13685 (N_13685,N_13350,N_13282);
or U13686 (N_13686,N_13171,N_13248);
nand U13687 (N_13687,N_12001,N_13223);
and U13688 (N_13688,N_13464,N_12319);
or U13689 (N_13689,N_13257,N_12181);
xnor U13690 (N_13690,N_12423,N_13179);
xnor U13691 (N_13691,N_12812,N_12736);
or U13692 (N_13692,N_12535,N_12654);
and U13693 (N_13693,N_12818,N_12996);
xor U13694 (N_13694,N_12127,N_12739);
and U13695 (N_13695,N_12347,N_12041);
or U13696 (N_13696,N_13424,N_12355);
nor U13697 (N_13697,N_13453,N_12185);
or U13698 (N_13698,N_12782,N_12485);
and U13699 (N_13699,N_12580,N_12212);
or U13700 (N_13700,N_13175,N_13323);
nand U13701 (N_13701,N_13053,N_13419);
and U13702 (N_13702,N_12505,N_12593);
and U13703 (N_13703,N_12177,N_13389);
and U13704 (N_13704,N_12594,N_13294);
and U13705 (N_13705,N_12720,N_12749);
and U13706 (N_13706,N_12012,N_12509);
or U13707 (N_13707,N_12569,N_13003);
nand U13708 (N_13708,N_12099,N_13237);
xnor U13709 (N_13709,N_12591,N_12150);
or U13710 (N_13710,N_12662,N_12661);
nand U13711 (N_13711,N_12928,N_12479);
or U13712 (N_13712,N_12339,N_12990);
nor U13713 (N_13713,N_12133,N_12898);
and U13714 (N_13714,N_13181,N_12881);
xor U13715 (N_13715,N_12961,N_13011);
nand U13716 (N_13716,N_12030,N_12734);
xor U13717 (N_13717,N_13336,N_12248);
xor U13718 (N_13718,N_12639,N_12373);
nand U13719 (N_13719,N_13266,N_12470);
xor U13720 (N_13720,N_12978,N_12259);
or U13721 (N_13721,N_12987,N_13400);
xnor U13722 (N_13722,N_12831,N_12758);
nand U13723 (N_13723,N_12908,N_12183);
xor U13724 (N_13724,N_12039,N_12751);
nor U13725 (N_13725,N_12469,N_12680);
nor U13726 (N_13726,N_13126,N_13238);
and U13727 (N_13727,N_12493,N_12273);
nor U13728 (N_13728,N_12584,N_12100);
and U13729 (N_13729,N_13412,N_12207);
and U13730 (N_13730,N_12480,N_13252);
nand U13731 (N_13731,N_12145,N_13348);
nand U13732 (N_13732,N_12779,N_12021);
and U13733 (N_13733,N_12210,N_12854);
nor U13734 (N_13734,N_12332,N_12272);
nand U13735 (N_13735,N_12304,N_12376);
nand U13736 (N_13736,N_12309,N_13450);
or U13737 (N_13737,N_12351,N_12560);
or U13738 (N_13738,N_13159,N_13274);
or U13739 (N_13739,N_13284,N_12026);
and U13740 (N_13740,N_12988,N_12551);
or U13741 (N_13741,N_13345,N_12947);
nand U13742 (N_13742,N_12354,N_12504);
or U13743 (N_13743,N_12194,N_12123);
or U13744 (N_13744,N_13123,N_13062);
nor U13745 (N_13745,N_13349,N_13012);
nor U13746 (N_13746,N_12523,N_12390);
and U13747 (N_13747,N_12155,N_13379);
and U13748 (N_13748,N_12323,N_13273);
xor U13749 (N_13749,N_12858,N_12905);
and U13750 (N_13750,N_12298,N_12705);
or U13751 (N_13751,N_12994,N_12287);
and U13752 (N_13752,N_12179,N_12602);
nand U13753 (N_13753,N_12703,N_12935);
or U13754 (N_13754,N_13161,N_12502);
nor U13755 (N_13755,N_12647,N_12603);
nor U13756 (N_13756,N_12760,N_13178);
and U13757 (N_13757,N_13269,N_12876);
nand U13758 (N_13758,N_13013,N_13408);
xor U13759 (N_13759,N_12621,N_12634);
xnor U13760 (N_13760,N_12315,N_12129);
nor U13761 (N_13761,N_12294,N_13344);
and U13762 (N_13762,N_13324,N_12839);
xor U13763 (N_13763,N_12198,N_13459);
nand U13764 (N_13764,N_12008,N_12490);
nor U13765 (N_13765,N_12477,N_12682);
or U13766 (N_13766,N_13202,N_12302);
nand U13767 (N_13767,N_12088,N_13197);
nor U13768 (N_13768,N_13032,N_12079);
nand U13769 (N_13769,N_13263,N_12635);
and U13770 (N_13770,N_12886,N_13329);
nor U13771 (N_13771,N_13092,N_13114);
and U13772 (N_13772,N_12579,N_12520);
nor U13773 (N_13773,N_12738,N_12576);
and U13774 (N_13774,N_13369,N_12274);
or U13775 (N_13775,N_12446,N_13157);
xor U13776 (N_13776,N_12057,N_13327);
and U13777 (N_13777,N_12723,N_12478);
nor U13778 (N_13778,N_13402,N_12265);
nor U13779 (N_13779,N_13116,N_12496);
nand U13780 (N_13780,N_12940,N_12536);
and U13781 (N_13781,N_12587,N_12731);
nand U13782 (N_13782,N_13456,N_13285);
nand U13783 (N_13783,N_12295,N_12859);
or U13784 (N_13784,N_13240,N_12081);
or U13785 (N_13785,N_13046,N_13265);
nor U13786 (N_13786,N_12395,N_12035);
nand U13787 (N_13787,N_13325,N_13130);
nor U13788 (N_13788,N_12513,N_12503);
and U13789 (N_13789,N_13145,N_12117);
nand U13790 (N_13790,N_12891,N_12540);
nand U13791 (N_13791,N_12400,N_13427);
or U13792 (N_13792,N_13319,N_12042);
nand U13793 (N_13793,N_12165,N_12773);
or U13794 (N_13794,N_12223,N_12387);
nor U13795 (N_13795,N_12065,N_13279);
nand U13796 (N_13796,N_12598,N_12828);
nor U13797 (N_13797,N_12056,N_12414);
or U13798 (N_13798,N_13027,N_12317);
nor U13799 (N_13799,N_12674,N_12620);
nand U13800 (N_13800,N_12942,N_13346);
and U13801 (N_13801,N_12219,N_12029);
or U13802 (N_13802,N_12855,N_13249);
xnor U13803 (N_13803,N_12225,N_12344);
or U13804 (N_13804,N_13481,N_12195);
and U13805 (N_13805,N_13088,N_12949);
and U13806 (N_13806,N_13472,N_12014);
nor U13807 (N_13807,N_12974,N_12067);
or U13808 (N_13808,N_12391,N_12313);
nand U13809 (N_13809,N_12368,N_12422);
nor U13810 (N_13810,N_12244,N_12281);
nand U13811 (N_13811,N_13124,N_13061);
or U13812 (N_13812,N_12328,N_12847);
xnor U13813 (N_13813,N_12548,N_13024);
xor U13814 (N_13814,N_13199,N_13125);
nor U13815 (N_13815,N_12016,N_12055);
or U13816 (N_13816,N_13217,N_12651);
nor U13817 (N_13817,N_12247,N_12856);
nand U13818 (N_13818,N_12506,N_12845);
or U13819 (N_13819,N_13339,N_12047);
nand U13820 (N_13820,N_12999,N_12482);
nor U13821 (N_13821,N_13195,N_12239);
and U13822 (N_13822,N_13048,N_12900);
xnor U13823 (N_13823,N_12401,N_12104);
xor U13824 (N_13824,N_12370,N_13216);
xor U13825 (N_13825,N_13056,N_13451);
nand U13826 (N_13826,N_12664,N_13364);
and U13827 (N_13827,N_12561,N_12359);
nor U13828 (N_13828,N_13387,N_12234);
or U13829 (N_13829,N_12329,N_13177);
and U13830 (N_13830,N_13401,N_13367);
nor U13831 (N_13831,N_12735,N_12192);
or U13832 (N_13832,N_13393,N_12937);
nor U13833 (N_13833,N_12346,N_13302);
nor U13834 (N_13834,N_13164,N_12280);
nand U13835 (N_13835,N_12226,N_12340);
or U13836 (N_13836,N_12380,N_12402);
nand U13837 (N_13837,N_12769,N_12726);
nand U13838 (N_13838,N_13328,N_13296);
and U13839 (N_13839,N_13070,N_13251);
or U13840 (N_13840,N_12419,N_12054);
and U13841 (N_13841,N_12953,N_12679);
xor U13842 (N_13842,N_13132,N_12396);
or U13843 (N_13843,N_13004,N_12683);
and U13844 (N_13844,N_12456,N_12852);
nand U13845 (N_13845,N_13270,N_13377);
and U13846 (N_13846,N_12526,N_12321);
nand U13847 (N_13847,N_13310,N_13452);
xor U13848 (N_13848,N_12750,N_12943);
and U13849 (N_13849,N_12211,N_12458);
or U13850 (N_13850,N_12562,N_12849);
xor U13851 (N_13851,N_12464,N_12742);
nand U13852 (N_13852,N_12973,N_12266);
and U13853 (N_13853,N_12965,N_12011);
and U13854 (N_13854,N_12737,N_12795);
or U13855 (N_13855,N_12241,N_12595);
nand U13856 (N_13856,N_13271,N_13366);
xnor U13857 (N_13857,N_12700,N_12916);
or U13858 (N_13858,N_12254,N_12417);
and U13859 (N_13859,N_12444,N_12119);
and U13860 (N_13860,N_12846,N_12072);
and U13861 (N_13861,N_13006,N_12589);
xnor U13862 (N_13862,N_12632,N_12770);
nand U13863 (N_13863,N_12369,N_12525);
xor U13864 (N_13864,N_12434,N_12448);
and U13865 (N_13865,N_12277,N_12796);
and U13866 (N_13866,N_12532,N_13099);
and U13867 (N_13867,N_12084,N_12252);
nand U13868 (N_13868,N_13313,N_12186);
xnor U13869 (N_13869,N_13022,N_12829);
xor U13870 (N_13870,N_12275,N_12570);
xor U13871 (N_13871,N_12963,N_13449);
nand U13872 (N_13872,N_12463,N_12841);
and U13873 (N_13873,N_12285,N_12832);
nand U13874 (N_13874,N_13170,N_12197);
and U13875 (N_13875,N_12430,N_12006);
or U13876 (N_13876,N_12172,N_13415);
or U13877 (N_13877,N_12964,N_12790);
and U13878 (N_13878,N_12336,N_12702);
and U13879 (N_13879,N_12495,N_12659);
nor U13880 (N_13880,N_12615,N_13468);
and U13881 (N_13881,N_12388,N_13108);
or U13882 (N_13882,N_12921,N_13470);
xnor U13883 (N_13883,N_13105,N_12384);
and U13884 (N_13884,N_13407,N_12544);
nand U13885 (N_13885,N_12371,N_13342);
nand U13886 (N_13886,N_13436,N_13010);
or U13887 (N_13887,N_12034,N_12524);
and U13888 (N_13888,N_13146,N_12060);
nand U13889 (N_13889,N_12164,N_12022);
or U13890 (N_13890,N_13074,N_12330);
xor U13891 (N_13891,N_12741,N_12406);
and U13892 (N_13892,N_13396,N_12094);
and U13893 (N_13893,N_13163,N_12644);
and U13894 (N_13894,N_12276,N_13156);
or U13895 (N_13895,N_12553,N_12222);
nor U13896 (N_13896,N_12138,N_13335);
xnor U13897 (N_13897,N_13106,N_12073);
xor U13898 (N_13898,N_12110,N_12394);
nor U13899 (N_13899,N_13281,N_12076);
nand U13900 (N_13900,N_12607,N_13141);
nand U13901 (N_13901,N_13250,N_13381);
xor U13902 (N_13902,N_12078,N_12498);
or U13903 (N_13903,N_12492,N_13432);
or U13904 (N_13904,N_13455,N_13136);
or U13905 (N_13905,N_12345,N_12343);
nand U13906 (N_13906,N_12160,N_12910);
or U13907 (N_13907,N_13245,N_12296);
xor U13908 (N_13908,N_13311,N_12971);
nor U13909 (N_13909,N_13474,N_13120);
nor U13910 (N_13910,N_12563,N_13026);
or U13911 (N_13911,N_12366,N_12920);
or U13912 (N_13912,N_12624,N_13283);
nand U13913 (N_13913,N_13084,N_12869);
nand U13914 (N_13914,N_13005,N_13227);
xor U13915 (N_13915,N_13465,N_12918);
nand U13916 (N_13916,N_13002,N_12062);
xnor U13917 (N_13917,N_13338,N_13276);
nor U13918 (N_13918,N_12801,N_12383);
and U13919 (N_13919,N_13077,N_13320);
or U13920 (N_13920,N_13028,N_13417);
xnor U13921 (N_13921,N_13034,N_12362);
nor U13922 (N_13922,N_13272,N_13307);
xnor U13923 (N_13923,N_12783,N_13212);
and U13924 (N_13924,N_12410,N_12894);
nand U13925 (N_13925,N_12638,N_12903);
and U13926 (N_13926,N_12257,N_13308);
nand U13927 (N_13927,N_12286,N_12692);
and U13928 (N_13928,N_12975,N_12472);
nor U13929 (N_13929,N_13318,N_12871);
and U13930 (N_13930,N_12676,N_12148);
nor U13931 (N_13931,N_12046,N_12066);
and U13932 (N_13932,N_13040,N_12176);
nand U13933 (N_13933,N_12815,N_13420);
nand U13934 (N_13934,N_13193,N_13370);
nor U13935 (N_13935,N_12653,N_13043);
or U13936 (N_13936,N_12824,N_13051);
nor U13937 (N_13937,N_13425,N_12069);
and U13938 (N_13938,N_12799,N_13430);
nor U13939 (N_13939,N_13305,N_13134);
and U13940 (N_13940,N_12631,N_12958);
nor U13941 (N_13941,N_12583,N_12432);
and U13942 (N_13942,N_12098,N_12967);
nor U13943 (N_13943,N_13267,N_12518);
or U13944 (N_13944,N_12018,N_12147);
nor U13945 (N_13945,N_12821,N_12435);
xor U13946 (N_13946,N_12521,N_12554);
nand U13947 (N_13947,N_12625,N_12061);
nand U13948 (N_13948,N_12695,N_13246);
or U13949 (N_13949,N_13352,N_12412);
and U13950 (N_13950,N_12743,N_13152);
nor U13951 (N_13951,N_12311,N_12774);
or U13952 (N_13952,N_13023,N_12019);
nand U13953 (N_13953,N_12696,N_12941);
and U13954 (N_13954,N_12460,N_12980);
nand U13955 (N_13955,N_12320,N_12240);
xor U13956 (N_13956,N_12107,N_13413);
nand U13957 (N_13957,N_12627,N_13309);
nor U13958 (N_13958,N_12694,N_12202);
nand U13959 (N_13959,N_12508,N_12087);
xor U13960 (N_13960,N_12045,N_12516);
nor U13961 (N_13961,N_13495,N_12514);
nor U13962 (N_13962,N_13461,N_12004);
xor U13963 (N_13963,N_12264,N_12669);
and U13964 (N_13964,N_13016,N_13333);
and U13965 (N_13965,N_13254,N_12451);
xnor U13966 (N_13966,N_13278,N_12232);
or U13967 (N_13967,N_12806,N_12698);
nor U13968 (N_13968,N_12468,N_12729);
or U13969 (N_13969,N_12555,N_13128);
or U13970 (N_13970,N_13434,N_13235);
or U13971 (N_13971,N_13093,N_12497);
nand U13972 (N_13972,N_12249,N_12243);
nand U13973 (N_13973,N_12697,N_12209);
nand U13974 (N_13974,N_13486,N_13458);
nor U13975 (N_13975,N_13143,N_13192);
or U13976 (N_13976,N_12166,N_13487);
nand U13977 (N_13977,N_13258,N_13484);
nand U13978 (N_13978,N_13466,N_12820);
or U13979 (N_13979,N_12709,N_13168);
nand U13980 (N_13980,N_12171,N_13047);
nand U13981 (N_13981,N_12484,N_12863);
xor U13982 (N_13982,N_12857,N_12230);
xor U13983 (N_13983,N_13131,N_13399);
and U13984 (N_13984,N_13103,N_13129);
nand U13985 (N_13985,N_12342,N_13150);
and U13986 (N_13986,N_12159,N_12227);
nor U13987 (N_13987,N_12310,N_12586);
and U13988 (N_13988,N_13045,N_13118);
xnor U13989 (N_13989,N_12216,N_12049);
or U13990 (N_13990,N_13490,N_13151);
or U13991 (N_13991,N_12873,N_13133);
or U13992 (N_13992,N_12268,N_12673);
nor U13993 (N_13993,N_12808,N_13423);
nor U13994 (N_13994,N_12086,N_12149);
nand U13995 (N_13995,N_12617,N_13068);
nand U13996 (N_13996,N_12253,N_13477);
or U13997 (N_13997,N_12409,N_12101);
or U13998 (N_13998,N_13362,N_13457);
or U13999 (N_13999,N_12324,N_13206);
or U14000 (N_14000,N_12443,N_13149);
and U14001 (N_14001,N_12092,N_13033);
and U14002 (N_14002,N_12636,N_12913);
or U14003 (N_14003,N_13388,N_13218);
nand U14004 (N_14004,N_12530,N_12708);
and U14005 (N_14005,N_13422,N_12686);
xnor U14006 (N_14006,N_12608,N_12578);
or U14007 (N_14007,N_12349,N_13483);
and U14008 (N_14008,N_12759,N_12840);
or U14009 (N_14009,N_13303,N_12425);
or U14010 (N_14010,N_12360,N_13264);
nand U14011 (N_14011,N_13211,N_13386);
or U14012 (N_14012,N_12835,N_13025);
xnor U14013 (N_14013,N_12059,N_13111);
nor U14014 (N_14014,N_13176,N_12215);
xor U14015 (N_14015,N_13017,N_13196);
nor U14016 (N_14016,N_13255,N_12577);
nand U14017 (N_14017,N_12125,N_12897);
or U14018 (N_14018,N_12454,N_12784);
nor U14019 (N_14019,N_12452,N_12727);
and U14020 (N_14020,N_12527,N_12701);
or U14021 (N_14021,N_12169,N_13355);
and U14022 (N_14022,N_12338,N_12361);
or U14023 (N_14023,N_12113,N_13448);
or U14024 (N_14024,N_12299,N_12064);
nor U14025 (N_14025,N_12861,N_12161);
and U14026 (N_14026,N_12292,N_13460);
nor U14027 (N_14027,N_13085,N_13290);
xnor U14028 (N_14028,N_13094,N_13442);
xnor U14029 (N_14029,N_12926,N_13390);
xor U14030 (N_14030,N_13234,N_12036);
or U14031 (N_14031,N_12972,N_12111);
nor U14032 (N_14032,N_13233,N_12875);
and U14033 (N_14033,N_12684,N_12263);
or U14034 (N_14034,N_12529,N_12693);
nand U14035 (N_14035,N_12044,N_12372);
or U14036 (N_14036,N_13169,N_12335);
or U14037 (N_14037,N_12622,N_12486);
nor U14038 (N_14038,N_12038,N_12231);
xor U14039 (N_14039,N_13244,N_13398);
nand U14040 (N_14040,N_13071,N_13138);
and U14041 (N_14041,N_12467,N_12752);
or U14042 (N_14042,N_12556,N_12888);
nor U14043 (N_14043,N_12599,N_13059);
or U14044 (N_14044,N_12794,N_13403);
nand U14045 (N_14045,N_13277,N_13469);
nand U14046 (N_14046,N_12642,N_12887);
xnor U14047 (N_14047,N_13316,N_13137);
nor U14048 (N_14048,N_12331,N_12763);
nor U14049 (N_14049,N_12261,N_13435);
xor U14050 (N_14050,N_12956,N_13089);
nor U14051 (N_14051,N_12660,N_12152);
nor U14052 (N_14052,N_12986,N_13064);
and U14053 (N_14053,N_12823,N_12334);
xnor U14054 (N_14054,N_12657,N_13213);
xnor U14055 (N_14055,N_12960,N_12834);
xnor U14056 (N_14056,N_13247,N_13165);
or U14057 (N_14057,N_12440,N_12408);
nand U14058 (N_14058,N_12995,N_12367);
nor U14059 (N_14059,N_12070,N_12977);
nor U14060 (N_14060,N_13036,N_13112);
and U14061 (N_14061,N_13014,N_12052);
nor U14062 (N_14062,N_13079,N_13378);
or U14063 (N_14063,N_12902,N_12883);
and U14064 (N_14064,N_12481,N_13063);
nand U14065 (N_14065,N_13188,N_13433);
and U14066 (N_14066,N_12427,N_12722);
or U14067 (N_14067,N_12778,N_12221);
nand U14068 (N_14068,N_13180,N_12473);
nand U14069 (N_14069,N_12713,N_12534);
nand U14070 (N_14070,N_12833,N_12681);
nor U14071 (N_14071,N_12416,N_13232);
xnor U14072 (N_14072,N_13037,N_12925);
or U14073 (N_14073,N_12890,N_13321);
nand U14074 (N_14074,N_12108,N_12628);
or U14075 (N_14075,N_12291,N_12175);
or U14076 (N_14076,N_12663,N_12707);
nor U14077 (N_14077,N_13172,N_12590);
nor U14078 (N_14078,N_12748,N_12091);
nand U14079 (N_14079,N_13498,N_12510);
nand U14080 (N_14080,N_12136,N_12080);
nor U14081 (N_14081,N_12768,N_12131);
and U14082 (N_14082,N_13383,N_12040);
nor U14083 (N_14083,N_12656,N_13215);
nor U14084 (N_14084,N_12733,N_12915);
nand U14085 (N_14085,N_12929,N_13374);
and U14086 (N_14086,N_13404,N_13340);
nor U14087 (N_14087,N_12494,N_13299);
and U14088 (N_14088,N_12453,N_12075);
xnor U14089 (N_14089,N_12229,N_13429);
nand U14090 (N_14090,N_12437,N_12582);
nand U14091 (N_14091,N_13280,N_12610);
nand U14092 (N_14092,N_12278,N_12868);
and U14093 (N_14093,N_12564,N_12575);
or U14094 (N_14094,N_12146,N_12297);
nor U14095 (N_14095,N_13009,N_12189);
and U14096 (N_14096,N_12993,N_12350);
nand U14097 (N_14097,N_12765,N_13373);
nand U14098 (N_14098,N_13122,N_13268);
and U14099 (N_14099,N_13322,N_12033);
xnor U14100 (N_14100,N_12932,N_12866);
and U14101 (N_14101,N_12144,N_13067);
or U14102 (N_14102,N_12862,N_13080);
and U14103 (N_14103,N_12691,N_13376);
nand U14104 (N_14104,N_12255,N_12365);
nor U14105 (N_14105,N_12405,N_12984);
or U14106 (N_14106,N_12997,N_12322);
xnor U14107 (N_14107,N_12431,N_13073);
nand U14108 (N_14108,N_13186,N_12867);
nand U14109 (N_14109,N_13315,N_13353);
or U14110 (N_14110,N_12982,N_12892);
or U14111 (N_14111,N_13317,N_12648);
xor U14112 (N_14112,N_12077,N_12447);
or U14113 (N_14113,N_12633,N_13082);
xor U14114 (N_14114,N_12753,N_13410);
and U14115 (N_14115,N_12991,N_13058);
nor U14116 (N_14116,N_13220,N_12288);
nand U14117 (N_14117,N_12236,N_13226);
nand U14118 (N_14118,N_12552,N_12786);
xor U14119 (N_14119,N_12217,N_13113);
and U14120 (N_14120,N_12912,N_12178);
and U14121 (N_14121,N_13431,N_13140);
xor U14122 (N_14122,N_13184,N_12568);
nand U14123 (N_14123,N_12906,N_13225);
xor U14124 (N_14124,N_13480,N_12668);
xnor U14125 (N_14125,N_12269,N_12196);
nor U14126 (N_14126,N_13454,N_12233);
nor U14127 (N_14127,N_13228,N_13210);
nand U14128 (N_14128,N_12600,N_12934);
or U14129 (N_14129,N_12250,N_12154);
or U14130 (N_14130,N_12754,N_13439);
and U14131 (N_14131,N_13300,N_13363);
and U14132 (N_14132,N_13031,N_12780);
or U14133 (N_14133,N_13096,N_12567);
nor U14134 (N_14134,N_13148,N_12063);
xnor U14135 (N_14135,N_12190,N_12364);
xnor U14136 (N_14136,N_12121,N_12983);
and U14137 (N_14137,N_12097,N_13395);
xnor U14138 (N_14138,N_12909,N_12007);
or U14139 (N_14139,N_12283,N_12704);
xor U14140 (N_14140,N_12630,N_12517);
nand U14141 (N_14141,N_13208,N_13021);
nor U14142 (N_14142,N_12715,N_12441);
nand U14143 (N_14143,N_12208,N_12333);
or U14144 (N_14144,N_12356,N_13331);
nor U14145 (N_14145,N_12170,N_12393);
nand U14146 (N_14146,N_12218,N_12675);
nand U14147 (N_14147,N_12206,N_13293);
and U14148 (N_14148,N_12788,N_13414);
xnor U14149 (N_14149,N_13015,N_13499);
nand U14150 (N_14150,N_12574,N_13030);
nand U14151 (N_14151,N_12102,N_12939);
nor U14152 (N_14152,N_13173,N_13230);
nor U14153 (N_14153,N_13115,N_13473);
nand U14154 (N_14154,N_12959,N_12489);
and U14155 (N_14155,N_13462,N_13358);
or U14156 (N_14156,N_12420,N_12706);
nor U14157 (N_14157,N_12802,N_12665);
or U14158 (N_14158,N_12341,N_12914);
nand U14159 (N_14159,N_13117,N_13104);
xor U14160 (N_14160,N_13087,N_12895);
nand U14161 (N_14161,N_13445,N_12242);
nor U14162 (N_14162,N_13242,N_13441);
xnor U14163 (N_14163,N_13314,N_13144);
xor U14164 (N_14164,N_13069,N_12411);
nor U14165 (N_14165,N_12672,N_12459);
and U14166 (N_14166,N_13256,N_12262);
nand U14167 (N_14167,N_13337,N_12714);
nand U14168 (N_14168,N_12985,N_12652);
xnor U14169 (N_14169,N_12403,N_12969);
nor U14170 (N_14170,N_13357,N_12641);
nand U14171 (N_14171,N_13326,N_13072);
nor U14172 (N_14172,N_12772,N_12618);
nor U14173 (N_14173,N_13330,N_12547);
nand U14174 (N_14174,N_12089,N_12182);
or U14175 (N_14175,N_12678,N_12301);
and U14176 (N_14176,N_12009,N_13375);
nor U14177 (N_14177,N_12813,N_13286);
and U14178 (N_14178,N_13222,N_12142);
and U14179 (N_14179,N_12153,N_12800);
nand U14180 (N_14180,N_12889,N_13287);
xnor U14181 (N_14181,N_13351,N_13038);
xnor U14182 (N_14182,N_12597,N_12566);
nand U14183 (N_14183,N_12074,N_12137);
and U14184 (N_14184,N_13497,N_12874);
xnor U14185 (N_14185,N_12203,N_13158);
xnor U14186 (N_14186,N_13050,N_12538);
xnor U14187 (N_14187,N_12237,N_12438);
nor U14188 (N_14188,N_12745,N_12927);
nor U14189 (N_14189,N_12377,N_12466);
nand U14190 (N_14190,N_12205,N_13261);
or U14191 (N_14191,N_12572,N_12666);
nor U14192 (N_14192,N_13057,N_12899);
xor U14193 (N_14193,N_12382,N_13097);
nand U14194 (N_14194,N_12718,N_13359);
nor U14195 (N_14195,N_12730,N_13478);
nor U14196 (N_14196,N_13368,N_13297);
nor U14197 (N_14197,N_12843,N_12981);
nand U14198 (N_14198,N_12337,N_12817);
nand U14199 (N_14199,N_13438,N_12764);
nor U14200 (N_14200,N_12637,N_12158);
or U14201 (N_14201,N_13185,N_13008);
nor U14202 (N_14202,N_12717,N_12433);
nand U14203 (N_14203,N_12785,N_12093);
nand U14204 (N_14204,N_12140,N_12528);
and U14205 (N_14205,N_12173,N_12671);
or U14206 (N_14206,N_13049,N_12114);
or U14207 (N_14207,N_12931,N_12549);
nor U14208 (N_14208,N_12581,N_13394);
nand U14209 (N_14209,N_12461,N_12623);
nor U14210 (N_14210,N_12687,N_13479);
nand U14211 (N_14211,N_12904,N_12418);
xor U14212 (N_14212,N_13007,N_12626);
nor U14213 (N_14213,N_13289,N_13054);
nand U14214 (N_14214,N_13147,N_12426);
nor U14215 (N_14215,N_12404,N_12822);
xnor U14216 (N_14216,N_12771,N_12793);
or U14217 (N_14217,N_12792,N_13361);
nor U14218 (N_14218,N_13204,N_12601);
xor U14219 (N_14219,N_13095,N_12725);
nor U14220 (N_14220,N_13275,N_12911);
and U14221 (N_14221,N_13437,N_12271);
or U14222 (N_14222,N_12655,N_12325);
xnor U14223 (N_14223,N_12157,N_12389);
nor U14224 (N_14224,N_12850,N_12307);
nor U14225 (N_14225,N_12962,N_12728);
and U14226 (N_14226,N_12122,N_13421);
nor U14227 (N_14227,N_13260,N_12830);
xor U14228 (N_14228,N_12141,N_13083);
nor U14229 (N_14229,N_12670,N_12413);
nor U14230 (N_14230,N_12825,N_13101);
nand U14231 (N_14231,N_13291,N_12757);
nand U14232 (N_14232,N_12130,N_13295);
or U14233 (N_14233,N_13166,N_12132);
or U14234 (N_14234,N_12746,N_12224);
nor U14235 (N_14235,N_12885,N_12352);
or U14236 (N_14236,N_12162,N_12187);
nor U14237 (N_14237,N_12688,N_12424);
and U14238 (N_14238,N_12168,N_12428);
xnor U14239 (N_14239,N_13042,N_12797);
or U14240 (N_14240,N_12923,N_13119);
xor U14241 (N_14241,N_13020,N_12450);
or U14242 (N_14242,N_12439,N_13334);
and U14243 (N_14243,N_12685,N_12267);
xnor U14244 (N_14244,N_12616,N_12870);
and U14245 (N_14245,N_13198,N_12071);
or U14246 (N_14246,N_13044,N_13482);
nand U14247 (N_14247,N_12592,N_12303);
nor U14248 (N_14248,N_12415,N_13489);
xnor U14249 (N_14249,N_12312,N_12487);
nor U14250 (N_14250,N_12481,N_13446);
nor U14251 (N_14251,N_13019,N_12037);
xnor U14252 (N_14252,N_12818,N_12974);
and U14253 (N_14253,N_13083,N_12298);
nand U14254 (N_14254,N_12339,N_13374);
or U14255 (N_14255,N_13425,N_12231);
nor U14256 (N_14256,N_12329,N_13140);
xor U14257 (N_14257,N_12248,N_12992);
nor U14258 (N_14258,N_12575,N_12550);
xor U14259 (N_14259,N_13023,N_13254);
nand U14260 (N_14260,N_12102,N_12008);
xnor U14261 (N_14261,N_13288,N_13045);
or U14262 (N_14262,N_12801,N_13077);
nor U14263 (N_14263,N_12340,N_12349);
or U14264 (N_14264,N_12948,N_12215);
nor U14265 (N_14265,N_12271,N_12107);
nor U14266 (N_14266,N_12264,N_12880);
xnor U14267 (N_14267,N_12310,N_13481);
and U14268 (N_14268,N_12193,N_13157);
or U14269 (N_14269,N_12083,N_12116);
and U14270 (N_14270,N_12409,N_12375);
or U14271 (N_14271,N_12809,N_12720);
xnor U14272 (N_14272,N_13435,N_13187);
nand U14273 (N_14273,N_13320,N_12224);
and U14274 (N_14274,N_12883,N_13241);
xnor U14275 (N_14275,N_12771,N_12355);
or U14276 (N_14276,N_13454,N_13451);
nand U14277 (N_14277,N_12306,N_12063);
or U14278 (N_14278,N_12194,N_12697);
nor U14279 (N_14279,N_13120,N_12393);
nor U14280 (N_14280,N_12360,N_12804);
or U14281 (N_14281,N_12644,N_13367);
or U14282 (N_14282,N_13053,N_13170);
nor U14283 (N_14283,N_12908,N_12803);
or U14284 (N_14284,N_12029,N_13338);
nand U14285 (N_14285,N_13126,N_13239);
xor U14286 (N_14286,N_12806,N_12781);
or U14287 (N_14287,N_13277,N_12372);
nand U14288 (N_14288,N_12627,N_12409);
nor U14289 (N_14289,N_13183,N_13184);
nand U14290 (N_14290,N_12536,N_13034);
or U14291 (N_14291,N_12247,N_12762);
nand U14292 (N_14292,N_12691,N_12555);
nor U14293 (N_14293,N_12492,N_12653);
nor U14294 (N_14294,N_12705,N_12874);
nor U14295 (N_14295,N_12016,N_12646);
xnor U14296 (N_14296,N_13398,N_12495);
xor U14297 (N_14297,N_13018,N_13342);
nor U14298 (N_14298,N_12023,N_12933);
nor U14299 (N_14299,N_12022,N_12966);
xnor U14300 (N_14300,N_12478,N_13202);
or U14301 (N_14301,N_13035,N_12896);
xor U14302 (N_14302,N_12444,N_13255);
nand U14303 (N_14303,N_12076,N_12150);
xor U14304 (N_14304,N_13085,N_13154);
nand U14305 (N_14305,N_13482,N_12239);
and U14306 (N_14306,N_12335,N_12101);
nand U14307 (N_14307,N_13465,N_12420);
nor U14308 (N_14308,N_12231,N_13170);
nand U14309 (N_14309,N_12572,N_13176);
and U14310 (N_14310,N_12857,N_12211);
nand U14311 (N_14311,N_12535,N_12730);
xor U14312 (N_14312,N_13471,N_12054);
xnor U14313 (N_14313,N_13170,N_12673);
nand U14314 (N_14314,N_13415,N_13450);
and U14315 (N_14315,N_12676,N_12060);
xnor U14316 (N_14316,N_13101,N_12797);
nand U14317 (N_14317,N_12143,N_12463);
nor U14318 (N_14318,N_13067,N_12803);
nand U14319 (N_14319,N_13487,N_13165);
nand U14320 (N_14320,N_13004,N_13321);
or U14321 (N_14321,N_13322,N_12839);
or U14322 (N_14322,N_12787,N_12422);
or U14323 (N_14323,N_13174,N_12111);
or U14324 (N_14324,N_13273,N_12421);
or U14325 (N_14325,N_13185,N_12720);
and U14326 (N_14326,N_12427,N_13163);
nor U14327 (N_14327,N_12597,N_12579);
nand U14328 (N_14328,N_13430,N_12895);
nor U14329 (N_14329,N_12333,N_13221);
and U14330 (N_14330,N_13019,N_12484);
and U14331 (N_14331,N_12540,N_12925);
xor U14332 (N_14332,N_12844,N_12293);
and U14333 (N_14333,N_13457,N_13120);
and U14334 (N_14334,N_12286,N_13439);
xor U14335 (N_14335,N_13352,N_13002);
xor U14336 (N_14336,N_12029,N_12688);
nand U14337 (N_14337,N_12304,N_12662);
and U14338 (N_14338,N_12671,N_12334);
nand U14339 (N_14339,N_13250,N_13020);
or U14340 (N_14340,N_12809,N_12124);
nand U14341 (N_14341,N_12575,N_12585);
nor U14342 (N_14342,N_13499,N_12685);
nand U14343 (N_14343,N_13444,N_13149);
xnor U14344 (N_14344,N_12465,N_13438);
nand U14345 (N_14345,N_13294,N_12953);
xor U14346 (N_14346,N_12281,N_13178);
nand U14347 (N_14347,N_12437,N_12399);
xnor U14348 (N_14348,N_12156,N_13067);
or U14349 (N_14349,N_12499,N_13429);
xnor U14350 (N_14350,N_12804,N_12700);
or U14351 (N_14351,N_12733,N_13104);
or U14352 (N_14352,N_13133,N_12156);
and U14353 (N_14353,N_12048,N_13096);
xnor U14354 (N_14354,N_12112,N_13497);
nand U14355 (N_14355,N_12888,N_13141);
nor U14356 (N_14356,N_12512,N_12778);
nor U14357 (N_14357,N_12545,N_12187);
or U14358 (N_14358,N_12849,N_12161);
nand U14359 (N_14359,N_12161,N_13457);
nor U14360 (N_14360,N_13379,N_12718);
and U14361 (N_14361,N_12415,N_12998);
xnor U14362 (N_14362,N_12714,N_12621);
nor U14363 (N_14363,N_12163,N_13168);
nor U14364 (N_14364,N_12168,N_12669);
xor U14365 (N_14365,N_12536,N_12239);
nor U14366 (N_14366,N_12778,N_12715);
nor U14367 (N_14367,N_12101,N_12818);
xnor U14368 (N_14368,N_13441,N_13468);
nand U14369 (N_14369,N_12473,N_12831);
nor U14370 (N_14370,N_12076,N_12197);
or U14371 (N_14371,N_13268,N_13399);
or U14372 (N_14372,N_13486,N_13244);
or U14373 (N_14373,N_12245,N_12704);
and U14374 (N_14374,N_12899,N_13080);
nand U14375 (N_14375,N_12392,N_13415);
or U14376 (N_14376,N_12609,N_12970);
and U14377 (N_14377,N_12266,N_12364);
nor U14378 (N_14378,N_13369,N_13289);
or U14379 (N_14379,N_13202,N_12707);
nand U14380 (N_14380,N_13187,N_12118);
xnor U14381 (N_14381,N_12055,N_12973);
nand U14382 (N_14382,N_13272,N_13314);
nand U14383 (N_14383,N_12108,N_12341);
xnor U14384 (N_14384,N_13396,N_12034);
nor U14385 (N_14385,N_12939,N_13447);
or U14386 (N_14386,N_13298,N_12118);
nand U14387 (N_14387,N_12244,N_12081);
and U14388 (N_14388,N_12966,N_13427);
nand U14389 (N_14389,N_12875,N_13472);
nor U14390 (N_14390,N_12349,N_13415);
and U14391 (N_14391,N_12908,N_12692);
nor U14392 (N_14392,N_12956,N_13215);
and U14393 (N_14393,N_13323,N_12996);
and U14394 (N_14394,N_12922,N_13157);
or U14395 (N_14395,N_13471,N_12649);
xor U14396 (N_14396,N_12658,N_12220);
nor U14397 (N_14397,N_12224,N_12584);
or U14398 (N_14398,N_13340,N_12507);
xor U14399 (N_14399,N_12454,N_13032);
nor U14400 (N_14400,N_12727,N_13198);
and U14401 (N_14401,N_13018,N_12223);
nor U14402 (N_14402,N_13193,N_12650);
xnor U14403 (N_14403,N_12106,N_12596);
nand U14404 (N_14404,N_12499,N_12615);
and U14405 (N_14405,N_13198,N_12414);
nand U14406 (N_14406,N_13071,N_12048);
nand U14407 (N_14407,N_12512,N_12085);
xnor U14408 (N_14408,N_13275,N_12979);
nand U14409 (N_14409,N_12774,N_12727);
and U14410 (N_14410,N_12666,N_12109);
xnor U14411 (N_14411,N_13280,N_12405);
nor U14412 (N_14412,N_12619,N_13410);
nand U14413 (N_14413,N_12874,N_12122);
or U14414 (N_14414,N_13375,N_12268);
and U14415 (N_14415,N_12982,N_12279);
nand U14416 (N_14416,N_12150,N_12431);
nand U14417 (N_14417,N_12636,N_13245);
nor U14418 (N_14418,N_12574,N_12139);
nand U14419 (N_14419,N_12936,N_12192);
or U14420 (N_14420,N_13209,N_13271);
nor U14421 (N_14421,N_13441,N_12305);
nor U14422 (N_14422,N_13356,N_13248);
nor U14423 (N_14423,N_12313,N_12695);
nor U14424 (N_14424,N_12229,N_13142);
nand U14425 (N_14425,N_13454,N_13375);
xor U14426 (N_14426,N_13428,N_12389);
nor U14427 (N_14427,N_13247,N_12994);
and U14428 (N_14428,N_13418,N_13312);
xnor U14429 (N_14429,N_12053,N_12890);
and U14430 (N_14430,N_12490,N_12904);
or U14431 (N_14431,N_13289,N_13039);
nor U14432 (N_14432,N_12123,N_13468);
and U14433 (N_14433,N_12866,N_12563);
nand U14434 (N_14434,N_12935,N_12637);
or U14435 (N_14435,N_12342,N_12773);
nor U14436 (N_14436,N_12603,N_13364);
or U14437 (N_14437,N_12890,N_12730);
xnor U14438 (N_14438,N_12234,N_12711);
xor U14439 (N_14439,N_12757,N_12355);
nand U14440 (N_14440,N_12549,N_12981);
nand U14441 (N_14441,N_12744,N_12559);
nand U14442 (N_14442,N_12800,N_12261);
and U14443 (N_14443,N_13012,N_12697);
or U14444 (N_14444,N_13401,N_13043);
nand U14445 (N_14445,N_12033,N_13246);
and U14446 (N_14446,N_13468,N_12461);
and U14447 (N_14447,N_13306,N_13489);
nor U14448 (N_14448,N_12404,N_12218);
nand U14449 (N_14449,N_13025,N_12460);
nor U14450 (N_14450,N_12284,N_13113);
and U14451 (N_14451,N_12451,N_13205);
or U14452 (N_14452,N_12466,N_13138);
and U14453 (N_14453,N_12510,N_13017);
and U14454 (N_14454,N_12050,N_13029);
nand U14455 (N_14455,N_12669,N_12973);
nor U14456 (N_14456,N_12088,N_13333);
and U14457 (N_14457,N_12517,N_12698);
and U14458 (N_14458,N_13028,N_13461);
and U14459 (N_14459,N_12348,N_12954);
or U14460 (N_14460,N_12886,N_13229);
xnor U14461 (N_14461,N_12429,N_12824);
xnor U14462 (N_14462,N_12069,N_12688);
nor U14463 (N_14463,N_12361,N_12905);
nand U14464 (N_14464,N_13283,N_13291);
xnor U14465 (N_14465,N_13198,N_12804);
nor U14466 (N_14466,N_12803,N_13290);
and U14467 (N_14467,N_12583,N_13435);
nor U14468 (N_14468,N_12869,N_12333);
or U14469 (N_14469,N_12764,N_12087);
nand U14470 (N_14470,N_12517,N_12290);
xor U14471 (N_14471,N_12136,N_13269);
and U14472 (N_14472,N_13120,N_13478);
xor U14473 (N_14473,N_12450,N_13253);
or U14474 (N_14474,N_12167,N_12873);
xor U14475 (N_14475,N_13278,N_13000);
or U14476 (N_14476,N_12644,N_13001);
nand U14477 (N_14477,N_12975,N_13258);
nor U14478 (N_14478,N_13335,N_12782);
or U14479 (N_14479,N_12014,N_13253);
nand U14480 (N_14480,N_12314,N_13252);
and U14481 (N_14481,N_12171,N_12642);
and U14482 (N_14482,N_12461,N_13129);
nand U14483 (N_14483,N_13258,N_13060);
and U14484 (N_14484,N_13077,N_12674);
xor U14485 (N_14485,N_12547,N_13362);
or U14486 (N_14486,N_13329,N_12118);
or U14487 (N_14487,N_13391,N_12852);
xnor U14488 (N_14488,N_12106,N_12584);
and U14489 (N_14489,N_13085,N_13371);
or U14490 (N_14490,N_12141,N_13154);
or U14491 (N_14491,N_13072,N_12897);
and U14492 (N_14492,N_12194,N_13408);
nand U14493 (N_14493,N_13062,N_13465);
xor U14494 (N_14494,N_13313,N_12800);
nor U14495 (N_14495,N_12162,N_12188);
nand U14496 (N_14496,N_13084,N_12891);
and U14497 (N_14497,N_12522,N_12436);
nor U14498 (N_14498,N_12965,N_12520);
nand U14499 (N_14499,N_12115,N_13441);
or U14500 (N_14500,N_13220,N_13050);
or U14501 (N_14501,N_13468,N_13236);
or U14502 (N_14502,N_13383,N_13126);
nor U14503 (N_14503,N_12490,N_12809);
nand U14504 (N_14504,N_13346,N_12983);
or U14505 (N_14505,N_12524,N_12275);
or U14506 (N_14506,N_13305,N_13267);
xor U14507 (N_14507,N_12723,N_12426);
and U14508 (N_14508,N_12770,N_12112);
or U14509 (N_14509,N_12620,N_13163);
and U14510 (N_14510,N_12862,N_12904);
or U14511 (N_14511,N_13054,N_13229);
and U14512 (N_14512,N_13198,N_12486);
xnor U14513 (N_14513,N_12294,N_12884);
nand U14514 (N_14514,N_12499,N_13170);
nand U14515 (N_14515,N_13392,N_12542);
nand U14516 (N_14516,N_12011,N_12012);
nor U14517 (N_14517,N_12749,N_12415);
nand U14518 (N_14518,N_13457,N_12145);
xnor U14519 (N_14519,N_13147,N_13021);
or U14520 (N_14520,N_12128,N_13293);
and U14521 (N_14521,N_12082,N_12505);
xor U14522 (N_14522,N_12548,N_12982);
nand U14523 (N_14523,N_13081,N_12200);
nor U14524 (N_14524,N_12791,N_12851);
or U14525 (N_14525,N_13475,N_12007);
xor U14526 (N_14526,N_13462,N_12907);
or U14527 (N_14527,N_12102,N_12249);
or U14528 (N_14528,N_13043,N_12551);
or U14529 (N_14529,N_13255,N_12140);
nor U14530 (N_14530,N_12363,N_12405);
and U14531 (N_14531,N_13217,N_13424);
xnor U14532 (N_14532,N_13120,N_12536);
nand U14533 (N_14533,N_12661,N_12684);
nand U14534 (N_14534,N_12526,N_13196);
xor U14535 (N_14535,N_13496,N_12463);
nand U14536 (N_14536,N_13127,N_12499);
or U14537 (N_14537,N_12259,N_13450);
xnor U14538 (N_14538,N_12458,N_13057);
xor U14539 (N_14539,N_13014,N_12738);
or U14540 (N_14540,N_12981,N_12034);
or U14541 (N_14541,N_12005,N_12082);
nor U14542 (N_14542,N_13467,N_12838);
xnor U14543 (N_14543,N_13209,N_13118);
nor U14544 (N_14544,N_13284,N_13075);
xnor U14545 (N_14545,N_12167,N_12434);
xnor U14546 (N_14546,N_12754,N_12257);
and U14547 (N_14547,N_12636,N_12416);
nand U14548 (N_14548,N_12879,N_13101);
xor U14549 (N_14549,N_12654,N_12371);
xor U14550 (N_14550,N_12342,N_13436);
xnor U14551 (N_14551,N_12314,N_13497);
nor U14552 (N_14552,N_12197,N_12840);
xor U14553 (N_14553,N_12279,N_12975);
or U14554 (N_14554,N_12140,N_13201);
and U14555 (N_14555,N_13344,N_12299);
or U14556 (N_14556,N_12202,N_12521);
nor U14557 (N_14557,N_13146,N_13314);
and U14558 (N_14558,N_13070,N_12112);
and U14559 (N_14559,N_13466,N_13105);
nor U14560 (N_14560,N_12424,N_12430);
nor U14561 (N_14561,N_12413,N_12388);
or U14562 (N_14562,N_12492,N_12564);
nand U14563 (N_14563,N_13246,N_13349);
or U14564 (N_14564,N_12382,N_12915);
and U14565 (N_14565,N_12578,N_12113);
nand U14566 (N_14566,N_12484,N_13047);
nand U14567 (N_14567,N_13091,N_12014);
and U14568 (N_14568,N_13292,N_12642);
or U14569 (N_14569,N_13426,N_13280);
nand U14570 (N_14570,N_12876,N_13046);
or U14571 (N_14571,N_12617,N_12804);
nand U14572 (N_14572,N_12527,N_12423);
or U14573 (N_14573,N_13156,N_12189);
or U14574 (N_14574,N_13358,N_13315);
and U14575 (N_14575,N_12464,N_13091);
nand U14576 (N_14576,N_13406,N_12400);
or U14577 (N_14577,N_12170,N_12093);
or U14578 (N_14578,N_12541,N_12356);
or U14579 (N_14579,N_12263,N_12532);
or U14580 (N_14580,N_13314,N_13402);
or U14581 (N_14581,N_12144,N_12545);
and U14582 (N_14582,N_13283,N_13047);
xor U14583 (N_14583,N_12119,N_12338);
or U14584 (N_14584,N_13159,N_13273);
xnor U14585 (N_14585,N_12058,N_12181);
and U14586 (N_14586,N_13341,N_13219);
xnor U14587 (N_14587,N_12635,N_13339);
and U14588 (N_14588,N_12298,N_12076);
nand U14589 (N_14589,N_12678,N_12055);
or U14590 (N_14590,N_13100,N_12661);
xor U14591 (N_14591,N_12692,N_12431);
or U14592 (N_14592,N_13085,N_12496);
or U14593 (N_14593,N_13004,N_12455);
nor U14594 (N_14594,N_12111,N_12479);
nor U14595 (N_14595,N_13270,N_13124);
nand U14596 (N_14596,N_13252,N_13186);
or U14597 (N_14597,N_13000,N_13386);
nor U14598 (N_14598,N_12974,N_12065);
nor U14599 (N_14599,N_12871,N_13226);
nor U14600 (N_14600,N_12680,N_13085);
and U14601 (N_14601,N_12102,N_13492);
xor U14602 (N_14602,N_12111,N_12173);
xnor U14603 (N_14603,N_12669,N_12156);
nand U14604 (N_14604,N_12623,N_12149);
and U14605 (N_14605,N_12863,N_12435);
nor U14606 (N_14606,N_12802,N_12770);
nand U14607 (N_14607,N_12593,N_12897);
and U14608 (N_14608,N_12401,N_12404);
xor U14609 (N_14609,N_13237,N_13182);
nand U14610 (N_14610,N_12205,N_13224);
nand U14611 (N_14611,N_13099,N_12621);
nor U14612 (N_14612,N_12592,N_13288);
xnor U14613 (N_14613,N_13012,N_12017);
xor U14614 (N_14614,N_12764,N_13061);
and U14615 (N_14615,N_12731,N_12582);
nand U14616 (N_14616,N_13022,N_12146);
and U14617 (N_14617,N_12112,N_12717);
or U14618 (N_14618,N_12578,N_12467);
and U14619 (N_14619,N_12929,N_12860);
and U14620 (N_14620,N_12052,N_12557);
and U14621 (N_14621,N_13064,N_12535);
xnor U14622 (N_14622,N_12632,N_12902);
xnor U14623 (N_14623,N_12569,N_12218);
nand U14624 (N_14624,N_13185,N_12894);
or U14625 (N_14625,N_13488,N_12405);
nor U14626 (N_14626,N_13385,N_12021);
xnor U14627 (N_14627,N_13132,N_12347);
or U14628 (N_14628,N_12220,N_12213);
nand U14629 (N_14629,N_12375,N_12688);
or U14630 (N_14630,N_13039,N_13120);
or U14631 (N_14631,N_12654,N_12290);
nor U14632 (N_14632,N_12921,N_12910);
or U14633 (N_14633,N_12031,N_12126);
nand U14634 (N_14634,N_12585,N_12170);
nand U14635 (N_14635,N_13243,N_12520);
and U14636 (N_14636,N_12812,N_12513);
xor U14637 (N_14637,N_13099,N_13368);
nor U14638 (N_14638,N_12652,N_13045);
nand U14639 (N_14639,N_13097,N_12686);
xnor U14640 (N_14640,N_12608,N_13134);
and U14641 (N_14641,N_13227,N_12931);
nor U14642 (N_14642,N_13237,N_12592);
nand U14643 (N_14643,N_13407,N_12764);
nand U14644 (N_14644,N_12325,N_12806);
and U14645 (N_14645,N_12374,N_13290);
or U14646 (N_14646,N_12342,N_12010);
and U14647 (N_14647,N_12405,N_12727);
nor U14648 (N_14648,N_12630,N_13208);
nor U14649 (N_14649,N_13101,N_12962);
nor U14650 (N_14650,N_12508,N_12870);
nor U14651 (N_14651,N_12341,N_12102);
xor U14652 (N_14652,N_12224,N_12975);
xor U14653 (N_14653,N_12765,N_12911);
nand U14654 (N_14654,N_12046,N_12270);
nand U14655 (N_14655,N_13367,N_12975);
or U14656 (N_14656,N_12668,N_13313);
or U14657 (N_14657,N_12070,N_12438);
nand U14658 (N_14658,N_13352,N_13014);
nand U14659 (N_14659,N_12671,N_12117);
or U14660 (N_14660,N_13281,N_13018);
xnor U14661 (N_14661,N_13430,N_12916);
xnor U14662 (N_14662,N_12621,N_13045);
nor U14663 (N_14663,N_13374,N_12659);
nor U14664 (N_14664,N_12619,N_12249);
xnor U14665 (N_14665,N_12708,N_13329);
nand U14666 (N_14666,N_13240,N_12816);
and U14667 (N_14667,N_13065,N_12322);
xnor U14668 (N_14668,N_12696,N_12603);
and U14669 (N_14669,N_12895,N_13247);
nor U14670 (N_14670,N_12438,N_13212);
or U14671 (N_14671,N_12429,N_13285);
xnor U14672 (N_14672,N_12742,N_12112);
nor U14673 (N_14673,N_12829,N_12509);
nand U14674 (N_14674,N_13018,N_12016);
nor U14675 (N_14675,N_12297,N_13184);
xor U14676 (N_14676,N_12706,N_12956);
and U14677 (N_14677,N_12922,N_12125);
nor U14678 (N_14678,N_13398,N_12432);
or U14679 (N_14679,N_13013,N_13292);
and U14680 (N_14680,N_12004,N_12079);
and U14681 (N_14681,N_12446,N_13010);
and U14682 (N_14682,N_13479,N_12878);
nor U14683 (N_14683,N_12618,N_13377);
xor U14684 (N_14684,N_12106,N_13394);
nand U14685 (N_14685,N_12326,N_12074);
nor U14686 (N_14686,N_12401,N_13465);
xnor U14687 (N_14687,N_12218,N_12627);
or U14688 (N_14688,N_12251,N_12581);
nor U14689 (N_14689,N_12309,N_13308);
xnor U14690 (N_14690,N_12255,N_12249);
nand U14691 (N_14691,N_12035,N_12456);
nor U14692 (N_14692,N_12390,N_12623);
xor U14693 (N_14693,N_12269,N_13075);
nand U14694 (N_14694,N_13366,N_13361);
and U14695 (N_14695,N_12535,N_12373);
xor U14696 (N_14696,N_12872,N_13196);
nor U14697 (N_14697,N_13015,N_13271);
nand U14698 (N_14698,N_12278,N_12831);
or U14699 (N_14699,N_12355,N_13310);
and U14700 (N_14700,N_12475,N_12644);
and U14701 (N_14701,N_12957,N_13129);
nor U14702 (N_14702,N_12173,N_12985);
nor U14703 (N_14703,N_12665,N_12946);
or U14704 (N_14704,N_12058,N_12963);
nor U14705 (N_14705,N_12601,N_12113);
or U14706 (N_14706,N_13346,N_12876);
nand U14707 (N_14707,N_12256,N_13217);
nor U14708 (N_14708,N_13071,N_13079);
and U14709 (N_14709,N_13286,N_12715);
or U14710 (N_14710,N_12658,N_13059);
nor U14711 (N_14711,N_12790,N_13077);
nor U14712 (N_14712,N_12006,N_12822);
and U14713 (N_14713,N_12478,N_13351);
nand U14714 (N_14714,N_12405,N_13028);
nor U14715 (N_14715,N_12849,N_12860);
or U14716 (N_14716,N_12489,N_12039);
nor U14717 (N_14717,N_12020,N_12380);
and U14718 (N_14718,N_13044,N_12198);
and U14719 (N_14719,N_12407,N_12243);
or U14720 (N_14720,N_12090,N_12984);
or U14721 (N_14721,N_12806,N_13493);
or U14722 (N_14722,N_12882,N_12723);
xor U14723 (N_14723,N_13439,N_12791);
and U14724 (N_14724,N_13365,N_13237);
and U14725 (N_14725,N_13367,N_13095);
and U14726 (N_14726,N_12047,N_12817);
xor U14727 (N_14727,N_12147,N_12596);
nor U14728 (N_14728,N_12872,N_13067);
and U14729 (N_14729,N_12004,N_12847);
xor U14730 (N_14730,N_13386,N_12384);
xnor U14731 (N_14731,N_13006,N_12423);
xnor U14732 (N_14732,N_12754,N_12990);
xor U14733 (N_14733,N_12400,N_12313);
xor U14734 (N_14734,N_12412,N_12389);
nand U14735 (N_14735,N_12799,N_12861);
xor U14736 (N_14736,N_13144,N_13287);
and U14737 (N_14737,N_12347,N_12093);
xor U14738 (N_14738,N_13118,N_12648);
nor U14739 (N_14739,N_12452,N_12334);
or U14740 (N_14740,N_12861,N_12123);
and U14741 (N_14741,N_12829,N_12622);
or U14742 (N_14742,N_12495,N_12741);
nand U14743 (N_14743,N_13129,N_13212);
or U14744 (N_14744,N_12463,N_12880);
nand U14745 (N_14745,N_13395,N_13071);
nor U14746 (N_14746,N_13320,N_13114);
and U14747 (N_14747,N_12476,N_12330);
nand U14748 (N_14748,N_12516,N_13280);
nand U14749 (N_14749,N_13291,N_12917);
nor U14750 (N_14750,N_12155,N_12185);
xor U14751 (N_14751,N_12755,N_12726);
or U14752 (N_14752,N_13236,N_13349);
nor U14753 (N_14753,N_13464,N_12685);
nor U14754 (N_14754,N_12946,N_12411);
or U14755 (N_14755,N_12232,N_12804);
xor U14756 (N_14756,N_13315,N_12477);
or U14757 (N_14757,N_13070,N_13494);
xor U14758 (N_14758,N_12431,N_13190);
or U14759 (N_14759,N_12284,N_13105);
and U14760 (N_14760,N_13142,N_13429);
xnor U14761 (N_14761,N_12043,N_13491);
and U14762 (N_14762,N_13178,N_12251);
nand U14763 (N_14763,N_13336,N_12969);
or U14764 (N_14764,N_13370,N_12015);
and U14765 (N_14765,N_12977,N_12207);
nor U14766 (N_14766,N_13103,N_13019);
xor U14767 (N_14767,N_12783,N_12579);
and U14768 (N_14768,N_12362,N_13229);
nor U14769 (N_14769,N_12311,N_13419);
and U14770 (N_14770,N_12099,N_12218);
nand U14771 (N_14771,N_12203,N_12728);
and U14772 (N_14772,N_13066,N_12701);
nand U14773 (N_14773,N_13059,N_12788);
nor U14774 (N_14774,N_13434,N_13214);
nor U14775 (N_14775,N_13081,N_13168);
nand U14776 (N_14776,N_13318,N_12470);
nand U14777 (N_14777,N_13386,N_12860);
and U14778 (N_14778,N_12860,N_12412);
nor U14779 (N_14779,N_13370,N_13150);
nand U14780 (N_14780,N_12090,N_13292);
or U14781 (N_14781,N_13191,N_12380);
xor U14782 (N_14782,N_13274,N_12628);
and U14783 (N_14783,N_12659,N_13377);
and U14784 (N_14784,N_12027,N_12092);
xnor U14785 (N_14785,N_13358,N_12455);
nor U14786 (N_14786,N_12460,N_13181);
xnor U14787 (N_14787,N_12794,N_13489);
nand U14788 (N_14788,N_13225,N_13457);
or U14789 (N_14789,N_12724,N_13261);
nor U14790 (N_14790,N_13252,N_12343);
nor U14791 (N_14791,N_13356,N_12440);
xor U14792 (N_14792,N_13004,N_12860);
nor U14793 (N_14793,N_12425,N_13064);
nor U14794 (N_14794,N_12824,N_12861);
and U14795 (N_14795,N_12400,N_13376);
and U14796 (N_14796,N_12627,N_12545);
and U14797 (N_14797,N_12690,N_12296);
nor U14798 (N_14798,N_13307,N_12435);
nor U14799 (N_14799,N_12064,N_12613);
or U14800 (N_14800,N_12937,N_12461);
nor U14801 (N_14801,N_12943,N_13241);
xor U14802 (N_14802,N_12983,N_12811);
xor U14803 (N_14803,N_12226,N_13153);
and U14804 (N_14804,N_13406,N_12089);
xor U14805 (N_14805,N_12229,N_12558);
xnor U14806 (N_14806,N_13385,N_12402);
xor U14807 (N_14807,N_13216,N_13298);
nand U14808 (N_14808,N_13495,N_13152);
or U14809 (N_14809,N_13271,N_12775);
nor U14810 (N_14810,N_12341,N_13326);
nand U14811 (N_14811,N_13456,N_12492);
nor U14812 (N_14812,N_12911,N_13239);
nand U14813 (N_14813,N_12470,N_12508);
and U14814 (N_14814,N_12077,N_12933);
nor U14815 (N_14815,N_13413,N_12067);
and U14816 (N_14816,N_12098,N_12030);
xnor U14817 (N_14817,N_12710,N_12228);
nor U14818 (N_14818,N_13035,N_12829);
xor U14819 (N_14819,N_12460,N_13170);
nor U14820 (N_14820,N_12128,N_12946);
nor U14821 (N_14821,N_12124,N_12049);
and U14822 (N_14822,N_13329,N_12618);
nand U14823 (N_14823,N_12407,N_12125);
or U14824 (N_14824,N_12693,N_13033);
or U14825 (N_14825,N_12056,N_12112);
xnor U14826 (N_14826,N_12946,N_12563);
nand U14827 (N_14827,N_13339,N_12680);
or U14828 (N_14828,N_12230,N_13008);
or U14829 (N_14829,N_13326,N_12888);
nor U14830 (N_14830,N_12447,N_12729);
nand U14831 (N_14831,N_12043,N_12126);
or U14832 (N_14832,N_12620,N_13307);
xor U14833 (N_14833,N_12715,N_12450);
xor U14834 (N_14834,N_12465,N_12627);
and U14835 (N_14835,N_12667,N_12147);
nand U14836 (N_14836,N_13362,N_13266);
xor U14837 (N_14837,N_12927,N_13474);
or U14838 (N_14838,N_12245,N_13430);
and U14839 (N_14839,N_12211,N_12123);
xnor U14840 (N_14840,N_13037,N_12309);
and U14841 (N_14841,N_12191,N_13320);
xor U14842 (N_14842,N_12356,N_12658);
nand U14843 (N_14843,N_13001,N_12212);
nor U14844 (N_14844,N_12533,N_12716);
xor U14845 (N_14845,N_12596,N_13084);
xor U14846 (N_14846,N_13391,N_12176);
xor U14847 (N_14847,N_13476,N_12420);
and U14848 (N_14848,N_13241,N_12053);
or U14849 (N_14849,N_13492,N_12259);
nand U14850 (N_14850,N_12737,N_12576);
or U14851 (N_14851,N_13073,N_13320);
nand U14852 (N_14852,N_13326,N_13354);
nand U14853 (N_14853,N_12927,N_13333);
nand U14854 (N_14854,N_12172,N_12680);
xor U14855 (N_14855,N_12445,N_12723);
nand U14856 (N_14856,N_12269,N_12093);
and U14857 (N_14857,N_12518,N_12044);
and U14858 (N_14858,N_13414,N_13204);
nor U14859 (N_14859,N_12675,N_12833);
or U14860 (N_14860,N_12684,N_13398);
xor U14861 (N_14861,N_12255,N_12257);
nand U14862 (N_14862,N_12537,N_13247);
and U14863 (N_14863,N_12512,N_12933);
or U14864 (N_14864,N_12028,N_12351);
or U14865 (N_14865,N_12624,N_12797);
nor U14866 (N_14866,N_12086,N_13248);
xor U14867 (N_14867,N_13212,N_12096);
nand U14868 (N_14868,N_13376,N_13222);
nor U14869 (N_14869,N_12129,N_12720);
nand U14870 (N_14870,N_12079,N_12103);
or U14871 (N_14871,N_13490,N_12012);
nor U14872 (N_14872,N_12420,N_12957);
nand U14873 (N_14873,N_12423,N_13284);
nand U14874 (N_14874,N_12037,N_13273);
and U14875 (N_14875,N_13024,N_12456);
nor U14876 (N_14876,N_13026,N_13447);
nand U14877 (N_14877,N_12221,N_12030);
and U14878 (N_14878,N_12533,N_13114);
xnor U14879 (N_14879,N_12932,N_12343);
nor U14880 (N_14880,N_13232,N_12588);
nor U14881 (N_14881,N_12803,N_12924);
or U14882 (N_14882,N_12088,N_12179);
or U14883 (N_14883,N_13115,N_12437);
or U14884 (N_14884,N_12522,N_12000);
nand U14885 (N_14885,N_12919,N_13000);
and U14886 (N_14886,N_12514,N_12572);
nor U14887 (N_14887,N_12100,N_12838);
xnor U14888 (N_14888,N_13447,N_12175);
and U14889 (N_14889,N_12616,N_12212);
and U14890 (N_14890,N_13421,N_12385);
nor U14891 (N_14891,N_13228,N_12030);
and U14892 (N_14892,N_12396,N_12364);
nand U14893 (N_14893,N_12375,N_12786);
and U14894 (N_14894,N_12135,N_12531);
or U14895 (N_14895,N_12894,N_12285);
nor U14896 (N_14896,N_13434,N_13304);
nand U14897 (N_14897,N_13157,N_12263);
xnor U14898 (N_14898,N_12601,N_12642);
nor U14899 (N_14899,N_12544,N_13293);
nand U14900 (N_14900,N_13149,N_12117);
or U14901 (N_14901,N_12867,N_12165);
or U14902 (N_14902,N_12133,N_13337);
nand U14903 (N_14903,N_12826,N_12723);
or U14904 (N_14904,N_12856,N_12545);
xnor U14905 (N_14905,N_12854,N_12030);
nand U14906 (N_14906,N_12400,N_13107);
nor U14907 (N_14907,N_12712,N_13391);
xor U14908 (N_14908,N_13390,N_13010);
xnor U14909 (N_14909,N_12518,N_13096);
nand U14910 (N_14910,N_12446,N_12328);
or U14911 (N_14911,N_12087,N_12791);
nor U14912 (N_14912,N_12266,N_12639);
and U14913 (N_14913,N_12632,N_12500);
nand U14914 (N_14914,N_12363,N_12570);
xor U14915 (N_14915,N_12131,N_12164);
or U14916 (N_14916,N_12076,N_12972);
or U14917 (N_14917,N_12399,N_12960);
xnor U14918 (N_14918,N_13344,N_12509);
and U14919 (N_14919,N_13221,N_12229);
or U14920 (N_14920,N_13176,N_12609);
xnor U14921 (N_14921,N_13156,N_12166);
nand U14922 (N_14922,N_12698,N_12868);
nor U14923 (N_14923,N_12516,N_12721);
nor U14924 (N_14924,N_12211,N_13452);
xor U14925 (N_14925,N_13052,N_12585);
and U14926 (N_14926,N_12424,N_12666);
or U14927 (N_14927,N_12776,N_12227);
nor U14928 (N_14928,N_13349,N_12435);
nor U14929 (N_14929,N_12524,N_12202);
nor U14930 (N_14930,N_13317,N_12904);
or U14931 (N_14931,N_12205,N_12199);
xnor U14932 (N_14932,N_12003,N_13477);
nor U14933 (N_14933,N_12352,N_13365);
or U14934 (N_14934,N_12830,N_12024);
nand U14935 (N_14935,N_12199,N_13360);
xor U14936 (N_14936,N_12522,N_12902);
nand U14937 (N_14937,N_12853,N_13416);
xor U14938 (N_14938,N_12956,N_12356);
xnor U14939 (N_14939,N_12685,N_13492);
and U14940 (N_14940,N_12582,N_12747);
and U14941 (N_14941,N_13042,N_12673);
xor U14942 (N_14942,N_13110,N_13253);
or U14943 (N_14943,N_12417,N_13472);
or U14944 (N_14944,N_12487,N_12399);
or U14945 (N_14945,N_12734,N_12599);
nor U14946 (N_14946,N_13401,N_13312);
nor U14947 (N_14947,N_13367,N_12776);
and U14948 (N_14948,N_12327,N_13127);
xor U14949 (N_14949,N_12418,N_12489);
nor U14950 (N_14950,N_13302,N_13183);
and U14951 (N_14951,N_12697,N_13263);
nor U14952 (N_14952,N_12901,N_13469);
or U14953 (N_14953,N_13162,N_12485);
xor U14954 (N_14954,N_12362,N_12836);
xor U14955 (N_14955,N_13294,N_12340);
or U14956 (N_14956,N_12913,N_13322);
or U14957 (N_14957,N_13377,N_12867);
xnor U14958 (N_14958,N_13490,N_12961);
or U14959 (N_14959,N_12944,N_13471);
nor U14960 (N_14960,N_13016,N_12153);
nor U14961 (N_14961,N_12810,N_12997);
or U14962 (N_14962,N_12636,N_12610);
and U14963 (N_14963,N_13366,N_13077);
or U14964 (N_14964,N_13077,N_12519);
nor U14965 (N_14965,N_12872,N_13323);
or U14966 (N_14966,N_13027,N_12883);
or U14967 (N_14967,N_12090,N_13176);
xnor U14968 (N_14968,N_12724,N_12770);
or U14969 (N_14969,N_13379,N_12940);
nand U14970 (N_14970,N_12654,N_13154);
or U14971 (N_14971,N_13048,N_12541);
or U14972 (N_14972,N_12849,N_13156);
nor U14973 (N_14973,N_12129,N_13360);
and U14974 (N_14974,N_12116,N_12395);
or U14975 (N_14975,N_12091,N_12790);
or U14976 (N_14976,N_12435,N_12362);
nor U14977 (N_14977,N_12870,N_12791);
xor U14978 (N_14978,N_13156,N_13112);
or U14979 (N_14979,N_13370,N_12644);
and U14980 (N_14980,N_12547,N_12849);
xor U14981 (N_14981,N_12822,N_12902);
and U14982 (N_14982,N_12834,N_13469);
and U14983 (N_14983,N_13096,N_12856);
xor U14984 (N_14984,N_12809,N_12370);
xnor U14985 (N_14985,N_12438,N_12145);
or U14986 (N_14986,N_12251,N_12952);
nand U14987 (N_14987,N_13397,N_12142);
nand U14988 (N_14988,N_12033,N_12660);
or U14989 (N_14989,N_12623,N_12517);
xor U14990 (N_14990,N_12016,N_12364);
nor U14991 (N_14991,N_12735,N_12671);
and U14992 (N_14992,N_12165,N_12536);
and U14993 (N_14993,N_13056,N_12873);
nor U14994 (N_14994,N_12910,N_12676);
nand U14995 (N_14995,N_13164,N_12533);
and U14996 (N_14996,N_13325,N_12596);
and U14997 (N_14997,N_13196,N_12867);
and U14998 (N_14998,N_12518,N_12241);
and U14999 (N_14999,N_12974,N_12512);
xor U15000 (N_15000,N_14287,N_13788);
and U15001 (N_15001,N_14518,N_13791);
nor U15002 (N_15002,N_14559,N_14045);
nand U15003 (N_15003,N_14561,N_13785);
nand U15004 (N_15004,N_14314,N_14322);
and U15005 (N_15005,N_13674,N_14244);
and U15006 (N_15006,N_14610,N_14732);
nor U15007 (N_15007,N_14250,N_13618);
xnor U15008 (N_15008,N_13699,N_13852);
and U15009 (N_15009,N_13625,N_13804);
nor U15010 (N_15010,N_13610,N_14246);
and U15011 (N_15011,N_13916,N_13657);
nor U15012 (N_15012,N_14071,N_14697);
or U15013 (N_15013,N_14640,N_14899);
xnor U15014 (N_15014,N_13752,N_14480);
and U15015 (N_15015,N_14613,N_13824);
or U15016 (N_15016,N_14509,N_14624);
and U15017 (N_15017,N_13567,N_14029);
nor U15018 (N_15018,N_14046,N_13570);
nand U15019 (N_15019,N_13997,N_13524);
xor U15020 (N_15020,N_13856,N_14028);
nand U15021 (N_15021,N_14762,N_14243);
nor U15022 (N_15022,N_13993,N_14931);
or U15023 (N_15023,N_13793,N_14930);
nor U15024 (N_15024,N_14196,N_14069);
nand U15025 (N_15025,N_14924,N_14748);
nor U15026 (N_15026,N_13628,N_13575);
xnor U15027 (N_15027,N_14147,N_14240);
nand U15028 (N_15028,N_13733,N_14964);
xnor U15029 (N_15029,N_14116,N_14160);
or U15030 (N_15030,N_14227,N_14721);
nand U15031 (N_15031,N_14991,N_14706);
xor U15032 (N_15032,N_14836,N_14918);
xor U15033 (N_15033,N_13779,N_14600);
or U15034 (N_15034,N_14718,N_14499);
or U15035 (N_15035,N_14114,N_14139);
and U15036 (N_15036,N_14895,N_14236);
and U15037 (N_15037,N_13763,N_14332);
xnor U15038 (N_15038,N_14126,N_13967);
or U15039 (N_15039,N_14966,N_13879);
nand U15040 (N_15040,N_14752,N_14411);
or U15041 (N_15041,N_13745,N_14214);
nor U15042 (N_15042,N_14472,N_13556);
nor U15043 (N_15043,N_14969,N_14271);
nand U15044 (N_15044,N_13663,N_13825);
nand U15045 (N_15045,N_13500,N_14002);
nor U15046 (N_15046,N_14475,N_14885);
xnor U15047 (N_15047,N_14565,N_14186);
or U15048 (N_15048,N_13917,N_13941);
nor U15049 (N_15049,N_14595,N_14377);
xnor U15050 (N_15050,N_14496,N_14837);
or U15051 (N_15051,N_14735,N_14450);
or U15052 (N_15052,N_14337,N_14746);
nor U15053 (N_15053,N_13768,N_13517);
nand U15054 (N_15054,N_14426,N_14357);
nor U15055 (N_15055,N_13778,N_14481);
nand U15056 (N_15056,N_14960,N_13980);
xor U15057 (N_15057,N_14184,N_14479);
and U15058 (N_15058,N_13645,N_14675);
and U15059 (N_15059,N_13678,N_13960);
and U15060 (N_15060,N_14761,N_13837);
xor U15061 (N_15061,N_14488,N_14188);
or U15062 (N_15062,N_14394,N_13787);
nand U15063 (N_15063,N_14474,N_14424);
xnor U15064 (N_15064,N_13953,N_13565);
xor U15065 (N_15065,N_13704,N_14004);
xnor U15066 (N_15066,N_13693,N_13713);
nor U15067 (N_15067,N_13795,N_13849);
xor U15068 (N_15068,N_14347,N_14290);
xnor U15069 (N_15069,N_14674,N_14129);
nor U15070 (N_15070,N_14744,N_13668);
or U15071 (N_15071,N_13571,N_14767);
or U15072 (N_15072,N_13650,N_14597);
or U15073 (N_15073,N_13594,N_13597);
and U15074 (N_15074,N_14128,N_13999);
nand U15075 (N_15075,N_14050,N_14660);
and U15076 (N_15076,N_14758,N_14995);
or U15077 (N_15077,N_14514,N_14389);
or U15078 (N_15078,N_14604,N_14493);
or U15079 (N_15079,N_13922,N_14201);
or U15080 (N_15080,N_14099,N_14221);
xor U15081 (N_15081,N_14096,N_13614);
or U15082 (N_15082,N_13990,N_14666);
and U15083 (N_15083,N_13928,N_14992);
nor U15084 (N_15084,N_14469,N_14652);
and U15085 (N_15085,N_14868,N_14256);
or U15086 (N_15086,N_14832,N_14462);
nand U15087 (N_15087,N_14405,N_13735);
and U15088 (N_15088,N_13782,N_14522);
xor U15089 (N_15089,N_14408,N_14520);
or U15090 (N_15090,N_13796,N_13858);
and U15091 (N_15091,N_14968,N_14294);
and U15092 (N_15092,N_14367,N_14344);
and U15093 (N_15093,N_13672,N_14861);
and U15094 (N_15094,N_13835,N_14775);
nand U15095 (N_15095,N_13660,N_14686);
nor U15096 (N_15096,N_13540,N_14125);
xor U15097 (N_15097,N_14026,N_13739);
nor U15098 (N_15098,N_14235,N_13840);
xor U15099 (N_15099,N_14451,N_13995);
or U15100 (N_15100,N_13921,N_14699);
or U15101 (N_15101,N_14193,N_14648);
nand U15102 (N_15102,N_14694,N_14875);
and U15103 (N_15103,N_13585,N_14629);
nand U15104 (N_15104,N_14315,N_14517);
nand U15105 (N_15105,N_14502,N_13714);
nor U15106 (N_15106,N_13780,N_13648);
xor U15107 (N_15107,N_14714,N_13562);
xnor U15108 (N_15108,N_13985,N_14533);
nor U15109 (N_15109,N_14289,N_14807);
xor U15110 (N_15110,N_13655,N_13792);
xor U15111 (N_15111,N_14503,N_14633);
nand U15112 (N_15112,N_13683,N_13894);
xnor U15113 (N_15113,N_13805,N_14811);
nand U15114 (N_15114,N_14871,N_13698);
nand U15115 (N_15115,N_14788,N_13584);
nor U15116 (N_15116,N_13537,N_14231);
xnor U15117 (N_15117,N_14635,N_14866);
nor U15118 (N_15118,N_13551,N_14204);
and U15119 (N_15119,N_13630,N_14141);
and U15120 (N_15120,N_14239,N_13865);
nor U15121 (N_15121,N_14453,N_14818);
nor U15122 (N_15122,N_14159,N_14265);
or U15123 (N_15123,N_14252,N_14262);
nor U15124 (N_15124,N_14275,N_14030);
xor U15125 (N_15125,N_14829,N_14420);
and U15126 (N_15126,N_14023,N_13632);
or U15127 (N_15127,N_14833,N_14162);
xnor U15128 (N_15128,N_14812,N_13661);
xnor U15129 (N_15129,N_13769,N_13890);
xnor U15130 (N_15130,N_14316,N_14335);
xor U15131 (N_15131,N_13725,N_14508);
and U15132 (N_15132,N_14485,N_13509);
nor U15133 (N_15133,N_14548,N_14189);
nor U15134 (N_15134,N_14407,N_14111);
xnor U15135 (N_15135,N_13918,N_14738);
nand U15136 (N_15136,N_14015,N_14932);
nor U15137 (N_15137,N_13587,N_13838);
xnor U15138 (N_15138,N_14847,N_13842);
xnor U15139 (N_15139,N_13577,N_14530);
or U15140 (N_15140,N_14531,N_14524);
xnor U15141 (N_15141,N_14580,N_13870);
nand U15142 (N_15142,N_14067,N_14908);
nor U15143 (N_15143,N_13919,N_14368);
xnor U15144 (N_15144,N_14471,N_14181);
and U15145 (N_15145,N_14606,N_14253);
and U15146 (N_15146,N_13955,N_14786);
and U15147 (N_15147,N_13957,N_14180);
xnor U15148 (N_15148,N_13749,N_14364);
or U15149 (N_15149,N_14005,N_13526);
nand U15150 (N_15150,N_13803,N_14276);
xnor U15151 (N_15151,N_13695,N_14435);
xor U15152 (N_15152,N_14140,N_14327);
nand U15153 (N_15153,N_13816,N_14563);
nand U15154 (N_15154,N_14100,N_14989);
or U15155 (N_15155,N_14720,N_13641);
xor U15156 (N_15156,N_14379,N_14219);
and U15157 (N_15157,N_13887,N_13836);
nor U15158 (N_15158,N_14813,N_14704);
nor U15159 (N_15159,N_14190,N_14272);
or U15160 (N_15160,N_14835,N_13984);
xnor U15161 (N_15161,N_14443,N_14766);
nand U15162 (N_15162,N_13864,N_14881);
xnor U15163 (N_15163,N_14320,N_14319);
or U15164 (N_15164,N_13964,N_14362);
xor U15165 (N_15165,N_14318,N_13621);
or U15166 (N_15166,N_14733,N_14896);
nand U15167 (N_15167,N_14799,N_14178);
nor U15168 (N_15168,N_14627,N_14370);
xnor U15169 (N_15169,N_13924,N_14566);
nor U15170 (N_15170,N_14959,N_14304);
nand U15171 (N_15171,N_14378,N_14343);
nor U15172 (N_15172,N_14061,N_13869);
nor U15173 (N_15173,N_14073,N_14088);
nand U15174 (N_15174,N_14809,N_13817);
xor U15175 (N_15175,N_14878,N_13596);
or U15176 (N_15176,N_14537,N_14556);
nor U15177 (N_15177,N_14406,N_13506);
nand U15178 (N_15178,N_14151,N_14954);
and U15179 (N_15179,N_14935,N_13776);
xor U15180 (N_15180,N_14890,N_14158);
nand U15181 (N_15181,N_14948,N_13667);
and U15182 (N_15182,N_14618,N_13937);
nor U15183 (N_15183,N_14007,N_13538);
xor U15184 (N_15184,N_13975,N_14080);
and U15185 (N_15185,N_13572,N_14927);
nand U15186 (N_15186,N_14584,N_14428);
or U15187 (N_15187,N_14630,N_13520);
or U15188 (N_15188,N_13766,N_14296);
nand U15189 (N_15189,N_13830,N_14552);
nor U15190 (N_15190,N_14467,N_14209);
xnor U15191 (N_15191,N_14905,N_13692);
xnor U15192 (N_15192,N_13811,N_13653);
and U15193 (N_15193,N_14555,N_14619);
or U15194 (N_15194,N_14662,N_14280);
xor U15195 (N_15195,N_14911,N_13612);
xor U15196 (N_15196,N_13911,N_13880);
xor U15197 (N_15197,N_13573,N_13731);
nor U15198 (N_15198,N_14498,N_14313);
or U15199 (N_15199,N_13883,N_13989);
or U15200 (N_15200,N_13715,N_14115);
xor U15201 (N_15201,N_14550,N_14000);
and U15202 (N_15202,N_13862,N_13754);
xnor U15203 (N_15203,N_14081,N_13746);
and U15204 (N_15204,N_14113,N_14669);
nor U15205 (N_15205,N_14928,N_14416);
nand U15206 (N_15206,N_13772,N_14354);
or U15207 (N_15207,N_14609,N_14737);
or U15208 (N_15208,N_13607,N_14459);
nand U15209 (N_15209,N_14210,N_13501);
xnor U15210 (N_15210,N_13868,N_13821);
and U15211 (N_15211,N_13589,N_14120);
or U15212 (N_15212,N_14505,N_13945);
and U15213 (N_15213,N_14458,N_14392);
or U15214 (N_15214,N_13898,N_14779);
or U15215 (N_15215,N_13765,N_14103);
nand U15216 (N_15216,N_13590,N_14900);
nand U15217 (N_15217,N_14292,N_13720);
or U15218 (N_15218,N_14990,N_14104);
or U15219 (N_15219,N_14303,N_13963);
nand U15220 (N_15220,N_14056,N_14751);
or U15221 (N_15221,N_14404,N_14047);
nand U15222 (N_15222,N_14078,N_14547);
xnor U15223 (N_15223,N_13734,N_14838);
nor U15224 (N_15224,N_14218,N_14685);
nor U15225 (N_15225,N_14489,N_14351);
and U15226 (N_15226,N_13664,N_13969);
nor U15227 (N_15227,N_13992,N_14288);
or U15228 (N_15228,N_13541,N_14864);
nor U15229 (N_15229,N_13806,N_14631);
nand U15230 (N_15230,N_13554,N_14677);
nand U15231 (N_15231,N_13759,N_14082);
xnor U15232 (N_15232,N_14187,N_14171);
xor U15233 (N_15233,N_14820,N_14170);
xnor U15234 (N_15234,N_13708,N_14795);
or U15235 (N_15235,N_13581,N_13951);
and U15236 (N_15236,N_14445,N_14632);
or U15237 (N_15237,N_14042,N_14637);
nand U15238 (N_15238,N_13876,N_14083);
nand U15239 (N_15239,N_14041,N_13936);
nor U15240 (N_15240,N_13929,N_14696);
xnor U15241 (N_15241,N_13710,N_14274);
xor U15242 (N_15242,N_14340,N_14817);
and U15243 (N_15243,N_13934,N_14345);
or U15244 (N_15244,N_14841,N_14473);
xor U15245 (N_15245,N_13751,N_14869);
and U15246 (N_15246,N_13712,N_14477);
and U15247 (N_15247,N_14585,N_14084);
nand U15248 (N_15248,N_14433,N_14242);
or U15249 (N_15249,N_14490,N_13557);
or U15250 (N_15250,N_13948,N_14019);
nand U15251 (N_15251,N_14179,N_14157);
and U15252 (N_15252,N_14329,N_13600);
nor U15253 (N_15253,N_14495,N_14800);
nand U15254 (N_15254,N_14057,N_14998);
or U15255 (N_15255,N_14543,N_13956);
xor U15256 (N_15256,N_14665,N_14386);
or U15257 (N_15257,N_14776,N_13603);
and U15258 (N_15258,N_13716,N_14554);
and U15259 (N_15259,N_14693,N_13671);
nand U15260 (N_15260,N_14785,N_14897);
and U15261 (N_15261,N_14300,N_13949);
nor U15262 (N_15262,N_14399,N_14577);
and U15263 (N_15263,N_14237,N_13820);
xor U15264 (N_15264,N_14700,N_13622);
nor U15265 (N_15265,N_14167,N_14311);
or U15266 (N_15266,N_13691,N_14657);
nor U15267 (N_15267,N_13823,N_13923);
and U15268 (N_15268,N_13659,N_14754);
xnor U15269 (N_15269,N_13748,N_14952);
and U15270 (N_15270,N_14447,N_13848);
nor U15271 (N_15271,N_14176,N_13552);
nand U15272 (N_15272,N_14064,N_14971);
or U15273 (N_15273,N_14174,N_14484);
xnor U15274 (N_15274,N_13818,N_14951);
nand U15275 (N_15275,N_14876,N_14544);
nand U15276 (N_15276,N_14153,N_14409);
nor U15277 (N_15277,N_13521,N_13617);
nand U15278 (N_15278,N_14279,N_14769);
nand U15279 (N_15279,N_14233,N_14202);
nor U15280 (N_15280,N_14622,N_14593);
and U15281 (N_15281,N_14594,N_14743);
xor U15282 (N_15282,N_14270,N_13750);
nor U15283 (N_15283,N_14805,N_13885);
or U15284 (N_15284,N_13874,N_13943);
xor U15285 (N_15285,N_14771,N_13684);
or U15286 (N_15286,N_13592,N_13611);
nor U15287 (N_15287,N_13901,N_13703);
or U15288 (N_15288,N_14097,N_14512);
or U15289 (N_15289,N_14446,N_13665);
and U15290 (N_15290,N_14623,N_14355);
and U15291 (N_15291,N_13938,N_13799);
and U15292 (N_15292,N_13599,N_13906);
and U15293 (N_15293,N_14123,N_14826);
and U15294 (N_15294,N_13832,N_14273);
xnor U15295 (N_15295,N_13784,N_13737);
and U15296 (N_15296,N_14612,N_13889);
xnor U15297 (N_15297,N_14172,N_14258);
nand U15298 (N_15298,N_14439,N_14915);
xnor U15299 (N_15299,N_13639,N_14557);
nand U15300 (N_15300,N_13853,N_14043);
or U15301 (N_15301,N_13504,N_14259);
xnor U15302 (N_15302,N_14014,N_14843);
or U15303 (N_15303,N_14325,N_14284);
and U15304 (N_15304,N_14092,N_14570);
nand U15305 (N_15305,N_14155,N_14143);
nand U15306 (N_15306,N_14317,N_14079);
and U15307 (N_15307,N_14821,N_13624);
or U15308 (N_15308,N_14033,N_13602);
nor U15309 (N_15309,N_14963,N_13550);
and U15310 (N_15310,N_14756,N_13535);
nand U15311 (N_15311,N_14255,N_14944);
or U15312 (N_15312,N_14538,N_13814);
and U15313 (N_15313,N_14797,N_14299);
or U15314 (N_15314,N_14049,N_13656);
and U15315 (N_15315,N_14412,N_14650);
nor U15316 (N_15316,N_13912,N_13544);
nor U15317 (N_15317,N_14150,N_14938);
xor U15318 (N_15318,N_14987,N_14796);
and U15319 (N_15319,N_14022,N_14937);
nand U15320 (N_15320,N_14972,N_14268);
nor U15321 (N_15321,N_14526,N_13828);
nor U15322 (N_15322,N_13508,N_14198);
or U15323 (N_15323,N_13512,N_13709);
xnor U15324 (N_15324,N_13635,N_14361);
or U15325 (N_15325,N_13987,N_14664);
or U15326 (N_15326,N_14719,N_13764);
nor U15327 (N_15327,N_14815,N_14961);
nor U15328 (N_15328,N_13642,N_13925);
or U15329 (N_15329,N_14238,N_14429);
and U15330 (N_15330,N_14919,N_14901);
or U15331 (N_15331,N_14909,N_14483);
and U15332 (N_15332,N_14572,N_14397);
nor U15333 (N_15333,N_13591,N_14614);
and U15334 (N_15334,N_13636,N_14427);
or U15335 (N_15335,N_14168,N_13813);
and U15336 (N_15336,N_14217,N_13702);
and U15337 (N_15337,N_14768,N_14546);
or U15338 (N_15338,N_14413,N_14814);
or U15339 (N_15339,N_14642,N_14182);
and U15340 (N_15340,N_13857,N_14551);
and U15341 (N_15341,N_14220,N_14468);
nor U15342 (N_15342,N_14295,N_14849);
xnor U15343 (N_15343,N_14525,N_13568);
nor U15344 (N_15344,N_13962,N_14857);
xor U15345 (N_15345,N_13877,N_14077);
or U15346 (N_15346,N_14855,N_14309);
xor U15347 (N_15347,N_14925,N_14777);
or U15348 (N_15348,N_13559,N_14321);
xor U15349 (N_15349,N_14926,N_13619);
nand U15350 (N_15350,N_13580,N_13904);
or U15351 (N_15351,N_14491,N_14310);
xor U15352 (N_15352,N_14349,N_14059);
nor U15353 (N_15353,N_14431,N_13644);
xnor U15354 (N_15354,N_13932,N_14791);
nor U15355 (N_15355,N_13843,N_14527);
nand U15356 (N_15356,N_14039,N_14009);
nor U15357 (N_15357,N_13950,N_14586);
xnor U15358 (N_15358,N_13847,N_14402);
and U15359 (N_15359,N_14144,N_14688);
nand U15360 (N_15360,N_14880,N_14605);
and U15361 (N_15361,N_14542,N_13786);
xnor U15362 (N_15362,N_13760,N_14553);
and U15363 (N_15363,N_14996,N_13767);
or U15364 (N_15364,N_13727,N_14156);
xnor U15365 (N_15365,N_14806,N_13991);
nand U15366 (N_15366,N_13643,N_14482);
or U15367 (N_15367,N_14740,N_13998);
and U15368 (N_15368,N_13681,N_14993);
nor U15369 (N_15369,N_14945,N_13629);
or U15370 (N_15370,N_14173,N_14245);
and U15371 (N_15371,N_14701,N_14840);
nand U15372 (N_15372,N_13971,N_14611);
xor U15373 (N_15373,N_14912,N_14017);
nand U15374 (N_15374,N_13696,N_14691);
or U15375 (N_15375,N_13502,N_13598);
and U15376 (N_15376,N_14454,N_14979);
nor U15377 (N_15377,N_14576,N_14305);
nor U15378 (N_15378,N_13680,N_14645);
and U15379 (N_15379,N_14234,N_14974);
nand U15380 (N_15380,N_14037,N_14138);
nor U15381 (N_15381,N_14667,N_14455);
nand U15382 (N_15382,N_14105,N_14387);
xnor U15383 (N_15383,N_14943,N_14656);
xnor U15384 (N_15384,N_13705,N_14093);
nand U15385 (N_15385,N_14985,N_14910);
xnor U15386 (N_15386,N_14904,N_14348);
or U15387 (N_15387,N_13790,N_14425);
and U15388 (N_15388,N_13891,N_14216);
nor U15389 (N_15389,N_14634,N_14363);
xnor U15390 (N_15390,N_13846,N_14649);
nand U15391 (N_15391,N_13913,N_14860);
xnor U15392 (N_15392,N_13819,N_13812);
xnor U15393 (N_15393,N_13810,N_14906);
and U15394 (N_15394,N_14916,N_14515);
xor U15395 (N_15395,N_14163,N_14124);
xnor U15396 (N_15396,N_14452,N_14154);
nor U15397 (N_15397,N_13841,N_14842);
nand U15398 (N_15398,N_14934,N_13976);
and U15399 (N_15399,N_14641,N_14755);
nor U15400 (N_15400,N_13944,N_14127);
nor U15401 (N_15401,N_13634,N_14072);
and U15402 (N_15402,N_14671,N_14651);
and U15403 (N_15403,N_14090,N_14819);
xor U15404 (N_15404,N_13519,N_14867);
and U15405 (N_15405,N_14194,N_14984);
or U15406 (N_15406,N_13626,N_13722);
or U15407 (N_15407,N_14856,N_14263);
nor U15408 (N_15408,N_14780,N_13531);
nand U15409 (N_15409,N_14678,N_14845);
nor U15410 (N_15410,N_14063,N_14307);
or U15411 (N_15411,N_14205,N_13873);
xor U15412 (N_15412,N_14089,N_14760);
nand U15413 (N_15413,N_14921,N_14646);
and U15414 (N_15414,N_14432,N_13882);
xor U15415 (N_15415,N_14494,N_14626);
nor U15416 (N_15416,N_14036,N_13578);
or U15417 (N_15417,N_13515,N_14027);
or U15418 (N_15418,N_14197,N_13546);
or U15419 (N_15419,N_13884,N_13706);
nand U15420 (N_15420,N_14684,N_13606);
and U15421 (N_15421,N_14278,N_13972);
nand U15422 (N_15422,N_13893,N_14852);
and U15423 (N_15423,N_14528,N_14628);
xnor U15424 (N_15424,N_13724,N_14747);
xor U15425 (N_15425,N_13637,N_14638);
nor U15426 (N_15426,N_13942,N_14010);
or U15427 (N_15427,N_14261,N_14942);
or U15428 (N_15428,N_14464,N_14687);
nand U15429 (N_15429,N_14923,N_13669);
or U15430 (N_15430,N_14887,N_14893);
or U15431 (N_15431,N_14682,N_14228);
nand U15432 (N_15432,N_14415,N_14013);
or U15433 (N_15433,N_14511,N_14581);
nor U15434 (N_15434,N_14802,N_14888);
nor U15435 (N_15435,N_13586,N_14247);
nand U15436 (N_15436,N_14146,N_14224);
or U15437 (N_15437,N_13569,N_14598);
nor U15438 (N_15438,N_14574,N_13730);
or U15439 (N_15439,N_13761,N_13888);
nor U15440 (N_15440,N_14331,N_14286);
nor U15441 (N_15441,N_14192,N_13595);
nand U15442 (N_15442,N_13822,N_14907);
nand U15443 (N_15443,N_14940,N_14728);
and U15444 (N_15444,N_14913,N_13940);
and U15445 (N_15445,N_14883,N_14195);
and U15446 (N_15446,N_13958,N_14715);
nor U15447 (N_15447,N_14858,N_14132);
nand U15448 (N_15448,N_14830,N_14264);
nor U15449 (N_15449,N_14568,N_13583);
nand U15450 (N_15450,N_14044,N_13563);
and U15451 (N_15451,N_13973,N_14025);
nand U15452 (N_15452,N_13886,N_14066);
nor U15453 (N_15453,N_14827,N_14729);
xor U15454 (N_15454,N_14388,N_14975);
or U15455 (N_15455,N_14573,N_14133);
xnor U15456 (N_15456,N_14532,N_14350);
nand U15457 (N_15457,N_14516,N_13627);
nand U15458 (N_15458,N_13994,N_14659);
xnor U15459 (N_15459,N_13827,N_14169);
nor U15460 (N_15460,N_13528,N_14380);
xor U15461 (N_15461,N_14596,N_13833);
and U15462 (N_15462,N_14251,N_13881);
and U15463 (N_15463,N_14884,N_14644);
xor U15464 (N_15464,N_14006,N_14395);
xor U15465 (N_15465,N_14101,N_13866);
or U15466 (N_15466,N_14958,N_14541);
or U15467 (N_15467,N_13553,N_14792);
xnor U15468 (N_15468,N_14591,N_14373);
nand U15469 (N_15469,N_13755,N_14465);
nand U15470 (N_15470,N_13861,N_14726);
xor U15471 (N_15471,N_14962,N_14297);
or U15472 (N_15472,N_13651,N_13687);
or U15473 (N_15473,N_13566,N_14862);
and U15474 (N_15474,N_14602,N_14834);
and U15475 (N_15475,N_14385,N_14643);
xnor U15476 (N_15476,N_14757,N_14293);
xnor U15477 (N_15477,N_14021,N_13959);
and U15478 (N_15478,N_14965,N_14248);
xor U15479 (N_15479,N_13996,N_14727);
xor U15480 (N_15480,N_13899,N_13723);
xnor U15481 (N_15481,N_13939,N_14803);
and U15482 (N_15482,N_14941,N_13673);
or U15483 (N_15483,N_14801,N_14707);
nor U15484 (N_15484,N_13927,N_13662);
or U15485 (N_15485,N_13815,N_13777);
nand U15486 (N_15486,N_13707,N_13633);
xor U15487 (N_15487,N_14933,N_14381);
nand U15488 (N_15488,N_14967,N_14997);
xnor U15489 (N_15489,N_14177,N_14571);
xnor U15490 (N_15490,N_14417,N_13522);
nand U15491 (N_15491,N_14708,N_14122);
or U15492 (N_15492,N_14476,N_14478);
or U15493 (N_15493,N_14460,N_14575);
nor U15494 (N_15494,N_13623,N_14110);
and U15495 (N_15495,N_14793,N_14410);
nand U15496 (N_15496,N_14668,N_13523);
or U15497 (N_15497,N_14312,N_14789);
or U15498 (N_15498,N_14564,N_14254);
and U15499 (N_15499,N_13775,N_14301);
xnor U15500 (N_15500,N_14698,N_13798);
and U15501 (N_15501,N_13679,N_14980);
and U15502 (N_15502,N_13564,N_13530);
or U15503 (N_15503,N_14074,N_14535);
or U15504 (N_15504,N_14655,N_14382);
or U15505 (N_15505,N_13601,N_14003);
nand U15506 (N_15506,N_14782,N_14200);
xnor U15507 (N_15507,N_13542,N_14653);
and U15508 (N_15508,N_14983,N_14712);
nand U15509 (N_15509,N_13677,N_13896);
and U15510 (N_15510,N_14257,N_14438);
and U15511 (N_15511,N_14504,N_14592);
or U15512 (N_15512,N_14745,N_14232);
xor U15513 (N_15513,N_14730,N_14589);
and U15514 (N_15514,N_13690,N_14011);
xnor U15515 (N_15515,N_14703,N_14298);
or U15516 (N_15516,N_14306,N_13738);
nand U15517 (N_15517,N_14185,N_14142);
xor U15518 (N_15518,N_14055,N_14810);
nand U15519 (N_15519,N_14567,N_14356);
nor U15520 (N_15520,N_14903,N_14330);
xor U15521 (N_15521,N_14366,N_14590);
or U15522 (N_15522,N_13910,N_14136);
nor U15523 (N_15523,N_14978,N_13802);
xor U15524 (N_15524,N_13860,N_13507);
and U15525 (N_15525,N_14889,N_13859);
nor U15526 (N_15526,N_14823,N_14442);
or U15527 (N_15527,N_14487,N_14342);
or U15528 (N_15528,N_14731,N_14095);
nor U15529 (N_15529,N_13549,N_14636);
or U15530 (N_15530,N_14323,N_14709);
nand U15531 (N_15531,N_14436,N_14051);
and U15532 (N_15532,N_14058,N_13654);
and U15533 (N_15533,N_14616,N_13961);
xnor U15534 (N_15534,N_13718,N_14421);
xnor U15535 (N_15535,N_14545,N_14781);
nand U15536 (N_15536,N_14988,N_13676);
or U15537 (N_15537,N_14839,N_14920);
xnor U15538 (N_15538,N_14440,N_13986);
nand U15539 (N_15539,N_14723,N_14661);
and U15540 (N_15540,N_14230,N_13966);
nand U15541 (N_15541,N_14763,N_13974);
nor U15542 (N_15542,N_13826,N_13988);
xor U15543 (N_15543,N_13757,N_14947);
nand U15544 (N_15544,N_13534,N_13505);
nand U15545 (N_15545,N_14500,N_13770);
and U15546 (N_15546,N_13605,N_13582);
and U15547 (N_15547,N_14949,N_14725);
xnor U15548 (N_15548,N_14336,N_14134);
xor U15549 (N_15549,N_14034,N_14396);
and U15550 (N_15550,N_14461,N_14716);
xnor U15551 (N_15551,N_14183,N_14121);
or U15552 (N_15552,N_14658,N_14119);
or U15553 (N_15553,N_14393,N_14759);
and U15554 (N_15554,N_13527,N_14444);
nand U15555 (N_15555,N_13903,N_13920);
nand U15556 (N_15556,N_14680,N_14956);
xor U15557 (N_15557,N_14076,N_14203);
and U15558 (N_15558,N_14223,N_14741);
nand U15559 (N_15559,N_13511,N_14283);
nand U15560 (N_15560,N_13732,N_13954);
or U15561 (N_15561,N_14497,N_14929);
and U15562 (N_15562,N_14222,N_14521);
xor U15563 (N_15563,N_14922,N_13915);
xor U15564 (N_15564,N_13638,N_13789);
nor U15565 (N_15565,N_14854,N_13543);
nor U15566 (N_15566,N_14578,N_13608);
or U15567 (N_15567,N_14790,N_14981);
and U15568 (N_15568,N_13532,N_13701);
and U15569 (N_15569,N_14012,N_13700);
xor U15570 (N_15570,N_14539,N_13947);
and U15571 (N_15571,N_14560,N_14341);
and U15572 (N_15572,N_13666,N_14492);
xor U15573 (N_15573,N_13900,N_14024);
xor U15574 (N_15574,N_13844,N_14976);
or U15575 (N_15575,N_14513,N_14955);
nand U15576 (N_15576,N_13574,N_14249);
nor U15577 (N_15577,N_14683,N_13834);
xor U15578 (N_15578,N_14434,N_13620);
nor U15579 (N_15579,N_13719,N_14326);
nand U15580 (N_15580,N_14957,N_14549);
xnor U15581 (N_15581,N_13548,N_13933);
nand U15582 (N_15582,N_13593,N_14062);
nand U15583 (N_15583,N_13682,N_14562);
nand U15584 (N_15584,N_14615,N_13970);
nor U15585 (N_15585,N_14621,N_14291);
nor U15586 (N_15586,N_14149,N_14001);
and U15587 (N_15587,N_13902,N_14086);
xor U15588 (N_15588,N_14376,N_14038);
nand U15589 (N_15589,N_14603,N_14828);
nand U15590 (N_15590,N_14466,N_14191);
xor U15591 (N_15591,N_14148,N_14285);
nand U15592 (N_15592,N_13740,N_14946);
or U15593 (N_15593,N_13875,N_13771);
and U15594 (N_15594,N_14774,N_14588);
or U15595 (N_15595,N_14365,N_14994);
nor U15596 (N_15596,N_14437,N_14229);
nor U15597 (N_15597,N_13747,N_14808);
xor U15598 (N_15598,N_14102,N_13863);
nand U15599 (N_15599,N_13717,N_13808);
xnor U15600 (N_15600,N_14569,N_14145);
and U15601 (N_15601,N_14999,N_13758);
xnor U15602 (N_15602,N_14783,N_14423);
or U15603 (N_15603,N_14470,N_14098);
and U15604 (N_15604,N_14844,N_14346);
or U15605 (N_15605,N_13907,N_13895);
nor U15606 (N_15606,N_14463,N_14441);
nor U15607 (N_15607,N_14371,N_13905);
nand U15608 (N_15608,N_14710,N_13604);
xnor U15609 (N_15609,N_14333,N_14787);
or U15610 (N_15610,N_14506,N_14040);
xor U15611 (N_15611,N_14798,N_14672);
or U15612 (N_15612,N_14020,N_14053);
or U15613 (N_15613,N_13831,N_13609);
nor U15614 (N_15614,N_14713,N_14383);
or U15615 (N_15615,N_14112,N_14898);
xor U15616 (N_15616,N_14717,N_13783);
xnor U15617 (N_15617,N_14874,N_14620);
and U15618 (N_15618,N_14282,N_14401);
xor U15619 (N_15619,N_14804,N_14352);
or U15620 (N_15620,N_14175,N_14068);
xnor U15621 (N_15621,N_14722,N_14052);
and U15622 (N_15622,N_14917,N_14765);
or U15623 (N_15623,N_14369,N_14772);
xor U15624 (N_15624,N_13756,N_13935);
and U15625 (N_15625,N_13850,N_14032);
and U15626 (N_15626,N_13694,N_14241);
xor U15627 (N_15627,N_13794,N_14870);
nand U15628 (N_15628,N_13839,N_14705);
or U15629 (N_15629,N_13867,N_14583);
xor U15630 (N_15630,N_14207,N_14663);
nand U15631 (N_15631,N_14166,N_13721);
nor U15632 (N_15632,N_13968,N_14384);
or U15633 (N_15633,N_14456,N_13965);
xnor U15634 (N_15634,N_14501,N_14390);
and U15635 (N_15635,N_14734,N_14165);
nand U15636 (N_15636,N_14208,N_14892);
xor U15637 (N_15637,N_14302,N_14486);
or U15638 (N_15638,N_13685,N_13982);
xor U15639 (N_15639,N_13981,N_13658);
and U15640 (N_15640,N_14939,N_13697);
nor U15641 (N_15641,N_13797,N_14048);
or U15642 (N_15642,N_14695,N_14702);
xor U15643 (N_15643,N_13525,N_14647);
nand U15644 (N_15644,N_14749,N_14773);
and U15645 (N_15645,N_14226,N_13675);
and U15646 (N_15646,N_14851,N_14085);
xnor U15647 (N_15647,N_14986,N_14225);
xnor U15648 (N_15648,N_14582,N_13631);
nor U15649 (N_15649,N_13930,N_14281);
and U15650 (N_15650,N_14886,N_13773);
nor U15651 (N_15651,N_13871,N_13613);
xor U15652 (N_15652,N_14414,N_14690);
nor U15653 (N_15653,N_14008,N_14859);
nand U15654 (N_15654,N_14711,N_13872);
nand U15655 (N_15655,N_14152,N_14070);
nand U15656 (N_15656,N_14865,N_13518);
or U15657 (N_15657,N_14135,N_13931);
nand U15658 (N_15658,N_13736,N_14936);
nor U15659 (N_15659,N_13558,N_14778);
nor U15660 (N_15660,N_14016,N_13742);
nor U15661 (N_15661,N_14853,N_14211);
or U15662 (N_15662,N_14617,N_14894);
or U15663 (N_15663,N_14891,N_14784);
and U15664 (N_15664,N_13729,N_14213);
xnor U15665 (N_15665,N_14457,N_13809);
nor U15666 (N_15666,N_13615,N_13652);
or U15667 (N_15667,N_14882,N_13800);
xor U15668 (N_15668,N_13914,N_13978);
xor U15669 (N_15669,N_13878,N_13908);
and U15670 (N_15670,N_13892,N_13983);
xor U15671 (N_15671,N_13909,N_13977);
and U15672 (N_15672,N_14212,N_14753);
xnor U15673 (N_15673,N_13547,N_14670);
or U15674 (N_15674,N_14065,N_13726);
nor U15675 (N_15675,N_14977,N_14267);
xnor U15676 (N_15676,N_14587,N_14607);
and U15677 (N_15677,N_14724,N_14794);
nor U15678 (N_15678,N_14816,N_13516);
nand U15679 (N_15679,N_14681,N_13555);
or U15680 (N_15680,N_13647,N_14161);
nand U15681 (N_15681,N_14164,N_14822);
nor U15682 (N_15682,N_14764,N_14353);
nand U15683 (N_15683,N_13539,N_14215);
nor U15684 (N_15684,N_13728,N_13744);
xnor U15685 (N_15685,N_13762,N_13851);
xnor U15686 (N_15686,N_13688,N_14540);
or U15687 (N_15687,N_14825,N_14679);
xor U15688 (N_15688,N_13503,N_14902);
xor U15689 (N_15689,N_14914,N_13536);
nand U15690 (N_15690,N_14422,N_14106);
nor U15691 (N_15691,N_14060,N_14130);
or U15692 (N_15692,N_14850,N_14872);
xnor U15693 (N_15693,N_14846,N_13646);
nor U15694 (N_15694,N_14824,N_14418);
and U15695 (N_15695,N_14529,N_14534);
or U15696 (N_15696,N_14510,N_13579);
nand U15697 (N_15697,N_13743,N_14391);
and U15698 (N_15698,N_13588,N_14973);
and U15699 (N_15699,N_14863,N_14419);
and U15700 (N_15700,N_13897,N_13774);
nand U15701 (N_15701,N_13781,N_14689);
and U15702 (N_15702,N_14770,N_14137);
nor U15703 (N_15703,N_14277,N_13855);
nor U15704 (N_15704,N_14953,N_14260);
and U15705 (N_15705,N_14739,N_13510);
and U15706 (N_15706,N_14091,N_14673);
xnor U15707 (N_15707,N_14109,N_13829);
and U15708 (N_15708,N_13560,N_14398);
xor U15709 (N_15709,N_13513,N_13807);
nor U15710 (N_15710,N_14018,N_14054);
nor U15711 (N_15711,N_14324,N_14448);
nand U15712 (N_15712,N_14848,N_14625);
xnor U15713 (N_15713,N_14692,N_14558);
nor U15714 (N_15714,N_14831,N_14269);
xnor U15715 (N_15715,N_14087,N_13576);
or U15716 (N_15716,N_14449,N_13946);
xor U15717 (N_15717,N_13711,N_13649);
nand U15718 (N_15718,N_14742,N_14736);
nand U15719 (N_15719,N_14400,N_14035);
and U15720 (N_15720,N_13854,N_14094);
nor U15721 (N_15721,N_14372,N_14266);
or U15722 (N_15722,N_14359,N_14879);
or U15723 (N_15723,N_14601,N_14334);
and U15724 (N_15724,N_14599,N_13529);
nand U15725 (N_15725,N_14131,N_14536);
nand U15726 (N_15726,N_14360,N_13545);
nor U15727 (N_15727,N_13741,N_14375);
nand U15728 (N_15728,N_14750,N_14877);
or U15729 (N_15729,N_14523,N_13979);
nor U15730 (N_15730,N_14579,N_14982);
nand U15731 (N_15731,N_14608,N_13640);
xor U15732 (N_15732,N_14118,N_14358);
nand U15733 (N_15733,N_14430,N_13801);
nor U15734 (N_15734,N_13686,N_14654);
and U15735 (N_15735,N_14374,N_14676);
nor U15736 (N_15736,N_14339,N_14970);
nor U15737 (N_15737,N_14075,N_14328);
and U15738 (N_15738,N_14507,N_13514);
and U15739 (N_15739,N_14199,N_14117);
nand U15740 (N_15740,N_13845,N_13533);
or U15741 (N_15741,N_13561,N_14950);
and U15742 (N_15742,N_14519,N_14108);
nand U15743 (N_15743,N_14206,N_14031);
nand U15744 (N_15744,N_14403,N_13689);
and U15745 (N_15745,N_14639,N_14107);
nand U15746 (N_15746,N_13670,N_14308);
xor U15747 (N_15747,N_14873,N_13952);
xnor U15748 (N_15748,N_13926,N_14338);
or U15749 (N_15749,N_13616,N_13753);
or U15750 (N_15750,N_14961,N_13894);
nor U15751 (N_15751,N_13825,N_14732);
nand U15752 (N_15752,N_13683,N_14697);
and U15753 (N_15753,N_14236,N_14797);
nand U15754 (N_15754,N_14708,N_14645);
nand U15755 (N_15755,N_14598,N_14968);
nand U15756 (N_15756,N_14854,N_13669);
nand U15757 (N_15757,N_14539,N_14780);
and U15758 (N_15758,N_13794,N_14736);
and U15759 (N_15759,N_14303,N_14511);
and U15760 (N_15760,N_14951,N_14408);
or U15761 (N_15761,N_14327,N_13653);
nand U15762 (N_15762,N_14797,N_14719);
nor U15763 (N_15763,N_13765,N_14148);
nor U15764 (N_15764,N_13651,N_14667);
or U15765 (N_15765,N_14948,N_14993);
nor U15766 (N_15766,N_14397,N_14922);
nand U15767 (N_15767,N_14585,N_14155);
xnor U15768 (N_15768,N_14087,N_14263);
xnor U15769 (N_15769,N_13762,N_14644);
nand U15770 (N_15770,N_13840,N_14984);
nand U15771 (N_15771,N_14119,N_14445);
nand U15772 (N_15772,N_13601,N_14561);
nand U15773 (N_15773,N_13678,N_14239);
nor U15774 (N_15774,N_14481,N_14544);
nor U15775 (N_15775,N_14522,N_14745);
and U15776 (N_15776,N_13879,N_14494);
and U15777 (N_15777,N_14110,N_14568);
and U15778 (N_15778,N_14680,N_13973);
or U15779 (N_15779,N_14294,N_14775);
xor U15780 (N_15780,N_14688,N_14205);
or U15781 (N_15781,N_14433,N_14248);
nand U15782 (N_15782,N_13523,N_13556);
and U15783 (N_15783,N_14618,N_13632);
xnor U15784 (N_15784,N_14943,N_14147);
or U15785 (N_15785,N_14540,N_14638);
and U15786 (N_15786,N_13796,N_14452);
xnor U15787 (N_15787,N_14588,N_13940);
or U15788 (N_15788,N_14746,N_14286);
nor U15789 (N_15789,N_14271,N_14872);
nor U15790 (N_15790,N_13690,N_14277);
and U15791 (N_15791,N_14008,N_14718);
nand U15792 (N_15792,N_13820,N_14186);
xnor U15793 (N_15793,N_13869,N_14901);
or U15794 (N_15794,N_14349,N_13715);
and U15795 (N_15795,N_14328,N_13871);
nor U15796 (N_15796,N_13575,N_14318);
xnor U15797 (N_15797,N_14232,N_14624);
and U15798 (N_15798,N_14503,N_13722);
or U15799 (N_15799,N_14941,N_13820);
and U15800 (N_15800,N_14069,N_14146);
or U15801 (N_15801,N_14237,N_14854);
nor U15802 (N_15802,N_14509,N_14690);
nand U15803 (N_15803,N_13796,N_14332);
and U15804 (N_15804,N_14465,N_14069);
nand U15805 (N_15805,N_14006,N_14781);
nand U15806 (N_15806,N_14917,N_13602);
and U15807 (N_15807,N_14381,N_13639);
nand U15808 (N_15808,N_13978,N_13863);
and U15809 (N_15809,N_13608,N_14079);
xor U15810 (N_15810,N_13652,N_13722);
and U15811 (N_15811,N_14519,N_14732);
and U15812 (N_15812,N_14704,N_14863);
and U15813 (N_15813,N_14561,N_14826);
xor U15814 (N_15814,N_14545,N_13921);
nor U15815 (N_15815,N_13528,N_14449);
xnor U15816 (N_15816,N_14754,N_14884);
nand U15817 (N_15817,N_14237,N_14232);
nor U15818 (N_15818,N_14658,N_14376);
nor U15819 (N_15819,N_14225,N_13830);
nand U15820 (N_15820,N_13601,N_13933);
xnor U15821 (N_15821,N_14706,N_14844);
xor U15822 (N_15822,N_14500,N_14201);
xnor U15823 (N_15823,N_13865,N_14593);
and U15824 (N_15824,N_13718,N_13596);
xnor U15825 (N_15825,N_14299,N_13840);
xor U15826 (N_15826,N_14149,N_13628);
nor U15827 (N_15827,N_14996,N_13823);
and U15828 (N_15828,N_14528,N_14676);
or U15829 (N_15829,N_14310,N_14299);
or U15830 (N_15830,N_13625,N_13819);
nor U15831 (N_15831,N_14632,N_14781);
nor U15832 (N_15832,N_14949,N_14497);
nor U15833 (N_15833,N_14596,N_13866);
nand U15834 (N_15834,N_14729,N_13648);
or U15835 (N_15835,N_13925,N_14896);
nor U15836 (N_15836,N_14140,N_13716);
and U15837 (N_15837,N_13938,N_14877);
nand U15838 (N_15838,N_14933,N_13838);
nor U15839 (N_15839,N_13725,N_14357);
nand U15840 (N_15840,N_14096,N_14046);
or U15841 (N_15841,N_14498,N_14416);
nand U15842 (N_15842,N_13979,N_14752);
nand U15843 (N_15843,N_14678,N_14858);
xnor U15844 (N_15844,N_13961,N_14571);
nor U15845 (N_15845,N_14374,N_14207);
and U15846 (N_15846,N_14872,N_14255);
or U15847 (N_15847,N_14619,N_14279);
xnor U15848 (N_15848,N_14258,N_13953);
or U15849 (N_15849,N_14947,N_13546);
or U15850 (N_15850,N_13731,N_14951);
xor U15851 (N_15851,N_13640,N_14217);
nor U15852 (N_15852,N_14925,N_14999);
xnor U15853 (N_15853,N_13634,N_14613);
nand U15854 (N_15854,N_14348,N_13653);
xnor U15855 (N_15855,N_14733,N_14486);
and U15856 (N_15856,N_14168,N_13978);
and U15857 (N_15857,N_14166,N_13632);
nand U15858 (N_15858,N_14157,N_14936);
or U15859 (N_15859,N_14837,N_14169);
nand U15860 (N_15860,N_14522,N_14643);
or U15861 (N_15861,N_13532,N_13631);
nor U15862 (N_15862,N_13899,N_14741);
and U15863 (N_15863,N_14687,N_13587);
xnor U15864 (N_15864,N_13880,N_14324);
nor U15865 (N_15865,N_13762,N_14689);
and U15866 (N_15866,N_13742,N_14070);
and U15867 (N_15867,N_14722,N_14359);
nand U15868 (N_15868,N_14610,N_13980);
nand U15869 (N_15869,N_14570,N_14237);
xor U15870 (N_15870,N_14128,N_14519);
or U15871 (N_15871,N_14446,N_14975);
nand U15872 (N_15872,N_14319,N_13889);
xor U15873 (N_15873,N_13875,N_14173);
xor U15874 (N_15874,N_13745,N_13705);
or U15875 (N_15875,N_14279,N_13859);
nor U15876 (N_15876,N_14125,N_13988);
nand U15877 (N_15877,N_14122,N_13697);
xor U15878 (N_15878,N_14203,N_13766);
nand U15879 (N_15879,N_14720,N_14731);
nand U15880 (N_15880,N_13758,N_13882);
xor U15881 (N_15881,N_14285,N_13929);
xnor U15882 (N_15882,N_14985,N_13926);
xor U15883 (N_15883,N_14275,N_14066);
or U15884 (N_15884,N_13631,N_14068);
nor U15885 (N_15885,N_14176,N_13627);
and U15886 (N_15886,N_14685,N_14394);
or U15887 (N_15887,N_13529,N_14325);
and U15888 (N_15888,N_14751,N_14122);
nor U15889 (N_15889,N_14210,N_13782);
or U15890 (N_15890,N_13742,N_14976);
nor U15891 (N_15891,N_14250,N_14590);
or U15892 (N_15892,N_14142,N_14759);
and U15893 (N_15893,N_14098,N_14140);
nand U15894 (N_15894,N_14855,N_13685);
nand U15895 (N_15895,N_14153,N_14546);
or U15896 (N_15896,N_14236,N_14296);
xnor U15897 (N_15897,N_14587,N_14497);
and U15898 (N_15898,N_14303,N_13959);
and U15899 (N_15899,N_14704,N_14617);
nor U15900 (N_15900,N_14967,N_14040);
xnor U15901 (N_15901,N_14232,N_13810);
or U15902 (N_15902,N_14786,N_14362);
or U15903 (N_15903,N_14830,N_14521);
xor U15904 (N_15904,N_14209,N_13689);
or U15905 (N_15905,N_14146,N_14182);
xnor U15906 (N_15906,N_14023,N_14103);
nor U15907 (N_15907,N_13702,N_13691);
or U15908 (N_15908,N_13769,N_14304);
or U15909 (N_15909,N_14862,N_13869);
nor U15910 (N_15910,N_13765,N_14401);
xnor U15911 (N_15911,N_13804,N_14683);
and U15912 (N_15912,N_14519,N_14011);
nand U15913 (N_15913,N_14742,N_13599);
or U15914 (N_15914,N_13730,N_14051);
nand U15915 (N_15915,N_13798,N_13843);
xor U15916 (N_15916,N_14858,N_14154);
nor U15917 (N_15917,N_14456,N_13825);
xnor U15918 (N_15918,N_13932,N_14922);
nand U15919 (N_15919,N_14458,N_14226);
xnor U15920 (N_15920,N_14076,N_14497);
nor U15921 (N_15921,N_14200,N_13539);
xnor U15922 (N_15922,N_14370,N_13657);
xnor U15923 (N_15923,N_14240,N_13737);
xor U15924 (N_15924,N_14593,N_13905);
or U15925 (N_15925,N_14551,N_14336);
or U15926 (N_15926,N_13864,N_14243);
nor U15927 (N_15927,N_13895,N_13926);
or U15928 (N_15928,N_14583,N_14184);
xnor U15929 (N_15929,N_14286,N_13653);
nor U15930 (N_15930,N_14631,N_14664);
nor U15931 (N_15931,N_13670,N_14623);
xor U15932 (N_15932,N_13844,N_14526);
or U15933 (N_15933,N_14407,N_13605);
nor U15934 (N_15934,N_14585,N_14752);
or U15935 (N_15935,N_14248,N_14954);
or U15936 (N_15936,N_14090,N_14954);
or U15937 (N_15937,N_13729,N_14806);
and U15938 (N_15938,N_14134,N_14075);
nor U15939 (N_15939,N_13543,N_13826);
or U15940 (N_15940,N_13880,N_14470);
nand U15941 (N_15941,N_14186,N_14448);
nand U15942 (N_15942,N_14577,N_14198);
nand U15943 (N_15943,N_14087,N_14899);
and U15944 (N_15944,N_14455,N_14639);
nor U15945 (N_15945,N_14042,N_13558);
or U15946 (N_15946,N_14293,N_13679);
xor U15947 (N_15947,N_14389,N_14121);
xor U15948 (N_15948,N_14968,N_14517);
xor U15949 (N_15949,N_14883,N_13647);
xnor U15950 (N_15950,N_14957,N_13652);
and U15951 (N_15951,N_14208,N_14513);
or U15952 (N_15952,N_13847,N_13965);
or U15953 (N_15953,N_14809,N_13839);
nor U15954 (N_15954,N_14659,N_14470);
nand U15955 (N_15955,N_14163,N_14194);
xor U15956 (N_15956,N_13534,N_13909);
or U15957 (N_15957,N_14546,N_14755);
nor U15958 (N_15958,N_14313,N_14108);
nor U15959 (N_15959,N_13927,N_13550);
xnor U15960 (N_15960,N_14110,N_13846);
or U15961 (N_15961,N_14323,N_14741);
xor U15962 (N_15962,N_14678,N_13582);
and U15963 (N_15963,N_14944,N_14566);
and U15964 (N_15964,N_13648,N_13667);
and U15965 (N_15965,N_14069,N_14726);
xnor U15966 (N_15966,N_14142,N_13525);
nor U15967 (N_15967,N_13554,N_13826);
nor U15968 (N_15968,N_14870,N_13599);
xnor U15969 (N_15969,N_14878,N_14962);
or U15970 (N_15970,N_14733,N_13783);
nor U15971 (N_15971,N_14543,N_14852);
or U15972 (N_15972,N_14045,N_14102);
nor U15973 (N_15973,N_13954,N_14950);
xnor U15974 (N_15974,N_14285,N_13768);
and U15975 (N_15975,N_14534,N_13573);
nand U15976 (N_15976,N_13540,N_14024);
or U15977 (N_15977,N_14853,N_14977);
nor U15978 (N_15978,N_14078,N_13853);
or U15979 (N_15979,N_13962,N_14611);
or U15980 (N_15980,N_14582,N_14491);
xor U15981 (N_15981,N_13540,N_14036);
nor U15982 (N_15982,N_13798,N_14719);
nand U15983 (N_15983,N_14977,N_14978);
or U15984 (N_15984,N_14972,N_14620);
nor U15985 (N_15985,N_13854,N_14837);
xnor U15986 (N_15986,N_14847,N_13518);
nand U15987 (N_15987,N_14374,N_14832);
nand U15988 (N_15988,N_13574,N_14974);
or U15989 (N_15989,N_14833,N_13695);
nor U15990 (N_15990,N_14684,N_14289);
nor U15991 (N_15991,N_14536,N_13996);
and U15992 (N_15992,N_14785,N_14201);
or U15993 (N_15993,N_14636,N_13762);
nand U15994 (N_15994,N_14392,N_13727);
or U15995 (N_15995,N_14376,N_14145);
nand U15996 (N_15996,N_14209,N_13912);
nor U15997 (N_15997,N_14846,N_13587);
and U15998 (N_15998,N_13677,N_13602);
and U15999 (N_15999,N_13565,N_14018);
and U16000 (N_16000,N_14402,N_14033);
nand U16001 (N_16001,N_13605,N_14122);
nand U16002 (N_16002,N_13620,N_13993);
or U16003 (N_16003,N_13608,N_14962);
xor U16004 (N_16004,N_14998,N_14304);
xnor U16005 (N_16005,N_14498,N_14874);
xor U16006 (N_16006,N_14076,N_14445);
xor U16007 (N_16007,N_13734,N_14444);
or U16008 (N_16008,N_14003,N_14749);
nand U16009 (N_16009,N_13742,N_14231);
or U16010 (N_16010,N_14596,N_14929);
and U16011 (N_16011,N_14084,N_13840);
nand U16012 (N_16012,N_13694,N_13673);
or U16013 (N_16013,N_13637,N_14234);
xor U16014 (N_16014,N_14119,N_14088);
nand U16015 (N_16015,N_14789,N_14674);
and U16016 (N_16016,N_14157,N_13555);
or U16017 (N_16017,N_14370,N_14524);
nand U16018 (N_16018,N_13888,N_13609);
and U16019 (N_16019,N_14287,N_14846);
and U16020 (N_16020,N_14373,N_14184);
or U16021 (N_16021,N_13507,N_14885);
and U16022 (N_16022,N_14217,N_13731);
or U16023 (N_16023,N_14410,N_14264);
and U16024 (N_16024,N_13501,N_14996);
nand U16025 (N_16025,N_13510,N_13707);
xnor U16026 (N_16026,N_13659,N_13829);
and U16027 (N_16027,N_14087,N_13598);
nand U16028 (N_16028,N_14652,N_14759);
xor U16029 (N_16029,N_13506,N_14676);
xnor U16030 (N_16030,N_14323,N_14612);
or U16031 (N_16031,N_13819,N_14544);
xnor U16032 (N_16032,N_14095,N_14532);
nand U16033 (N_16033,N_14598,N_14099);
xor U16034 (N_16034,N_13862,N_14328);
nand U16035 (N_16035,N_14498,N_14639);
nand U16036 (N_16036,N_13951,N_13738);
and U16037 (N_16037,N_13811,N_14256);
or U16038 (N_16038,N_13922,N_14986);
nor U16039 (N_16039,N_14959,N_14670);
nand U16040 (N_16040,N_13590,N_14080);
nand U16041 (N_16041,N_14384,N_14416);
nand U16042 (N_16042,N_14048,N_14259);
and U16043 (N_16043,N_13696,N_13804);
nand U16044 (N_16044,N_14629,N_14788);
and U16045 (N_16045,N_14704,N_14871);
nand U16046 (N_16046,N_13963,N_14706);
nor U16047 (N_16047,N_14241,N_14879);
nand U16048 (N_16048,N_14955,N_14349);
nand U16049 (N_16049,N_14348,N_14958);
and U16050 (N_16050,N_14337,N_14979);
nor U16051 (N_16051,N_14470,N_14569);
or U16052 (N_16052,N_14851,N_14075);
nor U16053 (N_16053,N_14504,N_14213);
or U16054 (N_16054,N_13851,N_13730);
and U16055 (N_16055,N_14432,N_13720);
xnor U16056 (N_16056,N_14573,N_13706);
xor U16057 (N_16057,N_14678,N_13741);
and U16058 (N_16058,N_13573,N_14628);
nand U16059 (N_16059,N_14797,N_14034);
or U16060 (N_16060,N_14757,N_13518);
or U16061 (N_16061,N_13785,N_14711);
or U16062 (N_16062,N_14359,N_14091);
xor U16063 (N_16063,N_13769,N_13818);
or U16064 (N_16064,N_14711,N_13813);
xor U16065 (N_16065,N_14379,N_13647);
and U16066 (N_16066,N_14059,N_13991);
xnor U16067 (N_16067,N_14982,N_14991);
nand U16068 (N_16068,N_13759,N_14332);
and U16069 (N_16069,N_14923,N_13935);
or U16070 (N_16070,N_13571,N_14631);
and U16071 (N_16071,N_13795,N_14667);
nand U16072 (N_16072,N_13739,N_14230);
nand U16073 (N_16073,N_14320,N_14745);
or U16074 (N_16074,N_14493,N_13686);
nor U16075 (N_16075,N_14528,N_14939);
xnor U16076 (N_16076,N_14738,N_14385);
and U16077 (N_16077,N_13565,N_14597);
xnor U16078 (N_16078,N_13947,N_14046);
nand U16079 (N_16079,N_14006,N_14053);
nor U16080 (N_16080,N_14739,N_14983);
nand U16081 (N_16081,N_13655,N_13587);
nor U16082 (N_16082,N_14891,N_13994);
and U16083 (N_16083,N_13799,N_13842);
nor U16084 (N_16084,N_13692,N_13734);
xnor U16085 (N_16085,N_14623,N_14065);
nor U16086 (N_16086,N_14971,N_13740);
xnor U16087 (N_16087,N_13872,N_13571);
nand U16088 (N_16088,N_14338,N_14641);
or U16089 (N_16089,N_14665,N_13745);
or U16090 (N_16090,N_14856,N_14055);
nor U16091 (N_16091,N_14994,N_13661);
nand U16092 (N_16092,N_14852,N_14653);
xnor U16093 (N_16093,N_14967,N_14880);
and U16094 (N_16094,N_13789,N_13633);
nor U16095 (N_16095,N_13747,N_14175);
nand U16096 (N_16096,N_13641,N_13989);
nor U16097 (N_16097,N_14896,N_13571);
or U16098 (N_16098,N_14779,N_14475);
and U16099 (N_16099,N_14798,N_13856);
xnor U16100 (N_16100,N_14012,N_14095);
nor U16101 (N_16101,N_13670,N_14754);
xor U16102 (N_16102,N_13637,N_13523);
or U16103 (N_16103,N_14848,N_14705);
and U16104 (N_16104,N_13731,N_14271);
or U16105 (N_16105,N_13604,N_13946);
xnor U16106 (N_16106,N_14212,N_14297);
nor U16107 (N_16107,N_13839,N_14640);
or U16108 (N_16108,N_14775,N_14641);
and U16109 (N_16109,N_14814,N_13721);
and U16110 (N_16110,N_13575,N_13676);
xnor U16111 (N_16111,N_14448,N_14981);
and U16112 (N_16112,N_14905,N_14172);
xor U16113 (N_16113,N_14551,N_14406);
nand U16114 (N_16114,N_14728,N_13547);
nand U16115 (N_16115,N_13522,N_13648);
nand U16116 (N_16116,N_14980,N_14052);
nor U16117 (N_16117,N_13597,N_14952);
nand U16118 (N_16118,N_14562,N_13780);
nand U16119 (N_16119,N_13855,N_14768);
and U16120 (N_16120,N_14996,N_13559);
and U16121 (N_16121,N_14580,N_14980);
nor U16122 (N_16122,N_14138,N_14901);
xnor U16123 (N_16123,N_14095,N_14053);
and U16124 (N_16124,N_14448,N_13779);
or U16125 (N_16125,N_14148,N_14697);
xor U16126 (N_16126,N_13512,N_13689);
nor U16127 (N_16127,N_14044,N_13877);
nor U16128 (N_16128,N_14691,N_14022);
nor U16129 (N_16129,N_13625,N_14703);
and U16130 (N_16130,N_13510,N_13545);
xnor U16131 (N_16131,N_14274,N_14497);
nor U16132 (N_16132,N_14675,N_14445);
and U16133 (N_16133,N_13831,N_13835);
nor U16134 (N_16134,N_14353,N_13615);
nor U16135 (N_16135,N_14077,N_14807);
nor U16136 (N_16136,N_14312,N_14690);
and U16137 (N_16137,N_14701,N_13805);
nor U16138 (N_16138,N_14244,N_14021);
or U16139 (N_16139,N_14594,N_14406);
or U16140 (N_16140,N_14496,N_14941);
and U16141 (N_16141,N_14495,N_14043);
and U16142 (N_16142,N_14263,N_13666);
and U16143 (N_16143,N_14000,N_13683);
nand U16144 (N_16144,N_14241,N_14010);
and U16145 (N_16145,N_13583,N_13663);
nor U16146 (N_16146,N_14786,N_13742);
or U16147 (N_16147,N_14167,N_14877);
nor U16148 (N_16148,N_13568,N_13518);
nand U16149 (N_16149,N_14155,N_14917);
nand U16150 (N_16150,N_13967,N_14609);
and U16151 (N_16151,N_14579,N_14493);
nand U16152 (N_16152,N_14728,N_13959);
nand U16153 (N_16153,N_14877,N_14600);
nand U16154 (N_16154,N_13730,N_14808);
and U16155 (N_16155,N_13511,N_14245);
nor U16156 (N_16156,N_13611,N_14786);
nand U16157 (N_16157,N_13638,N_14907);
xnor U16158 (N_16158,N_14130,N_14828);
and U16159 (N_16159,N_14089,N_14569);
or U16160 (N_16160,N_13959,N_13537);
xnor U16161 (N_16161,N_14100,N_14062);
and U16162 (N_16162,N_13609,N_14538);
nor U16163 (N_16163,N_14011,N_14761);
xnor U16164 (N_16164,N_13608,N_14651);
xor U16165 (N_16165,N_13700,N_13904);
nand U16166 (N_16166,N_14723,N_14160);
xor U16167 (N_16167,N_14481,N_14560);
or U16168 (N_16168,N_13837,N_13633);
and U16169 (N_16169,N_14929,N_14047);
or U16170 (N_16170,N_14433,N_14515);
xnor U16171 (N_16171,N_13723,N_14350);
or U16172 (N_16172,N_14560,N_14316);
or U16173 (N_16173,N_13607,N_14787);
nor U16174 (N_16174,N_14493,N_13893);
xor U16175 (N_16175,N_14707,N_14360);
or U16176 (N_16176,N_14362,N_14688);
xnor U16177 (N_16177,N_13636,N_13831);
or U16178 (N_16178,N_13653,N_14711);
xor U16179 (N_16179,N_13773,N_14805);
nand U16180 (N_16180,N_14730,N_14770);
nor U16181 (N_16181,N_14320,N_13687);
nor U16182 (N_16182,N_14894,N_14144);
nor U16183 (N_16183,N_14224,N_14265);
and U16184 (N_16184,N_13750,N_14161);
and U16185 (N_16185,N_13978,N_14965);
nor U16186 (N_16186,N_13760,N_14695);
nor U16187 (N_16187,N_14839,N_14982);
or U16188 (N_16188,N_13931,N_13659);
and U16189 (N_16189,N_13760,N_14526);
or U16190 (N_16190,N_14657,N_14356);
nor U16191 (N_16191,N_14086,N_14960);
nand U16192 (N_16192,N_13535,N_14561);
nand U16193 (N_16193,N_14120,N_13901);
xor U16194 (N_16194,N_14310,N_14839);
or U16195 (N_16195,N_14124,N_13663);
nor U16196 (N_16196,N_14390,N_13514);
or U16197 (N_16197,N_14609,N_14815);
xnor U16198 (N_16198,N_14308,N_13806);
and U16199 (N_16199,N_14408,N_13784);
and U16200 (N_16200,N_14490,N_14800);
nor U16201 (N_16201,N_13617,N_14368);
nand U16202 (N_16202,N_14919,N_14578);
nor U16203 (N_16203,N_14612,N_13601);
or U16204 (N_16204,N_14673,N_14965);
or U16205 (N_16205,N_13751,N_13893);
nor U16206 (N_16206,N_14298,N_13970);
and U16207 (N_16207,N_14282,N_14005);
xnor U16208 (N_16208,N_13994,N_14667);
xnor U16209 (N_16209,N_13739,N_14163);
nor U16210 (N_16210,N_14961,N_13971);
nor U16211 (N_16211,N_14813,N_14338);
or U16212 (N_16212,N_14704,N_13926);
and U16213 (N_16213,N_13862,N_14042);
xor U16214 (N_16214,N_13815,N_13761);
nand U16215 (N_16215,N_14632,N_13949);
and U16216 (N_16216,N_14995,N_13526);
or U16217 (N_16217,N_14302,N_14472);
nor U16218 (N_16218,N_14710,N_13509);
nor U16219 (N_16219,N_14934,N_13701);
or U16220 (N_16220,N_14548,N_13518);
xnor U16221 (N_16221,N_14904,N_14734);
and U16222 (N_16222,N_14051,N_14527);
nor U16223 (N_16223,N_13968,N_14303);
and U16224 (N_16224,N_14092,N_14031);
and U16225 (N_16225,N_14612,N_13865);
nand U16226 (N_16226,N_14877,N_13529);
nor U16227 (N_16227,N_14869,N_14522);
nand U16228 (N_16228,N_14837,N_14403);
nor U16229 (N_16229,N_14609,N_14767);
nor U16230 (N_16230,N_14074,N_14326);
nand U16231 (N_16231,N_14442,N_14953);
xnor U16232 (N_16232,N_14096,N_14368);
nand U16233 (N_16233,N_14718,N_14241);
xor U16234 (N_16234,N_14643,N_14293);
and U16235 (N_16235,N_13558,N_13974);
xnor U16236 (N_16236,N_13507,N_14623);
or U16237 (N_16237,N_13742,N_14544);
and U16238 (N_16238,N_13720,N_14437);
nand U16239 (N_16239,N_14764,N_13752);
and U16240 (N_16240,N_13613,N_14171);
nand U16241 (N_16241,N_14750,N_14629);
nor U16242 (N_16242,N_14998,N_13789);
nor U16243 (N_16243,N_14153,N_14476);
and U16244 (N_16244,N_13949,N_14708);
and U16245 (N_16245,N_13884,N_14566);
nor U16246 (N_16246,N_14234,N_14269);
nor U16247 (N_16247,N_14131,N_13626);
nor U16248 (N_16248,N_13887,N_14587);
and U16249 (N_16249,N_13714,N_14906);
nand U16250 (N_16250,N_14875,N_13535);
and U16251 (N_16251,N_14571,N_13632);
xor U16252 (N_16252,N_13743,N_14839);
and U16253 (N_16253,N_14953,N_14137);
nand U16254 (N_16254,N_14523,N_14478);
and U16255 (N_16255,N_14246,N_14467);
nor U16256 (N_16256,N_14810,N_14855);
nor U16257 (N_16257,N_14715,N_14064);
and U16258 (N_16258,N_14470,N_14199);
or U16259 (N_16259,N_14460,N_13582);
xnor U16260 (N_16260,N_13971,N_14988);
or U16261 (N_16261,N_14987,N_13541);
xnor U16262 (N_16262,N_14812,N_14649);
and U16263 (N_16263,N_14336,N_14365);
or U16264 (N_16264,N_14232,N_14733);
and U16265 (N_16265,N_14532,N_13902);
nand U16266 (N_16266,N_13840,N_13878);
nor U16267 (N_16267,N_14304,N_14845);
or U16268 (N_16268,N_13861,N_14583);
or U16269 (N_16269,N_14616,N_14220);
nand U16270 (N_16270,N_14537,N_14938);
or U16271 (N_16271,N_14960,N_13660);
nand U16272 (N_16272,N_14255,N_14264);
xnor U16273 (N_16273,N_14211,N_14369);
nand U16274 (N_16274,N_14592,N_14871);
nor U16275 (N_16275,N_14575,N_13791);
nor U16276 (N_16276,N_14837,N_13555);
or U16277 (N_16277,N_14542,N_13928);
nor U16278 (N_16278,N_13536,N_13971);
nand U16279 (N_16279,N_13596,N_14485);
and U16280 (N_16280,N_14052,N_13628);
nor U16281 (N_16281,N_14415,N_14502);
xor U16282 (N_16282,N_13618,N_14173);
nor U16283 (N_16283,N_14743,N_14805);
nor U16284 (N_16284,N_13653,N_13535);
nand U16285 (N_16285,N_14663,N_14356);
xor U16286 (N_16286,N_14774,N_14963);
xnor U16287 (N_16287,N_13720,N_14048);
and U16288 (N_16288,N_13740,N_14177);
nand U16289 (N_16289,N_14321,N_14993);
and U16290 (N_16290,N_14204,N_13589);
nor U16291 (N_16291,N_13908,N_14749);
nand U16292 (N_16292,N_13898,N_14941);
xor U16293 (N_16293,N_14531,N_14383);
or U16294 (N_16294,N_14419,N_14568);
and U16295 (N_16295,N_13936,N_13721);
or U16296 (N_16296,N_14304,N_14381);
or U16297 (N_16297,N_14270,N_14730);
nand U16298 (N_16298,N_13643,N_13529);
or U16299 (N_16299,N_13597,N_13541);
or U16300 (N_16300,N_14179,N_14576);
xnor U16301 (N_16301,N_13505,N_14028);
and U16302 (N_16302,N_14971,N_13547);
or U16303 (N_16303,N_13633,N_13903);
and U16304 (N_16304,N_13602,N_14232);
nor U16305 (N_16305,N_13944,N_14394);
and U16306 (N_16306,N_14928,N_13840);
and U16307 (N_16307,N_14023,N_13543);
and U16308 (N_16308,N_14761,N_14762);
nand U16309 (N_16309,N_14563,N_14726);
nor U16310 (N_16310,N_13723,N_14708);
and U16311 (N_16311,N_14055,N_14931);
or U16312 (N_16312,N_14797,N_14361);
nand U16313 (N_16313,N_14380,N_14921);
and U16314 (N_16314,N_14847,N_14157);
xnor U16315 (N_16315,N_13932,N_14532);
or U16316 (N_16316,N_14814,N_14110);
nor U16317 (N_16317,N_13870,N_14636);
and U16318 (N_16318,N_14822,N_13656);
nor U16319 (N_16319,N_14511,N_14680);
nand U16320 (N_16320,N_14550,N_14303);
nand U16321 (N_16321,N_14183,N_14829);
xnor U16322 (N_16322,N_14031,N_14628);
and U16323 (N_16323,N_14570,N_13607);
and U16324 (N_16324,N_14207,N_14263);
nand U16325 (N_16325,N_14328,N_13659);
and U16326 (N_16326,N_13512,N_14993);
xor U16327 (N_16327,N_14962,N_13821);
xnor U16328 (N_16328,N_14509,N_13585);
nand U16329 (N_16329,N_14398,N_14419);
or U16330 (N_16330,N_14242,N_14370);
nand U16331 (N_16331,N_14947,N_14938);
or U16332 (N_16332,N_14306,N_14424);
nand U16333 (N_16333,N_13563,N_14419);
nor U16334 (N_16334,N_13636,N_13960);
and U16335 (N_16335,N_14663,N_14362);
and U16336 (N_16336,N_14486,N_14412);
xnor U16337 (N_16337,N_14021,N_14732);
xnor U16338 (N_16338,N_14304,N_14612);
and U16339 (N_16339,N_14317,N_14946);
xor U16340 (N_16340,N_14220,N_14961);
nor U16341 (N_16341,N_14817,N_13673);
or U16342 (N_16342,N_14962,N_14537);
nand U16343 (N_16343,N_14681,N_14738);
or U16344 (N_16344,N_13660,N_13586);
nor U16345 (N_16345,N_14509,N_13867);
or U16346 (N_16346,N_14552,N_14401);
nand U16347 (N_16347,N_14719,N_13921);
or U16348 (N_16348,N_13594,N_14235);
or U16349 (N_16349,N_14391,N_14520);
nand U16350 (N_16350,N_14931,N_14037);
and U16351 (N_16351,N_14998,N_13620);
and U16352 (N_16352,N_13711,N_13628);
nor U16353 (N_16353,N_14031,N_14781);
and U16354 (N_16354,N_13716,N_14459);
nand U16355 (N_16355,N_14439,N_14958);
and U16356 (N_16356,N_14874,N_14006);
xor U16357 (N_16357,N_14344,N_14700);
or U16358 (N_16358,N_14242,N_14018);
and U16359 (N_16359,N_14638,N_13585);
and U16360 (N_16360,N_14268,N_13780);
or U16361 (N_16361,N_13895,N_14561);
nand U16362 (N_16362,N_14915,N_14892);
and U16363 (N_16363,N_14612,N_14309);
or U16364 (N_16364,N_14272,N_13521);
and U16365 (N_16365,N_14204,N_13966);
and U16366 (N_16366,N_14328,N_14417);
xnor U16367 (N_16367,N_14033,N_13915);
or U16368 (N_16368,N_13869,N_14690);
and U16369 (N_16369,N_14969,N_14420);
xor U16370 (N_16370,N_14693,N_13976);
and U16371 (N_16371,N_13539,N_13694);
xnor U16372 (N_16372,N_14877,N_13681);
xnor U16373 (N_16373,N_13542,N_14133);
nand U16374 (N_16374,N_14280,N_14188);
or U16375 (N_16375,N_14884,N_13589);
or U16376 (N_16376,N_14486,N_13930);
xor U16377 (N_16377,N_14383,N_14873);
xor U16378 (N_16378,N_14738,N_13916);
nor U16379 (N_16379,N_14765,N_14204);
and U16380 (N_16380,N_13797,N_13736);
xor U16381 (N_16381,N_14983,N_13526);
and U16382 (N_16382,N_14871,N_14821);
xor U16383 (N_16383,N_13575,N_14185);
or U16384 (N_16384,N_14005,N_14592);
nor U16385 (N_16385,N_14432,N_14462);
and U16386 (N_16386,N_13648,N_13755);
nor U16387 (N_16387,N_14418,N_13784);
nor U16388 (N_16388,N_13693,N_13581);
nand U16389 (N_16389,N_13806,N_14529);
and U16390 (N_16390,N_14860,N_14551);
nor U16391 (N_16391,N_14011,N_13552);
and U16392 (N_16392,N_13798,N_13853);
or U16393 (N_16393,N_14315,N_14017);
nand U16394 (N_16394,N_13685,N_13697);
xnor U16395 (N_16395,N_13681,N_14496);
and U16396 (N_16396,N_14844,N_13821);
xor U16397 (N_16397,N_14936,N_14947);
xor U16398 (N_16398,N_14814,N_13779);
nand U16399 (N_16399,N_13581,N_13686);
or U16400 (N_16400,N_13975,N_14841);
or U16401 (N_16401,N_14740,N_14248);
nand U16402 (N_16402,N_13640,N_14140);
nand U16403 (N_16403,N_14072,N_13806);
or U16404 (N_16404,N_13553,N_13721);
nor U16405 (N_16405,N_14262,N_14023);
or U16406 (N_16406,N_14828,N_14833);
xor U16407 (N_16407,N_14005,N_14710);
and U16408 (N_16408,N_14578,N_14926);
and U16409 (N_16409,N_14727,N_14369);
and U16410 (N_16410,N_14601,N_13773);
and U16411 (N_16411,N_14799,N_14346);
nor U16412 (N_16412,N_14884,N_13719);
or U16413 (N_16413,N_14927,N_14731);
xnor U16414 (N_16414,N_14579,N_14845);
or U16415 (N_16415,N_14540,N_14840);
xnor U16416 (N_16416,N_14501,N_13726);
nand U16417 (N_16417,N_14409,N_13631);
nor U16418 (N_16418,N_13714,N_14818);
nand U16419 (N_16419,N_14720,N_14895);
or U16420 (N_16420,N_14194,N_13730);
xnor U16421 (N_16421,N_14990,N_14475);
nand U16422 (N_16422,N_14379,N_14653);
or U16423 (N_16423,N_13991,N_14983);
and U16424 (N_16424,N_14760,N_13777);
nor U16425 (N_16425,N_14251,N_13769);
or U16426 (N_16426,N_13781,N_14752);
nand U16427 (N_16427,N_14272,N_14958);
nand U16428 (N_16428,N_14273,N_14197);
nor U16429 (N_16429,N_14233,N_14449);
nand U16430 (N_16430,N_13778,N_13756);
nand U16431 (N_16431,N_14262,N_14997);
nand U16432 (N_16432,N_13512,N_14883);
nand U16433 (N_16433,N_13873,N_14411);
nand U16434 (N_16434,N_14955,N_14169);
and U16435 (N_16435,N_13975,N_14273);
or U16436 (N_16436,N_14845,N_14345);
nand U16437 (N_16437,N_14968,N_14739);
and U16438 (N_16438,N_14351,N_13614);
nor U16439 (N_16439,N_14789,N_13513);
and U16440 (N_16440,N_14152,N_14905);
nor U16441 (N_16441,N_13779,N_14025);
and U16442 (N_16442,N_13575,N_13740);
and U16443 (N_16443,N_13518,N_14220);
and U16444 (N_16444,N_14494,N_13943);
nand U16445 (N_16445,N_14985,N_14311);
nand U16446 (N_16446,N_14704,N_14588);
and U16447 (N_16447,N_13647,N_14355);
or U16448 (N_16448,N_14523,N_14645);
or U16449 (N_16449,N_14289,N_13532);
or U16450 (N_16450,N_13828,N_14761);
or U16451 (N_16451,N_14229,N_14918);
xor U16452 (N_16452,N_14482,N_14659);
xor U16453 (N_16453,N_13604,N_14264);
nor U16454 (N_16454,N_13985,N_14539);
and U16455 (N_16455,N_13638,N_14994);
nor U16456 (N_16456,N_14970,N_13634);
or U16457 (N_16457,N_13701,N_14991);
nand U16458 (N_16458,N_13690,N_13838);
nor U16459 (N_16459,N_14869,N_14534);
or U16460 (N_16460,N_13836,N_14387);
or U16461 (N_16461,N_14212,N_14352);
xnor U16462 (N_16462,N_13678,N_14756);
nor U16463 (N_16463,N_14841,N_13717);
or U16464 (N_16464,N_14373,N_14842);
nor U16465 (N_16465,N_14313,N_14121);
and U16466 (N_16466,N_13837,N_14811);
nand U16467 (N_16467,N_14638,N_13628);
nand U16468 (N_16468,N_13629,N_13697);
nand U16469 (N_16469,N_14799,N_14017);
xor U16470 (N_16470,N_14351,N_14715);
and U16471 (N_16471,N_14637,N_13701);
nand U16472 (N_16472,N_13976,N_13668);
or U16473 (N_16473,N_14393,N_13585);
xnor U16474 (N_16474,N_14109,N_14046);
nor U16475 (N_16475,N_14095,N_14587);
and U16476 (N_16476,N_13522,N_14833);
nor U16477 (N_16477,N_14191,N_13889);
nor U16478 (N_16478,N_14490,N_13733);
nor U16479 (N_16479,N_14715,N_14229);
nor U16480 (N_16480,N_13752,N_13547);
xor U16481 (N_16481,N_14368,N_13670);
xnor U16482 (N_16482,N_14174,N_14984);
nor U16483 (N_16483,N_14439,N_14118);
or U16484 (N_16484,N_14393,N_14063);
nand U16485 (N_16485,N_14492,N_14532);
nor U16486 (N_16486,N_14430,N_14745);
nor U16487 (N_16487,N_14461,N_14445);
nor U16488 (N_16488,N_13882,N_13952);
or U16489 (N_16489,N_13597,N_14648);
nand U16490 (N_16490,N_14623,N_14070);
or U16491 (N_16491,N_14947,N_14771);
or U16492 (N_16492,N_13605,N_14883);
and U16493 (N_16493,N_14988,N_14698);
xnor U16494 (N_16494,N_14071,N_13557);
xnor U16495 (N_16495,N_14779,N_14612);
nor U16496 (N_16496,N_13804,N_14409);
nor U16497 (N_16497,N_14307,N_13714);
xor U16498 (N_16498,N_14596,N_14959);
and U16499 (N_16499,N_14613,N_14810);
and U16500 (N_16500,N_16129,N_16393);
nand U16501 (N_16501,N_16282,N_16356);
and U16502 (N_16502,N_16202,N_16091);
xnor U16503 (N_16503,N_15270,N_15868);
nand U16504 (N_16504,N_15106,N_16418);
nor U16505 (N_16505,N_15289,N_15817);
and U16506 (N_16506,N_16290,N_16402);
xnor U16507 (N_16507,N_15296,N_15521);
xnor U16508 (N_16508,N_15477,N_15355);
nor U16509 (N_16509,N_16030,N_15489);
nor U16510 (N_16510,N_15313,N_15615);
nand U16511 (N_16511,N_15042,N_16307);
and U16512 (N_16512,N_16012,N_15174);
nor U16513 (N_16513,N_15642,N_16027);
or U16514 (N_16514,N_16361,N_16032);
nor U16515 (N_16515,N_16241,N_16126);
nand U16516 (N_16516,N_15170,N_15865);
xnor U16517 (N_16517,N_16112,N_15483);
or U16518 (N_16518,N_15925,N_15882);
xor U16519 (N_16519,N_15857,N_15418);
nor U16520 (N_16520,N_15345,N_15485);
xor U16521 (N_16521,N_16158,N_15150);
xor U16522 (N_16522,N_15705,N_16131);
or U16523 (N_16523,N_15414,N_15332);
or U16524 (N_16524,N_15570,N_15140);
nor U16525 (N_16525,N_15420,N_16221);
xnor U16526 (N_16526,N_15660,N_16054);
xnor U16527 (N_16527,N_15717,N_15478);
and U16528 (N_16528,N_15018,N_16127);
nor U16529 (N_16529,N_15518,N_15305);
xor U16530 (N_16530,N_15585,N_15644);
nand U16531 (N_16531,N_15666,N_15275);
nand U16532 (N_16532,N_15513,N_16218);
nor U16533 (N_16533,N_16355,N_15233);
xnor U16534 (N_16534,N_15582,N_15895);
nand U16535 (N_16535,N_16094,N_15870);
nand U16536 (N_16536,N_16063,N_16020);
xnor U16537 (N_16537,N_15527,N_15331);
nor U16538 (N_16538,N_15720,N_16328);
or U16539 (N_16539,N_15954,N_15424);
nand U16540 (N_16540,N_16254,N_15864);
xor U16541 (N_16541,N_15415,N_15764);
nand U16542 (N_16542,N_16046,N_16024);
xor U16543 (N_16543,N_16234,N_15655);
nand U16544 (N_16544,N_15880,N_15781);
nand U16545 (N_16545,N_15184,N_15397);
nand U16546 (N_16546,N_16199,N_15543);
nor U16547 (N_16547,N_15109,N_15061);
nand U16548 (N_16548,N_15380,N_15166);
and U16549 (N_16549,N_15823,N_15710);
nand U16550 (N_16550,N_15886,N_15678);
xnor U16551 (N_16551,N_15283,N_15059);
nand U16552 (N_16552,N_16277,N_15921);
and U16553 (N_16553,N_15385,N_15529);
and U16554 (N_16554,N_16232,N_15923);
and U16555 (N_16555,N_15920,N_15135);
or U16556 (N_16556,N_16069,N_16117);
xnor U16557 (N_16557,N_16262,N_16476);
xnor U16558 (N_16558,N_16233,N_15503);
nand U16559 (N_16559,N_15645,N_16335);
and U16560 (N_16560,N_15721,N_15006);
nand U16561 (N_16561,N_16392,N_16439);
and U16562 (N_16562,N_15218,N_15494);
xor U16563 (N_16563,N_15152,N_16464);
and U16564 (N_16564,N_16193,N_16113);
and U16565 (N_16565,N_15968,N_15845);
and U16566 (N_16566,N_15984,N_15650);
xnor U16567 (N_16567,N_15099,N_15614);
or U16568 (N_16568,N_15171,N_15998);
or U16569 (N_16569,N_15671,N_15205);
nand U16570 (N_16570,N_16302,N_15287);
xor U16571 (N_16571,N_15439,N_15855);
xor U16572 (N_16572,N_16334,N_15773);
xor U16573 (N_16573,N_16106,N_16414);
nand U16574 (N_16574,N_15273,N_16263);
or U16575 (N_16575,N_16416,N_15123);
and U16576 (N_16576,N_15809,N_15336);
and U16577 (N_16577,N_15465,N_16330);
nand U16578 (N_16578,N_15079,N_15389);
or U16579 (N_16579,N_16042,N_15450);
xor U16580 (N_16580,N_15639,N_15481);
nor U16581 (N_16581,N_15366,N_16403);
nand U16582 (N_16582,N_15155,N_15219);
or U16583 (N_16583,N_15464,N_15738);
nor U16584 (N_16584,N_15442,N_15962);
nor U16585 (N_16585,N_15374,N_15511);
nor U16586 (N_16586,N_15101,N_16279);
or U16587 (N_16587,N_16051,N_15046);
xnor U16588 (N_16588,N_15975,N_16219);
and U16589 (N_16589,N_15593,N_15735);
xor U16590 (N_16590,N_15388,N_16323);
nand U16591 (N_16591,N_16327,N_15310);
nand U16592 (N_16592,N_15144,N_16246);
or U16593 (N_16593,N_16359,N_16107);
or U16594 (N_16594,N_16010,N_15510);
and U16595 (N_16595,N_15567,N_15762);
nand U16596 (N_16596,N_16070,N_15338);
or U16597 (N_16597,N_15562,N_16240);
nand U16598 (N_16598,N_15526,N_15149);
nand U16599 (N_16599,N_15005,N_15110);
or U16600 (N_16600,N_16137,N_15497);
xnor U16601 (N_16601,N_15492,N_15488);
xor U16602 (N_16602,N_15532,N_15276);
nor U16603 (N_16603,N_15167,N_15749);
xnor U16604 (N_16604,N_15300,N_15255);
nand U16605 (N_16605,N_15251,N_15800);
or U16606 (N_16606,N_16289,N_16001);
xnor U16607 (N_16607,N_16159,N_15253);
or U16608 (N_16608,N_15632,N_16130);
nor U16609 (N_16609,N_15182,N_15922);
and U16610 (N_16610,N_16034,N_15957);
and U16611 (N_16611,N_16157,N_15879);
or U16612 (N_16612,N_16469,N_16269);
nor U16613 (N_16613,N_16357,N_15020);
nand U16614 (N_16614,N_16381,N_15154);
and U16615 (N_16615,N_15223,N_16195);
nor U16616 (N_16616,N_15853,N_15832);
nor U16617 (N_16617,N_15986,N_15980);
or U16618 (N_16618,N_15785,N_16311);
and U16619 (N_16619,N_16405,N_15535);
or U16620 (N_16620,N_15556,N_15034);
nand U16621 (N_16621,N_15432,N_15151);
xor U16622 (N_16622,N_15618,N_15969);
and U16623 (N_16623,N_15824,N_15153);
xor U16624 (N_16624,N_16015,N_15209);
xor U16625 (N_16625,N_15013,N_16301);
xnor U16626 (N_16626,N_16033,N_15716);
nor U16627 (N_16627,N_15369,N_15896);
nand U16628 (N_16628,N_16152,N_15353);
xor U16629 (N_16629,N_15673,N_16337);
or U16630 (N_16630,N_15727,N_16205);
or U16631 (N_16631,N_15842,N_16297);
and U16632 (N_16632,N_15568,N_15105);
and U16633 (N_16633,N_15221,N_16494);
nand U16634 (N_16634,N_16299,N_15595);
nor U16635 (N_16635,N_15169,N_15337);
or U16636 (N_16636,N_15772,N_15675);
nor U16637 (N_16637,N_15804,N_16377);
and U16638 (N_16638,N_15220,N_16000);
nor U16639 (N_16639,N_15652,N_15944);
and U16640 (N_16640,N_15907,N_15071);
nand U16641 (N_16641,N_15473,N_16088);
or U16642 (N_16642,N_15722,N_15408);
and U16643 (N_16643,N_15905,N_15941);
or U16644 (N_16644,N_15542,N_15604);
xor U16645 (N_16645,N_16428,N_15016);
nor U16646 (N_16646,N_15976,N_16462);
and U16647 (N_16647,N_15426,N_16179);
nand U16648 (N_16648,N_15351,N_15158);
xor U16649 (N_16649,N_16211,N_15611);
xor U16650 (N_16650,N_15697,N_15288);
and U16651 (N_16651,N_16058,N_15558);
and U16652 (N_16652,N_16288,N_15217);
or U16653 (N_16653,N_15592,N_15603);
xor U16654 (N_16654,N_16076,N_16165);
or U16655 (N_16655,N_15316,N_16273);
nor U16656 (N_16656,N_16372,N_15779);
nor U16657 (N_16657,N_15041,N_15157);
nor U16658 (N_16658,N_15372,N_16135);
nand U16659 (N_16659,N_15656,N_15248);
nor U16660 (N_16660,N_15700,N_15999);
xor U16661 (N_16661,N_15234,N_15029);
xor U16662 (N_16662,N_15789,N_16200);
xor U16663 (N_16663,N_15767,N_15658);
nand U16664 (N_16664,N_15690,N_16090);
nor U16665 (N_16665,N_15928,N_16197);
nand U16666 (N_16666,N_15761,N_15214);
and U16667 (N_16667,N_15626,N_15757);
xor U16668 (N_16668,N_15956,N_15688);
or U16669 (N_16669,N_15576,N_15659);
and U16670 (N_16670,N_15092,N_16239);
or U16671 (N_16671,N_15378,N_15187);
or U16672 (N_16672,N_16400,N_15669);
nor U16673 (N_16673,N_15934,N_15959);
nand U16674 (N_16674,N_16343,N_16097);
xnor U16675 (N_16675,N_15851,N_16217);
nand U16676 (N_16676,N_16440,N_16110);
xor U16677 (N_16677,N_15193,N_15291);
nor U16678 (N_16678,N_16207,N_16248);
and U16679 (N_16679,N_15913,N_15130);
and U16680 (N_16680,N_16102,N_15502);
nand U16681 (N_16681,N_15243,N_16398);
nor U16682 (N_16682,N_16443,N_15884);
xor U16683 (N_16683,N_15327,N_15049);
xor U16684 (N_16684,N_15319,N_15458);
nor U16685 (N_16685,N_15329,N_15470);
or U16686 (N_16686,N_16445,N_16120);
nand U16687 (N_16687,N_15093,N_15814);
nor U16688 (N_16688,N_16116,N_15084);
and U16689 (N_16689,N_15080,N_15569);
or U16690 (N_16690,N_15955,N_15363);
xor U16691 (N_16691,N_15479,N_15294);
nor U16692 (N_16692,N_15280,N_16229);
or U16693 (N_16693,N_15131,N_15816);
or U16694 (N_16694,N_15699,N_15117);
nor U16695 (N_16695,N_15663,N_16118);
nand U16696 (N_16696,N_15204,N_15790);
xor U16697 (N_16697,N_16379,N_16480);
or U16698 (N_16698,N_15547,N_16085);
xor U16699 (N_16699,N_15566,N_16340);
or U16700 (N_16700,N_15958,N_16431);
and U16701 (N_16701,N_15398,N_16047);
nand U16702 (N_16702,N_15610,N_15197);
nor U16703 (N_16703,N_15083,N_16079);
nor U16704 (N_16704,N_16455,N_15805);
and U16705 (N_16705,N_15634,N_15691);
nand U16706 (N_16706,N_15917,N_16139);
or U16707 (N_16707,N_16250,N_16022);
nor U16708 (N_16708,N_16189,N_15755);
and U16709 (N_16709,N_15752,N_15891);
nor U16710 (N_16710,N_16201,N_15770);
and U16711 (N_16711,N_16108,N_15062);
and U16712 (N_16712,N_15517,N_16479);
nand U16713 (N_16713,N_15589,N_15578);
nand U16714 (N_16714,N_15443,N_15163);
nor U16715 (N_16715,N_15508,N_15377);
xor U16716 (N_16716,N_15862,N_15411);
and U16717 (N_16717,N_15616,N_15054);
xor U16718 (N_16718,N_15278,N_15127);
xnor U16719 (N_16719,N_15822,N_15040);
nand U16720 (N_16720,N_15893,N_15082);
or U16721 (N_16721,N_16364,N_16188);
xor U16722 (N_16722,N_16367,N_15608);
xor U16723 (N_16723,N_15146,N_15641);
and U16724 (N_16724,N_15739,N_15201);
and U16725 (N_16725,N_16489,N_15531);
and U16726 (N_16726,N_15022,N_16294);
xor U16727 (N_16727,N_16322,N_15929);
xnor U16728 (N_16728,N_16053,N_15583);
and U16729 (N_16729,N_16222,N_16083);
nor U16730 (N_16730,N_15431,N_15515);
nand U16731 (N_16731,N_15405,N_15269);
and U16732 (N_16732,N_16287,N_15676);
nand U16733 (N_16733,N_15438,N_16089);
nor U16734 (N_16734,N_15587,N_16174);
and U16735 (N_16735,N_15460,N_16345);
or U16736 (N_16736,N_15778,N_15224);
and U16737 (N_16737,N_16348,N_15745);
xnor U16738 (N_16738,N_15335,N_16134);
nor U16739 (N_16739,N_15445,N_16035);
nor U16740 (N_16740,N_15232,N_15088);
and U16741 (N_16741,N_16176,N_16087);
or U16742 (N_16742,N_15216,N_16452);
or U16743 (N_16743,N_16276,N_16007);
or U16744 (N_16744,N_16459,N_15620);
xor U16745 (N_16745,N_15964,N_16298);
or U16746 (N_16746,N_16427,N_16111);
and U16747 (N_16747,N_15407,N_16073);
nor U16748 (N_16748,N_16192,N_15298);
or U16749 (N_16749,N_16040,N_15982);
xnor U16750 (N_16750,N_15776,N_16314);
and U16751 (N_16751,N_16081,N_15831);
xnor U16752 (N_16752,N_15848,N_16317);
and U16753 (N_16753,N_16401,N_16397);
and U16754 (N_16754,N_15238,N_15134);
or U16755 (N_16755,N_16006,N_15333);
xnor U16756 (N_16756,N_16266,N_15413);
or U16757 (N_16757,N_15667,N_16434);
nor U16758 (N_16758,N_15452,N_15965);
xor U16759 (N_16759,N_15320,N_15534);
xor U16760 (N_16760,N_15113,N_15872);
and U16761 (N_16761,N_16346,N_15066);
and U16762 (N_16762,N_16238,N_15693);
or U16763 (N_16763,N_16306,N_15787);
nor U16764 (N_16764,N_15303,N_16169);
nand U16765 (N_16765,N_15813,N_16447);
nor U16766 (N_16766,N_16002,N_15860);
and U16767 (N_16767,N_15875,N_16429);
nand U16768 (N_16768,N_16438,N_16285);
nand U16769 (N_16769,N_15897,N_15729);
nor U16770 (N_16770,N_15318,N_15930);
and U16771 (N_16771,N_15322,N_15522);
xor U16772 (N_16772,N_15876,N_15933);
or U16773 (N_16773,N_15075,N_16100);
xnor U16774 (N_16774,N_15539,N_15836);
nand U16775 (N_16775,N_16312,N_15758);
nor U16776 (N_16776,N_15261,N_15188);
or U16777 (N_16777,N_16153,N_15635);
nor U16778 (N_16778,N_15132,N_15519);
nand U16779 (N_16779,N_15012,N_15212);
and U16780 (N_16780,N_15637,N_16454);
or U16781 (N_16781,N_15780,N_15695);
nor U16782 (N_16782,N_15048,N_15343);
xnor U16783 (N_16783,N_15357,N_15881);
and U16784 (N_16784,N_15803,N_15175);
nand U16785 (N_16785,N_15981,N_15812);
nor U16786 (N_16786,N_15081,N_15834);
xnor U16787 (N_16787,N_16300,N_15376);
and U16788 (N_16788,N_16164,N_15019);
and U16789 (N_16789,N_16442,N_15362);
nor U16790 (N_16790,N_16249,N_16458);
or U16791 (N_16791,N_16268,N_16213);
xor U16792 (N_16792,N_15948,N_15742);
xor U16793 (N_16793,N_15926,N_16077);
and U16794 (N_16794,N_16471,N_15902);
xor U16795 (N_16795,N_16062,N_16064);
and U16796 (N_16796,N_16286,N_15446);
nor U16797 (N_16797,N_16391,N_15936);
nor U16798 (N_16798,N_15708,N_16061);
nand U16799 (N_16799,N_15456,N_16292);
or U16800 (N_16800,N_15723,N_15119);
nor U16801 (N_16801,N_15242,N_16162);
or U16802 (N_16802,N_16466,N_15306);
nor U16803 (N_16803,N_15683,N_16316);
nand U16804 (N_16804,N_16368,N_16426);
nor U16805 (N_16805,N_16208,N_15874);
xor U16806 (N_16806,N_15108,N_15256);
nor U16807 (N_16807,N_15025,N_16242);
or U16808 (N_16808,N_16272,N_15178);
or U16809 (N_16809,N_15828,N_16291);
or U16810 (N_16810,N_15186,N_16161);
nor U16811 (N_16811,N_16399,N_15472);
and U16812 (N_16812,N_16123,N_15590);
nor U16813 (N_16813,N_15441,N_15661);
and U16814 (N_16814,N_16320,N_15349);
or U16815 (N_16815,N_16407,N_15994);
nor U16816 (N_16816,N_15194,N_15286);
xor U16817 (N_16817,N_15943,N_16339);
nor U16818 (N_16818,N_15989,N_16460);
xnor U16819 (N_16819,N_15867,N_15859);
xnor U16820 (N_16820,N_15509,N_15487);
and U16821 (N_16821,N_16499,N_15039);
nand U16822 (N_16822,N_15401,N_15885);
and U16823 (N_16823,N_15474,N_15341);
or U16824 (N_16824,N_16244,N_15403);
and U16825 (N_16825,N_15903,N_15490);
nor U16826 (N_16826,N_16037,N_16004);
nor U16827 (N_16827,N_15706,N_15577);
nor U16828 (N_16828,N_15475,N_16009);
nor U16829 (N_16829,N_15138,N_15505);
and U16830 (N_16830,N_16347,N_15978);
xnor U16831 (N_16831,N_16421,N_15966);
nor U16832 (N_16832,N_15364,N_16257);
nor U16833 (N_16833,N_15172,N_15765);
xor U16834 (N_16834,N_15370,N_15808);
xor U16835 (N_16835,N_15588,N_15074);
or U16836 (N_16836,N_15674,N_15581);
and U16837 (N_16837,N_16114,N_16374);
xor U16838 (N_16838,N_15001,N_15326);
or U16839 (N_16839,N_16470,N_15392);
nor U16840 (N_16840,N_15686,N_15419);
xnor U16841 (N_16841,N_16016,N_15584);
xnor U16842 (N_16842,N_15866,N_15440);
xor U16843 (N_16843,N_16336,N_16492);
and U16844 (N_16844,N_15199,N_15546);
or U16845 (N_16845,N_15116,N_15493);
nand U16846 (N_16846,N_16080,N_15908);
nand U16847 (N_16847,N_15334,N_15664);
nand U16848 (N_16848,N_15536,N_16209);
or U16849 (N_16849,N_15878,N_16082);
nand U16850 (N_16850,N_15476,N_15843);
nor U16851 (N_16851,N_15340,N_16332);
xnor U16852 (N_16852,N_16166,N_15679);
or U16853 (N_16853,N_15931,N_15602);
or U16854 (N_16854,N_15670,N_15121);
nand U16855 (N_16855,N_15753,N_15871);
or U16856 (N_16856,N_15798,N_15555);
nand U16857 (N_16857,N_15990,N_16256);
nand U16858 (N_16858,N_15246,N_15628);
and U16859 (N_16859,N_16086,N_16408);
or U16860 (N_16860,N_15680,N_15482);
and U16861 (N_16861,N_15573,N_15837);
xnor U16862 (N_16862,N_15266,N_16358);
nand U16863 (N_16863,N_16493,N_15324);
or U16864 (N_16864,N_16338,N_15709);
nor U16865 (N_16865,N_15947,N_15077);
nor U16866 (N_16866,N_15437,N_15356);
or U16867 (N_16867,N_16145,N_16321);
nor U16868 (N_16868,N_16142,N_15942);
nand U16869 (N_16869,N_15821,N_15299);
and U16870 (N_16870,N_15888,N_15089);
and U16871 (N_16871,N_15972,N_15231);
xor U16872 (N_16872,N_15346,N_15451);
nor U16873 (N_16873,N_16215,N_15330);
nand U16874 (N_16874,N_16092,N_16423);
nand U16875 (N_16875,N_15838,N_15030);
or U16876 (N_16876,N_15466,N_15284);
xor U16877 (N_16877,N_16052,N_15008);
nor U16878 (N_16878,N_15459,N_15643);
xnor U16879 (N_16879,N_15685,N_15455);
nor U16880 (N_16880,N_16183,N_15128);
nand U16881 (N_16881,N_15198,N_16160);
nor U16882 (N_16882,N_15094,N_15560);
xnor U16883 (N_16883,N_15057,N_15003);
nor U16884 (N_16884,N_16031,N_15987);
or U16885 (N_16885,N_15579,N_16444);
nor U16886 (N_16886,N_16147,N_16206);
or U16887 (N_16887,N_15394,N_15145);
or U16888 (N_16888,N_16333,N_15367);
nand U16889 (N_16889,N_15185,N_15382);
nand U16890 (N_16890,N_16072,N_15846);
nand U16891 (N_16891,N_15501,N_16017);
nor U16892 (N_16892,N_16475,N_16484);
or U16893 (N_16893,N_15937,N_15953);
or U16894 (N_16894,N_16156,N_15468);
or U16895 (N_16895,N_15741,N_15599);
and U16896 (N_16896,N_15997,N_15769);
and U16897 (N_16897,N_15010,N_15391);
xor U16898 (N_16898,N_15651,N_15436);
xnor U16899 (N_16899,N_15000,N_15743);
and U16900 (N_16900,N_15347,N_15935);
or U16901 (N_16901,N_15533,N_15354);
nor U16902 (N_16902,N_16225,N_16406);
xor U16903 (N_16903,N_15156,N_15317);
nor U16904 (N_16904,N_16280,N_15839);
nor U16905 (N_16905,N_16253,N_15596);
nor U16906 (N_16906,N_16498,N_15085);
xnor U16907 (N_16907,N_15967,N_15811);
and U16908 (N_16908,N_16212,N_15552);
or U16909 (N_16909,N_15726,N_15551);
nor U16910 (N_16910,N_15133,N_15429);
xnor U16911 (N_16911,N_15033,N_15946);
or U16912 (N_16912,N_15028,N_15325);
and U16913 (N_16913,N_15572,N_16275);
nand U16914 (N_16914,N_16132,N_16141);
nand U16915 (N_16915,N_15919,N_15538);
nand U16916 (N_16916,N_15307,N_15985);
and U16917 (N_16917,N_15023,N_16191);
and U16918 (N_16918,N_16260,N_16483);
and U16919 (N_16919,N_15629,N_16344);
or U16920 (N_16920,N_15906,N_15229);
xnor U16921 (N_16921,N_15350,N_15754);
xnor U16922 (N_16922,N_15909,N_15724);
nand U16923 (N_16923,N_15203,N_16420);
xnor U16924 (N_16924,N_15236,N_16468);
and U16925 (N_16925,N_16023,N_15107);
xor U16926 (N_16926,N_15887,N_15207);
nor U16927 (N_16927,N_15952,N_16048);
nand U16928 (N_16928,N_16055,N_15949);
nor U16929 (N_16929,N_15196,N_15715);
nand U16930 (N_16930,N_16038,N_15177);
nand U16931 (N_16931,N_16425,N_15621);
nor U16932 (N_16932,N_16236,N_15444);
nor U16933 (N_16933,N_15496,N_15889);
nor U16934 (N_16934,N_15574,N_16382);
nor U16935 (N_16935,N_16371,N_15321);
and U16936 (N_16936,N_16119,N_15063);
or U16937 (N_16937,N_15247,N_15262);
nor U16938 (N_16938,N_15545,N_15924);
nor U16939 (N_16939,N_15192,N_15227);
or U16940 (N_16940,N_16295,N_16284);
or U16941 (N_16941,N_15512,N_15662);
or U16942 (N_16942,N_16021,N_15282);
nor U16943 (N_16943,N_15375,N_15737);
nand U16944 (N_16944,N_15802,N_16411);
nor U16945 (N_16945,N_15544,N_16384);
and U16946 (N_16946,N_15179,N_15939);
nor U16947 (N_16947,N_16354,N_16180);
nand U16948 (N_16948,N_15553,N_16036);
and U16949 (N_16949,N_16049,N_15598);
or U16950 (N_16950,N_16331,N_15250);
nor U16951 (N_16951,N_15368,N_15387);
or U16952 (N_16952,N_16496,N_16005);
nor U16953 (N_16953,N_15974,N_15359);
nand U16954 (N_16954,N_15344,N_15215);
xor U16955 (N_16955,N_15036,N_15180);
or U16956 (N_16956,N_16151,N_15731);
xnor U16957 (N_16957,N_15206,N_16025);
or U16958 (N_16958,N_15393,N_15744);
nand U16959 (N_16959,N_15076,N_16278);
xor U16960 (N_16960,N_15467,N_16366);
and U16961 (N_16961,N_15580,N_15308);
xnor U16962 (N_16962,N_16437,N_16148);
nor U16963 (N_16963,N_15225,N_15711);
xnor U16964 (N_16964,N_15993,N_16318);
nand U16965 (N_16965,N_16430,N_16274);
xor U16966 (N_16966,N_15636,N_16448);
nor U16967 (N_16967,N_15771,N_16446);
nand U16968 (N_16968,N_15449,N_16154);
nand U16969 (N_16969,N_15073,N_15830);
and U16970 (N_16970,N_15396,N_15672);
or U16971 (N_16971,N_16303,N_16495);
or U16972 (N_16972,N_15486,N_16243);
nor U16973 (N_16973,N_15202,N_16473);
or U16974 (N_16974,N_15373,N_16133);
and U16975 (N_16975,N_16231,N_16043);
or U16976 (N_16976,N_15181,N_15649);
nor U16977 (N_16977,N_16067,N_15165);
xor U16978 (N_16978,N_15654,N_15264);
and U16979 (N_16979,N_15302,N_15021);
nor U16980 (N_16980,N_15624,N_16435);
xor U16981 (N_16981,N_15122,N_15435);
and U16982 (N_16982,N_15383,N_15379);
nand U16983 (N_16983,N_16283,N_16390);
or U16984 (N_16984,N_15918,N_15323);
nor U16985 (N_16985,N_15070,N_16074);
nand U16986 (N_16986,N_15759,N_16095);
or U16987 (N_16987,N_15960,N_15714);
and U16988 (N_16988,N_15096,N_15694);
nand U16989 (N_16989,N_15314,N_15945);
and U16990 (N_16990,N_15254,N_16039);
or U16991 (N_16991,N_15024,N_15239);
nor U16992 (N_16992,N_16351,N_15058);
or U16993 (N_16993,N_15491,N_15554);
or U16994 (N_16994,N_15516,N_15665);
and U16995 (N_16995,N_15916,N_15883);
nand U16996 (N_16996,N_16224,N_15687);
or U16997 (N_16997,N_15890,N_15850);
nand U16998 (N_16998,N_15453,N_15794);
nor U16999 (N_16999,N_15591,N_15235);
xnor U17000 (N_17000,N_15733,N_15430);
nor U17001 (N_17001,N_15801,N_15064);
and U17002 (N_17002,N_16395,N_15126);
and U17003 (N_17003,N_16014,N_15384);
and U17004 (N_17004,N_15480,N_15523);
nand U17005 (N_17005,N_15069,N_16325);
and U17006 (N_17006,N_15258,N_16228);
and U17007 (N_17007,N_16456,N_16171);
nor U17008 (N_17008,N_15015,N_15617);
or U17009 (N_17009,N_16143,N_15011);
or U17010 (N_17010,N_15970,N_15124);
nor U17011 (N_17011,N_15348,N_16210);
or U17012 (N_17012,N_16011,N_16150);
nor U17013 (N_17013,N_15200,N_15563);
nand U17014 (N_17014,N_15259,N_15506);
nand U17015 (N_17015,N_15448,N_16363);
or U17016 (N_17016,N_15400,N_15065);
and U17017 (N_17017,N_15777,N_16124);
or U17018 (N_17018,N_15051,N_16223);
and U17019 (N_17019,N_15858,N_16194);
nand U17020 (N_17020,N_16178,N_16305);
nor U17021 (N_17021,N_15940,N_15007);
or U17022 (N_17022,N_16182,N_16230);
nor U17023 (N_17023,N_15528,N_16168);
or U17024 (N_17024,N_15597,N_15026);
or U17025 (N_17025,N_16060,N_15899);
and U17026 (N_17026,N_15702,N_15009);
and U17027 (N_17027,N_16387,N_15274);
nor U17028 (N_17028,N_15237,N_15315);
and U17029 (N_17029,N_15103,N_16270);
nor U17030 (N_17030,N_15416,N_16172);
or U17031 (N_17031,N_15718,N_16487);
nand U17032 (N_17032,N_16422,N_15586);
or U17033 (N_17033,N_16170,N_15991);
and U17034 (N_17034,N_16370,N_15728);
and U17035 (N_17035,N_15748,N_15190);
nand U17036 (N_17036,N_16412,N_16045);
nor U17037 (N_17037,N_15756,N_15995);
nor U17038 (N_17038,N_15090,N_16026);
xnor U17039 (N_17039,N_15060,N_16383);
nor U17040 (N_17040,N_16463,N_15004);
xnor U17041 (N_17041,N_16167,N_15027);
and U17042 (N_17042,N_15160,N_15495);
nand U17043 (N_17043,N_15409,N_16245);
and U17044 (N_17044,N_15210,N_15244);
nor U17045 (N_17045,N_16093,N_16068);
or U17046 (N_17046,N_15703,N_15784);
nor U17047 (N_17047,N_15736,N_16410);
nor U17048 (N_17048,N_15447,N_15386);
nand U17049 (N_17049,N_16293,N_15252);
and U17050 (N_17050,N_15938,N_16296);
nor U17051 (N_17051,N_16103,N_15782);
nor U17052 (N_17052,N_15631,N_16378);
nand U17053 (N_17053,N_15228,N_15898);
or U17054 (N_17054,N_15044,N_15607);
nand U17055 (N_17055,N_15281,N_15788);
xor U17056 (N_17056,N_16226,N_16474);
xnor U17057 (N_17057,N_15017,N_16365);
nand U17058 (N_17058,N_15055,N_16419);
nand U17059 (N_17059,N_15600,N_15311);
xor U17060 (N_17060,N_15304,N_15825);
nand U17061 (N_17061,N_15100,N_16096);
nand U17062 (N_17062,N_15454,N_16477);
or U17063 (N_17063,N_16220,N_16404);
or U17064 (N_17064,N_16105,N_15091);
xor U17065 (N_17065,N_15550,N_15050);
xnor U17066 (N_17066,N_16450,N_15358);
nor U17067 (N_17067,N_16252,N_16491);
nand U17068 (N_17068,N_15499,N_15775);
or U17069 (N_17069,N_16056,N_16057);
nand U17070 (N_17070,N_15806,N_15712);
and U17071 (N_17071,N_15078,N_16163);
and U17072 (N_17072,N_15498,N_16441);
or U17073 (N_17073,N_15087,N_16104);
or U17074 (N_17074,N_15425,N_15719);
xor U17075 (N_17075,N_15613,N_15068);
and U17076 (N_17076,N_16071,N_16115);
xnor U17077 (N_17077,N_15161,N_15818);
xnor U17078 (N_17078,N_15265,N_15565);
nor U17079 (N_17079,N_16353,N_15471);
nand U17080 (N_17080,N_16313,N_15098);
xnor U17081 (N_17081,N_15977,N_16432);
or U17082 (N_17082,N_16101,N_16281);
nand U17083 (N_17083,N_15912,N_16138);
nor U17084 (N_17084,N_16457,N_16267);
xnor U17085 (N_17085,N_15877,N_16013);
and U17086 (N_17086,N_15633,N_15272);
or U17087 (N_17087,N_15035,N_16319);
nand U17088 (N_17088,N_15423,N_15575);
and U17089 (N_17089,N_15342,N_15541);
or U17090 (N_17090,N_15136,N_15162);
and U17091 (N_17091,N_16409,N_15681);
nand U17092 (N_17092,N_15961,N_15740);
and U17093 (N_17093,N_15285,N_15840);
xor U17094 (N_17094,N_15873,N_15390);
or U17095 (N_17095,N_15293,N_15211);
and U17096 (N_17096,N_16385,N_15072);
nand U17097 (N_17097,N_15240,N_15623);
or U17098 (N_17098,N_15783,N_16149);
nor U17099 (N_17099,N_15601,N_15692);
and U17100 (N_17100,N_16050,N_16465);
nor U17101 (N_17101,N_16352,N_16486);
or U17102 (N_17102,N_16315,N_15625);
or U17103 (N_17103,N_16258,N_15910);
and U17104 (N_17104,N_15869,N_15704);
or U17105 (N_17105,N_15746,N_15829);
or U17106 (N_17106,N_16375,N_15469);
xor U17107 (N_17107,N_16019,N_16227);
and U17108 (N_17108,N_16360,N_15786);
nor U17109 (N_17109,N_15612,N_15421);
and U17110 (N_17110,N_15295,N_15992);
nand U17111 (N_17111,N_16041,N_16264);
and U17112 (N_17112,N_16350,N_16436);
or U17113 (N_17113,N_16326,N_15914);
nor U17114 (N_17114,N_15297,N_15530);
nand U17115 (N_17115,N_15856,N_16304);
and U17116 (N_17116,N_16481,N_16247);
or U17117 (N_17117,N_16214,N_16388);
and U17118 (N_17118,N_15118,N_16451);
nor U17119 (N_17119,N_15988,N_16413);
nand U17120 (N_17120,N_15653,N_16028);
xor U17121 (N_17121,N_15932,N_15120);
nor U17122 (N_17122,N_15263,N_16467);
and U17123 (N_17123,N_15067,N_16485);
and U17124 (N_17124,N_15963,N_15352);
or U17125 (N_17125,N_16204,N_16261);
nor U17126 (N_17126,N_15525,N_16109);
and U17127 (N_17127,N_15996,N_15365);
nand U17128 (N_17128,N_16380,N_16065);
and U17129 (N_17129,N_16078,N_15309);
xor U17130 (N_17130,N_15139,N_15861);
or U17131 (N_17131,N_15630,N_15422);
or U17132 (N_17132,N_15461,N_15114);
nor U17133 (N_17133,N_15434,N_15627);
nor U17134 (N_17134,N_15484,N_15176);
or U17135 (N_17135,N_16198,N_16084);
xor U17136 (N_17136,N_16185,N_16324);
nand U17137 (N_17137,N_15226,N_15399);
nor U17138 (N_17138,N_16008,N_15751);
nor U17139 (N_17139,N_15950,N_15915);
and U17140 (N_17140,N_15412,N_15852);
nor U17141 (N_17141,N_15820,N_15810);
or U17142 (N_17142,N_15143,N_15189);
and U17143 (N_17143,N_15701,N_15183);
xnor U17144 (N_17144,N_16173,N_15609);
and U17145 (N_17145,N_16373,N_15951);
xor U17146 (N_17146,N_16376,N_15605);
xnor U17147 (N_17147,N_15086,N_15164);
nor U17148 (N_17148,N_15047,N_15520);
or U17149 (N_17149,N_15863,N_15561);
nand U17150 (N_17150,N_15147,N_15173);
xnor U17151 (N_17151,N_15222,N_15507);
nand U17152 (N_17152,N_15504,N_15230);
xor U17153 (N_17153,N_15819,N_15260);
xor U17154 (N_17154,N_15797,N_16424);
or U17155 (N_17155,N_16140,N_15301);
xor U17156 (N_17156,N_16203,N_16478);
xnor U17157 (N_17157,N_15031,N_16329);
or U17158 (N_17158,N_16389,N_15406);
and U17159 (N_17159,N_16415,N_15833);
and U17160 (N_17160,N_15032,N_15622);
nand U17161 (N_17161,N_15524,N_16144);
nand U17162 (N_17162,N_15142,N_15971);
xor U17163 (N_17163,N_15619,N_15844);
nand U17164 (N_17164,N_16453,N_16308);
xor U17165 (N_17165,N_16235,N_15594);
nor U17166 (N_17166,N_15129,N_15646);
and U17167 (N_17167,N_16122,N_15807);
and U17168 (N_17168,N_15677,N_15268);
nor U17169 (N_17169,N_16099,N_15112);
nand U17170 (N_17170,N_15371,N_15973);
or U17171 (N_17171,N_15795,N_15847);
or U17172 (N_17172,N_15002,N_16146);
xnor U17173 (N_17173,N_15500,N_16184);
and U17174 (N_17174,N_15514,N_15647);
nor U17175 (N_17175,N_15417,N_15606);
nor U17176 (N_17176,N_16121,N_15540);
nand U17177 (N_17177,N_15095,N_15768);
and U17178 (N_17178,N_15900,N_15168);
and U17179 (N_17179,N_15796,N_16128);
or U17180 (N_17180,N_15684,N_16136);
and U17181 (N_17181,N_16251,N_15835);
nand U17182 (N_17182,N_16265,N_16490);
nand U17183 (N_17183,N_16059,N_15045);
nand U17184 (N_17184,N_16190,N_16044);
xnor U17185 (N_17185,N_15195,N_15462);
nand U17186 (N_17186,N_15395,N_15564);
or U17187 (N_17187,N_15292,N_15463);
nand U17188 (N_17188,N_15404,N_15557);
and U17189 (N_17189,N_16003,N_15698);
or U17190 (N_17190,N_15792,N_16461);
nor U17191 (N_17191,N_15115,N_15097);
and U17192 (N_17192,N_15548,N_15267);
or U17193 (N_17193,N_15249,N_15559);
or U17194 (N_17194,N_15713,N_15760);
xor U17195 (N_17195,N_15312,N_16417);
nor U17196 (N_17196,N_15732,N_16396);
xor U17197 (N_17197,N_16255,N_15793);
nor U17198 (N_17198,N_16259,N_15640);
nand U17199 (N_17199,N_15433,N_16488);
xnor U17200 (N_17200,N_16018,N_15826);
xnor U17201 (N_17201,N_16175,N_16369);
and U17202 (N_17202,N_16386,N_16125);
nand U17203 (N_17203,N_15892,N_16349);
and U17204 (N_17204,N_16482,N_16196);
nor U17205 (N_17205,N_15111,N_16394);
or U17206 (N_17206,N_15381,N_15056);
and U17207 (N_17207,N_16216,N_16341);
nand U17208 (N_17208,N_15750,N_15102);
nor U17209 (N_17209,N_16029,N_15137);
or U17210 (N_17210,N_15052,N_15696);
xnor U17211 (N_17211,N_15841,N_15290);
xor U17212 (N_17212,N_15571,N_15766);
or U17213 (N_17213,N_15427,N_15410);
and U17214 (N_17214,N_16066,N_15037);
xor U17215 (N_17215,N_15428,N_16155);
or U17216 (N_17216,N_15682,N_15043);
or U17217 (N_17217,N_15983,N_16342);
nand U17218 (N_17218,N_15815,N_15339);
or U17219 (N_17219,N_16187,N_15763);
and U17220 (N_17220,N_15668,N_15799);
xor U17221 (N_17221,N_15241,N_15747);
and U17222 (N_17222,N_16497,N_16271);
nor U17223 (N_17223,N_16186,N_15689);
or U17224 (N_17224,N_15279,N_15402);
xor U17225 (N_17225,N_15148,N_15104);
nor U17226 (N_17226,N_15774,N_15328);
xor U17227 (N_17227,N_15979,N_15141);
and U17228 (N_17228,N_15257,N_16181);
nor U17229 (N_17229,N_16075,N_16098);
xnor U17230 (N_17230,N_15213,N_15549);
nor U17231 (N_17231,N_16362,N_16237);
nor U17232 (N_17232,N_15457,N_15725);
xor U17233 (N_17233,N_15638,N_15014);
or U17234 (N_17234,N_15904,N_15849);
nor U17235 (N_17235,N_15361,N_16309);
or U17236 (N_17236,N_15730,N_15894);
nand U17237 (N_17237,N_15245,N_15159);
nor U17238 (N_17238,N_16310,N_15734);
xor U17239 (N_17239,N_15271,N_15208);
nand U17240 (N_17240,N_16449,N_15053);
nor U17241 (N_17241,N_15537,N_15648);
or U17242 (N_17242,N_15707,N_16472);
xor U17243 (N_17243,N_15360,N_15277);
nor U17244 (N_17244,N_16177,N_15038);
xor U17245 (N_17245,N_15901,N_15827);
or U17246 (N_17246,N_15125,N_15911);
xnor U17247 (N_17247,N_15191,N_15927);
nor U17248 (N_17248,N_15854,N_15657);
and U17249 (N_17249,N_16433,N_15791);
nand U17250 (N_17250,N_15954,N_15383);
or U17251 (N_17251,N_16070,N_15829);
and U17252 (N_17252,N_15449,N_16304);
or U17253 (N_17253,N_15172,N_15358);
and U17254 (N_17254,N_16338,N_15166);
and U17255 (N_17255,N_15730,N_16084);
and U17256 (N_17256,N_16394,N_16291);
or U17257 (N_17257,N_15003,N_15024);
nor U17258 (N_17258,N_15545,N_15664);
nor U17259 (N_17259,N_15829,N_15784);
nor U17260 (N_17260,N_15108,N_15495);
and U17261 (N_17261,N_15396,N_16421);
or U17262 (N_17262,N_15314,N_16136);
and U17263 (N_17263,N_15616,N_15644);
or U17264 (N_17264,N_15110,N_16337);
nor U17265 (N_17265,N_15390,N_15062);
or U17266 (N_17266,N_15977,N_15576);
nor U17267 (N_17267,N_16294,N_15098);
nor U17268 (N_17268,N_16073,N_16378);
or U17269 (N_17269,N_15220,N_16211);
and U17270 (N_17270,N_15110,N_16399);
xnor U17271 (N_17271,N_15566,N_16431);
and U17272 (N_17272,N_15701,N_15203);
nor U17273 (N_17273,N_15148,N_15081);
and U17274 (N_17274,N_16083,N_15920);
nand U17275 (N_17275,N_15949,N_16244);
and U17276 (N_17276,N_15802,N_15097);
xnor U17277 (N_17277,N_15858,N_16315);
and U17278 (N_17278,N_15174,N_15391);
or U17279 (N_17279,N_15438,N_15799);
nand U17280 (N_17280,N_15833,N_15502);
or U17281 (N_17281,N_15741,N_15207);
nor U17282 (N_17282,N_16275,N_15202);
xnor U17283 (N_17283,N_15776,N_16332);
nor U17284 (N_17284,N_15746,N_16376);
or U17285 (N_17285,N_15892,N_16300);
nor U17286 (N_17286,N_15077,N_15201);
xnor U17287 (N_17287,N_15013,N_15012);
nand U17288 (N_17288,N_15448,N_16468);
xnor U17289 (N_17289,N_15979,N_15252);
nor U17290 (N_17290,N_15729,N_15232);
or U17291 (N_17291,N_15947,N_15203);
or U17292 (N_17292,N_16117,N_16243);
nor U17293 (N_17293,N_15587,N_15284);
nor U17294 (N_17294,N_15056,N_16279);
or U17295 (N_17295,N_15270,N_15027);
and U17296 (N_17296,N_16325,N_15679);
xnor U17297 (N_17297,N_15668,N_15524);
and U17298 (N_17298,N_16313,N_15288);
nand U17299 (N_17299,N_16339,N_16193);
or U17300 (N_17300,N_15655,N_15880);
or U17301 (N_17301,N_15186,N_15992);
nand U17302 (N_17302,N_15912,N_15368);
nor U17303 (N_17303,N_16338,N_15161);
xor U17304 (N_17304,N_15402,N_15400);
and U17305 (N_17305,N_16138,N_15755);
nand U17306 (N_17306,N_16070,N_15608);
and U17307 (N_17307,N_16193,N_16471);
nand U17308 (N_17308,N_16000,N_16316);
xor U17309 (N_17309,N_16170,N_15510);
xor U17310 (N_17310,N_16104,N_15827);
or U17311 (N_17311,N_15200,N_15765);
nand U17312 (N_17312,N_16193,N_16156);
nand U17313 (N_17313,N_16057,N_15002);
xor U17314 (N_17314,N_16012,N_15592);
and U17315 (N_17315,N_16324,N_15155);
nand U17316 (N_17316,N_16022,N_16493);
and U17317 (N_17317,N_16146,N_15788);
nor U17318 (N_17318,N_15927,N_15432);
or U17319 (N_17319,N_15543,N_16012);
nor U17320 (N_17320,N_16301,N_16385);
and U17321 (N_17321,N_15737,N_16348);
nor U17322 (N_17322,N_15462,N_16090);
nor U17323 (N_17323,N_16135,N_15105);
and U17324 (N_17324,N_15982,N_15901);
nand U17325 (N_17325,N_16377,N_15182);
xnor U17326 (N_17326,N_16260,N_15949);
and U17327 (N_17327,N_15365,N_16470);
or U17328 (N_17328,N_15521,N_16261);
xnor U17329 (N_17329,N_15028,N_15471);
or U17330 (N_17330,N_16190,N_15935);
xor U17331 (N_17331,N_16265,N_15438);
and U17332 (N_17332,N_15272,N_16228);
nand U17333 (N_17333,N_15892,N_16004);
xor U17334 (N_17334,N_15922,N_15591);
xor U17335 (N_17335,N_15122,N_15603);
and U17336 (N_17336,N_16272,N_15976);
and U17337 (N_17337,N_15333,N_15457);
nand U17338 (N_17338,N_15200,N_15727);
and U17339 (N_17339,N_16276,N_15725);
xor U17340 (N_17340,N_15634,N_16262);
nor U17341 (N_17341,N_16441,N_16306);
nand U17342 (N_17342,N_15956,N_15580);
xor U17343 (N_17343,N_15607,N_15144);
or U17344 (N_17344,N_16491,N_15937);
nand U17345 (N_17345,N_15685,N_16203);
nor U17346 (N_17346,N_15268,N_15021);
xnor U17347 (N_17347,N_15737,N_15615);
nor U17348 (N_17348,N_15939,N_15707);
and U17349 (N_17349,N_16101,N_15878);
or U17350 (N_17350,N_15082,N_16133);
nor U17351 (N_17351,N_16321,N_15400);
and U17352 (N_17352,N_16443,N_15066);
nor U17353 (N_17353,N_15993,N_15633);
xor U17354 (N_17354,N_15111,N_15054);
nand U17355 (N_17355,N_15839,N_16003);
and U17356 (N_17356,N_16453,N_16229);
or U17357 (N_17357,N_15734,N_15095);
nand U17358 (N_17358,N_16269,N_15106);
nor U17359 (N_17359,N_15210,N_16365);
nand U17360 (N_17360,N_15635,N_16246);
nor U17361 (N_17361,N_15575,N_16029);
nor U17362 (N_17362,N_15395,N_16464);
or U17363 (N_17363,N_16177,N_15006);
nand U17364 (N_17364,N_15790,N_15647);
and U17365 (N_17365,N_15293,N_16446);
or U17366 (N_17366,N_16456,N_15424);
nand U17367 (N_17367,N_16025,N_15802);
and U17368 (N_17368,N_15563,N_15628);
xnor U17369 (N_17369,N_15665,N_15769);
xnor U17370 (N_17370,N_15757,N_15957);
or U17371 (N_17371,N_15706,N_16295);
nand U17372 (N_17372,N_15869,N_15845);
xnor U17373 (N_17373,N_15337,N_15587);
xnor U17374 (N_17374,N_15171,N_15774);
nor U17375 (N_17375,N_15660,N_15520);
nor U17376 (N_17376,N_15238,N_15215);
and U17377 (N_17377,N_15828,N_16190);
xor U17378 (N_17378,N_15224,N_15177);
nand U17379 (N_17379,N_15371,N_15481);
nor U17380 (N_17380,N_16057,N_15875);
or U17381 (N_17381,N_15474,N_16050);
xnor U17382 (N_17382,N_15238,N_15965);
nor U17383 (N_17383,N_15323,N_15917);
or U17384 (N_17384,N_15625,N_15844);
xnor U17385 (N_17385,N_16472,N_15957);
nor U17386 (N_17386,N_15404,N_16368);
or U17387 (N_17387,N_15425,N_15809);
or U17388 (N_17388,N_16486,N_15438);
nand U17389 (N_17389,N_15444,N_15078);
or U17390 (N_17390,N_15482,N_15456);
or U17391 (N_17391,N_15773,N_15059);
or U17392 (N_17392,N_15061,N_15494);
nor U17393 (N_17393,N_15511,N_15189);
and U17394 (N_17394,N_15837,N_16388);
xnor U17395 (N_17395,N_15364,N_15682);
or U17396 (N_17396,N_16092,N_16376);
xnor U17397 (N_17397,N_15346,N_16491);
and U17398 (N_17398,N_16305,N_15545);
and U17399 (N_17399,N_15694,N_15835);
or U17400 (N_17400,N_15557,N_15730);
and U17401 (N_17401,N_15945,N_16481);
nand U17402 (N_17402,N_15952,N_15620);
xor U17403 (N_17403,N_16289,N_15532);
and U17404 (N_17404,N_15547,N_16449);
and U17405 (N_17405,N_15883,N_16186);
nor U17406 (N_17406,N_15704,N_16431);
or U17407 (N_17407,N_15738,N_15080);
nand U17408 (N_17408,N_15647,N_15159);
xor U17409 (N_17409,N_16165,N_15200);
nor U17410 (N_17410,N_15965,N_15444);
nor U17411 (N_17411,N_16313,N_15585);
or U17412 (N_17412,N_16044,N_15196);
nor U17413 (N_17413,N_15770,N_16011);
nand U17414 (N_17414,N_16282,N_16412);
or U17415 (N_17415,N_16246,N_16133);
and U17416 (N_17416,N_15060,N_15071);
xnor U17417 (N_17417,N_15219,N_16481);
xnor U17418 (N_17418,N_16136,N_16386);
nand U17419 (N_17419,N_16228,N_16327);
and U17420 (N_17420,N_15574,N_16294);
nor U17421 (N_17421,N_15115,N_16241);
nand U17422 (N_17422,N_16303,N_15952);
and U17423 (N_17423,N_15204,N_15292);
nand U17424 (N_17424,N_15863,N_15491);
and U17425 (N_17425,N_16163,N_16139);
nor U17426 (N_17426,N_15472,N_16174);
and U17427 (N_17427,N_16213,N_16405);
xor U17428 (N_17428,N_15475,N_15798);
nand U17429 (N_17429,N_15386,N_16130);
xor U17430 (N_17430,N_15263,N_15397);
or U17431 (N_17431,N_15557,N_15972);
xor U17432 (N_17432,N_15082,N_15591);
or U17433 (N_17433,N_15187,N_16074);
xnor U17434 (N_17434,N_16238,N_15519);
or U17435 (N_17435,N_15578,N_15927);
nor U17436 (N_17436,N_16281,N_15473);
and U17437 (N_17437,N_15459,N_15022);
xor U17438 (N_17438,N_15795,N_15020);
or U17439 (N_17439,N_15632,N_15614);
nor U17440 (N_17440,N_16068,N_16278);
or U17441 (N_17441,N_16199,N_15845);
nand U17442 (N_17442,N_16414,N_16005);
nand U17443 (N_17443,N_15499,N_15047);
xor U17444 (N_17444,N_15748,N_15000);
nand U17445 (N_17445,N_15270,N_15058);
and U17446 (N_17446,N_15478,N_15491);
or U17447 (N_17447,N_15175,N_16400);
nand U17448 (N_17448,N_15781,N_16457);
and U17449 (N_17449,N_16468,N_15266);
nand U17450 (N_17450,N_16317,N_15824);
and U17451 (N_17451,N_16401,N_16415);
and U17452 (N_17452,N_15887,N_15938);
or U17453 (N_17453,N_16166,N_16389);
or U17454 (N_17454,N_16438,N_16375);
nand U17455 (N_17455,N_15334,N_15793);
nor U17456 (N_17456,N_16199,N_16339);
xor U17457 (N_17457,N_15413,N_15974);
nand U17458 (N_17458,N_16149,N_15211);
and U17459 (N_17459,N_16340,N_15305);
xnor U17460 (N_17460,N_15955,N_15397);
nor U17461 (N_17461,N_15129,N_16353);
nor U17462 (N_17462,N_15417,N_15197);
xor U17463 (N_17463,N_15696,N_15470);
or U17464 (N_17464,N_16018,N_15605);
xnor U17465 (N_17465,N_16275,N_15771);
nor U17466 (N_17466,N_15269,N_16016);
or U17467 (N_17467,N_15017,N_16138);
and U17468 (N_17468,N_15250,N_15934);
or U17469 (N_17469,N_16022,N_15328);
nand U17470 (N_17470,N_15033,N_16400);
or U17471 (N_17471,N_15369,N_15054);
or U17472 (N_17472,N_15539,N_16468);
nor U17473 (N_17473,N_16150,N_15721);
or U17474 (N_17474,N_16247,N_15024);
nor U17475 (N_17475,N_15020,N_16434);
xor U17476 (N_17476,N_15634,N_15172);
or U17477 (N_17477,N_16011,N_16126);
xor U17478 (N_17478,N_15285,N_15429);
xor U17479 (N_17479,N_16081,N_15466);
xor U17480 (N_17480,N_16499,N_15400);
xnor U17481 (N_17481,N_16465,N_15341);
nor U17482 (N_17482,N_15308,N_16222);
or U17483 (N_17483,N_15309,N_16284);
nor U17484 (N_17484,N_15948,N_16087);
or U17485 (N_17485,N_15593,N_15338);
nor U17486 (N_17486,N_16005,N_15977);
or U17487 (N_17487,N_16149,N_16202);
nand U17488 (N_17488,N_15000,N_15227);
nand U17489 (N_17489,N_15241,N_15683);
nor U17490 (N_17490,N_15735,N_15687);
and U17491 (N_17491,N_16240,N_15245);
and U17492 (N_17492,N_16483,N_15006);
nand U17493 (N_17493,N_15248,N_15076);
xnor U17494 (N_17494,N_16035,N_15402);
nor U17495 (N_17495,N_15389,N_15904);
and U17496 (N_17496,N_15114,N_16316);
or U17497 (N_17497,N_16305,N_15789);
and U17498 (N_17498,N_15490,N_16219);
xor U17499 (N_17499,N_16132,N_16293);
and U17500 (N_17500,N_15249,N_16261);
nor U17501 (N_17501,N_16156,N_15517);
nor U17502 (N_17502,N_15110,N_15528);
and U17503 (N_17503,N_15355,N_16191);
nor U17504 (N_17504,N_15430,N_15524);
xor U17505 (N_17505,N_15003,N_15645);
or U17506 (N_17506,N_15833,N_16151);
xor U17507 (N_17507,N_15325,N_15433);
xor U17508 (N_17508,N_15965,N_15548);
xor U17509 (N_17509,N_16104,N_15762);
or U17510 (N_17510,N_16411,N_16073);
or U17511 (N_17511,N_16167,N_16074);
or U17512 (N_17512,N_15811,N_16423);
nand U17513 (N_17513,N_16234,N_16370);
nor U17514 (N_17514,N_16320,N_16102);
nor U17515 (N_17515,N_16043,N_15084);
or U17516 (N_17516,N_15754,N_16074);
xor U17517 (N_17517,N_16448,N_16471);
xor U17518 (N_17518,N_15685,N_15069);
or U17519 (N_17519,N_15270,N_16048);
and U17520 (N_17520,N_15220,N_16366);
or U17521 (N_17521,N_16472,N_16473);
xor U17522 (N_17522,N_15079,N_16334);
nand U17523 (N_17523,N_15236,N_16132);
or U17524 (N_17524,N_15522,N_15629);
and U17525 (N_17525,N_15392,N_15000);
or U17526 (N_17526,N_16245,N_16066);
nor U17527 (N_17527,N_15405,N_15406);
or U17528 (N_17528,N_15108,N_16033);
and U17529 (N_17529,N_16306,N_15178);
nor U17530 (N_17530,N_16138,N_16108);
nand U17531 (N_17531,N_16198,N_15209);
nand U17532 (N_17532,N_15226,N_15625);
nor U17533 (N_17533,N_15368,N_16009);
or U17534 (N_17534,N_15460,N_15272);
nand U17535 (N_17535,N_16400,N_15576);
or U17536 (N_17536,N_15154,N_16272);
nand U17537 (N_17537,N_15777,N_16181);
xnor U17538 (N_17538,N_15634,N_15660);
nand U17539 (N_17539,N_16185,N_16189);
or U17540 (N_17540,N_15616,N_15272);
xnor U17541 (N_17541,N_16436,N_16198);
nor U17542 (N_17542,N_15795,N_15186);
or U17543 (N_17543,N_16038,N_16143);
nor U17544 (N_17544,N_16311,N_15955);
or U17545 (N_17545,N_15836,N_15473);
xor U17546 (N_17546,N_15947,N_15341);
or U17547 (N_17547,N_15826,N_15079);
and U17548 (N_17548,N_16268,N_15518);
xor U17549 (N_17549,N_15398,N_15537);
nand U17550 (N_17550,N_15909,N_16297);
nand U17551 (N_17551,N_15822,N_15110);
or U17552 (N_17552,N_15644,N_16410);
nor U17553 (N_17553,N_15837,N_15836);
or U17554 (N_17554,N_15438,N_15921);
nand U17555 (N_17555,N_16305,N_15018);
and U17556 (N_17556,N_15827,N_16373);
or U17557 (N_17557,N_15260,N_15299);
nor U17558 (N_17558,N_16203,N_15741);
nand U17559 (N_17559,N_16137,N_15622);
nor U17560 (N_17560,N_15624,N_15203);
nand U17561 (N_17561,N_15927,N_16285);
nor U17562 (N_17562,N_16148,N_15689);
and U17563 (N_17563,N_15222,N_16111);
nand U17564 (N_17564,N_15061,N_16352);
or U17565 (N_17565,N_16474,N_15987);
nor U17566 (N_17566,N_15981,N_15964);
nand U17567 (N_17567,N_15556,N_15494);
nand U17568 (N_17568,N_15200,N_15814);
or U17569 (N_17569,N_15384,N_15205);
and U17570 (N_17570,N_16078,N_15084);
and U17571 (N_17571,N_16433,N_15654);
xnor U17572 (N_17572,N_16430,N_15668);
nand U17573 (N_17573,N_16163,N_16187);
and U17574 (N_17574,N_16149,N_15391);
and U17575 (N_17575,N_15314,N_15675);
nand U17576 (N_17576,N_15936,N_15152);
nor U17577 (N_17577,N_15022,N_15354);
and U17578 (N_17578,N_15856,N_15408);
xor U17579 (N_17579,N_15229,N_16021);
and U17580 (N_17580,N_15772,N_15843);
and U17581 (N_17581,N_16277,N_15999);
xnor U17582 (N_17582,N_16052,N_15791);
xnor U17583 (N_17583,N_15582,N_15101);
nor U17584 (N_17584,N_15981,N_15650);
xor U17585 (N_17585,N_15929,N_15408);
and U17586 (N_17586,N_16034,N_15818);
nor U17587 (N_17587,N_16057,N_16450);
and U17588 (N_17588,N_16415,N_15931);
nor U17589 (N_17589,N_16158,N_15478);
nand U17590 (N_17590,N_15723,N_15474);
xor U17591 (N_17591,N_15518,N_16301);
nor U17592 (N_17592,N_16349,N_15435);
or U17593 (N_17593,N_15868,N_15815);
nor U17594 (N_17594,N_16383,N_16147);
nor U17595 (N_17595,N_15301,N_15664);
nand U17596 (N_17596,N_16338,N_16319);
nand U17597 (N_17597,N_15047,N_15096);
or U17598 (N_17598,N_15534,N_16403);
nor U17599 (N_17599,N_15511,N_16211);
nor U17600 (N_17600,N_16026,N_15341);
and U17601 (N_17601,N_15267,N_15147);
nand U17602 (N_17602,N_15855,N_16487);
or U17603 (N_17603,N_15115,N_16079);
nand U17604 (N_17604,N_16497,N_15898);
xnor U17605 (N_17605,N_16253,N_16029);
xnor U17606 (N_17606,N_15265,N_15193);
nand U17607 (N_17607,N_15407,N_15713);
or U17608 (N_17608,N_16490,N_15551);
nor U17609 (N_17609,N_15420,N_16194);
or U17610 (N_17610,N_15868,N_16217);
nor U17611 (N_17611,N_16181,N_16175);
nor U17612 (N_17612,N_15007,N_15998);
xnor U17613 (N_17613,N_15797,N_16251);
and U17614 (N_17614,N_15468,N_15126);
or U17615 (N_17615,N_16300,N_15125);
and U17616 (N_17616,N_16057,N_15082);
nor U17617 (N_17617,N_15075,N_15870);
xor U17618 (N_17618,N_16490,N_16277);
or U17619 (N_17619,N_15968,N_15168);
xor U17620 (N_17620,N_16237,N_16111);
nor U17621 (N_17621,N_15435,N_15018);
nand U17622 (N_17622,N_15713,N_15654);
nand U17623 (N_17623,N_15021,N_15134);
nor U17624 (N_17624,N_16357,N_15795);
and U17625 (N_17625,N_15678,N_15685);
xnor U17626 (N_17626,N_15475,N_16175);
nand U17627 (N_17627,N_16132,N_16324);
and U17628 (N_17628,N_15196,N_16472);
nand U17629 (N_17629,N_15894,N_15351);
nor U17630 (N_17630,N_15270,N_15169);
or U17631 (N_17631,N_15879,N_16475);
xnor U17632 (N_17632,N_15065,N_15549);
xor U17633 (N_17633,N_15486,N_15895);
and U17634 (N_17634,N_15317,N_15268);
or U17635 (N_17635,N_15281,N_15441);
xor U17636 (N_17636,N_15138,N_16020);
nand U17637 (N_17637,N_15416,N_15200);
xnor U17638 (N_17638,N_16131,N_15842);
or U17639 (N_17639,N_15872,N_15558);
xor U17640 (N_17640,N_15811,N_15235);
xnor U17641 (N_17641,N_15346,N_16061);
and U17642 (N_17642,N_15166,N_15687);
or U17643 (N_17643,N_15877,N_15925);
or U17644 (N_17644,N_16277,N_15337);
xor U17645 (N_17645,N_15174,N_15661);
nand U17646 (N_17646,N_16036,N_15686);
xor U17647 (N_17647,N_16395,N_15716);
or U17648 (N_17648,N_15337,N_15413);
nand U17649 (N_17649,N_15213,N_15795);
xnor U17650 (N_17650,N_16229,N_15657);
xnor U17651 (N_17651,N_15801,N_15825);
nand U17652 (N_17652,N_15107,N_15229);
and U17653 (N_17653,N_16367,N_15804);
nor U17654 (N_17654,N_16224,N_15467);
nor U17655 (N_17655,N_15618,N_16295);
xor U17656 (N_17656,N_15186,N_15548);
and U17657 (N_17657,N_15325,N_15851);
nor U17658 (N_17658,N_15504,N_16427);
or U17659 (N_17659,N_15539,N_15621);
nor U17660 (N_17660,N_16202,N_15915);
nor U17661 (N_17661,N_15003,N_15630);
xnor U17662 (N_17662,N_16271,N_15653);
nor U17663 (N_17663,N_15401,N_15950);
or U17664 (N_17664,N_15593,N_15126);
xor U17665 (N_17665,N_16088,N_15844);
xor U17666 (N_17666,N_16287,N_15899);
xnor U17667 (N_17667,N_16104,N_15391);
nand U17668 (N_17668,N_16219,N_16437);
and U17669 (N_17669,N_15255,N_16133);
xor U17670 (N_17670,N_16467,N_15136);
nand U17671 (N_17671,N_15850,N_16115);
or U17672 (N_17672,N_16192,N_15749);
and U17673 (N_17673,N_15431,N_15540);
nor U17674 (N_17674,N_15551,N_16034);
nor U17675 (N_17675,N_15937,N_15921);
nor U17676 (N_17676,N_16233,N_15728);
nor U17677 (N_17677,N_16442,N_15112);
xor U17678 (N_17678,N_15562,N_16094);
nor U17679 (N_17679,N_16259,N_15323);
and U17680 (N_17680,N_15461,N_15741);
or U17681 (N_17681,N_15920,N_15260);
nand U17682 (N_17682,N_15563,N_16026);
xor U17683 (N_17683,N_16159,N_16396);
or U17684 (N_17684,N_16460,N_15067);
and U17685 (N_17685,N_15405,N_15124);
xnor U17686 (N_17686,N_15628,N_16015);
or U17687 (N_17687,N_16357,N_15554);
nand U17688 (N_17688,N_16254,N_15691);
and U17689 (N_17689,N_15227,N_15753);
and U17690 (N_17690,N_15847,N_15715);
xnor U17691 (N_17691,N_16395,N_15665);
or U17692 (N_17692,N_15569,N_16061);
or U17693 (N_17693,N_15649,N_15308);
nand U17694 (N_17694,N_16349,N_15191);
and U17695 (N_17695,N_15168,N_16138);
nor U17696 (N_17696,N_16386,N_16019);
or U17697 (N_17697,N_16487,N_16187);
and U17698 (N_17698,N_15633,N_15451);
nor U17699 (N_17699,N_15722,N_16364);
or U17700 (N_17700,N_16070,N_16257);
or U17701 (N_17701,N_15454,N_15653);
nor U17702 (N_17702,N_15236,N_15949);
nor U17703 (N_17703,N_15435,N_15783);
xor U17704 (N_17704,N_15844,N_15033);
nand U17705 (N_17705,N_15420,N_15828);
or U17706 (N_17706,N_15486,N_15164);
or U17707 (N_17707,N_16162,N_15415);
xnor U17708 (N_17708,N_15747,N_15465);
or U17709 (N_17709,N_16422,N_16029);
xnor U17710 (N_17710,N_16304,N_15511);
or U17711 (N_17711,N_16049,N_15295);
nor U17712 (N_17712,N_15230,N_16422);
nor U17713 (N_17713,N_15701,N_15303);
nand U17714 (N_17714,N_15360,N_15571);
nand U17715 (N_17715,N_15533,N_15719);
xor U17716 (N_17716,N_16291,N_16205);
nor U17717 (N_17717,N_15228,N_15802);
nand U17718 (N_17718,N_16163,N_15169);
and U17719 (N_17719,N_15138,N_15946);
and U17720 (N_17720,N_15791,N_15715);
or U17721 (N_17721,N_15771,N_15513);
and U17722 (N_17722,N_15821,N_15138);
and U17723 (N_17723,N_15235,N_16163);
and U17724 (N_17724,N_16356,N_16280);
xor U17725 (N_17725,N_15553,N_15591);
nand U17726 (N_17726,N_16148,N_16200);
or U17727 (N_17727,N_15837,N_16070);
xor U17728 (N_17728,N_15400,N_16013);
or U17729 (N_17729,N_15789,N_16262);
nor U17730 (N_17730,N_16449,N_16314);
or U17731 (N_17731,N_15207,N_15610);
or U17732 (N_17732,N_15259,N_15689);
nor U17733 (N_17733,N_15569,N_15362);
nand U17734 (N_17734,N_15513,N_16299);
or U17735 (N_17735,N_15162,N_15764);
xor U17736 (N_17736,N_15068,N_15484);
xnor U17737 (N_17737,N_15337,N_15267);
and U17738 (N_17738,N_16154,N_15445);
or U17739 (N_17739,N_15263,N_15181);
or U17740 (N_17740,N_16088,N_15824);
nand U17741 (N_17741,N_15858,N_16154);
xnor U17742 (N_17742,N_15986,N_15370);
xnor U17743 (N_17743,N_15465,N_15402);
and U17744 (N_17744,N_15881,N_16478);
nand U17745 (N_17745,N_16478,N_15761);
and U17746 (N_17746,N_16044,N_15349);
nor U17747 (N_17747,N_16351,N_16156);
nand U17748 (N_17748,N_16010,N_15616);
xnor U17749 (N_17749,N_15396,N_15622);
and U17750 (N_17750,N_16040,N_15153);
or U17751 (N_17751,N_15244,N_16071);
and U17752 (N_17752,N_16476,N_15164);
or U17753 (N_17753,N_16380,N_16259);
and U17754 (N_17754,N_15470,N_15364);
nand U17755 (N_17755,N_15618,N_15077);
or U17756 (N_17756,N_16051,N_16338);
nor U17757 (N_17757,N_15190,N_15238);
nand U17758 (N_17758,N_15511,N_15463);
xnor U17759 (N_17759,N_16265,N_15595);
xor U17760 (N_17760,N_16292,N_15109);
nor U17761 (N_17761,N_15750,N_15050);
xor U17762 (N_17762,N_15572,N_16196);
nor U17763 (N_17763,N_15745,N_15710);
nor U17764 (N_17764,N_16289,N_15415);
xor U17765 (N_17765,N_16496,N_16033);
or U17766 (N_17766,N_15116,N_15221);
nor U17767 (N_17767,N_15455,N_15720);
and U17768 (N_17768,N_15655,N_16199);
or U17769 (N_17769,N_15327,N_16315);
nand U17770 (N_17770,N_15970,N_16414);
xnor U17771 (N_17771,N_15765,N_15441);
and U17772 (N_17772,N_16421,N_15885);
xor U17773 (N_17773,N_15372,N_16346);
or U17774 (N_17774,N_15004,N_16256);
xor U17775 (N_17775,N_15351,N_15181);
nand U17776 (N_17776,N_16041,N_15963);
xnor U17777 (N_17777,N_15979,N_15222);
and U17778 (N_17778,N_15429,N_15193);
nand U17779 (N_17779,N_15677,N_15295);
or U17780 (N_17780,N_15575,N_15213);
or U17781 (N_17781,N_15806,N_16101);
or U17782 (N_17782,N_15556,N_16438);
nand U17783 (N_17783,N_16264,N_15394);
nor U17784 (N_17784,N_16342,N_15928);
and U17785 (N_17785,N_16112,N_16229);
or U17786 (N_17786,N_16400,N_15766);
xor U17787 (N_17787,N_15862,N_16272);
and U17788 (N_17788,N_15566,N_16402);
or U17789 (N_17789,N_15986,N_15735);
and U17790 (N_17790,N_15549,N_15221);
xnor U17791 (N_17791,N_16014,N_15257);
and U17792 (N_17792,N_15171,N_16264);
or U17793 (N_17793,N_16098,N_16487);
xor U17794 (N_17794,N_16260,N_15289);
and U17795 (N_17795,N_15390,N_15512);
nand U17796 (N_17796,N_15260,N_16073);
or U17797 (N_17797,N_16323,N_15704);
xor U17798 (N_17798,N_16157,N_15826);
or U17799 (N_17799,N_16402,N_15086);
xor U17800 (N_17800,N_15509,N_15924);
nor U17801 (N_17801,N_15174,N_15283);
nand U17802 (N_17802,N_16367,N_15556);
or U17803 (N_17803,N_16202,N_15675);
nand U17804 (N_17804,N_15033,N_15118);
or U17805 (N_17805,N_15065,N_15498);
xor U17806 (N_17806,N_16172,N_15484);
nor U17807 (N_17807,N_15894,N_16106);
nor U17808 (N_17808,N_15352,N_16479);
or U17809 (N_17809,N_15257,N_15012);
nand U17810 (N_17810,N_16002,N_15149);
and U17811 (N_17811,N_15739,N_16026);
nand U17812 (N_17812,N_15393,N_16164);
or U17813 (N_17813,N_15267,N_16145);
and U17814 (N_17814,N_16331,N_16042);
xor U17815 (N_17815,N_15908,N_15374);
xor U17816 (N_17816,N_15275,N_15783);
and U17817 (N_17817,N_15294,N_15160);
and U17818 (N_17818,N_15420,N_15226);
nor U17819 (N_17819,N_15714,N_15827);
and U17820 (N_17820,N_15241,N_16135);
and U17821 (N_17821,N_16178,N_15836);
nand U17822 (N_17822,N_16153,N_15869);
xor U17823 (N_17823,N_16373,N_15822);
or U17824 (N_17824,N_15531,N_15234);
or U17825 (N_17825,N_15247,N_15675);
and U17826 (N_17826,N_15465,N_15421);
xor U17827 (N_17827,N_15432,N_15956);
nand U17828 (N_17828,N_16360,N_16150);
and U17829 (N_17829,N_16022,N_15725);
nor U17830 (N_17830,N_15020,N_16200);
nor U17831 (N_17831,N_15274,N_16021);
nand U17832 (N_17832,N_15366,N_15707);
nor U17833 (N_17833,N_16056,N_16296);
xor U17834 (N_17834,N_15349,N_15945);
and U17835 (N_17835,N_16101,N_15969);
nor U17836 (N_17836,N_16099,N_15581);
xnor U17837 (N_17837,N_15659,N_16441);
or U17838 (N_17838,N_15183,N_15966);
xor U17839 (N_17839,N_15133,N_15435);
xnor U17840 (N_17840,N_15741,N_15506);
or U17841 (N_17841,N_15714,N_16094);
and U17842 (N_17842,N_15780,N_15205);
and U17843 (N_17843,N_15361,N_15556);
and U17844 (N_17844,N_16092,N_16032);
nand U17845 (N_17845,N_16229,N_16143);
nor U17846 (N_17846,N_15226,N_16158);
or U17847 (N_17847,N_15470,N_15894);
nor U17848 (N_17848,N_16107,N_15667);
xnor U17849 (N_17849,N_15986,N_15279);
and U17850 (N_17850,N_15024,N_15553);
and U17851 (N_17851,N_15786,N_16182);
xor U17852 (N_17852,N_16294,N_15302);
nand U17853 (N_17853,N_15286,N_16123);
and U17854 (N_17854,N_15082,N_15648);
nor U17855 (N_17855,N_16088,N_15359);
or U17856 (N_17856,N_15511,N_16073);
or U17857 (N_17857,N_15645,N_16024);
or U17858 (N_17858,N_15360,N_16246);
and U17859 (N_17859,N_15098,N_16169);
nand U17860 (N_17860,N_15848,N_16356);
nand U17861 (N_17861,N_16088,N_16302);
or U17862 (N_17862,N_15149,N_15011);
or U17863 (N_17863,N_15823,N_16103);
nand U17864 (N_17864,N_15164,N_16291);
xor U17865 (N_17865,N_16475,N_16218);
or U17866 (N_17866,N_16413,N_15353);
or U17867 (N_17867,N_15123,N_15003);
and U17868 (N_17868,N_16117,N_15074);
or U17869 (N_17869,N_15621,N_15989);
or U17870 (N_17870,N_15899,N_15486);
and U17871 (N_17871,N_15539,N_16160);
xor U17872 (N_17872,N_15274,N_15079);
nand U17873 (N_17873,N_15357,N_16328);
xnor U17874 (N_17874,N_16382,N_16427);
nand U17875 (N_17875,N_16214,N_15233);
nand U17876 (N_17876,N_16357,N_15856);
or U17877 (N_17877,N_16442,N_15486);
nor U17878 (N_17878,N_15294,N_15402);
xor U17879 (N_17879,N_15734,N_15562);
xor U17880 (N_17880,N_15339,N_16047);
or U17881 (N_17881,N_15397,N_15571);
xor U17882 (N_17882,N_15820,N_15532);
xnor U17883 (N_17883,N_16005,N_15237);
or U17884 (N_17884,N_16021,N_15498);
xnor U17885 (N_17885,N_15993,N_15941);
nor U17886 (N_17886,N_15940,N_15656);
nand U17887 (N_17887,N_15385,N_16474);
xnor U17888 (N_17888,N_15724,N_15461);
and U17889 (N_17889,N_15207,N_16332);
nand U17890 (N_17890,N_16022,N_15243);
or U17891 (N_17891,N_15234,N_15055);
xor U17892 (N_17892,N_16265,N_15801);
or U17893 (N_17893,N_15415,N_15849);
or U17894 (N_17894,N_15257,N_16461);
or U17895 (N_17895,N_15832,N_15014);
and U17896 (N_17896,N_15800,N_16234);
nor U17897 (N_17897,N_16386,N_15420);
nand U17898 (N_17898,N_16481,N_16105);
and U17899 (N_17899,N_15201,N_16330);
nand U17900 (N_17900,N_16247,N_16296);
xor U17901 (N_17901,N_15345,N_15552);
nand U17902 (N_17902,N_16487,N_15432);
or U17903 (N_17903,N_15750,N_15853);
or U17904 (N_17904,N_15341,N_15386);
and U17905 (N_17905,N_16264,N_15918);
xor U17906 (N_17906,N_15242,N_16441);
and U17907 (N_17907,N_15679,N_15215);
xnor U17908 (N_17908,N_15903,N_15191);
xnor U17909 (N_17909,N_16183,N_15810);
or U17910 (N_17910,N_15147,N_16034);
or U17911 (N_17911,N_15021,N_16222);
or U17912 (N_17912,N_15352,N_15074);
nor U17913 (N_17913,N_15275,N_15004);
xor U17914 (N_17914,N_16166,N_15087);
nor U17915 (N_17915,N_15045,N_15439);
xnor U17916 (N_17916,N_15043,N_16122);
xnor U17917 (N_17917,N_15174,N_15611);
nand U17918 (N_17918,N_16099,N_15958);
nand U17919 (N_17919,N_16215,N_15480);
xor U17920 (N_17920,N_16117,N_15840);
nand U17921 (N_17921,N_15933,N_16090);
nand U17922 (N_17922,N_15370,N_16421);
or U17923 (N_17923,N_15863,N_15531);
nand U17924 (N_17924,N_15599,N_16087);
nand U17925 (N_17925,N_16135,N_15424);
nor U17926 (N_17926,N_15154,N_16198);
nand U17927 (N_17927,N_15535,N_15124);
or U17928 (N_17928,N_15575,N_15941);
and U17929 (N_17929,N_15423,N_16376);
xor U17930 (N_17930,N_15125,N_15376);
xnor U17931 (N_17931,N_15868,N_16264);
nor U17932 (N_17932,N_15562,N_15334);
xor U17933 (N_17933,N_15982,N_15028);
or U17934 (N_17934,N_16062,N_16002);
xnor U17935 (N_17935,N_15160,N_15037);
nor U17936 (N_17936,N_15734,N_15280);
or U17937 (N_17937,N_15184,N_16328);
xor U17938 (N_17938,N_16101,N_15877);
or U17939 (N_17939,N_15932,N_16107);
or U17940 (N_17940,N_16019,N_15879);
or U17941 (N_17941,N_15628,N_15745);
and U17942 (N_17942,N_15064,N_15672);
xor U17943 (N_17943,N_15582,N_16184);
or U17944 (N_17944,N_15357,N_16023);
nand U17945 (N_17945,N_15219,N_16245);
nor U17946 (N_17946,N_16051,N_16033);
and U17947 (N_17947,N_15888,N_15120);
xnor U17948 (N_17948,N_15811,N_15225);
or U17949 (N_17949,N_15348,N_15064);
nand U17950 (N_17950,N_16300,N_15894);
nor U17951 (N_17951,N_15203,N_16076);
nor U17952 (N_17952,N_15212,N_15211);
or U17953 (N_17953,N_15931,N_16203);
xnor U17954 (N_17954,N_15710,N_16462);
nor U17955 (N_17955,N_15084,N_15871);
nand U17956 (N_17956,N_15455,N_15866);
and U17957 (N_17957,N_16024,N_16051);
and U17958 (N_17958,N_15158,N_15278);
nor U17959 (N_17959,N_15250,N_16428);
nand U17960 (N_17960,N_15058,N_15776);
and U17961 (N_17961,N_15152,N_16446);
nand U17962 (N_17962,N_15875,N_15442);
xor U17963 (N_17963,N_15942,N_16422);
nand U17964 (N_17964,N_15493,N_15672);
nor U17965 (N_17965,N_15477,N_15523);
nand U17966 (N_17966,N_15645,N_15960);
or U17967 (N_17967,N_15858,N_15227);
and U17968 (N_17968,N_16300,N_16071);
xnor U17969 (N_17969,N_15902,N_15624);
nor U17970 (N_17970,N_15683,N_15248);
and U17971 (N_17971,N_15096,N_15679);
or U17972 (N_17972,N_15657,N_16375);
or U17973 (N_17973,N_16369,N_15495);
nor U17974 (N_17974,N_15481,N_16046);
xnor U17975 (N_17975,N_16204,N_15053);
nor U17976 (N_17976,N_15828,N_16414);
xnor U17977 (N_17977,N_15385,N_16115);
nor U17978 (N_17978,N_16083,N_15568);
xnor U17979 (N_17979,N_16400,N_15288);
xnor U17980 (N_17980,N_15403,N_15336);
xor U17981 (N_17981,N_15788,N_16229);
xor U17982 (N_17982,N_15538,N_16238);
nand U17983 (N_17983,N_16061,N_15046);
or U17984 (N_17984,N_15983,N_16359);
and U17985 (N_17985,N_16117,N_15839);
xnor U17986 (N_17986,N_16139,N_15976);
nor U17987 (N_17987,N_16490,N_15550);
nor U17988 (N_17988,N_16305,N_16182);
nand U17989 (N_17989,N_15579,N_15717);
and U17990 (N_17990,N_15774,N_15353);
nand U17991 (N_17991,N_16029,N_16308);
xnor U17992 (N_17992,N_15320,N_15074);
and U17993 (N_17993,N_15951,N_16186);
xnor U17994 (N_17994,N_15458,N_16419);
xnor U17995 (N_17995,N_15557,N_16418);
nor U17996 (N_17996,N_15988,N_16258);
and U17997 (N_17997,N_16020,N_15652);
nand U17998 (N_17998,N_15722,N_15288);
xor U17999 (N_17999,N_15297,N_15777);
xor U18000 (N_18000,N_17932,N_16560);
and U18001 (N_18001,N_16950,N_17651);
nand U18002 (N_18002,N_17196,N_17700);
and U18003 (N_18003,N_17789,N_17454);
nand U18004 (N_18004,N_17614,N_17112);
xor U18005 (N_18005,N_16531,N_17904);
nand U18006 (N_18006,N_17599,N_16627);
or U18007 (N_18007,N_17480,N_17348);
or U18008 (N_18008,N_17251,N_17858);
and U18009 (N_18009,N_16628,N_17911);
and U18010 (N_18010,N_16926,N_17177);
or U18011 (N_18011,N_16725,N_17515);
and U18012 (N_18012,N_16651,N_17520);
xnor U18013 (N_18013,N_16665,N_16849);
nand U18014 (N_18014,N_16896,N_16608);
or U18015 (N_18015,N_17108,N_16835);
and U18016 (N_18016,N_17968,N_16749);
and U18017 (N_18017,N_17323,N_16808);
nand U18018 (N_18018,N_16523,N_17568);
and U18019 (N_18019,N_17105,N_17610);
and U18020 (N_18020,N_16700,N_16895);
nand U18021 (N_18021,N_17114,N_17535);
or U18022 (N_18022,N_17688,N_16629);
nor U18023 (N_18023,N_17237,N_17181);
xnor U18024 (N_18024,N_17538,N_17376);
nand U18025 (N_18025,N_17053,N_16557);
xnor U18026 (N_18026,N_16880,N_17365);
and U18027 (N_18027,N_16988,N_16780);
nor U18028 (N_18028,N_17756,N_17748);
nand U18029 (N_18029,N_16690,N_16512);
or U18030 (N_18030,N_17987,N_16830);
nor U18031 (N_18031,N_17083,N_16980);
xnor U18032 (N_18032,N_16846,N_16589);
nand U18033 (N_18033,N_16816,N_16774);
or U18034 (N_18034,N_16652,N_17195);
and U18035 (N_18035,N_17971,N_16909);
and U18036 (N_18036,N_16504,N_16614);
xor U18037 (N_18037,N_17673,N_17357);
nand U18038 (N_18038,N_17386,N_17902);
nor U18039 (N_18039,N_16738,N_16593);
nor U18040 (N_18040,N_17206,N_16607);
nand U18041 (N_18041,N_17295,N_17256);
nand U18042 (N_18042,N_17872,N_17464);
and U18043 (N_18043,N_17328,N_17723);
and U18044 (N_18044,N_17644,N_16932);
or U18045 (N_18045,N_17032,N_17793);
and U18046 (N_18046,N_16685,N_17084);
nor U18047 (N_18047,N_16916,N_17836);
or U18048 (N_18048,N_17071,N_16555);
xnor U18049 (N_18049,N_17353,N_16852);
xnor U18050 (N_18050,N_17235,N_17578);
xnor U18051 (N_18051,N_17134,N_16992);
and U18052 (N_18052,N_16732,N_17419);
nor U18053 (N_18053,N_17097,N_17199);
xnor U18054 (N_18054,N_17269,N_17065);
and U18055 (N_18055,N_17270,N_16990);
or U18056 (N_18056,N_17524,N_17602);
xor U18057 (N_18057,N_16966,N_17895);
nand U18058 (N_18058,N_17654,N_17173);
and U18059 (N_18059,N_17178,N_16914);
xnor U18060 (N_18060,N_17989,N_17795);
nand U18061 (N_18061,N_17582,N_16847);
and U18062 (N_18062,N_16807,N_16925);
xnor U18063 (N_18063,N_16899,N_17893);
or U18064 (N_18064,N_16995,N_16977);
xor U18065 (N_18065,N_17714,N_17507);
and U18066 (N_18066,N_17119,N_16656);
or U18067 (N_18067,N_16902,N_17806);
or U18068 (N_18068,N_17660,N_17122);
xor U18069 (N_18069,N_17991,N_17068);
or U18070 (N_18070,N_17655,N_16944);
nand U18071 (N_18071,N_17819,N_16753);
nor U18072 (N_18072,N_17483,N_17788);
or U18073 (N_18073,N_16576,N_17567);
and U18074 (N_18074,N_16982,N_16919);
and U18075 (N_18075,N_17226,N_17824);
and U18076 (N_18076,N_16781,N_16859);
or U18077 (N_18077,N_17924,N_17728);
nor U18078 (N_18078,N_17208,N_16826);
nor U18079 (N_18079,N_16979,N_17049);
nand U18080 (N_18080,N_17048,N_17790);
xor U18081 (N_18081,N_17865,N_17609);
and U18082 (N_18082,N_16963,N_17772);
xor U18083 (N_18083,N_17505,N_17000);
or U18084 (N_18084,N_16953,N_17658);
or U18085 (N_18085,N_17504,N_17404);
and U18086 (N_18086,N_17549,N_17639);
nor U18087 (N_18087,N_17922,N_17211);
nor U18088 (N_18088,N_17992,N_17448);
or U18089 (N_18089,N_17413,N_16959);
and U18090 (N_18090,N_16657,N_17730);
xnor U18091 (N_18091,N_17244,N_17783);
xor U18092 (N_18092,N_17209,N_16567);
xor U18093 (N_18093,N_16720,N_17884);
and U18094 (N_18094,N_17689,N_17213);
xor U18095 (N_18095,N_17970,N_17521);
or U18096 (N_18096,N_16583,N_17290);
xor U18097 (N_18097,N_17394,N_16621);
or U18098 (N_18098,N_17111,N_16615);
xor U18099 (N_18099,N_17456,N_17947);
nor U18100 (N_18100,N_17481,N_17368);
nand U18101 (N_18101,N_17336,N_17030);
nand U18102 (N_18102,N_17337,N_17729);
xor U18103 (N_18103,N_16891,N_17476);
and U18104 (N_18104,N_17013,N_17821);
nand U18105 (N_18105,N_16778,N_17377);
and U18106 (N_18106,N_17154,N_17937);
nand U18107 (N_18107,N_17408,N_17581);
nand U18108 (N_18108,N_17741,N_17167);
xnor U18109 (N_18109,N_16693,N_16622);
or U18110 (N_18110,N_17072,N_17469);
nor U18111 (N_18111,N_17045,N_16987);
xnor U18112 (N_18112,N_16554,N_17548);
nor U18113 (N_18113,N_17558,N_16930);
nand U18114 (N_18114,N_17364,N_17636);
nand U18115 (N_18115,N_17063,N_17144);
or U18116 (N_18116,N_17038,N_16506);
nand U18117 (N_18117,N_17852,N_16955);
xor U18118 (N_18118,N_17981,N_16812);
nor U18119 (N_18119,N_17841,N_17798);
xnor U18120 (N_18120,N_17054,N_17896);
or U18121 (N_18121,N_16773,N_17215);
xnor U18122 (N_18122,N_17466,N_17274);
nor U18123 (N_18123,N_17875,N_17238);
or U18124 (N_18124,N_16864,N_17601);
nand U18125 (N_18125,N_16658,N_17052);
nand U18126 (N_18126,N_17802,N_17482);
nor U18127 (N_18127,N_17839,N_17387);
or U18128 (N_18128,N_17287,N_16514);
nand U18129 (N_18129,N_17935,N_17950);
xor U18130 (N_18130,N_17853,N_17533);
and U18131 (N_18131,N_17130,N_17489);
xnor U18132 (N_18132,N_16619,N_16716);
and U18133 (N_18133,N_16637,N_16569);
and U18134 (N_18134,N_17620,N_17585);
nand U18135 (N_18135,N_16533,N_17917);
xor U18136 (N_18136,N_16888,N_17008);
or U18137 (N_18137,N_17069,N_16522);
xor U18138 (N_18138,N_16603,N_17305);
nand U18139 (N_18139,N_16537,N_17534);
nor U18140 (N_18140,N_16655,N_17266);
and U18141 (N_18141,N_16827,N_17557);
and U18142 (N_18142,N_17358,N_16927);
and U18143 (N_18143,N_16551,N_17550);
and U18144 (N_18144,N_17418,N_16815);
xnor U18145 (N_18145,N_17869,N_17471);
nor U18146 (N_18146,N_17747,N_17960);
or U18147 (N_18147,N_17147,N_17864);
and U18148 (N_18148,N_16819,N_17951);
or U18149 (N_18149,N_17701,N_17663);
nand U18150 (N_18150,N_16636,N_17706);
or U18151 (N_18151,N_17109,N_17443);
or U18152 (N_18152,N_16737,N_17682);
or U18153 (N_18153,N_16702,N_16884);
or U18154 (N_18154,N_16735,N_17647);
nand U18155 (N_18155,N_16626,N_17145);
nand U18156 (N_18156,N_16724,N_17612);
nand U18157 (N_18157,N_16727,N_17234);
or U18158 (N_18158,N_17894,N_16989);
nand U18159 (N_18159,N_17670,N_17859);
nand U18160 (N_18160,N_17303,N_17265);
or U18161 (N_18161,N_17009,N_17955);
and U18162 (N_18162,N_17829,N_17967);
xnor U18163 (N_18163,N_17889,N_17015);
nand U18164 (N_18164,N_17997,N_16596);
or U18165 (N_18165,N_17439,N_17596);
nor U18166 (N_18166,N_17734,N_17152);
xor U18167 (N_18167,N_17746,N_17531);
nand U18168 (N_18168,N_17468,N_17845);
or U18169 (N_18169,N_17933,N_17914);
nor U18170 (N_18170,N_17705,N_17098);
xor U18171 (N_18171,N_17509,N_16632);
or U18172 (N_18172,N_17207,N_16784);
nor U18173 (N_18173,N_16984,N_16670);
and U18174 (N_18174,N_17311,N_16779);
xnor U18175 (N_18175,N_17276,N_17382);
and U18176 (N_18176,N_16829,N_17735);
and U18177 (N_18177,N_17056,N_16936);
nand U18178 (N_18178,N_17343,N_17133);
xor U18179 (N_18179,N_17964,N_16825);
and U18180 (N_18180,N_16613,N_16832);
and U18181 (N_18181,N_16543,N_16680);
nand U18182 (N_18182,N_17794,N_17285);
nor U18183 (N_18183,N_16726,N_17868);
and U18184 (N_18184,N_16933,N_17915);
nor U18185 (N_18185,N_16601,N_17813);
nor U18186 (N_18186,N_16804,N_16873);
and U18187 (N_18187,N_17577,N_17283);
and U18188 (N_18188,N_17246,N_16920);
or U18189 (N_18189,N_17399,N_17551);
or U18190 (N_18190,N_17021,N_17099);
or U18191 (N_18191,N_16752,N_17477);
and U18192 (N_18192,N_17784,N_16841);
or U18193 (N_18193,N_17406,N_17522);
xnor U18194 (N_18194,N_16631,N_17959);
xor U18195 (N_18195,N_16878,N_17427);
nand U18196 (N_18196,N_16581,N_16762);
nand U18197 (N_18197,N_17087,N_17062);
and U18198 (N_18198,N_17275,N_17724);
nand U18199 (N_18199,N_17943,N_17241);
xor U18200 (N_18200,N_17395,N_17416);
nor U18201 (N_18201,N_17020,N_17070);
xnor U18202 (N_18202,N_16794,N_17961);
and U18203 (N_18203,N_17566,N_17397);
or U18204 (N_18204,N_17318,N_17139);
nor U18205 (N_18205,N_17239,N_17478);
nor U18206 (N_18206,N_16917,N_17268);
and U18207 (N_18207,N_17230,N_17057);
nor U18208 (N_18208,N_17523,N_17179);
xnor U18209 (N_18209,N_16659,N_16714);
nor U18210 (N_18210,N_17007,N_16529);
or U18211 (N_18211,N_17768,N_17499);
or U18212 (N_18212,N_17738,N_17646);
nor U18213 (N_18213,N_17591,N_17085);
or U18214 (N_18214,N_16556,N_17229);
nand U18215 (N_18215,N_17722,N_16840);
nand U18216 (N_18216,N_17405,N_17539);
or U18217 (N_18217,N_16772,N_17342);
nor U18218 (N_18218,N_16810,N_16706);
or U18219 (N_18219,N_17172,N_17155);
or U18220 (N_18220,N_17488,N_16566);
xor U18221 (N_18221,N_17224,N_17197);
nand U18222 (N_18222,N_16974,N_16759);
xor U18223 (N_18223,N_17010,N_17586);
xnor U18224 (N_18224,N_16954,N_17580);
and U18225 (N_18225,N_17983,N_16578);
nand U18226 (N_18226,N_17707,N_17374);
xnor U18227 (N_18227,N_17606,N_17017);
xor U18228 (N_18228,N_16718,N_17263);
nor U18229 (N_18229,N_17905,N_17240);
nand U18230 (N_18230,N_17528,N_17366);
xor U18231 (N_18231,N_17352,N_16814);
xnor U18232 (N_18232,N_17711,N_17322);
or U18233 (N_18233,N_17247,N_17390);
nor U18234 (N_18234,N_16769,N_17327);
and U18235 (N_18235,N_16922,N_17255);
xor U18236 (N_18236,N_16610,N_17838);
xor U18237 (N_18237,N_17543,N_17605);
and U18238 (N_18238,N_16580,N_17774);
nand U18239 (N_18239,N_17760,N_16515);
xor U18240 (N_18240,N_17158,N_16837);
nand U18241 (N_18241,N_17361,N_16863);
nand U18242 (N_18242,N_17990,N_17622);
nand U18243 (N_18243,N_16536,N_17389);
xnor U18244 (N_18244,N_17036,N_17479);
nor U18245 (N_18245,N_17107,N_17383);
xnor U18246 (N_18246,N_16777,N_17720);
nand U18247 (N_18247,N_17339,N_17993);
nor U18248 (N_18248,N_16918,N_17319);
or U18249 (N_18249,N_17833,N_16683);
and U18250 (N_18250,N_17718,N_16860);
nor U18251 (N_18251,N_16881,N_16964);
and U18252 (N_18252,N_17598,N_17850);
nor U18253 (N_18253,N_16865,N_17681);
nand U18254 (N_18254,N_17751,N_17051);
and U18255 (N_18255,N_17667,N_17284);
xor U18256 (N_18256,N_17946,N_17686);
and U18257 (N_18257,N_16886,N_17762);
xor U18258 (N_18258,N_17288,N_17378);
nor U18259 (N_18259,N_17925,N_17671);
nand U18260 (N_18260,N_17764,N_17047);
and U18261 (N_18261,N_17225,N_17082);
nand U18262 (N_18262,N_17676,N_16998);
nor U18263 (N_18263,N_17820,N_17856);
or U18264 (N_18264,N_16904,N_17228);
nor U18265 (N_18265,N_16876,N_17590);
or U18266 (N_18266,N_17680,N_17776);
and U18267 (N_18267,N_17526,N_16870);
and U18268 (N_18268,N_17778,N_17882);
xnor U18269 (N_18269,N_17907,N_16633);
nor U18270 (N_18270,N_16801,N_17497);
nand U18271 (N_18271,N_17976,N_17725);
xnor U18272 (N_18272,N_17424,N_16911);
xnor U18273 (N_18273,N_16600,N_16511);
or U18274 (N_18274,N_16586,N_16943);
xor U18275 (N_18275,N_17678,N_17912);
and U18276 (N_18276,N_17279,N_17828);
nor U18277 (N_18277,N_17326,N_17079);
xnor U18278 (N_18278,N_17183,N_17106);
xor U18279 (N_18279,N_17587,N_17330);
and U18280 (N_18280,N_17116,N_17782);
nand U18281 (N_18281,N_17035,N_17867);
nor U18282 (N_18282,N_17452,N_17002);
nor U18283 (N_18283,N_16986,N_16676);
xor U18284 (N_18284,N_16746,N_16711);
nor U18285 (N_18285,N_17851,N_16901);
nand U18286 (N_18286,N_17608,N_17184);
and U18287 (N_18287,N_17617,N_16679);
or U18288 (N_18288,N_16575,N_16571);
or U18289 (N_18289,N_17267,N_17450);
nand U18290 (N_18290,N_16822,N_17843);
nand U18291 (N_18291,N_17630,N_17963);
or U18292 (N_18292,N_17755,N_17687);
nand U18293 (N_18293,N_16775,N_17113);
or U18294 (N_18294,N_17385,N_17835);
or U18295 (N_18295,N_16649,N_17544);
nand U18296 (N_18296,N_17102,N_17236);
and U18297 (N_18297,N_17034,N_16811);
and U18298 (N_18298,N_17721,N_17315);
and U18299 (N_18299,N_17506,N_17977);
and U18300 (N_18300,N_17939,N_17641);
nand U18301 (N_18301,N_16809,N_16708);
and U18302 (N_18302,N_17910,N_16518);
nor U18303 (N_18303,N_17623,N_16574);
nor U18304 (N_18304,N_16820,N_17121);
or U18305 (N_18305,N_17805,N_16584);
or U18306 (N_18306,N_17187,N_17530);
nand U18307 (N_18307,N_17649,N_16760);
xor U18308 (N_18308,N_17391,N_17059);
and U18309 (N_18309,N_17250,N_17103);
nor U18310 (N_18310,N_17449,N_17412);
nor U18311 (N_18311,N_16565,N_17463);
nor U18312 (N_18312,N_16877,N_17659);
or U18313 (N_18313,N_16516,N_16931);
nor U18314 (N_18314,N_16912,N_17611);
nor U18315 (N_18315,N_17050,N_17086);
and U18316 (N_18316,N_17818,N_16579);
or U18317 (N_18317,N_16736,N_16806);
and U18318 (N_18318,N_17414,N_17677);
xor U18319 (N_18319,N_17362,N_17262);
xor U18320 (N_18320,N_17492,N_16666);
nor U18321 (N_18321,N_17161,N_17486);
nand U18322 (N_18322,N_17029,N_17307);
nand U18323 (N_18323,N_16501,N_17870);
or U18324 (N_18324,N_17160,N_17415);
or U18325 (N_18325,N_17088,N_17398);
nor U18326 (N_18326,N_17411,N_17485);
nand U18327 (N_18327,N_17191,N_16671);
nand U18328 (N_18328,N_17675,N_17842);
and U18329 (N_18329,N_17118,N_16791);
xor U18330 (N_18330,N_16818,N_17494);
xor U18331 (N_18331,N_16634,N_16642);
nor U18332 (N_18332,N_17825,N_17138);
nand U18333 (N_18333,N_16898,N_17260);
nor U18334 (N_18334,N_17702,N_17074);
nand U18335 (N_18335,N_17973,N_17708);
or U18336 (N_18336,N_16729,N_17938);
nand U18337 (N_18337,N_17217,N_16715);
xnor U18338 (N_18338,N_17848,N_17042);
xor U18339 (N_18339,N_16962,N_17136);
nand U18340 (N_18340,N_17300,N_16947);
or U18341 (N_18341,N_17001,N_16598);
nand U18342 (N_18342,N_17791,N_17500);
or U18343 (N_18343,N_17978,N_16887);
and U18344 (N_18344,N_16782,N_16973);
xor U18345 (N_18345,N_16564,N_17634);
xnor U18346 (N_18346,N_17115,N_17874);
xor U18347 (N_18347,N_16915,N_17324);
or U18348 (N_18348,N_17192,N_16903);
and U18349 (N_18349,N_17461,N_16611);
or U18350 (N_18350,N_16952,N_17901);
and U18351 (N_18351,N_17501,N_16675);
and U18352 (N_18352,N_17186,N_17465);
nand U18353 (N_18353,N_17638,N_17135);
and U18354 (N_18354,N_17493,N_16764);
nand U18355 (N_18355,N_16833,N_17198);
and U18356 (N_18356,N_16524,N_16941);
nand U18357 (N_18357,N_17446,N_16838);
and U18358 (N_18358,N_17553,N_17831);
nand U18359 (N_18359,N_17407,N_17278);
or U18360 (N_18360,N_17525,N_16790);
xor U18361 (N_18361,N_17438,N_16905);
or U18362 (N_18362,N_17472,N_17297);
xnor U18363 (N_18363,N_16572,N_17926);
nor U18364 (N_18364,N_17913,N_16520);
nor U18365 (N_18365,N_17518,N_16590);
or U18366 (N_18366,N_17457,N_17883);
nand U18367 (N_18367,N_17402,N_16527);
nor U18368 (N_18368,N_17684,N_16798);
nor U18369 (N_18369,N_17652,N_16743);
and U18370 (N_18370,N_17559,N_17801);
xnor U18371 (N_18371,N_16795,N_17787);
and U18372 (N_18372,N_16616,N_17949);
xor U18373 (N_18373,N_17727,N_16800);
or U18374 (N_18374,N_17994,N_17249);
nand U18375 (N_18375,N_16856,N_17900);
nor U18376 (N_18376,N_17189,N_16547);
or U18377 (N_18377,N_16836,N_17830);
or U18378 (N_18378,N_17204,N_17555);
or U18379 (N_18379,N_17129,N_17541);
xor U18380 (N_18380,N_17556,N_17569);
nor U18381 (N_18381,N_17502,N_17373);
or U18382 (N_18382,N_17713,N_17890);
nand U18383 (N_18383,N_17321,N_17753);
nand U18384 (N_18384,N_17370,N_17137);
xnor U18385 (N_18385,N_17574,N_17312);
and U18386 (N_18386,N_16599,N_17621);
or U18387 (N_18387,N_16562,N_17576);
nor U18388 (N_18388,N_17930,N_16882);
and U18389 (N_18389,N_17495,N_17076);
nor U18390 (N_18390,N_16894,N_17733);
xnor U18391 (N_18391,N_17299,N_17732);
and U18392 (N_18392,N_17019,N_17906);
xor U18393 (N_18393,N_16907,N_16935);
and U18394 (N_18394,N_17094,N_17359);
nand U18395 (N_18395,N_17908,N_17618);
and U18396 (N_18396,N_17811,N_17203);
and U18397 (N_18397,N_17771,N_17745);
nor U18398 (N_18398,N_16981,N_16889);
or U18399 (N_18399,N_17281,N_16970);
xor U18400 (N_18400,N_17037,N_16528);
and U18401 (N_18401,N_17785,N_16834);
and U18402 (N_18402,N_16545,N_17840);
nor U18403 (N_18403,N_17985,N_17159);
nor U18404 (N_18404,N_17816,N_17248);
nand U18405 (N_18405,N_17141,N_16544);
or U18406 (N_18406,N_17613,N_17081);
or U18407 (N_18407,N_16688,N_16824);
xnor U18408 (N_18408,N_17731,N_16946);
xor U18409 (N_18409,N_17055,N_16673);
or U18410 (N_18410,N_17346,N_16910);
xor U18411 (N_18411,N_16908,N_17458);
or U18412 (N_18412,N_16993,N_16872);
or U18413 (N_18413,N_16843,N_17075);
or U18414 (N_18414,N_17583,N_17096);
xor U18415 (N_18415,N_17934,N_17176);
xor U18416 (N_18416,N_17104,N_16845);
and U18417 (N_18417,N_17749,N_17562);
nand U18418 (N_18418,N_17254,N_17291);
or U18419 (N_18419,N_17879,N_17542);
xor U18420 (N_18420,N_17264,N_17006);
nor U18421 (N_18421,N_17171,N_16591);
nor U18422 (N_18422,N_16937,N_16617);
xnor U18423 (N_18423,N_17245,N_17221);
and U18424 (N_18424,N_16661,N_16850);
xor U18425 (N_18425,N_16789,N_16858);
nor U18426 (N_18426,N_17761,N_16960);
nor U18427 (N_18427,N_17375,N_17156);
nor U18428 (N_18428,N_17999,N_16793);
nand U18429 (N_18429,N_17462,N_17040);
nand U18430 (N_18430,N_17897,N_16728);
or U18431 (N_18431,N_16745,N_17832);
nor U18432 (N_18432,N_17899,N_17632);
nand U18433 (N_18433,N_16997,N_16540);
nor U18434 (N_18434,N_17892,N_17403);
nor U18435 (N_18435,N_16742,N_16568);
or U18436 (N_18436,N_16606,N_16505);
nand U18437 (N_18437,N_16975,N_16740);
nand U18438 (N_18438,N_17554,N_17475);
or U18439 (N_18439,N_17164,N_17703);
or U18440 (N_18440,N_17344,N_16999);
nand U18441 (N_18441,N_16761,N_17662);
xor U18442 (N_18442,N_17496,N_17100);
nor U18443 (N_18443,N_17372,N_17182);
or U18444 (N_18444,N_17928,N_17588);
nor U18445 (N_18445,N_17292,N_17282);
xnor U18446 (N_18446,N_17393,N_17736);
nor U18447 (N_18447,N_17565,N_16766);
or U18448 (N_18448,N_16768,N_17027);
nor U18449 (N_18449,N_17529,N_17043);
and U18450 (N_18450,N_16539,N_17442);
or U18451 (N_18451,N_17827,N_17329);
and U18452 (N_18452,N_17261,N_17193);
nor U18453 (N_18453,N_16672,N_16502);
nand U18454 (N_18454,N_17243,N_16563);
nor U18455 (N_18455,N_17126,N_17441);
xor U18456 (N_18456,N_16853,N_16797);
and U18457 (N_18457,N_17258,N_17837);
and U18458 (N_18458,N_17331,N_17132);
and U18459 (N_18459,N_16967,N_16707);
nand U18460 (N_18460,N_17423,N_17826);
or U18461 (N_18461,N_17710,N_16996);
nor U18462 (N_18462,N_17754,N_17527);
and U18463 (N_18463,N_16939,N_17046);
nand U18464 (N_18464,N_17979,N_16689);
or U18465 (N_18465,N_16667,N_16821);
and U18466 (N_18466,N_17898,N_16842);
or U18467 (N_18467,N_17440,N_16558);
xnor U18468 (N_18468,N_17409,N_17363);
xnor U18469 (N_18469,N_16709,N_16592);
and U18470 (N_18470,N_17797,N_16785);
nand U18471 (N_18471,N_17594,N_16875);
or U18472 (N_18472,N_17800,N_17093);
nor U18473 (N_18473,N_16526,N_16653);
or U18474 (N_18474,N_16694,N_17616);
and U18475 (N_18475,N_17162,N_17123);
or U18476 (N_18476,N_16570,N_17447);
nand U18477 (N_18477,N_17124,N_17592);
nand U18478 (N_18478,N_17699,N_17624);
or U18479 (N_18479,N_17759,N_17857);
nor U18480 (N_18480,N_17210,N_17271);
or U18481 (N_18481,N_17381,N_16561);
and U18482 (N_18482,N_17277,N_16906);
and U18483 (N_18483,N_17490,N_17674);
nand U18484 (N_18484,N_16664,N_16552);
and U18485 (N_18485,N_16638,N_16582);
and U18486 (N_18486,N_17273,N_16731);
or U18487 (N_18487,N_17780,N_17175);
and U18488 (N_18488,N_17861,N_17143);
nor U18489 (N_18489,N_17719,N_17431);
nor U18490 (N_18490,N_17631,N_17163);
nand U18491 (N_18491,N_17400,N_17354);
nor U18492 (N_18492,N_17936,N_17012);
or U18493 (N_18493,N_17871,N_17563);
or U18494 (N_18494,N_17272,N_16549);
and U18495 (N_18495,N_17807,N_17957);
and U18496 (N_18496,N_17024,N_16788);
nor U18497 (N_18497,N_16703,N_16730);
xor U18498 (N_18498,N_16978,N_16929);
and U18499 (N_18499,N_17369,N_17350);
and U18500 (N_18500,N_17433,N_17693);
nand U18501 (N_18501,N_17218,N_16756);
nor U18502 (N_18502,N_17232,N_17920);
nand U18503 (N_18503,N_16879,N_17716);
nand U18504 (N_18504,N_16721,N_16594);
nor U18505 (N_18505,N_17168,N_17380);
and U18506 (N_18506,N_16719,N_16588);
or U18507 (N_18507,N_17803,N_16517);
or U18508 (N_18508,N_17513,N_17607);
nand U18509 (N_18509,N_16971,N_17028);
xnor U18510 (N_18510,N_17294,N_16602);
and U18511 (N_18511,N_16604,N_16839);
or U18512 (N_18512,N_17474,N_17110);
xor U18513 (N_18513,N_16663,N_17597);
and U18514 (N_18514,N_17039,N_17095);
or U18515 (N_18515,N_17080,N_17148);
and U18516 (N_18516,N_17286,N_16969);
or U18517 (N_18517,N_17165,N_17923);
xor U18518 (N_18518,N_17635,N_16510);
and U18519 (N_18519,N_17222,N_17066);
or U18520 (N_18520,N_17672,N_17202);
nor U18521 (N_18521,N_17692,N_17508);
or U18522 (N_18522,N_17313,N_17436);
and U18523 (N_18523,N_17691,N_16828);
nand U18524 (N_18524,N_17579,N_16813);
nand U18525 (N_18525,N_17090,N_17604);
xor U18526 (N_18526,N_17023,N_16869);
xnor U18527 (N_18527,N_17227,N_16691);
and U18528 (N_18528,N_16739,N_16991);
or U18529 (N_18529,N_17712,N_17306);
and U18530 (N_18530,N_17334,N_17432);
and U18531 (N_18531,N_17786,N_17293);
or U18532 (N_18532,N_16776,N_17131);
and U18533 (N_18533,N_16548,N_16640);
or U18534 (N_18534,N_16646,N_17435);
and U18535 (N_18535,N_17685,N_17201);
xor U18536 (N_18536,N_17031,N_17242);
nand U18537 (N_18537,N_17016,N_16744);
xnor U18538 (N_18538,N_17517,N_17120);
nand U18539 (N_18539,N_16900,N_17058);
xor U18540 (N_18540,N_17428,N_16595);
and U18541 (N_18541,N_17379,N_17571);
xor U18542 (N_18542,N_16684,N_16948);
nor U18543 (N_18543,N_17808,N_17881);
xor U18544 (N_18544,N_17704,N_17996);
or U18545 (N_18545,N_17392,N_16805);
nor U18546 (N_18546,N_16758,N_16961);
and U18547 (N_18547,N_17026,N_16934);
nor U18548 (N_18548,N_16541,N_17341);
nand U18549 (N_18549,N_17929,N_16802);
xor U18550 (N_18550,N_17078,N_17593);
and U18551 (N_18551,N_17877,N_17921);
nand U18552 (N_18552,N_17190,N_17765);
xor U18553 (N_18553,N_16763,N_17615);
nand U18554 (N_18554,N_16958,N_17540);
or U18555 (N_18555,N_17194,N_16687);
and U18556 (N_18556,N_17643,N_17220);
xor U18557 (N_18557,N_16786,N_17169);
and U18558 (N_18558,N_16857,N_17301);
nor U18559 (N_18559,N_17340,N_17092);
or U18560 (N_18560,N_17855,N_16748);
xor U18561 (N_18561,N_16553,N_16623);
xor U18562 (N_18562,N_16741,N_17998);
nor U18563 (N_18563,N_17742,N_17664);
or U18564 (N_18564,N_17073,N_17876);
nor U18565 (N_18565,N_17200,N_16500);
or U18566 (N_18566,N_17942,N_16644);
and U18567 (N_18567,N_17944,N_16754);
xor U18568 (N_18568,N_16681,N_17657);
nor U18569 (N_18569,N_17335,N_17174);
nand U18570 (N_18570,N_16686,N_17885);
or U18571 (N_18571,N_16669,N_16698);
nor U18572 (N_18572,N_17510,N_17257);
nand U18573 (N_18573,N_16871,N_16722);
or U18574 (N_18574,N_16734,N_17445);
nor U18575 (N_18575,N_17799,N_17537);
or U18576 (N_18576,N_17969,N_17941);
nor U18577 (N_18577,N_17860,N_17212);
nor U18578 (N_18578,N_16994,N_16750);
nor U18579 (N_18579,N_17975,N_16897);
nand U18580 (N_18580,N_17866,N_17709);
and U18581 (N_18581,N_16643,N_16662);
nand U18582 (N_18582,N_16848,N_17642);
xor U18583 (N_18583,N_17018,N_17640);
and U18584 (N_18584,N_17595,N_17309);
or U18585 (N_18585,N_16892,N_16938);
and U18586 (N_18586,N_17421,N_17603);
and U18587 (N_18587,N_17763,N_16668);
and U18588 (N_18588,N_17214,N_16625);
nand U18589 (N_18589,N_17296,N_17698);
xnor U18590 (N_18590,N_17349,N_16717);
xor U18591 (N_18591,N_16577,N_17180);
and U18592 (N_18592,N_17231,N_17965);
or U18593 (N_18593,N_17637,N_16968);
xnor U18594 (N_18594,N_17986,N_16972);
or U18595 (N_18595,N_17766,N_16530);
nand U18596 (N_18596,N_17188,N_16965);
and U18597 (N_18597,N_16630,N_16546);
or U18598 (N_18598,N_17401,N_16851);
nor U18599 (N_18599,N_17157,N_17849);
nor U18600 (N_18600,N_16550,N_17619);
or U18601 (N_18601,N_16951,N_17945);
nand U18602 (N_18602,N_17338,N_17410);
and U18603 (N_18603,N_17166,N_16682);
and U18604 (N_18604,N_17470,N_16866);
xnor U18605 (N_18605,N_16723,N_17846);
xnor U18606 (N_18606,N_17697,N_17980);
nand U18607 (N_18607,N_17426,N_17815);
and U18608 (N_18608,N_17417,N_17140);
xnor U18609 (N_18609,N_17005,N_17744);
nor U18610 (N_18610,N_17185,N_16767);
xor U18611 (N_18611,N_17101,N_16956);
and U18612 (N_18612,N_16641,N_17552);
xnor U18613 (N_18613,N_17487,N_16705);
nand U18614 (N_18614,N_16519,N_16647);
and U18615 (N_18615,N_17974,N_16712);
and U18616 (N_18616,N_17437,N_17253);
or U18617 (N_18617,N_17044,N_16532);
nor U18618 (N_18618,N_16503,N_17862);
and U18619 (N_18619,N_16534,N_16713);
xnor U18620 (N_18620,N_17972,N_16874);
xor U18621 (N_18621,N_17304,N_16674);
and U18622 (N_18622,N_16559,N_17777);
or U18623 (N_18623,N_17844,N_17355);
and U18624 (N_18624,N_17351,N_17792);
nand U18625 (N_18625,N_16654,N_17061);
xor U18626 (N_18626,N_17823,N_17834);
xor U18627 (N_18627,N_16831,N_16770);
xor U18628 (N_18628,N_17694,N_16861);
or U18629 (N_18629,N_17575,N_17396);
nand U18630 (N_18630,N_16538,N_17459);
or U18631 (N_18631,N_17810,N_17289);
and U18632 (N_18632,N_17420,N_16677);
xnor U18633 (N_18633,N_17205,N_16542);
nand U18634 (N_18634,N_17484,N_17511);
or U18635 (N_18635,N_17316,N_16639);
and U18636 (N_18636,N_17014,N_16923);
xnor U18637 (N_18637,N_17653,N_16796);
nor U18638 (N_18638,N_17589,N_16692);
xor U18639 (N_18639,N_16678,N_17546);
nand U18640 (N_18640,N_17822,N_17325);
nor U18641 (N_18641,N_16928,N_17444);
or U18642 (N_18642,N_17150,N_17060);
nand U18643 (N_18643,N_17453,N_17695);
nor U18644 (N_18644,N_16985,N_16508);
and U18645 (N_18645,N_17666,N_17561);
or U18646 (N_18646,N_17127,N_16799);
nand U18647 (N_18647,N_16844,N_17041);
nor U18648 (N_18648,N_17503,N_17891);
nand U18649 (N_18649,N_17388,N_17033);
xor U18650 (N_18650,N_17564,N_17750);
nand U18651 (N_18651,N_17954,N_16890);
xnor U18652 (N_18652,N_16855,N_17931);
nor U18653 (N_18653,N_17690,N_17514);
nor U18654 (N_18654,N_16609,N_17302);
and U18655 (N_18655,N_17773,N_17648);
xor U18656 (N_18656,N_16699,N_17909);
and U18657 (N_18657,N_16757,N_17661);
or U18658 (N_18658,N_17003,N_17460);
xnor U18659 (N_18659,N_17873,N_17903);
nand U18660 (N_18660,N_16695,N_17356);
nand U18661 (N_18661,N_17280,N_16854);
nand U18662 (N_18662,N_17252,N_17425);
or U18663 (N_18663,N_17532,N_17422);
nor U18664 (N_18664,N_17817,N_16755);
nor U18665 (N_18665,N_17650,N_16787);
xnor U18666 (N_18666,N_16771,N_17679);
or U18667 (N_18667,N_17345,N_17570);
xnor U18668 (N_18668,N_17752,N_17512);
nand U18669 (N_18669,N_17434,N_17149);
and U18670 (N_18670,N_17371,N_16733);
xnor U18671 (N_18671,N_17758,N_16710);
xor U18672 (N_18672,N_17918,N_16957);
or U18673 (N_18673,N_16525,N_16765);
nand U18674 (N_18674,N_16868,N_17668);
or U18675 (N_18675,N_16893,N_16573);
and U18676 (N_18676,N_17781,N_17878);
xnor U18677 (N_18677,N_16618,N_17560);
nor U18678 (N_18678,N_16862,N_17153);
nor U18679 (N_18679,N_17142,N_17384);
and U18680 (N_18680,N_16792,N_16697);
xnor U18681 (N_18681,N_17536,N_16823);
and U18682 (N_18682,N_17880,N_17814);
or U18683 (N_18683,N_17429,N_17347);
nand U18684 (N_18684,N_17519,N_17854);
xor U18685 (N_18685,N_17984,N_17948);
nor U18686 (N_18686,N_17310,N_17962);
nor U18687 (N_18687,N_17886,N_16605);
nand U18688 (N_18688,N_16507,N_17146);
nor U18689 (N_18689,N_17022,N_17770);
nand U18690 (N_18690,N_17491,N_17958);
nor U18691 (N_18691,N_17332,N_17717);
and U18692 (N_18692,N_17769,N_17927);
xor U18693 (N_18693,N_17847,N_17117);
or U18694 (N_18694,N_17219,N_17887);
or U18695 (N_18695,N_17669,N_16803);
and U18696 (N_18696,N_17573,N_16983);
xor U18697 (N_18697,N_17779,N_17626);
nand U18698 (N_18698,N_17089,N_16949);
xor U18699 (N_18699,N_17809,N_16817);
nor U18700 (N_18700,N_17455,N_17584);
or U18701 (N_18701,N_16624,N_16660);
nand U18702 (N_18702,N_17467,N_17696);
and U18703 (N_18703,N_16535,N_16924);
nand U18704 (N_18704,N_17940,N_16635);
xor U18705 (N_18705,N_16783,N_17966);
and U18706 (N_18706,N_16704,N_17516);
nand U18707 (N_18707,N_16509,N_17916);
nand U18708 (N_18708,N_16620,N_17011);
or U18709 (N_18709,N_17216,N_16867);
and U18710 (N_18710,N_17333,N_16645);
and U18711 (N_18711,N_17308,N_17988);
nand U18712 (N_18712,N_17004,N_17314);
xor U18713 (N_18713,N_16751,N_17952);
nand U18714 (N_18714,N_17737,N_16747);
or U18715 (N_18715,N_17077,N_16585);
and U18716 (N_18716,N_17600,N_17726);
and U18717 (N_18717,N_17812,N_16612);
nand U18718 (N_18718,N_17259,N_16942);
or U18719 (N_18719,N_16513,N_16921);
nor U18720 (N_18720,N_16945,N_17956);
xnor U18721 (N_18721,N_16940,N_17715);
xor U18722 (N_18722,N_17320,N_17025);
and U18723 (N_18723,N_17796,N_17633);
and U18724 (N_18724,N_17367,N_17645);
xnor U18725 (N_18725,N_16976,N_17430);
xor U18726 (N_18726,N_17888,N_16883);
or U18727 (N_18727,N_17767,N_17804);
and U18728 (N_18728,N_17545,N_17627);
xnor U18729 (N_18729,N_17067,N_16521);
and U18730 (N_18730,N_17473,N_16696);
xor U18731 (N_18731,N_17656,N_17739);
nor U18732 (N_18732,N_17919,N_17223);
or U18733 (N_18733,N_17125,N_17757);
xnor U18734 (N_18734,N_17233,N_16587);
and U18735 (N_18735,N_17995,N_17170);
nand U18736 (N_18736,N_16650,N_16913);
and U18737 (N_18737,N_17128,N_17151);
or U18738 (N_18738,N_17863,N_17498);
and U18739 (N_18739,N_17743,N_16597);
nor U18740 (N_18740,N_17683,N_17360);
xor U18741 (N_18741,N_17572,N_17629);
or U18742 (N_18742,N_17775,N_17317);
and U18743 (N_18743,N_17982,N_17547);
nand U18744 (N_18744,N_17628,N_17091);
nor U18745 (N_18745,N_17665,N_16701);
or U18746 (N_18746,N_17625,N_17298);
nor U18747 (N_18747,N_17451,N_17740);
or U18748 (N_18748,N_16648,N_16885);
xor U18749 (N_18749,N_17064,N_17953);
and U18750 (N_18750,N_17799,N_17082);
nand U18751 (N_18751,N_16779,N_16951);
and U18752 (N_18752,N_17141,N_16897);
xor U18753 (N_18753,N_16589,N_17187);
xor U18754 (N_18754,N_16858,N_16707);
or U18755 (N_18755,N_17831,N_17662);
nor U18756 (N_18756,N_17454,N_17398);
xor U18757 (N_18757,N_17023,N_17313);
nor U18758 (N_18758,N_17803,N_16953);
xnor U18759 (N_18759,N_16913,N_17456);
or U18760 (N_18760,N_16818,N_17269);
nor U18761 (N_18761,N_17392,N_17557);
nand U18762 (N_18762,N_16645,N_17937);
nor U18763 (N_18763,N_17311,N_17020);
and U18764 (N_18764,N_16652,N_17048);
nor U18765 (N_18765,N_17499,N_16806);
and U18766 (N_18766,N_17794,N_16911);
nor U18767 (N_18767,N_16794,N_16902);
and U18768 (N_18768,N_17882,N_17341);
and U18769 (N_18769,N_17822,N_17253);
nand U18770 (N_18770,N_17889,N_16670);
nor U18771 (N_18771,N_17046,N_17259);
nand U18772 (N_18772,N_17930,N_17697);
and U18773 (N_18773,N_16869,N_16931);
or U18774 (N_18774,N_17575,N_17630);
and U18775 (N_18775,N_17708,N_16531);
xnor U18776 (N_18776,N_17584,N_16873);
nand U18777 (N_18777,N_17225,N_17627);
xor U18778 (N_18778,N_17104,N_16570);
nor U18779 (N_18779,N_16728,N_17299);
nand U18780 (N_18780,N_17711,N_17206);
and U18781 (N_18781,N_16871,N_16892);
or U18782 (N_18782,N_17579,N_16657);
and U18783 (N_18783,N_17862,N_17591);
xnor U18784 (N_18784,N_17129,N_17011);
xnor U18785 (N_18785,N_17717,N_16782);
xnor U18786 (N_18786,N_17830,N_17769);
xor U18787 (N_18787,N_17348,N_16714);
and U18788 (N_18788,N_17400,N_16998);
and U18789 (N_18789,N_17609,N_17953);
and U18790 (N_18790,N_17990,N_17610);
and U18791 (N_18791,N_17023,N_17538);
or U18792 (N_18792,N_17545,N_16737);
nand U18793 (N_18793,N_17760,N_17497);
xor U18794 (N_18794,N_17761,N_17707);
nor U18795 (N_18795,N_17618,N_17941);
nand U18796 (N_18796,N_17859,N_17907);
and U18797 (N_18797,N_17726,N_17801);
or U18798 (N_18798,N_17391,N_17052);
xor U18799 (N_18799,N_17575,N_17316);
xnor U18800 (N_18800,N_16834,N_16534);
and U18801 (N_18801,N_16980,N_16624);
nand U18802 (N_18802,N_16975,N_16818);
and U18803 (N_18803,N_16862,N_16913);
xnor U18804 (N_18804,N_16786,N_16932);
nand U18805 (N_18805,N_17464,N_17376);
nor U18806 (N_18806,N_16731,N_16620);
or U18807 (N_18807,N_17310,N_16863);
xnor U18808 (N_18808,N_17955,N_16564);
nand U18809 (N_18809,N_17106,N_17616);
nand U18810 (N_18810,N_17448,N_17132);
and U18811 (N_18811,N_17018,N_16506);
nor U18812 (N_18812,N_17963,N_17438);
or U18813 (N_18813,N_16635,N_17031);
or U18814 (N_18814,N_17629,N_17953);
nor U18815 (N_18815,N_17186,N_17946);
nand U18816 (N_18816,N_17646,N_16775);
or U18817 (N_18817,N_17426,N_16671);
nor U18818 (N_18818,N_17921,N_17183);
xnor U18819 (N_18819,N_17057,N_16882);
or U18820 (N_18820,N_17303,N_17688);
xnor U18821 (N_18821,N_17256,N_17290);
xnor U18822 (N_18822,N_16507,N_16659);
nand U18823 (N_18823,N_17770,N_16815);
xnor U18824 (N_18824,N_17817,N_17336);
and U18825 (N_18825,N_16700,N_17968);
nor U18826 (N_18826,N_17135,N_16661);
or U18827 (N_18827,N_17087,N_16708);
nand U18828 (N_18828,N_17449,N_16916);
or U18829 (N_18829,N_17255,N_16904);
nor U18830 (N_18830,N_17631,N_17915);
or U18831 (N_18831,N_16888,N_16565);
or U18832 (N_18832,N_17339,N_16511);
nor U18833 (N_18833,N_17733,N_17783);
and U18834 (N_18834,N_17969,N_16580);
nand U18835 (N_18835,N_17112,N_17308);
or U18836 (N_18836,N_17470,N_16918);
or U18837 (N_18837,N_17807,N_17362);
nor U18838 (N_18838,N_17026,N_16801);
or U18839 (N_18839,N_17025,N_17529);
and U18840 (N_18840,N_16829,N_16904);
or U18841 (N_18841,N_16934,N_16604);
or U18842 (N_18842,N_16525,N_17216);
xor U18843 (N_18843,N_17690,N_16985);
nor U18844 (N_18844,N_17454,N_17199);
or U18845 (N_18845,N_17646,N_16927);
nor U18846 (N_18846,N_17908,N_17038);
or U18847 (N_18847,N_16853,N_17073);
xor U18848 (N_18848,N_17358,N_17448);
nor U18849 (N_18849,N_16895,N_16663);
and U18850 (N_18850,N_16595,N_17020);
xnor U18851 (N_18851,N_16905,N_16671);
or U18852 (N_18852,N_16753,N_17196);
or U18853 (N_18853,N_17213,N_17058);
nor U18854 (N_18854,N_16608,N_17243);
nor U18855 (N_18855,N_17516,N_17144);
nand U18856 (N_18856,N_17495,N_17397);
nand U18857 (N_18857,N_17876,N_17918);
or U18858 (N_18858,N_16898,N_17318);
xor U18859 (N_18859,N_17924,N_16977);
nor U18860 (N_18860,N_17197,N_17752);
and U18861 (N_18861,N_17045,N_17734);
and U18862 (N_18862,N_17267,N_16719);
nor U18863 (N_18863,N_16906,N_16973);
nand U18864 (N_18864,N_17217,N_17174);
nor U18865 (N_18865,N_16833,N_17674);
and U18866 (N_18866,N_16965,N_17402);
nor U18867 (N_18867,N_17516,N_17735);
and U18868 (N_18868,N_17119,N_17517);
and U18869 (N_18869,N_17116,N_17473);
nand U18870 (N_18870,N_17164,N_17454);
nand U18871 (N_18871,N_17497,N_17813);
nand U18872 (N_18872,N_16912,N_17679);
or U18873 (N_18873,N_17598,N_17808);
and U18874 (N_18874,N_17690,N_17931);
nand U18875 (N_18875,N_16628,N_17455);
or U18876 (N_18876,N_17889,N_16589);
xnor U18877 (N_18877,N_16569,N_17027);
nand U18878 (N_18878,N_17144,N_16934);
or U18879 (N_18879,N_17656,N_17819);
or U18880 (N_18880,N_16534,N_16756);
xnor U18881 (N_18881,N_17536,N_16811);
and U18882 (N_18882,N_17939,N_17494);
or U18883 (N_18883,N_17847,N_17716);
xnor U18884 (N_18884,N_16571,N_17182);
nand U18885 (N_18885,N_16720,N_17062);
nor U18886 (N_18886,N_17339,N_17638);
nor U18887 (N_18887,N_17566,N_17947);
nor U18888 (N_18888,N_17696,N_17958);
xnor U18889 (N_18889,N_17155,N_16612);
xnor U18890 (N_18890,N_17088,N_17021);
nor U18891 (N_18891,N_17387,N_17826);
xor U18892 (N_18892,N_17947,N_17341);
and U18893 (N_18893,N_17050,N_17598);
nand U18894 (N_18894,N_17277,N_17549);
xnor U18895 (N_18895,N_17750,N_17620);
nand U18896 (N_18896,N_17842,N_17653);
xor U18897 (N_18897,N_17153,N_17440);
nand U18898 (N_18898,N_17012,N_17712);
or U18899 (N_18899,N_17839,N_17719);
or U18900 (N_18900,N_17081,N_16548);
nand U18901 (N_18901,N_17671,N_16681);
xor U18902 (N_18902,N_17970,N_17830);
or U18903 (N_18903,N_17917,N_17590);
nor U18904 (N_18904,N_17102,N_17184);
nor U18905 (N_18905,N_17739,N_17735);
nor U18906 (N_18906,N_17294,N_17442);
nor U18907 (N_18907,N_17200,N_17606);
nor U18908 (N_18908,N_17870,N_17387);
xnor U18909 (N_18909,N_16913,N_16664);
and U18910 (N_18910,N_16876,N_16839);
or U18911 (N_18911,N_17965,N_16546);
nor U18912 (N_18912,N_16779,N_16515);
nand U18913 (N_18913,N_16933,N_16503);
xnor U18914 (N_18914,N_16904,N_16612);
nor U18915 (N_18915,N_17524,N_17289);
xor U18916 (N_18916,N_16855,N_17828);
and U18917 (N_18917,N_17988,N_16739);
nor U18918 (N_18918,N_17945,N_17593);
or U18919 (N_18919,N_17028,N_17882);
and U18920 (N_18920,N_16649,N_16576);
and U18921 (N_18921,N_16680,N_16654);
or U18922 (N_18922,N_16841,N_17202);
nor U18923 (N_18923,N_16765,N_17186);
nor U18924 (N_18924,N_17187,N_17897);
nand U18925 (N_18925,N_16892,N_16849);
or U18926 (N_18926,N_16913,N_16905);
nand U18927 (N_18927,N_17174,N_17259);
and U18928 (N_18928,N_17537,N_16864);
xnor U18929 (N_18929,N_17442,N_17608);
nand U18930 (N_18930,N_17765,N_16564);
nor U18931 (N_18931,N_16701,N_17408);
or U18932 (N_18932,N_17923,N_16508);
nor U18933 (N_18933,N_17747,N_17053);
nand U18934 (N_18934,N_16664,N_17443);
or U18935 (N_18935,N_17364,N_16984);
or U18936 (N_18936,N_17806,N_16749);
nand U18937 (N_18937,N_16638,N_16589);
or U18938 (N_18938,N_17566,N_17217);
xor U18939 (N_18939,N_17900,N_17023);
nand U18940 (N_18940,N_17255,N_17629);
nand U18941 (N_18941,N_17429,N_16899);
xnor U18942 (N_18942,N_16963,N_17281);
or U18943 (N_18943,N_17438,N_16962);
nand U18944 (N_18944,N_17844,N_17559);
nand U18945 (N_18945,N_16853,N_17227);
nand U18946 (N_18946,N_16662,N_17459);
and U18947 (N_18947,N_17193,N_17365);
nor U18948 (N_18948,N_17492,N_17034);
nand U18949 (N_18949,N_17894,N_17439);
or U18950 (N_18950,N_16834,N_16926);
nor U18951 (N_18951,N_16536,N_17212);
or U18952 (N_18952,N_17111,N_17300);
nor U18953 (N_18953,N_16793,N_16643);
and U18954 (N_18954,N_17459,N_17201);
nand U18955 (N_18955,N_16773,N_16812);
or U18956 (N_18956,N_16501,N_16817);
xor U18957 (N_18957,N_17810,N_17278);
or U18958 (N_18958,N_17266,N_17694);
xor U18959 (N_18959,N_17732,N_16939);
xor U18960 (N_18960,N_17963,N_16682);
nand U18961 (N_18961,N_17423,N_17528);
or U18962 (N_18962,N_16743,N_17595);
nand U18963 (N_18963,N_16955,N_16700);
nand U18964 (N_18964,N_17652,N_17897);
nor U18965 (N_18965,N_16610,N_16938);
nor U18966 (N_18966,N_17656,N_17585);
xor U18967 (N_18967,N_17686,N_17891);
nor U18968 (N_18968,N_17473,N_17785);
nand U18969 (N_18969,N_17322,N_17126);
nor U18970 (N_18970,N_17439,N_16974);
or U18971 (N_18971,N_16960,N_17942);
nor U18972 (N_18972,N_17873,N_16504);
and U18973 (N_18973,N_17767,N_17679);
nor U18974 (N_18974,N_16838,N_17305);
and U18975 (N_18975,N_16550,N_17163);
and U18976 (N_18976,N_17472,N_16785);
nand U18977 (N_18977,N_17486,N_17047);
and U18978 (N_18978,N_17802,N_16651);
nor U18979 (N_18979,N_16579,N_17150);
or U18980 (N_18980,N_17519,N_16894);
nand U18981 (N_18981,N_17682,N_16973);
xor U18982 (N_18982,N_17678,N_17444);
nor U18983 (N_18983,N_17824,N_17744);
or U18984 (N_18984,N_17784,N_17917);
nor U18985 (N_18985,N_16563,N_17275);
nor U18986 (N_18986,N_17244,N_17026);
and U18987 (N_18987,N_17965,N_17222);
or U18988 (N_18988,N_17196,N_17578);
nand U18989 (N_18989,N_17158,N_17526);
and U18990 (N_18990,N_17880,N_16988);
and U18991 (N_18991,N_16748,N_17302);
nand U18992 (N_18992,N_17853,N_17616);
nand U18993 (N_18993,N_17675,N_17910);
nand U18994 (N_18994,N_16677,N_17961);
xnor U18995 (N_18995,N_17098,N_17191);
nand U18996 (N_18996,N_16893,N_16930);
nand U18997 (N_18997,N_17653,N_16704);
nor U18998 (N_18998,N_17256,N_16750);
xnor U18999 (N_18999,N_16851,N_16637);
and U19000 (N_19000,N_17776,N_17230);
or U19001 (N_19001,N_17449,N_17545);
or U19002 (N_19002,N_16695,N_17969);
and U19003 (N_19003,N_17280,N_17278);
nor U19004 (N_19004,N_17273,N_17197);
and U19005 (N_19005,N_17823,N_17582);
nor U19006 (N_19006,N_16955,N_17783);
or U19007 (N_19007,N_17756,N_16505);
or U19008 (N_19008,N_17849,N_17318);
nand U19009 (N_19009,N_16591,N_16794);
nand U19010 (N_19010,N_16531,N_16681);
and U19011 (N_19011,N_17925,N_17259);
xor U19012 (N_19012,N_17330,N_17059);
or U19013 (N_19013,N_17744,N_16941);
nand U19014 (N_19014,N_16657,N_17507);
or U19015 (N_19015,N_16700,N_16712);
xnor U19016 (N_19016,N_17952,N_17487);
and U19017 (N_19017,N_17097,N_16761);
nand U19018 (N_19018,N_16906,N_16503);
nor U19019 (N_19019,N_17161,N_17950);
nor U19020 (N_19020,N_17156,N_16544);
and U19021 (N_19021,N_17240,N_17981);
or U19022 (N_19022,N_17707,N_17523);
xor U19023 (N_19023,N_16755,N_16832);
nand U19024 (N_19024,N_16993,N_17364);
and U19025 (N_19025,N_17466,N_16821);
or U19026 (N_19026,N_17112,N_17295);
nand U19027 (N_19027,N_16525,N_17181);
or U19028 (N_19028,N_17652,N_16813);
nor U19029 (N_19029,N_16756,N_16673);
nor U19030 (N_19030,N_16931,N_17159);
nor U19031 (N_19031,N_17199,N_17859);
nand U19032 (N_19032,N_16850,N_17493);
and U19033 (N_19033,N_17690,N_17987);
or U19034 (N_19034,N_16754,N_16941);
and U19035 (N_19035,N_17857,N_17291);
nor U19036 (N_19036,N_16932,N_17725);
and U19037 (N_19037,N_17351,N_17388);
or U19038 (N_19038,N_17578,N_17922);
xor U19039 (N_19039,N_17400,N_16891);
nand U19040 (N_19040,N_17160,N_17304);
and U19041 (N_19041,N_16535,N_16760);
and U19042 (N_19042,N_16512,N_17585);
nand U19043 (N_19043,N_17590,N_17546);
xor U19044 (N_19044,N_16920,N_17990);
nand U19045 (N_19045,N_17050,N_16604);
nand U19046 (N_19046,N_17266,N_16955);
and U19047 (N_19047,N_17295,N_17823);
nor U19048 (N_19048,N_17110,N_17433);
or U19049 (N_19049,N_17751,N_17689);
or U19050 (N_19050,N_16706,N_16898);
and U19051 (N_19051,N_16519,N_16662);
and U19052 (N_19052,N_17916,N_17846);
or U19053 (N_19053,N_17377,N_17360);
nor U19054 (N_19054,N_17919,N_16641);
nand U19055 (N_19055,N_17980,N_16615);
nor U19056 (N_19056,N_16857,N_17369);
and U19057 (N_19057,N_17775,N_16592);
nor U19058 (N_19058,N_17112,N_17976);
xor U19059 (N_19059,N_17402,N_16976);
or U19060 (N_19060,N_17880,N_16523);
xor U19061 (N_19061,N_17434,N_17201);
or U19062 (N_19062,N_17697,N_17148);
nand U19063 (N_19063,N_16924,N_17079);
nor U19064 (N_19064,N_16580,N_16803);
or U19065 (N_19065,N_16938,N_17061);
nand U19066 (N_19066,N_17738,N_17812);
or U19067 (N_19067,N_17044,N_16788);
and U19068 (N_19068,N_17904,N_17729);
and U19069 (N_19069,N_16639,N_16515);
nor U19070 (N_19070,N_17354,N_16626);
or U19071 (N_19071,N_16894,N_17674);
nor U19072 (N_19072,N_17383,N_16614);
nor U19073 (N_19073,N_16931,N_17768);
nor U19074 (N_19074,N_17478,N_17007);
xor U19075 (N_19075,N_17219,N_17617);
nor U19076 (N_19076,N_17448,N_17837);
and U19077 (N_19077,N_16881,N_17784);
nor U19078 (N_19078,N_17204,N_17146);
nand U19079 (N_19079,N_17898,N_17816);
nand U19080 (N_19080,N_16789,N_17557);
or U19081 (N_19081,N_17192,N_16938);
nand U19082 (N_19082,N_17716,N_16566);
and U19083 (N_19083,N_16880,N_17262);
xnor U19084 (N_19084,N_17958,N_17205);
and U19085 (N_19085,N_17601,N_16682);
or U19086 (N_19086,N_16854,N_17515);
and U19087 (N_19087,N_17551,N_17356);
xnor U19088 (N_19088,N_17816,N_17894);
and U19089 (N_19089,N_16921,N_17860);
nor U19090 (N_19090,N_16579,N_16802);
or U19091 (N_19091,N_16669,N_16976);
nor U19092 (N_19092,N_17006,N_16983);
nor U19093 (N_19093,N_17837,N_17152);
or U19094 (N_19094,N_17415,N_17648);
nor U19095 (N_19095,N_17589,N_16728);
or U19096 (N_19096,N_17223,N_17605);
nor U19097 (N_19097,N_17489,N_16960);
nor U19098 (N_19098,N_17934,N_17920);
nand U19099 (N_19099,N_17699,N_16767);
nor U19100 (N_19100,N_17560,N_17706);
and U19101 (N_19101,N_16681,N_16539);
nand U19102 (N_19102,N_17245,N_17144);
nand U19103 (N_19103,N_16658,N_17476);
and U19104 (N_19104,N_17898,N_17958);
and U19105 (N_19105,N_17990,N_16865);
xnor U19106 (N_19106,N_17315,N_17961);
or U19107 (N_19107,N_16803,N_17597);
or U19108 (N_19108,N_17610,N_16540);
nand U19109 (N_19109,N_17056,N_17895);
nor U19110 (N_19110,N_17213,N_16538);
or U19111 (N_19111,N_17141,N_16613);
xor U19112 (N_19112,N_17013,N_17197);
or U19113 (N_19113,N_17248,N_17383);
and U19114 (N_19114,N_17770,N_16632);
nand U19115 (N_19115,N_16762,N_17510);
nor U19116 (N_19116,N_17328,N_16773);
or U19117 (N_19117,N_17647,N_16554);
nand U19118 (N_19118,N_17700,N_16779);
and U19119 (N_19119,N_16896,N_16552);
or U19120 (N_19120,N_16887,N_17692);
nand U19121 (N_19121,N_17250,N_17315);
or U19122 (N_19122,N_17780,N_17131);
xnor U19123 (N_19123,N_16752,N_16566);
nor U19124 (N_19124,N_17043,N_17699);
and U19125 (N_19125,N_17059,N_16668);
and U19126 (N_19126,N_16979,N_16958);
and U19127 (N_19127,N_17710,N_16993);
and U19128 (N_19128,N_16506,N_17529);
or U19129 (N_19129,N_17748,N_16969);
nor U19130 (N_19130,N_17596,N_17631);
nand U19131 (N_19131,N_17892,N_17185);
xor U19132 (N_19132,N_17789,N_17386);
xnor U19133 (N_19133,N_17309,N_17797);
nor U19134 (N_19134,N_16726,N_17687);
nand U19135 (N_19135,N_17354,N_16699);
and U19136 (N_19136,N_16698,N_17714);
xnor U19137 (N_19137,N_17120,N_17456);
and U19138 (N_19138,N_16945,N_17719);
or U19139 (N_19139,N_17142,N_17177);
or U19140 (N_19140,N_17553,N_17558);
or U19141 (N_19141,N_17649,N_17349);
nor U19142 (N_19142,N_17804,N_17046);
or U19143 (N_19143,N_17245,N_17051);
nand U19144 (N_19144,N_16553,N_17214);
nand U19145 (N_19145,N_17271,N_16598);
or U19146 (N_19146,N_17268,N_17312);
or U19147 (N_19147,N_17507,N_16836);
xnor U19148 (N_19148,N_17223,N_16722);
nand U19149 (N_19149,N_16848,N_17815);
or U19150 (N_19150,N_17729,N_16909);
nand U19151 (N_19151,N_17415,N_17572);
or U19152 (N_19152,N_16758,N_17508);
xnor U19153 (N_19153,N_17426,N_16941);
nand U19154 (N_19154,N_17168,N_17446);
and U19155 (N_19155,N_17299,N_17131);
xor U19156 (N_19156,N_17519,N_16997);
and U19157 (N_19157,N_16948,N_16592);
and U19158 (N_19158,N_17094,N_17185);
or U19159 (N_19159,N_17104,N_17172);
nand U19160 (N_19160,N_17490,N_17082);
or U19161 (N_19161,N_17815,N_17160);
nor U19162 (N_19162,N_17157,N_17299);
nor U19163 (N_19163,N_17631,N_17143);
and U19164 (N_19164,N_17807,N_17925);
nor U19165 (N_19165,N_17418,N_17319);
or U19166 (N_19166,N_17670,N_17220);
and U19167 (N_19167,N_17496,N_17123);
or U19168 (N_19168,N_17373,N_16855);
nor U19169 (N_19169,N_16508,N_17117);
nor U19170 (N_19170,N_17342,N_16896);
nor U19171 (N_19171,N_17678,N_17172);
and U19172 (N_19172,N_17663,N_16584);
and U19173 (N_19173,N_17056,N_17047);
xor U19174 (N_19174,N_17826,N_17081);
or U19175 (N_19175,N_17403,N_17718);
and U19176 (N_19176,N_17373,N_17914);
or U19177 (N_19177,N_17190,N_17165);
and U19178 (N_19178,N_17354,N_16742);
or U19179 (N_19179,N_16881,N_17628);
xor U19180 (N_19180,N_17936,N_16783);
xnor U19181 (N_19181,N_16749,N_16860);
nor U19182 (N_19182,N_17999,N_17743);
nand U19183 (N_19183,N_16576,N_17018);
nand U19184 (N_19184,N_17595,N_17024);
nand U19185 (N_19185,N_17674,N_17966);
nand U19186 (N_19186,N_17500,N_17358);
and U19187 (N_19187,N_17525,N_17900);
or U19188 (N_19188,N_16858,N_17848);
and U19189 (N_19189,N_17997,N_17078);
xnor U19190 (N_19190,N_17529,N_16990);
or U19191 (N_19191,N_17442,N_17157);
nand U19192 (N_19192,N_17853,N_17477);
xor U19193 (N_19193,N_17675,N_17325);
xor U19194 (N_19194,N_17924,N_17701);
xnor U19195 (N_19195,N_17288,N_17978);
xor U19196 (N_19196,N_16937,N_17722);
or U19197 (N_19197,N_16662,N_17533);
or U19198 (N_19198,N_17954,N_17045);
and U19199 (N_19199,N_17861,N_17745);
nor U19200 (N_19200,N_17031,N_17173);
xnor U19201 (N_19201,N_17004,N_17472);
nand U19202 (N_19202,N_16803,N_17733);
nor U19203 (N_19203,N_17607,N_16717);
xor U19204 (N_19204,N_17875,N_17125);
nor U19205 (N_19205,N_17555,N_16839);
nor U19206 (N_19206,N_16771,N_16654);
and U19207 (N_19207,N_16646,N_17986);
nand U19208 (N_19208,N_17185,N_16696);
nand U19209 (N_19209,N_17815,N_16775);
xnor U19210 (N_19210,N_17374,N_17976);
and U19211 (N_19211,N_17608,N_16540);
nor U19212 (N_19212,N_17630,N_16699);
xor U19213 (N_19213,N_17288,N_17437);
nand U19214 (N_19214,N_16725,N_17560);
xnor U19215 (N_19215,N_17855,N_17804);
xnor U19216 (N_19216,N_16837,N_17519);
nand U19217 (N_19217,N_17945,N_17824);
xnor U19218 (N_19218,N_16703,N_17043);
nand U19219 (N_19219,N_17874,N_16588);
and U19220 (N_19220,N_17840,N_16528);
nor U19221 (N_19221,N_17736,N_16708);
nand U19222 (N_19222,N_17721,N_17415);
and U19223 (N_19223,N_17354,N_16610);
nand U19224 (N_19224,N_16552,N_17210);
and U19225 (N_19225,N_17657,N_16713);
nor U19226 (N_19226,N_16540,N_16551);
or U19227 (N_19227,N_17256,N_17280);
or U19228 (N_19228,N_17236,N_16862);
or U19229 (N_19229,N_16806,N_17072);
and U19230 (N_19230,N_17820,N_17566);
and U19231 (N_19231,N_17476,N_16771);
xor U19232 (N_19232,N_16789,N_17574);
nor U19233 (N_19233,N_16678,N_16628);
nand U19234 (N_19234,N_17610,N_16788);
nor U19235 (N_19235,N_17760,N_16576);
and U19236 (N_19236,N_16747,N_16704);
and U19237 (N_19237,N_16645,N_17384);
and U19238 (N_19238,N_16684,N_16682);
or U19239 (N_19239,N_17539,N_17674);
or U19240 (N_19240,N_17001,N_16636);
nor U19241 (N_19241,N_17267,N_17160);
nor U19242 (N_19242,N_17782,N_16587);
xor U19243 (N_19243,N_17558,N_16679);
xor U19244 (N_19244,N_16803,N_17544);
nand U19245 (N_19245,N_17798,N_17922);
and U19246 (N_19246,N_16718,N_17799);
xnor U19247 (N_19247,N_16703,N_17280);
or U19248 (N_19248,N_16729,N_16682);
nand U19249 (N_19249,N_17116,N_17200);
and U19250 (N_19250,N_16507,N_17528);
nor U19251 (N_19251,N_16881,N_17364);
nor U19252 (N_19252,N_17269,N_16576);
nor U19253 (N_19253,N_17435,N_17595);
or U19254 (N_19254,N_17231,N_17101);
nand U19255 (N_19255,N_16633,N_17939);
and U19256 (N_19256,N_17185,N_16887);
nor U19257 (N_19257,N_17030,N_17128);
and U19258 (N_19258,N_16778,N_17601);
or U19259 (N_19259,N_17652,N_17265);
nand U19260 (N_19260,N_16820,N_17229);
or U19261 (N_19261,N_17742,N_17498);
or U19262 (N_19262,N_17599,N_16520);
nor U19263 (N_19263,N_16614,N_16584);
and U19264 (N_19264,N_17227,N_16563);
nor U19265 (N_19265,N_17764,N_17267);
nor U19266 (N_19266,N_17797,N_17208);
nor U19267 (N_19267,N_17387,N_16589);
nand U19268 (N_19268,N_17299,N_16514);
or U19269 (N_19269,N_16957,N_17482);
xnor U19270 (N_19270,N_17814,N_17355);
or U19271 (N_19271,N_17158,N_17309);
nor U19272 (N_19272,N_17634,N_17400);
nor U19273 (N_19273,N_17502,N_17321);
nor U19274 (N_19274,N_17819,N_16689);
nor U19275 (N_19275,N_16924,N_17189);
nand U19276 (N_19276,N_17938,N_17727);
xnor U19277 (N_19277,N_17671,N_16974);
nand U19278 (N_19278,N_17928,N_16501);
and U19279 (N_19279,N_16680,N_17645);
or U19280 (N_19280,N_17235,N_16891);
and U19281 (N_19281,N_17978,N_17621);
or U19282 (N_19282,N_16513,N_17671);
nor U19283 (N_19283,N_16884,N_16792);
nor U19284 (N_19284,N_17795,N_17246);
xnor U19285 (N_19285,N_17946,N_16653);
and U19286 (N_19286,N_17376,N_17583);
nand U19287 (N_19287,N_17310,N_17562);
xor U19288 (N_19288,N_16715,N_16647);
nor U19289 (N_19289,N_17297,N_16514);
nand U19290 (N_19290,N_16764,N_16797);
xor U19291 (N_19291,N_16870,N_17675);
nor U19292 (N_19292,N_17093,N_17916);
and U19293 (N_19293,N_17983,N_16559);
and U19294 (N_19294,N_17644,N_16571);
xnor U19295 (N_19295,N_17534,N_16664);
nand U19296 (N_19296,N_17087,N_16564);
nand U19297 (N_19297,N_17024,N_17730);
xnor U19298 (N_19298,N_16574,N_17784);
nand U19299 (N_19299,N_16524,N_16727);
nand U19300 (N_19300,N_17845,N_17250);
nand U19301 (N_19301,N_17514,N_17574);
xor U19302 (N_19302,N_16928,N_17501);
nand U19303 (N_19303,N_16988,N_17975);
xor U19304 (N_19304,N_16799,N_16641);
xnor U19305 (N_19305,N_17875,N_17567);
nand U19306 (N_19306,N_17593,N_16898);
nor U19307 (N_19307,N_16801,N_17542);
and U19308 (N_19308,N_17280,N_17955);
nand U19309 (N_19309,N_17703,N_17460);
nand U19310 (N_19310,N_17306,N_17060);
nand U19311 (N_19311,N_17861,N_17800);
and U19312 (N_19312,N_17102,N_17006);
nor U19313 (N_19313,N_17576,N_17529);
nand U19314 (N_19314,N_17760,N_17134);
and U19315 (N_19315,N_17495,N_17385);
nor U19316 (N_19316,N_16849,N_16740);
nor U19317 (N_19317,N_17044,N_16519);
or U19318 (N_19318,N_17750,N_17454);
or U19319 (N_19319,N_16683,N_16518);
nor U19320 (N_19320,N_17373,N_17947);
xor U19321 (N_19321,N_17786,N_17261);
xnor U19322 (N_19322,N_16631,N_17773);
nor U19323 (N_19323,N_17196,N_17829);
xor U19324 (N_19324,N_16765,N_16844);
and U19325 (N_19325,N_17559,N_16845);
nor U19326 (N_19326,N_17842,N_17281);
or U19327 (N_19327,N_16833,N_16926);
or U19328 (N_19328,N_16710,N_17852);
nor U19329 (N_19329,N_17107,N_17608);
nand U19330 (N_19330,N_17670,N_17591);
and U19331 (N_19331,N_16835,N_17109);
nand U19332 (N_19332,N_17063,N_17116);
nor U19333 (N_19333,N_17094,N_17089);
nand U19334 (N_19334,N_17956,N_16811);
nor U19335 (N_19335,N_16578,N_16828);
or U19336 (N_19336,N_17589,N_17779);
and U19337 (N_19337,N_17565,N_16638);
nand U19338 (N_19338,N_17495,N_17580);
xnor U19339 (N_19339,N_17649,N_16673);
and U19340 (N_19340,N_17519,N_17180);
nor U19341 (N_19341,N_17934,N_16758);
or U19342 (N_19342,N_16919,N_17784);
or U19343 (N_19343,N_17011,N_17851);
xor U19344 (N_19344,N_17037,N_16587);
and U19345 (N_19345,N_17007,N_16929);
or U19346 (N_19346,N_17586,N_17479);
and U19347 (N_19347,N_17644,N_17342);
nand U19348 (N_19348,N_17755,N_16526);
and U19349 (N_19349,N_17969,N_17123);
nor U19350 (N_19350,N_17443,N_17000);
xor U19351 (N_19351,N_17004,N_17239);
nand U19352 (N_19352,N_17819,N_17071);
and U19353 (N_19353,N_17253,N_16792);
nor U19354 (N_19354,N_16668,N_17144);
xnor U19355 (N_19355,N_17089,N_16766);
nand U19356 (N_19356,N_17152,N_17882);
xor U19357 (N_19357,N_17490,N_16991);
nand U19358 (N_19358,N_17793,N_16612);
xor U19359 (N_19359,N_17788,N_17052);
nand U19360 (N_19360,N_17769,N_16688);
and U19361 (N_19361,N_17784,N_17418);
or U19362 (N_19362,N_16807,N_16573);
or U19363 (N_19363,N_17748,N_16594);
nor U19364 (N_19364,N_17866,N_17661);
and U19365 (N_19365,N_16833,N_17519);
and U19366 (N_19366,N_16861,N_17666);
nor U19367 (N_19367,N_17643,N_17061);
and U19368 (N_19368,N_17922,N_17972);
or U19369 (N_19369,N_16782,N_17475);
xnor U19370 (N_19370,N_17744,N_17419);
and U19371 (N_19371,N_17970,N_17009);
and U19372 (N_19372,N_17941,N_17195);
or U19373 (N_19373,N_16738,N_16505);
nor U19374 (N_19374,N_16678,N_16627);
and U19375 (N_19375,N_17412,N_17441);
and U19376 (N_19376,N_17353,N_17502);
or U19377 (N_19377,N_17791,N_17020);
or U19378 (N_19378,N_17539,N_16820);
or U19379 (N_19379,N_17736,N_17333);
and U19380 (N_19380,N_17427,N_16610);
and U19381 (N_19381,N_17950,N_17559);
nor U19382 (N_19382,N_17990,N_16820);
and U19383 (N_19383,N_16859,N_16920);
and U19384 (N_19384,N_17613,N_17284);
nand U19385 (N_19385,N_17511,N_17325);
or U19386 (N_19386,N_17637,N_17213);
xor U19387 (N_19387,N_16805,N_17550);
nor U19388 (N_19388,N_17022,N_16718);
nor U19389 (N_19389,N_16648,N_16832);
or U19390 (N_19390,N_16976,N_17239);
or U19391 (N_19391,N_17785,N_17922);
xnor U19392 (N_19392,N_17664,N_17204);
and U19393 (N_19393,N_16531,N_17420);
xnor U19394 (N_19394,N_16787,N_16561);
nor U19395 (N_19395,N_17817,N_17679);
nand U19396 (N_19396,N_17279,N_17030);
or U19397 (N_19397,N_16795,N_17490);
nand U19398 (N_19398,N_17291,N_16775);
and U19399 (N_19399,N_16853,N_17539);
xor U19400 (N_19400,N_17392,N_17788);
nor U19401 (N_19401,N_16780,N_17347);
nor U19402 (N_19402,N_17423,N_16511);
xnor U19403 (N_19403,N_17152,N_17380);
nor U19404 (N_19404,N_17077,N_16960);
nor U19405 (N_19405,N_17489,N_16920);
and U19406 (N_19406,N_17398,N_17216);
nor U19407 (N_19407,N_17272,N_17444);
xnor U19408 (N_19408,N_16619,N_17322);
xor U19409 (N_19409,N_17809,N_17663);
or U19410 (N_19410,N_17854,N_16968);
or U19411 (N_19411,N_17104,N_17588);
nand U19412 (N_19412,N_16993,N_17987);
nand U19413 (N_19413,N_17913,N_16636);
and U19414 (N_19414,N_17584,N_17049);
xnor U19415 (N_19415,N_17304,N_16729);
nor U19416 (N_19416,N_17965,N_16669);
nand U19417 (N_19417,N_17971,N_16713);
or U19418 (N_19418,N_16753,N_17111);
nand U19419 (N_19419,N_16515,N_16806);
nor U19420 (N_19420,N_16782,N_17334);
or U19421 (N_19421,N_16505,N_16546);
xnor U19422 (N_19422,N_16640,N_17427);
xor U19423 (N_19423,N_17447,N_16605);
and U19424 (N_19424,N_16851,N_16556);
nand U19425 (N_19425,N_17300,N_16650);
nor U19426 (N_19426,N_17999,N_17310);
nor U19427 (N_19427,N_16827,N_17896);
and U19428 (N_19428,N_16546,N_17152);
nand U19429 (N_19429,N_17686,N_17519);
or U19430 (N_19430,N_17004,N_17550);
and U19431 (N_19431,N_17435,N_16894);
or U19432 (N_19432,N_17758,N_17117);
or U19433 (N_19433,N_17955,N_16790);
nor U19434 (N_19434,N_17539,N_17296);
and U19435 (N_19435,N_17542,N_16849);
and U19436 (N_19436,N_17909,N_17355);
xor U19437 (N_19437,N_16902,N_17574);
nor U19438 (N_19438,N_16686,N_17449);
and U19439 (N_19439,N_16882,N_17488);
and U19440 (N_19440,N_17430,N_17407);
xnor U19441 (N_19441,N_17476,N_17573);
xnor U19442 (N_19442,N_17709,N_17064);
and U19443 (N_19443,N_17364,N_17605);
nand U19444 (N_19444,N_17184,N_16832);
xor U19445 (N_19445,N_16752,N_17863);
or U19446 (N_19446,N_17038,N_16545);
nand U19447 (N_19447,N_16791,N_17299);
nor U19448 (N_19448,N_17843,N_16705);
xor U19449 (N_19449,N_17903,N_17489);
xnor U19450 (N_19450,N_17294,N_17548);
nand U19451 (N_19451,N_16864,N_17547);
nand U19452 (N_19452,N_16853,N_17958);
or U19453 (N_19453,N_17173,N_16962);
or U19454 (N_19454,N_17067,N_17137);
and U19455 (N_19455,N_16675,N_17527);
xnor U19456 (N_19456,N_17442,N_17712);
or U19457 (N_19457,N_17215,N_17152);
nand U19458 (N_19458,N_17333,N_17389);
and U19459 (N_19459,N_16687,N_17472);
xor U19460 (N_19460,N_17734,N_17949);
xor U19461 (N_19461,N_17368,N_16663);
xor U19462 (N_19462,N_17992,N_17082);
xnor U19463 (N_19463,N_17327,N_16583);
and U19464 (N_19464,N_17761,N_17819);
xnor U19465 (N_19465,N_16816,N_17393);
nand U19466 (N_19466,N_16853,N_17269);
nand U19467 (N_19467,N_16608,N_17473);
nor U19468 (N_19468,N_16732,N_17598);
nand U19469 (N_19469,N_16600,N_17123);
xnor U19470 (N_19470,N_17981,N_17267);
xnor U19471 (N_19471,N_16646,N_17518);
nand U19472 (N_19472,N_16901,N_16992);
or U19473 (N_19473,N_17443,N_17809);
nor U19474 (N_19474,N_17049,N_17529);
or U19475 (N_19475,N_16962,N_17892);
nand U19476 (N_19476,N_16814,N_16630);
or U19477 (N_19477,N_17803,N_16674);
nor U19478 (N_19478,N_17139,N_16592);
or U19479 (N_19479,N_17274,N_16907);
and U19480 (N_19480,N_16702,N_16840);
nand U19481 (N_19481,N_16691,N_17810);
xor U19482 (N_19482,N_16821,N_17100);
nor U19483 (N_19483,N_17688,N_16984);
nor U19484 (N_19484,N_17839,N_17053);
or U19485 (N_19485,N_17345,N_17917);
nand U19486 (N_19486,N_17907,N_17941);
xor U19487 (N_19487,N_17128,N_17896);
xor U19488 (N_19488,N_17620,N_17420);
nor U19489 (N_19489,N_17014,N_17751);
and U19490 (N_19490,N_17508,N_17712);
xor U19491 (N_19491,N_17091,N_16908);
nand U19492 (N_19492,N_17105,N_16987);
or U19493 (N_19493,N_17354,N_17950);
xor U19494 (N_19494,N_17771,N_17139);
xnor U19495 (N_19495,N_16911,N_17155);
nor U19496 (N_19496,N_17866,N_17045);
and U19497 (N_19497,N_17230,N_17245);
and U19498 (N_19498,N_16599,N_16626);
nand U19499 (N_19499,N_16773,N_17934);
and U19500 (N_19500,N_18176,N_19284);
nand U19501 (N_19501,N_19371,N_19403);
or U19502 (N_19502,N_19181,N_19354);
nand U19503 (N_19503,N_19246,N_18458);
or U19504 (N_19504,N_18929,N_19092);
or U19505 (N_19505,N_18477,N_18851);
nor U19506 (N_19506,N_18250,N_19080);
nand U19507 (N_19507,N_18305,N_18094);
xnor U19508 (N_19508,N_19227,N_18597);
nor U19509 (N_19509,N_18718,N_18807);
nand U19510 (N_19510,N_18843,N_18616);
nor U19511 (N_19511,N_18328,N_19245);
and U19512 (N_19512,N_18419,N_18549);
nand U19513 (N_19513,N_18714,N_19226);
nor U19514 (N_19514,N_18375,N_18555);
or U19515 (N_19515,N_18456,N_19074);
nand U19516 (N_19516,N_18591,N_18253);
nor U19517 (N_19517,N_19028,N_18225);
xnor U19518 (N_19518,N_18287,N_18845);
or U19519 (N_19519,N_18904,N_18018);
xor U19520 (N_19520,N_19414,N_18613);
or U19521 (N_19521,N_19203,N_18471);
or U19522 (N_19522,N_18890,N_18234);
and U19523 (N_19523,N_18838,N_18277);
and U19524 (N_19524,N_18876,N_18457);
nor U19525 (N_19525,N_19138,N_19348);
or U19526 (N_19526,N_19094,N_18294);
or U19527 (N_19527,N_18619,N_18697);
or U19528 (N_19528,N_18648,N_18233);
nand U19529 (N_19529,N_18262,N_18667);
and U19530 (N_19530,N_18396,N_19449);
nor U19531 (N_19531,N_18207,N_18196);
or U19532 (N_19532,N_19276,N_18045);
and U19533 (N_19533,N_19438,N_18254);
and U19534 (N_19534,N_19002,N_18126);
and U19535 (N_19535,N_18425,N_19247);
nand U19536 (N_19536,N_19385,N_18765);
nand U19537 (N_19537,N_18923,N_19440);
xnor U19538 (N_19538,N_18461,N_19307);
nor U19539 (N_19539,N_18275,N_18687);
or U19540 (N_19540,N_19287,N_18785);
xor U19541 (N_19541,N_18829,N_19162);
xor U19542 (N_19542,N_18455,N_19019);
or U19543 (N_19543,N_18265,N_18166);
or U19544 (N_19544,N_18654,N_18758);
or U19545 (N_19545,N_18775,N_18139);
nand U19546 (N_19546,N_18053,N_18342);
or U19547 (N_19547,N_18335,N_18147);
nor U19548 (N_19548,N_18823,N_18700);
or U19549 (N_19549,N_19294,N_18332);
xnor U19550 (N_19550,N_19105,N_19353);
and U19551 (N_19551,N_19048,N_18570);
nor U19552 (N_19552,N_18189,N_18232);
nand U19553 (N_19553,N_18681,N_19462);
nor U19554 (N_19554,N_18204,N_18801);
nand U19555 (N_19555,N_19335,N_18727);
or U19556 (N_19556,N_18058,N_19429);
or U19557 (N_19557,N_18793,N_19248);
nand U19558 (N_19558,N_19163,N_18357);
or U19559 (N_19559,N_18214,N_18051);
or U19560 (N_19560,N_18966,N_18003);
or U19561 (N_19561,N_18552,N_18603);
and U19562 (N_19562,N_18329,N_18343);
nand U19563 (N_19563,N_19046,N_18574);
and U19564 (N_19564,N_19321,N_18997);
and U19565 (N_19565,N_18097,N_19278);
nor U19566 (N_19566,N_18208,N_18693);
nor U19567 (N_19567,N_18231,N_18959);
nor U19568 (N_19568,N_18363,N_18739);
xor U19569 (N_19569,N_18142,N_18780);
or U19570 (N_19570,N_18686,N_18792);
and U19571 (N_19571,N_19139,N_19198);
and U19572 (N_19572,N_18649,N_19180);
nand U19573 (N_19573,N_18964,N_18881);
or U19574 (N_19574,N_18917,N_19154);
xor U19575 (N_19575,N_18952,N_18355);
nor U19576 (N_19576,N_18995,N_19086);
or U19577 (N_19577,N_19450,N_18816);
nor U19578 (N_19578,N_18704,N_18398);
xor U19579 (N_19579,N_18941,N_19067);
nor U19580 (N_19580,N_18263,N_18604);
nand U19581 (N_19581,N_18152,N_18651);
nor U19582 (N_19582,N_18559,N_18293);
or U19583 (N_19583,N_18182,N_18599);
or U19584 (N_19584,N_19223,N_18715);
nand U19585 (N_19585,N_19430,N_18230);
nand U19586 (N_19586,N_18537,N_19254);
nand U19587 (N_19587,N_18588,N_19336);
xnor U19588 (N_19588,N_18626,N_19265);
xnor U19589 (N_19589,N_18840,N_18144);
nand U19590 (N_19590,N_19137,N_19295);
nor U19591 (N_19591,N_18089,N_19412);
xnor U19592 (N_19592,N_18406,N_18819);
nand U19593 (N_19593,N_19292,N_19487);
xnor U19594 (N_19594,N_18276,N_18857);
nor U19595 (N_19595,N_18492,N_18728);
xnor U19596 (N_19596,N_19471,N_19442);
xnor U19597 (N_19597,N_18595,N_18578);
and U19598 (N_19598,N_18072,N_18159);
nand U19599 (N_19599,N_18174,N_18005);
nand U19600 (N_19600,N_19083,N_19328);
nand U19601 (N_19601,N_18397,N_18642);
and U19602 (N_19602,N_19061,N_19362);
nand U19603 (N_19603,N_18273,N_18435);
nor U19604 (N_19604,N_19050,N_18988);
nor U19605 (N_19605,N_19087,N_18169);
and U19606 (N_19606,N_18928,N_19457);
xnor U19607 (N_19607,N_18321,N_18405);
nand U19608 (N_19608,N_19179,N_18060);
xnor U19609 (N_19609,N_18082,N_18926);
nor U19610 (N_19610,N_18799,N_18035);
nor U19611 (N_19611,N_18924,N_18865);
nor U19612 (N_19612,N_18307,N_18830);
and U19613 (N_19613,N_18772,N_18659);
xor U19614 (N_19614,N_18490,N_19342);
nand U19615 (N_19615,N_18165,N_19122);
xor U19616 (N_19616,N_19026,N_18194);
and U19617 (N_19617,N_19047,N_18965);
or U19618 (N_19618,N_18576,N_18711);
and U19619 (N_19619,N_18374,N_19463);
nor U19620 (N_19620,N_18245,N_18179);
and U19621 (N_19621,N_18976,N_19402);
nor U19622 (N_19622,N_18701,N_18487);
nand U19623 (N_19623,N_19062,N_19123);
xor U19624 (N_19624,N_18212,N_18021);
and U19625 (N_19625,N_18602,N_18688);
xor U19626 (N_19626,N_19459,N_19044);
and U19627 (N_19627,N_18810,N_18842);
xnor U19628 (N_19628,N_19455,N_18579);
xor U19629 (N_19629,N_19493,N_18480);
and U19630 (N_19630,N_19470,N_19452);
and U19631 (N_19631,N_18643,N_18331);
nor U19632 (N_19632,N_18892,N_18309);
nor U19633 (N_19633,N_18956,N_18408);
or U19634 (N_19634,N_18338,N_18101);
xor U19635 (N_19635,N_18109,N_18114);
xnor U19636 (N_19636,N_18133,N_19021);
nor U19637 (N_19637,N_19421,N_18521);
nand U19638 (N_19638,N_18957,N_18614);
xor U19639 (N_19639,N_18900,N_19182);
or U19640 (N_19640,N_18171,N_19489);
and U19641 (N_19641,N_19060,N_18349);
and U19642 (N_19642,N_19168,N_18107);
or U19643 (N_19643,N_18111,N_18125);
xor U19644 (N_19644,N_18036,N_18726);
nand U19645 (N_19645,N_18695,N_18503);
nor U19646 (N_19646,N_18994,N_18079);
xnor U19647 (N_19647,N_18304,N_18543);
nand U19648 (N_19648,N_18970,N_19127);
and U19649 (N_19649,N_18259,N_18895);
nand U19650 (N_19650,N_18317,N_18783);
or U19651 (N_19651,N_18404,N_19089);
nand U19652 (N_19652,N_18081,N_18962);
and U19653 (N_19653,N_18495,N_18615);
nor U19654 (N_19654,N_19054,N_18380);
xnor U19655 (N_19655,N_18870,N_19055);
and U19656 (N_19656,N_19215,N_19078);
and U19657 (N_19657,N_18824,N_18633);
nor U19658 (N_19658,N_18149,N_19129);
or U19659 (N_19659,N_19184,N_18943);
and U19660 (N_19660,N_18270,N_19386);
nor U19661 (N_19661,N_18912,N_19355);
nand U19662 (N_19662,N_18638,N_18135);
xor U19663 (N_19663,N_18716,N_18175);
xnor U19664 (N_19664,N_18848,N_18157);
xnor U19665 (N_19665,N_19419,N_18907);
nor U19666 (N_19666,N_18562,N_18940);
nand U19667 (N_19667,N_18963,N_18533);
xor U19668 (N_19668,N_19120,N_19024);
and U19669 (N_19669,N_18049,N_18835);
nand U19670 (N_19670,N_18846,N_18439);
or U19671 (N_19671,N_18937,N_19305);
nor U19672 (N_19672,N_19111,N_19316);
and U19673 (N_19673,N_19326,N_18143);
nor U19674 (N_19674,N_19236,N_19464);
nand U19675 (N_19675,N_19498,N_19218);
xor U19676 (N_19676,N_18763,N_19253);
xnor U19677 (N_19677,N_18608,N_18489);
and U19678 (N_19678,N_18430,N_18195);
xor U19679 (N_19679,N_19155,N_18925);
nand U19680 (N_19680,N_19374,N_18589);
and U19681 (N_19681,N_18528,N_18779);
nor U19682 (N_19682,N_18110,N_19368);
xnor U19683 (N_19683,N_18413,N_18764);
xnor U19684 (N_19684,N_19206,N_19043);
or U19685 (N_19685,N_18223,N_18326);
nor U19686 (N_19686,N_19020,N_18510);
nand U19687 (N_19687,N_18462,N_18102);
or U19688 (N_19688,N_18128,N_19389);
nor U19689 (N_19689,N_19159,N_18782);
and U19690 (N_19690,N_18628,N_18736);
nand U19691 (N_19691,N_19369,N_18272);
nand U19692 (N_19692,N_19327,N_18580);
xor U19693 (N_19693,N_19366,N_18600);
xor U19694 (N_19694,N_19103,N_19322);
nor U19695 (N_19695,N_19204,N_19045);
nor U19696 (N_19696,N_18669,N_18771);
and U19697 (N_19697,N_19040,N_18366);
and U19698 (N_19698,N_19499,N_18820);
nor U19699 (N_19699,N_19263,N_18306);
nand U19700 (N_19700,N_18909,N_18703);
and U19701 (N_19701,N_18506,N_19271);
nor U19702 (N_19702,N_18861,N_18444);
nor U19703 (N_19703,N_18889,N_18817);
xnor U19704 (N_19704,N_18505,N_18450);
nand U19705 (N_19705,N_19017,N_18577);
xor U19706 (N_19706,N_19351,N_18414);
and U19707 (N_19707,N_18844,N_18942);
xnor U19708 (N_19708,N_18327,N_18369);
xor U19709 (N_19709,N_18787,N_18971);
xnor U19710 (N_19710,N_18394,N_18958);
nor U19711 (N_19711,N_18446,N_18993);
and U19712 (N_19712,N_18516,N_18808);
and U19713 (N_19713,N_18502,N_18227);
xor U19714 (N_19714,N_19004,N_18421);
nand U19715 (N_19715,N_18518,N_18316);
nor U19716 (N_19716,N_18154,N_18690);
or U19717 (N_19717,N_19082,N_19077);
nor U19718 (N_19718,N_18884,N_18496);
nand U19719 (N_19719,N_19497,N_19121);
nand U19720 (N_19720,N_18407,N_18044);
xnor U19721 (N_19721,N_18888,N_19210);
xnor U19722 (N_19722,N_18762,N_18008);
or U19723 (N_19723,N_18809,N_18735);
or U19724 (N_19724,N_19071,N_18353);
and U19725 (N_19725,N_19437,N_18065);
xor U19726 (N_19726,N_19041,N_18948);
and U19727 (N_19727,N_18730,N_19480);
xnor U19728 (N_19728,N_19349,N_18826);
nor U19729 (N_19729,N_18371,N_18300);
and U19730 (N_19730,N_19290,N_19474);
nand U19731 (N_19731,N_18443,N_19289);
or U19732 (N_19732,N_18584,N_18757);
xnor U19733 (N_19733,N_18136,N_19436);
and U19734 (N_19734,N_18850,N_18754);
nor U19735 (N_19735,N_18393,N_19214);
nor U19736 (N_19736,N_18662,N_18163);
and U19737 (N_19737,N_18977,N_19051);
nor U19738 (N_19738,N_18409,N_19472);
and U19739 (N_19739,N_18281,N_18705);
nand U19740 (N_19740,N_19352,N_18781);
or U19741 (N_19741,N_18575,N_18547);
nor U19742 (N_19742,N_18680,N_19264);
xor U19743 (N_19743,N_19257,N_18238);
nand U19744 (N_19744,N_18665,N_18512);
and U19745 (N_19745,N_18655,N_19230);
nor U19746 (N_19746,N_18198,N_18348);
nand U19747 (N_19747,N_18975,N_18702);
xnor U19748 (N_19748,N_18864,N_19022);
xnor U19749 (N_19749,N_18180,N_18949);
nand U19750 (N_19750,N_18322,N_18145);
or U19751 (N_19751,N_18067,N_19364);
or U19752 (N_19752,N_18791,N_18517);
and U19753 (N_19753,N_19454,N_18488);
nor U19754 (N_19754,N_19484,N_19458);
nor U19755 (N_19755,N_19208,N_19173);
or U19756 (N_19756,N_19134,N_18837);
nor U19757 (N_19757,N_18085,N_19239);
or U19758 (N_19758,N_19310,N_18137);
and U19759 (N_19759,N_18183,N_19073);
nor U19760 (N_19760,N_18386,N_18034);
nand U19761 (N_19761,N_18310,N_18811);
nand U19762 (N_19762,N_18919,N_19379);
or U19763 (N_19763,N_18001,N_19104);
nor U19764 (N_19764,N_18664,N_19191);
nor U19765 (N_19765,N_19390,N_18161);
and U19766 (N_19766,N_19197,N_18950);
nor U19767 (N_19767,N_18531,N_18295);
or U19768 (N_19768,N_19394,N_18216);
nor U19769 (N_19769,N_18241,N_18084);
nor U19770 (N_19770,N_18077,N_18676);
or U19771 (N_19771,N_18151,N_18563);
xnor U19772 (N_19772,N_19220,N_18637);
or U19773 (N_19773,N_18747,N_18382);
nand U19774 (N_19774,N_18813,N_18346);
nand U19775 (N_19775,N_18869,N_19075);
nand U19776 (N_19776,N_18160,N_18285);
xor U19777 (N_19777,N_18646,N_19494);
nand U19778 (N_19778,N_18769,N_18596);
nand U19779 (N_19779,N_18894,N_19177);
or U19780 (N_19780,N_19126,N_19076);
nor U19781 (N_19781,N_19415,N_19387);
nor U19782 (N_19782,N_18478,N_18539);
and U19783 (N_19783,N_18029,N_18678);
nor U19784 (N_19784,N_18090,N_18377);
nor U19785 (N_19785,N_18028,N_18939);
or U19786 (N_19786,N_19166,N_18789);
nand U19787 (N_19787,N_18056,N_18699);
or U19788 (N_19788,N_19275,N_18587);
xnor U19789 (N_19789,N_19216,N_19240);
and U19790 (N_19790,N_18542,N_18199);
xor U19791 (N_19791,N_18571,N_18150);
xor U19792 (N_19792,N_19217,N_18607);
nand U19793 (N_19793,N_18432,N_19003);
and U19794 (N_19794,N_19016,N_18636);
xor U19795 (N_19795,N_18087,N_18930);
nand U19796 (N_19796,N_19341,N_18124);
nor U19797 (N_19797,N_18330,N_18979);
nand U19798 (N_19798,N_18205,N_19229);
nand U19799 (N_19799,N_18451,N_19426);
or U19800 (N_19800,N_19400,N_18069);
nand U19801 (N_19801,N_18558,N_19378);
and U19802 (N_19802,N_19033,N_18656);
xor U19803 (N_19803,N_18311,N_19135);
xor U19804 (N_19804,N_18709,N_19145);
nor U19805 (N_19805,N_19444,N_19178);
or U19806 (N_19806,N_18141,N_18960);
or U19807 (N_19807,N_18376,N_18268);
nor U19808 (N_19808,N_18298,N_18743);
and U19809 (N_19809,N_19252,N_18751);
nor U19810 (N_19810,N_18668,N_18383);
nand U19811 (N_19811,N_18491,N_19189);
nor U19812 (N_19812,N_18913,N_19404);
xor U19813 (N_19813,N_19286,N_18724);
nor U19814 (N_19814,N_18220,N_19491);
or U19815 (N_19815,N_18209,N_18692);
nand U19816 (N_19816,N_18732,N_18256);
and U19817 (N_19817,N_18798,N_18998);
nand U19818 (N_19818,N_18373,N_18368);
nand U19819 (N_19819,N_18748,N_19143);
and U19820 (N_19820,N_19338,N_18610);
nor U19821 (N_19821,N_18352,N_18514);
nand U19822 (N_19822,N_18855,N_18802);
nand U19823 (N_19823,N_18178,N_18803);
xor U19824 (N_19824,N_18422,N_19408);
nor U19825 (N_19825,N_18741,N_18236);
or U19826 (N_19826,N_18459,N_18301);
and U19827 (N_19827,N_18706,N_19288);
nor U19828 (N_19828,N_18206,N_18117);
nand U19829 (N_19829,N_18025,N_18266);
xnor U19830 (N_19830,N_19317,N_18553);
xnor U19831 (N_19831,N_18671,N_18887);
xnor U19832 (N_19832,N_18027,N_18370);
xnor U19833 (N_19833,N_18786,N_18974);
xnor U19834 (N_19834,N_19243,N_19432);
nor U19835 (N_19835,N_18550,N_19015);
and U19836 (N_19836,N_19175,N_19030);
nor U19837 (N_19837,N_19232,N_18916);
nor U19838 (N_19838,N_18847,N_18752);
xnor U19839 (N_19839,N_18658,N_18410);
xor U19840 (N_19840,N_18011,N_18063);
nand U19841 (N_19841,N_19152,N_18200);
or U19842 (N_19842,N_18184,N_19234);
xnor U19843 (N_19843,N_18713,N_18629);
nor U19844 (N_19844,N_18350,N_18815);
and U19845 (N_19845,N_19113,N_19311);
or U19846 (N_19846,N_19283,N_19202);
nor U19847 (N_19847,N_19225,N_18622);
or U19848 (N_19848,N_18486,N_18663);
or U19849 (N_19849,N_18454,N_18479);
xnor U19850 (N_19850,N_18841,N_19468);
nor U19851 (N_19851,N_19150,N_18080);
nand U19852 (N_19852,N_19029,N_18945);
nor U19853 (N_19853,N_18426,N_18291);
xor U19854 (N_19854,N_18523,N_18362);
nand U19855 (N_19855,N_19270,N_19382);
nand U19856 (N_19856,N_18684,N_18391);
nor U19857 (N_19857,N_18903,N_19381);
xnor U19858 (N_19858,N_19256,N_19488);
or U19859 (N_19859,N_19274,N_18914);
nor U19860 (N_19860,N_18379,N_19279);
and U19861 (N_19861,N_19224,N_19237);
nor U19862 (N_19862,N_19081,N_18719);
nand U19863 (N_19863,N_18606,N_18593);
xor U19864 (N_19864,N_18416,N_19034);
and U19865 (N_19865,N_19465,N_19099);
and U19866 (N_19866,N_19141,N_18221);
xor U19867 (N_19867,N_19096,N_18155);
nor U19868 (N_19868,N_18336,N_18991);
nand U19869 (N_19869,N_18901,N_19291);
xor U19870 (N_19870,N_18134,N_18873);
xnor U19871 (N_19871,N_19065,N_18113);
or U19872 (N_19872,N_18548,N_19193);
nand U19873 (N_19873,N_19435,N_19142);
nand U19874 (N_19874,N_19388,N_18640);
xnor U19875 (N_19875,N_18123,N_19124);
and U19876 (N_19876,N_18465,N_18038);
and U19877 (N_19877,N_18341,N_18712);
xor U19878 (N_19878,N_18269,N_18777);
or U19879 (N_19879,N_18770,N_18832);
and U19880 (N_19880,N_18645,N_18260);
and U19881 (N_19881,N_18438,N_18282);
and U19882 (N_19882,N_18592,N_19188);
and U19883 (N_19883,N_18922,N_18698);
or U19884 (N_19884,N_19300,N_19157);
nor U19885 (N_19885,N_18583,N_18303);
or U19886 (N_19886,N_19413,N_19428);
or U19887 (N_19887,N_18140,N_18883);
and U19888 (N_19888,N_18825,N_18598);
nor U19889 (N_19889,N_18527,N_19106);
nor U19890 (N_19890,N_19280,N_18635);
and U19891 (N_19891,N_19007,N_18239);
or U19892 (N_19892,N_19091,N_18433);
nor U19893 (N_19893,N_19068,N_19012);
xnor U19894 (N_19894,N_18116,N_19063);
or U19895 (N_19895,N_18390,N_18611);
or U19896 (N_19896,N_19431,N_18417);
xnor U19897 (N_19897,N_19446,N_19130);
and U19898 (N_19898,N_19231,N_19466);
nand U19899 (N_19899,N_18696,N_18532);
nand U19900 (N_19900,N_18955,N_18340);
and U19901 (N_19901,N_19360,N_18292);
and U19902 (N_19902,N_18566,N_18138);
or U19903 (N_19903,N_18530,N_18014);
or U19904 (N_19904,N_19417,N_18749);
nand U19905 (N_19905,N_18315,N_19395);
nand U19906 (N_19906,N_18672,N_18880);
nand U19907 (N_19907,N_19377,N_18882);
or U19908 (N_19908,N_19476,N_18745);
or U19909 (N_19909,N_18037,N_18334);
nor U19910 (N_19910,N_19014,N_18657);
nor U19911 (N_19911,N_18674,N_18852);
or U19912 (N_19912,N_19461,N_18573);
nor U19913 (N_19913,N_19170,N_18720);
and U19914 (N_19914,N_18774,N_18794);
nand U19915 (N_19915,N_18467,N_18359);
xor U19916 (N_19916,N_18630,N_18015);
xor U19917 (N_19917,N_18188,N_19058);
xnor U19918 (N_19918,N_18240,N_18388);
nor U19919 (N_19919,N_19221,N_18946);
xnor U19920 (N_19920,N_18384,N_19042);
nor U19921 (N_19921,N_18318,N_18218);
nand U19922 (N_19922,N_18022,N_18984);
or U19923 (N_19923,N_18908,N_18429);
nor U19924 (N_19924,N_19314,N_18981);
and U19925 (N_19925,N_19031,N_19085);
or U19926 (N_19926,N_19219,N_19315);
and U19927 (N_19927,N_19114,N_18224);
nor U19928 (N_19928,N_18076,N_18800);
or U19929 (N_19929,N_18000,N_18731);
or U19930 (N_19930,N_19392,N_18644);
nand U19931 (N_19931,N_18954,N_18511);
or U19932 (N_19932,N_18653,N_19433);
or U19933 (N_19933,N_19161,N_18290);
xnor U19934 (N_19934,N_18814,N_18392);
nor U19935 (N_19935,N_18729,N_18627);
or U19936 (N_19936,N_19424,N_19273);
and U19937 (N_19937,N_19151,N_19319);
xnor U19938 (N_19938,N_18009,N_19205);
xor U19939 (N_19939,N_19235,N_18560);
and U19940 (N_19940,N_18100,N_18248);
and U19941 (N_19941,N_19496,N_19090);
nor U19942 (N_19942,N_18046,N_18938);
nor U19943 (N_19943,N_19095,N_18968);
xnor U19944 (N_19944,N_18324,N_18474);
or U19945 (N_19945,N_18557,N_19456);
nand U19946 (N_19946,N_18121,N_18561);
nand U19947 (N_19947,N_19345,N_18091);
nor U19948 (N_19948,N_18618,N_18059);
xor U19949 (N_19949,N_19267,N_18401);
or U19950 (N_19950,N_18202,N_18725);
nor U19951 (N_19951,N_18278,N_19153);
and U19952 (N_19952,N_19027,N_19298);
xor U19953 (N_19953,N_19448,N_18185);
and U19954 (N_19954,N_18052,N_18524);
nand U19955 (N_19955,N_19006,N_18428);
and U19956 (N_19956,N_18190,N_18460);
nand U19957 (N_19957,N_18086,N_19358);
nand U19958 (N_19958,N_18906,N_18337);
or U19959 (N_19959,N_18918,N_19405);
and U19960 (N_19960,N_18083,N_18915);
nand U19961 (N_19961,N_19434,N_19025);
and U19962 (N_19962,N_18828,N_18319);
or U19963 (N_19963,N_18581,N_18675);
or U19964 (N_19964,N_19084,N_18609);
nor U19965 (N_19965,N_19406,N_18466);
nor U19966 (N_19966,N_19482,N_19196);
and U19967 (N_19967,N_19346,N_18118);
nand U19968 (N_19968,N_18132,N_19399);
nand U19969 (N_19969,N_18017,N_19250);
xor U19970 (N_19970,N_18546,N_18283);
nor U19971 (N_19971,N_18879,N_18257);
and U19972 (N_19972,N_18481,N_18361);
and U19973 (N_19973,N_18264,N_19109);
or U19974 (N_19974,N_19119,N_19148);
and U19975 (N_19975,N_18594,N_19486);
nand U19976 (N_19976,N_18862,N_18367);
nand U19977 (N_19977,N_19393,N_18007);
xnor U19978 (N_19978,N_18911,N_18891);
nand U19979 (N_19979,N_19479,N_19110);
xnor U19980 (N_19980,N_19383,N_18740);
nand U19981 (N_19981,N_18267,N_18866);
and U19982 (N_19982,N_19475,N_19309);
or U19983 (N_19983,N_18279,N_18859);
xor U19984 (N_19984,N_18875,N_19116);
nor U19985 (N_19985,N_19183,N_18839);
nor U19986 (N_19986,N_18469,N_18192);
xor U19987 (N_19987,N_19115,N_19133);
and U19988 (N_19988,N_18565,N_18812);
nor U19989 (N_19989,N_19222,N_18156);
nand U19990 (N_19990,N_18119,N_19451);
nand U19991 (N_19991,N_18673,N_18016);
xnor U19992 (N_19992,N_19066,N_19233);
xnor U19993 (N_19993,N_18484,N_19213);
nand U19994 (N_19994,N_18494,N_19107);
and U19995 (N_19995,N_19485,N_19477);
and U19996 (N_19996,N_18858,N_18987);
nor U19997 (N_19997,N_18742,N_18605);
and U19998 (N_19998,N_18288,N_18737);
nand U19999 (N_19999,N_19190,N_19422);
xor U20000 (N_20000,N_18972,N_19258);
or U20001 (N_20001,N_19036,N_18723);
nand U20002 (N_20002,N_19323,N_19490);
nand U20003 (N_20003,N_18493,N_18447);
xor U20004 (N_20004,N_18834,N_19423);
nor U20005 (N_20005,N_18041,N_19000);
xor U20006 (N_20006,N_19340,N_18586);
or U20007 (N_20007,N_18641,N_18186);
xnor U20008 (N_20008,N_18483,N_18980);
and U20009 (N_20009,N_19251,N_18042);
or U20010 (N_20010,N_19411,N_18222);
and U20011 (N_20011,N_18098,N_19195);
xor U20012 (N_20012,N_18536,N_19318);
or U20013 (N_20013,N_18677,N_18755);
and U20014 (N_20014,N_18020,N_19339);
nor U20015 (N_20015,N_19409,N_18070);
or U20016 (N_20016,N_18768,N_18026);
xor U20017 (N_20017,N_18078,N_19144);
or U20018 (N_20018,N_18402,N_18164);
and U20019 (N_20019,N_19070,N_19427);
xor U20020 (N_20020,N_18243,N_19131);
or U20021 (N_20021,N_19268,N_18796);
nor U20022 (N_20022,N_18682,N_18242);
xnor U20023 (N_20023,N_18953,N_18215);
nand U20024 (N_20024,N_19416,N_18030);
xnor U20025 (N_20025,N_18612,N_19136);
and U20026 (N_20026,N_19097,N_19334);
and U20027 (N_20027,N_19420,N_18766);
nand U20028 (N_20028,N_18255,N_19165);
nor U20029 (N_20029,N_18973,N_18389);
xnor U20030 (N_20030,N_18985,N_18071);
xor U20031 (N_20031,N_19344,N_18624);
nor U20032 (N_20032,N_19469,N_18228);
xnor U20033 (N_20033,N_18936,N_18515);
xor U20034 (N_20034,N_18898,N_19302);
nor U20035 (N_20035,N_18284,N_18167);
or U20036 (N_20036,N_18130,N_18010);
and U20037 (N_20037,N_18499,N_18299);
xor U20038 (N_20038,N_18187,N_18177);
nand U20039 (N_20039,N_18023,N_18685);
xor U20040 (N_20040,N_18744,N_18717);
xnor U20041 (N_20041,N_19255,N_18385);
and U20042 (N_20042,N_18652,N_18431);
or U20043 (N_20043,N_19156,N_18854);
xnor U20044 (N_20044,N_18068,N_19052);
nand U20045 (N_20045,N_19212,N_18797);
or U20046 (N_20046,N_18399,N_19008);
nand U20047 (N_20047,N_18933,N_19039);
nand U20048 (N_20048,N_19118,N_18364);
or U20049 (N_20049,N_19200,N_18449);
xor U20050 (N_20050,N_18127,N_19376);
or U20051 (N_20051,N_19359,N_18064);
xnor U20052 (N_20052,N_18170,N_19102);
or U20053 (N_20053,N_19332,N_18043);
nand U20054 (N_20054,N_18424,N_18115);
nand U20055 (N_20055,N_19396,N_18520);
nand U20056 (N_20056,N_19308,N_19439);
nand U20057 (N_20057,N_19035,N_18778);
and U20058 (N_20058,N_18345,N_19088);
nand U20059 (N_20059,N_18012,N_18585);
or U20060 (N_20060,N_18513,N_18297);
and U20061 (N_20061,N_18572,N_18497);
or U20062 (N_20062,N_18931,N_18210);
or U20063 (N_20063,N_18921,N_18252);
or U20064 (N_20064,N_18271,N_18258);
or U20065 (N_20065,N_19373,N_18333);
nand U20066 (N_20066,N_19303,N_18867);
xnor U20067 (N_20067,N_18554,N_18464);
or U20068 (N_20068,N_18582,N_18509);
xnor U20069 (N_20069,N_18289,N_19164);
xor U20070 (N_20070,N_18411,N_18463);
and U20071 (N_20071,N_18986,N_18280);
and U20072 (N_20072,N_18173,N_18440);
and U20073 (N_20073,N_19117,N_18358);
nand U20074 (N_20074,N_18634,N_18897);
nand U20075 (N_20075,N_18013,N_18773);
nand U20076 (N_20076,N_19407,N_19418);
nor U20077 (N_20077,N_19325,N_19069);
xor U20078 (N_20078,N_18761,N_18750);
and U20079 (N_20079,N_18670,N_18286);
and U20080 (N_20080,N_18871,N_18525);
xor U20081 (N_20081,N_18193,N_19192);
nand U20082 (N_20082,N_18831,N_19112);
nand U20083 (N_20083,N_18365,N_18877);
or U20084 (N_20084,N_19356,N_18302);
or U20085 (N_20085,N_18162,N_19285);
xor U20086 (N_20086,N_18526,N_18788);
nor U20087 (N_20087,N_18476,N_18733);
nor U20088 (N_20088,N_18849,N_18418);
nand U20089 (N_20089,N_18853,N_18339);
xnor U20090 (N_20090,N_18006,N_19032);
nor U20091 (N_20091,N_18104,N_18093);
or U20092 (N_20092,N_19473,N_19001);
and U20093 (N_20093,N_18896,N_18689);
nor U20094 (N_20094,N_19492,N_19158);
nand U20095 (N_20095,N_18568,N_18040);
xnor U20096 (N_20096,N_19391,N_18448);
or U20097 (N_20097,N_18103,N_19333);
and U20098 (N_20098,N_18999,N_18694);
nor U20099 (N_20099,N_18387,N_18099);
xor U20100 (N_20100,N_18400,N_19259);
or U20101 (N_20101,N_19445,N_19169);
xnor U20102 (N_20102,N_18856,N_18621);
and U20103 (N_20103,N_19160,N_19372);
nor U20104 (N_20104,N_18660,N_18445);
nand U20105 (N_20105,N_18529,N_18590);
nand U20106 (N_20106,N_18061,N_18498);
and U20107 (N_20107,N_19064,N_19010);
nor U20108 (N_20108,N_19363,N_18899);
nand U20109 (N_20109,N_19301,N_18092);
or U20110 (N_20110,N_18217,N_19023);
xor U20111 (N_20111,N_19098,N_18538);
nand U20112 (N_20112,N_18541,N_19370);
nor U20113 (N_20113,N_18564,N_18002);
nand U20114 (N_20114,N_18874,N_19261);
nand U20115 (N_20115,N_19005,N_18623);
and U20116 (N_20116,N_19296,N_18095);
or U20117 (N_20117,N_19478,N_18325);
nor U20118 (N_20118,N_18033,N_19447);
xnor U20119 (N_20119,N_18482,N_18434);
and U20120 (N_20120,N_18201,N_19441);
and U20121 (N_20121,N_19304,N_19176);
nand U20122 (N_20122,N_18666,N_18122);
and U20123 (N_20123,N_18996,N_19282);
xnor U20124 (N_20124,N_19128,N_18055);
or U20125 (N_20125,N_18863,N_18213);
xor U20126 (N_20126,N_18760,N_18540);
or U20127 (N_20127,N_19186,N_18191);
xnor U20128 (N_20128,N_19329,N_18031);
and U20129 (N_20129,N_19211,N_19361);
xnor U20130 (N_20130,N_18632,N_18108);
and U20131 (N_20131,N_18990,N_19194);
and U20132 (N_20132,N_18146,N_18934);
or U20133 (N_20133,N_19228,N_18039);
and U20134 (N_20134,N_18244,N_18522);
xor U20135 (N_20135,N_18910,N_19331);
and U20136 (N_20136,N_19167,N_19320);
or U20137 (N_20137,N_18544,N_18650);
nor U20138 (N_20138,N_19347,N_19330);
nor U20139 (N_20139,N_19266,N_18203);
and U20140 (N_20140,N_18312,N_19313);
and U20141 (N_20141,N_18567,N_19241);
and U20142 (N_20142,N_18120,N_18237);
nor U20143 (N_20143,N_19460,N_18683);
and U20144 (N_20144,N_18967,N_18776);
and U20145 (N_20145,N_19209,N_18308);
nor U20146 (N_20146,N_18982,N_18485);
and U20147 (N_20147,N_19049,N_18235);
and U20148 (N_20148,N_19140,N_19108);
nor U20149 (N_20149,N_18738,N_18969);
nor U20150 (N_20150,N_19059,N_19009);
or U20151 (N_20151,N_18148,N_18872);
nor U20152 (N_20152,N_18868,N_18075);
and U20153 (N_20153,N_19201,N_18246);
or U20154 (N_20154,N_19100,N_19013);
or U20155 (N_20155,N_18886,N_19187);
nor U20156 (N_20156,N_19357,N_18992);
and U20157 (N_20157,N_18679,N_18032);
nand U20158 (N_20158,N_18617,N_18452);
or U20159 (N_20159,N_18818,N_18153);
or U20160 (N_20160,N_18470,N_19185);
nor U20161 (N_20161,N_18197,N_18806);
nor U20162 (N_20162,N_18131,N_19101);
nor U20163 (N_20163,N_18468,N_19367);
nor U20164 (N_20164,N_18249,N_18734);
or U20165 (N_20165,N_18378,N_18112);
nand U20166 (N_20166,N_19350,N_18403);
nand U20167 (N_20167,N_18983,N_19149);
or U20168 (N_20168,N_18944,N_18759);
or U20169 (N_20169,N_18722,N_18074);
and U20170 (N_20170,N_19238,N_18902);
xor U20171 (N_20171,N_18710,N_18473);
nor U20172 (N_20172,N_18631,N_18795);
nand U20173 (N_20173,N_19281,N_18229);
nor U20174 (N_20174,N_18320,N_18181);
or U20175 (N_20175,N_18639,N_18519);
nand U20176 (N_20176,N_19018,N_19380);
nand U20177 (N_20177,N_18932,N_18219);
and U20178 (N_20178,N_18504,N_18314);
or U20179 (N_20179,N_19132,N_18707);
nand U20180 (N_20180,N_18822,N_18247);
nor U20181 (N_20181,N_18351,N_18211);
and U20182 (N_20182,N_18048,N_18927);
or U20183 (N_20183,N_19244,N_19146);
nor U20184 (N_20184,N_19481,N_19072);
and U20185 (N_20185,N_18261,N_18535);
nor U20186 (N_20186,N_18381,N_18556);
nand U20187 (N_20187,N_18893,N_18821);
and U20188 (N_20188,N_18545,N_19125);
nor U20189 (N_20189,N_18978,N_19053);
xor U20190 (N_20190,N_18790,N_19172);
or U20191 (N_20191,N_19337,N_18441);
or U20192 (N_20192,N_19312,N_19299);
nand U20193 (N_20193,N_18753,N_18073);
nand U20194 (N_20194,N_18708,N_18804);
nand U20195 (N_20195,N_18647,N_18054);
nor U20196 (N_20196,N_18168,N_18313);
nand U20197 (N_20197,N_18827,N_18620);
nor U20198 (N_20198,N_18356,N_19401);
and U20199 (N_20199,N_19242,N_18057);
nor U20200 (N_20200,N_18296,N_19443);
nand U20201 (N_20201,N_18062,N_19453);
xnor U20202 (N_20202,N_18423,N_18004);
or U20203 (N_20203,N_18442,N_18415);
or U20204 (N_20204,N_18360,N_19093);
and U20205 (N_20205,N_18019,N_18475);
and U20206 (N_20206,N_18691,N_19272);
nand U20207 (N_20207,N_18047,N_18105);
nor U20208 (N_20208,N_18833,N_18569);
and U20209 (N_20209,N_19199,N_19306);
and U20210 (N_20210,N_18951,N_18508);
nor U20211 (N_20211,N_18507,N_18106);
nor U20212 (N_20212,N_18251,N_19293);
and U20213 (N_20213,N_18437,N_18436);
xor U20214 (N_20214,N_19249,N_18323);
and U20215 (N_20215,N_18534,N_18961);
nor U20216 (N_20216,N_18805,N_18274);
nor U20217 (N_20217,N_18947,N_18551);
nand U20218 (N_20218,N_18129,N_19011);
or U20219 (N_20219,N_19260,N_18096);
or U20220 (N_20220,N_18920,N_18395);
and U20221 (N_20221,N_18412,N_19467);
xnor U20222 (N_20222,N_18885,N_19262);
or U20223 (N_20223,N_18066,N_18088);
nor U20224 (N_20224,N_19397,N_18905);
or U20225 (N_20225,N_18784,N_19425);
xor U20226 (N_20226,N_19057,N_19147);
or U20227 (N_20227,N_19495,N_18661);
nor U20228 (N_20228,N_18767,N_19398);
nand U20229 (N_20229,N_18756,N_19079);
or U20230 (N_20230,N_18172,N_18354);
nor U20231 (N_20231,N_19269,N_18601);
or U20232 (N_20232,N_19171,N_18836);
and U20233 (N_20233,N_18501,N_19384);
nand U20234 (N_20234,N_18347,N_18860);
nand U20235 (N_20235,N_18746,N_19324);
and U20236 (N_20236,N_19297,N_18935);
xnor U20237 (N_20237,N_18989,N_19483);
nand U20238 (N_20238,N_18427,N_18625);
or U20239 (N_20239,N_19038,N_19343);
nor U20240 (N_20240,N_19277,N_18372);
xor U20241 (N_20241,N_19037,N_18472);
xor U20242 (N_20242,N_18344,N_18226);
xnor U20243 (N_20243,N_19207,N_18453);
and U20244 (N_20244,N_18721,N_19410);
nor U20245 (N_20245,N_18500,N_18024);
xor U20246 (N_20246,N_18878,N_18050);
nor U20247 (N_20247,N_18420,N_19056);
nor U20248 (N_20248,N_19365,N_18158);
nor U20249 (N_20249,N_19174,N_19375);
or U20250 (N_20250,N_19458,N_18423);
xnor U20251 (N_20251,N_18216,N_18759);
and U20252 (N_20252,N_18870,N_19207);
xnor U20253 (N_20253,N_18151,N_18979);
or U20254 (N_20254,N_18827,N_18146);
or U20255 (N_20255,N_18408,N_18213);
or U20256 (N_20256,N_19266,N_19179);
or U20257 (N_20257,N_18381,N_19025);
xor U20258 (N_20258,N_18849,N_18899);
nand U20259 (N_20259,N_19183,N_18117);
xnor U20260 (N_20260,N_18714,N_19460);
or U20261 (N_20261,N_19013,N_18158);
nand U20262 (N_20262,N_18036,N_19214);
nand U20263 (N_20263,N_18438,N_19014);
xnor U20264 (N_20264,N_18816,N_18570);
xnor U20265 (N_20265,N_19086,N_18959);
or U20266 (N_20266,N_18664,N_18887);
or U20267 (N_20267,N_18855,N_18666);
xnor U20268 (N_20268,N_18005,N_18064);
nand U20269 (N_20269,N_18876,N_18091);
or U20270 (N_20270,N_18036,N_18652);
nand U20271 (N_20271,N_18957,N_19467);
xnor U20272 (N_20272,N_18545,N_18730);
or U20273 (N_20273,N_18133,N_18122);
nand U20274 (N_20274,N_18411,N_18999);
nor U20275 (N_20275,N_18174,N_18935);
and U20276 (N_20276,N_19351,N_18917);
and U20277 (N_20277,N_18600,N_18382);
and U20278 (N_20278,N_19287,N_19383);
and U20279 (N_20279,N_18320,N_18364);
nor U20280 (N_20280,N_18799,N_18229);
nor U20281 (N_20281,N_19245,N_18531);
nand U20282 (N_20282,N_19154,N_18131);
nand U20283 (N_20283,N_18360,N_18283);
and U20284 (N_20284,N_19312,N_18724);
or U20285 (N_20285,N_19092,N_19364);
or U20286 (N_20286,N_19429,N_19414);
and U20287 (N_20287,N_18892,N_18938);
nor U20288 (N_20288,N_18136,N_18476);
nand U20289 (N_20289,N_19206,N_19008);
and U20290 (N_20290,N_18420,N_18962);
and U20291 (N_20291,N_18071,N_18069);
nand U20292 (N_20292,N_18842,N_19191);
xnor U20293 (N_20293,N_18811,N_18661);
and U20294 (N_20294,N_18731,N_19310);
nor U20295 (N_20295,N_19168,N_19323);
and U20296 (N_20296,N_18678,N_18961);
nor U20297 (N_20297,N_18808,N_18648);
xnor U20298 (N_20298,N_18720,N_18820);
xor U20299 (N_20299,N_19143,N_19462);
or U20300 (N_20300,N_19486,N_18760);
nand U20301 (N_20301,N_18762,N_19004);
xor U20302 (N_20302,N_19280,N_18186);
xnor U20303 (N_20303,N_19299,N_18662);
nor U20304 (N_20304,N_19015,N_18109);
nand U20305 (N_20305,N_18111,N_18344);
xor U20306 (N_20306,N_18802,N_18051);
nand U20307 (N_20307,N_18187,N_18348);
xnor U20308 (N_20308,N_18802,N_19230);
nor U20309 (N_20309,N_18193,N_18682);
or U20310 (N_20310,N_18924,N_18556);
nand U20311 (N_20311,N_18167,N_18080);
xor U20312 (N_20312,N_18368,N_19325);
nand U20313 (N_20313,N_18221,N_19229);
xnor U20314 (N_20314,N_18010,N_18456);
nor U20315 (N_20315,N_18794,N_18937);
nand U20316 (N_20316,N_18441,N_19271);
nand U20317 (N_20317,N_18433,N_18975);
nor U20318 (N_20318,N_18677,N_19294);
or U20319 (N_20319,N_18093,N_19417);
and U20320 (N_20320,N_19486,N_18140);
and U20321 (N_20321,N_18054,N_19316);
nand U20322 (N_20322,N_19498,N_18885);
nand U20323 (N_20323,N_19407,N_18881);
nor U20324 (N_20324,N_19246,N_18451);
nor U20325 (N_20325,N_19261,N_19482);
and U20326 (N_20326,N_19071,N_19150);
nand U20327 (N_20327,N_18974,N_18797);
or U20328 (N_20328,N_18447,N_18872);
nand U20329 (N_20329,N_19058,N_19373);
or U20330 (N_20330,N_19007,N_18502);
and U20331 (N_20331,N_19014,N_19412);
or U20332 (N_20332,N_19190,N_18713);
xor U20333 (N_20333,N_18242,N_19275);
xor U20334 (N_20334,N_19452,N_19116);
xnor U20335 (N_20335,N_18253,N_18973);
xnor U20336 (N_20336,N_18878,N_19250);
nor U20337 (N_20337,N_19248,N_18263);
nor U20338 (N_20338,N_18015,N_19074);
nor U20339 (N_20339,N_18987,N_18584);
or U20340 (N_20340,N_19426,N_18350);
nand U20341 (N_20341,N_18868,N_18454);
nand U20342 (N_20342,N_19178,N_18663);
xor U20343 (N_20343,N_18664,N_18279);
nand U20344 (N_20344,N_18161,N_18057);
or U20345 (N_20345,N_18234,N_19420);
nor U20346 (N_20346,N_18956,N_18642);
nand U20347 (N_20347,N_18062,N_18642);
or U20348 (N_20348,N_19493,N_19245);
nor U20349 (N_20349,N_18099,N_19300);
or U20350 (N_20350,N_18664,N_18764);
nand U20351 (N_20351,N_18283,N_18988);
nor U20352 (N_20352,N_18131,N_18049);
nor U20353 (N_20353,N_19448,N_18245);
nor U20354 (N_20354,N_19304,N_18716);
and U20355 (N_20355,N_18986,N_19006);
nor U20356 (N_20356,N_18286,N_18243);
nand U20357 (N_20357,N_18969,N_18074);
nor U20358 (N_20358,N_18045,N_19135);
xnor U20359 (N_20359,N_19010,N_18643);
or U20360 (N_20360,N_19247,N_18526);
and U20361 (N_20361,N_18168,N_18008);
xor U20362 (N_20362,N_19469,N_19204);
xor U20363 (N_20363,N_18042,N_19118);
nand U20364 (N_20364,N_19188,N_18494);
and U20365 (N_20365,N_19250,N_19397);
xnor U20366 (N_20366,N_18869,N_19158);
nand U20367 (N_20367,N_18344,N_19444);
or U20368 (N_20368,N_18165,N_18510);
nor U20369 (N_20369,N_18802,N_18552);
xnor U20370 (N_20370,N_19440,N_18552);
and U20371 (N_20371,N_18402,N_18426);
xor U20372 (N_20372,N_18690,N_19086);
nor U20373 (N_20373,N_18026,N_18501);
nand U20374 (N_20374,N_18492,N_18634);
or U20375 (N_20375,N_19101,N_18325);
and U20376 (N_20376,N_18157,N_19133);
or U20377 (N_20377,N_18609,N_18014);
or U20378 (N_20378,N_18483,N_18585);
or U20379 (N_20379,N_19174,N_19398);
nand U20380 (N_20380,N_18382,N_18353);
xnor U20381 (N_20381,N_18144,N_18106);
nor U20382 (N_20382,N_18563,N_18215);
and U20383 (N_20383,N_18498,N_18211);
nor U20384 (N_20384,N_18417,N_19408);
nor U20385 (N_20385,N_19440,N_18942);
or U20386 (N_20386,N_18587,N_18950);
nor U20387 (N_20387,N_18587,N_18571);
xnor U20388 (N_20388,N_19123,N_19019);
nor U20389 (N_20389,N_19290,N_18103);
nand U20390 (N_20390,N_18143,N_19289);
xnor U20391 (N_20391,N_19439,N_18117);
xnor U20392 (N_20392,N_19299,N_18660);
and U20393 (N_20393,N_18305,N_18393);
and U20394 (N_20394,N_19212,N_19264);
and U20395 (N_20395,N_18017,N_18083);
or U20396 (N_20396,N_19492,N_19159);
or U20397 (N_20397,N_18798,N_18862);
xor U20398 (N_20398,N_18332,N_18635);
nor U20399 (N_20399,N_18035,N_19242);
and U20400 (N_20400,N_19355,N_19415);
nor U20401 (N_20401,N_18580,N_19068);
and U20402 (N_20402,N_18815,N_19376);
and U20403 (N_20403,N_18521,N_18686);
nor U20404 (N_20404,N_19374,N_19059);
nand U20405 (N_20405,N_18755,N_18303);
nor U20406 (N_20406,N_18635,N_19076);
and U20407 (N_20407,N_18628,N_18121);
xnor U20408 (N_20408,N_18854,N_18956);
nor U20409 (N_20409,N_18713,N_18384);
nand U20410 (N_20410,N_18537,N_18409);
or U20411 (N_20411,N_18575,N_18693);
and U20412 (N_20412,N_19289,N_18198);
and U20413 (N_20413,N_19154,N_19106);
and U20414 (N_20414,N_18558,N_18581);
xnor U20415 (N_20415,N_18152,N_19290);
nand U20416 (N_20416,N_18015,N_18675);
nor U20417 (N_20417,N_18780,N_18575);
nor U20418 (N_20418,N_18505,N_19138);
xnor U20419 (N_20419,N_18727,N_19264);
nand U20420 (N_20420,N_18138,N_18214);
xor U20421 (N_20421,N_19244,N_18793);
or U20422 (N_20422,N_18017,N_18998);
nor U20423 (N_20423,N_18059,N_18522);
and U20424 (N_20424,N_18767,N_18859);
and U20425 (N_20425,N_18942,N_19126);
or U20426 (N_20426,N_18746,N_18982);
and U20427 (N_20427,N_19448,N_18934);
xnor U20428 (N_20428,N_18152,N_18085);
nand U20429 (N_20429,N_18269,N_18171);
nor U20430 (N_20430,N_18450,N_18949);
xnor U20431 (N_20431,N_18390,N_18414);
xor U20432 (N_20432,N_19272,N_18224);
xor U20433 (N_20433,N_18121,N_18128);
nand U20434 (N_20434,N_19286,N_18601);
nand U20435 (N_20435,N_18121,N_18587);
xor U20436 (N_20436,N_19315,N_18127);
and U20437 (N_20437,N_19117,N_18834);
nor U20438 (N_20438,N_18459,N_18562);
nand U20439 (N_20439,N_18998,N_18984);
and U20440 (N_20440,N_18231,N_18838);
xnor U20441 (N_20441,N_18540,N_19446);
xnor U20442 (N_20442,N_18735,N_19352);
xor U20443 (N_20443,N_18547,N_18261);
and U20444 (N_20444,N_18844,N_18997);
nand U20445 (N_20445,N_18319,N_19308);
and U20446 (N_20446,N_19247,N_18307);
or U20447 (N_20447,N_18816,N_18632);
and U20448 (N_20448,N_19080,N_19411);
nor U20449 (N_20449,N_18698,N_18444);
xnor U20450 (N_20450,N_18333,N_18865);
or U20451 (N_20451,N_18347,N_19446);
and U20452 (N_20452,N_18182,N_18521);
nor U20453 (N_20453,N_18800,N_18129);
nor U20454 (N_20454,N_18050,N_18600);
nor U20455 (N_20455,N_18178,N_19128);
nand U20456 (N_20456,N_18976,N_18432);
xnor U20457 (N_20457,N_19117,N_18653);
and U20458 (N_20458,N_18773,N_18613);
or U20459 (N_20459,N_19089,N_18786);
nor U20460 (N_20460,N_18791,N_18132);
nor U20461 (N_20461,N_19190,N_18069);
or U20462 (N_20462,N_18111,N_19141);
or U20463 (N_20463,N_19024,N_18228);
or U20464 (N_20464,N_18081,N_18441);
and U20465 (N_20465,N_19054,N_18767);
nand U20466 (N_20466,N_18548,N_18665);
nand U20467 (N_20467,N_18174,N_19337);
and U20468 (N_20468,N_19250,N_19261);
nand U20469 (N_20469,N_19380,N_19253);
xnor U20470 (N_20470,N_18342,N_18742);
and U20471 (N_20471,N_18518,N_19118);
xor U20472 (N_20472,N_18523,N_18743);
nor U20473 (N_20473,N_19456,N_18570);
or U20474 (N_20474,N_19433,N_19057);
or U20475 (N_20475,N_18073,N_18815);
nand U20476 (N_20476,N_19075,N_19021);
xnor U20477 (N_20477,N_18729,N_19455);
or U20478 (N_20478,N_18920,N_19296);
xnor U20479 (N_20479,N_18017,N_19471);
nand U20480 (N_20480,N_18513,N_18225);
nand U20481 (N_20481,N_18046,N_18091);
nand U20482 (N_20482,N_18518,N_18992);
nor U20483 (N_20483,N_19082,N_18784);
nor U20484 (N_20484,N_18342,N_19027);
nand U20485 (N_20485,N_18669,N_18865);
and U20486 (N_20486,N_19218,N_18223);
nor U20487 (N_20487,N_19190,N_19449);
or U20488 (N_20488,N_18051,N_19009);
and U20489 (N_20489,N_19250,N_18145);
and U20490 (N_20490,N_18384,N_18274);
or U20491 (N_20491,N_19321,N_18859);
nor U20492 (N_20492,N_18775,N_18161);
xnor U20493 (N_20493,N_18384,N_18176);
nor U20494 (N_20494,N_18807,N_19099);
nand U20495 (N_20495,N_18042,N_19242);
xnor U20496 (N_20496,N_18524,N_18201);
nand U20497 (N_20497,N_18615,N_18597);
nand U20498 (N_20498,N_19327,N_19161);
and U20499 (N_20499,N_18617,N_18120);
xor U20500 (N_20500,N_18601,N_18666);
xnor U20501 (N_20501,N_19083,N_18793);
and U20502 (N_20502,N_19256,N_18179);
and U20503 (N_20503,N_18840,N_18024);
and U20504 (N_20504,N_18347,N_18875);
nand U20505 (N_20505,N_19378,N_18391);
or U20506 (N_20506,N_19027,N_19464);
and U20507 (N_20507,N_19128,N_19125);
nor U20508 (N_20508,N_18893,N_18399);
or U20509 (N_20509,N_18349,N_19280);
or U20510 (N_20510,N_19186,N_18621);
nor U20511 (N_20511,N_18850,N_19052);
nand U20512 (N_20512,N_19498,N_18341);
and U20513 (N_20513,N_18081,N_18431);
and U20514 (N_20514,N_19477,N_19054);
or U20515 (N_20515,N_19398,N_18917);
nand U20516 (N_20516,N_19365,N_19393);
nand U20517 (N_20517,N_18380,N_19077);
xnor U20518 (N_20518,N_19432,N_19402);
or U20519 (N_20519,N_18967,N_18597);
nand U20520 (N_20520,N_18923,N_18514);
xnor U20521 (N_20521,N_18173,N_18388);
and U20522 (N_20522,N_18048,N_18202);
nor U20523 (N_20523,N_18393,N_18364);
nor U20524 (N_20524,N_19131,N_18082);
or U20525 (N_20525,N_18263,N_18141);
nor U20526 (N_20526,N_18382,N_18012);
and U20527 (N_20527,N_19486,N_18591);
xnor U20528 (N_20528,N_19068,N_18255);
and U20529 (N_20529,N_18724,N_18037);
and U20530 (N_20530,N_18208,N_19423);
or U20531 (N_20531,N_19461,N_19372);
nor U20532 (N_20532,N_19158,N_19486);
nand U20533 (N_20533,N_19248,N_18703);
and U20534 (N_20534,N_19367,N_19446);
or U20535 (N_20535,N_18108,N_19318);
nand U20536 (N_20536,N_19262,N_19043);
xnor U20537 (N_20537,N_19104,N_18635);
or U20538 (N_20538,N_19271,N_18618);
xor U20539 (N_20539,N_18804,N_19352);
xnor U20540 (N_20540,N_19160,N_19238);
nand U20541 (N_20541,N_19314,N_18426);
or U20542 (N_20542,N_18586,N_18959);
xor U20543 (N_20543,N_18264,N_19324);
or U20544 (N_20544,N_19474,N_18516);
nor U20545 (N_20545,N_19009,N_18234);
nand U20546 (N_20546,N_18400,N_18409);
xor U20547 (N_20547,N_19253,N_18112);
nand U20548 (N_20548,N_18050,N_18626);
or U20549 (N_20549,N_18570,N_18200);
nand U20550 (N_20550,N_18191,N_18949);
nor U20551 (N_20551,N_18039,N_18237);
nor U20552 (N_20552,N_19123,N_19060);
and U20553 (N_20553,N_18809,N_18778);
nand U20554 (N_20554,N_18914,N_18243);
and U20555 (N_20555,N_18424,N_18418);
and U20556 (N_20556,N_18073,N_18759);
and U20557 (N_20557,N_19251,N_18005);
and U20558 (N_20558,N_18677,N_19386);
xor U20559 (N_20559,N_18911,N_19474);
or U20560 (N_20560,N_18881,N_18788);
nor U20561 (N_20561,N_18547,N_19421);
nor U20562 (N_20562,N_19226,N_18191);
xor U20563 (N_20563,N_19359,N_18896);
nand U20564 (N_20564,N_18899,N_19335);
xnor U20565 (N_20565,N_18190,N_18882);
nand U20566 (N_20566,N_19342,N_18363);
xor U20567 (N_20567,N_18018,N_19406);
or U20568 (N_20568,N_18280,N_18334);
xor U20569 (N_20569,N_19234,N_18000);
and U20570 (N_20570,N_19401,N_18241);
nor U20571 (N_20571,N_19046,N_19105);
nor U20572 (N_20572,N_18683,N_19209);
nor U20573 (N_20573,N_18588,N_19443);
nor U20574 (N_20574,N_18295,N_18975);
and U20575 (N_20575,N_18186,N_18010);
and U20576 (N_20576,N_18526,N_19471);
and U20577 (N_20577,N_18020,N_19119);
and U20578 (N_20578,N_18314,N_18428);
or U20579 (N_20579,N_19071,N_18311);
and U20580 (N_20580,N_19169,N_18397);
and U20581 (N_20581,N_19010,N_18259);
or U20582 (N_20582,N_18405,N_19073);
or U20583 (N_20583,N_18694,N_18708);
xnor U20584 (N_20584,N_19257,N_18518);
nand U20585 (N_20585,N_19161,N_18017);
nor U20586 (N_20586,N_18070,N_18792);
nand U20587 (N_20587,N_19322,N_18444);
nor U20588 (N_20588,N_18642,N_18689);
and U20589 (N_20589,N_19059,N_19415);
nand U20590 (N_20590,N_18818,N_19042);
xor U20591 (N_20591,N_18125,N_19032);
nand U20592 (N_20592,N_18963,N_19490);
nand U20593 (N_20593,N_18023,N_18267);
xnor U20594 (N_20594,N_18985,N_18222);
xnor U20595 (N_20595,N_18163,N_18862);
or U20596 (N_20596,N_18980,N_19358);
nor U20597 (N_20597,N_18091,N_19149);
or U20598 (N_20598,N_19184,N_18158);
nand U20599 (N_20599,N_18767,N_18092);
xnor U20600 (N_20600,N_18717,N_18707);
nor U20601 (N_20601,N_18295,N_19028);
and U20602 (N_20602,N_18396,N_19430);
nor U20603 (N_20603,N_18985,N_19025);
xor U20604 (N_20604,N_19059,N_18342);
nand U20605 (N_20605,N_18619,N_18437);
nor U20606 (N_20606,N_18129,N_18288);
or U20607 (N_20607,N_19304,N_19114);
and U20608 (N_20608,N_19357,N_18056);
and U20609 (N_20609,N_18298,N_18814);
nand U20610 (N_20610,N_19227,N_18279);
xor U20611 (N_20611,N_19081,N_18555);
and U20612 (N_20612,N_19334,N_19039);
or U20613 (N_20613,N_19496,N_18029);
xor U20614 (N_20614,N_18043,N_18575);
or U20615 (N_20615,N_18679,N_19364);
and U20616 (N_20616,N_18564,N_18894);
nand U20617 (N_20617,N_18395,N_18363);
or U20618 (N_20618,N_18891,N_18144);
nor U20619 (N_20619,N_18026,N_18300);
xor U20620 (N_20620,N_19430,N_19028);
nand U20621 (N_20621,N_18317,N_18930);
or U20622 (N_20622,N_18064,N_18541);
and U20623 (N_20623,N_19315,N_19488);
xor U20624 (N_20624,N_18125,N_19480);
nand U20625 (N_20625,N_18761,N_19326);
nor U20626 (N_20626,N_19084,N_18290);
nand U20627 (N_20627,N_19183,N_19377);
xnor U20628 (N_20628,N_18011,N_18424);
or U20629 (N_20629,N_18301,N_18056);
xor U20630 (N_20630,N_19309,N_19125);
and U20631 (N_20631,N_18949,N_18024);
or U20632 (N_20632,N_19338,N_18834);
nand U20633 (N_20633,N_18642,N_18607);
or U20634 (N_20634,N_18667,N_18111);
and U20635 (N_20635,N_19323,N_19496);
xnor U20636 (N_20636,N_18733,N_19273);
or U20637 (N_20637,N_18922,N_19305);
and U20638 (N_20638,N_18916,N_18145);
xnor U20639 (N_20639,N_18364,N_18138);
or U20640 (N_20640,N_18702,N_19307);
nand U20641 (N_20641,N_18311,N_19407);
nand U20642 (N_20642,N_18681,N_18962);
nand U20643 (N_20643,N_19027,N_18019);
and U20644 (N_20644,N_18507,N_18583);
or U20645 (N_20645,N_18223,N_19121);
xor U20646 (N_20646,N_18193,N_18312);
or U20647 (N_20647,N_18038,N_18339);
xor U20648 (N_20648,N_18156,N_18824);
nand U20649 (N_20649,N_19333,N_18834);
nand U20650 (N_20650,N_19457,N_18458);
xnor U20651 (N_20651,N_18766,N_18460);
xnor U20652 (N_20652,N_18914,N_18777);
nor U20653 (N_20653,N_19001,N_19078);
and U20654 (N_20654,N_18258,N_19188);
xnor U20655 (N_20655,N_18670,N_19000);
or U20656 (N_20656,N_19105,N_18968);
and U20657 (N_20657,N_18557,N_18163);
xnor U20658 (N_20658,N_19304,N_18498);
and U20659 (N_20659,N_18981,N_18172);
or U20660 (N_20660,N_18302,N_18003);
nand U20661 (N_20661,N_18421,N_18034);
and U20662 (N_20662,N_18936,N_18693);
nand U20663 (N_20663,N_18429,N_18864);
and U20664 (N_20664,N_18702,N_18799);
nand U20665 (N_20665,N_18273,N_18613);
nand U20666 (N_20666,N_18285,N_19028);
nor U20667 (N_20667,N_18985,N_18597);
and U20668 (N_20668,N_18171,N_19459);
nand U20669 (N_20669,N_18413,N_18823);
xnor U20670 (N_20670,N_18910,N_18608);
or U20671 (N_20671,N_19210,N_19499);
and U20672 (N_20672,N_18497,N_18255);
and U20673 (N_20673,N_18324,N_19187);
nand U20674 (N_20674,N_19264,N_18174);
nor U20675 (N_20675,N_18911,N_18462);
nand U20676 (N_20676,N_18123,N_19154);
nor U20677 (N_20677,N_18412,N_18570);
and U20678 (N_20678,N_19094,N_18582);
or U20679 (N_20679,N_18830,N_18736);
xor U20680 (N_20680,N_18544,N_18562);
nor U20681 (N_20681,N_18668,N_18903);
nand U20682 (N_20682,N_18733,N_18514);
xnor U20683 (N_20683,N_18895,N_18228);
and U20684 (N_20684,N_18958,N_18880);
nand U20685 (N_20685,N_18092,N_18465);
nand U20686 (N_20686,N_19012,N_19218);
and U20687 (N_20687,N_18914,N_18753);
nor U20688 (N_20688,N_18809,N_19106);
xnor U20689 (N_20689,N_18812,N_18085);
and U20690 (N_20690,N_18029,N_19403);
and U20691 (N_20691,N_18439,N_19468);
nand U20692 (N_20692,N_19477,N_18384);
or U20693 (N_20693,N_18663,N_18341);
and U20694 (N_20694,N_18750,N_18086);
xnor U20695 (N_20695,N_18163,N_18432);
xnor U20696 (N_20696,N_19413,N_19067);
nor U20697 (N_20697,N_19121,N_18421);
nor U20698 (N_20698,N_19316,N_18071);
nand U20699 (N_20699,N_18523,N_18093);
or U20700 (N_20700,N_18776,N_19128);
xor U20701 (N_20701,N_18010,N_18183);
and U20702 (N_20702,N_19390,N_18876);
xor U20703 (N_20703,N_18466,N_19471);
nor U20704 (N_20704,N_18119,N_19278);
nor U20705 (N_20705,N_19023,N_19059);
and U20706 (N_20706,N_19251,N_19433);
or U20707 (N_20707,N_18413,N_18476);
nor U20708 (N_20708,N_18906,N_19448);
and U20709 (N_20709,N_18089,N_18580);
nand U20710 (N_20710,N_19322,N_18165);
xor U20711 (N_20711,N_19298,N_19225);
and U20712 (N_20712,N_18392,N_18047);
nand U20713 (N_20713,N_18358,N_18331);
and U20714 (N_20714,N_18238,N_19452);
xnor U20715 (N_20715,N_19294,N_18344);
nor U20716 (N_20716,N_18433,N_18247);
nor U20717 (N_20717,N_18906,N_19445);
or U20718 (N_20718,N_19070,N_19470);
nor U20719 (N_20719,N_18721,N_19273);
nor U20720 (N_20720,N_18489,N_18613);
xnor U20721 (N_20721,N_18681,N_19311);
or U20722 (N_20722,N_18236,N_19252);
or U20723 (N_20723,N_18792,N_18799);
or U20724 (N_20724,N_19013,N_18261);
and U20725 (N_20725,N_18856,N_18388);
and U20726 (N_20726,N_19150,N_18279);
and U20727 (N_20727,N_19335,N_19125);
xnor U20728 (N_20728,N_18769,N_19190);
nand U20729 (N_20729,N_18246,N_18632);
and U20730 (N_20730,N_18065,N_18019);
xnor U20731 (N_20731,N_18798,N_18250);
and U20732 (N_20732,N_18911,N_18301);
nand U20733 (N_20733,N_19195,N_18839);
xor U20734 (N_20734,N_18369,N_19393);
or U20735 (N_20735,N_18970,N_19268);
or U20736 (N_20736,N_18442,N_18909);
nor U20737 (N_20737,N_18567,N_19161);
xnor U20738 (N_20738,N_19468,N_19494);
nand U20739 (N_20739,N_18481,N_18225);
nand U20740 (N_20740,N_19005,N_18628);
nor U20741 (N_20741,N_19190,N_18930);
xor U20742 (N_20742,N_19368,N_18674);
and U20743 (N_20743,N_19278,N_18837);
nand U20744 (N_20744,N_18484,N_18233);
nand U20745 (N_20745,N_18634,N_19191);
nor U20746 (N_20746,N_19403,N_18602);
nand U20747 (N_20747,N_18971,N_18937);
nor U20748 (N_20748,N_18774,N_19078);
and U20749 (N_20749,N_18372,N_18239);
nor U20750 (N_20750,N_19445,N_18669);
or U20751 (N_20751,N_18629,N_19334);
or U20752 (N_20752,N_19107,N_19309);
nand U20753 (N_20753,N_19035,N_19420);
xor U20754 (N_20754,N_19309,N_18348);
xnor U20755 (N_20755,N_19262,N_19002);
xor U20756 (N_20756,N_18913,N_18030);
nor U20757 (N_20757,N_18775,N_19043);
nor U20758 (N_20758,N_19175,N_19478);
xnor U20759 (N_20759,N_19024,N_18629);
nor U20760 (N_20760,N_18285,N_18062);
xnor U20761 (N_20761,N_18686,N_18754);
nand U20762 (N_20762,N_19493,N_18637);
and U20763 (N_20763,N_19476,N_18580);
and U20764 (N_20764,N_19380,N_19355);
xor U20765 (N_20765,N_18853,N_19307);
nand U20766 (N_20766,N_18925,N_18478);
nor U20767 (N_20767,N_19415,N_19417);
nor U20768 (N_20768,N_19129,N_18668);
xnor U20769 (N_20769,N_18405,N_18041);
xnor U20770 (N_20770,N_18605,N_18949);
nor U20771 (N_20771,N_19372,N_18907);
or U20772 (N_20772,N_18207,N_18914);
nor U20773 (N_20773,N_18339,N_18614);
xnor U20774 (N_20774,N_18560,N_19207);
nor U20775 (N_20775,N_18965,N_18247);
and U20776 (N_20776,N_18379,N_18192);
or U20777 (N_20777,N_18872,N_18689);
nor U20778 (N_20778,N_18516,N_18617);
or U20779 (N_20779,N_18053,N_18231);
nand U20780 (N_20780,N_19457,N_19005);
and U20781 (N_20781,N_18350,N_18559);
xnor U20782 (N_20782,N_18745,N_19370);
or U20783 (N_20783,N_19381,N_18643);
and U20784 (N_20784,N_18748,N_18551);
xnor U20785 (N_20785,N_18127,N_18071);
or U20786 (N_20786,N_18817,N_19422);
xnor U20787 (N_20787,N_18312,N_18373);
and U20788 (N_20788,N_18327,N_19175);
and U20789 (N_20789,N_19152,N_19257);
nor U20790 (N_20790,N_19091,N_19346);
xor U20791 (N_20791,N_19335,N_18544);
and U20792 (N_20792,N_18393,N_18778);
xnor U20793 (N_20793,N_18571,N_18202);
xor U20794 (N_20794,N_18270,N_18361);
or U20795 (N_20795,N_18711,N_18848);
or U20796 (N_20796,N_18771,N_19162);
and U20797 (N_20797,N_18216,N_19307);
or U20798 (N_20798,N_19277,N_18092);
nor U20799 (N_20799,N_18411,N_18454);
or U20800 (N_20800,N_18935,N_19010);
nand U20801 (N_20801,N_18044,N_18316);
nor U20802 (N_20802,N_18487,N_19047);
or U20803 (N_20803,N_18660,N_18241);
or U20804 (N_20804,N_18763,N_18299);
or U20805 (N_20805,N_18606,N_19015);
nand U20806 (N_20806,N_18025,N_19490);
and U20807 (N_20807,N_19052,N_18125);
or U20808 (N_20808,N_18727,N_18857);
nor U20809 (N_20809,N_18934,N_18530);
or U20810 (N_20810,N_18263,N_18625);
nor U20811 (N_20811,N_18852,N_18398);
and U20812 (N_20812,N_19013,N_19303);
and U20813 (N_20813,N_18384,N_18115);
and U20814 (N_20814,N_18673,N_19311);
xnor U20815 (N_20815,N_18952,N_19198);
or U20816 (N_20816,N_18267,N_18278);
xnor U20817 (N_20817,N_19346,N_18162);
xnor U20818 (N_20818,N_19321,N_19217);
xnor U20819 (N_20819,N_18205,N_19466);
or U20820 (N_20820,N_18223,N_18609);
nor U20821 (N_20821,N_19343,N_18008);
nand U20822 (N_20822,N_18185,N_19150);
xor U20823 (N_20823,N_18815,N_18987);
nand U20824 (N_20824,N_18648,N_18655);
and U20825 (N_20825,N_19036,N_19486);
and U20826 (N_20826,N_18841,N_18753);
xor U20827 (N_20827,N_18452,N_18999);
nor U20828 (N_20828,N_18548,N_19101);
nor U20829 (N_20829,N_18358,N_19219);
and U20830 (N_20830,N_19226,N_19335);
xor U20831 (N_20831,N_18177,N_18642);
and U20832 (N_20832,N_18167,N_18762);
and U20833 (N_20833,N_19486,N_18024);
or U20834 (N_20834,N_18431,N_18289);
nor U20835 (N_20835,N_18302,N_19484);
nand U20836 (N_20836,N_19217,N_18755);
nand U20837 (N_20837,N_19179,N_18881);
xor U20838 (N_20838,N_18686,N_19346);
xnor U20839 (N_20839,N_18217,N_19109);
and U20840 (N_20840,N_18203,N_18350);
or U20841 (N_20841,N_19259,N_18103);
nand U20842 (N_20842,N_19272,N_19042);
nor U20843 (N_20843,N_18828,N_18383);
xnor U20844 (N_20844,N_18271,N_18940);
and U20845 (N_20845,N_18838,N_19477);
nand U20846 (N_20846,N_18897,N_18789);
and U20847 (N_20847,N_18647,N_19212);
or U20848 (N_20848,N_19468,N_18249);
nor U20849 (N_20849,N_18480,N_19492);
nor U20850 (N_20850,N_19359,N_18978);
nand U20851 (N_20851,N_19240,N_18156);
or U20852 (N_20852,N_18652,N_19097);
or U20853 (N_20853,N_18380,N_18778);
nor U20854 (N_20854,N_19396,N_19442);
xor U20855 (N_20855,N_18421,N_18161);
or U20856 (N_20856,N_18491,N_18459);
nand U20857 (N_20857,N_19203,N_18251);
and U20858 (N_20858,N_19210,N_19226);
xor U20859 (N_20859,N_18856,N_18339);
nor U20860 (N_20860,N_19240,N_18403);
nand U20861 (N_20861,N_18931,N_18082);
or U20862 (N_20862,N_19408,N_19320);
or U20863 (N_20863,N_19248,N_19071);
nor U20864 (N_20864,N_18394,N_18751);
nand U20865 (N_20865,N_18978,N_19156);
xor U20866 (N_20866,N_19203,N_18667);
and U20867 (N_20867,N_18051,N_18818);
and U20868 (N_20868,N_18824,N_18095);
and U20869 (N_20869,N_19423,N_18252);
nand U20870 (N_20870,N_18288,N_19400);
and U20871 (N_20871,N_18269,N_19079);
or U20872 (N_20872,N_18736,N_19292);
nand U20873 (N_20873,N_18774,N_18495);
nor U20874 (N_20874,N_18015,N_19400);
xnor U20875 (N_20875,N_18394,N_18063);
nand U20876 (N_20876,N_18917,N_18001);
xor U20877 (N_20877,N_18139,N_19344);
nor U20878 (N_20878,N_18302,N_18688);
nand U20879 (N_20879,N_18233,N_18641);
xor U20880 (N_20880,N_19275,N_19073);
or U20881 (N_20881,N_18284,N_18836);
and U20882 (N_20882,N_19257,N_18098);
or U20883 (N_20883,N_18789,N_18548);
or U20884 (N_20884,N_18226,N_18987);
nor U20885 (N_20885,N_18482,N_18879);
or U20886 (N_20886,N_18869,N_18968);
nor U20887 (N_20887,N_18111,N_18084);
or U20888 (N_20888,N_19259,N_18774);
nand U20889 (N_20889,N_18249,N_19157);
and U20890 (N_20890,N_18828,N_18482);
nand U20891 (N_20891,N_18387,N_19422);
and U20892 (N_20892,N_18678,N_18917);
xnor U20893 (N_20893,N_19489,N_18445);
and U20894 (N_20894,N_18667,N_19086);
nor U20895 (N_20895,N_19074,N_18934);
nand U20896 (N_20896,N_19466,N_18517);
or U20897 (N_20897,N_18307,N_18130);
and U20898 (N_20898,N_18302,N_18384);
nand U20899 (N_20899,N_18392,N_18496);
nand U20900 (N_20900,N_18095,N_18280);
nand U20901 (N_20901,N_18408,N_19083);
nand U20902 (N_20902,N_18928,N_19331);
or U20903 (N_20903,N_18189,N_18782);
xnor U20904 (N_20904,N_18644,N_18938);
or U20905 (N_20905,N_18854,N_18363);
or U20906 (N_20906,N_18949,N_18458);
nor U20907 (N_20907,N_19279,N_18799);
and U20908 (N_20908,N_18380,N_19208);
and U20909 (N_20909,N_19357,N_18108);
and U20910 (N_20910,N_18640,N_18691);
nor U20911 (N_20911,N_19160,N_19020);
xor U20912 (N_20912,N_18333,N_18553);
nand U20913 (N_20913,N_18048,N_18088);
nor U20914 (N_20914,N_19254,N_18275);
nand U20915 (N_20915,N_18568,N_19014);
xnor U20916 (N_20916,N_18881,N_18612);
nor U20917 (N_20917,N_18990,N_19324);
or U20918 (N_20918,N_18941,N_18228);
and U20919 (N_20919,N_19162,N_18128);
and U20920 (N_20920,N_19424,N_18264);
nand U20921 (N_20921,N_18204,N_19470);
nand U20922 (N_20922,N_18718,N_19339);
or U20923 (N_20923,N_19157,N_18996);
nand U20924 (N_20924,N_18085,N_18238);
or U20925 (N_20925,N_19257,N_18038);
and U20926 (N_20926,N_19142,N_18304);
nor U20927 (N_20927,N_19256,N_18134);
and U20928 (N_20928,N_18686,N_19499);
and U20929 (N_20929,N_18809,N_18197);
and U20930 (N_20930,N_18211,N_18680);
xor U20931 (N_20931,N_18843,N_19217);
and U20932 (N_20932,N_18205,N_18746);
and U20933 (N_20933,N_18546,N_18975);
nor U20934 (N_20934,N_18568,N_18136);
xnor U20935 (N_20935,N_19419,N_18605);
and U20936 (N_20936,N_18713,N_18780);
nand U20937 (N_20937,N_18533,N_18518);
and U20938 (N_20938,N_19367,N_19178);
xnor U20939 (N_20939,N_18658,N_18434);
nor U20940 (N_20940,N_19293,N_18048);
and U20941 (N_20941,N_18933,N_18638);
nor U20942 (N_20942,N_18633,N_18873);
xor U20943 (N_20943,N_19277,N_19312);
or U20944 (N_20944,N_19367,N_18319);
xor U20945 (N_20945,N_18126,N_18437);
nand U20946 (N_20946,N_18357,N_18697);
and U20947 (N_20947,N_18484,N_18088);
nor U20948 (N_20948,N_18253,N_18660);
nand U20949 (N_20949,N_18855,N_18267);
or U20950 (N_20950,N_18853,N_19218);
or U20951 (N_20951,N_18365,N_18278);
nand U20952 (N_20952,N_18565,N_18087);
nand U20953 (N_20953,N_18459,N_18552);
or U20954 (N_20954,N_18711,N_19122);
and U20955 (N_20955,N_19146,N_18364);
or U20956 (N_20956,N_19210,N_18591);
or U20957 (N_20957,N_18071,N_18577);
or U20958 (N_20958,N_18897,N_18032);
xor U20959 (N_20959,N_19462,N_18220);
nor U20960 (N_20960,N_18793,N_19331);
xnor U20961 (N_20961,N_18175,N_18793);
nand U20962 (N_20962,N_18565,N_19452);
nor U20963 (N_20963,N_18504,N_18017);
xor U20964 (N_20964,N_19168,N_18815);
nand U20965 (N_20965,N_19013,N_18236);
xor U20966 (N_20966,N_18915,N_19086);
nand U20967 (N_20967,N_19114,N_18345);
xor U20968 (N_20968,N_18877,N_18026);
nand U20969 (N_20969,N_18116,N_18497);
xnor U20970 (N_20970,N_18601,N_18676);
nor U20971 (N_20971,N_19414,N_18736);
nand U20972 (N_20972,N_18364,N_18299);
and U20973 (N_20973,N_18161,N_18872);
xnor U20974 (N_20974,N_19112,N_19310);
nand U20975 (N_20975,N_18826,N_18164);
nand U20976 (N_20976,N_19197,N_18360);
or U20977 (N_20977,N_19296,N_19446);
xnor U20978 (N_20978,N_19178,N_18709);
xnor U20979 (N_20979,N_19282,N_18468);
or U20980 (N_20980,N_18581,N_18179);
nor U20981 (N_20981,N_18339,N_18502);
nand U20982 (N_20982,N_18996,N_18722);
or U20983 (N_20983,N_18753,N_18924);
nor U20984 (N_20984,N_18697,N_18095);
nand U20985 (N_20985,N_18347,N_18618);
or U20986 (N_20986,N_19154,N_18609);
nor U20987 (N_20987,N_19066,N_18488);
or U20988 (N_20988,N_18413,N_18560);
nor U20989 (N_20989,N_18768,N_18878);
or U20990 (N_20990,N_18038,N_18015);
nor U20991 (N_20991,N_19074,N_18931);
nand U20992 (N_20992,N_18026,N_18234);
or U20993 (N_20993,N_18702,N_18902);
xnor U20994 (N_20994,N_19485,N_19424);
or U20995 (N_20995,N_19440,N_18457);
nor U20996 (N_20996,N_18258,N_18610);
xor U20997 (N_20997,N_19281,N_18390);
and U20998 (N_20998,N_18296,N_18314);
nor U20999 (N_20999,N_19115,N_18646);
nand U21000 (N_21000,N_20000,N_20143);
nor U21001 (N_21001,N_20583,N_19796);
nor U21002 (N_21002,N_20633,N_19797);
and U21003 (N_21003,N_20504,N_20398);
nor U21004 (N_21004,N_20196,N_20031);
or U21005 (N_21005,N_20912,N_19750);
nor U21006 (N_21006,N_20709,N_19781);
nand U21007 (N_21007,N_19887,N_20509);
or U21008 (N_21008,N_20058,N_20466);
or U21009 (N_21009,N_20775,N_20636);
or U21010 (N_21010,N_20754,N_19705);
xnor U21011 (N_21011,N_20669,N_20538);
or U21012 (N_21012,N_20543,N_19970);
nor U21013 (N_21013,N_19587,N_20678);
and U21014 (N_21014,N_20873,N_19996);
nand U21015 (N_21015,N_20406,N_19643);
xor U21016 (N_21016,N_19920,N_19949);
and U21017 (N_21017,N_20209,N_20672);
or U21018 (N_21018,N_20213,N_20199);
nand U21019 (N_21019,N_19672,N_20207);
xor U21020 (N_21020,N_19671,N_20751);
nor U21021 (N_21021,N_20387,N_20973);
or U21022 (N_21022,N_20277,N_20424);
xnor U21023 (N_21023,N_19676,N_20476);
xnor U21024 (N_21024,N_19971,N_20298);
nand U21025 (N_21025,N_19967,N_20408);
or U21026 (N_21026,N_20148,N_20690);
xor U21027 (N_21027,N_20378,N_20667);
nor U21028 (N_21028,N_20625,N_19853);
nor U21029 (N_21029,N_20311,N_20262);
nand U21030 (N_21030,N_20698,N_19859);
nor U21031 (N_21031,N_19696,N_19823);
or U21032 (N_21032,N_20452,N_20574);
xor U21033 (N_21033,N_20887,N_20901);
and U21034 (N_21034,N_19885,N_20844);
nand U21035 (N_21035,N_19727,N_20117);
nand U21036 (N_21036,N_20150,N_20315);
xor U21037 (N_21037,N_19907,N_19800);
or U21038 (N_21038,N_20488,N_20962);
or U21039 (N_21039,N_20727,N_20581);
nor U21040 (N_21040,N_20038,N_20511);
nor U21041 (N_21041,N_19819,N_20449);
nand U21042 (N_21042,N_20788,N_20297);
xor U21043 (N_21043,N_20149,N_20464);
xnor U21044 (N_21044,N_19947,N_20187);
nand U21045 (N_21045,N_20125,N_20024);
nor U21046 (N_21046,N_20659,N_20080);
xor U21047 (N_21047,N_20145,N_20542);
and U21048 (N_21048,N_20307,N_20022);
or U21049 (N_21049,N_19906,N_20318);
or U21050 (N_21050,N_20358,N_19986);
nand U21051 (N_21051,N_19846,N_20256);
nand U21052 (N_21052,N_20180,N_20789);
xor U21053 (N_21053,N_19769,N_19863);
nand U21054 (N_21054,N_20655,N_20591);
nand U21055 (N_21055,N_20760,N_20028);
nor U21056 (N_21056,N_19928,N_19686);
xnor U21057 (N_21057,N_20457,N_20558);
and U21058 (N_21058,N_19932,N_20853);
nand U21059 (N_21059,N_20287,N_20520);
nor U21060 (N_21060,N_20579,N_20162);
xnor U21061 (N_21061,N_20649,N_20205);
nand U21062 (N_21062,N_19849,N_19974);
nor U21063 (N_21063,N_20312,N_20878);
nor U21064 (N_21064,N_20093,N_20228);
nor U21065 (N_21065,N_20769,N_20984);
nor U21066 (N_21066,N_20922,N_19555);
xnor U21067 (N_21067,N_19650,N_20498);
and U21068 (N_21068,N_20666,N_19921);
nand U21069 (N_21069,N_20020,N_20695);
or U21070 (N_21070,N_19709,N_20065);
or U21071 (N_21071,N_19662,N_20147);
or U21072 (N_21072,N_20451,N_19680);
and U21073 (N_21073,N_19687,N_20053);
and U21074 (N_21074,N_19597,N_19802);
nor U21075 (N_21075,N_20516,N_20793);
or U21076 (N_21076,N_19673,N_20577);
nor U21077 (N_21077,N_19898,N_19565);
and U21078 (N_21078,N_20338,N_20578);
nor U21079 (N_21079,N_19882,N_20154);
nand U21080 (N_21080,N_20302,N_20238);
xor U21081 (N_21081,N_20765,N_19765);
xnor U21082 (N_21082,N_20160,N_19504);
nor U21083 (N_21083,N_20725,N_19682);
nand U21084 (N_21084,N_20501,N_20391);
or U21085 (N_21085,N_20414,N_19798);
nand U21086 (N_21086,N_20336,N_19814);
xnor U21087 (N_21087,N_19511,N_19522);
and U21088 (N_21088,N_20415,N_20253);
nor U21089 (N_21089,N_20546,N_20816);
and U21090 (N_21090,N_20141,N_20272);
and U21091 (N_21091,N_19507,N_20433);
or U21092 (N_21092,N_20411,N_20771);
and U21093 (N_21093,N_19752,N_19985);
xor U21094 (N_21094,N_19848,N_19837);
nand U21095 (N_21095,N_19799,N_20942);
xnor U21096 (N_21096,N_20936,N_20927);
xor U21097 (N_21097,N_20182,N_19713);
nand U21098 (N_21098,N_19659,N_20326);
nor U21099 (N_21099,N_20100,N_20774);
nor U21100 (N_21100,N_20335,N_19780);
or U21101 (N_21101,N_19722,N_19710);
or U21102 (N_21102,N_20136,N_19707);
or U21103 (N_21103,N_19564,N_19877);
xnor U21104 (N_21104,N_20337,N_20190);
and U21105 (N_21105,N_19913,N_19989);
or U21106 (N_21106,N_20903,N_20316);
nand U21107 (N_21107,N_19935,N_19642);
nand U21108 (N_21108,N_19810,N_20171);
or U21109 (N_21109,N_20214,N_19903);
xor U21110 (N_21110,N_20797,N_19517);
nor U21111 (N_21111,N_19604,N_20385);
xor U21112 (N_21112,N_19841,N_20593);
nand U21113 (N_21113,N_19585,N_20274);
nand U21114 (N_21114,N_20273,N_20620);
nor U21115 (N_21115,N_20185,N_20996);
nand U21116 (N_21116,N_19870,N_20514);
xor U21117 (N_21117,N_20071,N_20462);
nor U21118 (N_21118,N_20327,N_20132);
and U21119 (N_21119,N_19683,N_19776);
nor U21120 (N_21120,N_20393,N_20268);
nand U21121 (N_21121,N_19795,N_19599);
or U21122 (N_21122,N_19622,N_20468);
nand U21123 (N_21123,N_19994,N_20367);
nand U21124 (N_21124,N_20060,N_20242);
and U21125 (N_21125,N_20191,N_20568);
nand U21126 (N_21126,N_20714,N_19843);
and U21127 (N_21127,N_19987,N_19567);
nand U21128 (N_21128,N_20142,N_20308);
nor U21129 (N_21129,N_20941,N_20747);
nand U21130 (N_21130,N_20544,N_20934);
nand U21131 (N_21131,N_19964,N_20164);
or U21132 (N_21132,N_20953,N_20907);
nor U21133 (N_21133,N_20881,N_19602);
or U21134 (N_21134,N_20281,N_20513);
nand U21135 (N_21135,N_20805,N_19806);
xor U21136 (N_21136,N_20267,N_20499);
nand U21137 (N_21137,N_20134,N_20626);
xnor U21138 (N_21138,N_20561,N_19852);
and U21139 (N_21139,N_19756,N_20194);
nor U21140 (N_21140,N_19824,N_20264);
and U21141 (N_21141,N_20928,N_19976);
and U21142 (N_21142,N_20054,N_20215);
and U21143 (N_21143,N_20710,N_20061);
nor U21144 (N_21144,N_20342,N_19689);
and U21145 (N_21145,N_20245,N_20988);
nand U21146 (N_21146,N_20410,N_20004);
or U21147 (N_21147,N_20906,N_20119);
and U21148 (N_21148,N_20838,N_20564);
and U21149 (N_21149,N_19657,N_20346);
nor U21150 (N_21150,N_20115,N_19603);
xnor U21151 (N_21151,N_20833,N_20369);
nor U21152 (N_21152,N_20465,N_19944);
nor U21153 (N_21153,N_20560,N_20001);
xnor U21154 (N_21154,N_20192,N_19869);
nor U21155 (N_21155,N_20949,N_20374);
xnor U21156 (N_21156,N_20653,N_20402);
and U21157 (N_21157,N_19547,N_20777);
nor U21158 (N_21158,N_20703,N_20699);
xnor U21159 (N_21159,N_20434,N_20550);
nand U21160 (N_21160,N_20014,N_19918);
xor U21161 (N_21161,N_20938,N_20379);
or U21162 (N_21162,N_20068,N_20761);
xor U21163 (N_21163,N_20753,N_20758);
or U21164 (N_21164,N_20189,N_20331);
nor U21165 (N_21165,N_19850,N_20631);
or U21166 (N_21166,N_20682,N_20787);
xor U21167 (N_21167,N_19884,N_19988);
or U21168 (N_21168,N_19541,N_20220);
nand U21169 (N_21169,N_20894,N_20131);
or U21170 (N_21170,N_20656,N_20198);
nand U21171 (N_21171,N_19694,N_20045);
xor U21172 (N_21172,N_20744,N_19627);
and U21173 (N_21173,N_20419,N_20517);
or U21174 (N_21174,N_19891,N_20010);
nor U21175 (N_21175,N_19514,N_20594);
nand U21176 (N_21176,N_20485,N_20535);
xor U21177 (N_21177,N_20964,N_20944);
xnor U21178 (N_21178,N_20982,N_20258);
nand U21179 (N_21179,N_19701,N_20899);
and U21180 (N_21180,N_19613,N_19724);
or U21181 (N_21181,N_19542,N_19847);
or U21182 (N_21182,N_19930,N_20027);
nor U21183 (N_21183,N_20124,N_20723);
and U21184 (N_21184,N_19699,N_20321);
or U21185 (N_21185,N_20224,N_19502);
or U21186 (N_21186,N_20586,N_20704);
nor U21187 (N_21187,N_19592,N_19580);
xor U21188 (N_21188,N_20846,N_20324);
or U21189 (N_21189,N_20354,N_20943);
nand U21190 (N_21190,N_19621,N_20933);
nor U21191 (N_21191,N_20279,N_19741);
nor U21192 (N_21192,N_20435,N_20985);
or U21193 (N_21193,N_20286,N_20417);
nor U21194 (N_21194,N_20389,N_20929);
and U21195 (N_21195,N_20939,N_20856);
xnor U21196 (N_21196,N_20382,N_20319);
and U21197 (N_21197,N_19791,N_19833);
nor U21198 (N_21198,N_20571,N_19739);
nor U21199 (N_21199,N_19808,N_20343);
or U21200 (N_21200,N_20030,N_20862);
nor U21201 (N_21201,N_19904,N_19665);
or U21202 (N_21202,N_20486,N_19677);
or U21203 (N_21203,N_19737,N_19844);
and U21204 (N_21204,N_20737,N_20497);
and U21205 (N_21205,N_20019,N_20102);
or U21206 (N_21206,N_20876,N_19829);
xnor U21207 (N_21207,N_19982,N_20694);
or U21208 (N_21208,N_20200,N_20619);
nor U21209 (N_21209,N_19572,N_20521);
or U21210 (N_21210,N_20176,N_19723);
xor U21211 (N_21211,N_19997,N_20233);
xnor U21212 (N_21212,N_20650,N_20240);
nand U21213 (N_21213,N_20551,N_20158);
nand U21214 (N_21214,N_20810,N_20958);
and U21215 (N_21215,N_20735,N_20114);
and U21216 (N_21216,N_19530,N_19893);
xor U21217 (N_21217,N_19998,N_20992);
nand U21218 (N_21218,N_20105,N_20891);
xnor U21219 (N_21219,N_19864,N_19901);
xnor U21220 (N_21220,N_20193,N_19826);
nor U21221 (N_21221,N_20490,N_20721);
and U21222 (N_21222,N_20040,N_19539);
or U21223 (N_21223,N_19560,N_20701);
or U21224 (N_21224,N_20015,N_19733);
or U21225 (N_21225,N_20884,N_20645);
xnor U21226 (N_21226,N_20799,N_20373);
and U21227 (N_21227,N_20403,N_20585);
nand U21228 (N_21228,N_20768,N_20333);
or U21229 (N_21229,N_20370,N_20155);
nand U21230 (N_21230,N_20877,N_20975);
xor U21231 (N_21231,N_19927,N_19693);
or U21232 (N_21232,N_20763,N_19936);
and U21233 (N_21233,N_20118,N_20536);
or U21234 (N_21234,N_19740,N_20914);
and U21235 (N_21235,N_20622,N_19612);
nand U21236 (N_21236,N_20815,N_20186);
or U21237 (N_21237,N_19559,N_20248);
nand U21238 (N_21238,N_20400,N_19678);
and U21239 (N_21239,N_19544,N_20955);
nand U21240 (N_21240,N_19570,N_20526);
or U21241 (N_21241,N_20492,N_19758);
xnor U21242 (N_21242,N_20051,N_20047);
nor U21243 (N_21243,N_20270,N_20880);
or U21244 (N_21244,N_19748,N_20073);
nor U21245 (N_21245,N_20418,N_20288);
or U21246 (N_21246,N_19792,N_20557);
nor U21247 (N_21247,N_20607,N_20099);
nand U21248 (N_21248,N_20685,N_20658);
xnor U21249 (N_21249,N_19875,N_20084);
or U21250 (N_21250,N_20712,N_20066);
nor U21251 (N_21251,N_20580,N_20037);
xor U21252 (N_21252,N_20641,N_20652);
nand U21253 (N_21253,N_20018,N_20831);
nor U21254 (N_21254,N_20630,N_19924);
nor U21255 (N_21255,N_20860,N_19946);
and U21256 (N_21256,N_19888,N_20861);
nand U21257 (N_21257,N_20533,N_20610);
nor U21258 (N_21258,N_20826,N_20423);
or U21259 (N_21259,N_20879,N_20266);
or U21260 (N_21260,N_19933,N_19611);
nand U21261 (N_21261,N_20121,N_19979);
and U21262 (N_21262,N_20979,N_19744);
or U21263 (N_21263,N_20328,N_19708);
and U21264 (N_21264,N_20217,N_19973);
or U21265 (N_21265,N_19834,N_20998);
nor U21266 (N_21266,N_20991,N_20063);
nand U21267 (N_21267,N_19556,N_20743);
nor U21268 (N_21268,N_20919,N_19649);
xor U21269 (N_21269,N_20113,N_19968);
xnor U21270 (N_21270,N_19557,N_20866);
nor U21271 (N_21271,N_20857,N_19984);
or U21272 (N_21272,N_20009,N_20494);
nor U21273 (N_21273,N_20251,N_19905);
xnor U21274 (N_21274,N_20478,N_20183);
xnor U21275 (N_21275,N_20886,N_20265);
nand U21276 (N_21276,N_19719,N_20915);
nor U21277 (N_21277,N_20830,N_20752);
nand U21278 (N_21278,N_20983,N_20791);
nor U21279 (N_21279,N_20239,N_20522);
nor U21280 (N_21280,N_20083,N_19575);
nor U21281 (N_21281,N_20657,N_20697);
nor U21282 (N_21282,N_20139,N_20295);
or U21283 (N_21283,N_19871,N_20340);
and U21284 (N_21284,N_19595,N_20104);
nor U21285 (N_21285,N_20582,N_20827);
or U21286 (N_21286,N_20250,N_20260);
nand U21287 (N_21287,N_20569,N_19931);
and U21288 (N_21288,N_20849,N_20234);
nand U21289 (N_21289,N_19660,N_20129);
xnor U21290 (N_21290,N_19892,N_19716);
nand U21291 (N_21291,N_20629,N_20314);
nor U21292 (N_21292,N_19588,N_19851);
xor U21293 (N_21293,N_20440,N_19745);
xor U21294 (N_21294,N_20720,N_19573);
or U21295 (N_21295,N_19540,N_19582);
and U21296 (N_21296,N_20588,N_19993);
and U21297 (N_21297,N_20165,N_20924);
nor U21298 (N_21298,N_20458,N_20227);
or U21299 (N_21299,N_19895,N_20895);
xor U21300 (N_21300,N_19938,N_20638);
xor U21301 (N_21301,N_20705,N_19536);
xor U21302 (N_21302,N_20885,N_19690);
xnor U21303 (N_21303,N_20688,N_20459);
and U21304 (N_21304,N_19983,N_20383);
or U21305 (N_21305,N_20643,N_19711);
nor U21306 (N_21306,N_20823,N_20980);
and U21307 (N_21307,N_20177,N_20202);
nor U21308 (N_21308,N_19598,N_19773);
or U21309 (N_21309,N_20802,N_20219);
nand U21310 (N_21310,N_20252,N_19914);
and U21311 (N_21311,N_20332,N_20282);
xor U21312 (N_21312,N_19784,N_20668);
nor U21313 (N_21313,N_20604,N_19910);
and U21314 (N_21314,N_19509,N_20510);
nor U21315 (N_21315,N_20767,N_20293);
or U21316 (N_21316,N_19520,N_20553);
xor U21317 (N_21317,N_20197,N_20056);
nand U21318 (N_21318,N_20341,N_20280);
and U21319 (N_21319,N_20044,N_19576);
and U21320 (N_21320,N_19960,N_20587);
and U21321 (N_21321,N_20855,N_20707);
xnor U21322 (N_21322,N_20808,N_20796);
xnor U21323 (N_21323,N_19647,N_20127);
nor U21324 (N_21324,N_19515,N_20702);
and U21325 (N_21325,N_20310,N_20064);
nor U21326 (N_21326,N_20003,N_20750);
xnor U21327 (N_21327,N_20070,N_20072);
or U21328 (N_21328,N_19809,N_20531);
or U21329 (N_21329,N_19558,N_20493);
nand U21330 (N_21330,N_20012,N_20993);
nor U21331 (N_21331,N_19785,N_19666);
or U21332 (N_21332,N_20898,N_19977);
xnor U21333 (N_21333,N_19753,N_19929);
or U21334 (N_21334,N_20026,N_20970);
nand U21335 (N_21335,N_20088,N_19735);
and U21336 (N_21336,N_20330,N_20969);
and U21337 (N_21337,N_20595,N_20572);
and U21338 (N_21338,N_20111,N_20078);
xnor U21339 (N_21339,N_19959,N_20573);
and U21340 (N_21340,N_20930,N_20746);
and U21341 (N_21341,N_20029,N_20352);
nor U21342 (N_21342,N_20313,N_20505);
or U21343 (N_21343,N_19793,N_20103);
nor U21344 (N_21344,N_20592,N_20470);
and U21345 (N_21345,N_20997,N_20717);
and U21346 (N_21346,N_20085,N_20686);
nand U21347 (N_21347,N_20447,N_19633);
and U21348 (N_21348,N_20317,N_20195);
xnor U21349 (N_21349,N_20122,N_19881);
and U21350 (N_21350,N_19635,N_20820);
nor U21351 (N_21351,N_19941,N_19902);
xnor U21352 (N_21352,N_20231,N_20495);
nor U21353 (N_21353,N_20832,N_20842);
or U21354 (N_21354,N_20642,N_20968);
nor U21355 (N_21355,N_20247,N_19721);
and U21356 (N_21356,N_20782,N_19860);
nand U21357 (N_21357,N_19790,N_20684);
nand U21358 (N_21358,N_20299,N_20790);
xor U21359 (N_21359,N_19574,N_20430);
nand U21360 (N_21360,N_20174,N_19610);
nand U21361 (N_21361,N_20537,N_20107);
nor U21362 (N_21362,N_19518,N_20396);
or U21363 (N_21363,N_19821,N_19763);
nand U21364 (N_21364,N_20963,N_20563);
nand U21365 (N_21365,N_20216,N_20598);
xnor U21366 (N_21366,N_19766,N_20995);
xor U21367 (N_21367,N_20422,N_19743);
or U21368 (N_21368,N_20813,N_19855);
or U21369 (N_21369,N_19655,N_20011);
nor U21370 (N_21370,N_19962,N_20648);
nor U21371 (N_21371,N_20967,N_20301);
nand U21372 (N_21372,N_19531,N_20098);
nand U21373 (N_21373,N_20320,N_20940);
nor U21374 (N_21374,N_20916,N_20990);
or U21375 (N_21375,N_20218,N_20461);
nand U21376 (N_21376,N_20848,N_20547);
and U21377 (N_21377,N_19779,N_20357);
nor U21378 (N_21378,N_20603,N_20455);
or U21379 (N_21379,N_19957,N_20730);
nor U21380 (N_21380,N_19912,N_20713);
nand U21381 (N_21381,N_20739,N_20670);
nor U21382 (N_21382,N_19950,N_20960);
and U21383 (N_21383,N_19729,N_20905);
nor U21384 (N_21384,N_20523,N_19527);
and U21385 (N_21385,N_20819,N_19616);
nor U21386 (N_21386,N_20168,N_20188);
and U21387 (N_21387,N_20994,N_20473);
and U21388 (N_21388,N_20362,N_20052);
nor U21389 (N_21389,N_19896,N_20166);
xor U21390 (N_21390,N_20840,N_20005);
nand U21391 (N_21391,N_20904,N_20161);
xor U21392 (N_21392,N_19754,N_20444);
nor U21393 (N_21393,N_19955,N_19537);
nand U21394 (N_21394,N_20057,N_20173);
nand U21395 (N_21395,N_19925,N_19545);
or U21396 (N_21396,N_20539,N_20824);
nor U21397 (N_21397,N_20809,N_20618);
xor U21398 (N_21398,N_20947,N_19579);
xnor U21399 (N_21399,N_20079,N_19513);
or U21400 (N_21400,N_20261,N_20828);
or U21401 (N_21401,N_20178,N_20210);
nand U21402 (N_21402,N_19839,N_19873);
nor U21403 (N_21403,N_20851,N_20092);
and U21404 (N_21404,N_19897,N_19553);
and U21405 (N_21405,N_20184,N_19835);
or U21406 (N_21406,N_20951,N_20706);
nand U21407 (N_21407,N_20781,N_20566);
or U21408 (N_21408,N_19681,N_20965);
nand U21409 (N_21409,N_20397,N_19641);
nor U21410 (N_21410,N_20654,N_20025);
or U21411 (N_21411,N_20978,N_19838);
nand U21412 (N_21412,N_20764,N_20345);
and U21413 (N_21413,N_20138,N_20436);
xor U21414 (N_21414,N_20017,N_19638);
and U21415 (N_21415,N_20463,N_20007);
nor U21416 (N_21416,N_20212,N_20039);
nand U21417 (N_21417,N_19771,N_20091);
xor U21418 (N_21418,N_19503,N_19783);
nand U21419 (N_21419,N_19794,N_19568);
nand U21420 (N_21420,N_19939,N_20617);
nor U21421 (N_21421,N_20507,N_20128);
nand U21422 (N_21422,N_19807,N_19764);
xnor U21423 (N_21423,N_20926,N_19630);
or U21424 (N_21424,N_20472,N_20095);
and U21425 (N_21425,N_20614,N_19712);
nand U21426 (N_21426,N_19767,N_20680);
xor U21427 (N_21427,N_20718,N_20441);
nor U21428 (N_21428,N_20729,N_19916);
xnor U21429 (N_21429,N_20515,N_19629);
and U21430 (N_21430,N_19731,N_20867);
and U21431 (N_21431,N_19919,N_19639);
nand U21432 (N_21432,N_19679,N_19631);
xor U21433 (N_21433,N_20048,N_19620);
xnor U21434 (N_21434,N_19782,N_20628);
and U21435 (N_21435,N_19697,N_20850);
nor U21436 (N_21436,N_20911,N_19619);
nor U21437 (N_21437,N_20502,N_20394);
nand U21438 (N_21438,N_20794,N_20376);
nor U21439 (N_21439,N_20681,N_20783);
nand U21440 (N_21440,N_19822,N_20637);
or U21441 (N_21441,N_19519,N_19501);
nand U21442 (N_21442,N_20806,N_20624);
and U21443 (N_21443,N_20778,N_20892);
nand U21444 (N_21444,N_20632,N_20016);
nor U21445 (N_21445,N_19644,N_20576);
nor U21446 (N_21446,N_19563,N_19991);
nor U21447 (N_21447,N_20425,N_19880);
or U21448 (N_21448,N_19963,N_19804);
nand U21449 (N_21449,N_19732,N_20693);
nand U21450 (N_21450,N_20259,N_20069);
nor U21451 (N_21451,N_20987,N_20590);
or U21452 (N_21452,N_19972,N_19915);
nor U21453 (N_21453,N_19692,N_19815);
and U21454 (N_21454,N_20971,N_19828);
nor U21455 (N_21455,N_20976,N_20269);
xnor U21456 (N_21456,N_19548,N_20770);
nor U21457 (N_21457,N_20475,N_19854);
xnor U21458 (N_21458,N_20241,N_20865);
nand U21459 (N_21459,N_20530,N_20913);
xnor U21460 (N_21460,N_20109,N_19601);
xnor U21461 (N_21461,N_20169,N_20596);
xnor U21462 (N_21462,N_20294,N_19755);
and U21463 (N_21463,N_20825,N_20917);
and U21464 (N_21464,N_19589,N_20243);
or U21465 (N_21465,N_20225,N_19698);
nand U21466 (N_21466,N_20822,N_20323);
nor U21467 (N_21467,N_20067,N_20945);
or U21468 (N_21468,N_19831,N_20874);
and U21469 (N_21469,N_20671,N_20818);
nor U21470 (N_21470,N_19969,N_20471);
nand U21471 (N_21471,N_19695,N_20407);
nor U21472 (N_21472,N_19674,N_20554);
nor U21473 (N_21473,N_19534,N_19861);
nand U21474 (N_21474,N_20223,N_20484);
nor U21475 (N_21475,N_20900,N_19561);
xor U21476 (N_21476,N_20329,N_20803);
and U21477 (N_21477,N_19942,N_20276);
nand U21478 (N_21478,N_19866,N_19512);
nand U21479 (N_21479,N_20439,N_20662);
nor U21480 (N_21480,N_20716,N_20918);
nor U21481 (N_21481,N_19757,N_20605);
or U21482 (N_21482,N_19648,N_19606);
xor U21483 (N_21483,N_20283,N_20766);
nand U21484 (N_21484,N_20401,N_20602);
and U21485 (N_21485,N_20146,N_20094);
nor U21486 (N_21486,N_19554,N_19500);
nor U21487 (N_21487,N_19725,N_20023);
xnor U21488 (N_21488,N_19948,N_20519);
or U21489 (N_21489,N_20201,N_20181);
nand U21490 (N_21490,N_20404,N_20742);
nor U21491 (N_21491,N_19749,N_20204);
and U21492 (N_21492,N_20896,N_20600);
or U21493 (N_21493,N_20700,N_19590);
nand U21494 (N_21494,N_20613,N_19529);
nand U21495 (N_21495,N_19614,N_19842);
and U21496 (N_21496,N_20405,N_20841);
or U21497 (N_21497,N_19981,N_19654);
or U21498 (N_21498,N_20303,N_20731);
xor U21499 (N_21499,N_20428,N_19715);
nand U21500 (N_21500,N_20361,N_20110);
xor U21501 (N_21501,N_19857,N_20371);
or U21502 (N_21502,N_20480,N_20496);
nand U21503 (N_21503,N_20772,N_19868);
nand U21504 (N_21504,N_20935,N_20956);
or U21505 (N_21505,N_20722,N_19626);
nand U21506 (N_21506,N_20413,N_20640);
nand U21507 (N_21507,N_20966,N_20368);
or U21508 (N_21508,N_20599,N_20555);
or U21509 (N_21509,N_19805,N_19736);
or U21510 (N_21510,N_20888,N_20524);
nand U21511 (N_21511,N_20042,N_20445);
nand U21512 (N_21512,N_20130,N_20167);
or U21513 (N_21513,N_20206,N_19811);
or U21514 (N_21514,N_20448,N_19894);
xor U21515 (N_21515,N_20661,N_20647);
nand U21516 (N_21516,N_19865,N_20759);
or U21517 (N_21517,N_19867,N_20801);
xor U21518 (N_21518,N_20046,N_19958);
nor U21519 (N_21519,N_20236,N_19953);
or U21520 (N_21520,N_19751,N_20365);
or U21521 (N_21521,N_20858,N_20123);
nand U21522 (N_21522,N_19817,N_19717);
and U21523 (N_21523,N_20925,N_19760);
xor U21524 (N_21524,N_19508,N_19670);
nor U21525 (N_21525,N_19516,N_19628);
and U21526 (N_21526,N_19874,N_19634);
nor U21527 (N_21527,N_20757,N_20676);
nand U21528 (N_21528,N_20562,N_20420);
xnor U21529 (N_21529,N_20137,N_19954);
and U21530 (N_21530,N_20359,N_20749);
nand U21531 (N_21531,N_20724,N_19664);
nor U21532 (N_21532,N_19618,N_19816);
xnor U21533 (N_21533,N_20589,N_19789);
and U21534 (N_21534,N_19812,N_19738);
nand U21535 (N_21535,N_19830,N_20392);
or U21536 (N_21536,N_20923,N_20049);
nand U21537 (N_21537,N_19818,N_20479);
nor U21538 (N_21538,N_20467,N_20549);
xnor U21539 (N_21539,N_20290,N_20780);
and U21540 (N_21540,N_20453,N_20347);
xnor U21541 (N_21541,N_20601,N_19583);
xor U21542 (N_21542,N_20431,N_20518);
or U21543 (N_21543,N_20263,N_20959);
nor U21544 (N_21544,N_20612,N_20356);
and U21545 (N_21545,N_19615,N_19549);
and U21546 (N_21546,N_20937,N_20390);
nand U21547 (N_21547,N_19691,N_19562);
or U21548 (N_21548,N_20798,N_19820);
and U21549 (N_21549,N_19747,N_20525);
xor U21550 (N_21550,N_19840,N_20300);
nand U21551 (N_21551,N_19646,N_20322);
and U21552 (N_21552,N_20304,N_20353);
nand U21553 (N_21553,N_20784,N_20665);
nand U21554 (N_21554,N_20773,N_19889);
and U21555 (N_21555,N_20529,N_19787);
xor U21556 (N_21556,N_20909,N_20172);
nor U21557 (N_21557,N_20508,N_20108);
xor U21558 (N_21558,N_19538,N_20890);
or U21559 (N_21559,N_20450,N_20950);
xnor U21560 (N_21560,N_19703,N_20883);
or U21561 (N_21561,N_20421,N_20696);
xnor U21562 (N_21562,N_20795,N_20489);
or U21563 (N_21563,N_19645,N_19600);
or U21564 (N_21564,N_20325,N_20082);
and U21565 (N_21565,N_20438,N_19714);
nand U21566 (N_21566,N_19581,N_20957);
nor U21567 (N_21567,N_20284,N_19718);
nand U21568 (N_21568,N_20882,N_19934);
xor U21569 (N_21569,N_19532,N_20584);
xor U21570 (N_21570,N_19656,N_19759);
or U21571 (N_21571,N_20732,N_19762);
nor U21572 (N_21572,N_20375,N_20635);
nand U21573 (N_21573,N_20278,N_19663);
nand U21574 (N_21574,N_20999,N_20101);
nor U21575 (N_21575,N_20621,N_19945);
nor U21576 (N_21576,N_19546,N_20355);
or U21577 (N_21577,N_19625,N_19668);
xnor U21578 (N_21578,N_20852,N_20512);
or U21579 (N_21579,N_20254,N_19586);
nor U21580 (N_21580,N_20675,N_20377);
or U21581 (N_21581,N_20426,N_19569);
nor U21582 (N_21582,N_20864,N_20932);
nand U21583 (N_21583,N_20372,N_19788);
xor U21584 (N_21584,N_20677,N_19999);
or U21585 (N_21585,N_20835,N_19624);
or U21586 (N_21586,N_20454,N_20106);
xor U21587 (N_21587,N_20235,N_20921);
or U21588 (N_21588,N_20364,N_20032);
nor U21589 (N_21589,N_20437,N_19566);
or U21590 (N_21590,N_20296,N_20384);
nor U21591 (N_21591,N_20386,N_20446);
or U21592 (N_21592,N_20615,N_19578);
nor U21593 (N_21593,N_19862,N_19909);
and U21594 (N_21594,N_20034,N_20817);
and U21595 (N_21595,N_20946,N_19858);
and U21596 (N_21596,N_20481,N_20503);
nor U21597 (N_21597,N_19943,N_19510);
nand U21598 (N_21598,N_20989,N_20474);
or U21599 (N_21599,N_20908,N_19786);
xnor U21600 (N_21600,N_20334,N_19952);
nand U21601 (N_21601,N_19978,N_19653);
and U21602 (N_21602,N_20961,N_19720);
nand U21603 (N_21603,N_20733,N_20443);
nor U21604 (N_21604,N_20087,N_20257);
and U21605 (N_21605,N_20800,N_19726);
nor U21606 (N_21606,N_20395,N_20175);
or U21607 (N_21607,N_20179,N_20388);
nor U21608 (N_21608,N_20077,N_19734);
nor U21609 (N_21609,N_20756,N_19608);
and U21610 (N_21610,N_20221,N_20432);
or U21611 (N_21611,N_20986,N_20151);
nor U21612 (N_21612,N_20977,N_20556);
xor U21613 (N_21613,N_19617,N_19926);
and U21614 (N_21614,N_20409,N_20863);
nand U21615 (N_21615,N_19730,N_19803);
nand U21616 (N_21616,N_19992,N_20360);
and U21617 (N_21617,N_20081,N_20575);
and U21618 (N_21618,N_19596,N_20762);
nor U21619 (N_21619,N_19623,N_20893);
and U21620 (N_21620,N_20740,N_19937);
and U21621 (N_21621,N_20736,N_20541);
nor U21622 (N_21622,N_20674,N_20689);
nor U21623 (N_21623,N_20528,N_20974);
or U21624 (N_21624,N_19778,N_19684);
or U21625 (N_21625,N_19836,N_20755);
nor U21626 (N_21626,N_20008,N_20646);
xnor U21627 (N_21627,N_19742,N_19505);
or U21628 (N_21628,N_20429,N_19890);
and U21629 (N_21629,N_20506,N_20033);
nand U21630 (N_21630,N_20532,N_19526);
nand U21631 (N_21631,N_19636,N_20540);
and U21632 (N_21632,N_19951,N_20133);
nor U21633 (N_21633,N_19609,N_20339);
xnor U21634 (N_21634,N_20812,N_20875);
or U21635 (N_21635,N_20843,N_20847);
and U21636 (N_21636,N_20627,N_19911);
or U21637 (N_21637,N_19571,N_20785);
xnor U21638 (N_21638,N_20144,N_19593);
or U21639 (N_21639,N_19506,N_20116);
xor U21640 (N_21640,N_20229,N_19966);
nor U21641 (N_21641,N_19667,N_19584);
nor U21642 (N_21642,N_20427,N_19524);
xor U21643 (N_21643,N_19922,N_20836);
and U21644 (N_21644,N_20059,N_20306);
or U21645 (N_21645,N_20289,N_20952);
or U21646 (N_21646,N_20055,N_19975);
and U21647 (N_21647,N_20271,N_20366);
or U21648 (N_21648,N_20859,N_20112);
nor U21649 (N_21649,N_20548,N_19900);
and U21650 (N_21650,N_20291,N_20821);
or U21651 (N_21651,N_20159,N_20041);
and U21652 (N_21652,N_20814,N_19728);
nor U21653 (N_21653,N_20776,N_19552);
nand U21654 (N_21654,N_20870,N_19825);
or U21655 (N_21655,N_20611,N_19856);
or U21656 (N_21656,N_19632,N_20062);
and U21657 (N_21657,N_20275,N_19980);
or U21658 (N_21658,N_20792,N_20639);
nand U21659 (N_21659,N_20363,N_20552);
xnor U21660 (N_21660,N_20811,N_20482);
nor U21661 (N_21661,N_19637,N_19772);
and U21662 (N_21662,N_20255,N_19770);
xor U21663 (N_21663,N_19832,N_19523);
nor U21664 (N_21664,N_20559,N_20829);
xnor U21665 (N_21665,N_20845,N_20226);
and U21666 (N_21666,N_20399,N_20469);
nand U21667 (N_21667,N_20807,N_19669);
xnor U21668 (N_21668,N_20897,N_19886);
nor U21669 (N_21669,N_20902,N_20745);
nor U21670 (N_21670,N_19990,N_20708);
nand U21671 (N_21671,N_20834,N_19961);
xor U21672 (N_21672,N_20889,N_19883);
or U21673 (N_21673,N_20090,N_20002);
or U21674 (N_21674,N_19685,N_20748);
xnor U21675 (N_21675,N_19917,N_20786);
or U21676 (N_21676,N_20456,N_20837);
xor U21677 (N_21677,N_19876,N_20120);
or U21678 (N_21678,N_19535,N_19702);
or U21679 (N_21679,N_20719,N_20292);
xnor U21680 (N_21680,N_20608,N_20741);
and U21681 (N_21681,N_20715,N_19533);
or U21682 (N_21682,N_20910,N_19746);
xor U21683 (N_21683,N_20074,N_20634);
nor U21684 (N_21684,N_20673,N_20839);
and U21685 (N_21685,N_20460,N_20869);
nor U21686 (N_21686,N_19525,N_20076);
nand U21687 (N_21687,N_20156,N_20140);
or U21688 (N_21688,N_19688,N_19777);
and U21689 (N_21689,N_19813,N_19879);
and U21690 (N_21690,N_20691,N_20931);
and U21691 (N_21691,N_20565,N_20606);
nor U21692 (N_21692,N_20854,N_20477);
xnor U21693 (N_21693,N_20249,N_20527);
nand U21694 (N_21694,N_20086,N_19899);
nor U21695 (N_21695,N_19940,N_19908);
and U21696 (N_21696,N_20021,N_20211);
and U21697 (N_21697,N_20203,N_20152);
xnor U21698 (N_21698,N_20804,N_20483);
or U21699 (N_21699,N_20491,N_20135);
or U21700 (N_21700,N_20163,N_20711);
nor U21701 (N_21701,N_19878,N_20222);
nor U21702 (N_21702,N_20153,N_20660);
or U21703 (N_21703,N_19700,N_20683);
nor U21704 (N_21704,N_19652,N_20728);
nand U21705 (N_21705,N_19607,N_20920);
nor U21706 (N_21706,N_20871,N_20170);
nand U21707 (N_21707,N_19550,N_20734);
nor U21708 (N_21708,N_20692,N_20545);
nand U21709 (N_21709,N_20651,N_19775);
nor U21710 (N_21710,N_20948,N_20534);
and U21711 (N_21711,N_20013,N_20350);
nor U21712 (N_21712,N_20981,N_20096);
nand U21713 (N_21713,N_20035,N_20609);
nand U21714 (N_21714,N_20232,N_20036);
nand U21715 (N_21715,N_20246,N_19543);
and U21716 (N_21716,N_20597,N_19965);
xor U21717 (N_21717,N_20570,N_19801);
nor U21718 (N_21718,N_20285,N_20381);
nand U21719 (N_21719,N_20380,N_20779);
nand U21720 (N_21720,N_19704,N_19661);
or U21721 (N_21721,N_20126,N_19675);
and U21722 (N_21722,N_20244,N_20050);
nand U21723 (N_21723,N_19551,N_20487);
or U21724 (N_21724,N_20663,N_19845);
nand U21725 (N_21725,N_19956,N_20972);
and U21726 (N_21726,N_19605,N_20616);
nand U21727 (N_21727,N_19577,N_20567);
nor U21728 (N_21728,N_20348,N_20679);
and U21729 (N_21729,N_20075,N_19768);
or U21730 (N_21730,N_20687,N_19827);
nand U21731 (N_21731,N_19995,N_20872);
nand U21732 (N_21732,N_19521,N_19872);
or U21733 (N_21733,N_20309,N_20623);
xor U21734 (N_21734,N_19591,N_20868);
or U21735 (N_21735,N_20644,N_20442);
nor U21736 (N_21736,N_20412,N_20089);
nand U21737 (N_21737,N_19658,N_20954);
or U21738 (N_21738,N_20237,N_20006);
and U21739 (N_21739,N_19528,N_20208);
nor U21740 (N_21740,N_20664,N_19774);
xor U21741 (N_21741,N_19923,N_19761);
nand U21742 (N_21742,N_20157,N_20043);
nor U21743 (N_21743,N_20416,N_20305);
nor U21744 (N_21744,N_20351,N_19706);
nand U21745 (N_21745,N_20230,N_20500);
xor U21746 (N_21746,N_19651,N_19594);
xor U21747 (N_21747,N_20097,N_19640);
nand U21748 (N_21748,N_20349,N_20738);
nand U21749 (N_21749,N_20726,N_20344);
and U21750 (N_21750,N_19613,N_20921);
xnor U21751 (N_21751,N_20839,N_20707);
nand U21752 (N_21752,N_20095,N_20091);
nor U21753 (N_21753,N_20987,N_20266);
and U21754 (N_21754,N_19976,N_20748);
and U21755 (N_21755,N_19605,N_20387);
or U21756 (N_21756,N_19947,N_19677);
nand U21757 (N_21757,N_20647,N_19666);
or U21758 (N_21758,N_20592,N_20133);
xor U21759 (N_21759,N_20915,N_20027);
nand U21760 (N_21760,N_20259,N_20811);
nand U21761 (N_21761,N_20888,N_20822);
xor U21762 (N_21762,N_20832,N_20027);
or U21763 (N_21763,N_20699,N_19662);
or U21764 (N_21764,N_19537,N_19564);
nor U21765 (N_21765,N_19997,N_20810);
nor U21766 (N_21766,N_20932,N_20755);
nand U21767 (N_21767,N_20190,N_20210);
nand U21768 (N_21768,N_20720,N_19932);
and U21769 (N_21769,N_19667,N_20205);
xor U21770 (N_21770,N_20680,N_20187);
and U21771 (N_21771,N_19655,N_20266);
and U21772 (N_21772,N_20847,N_20103);
and U21773 (N_21773,N_20126,N_20389);
xnor U21774 (N_21774,N_20153,N_19636);
nand U21775 (N_21775,N_20788,N_19506);
or U21776 (N_21776,N_20382,N_20941);
or U21777 (N_21777,N_19591,N_20860);
or U21778 (N_21778,N_19557,N_19678);
xor U21779 (N_21779,N_20081,N_19682);
xnor U21780 (N_21780,N_20128,N_20633);
and U21781 (N_21781,N_20705,N_20985);
nor U21782 (N_21782,N_20768,N_20586);
nand U21783 (N_21783,N_19569,N_20756);
xor U21784 (N_21784,N_20827,N_19955);
xnor U21785 (N_21785,N_20647,N_20530);
nand U21786 (N_21786,N_19835,N_20367);
nor U21787 (N_21787,N_20277,N_20290);
nor U21788 (N_21788,N_20061,N_20753);
and U21789 (N_21789,N_20515,N_19812);
nand U21790 (N_21790,N_20623,N_20332);
and U21791 (N_21791,N_20742,N_20287);
and U21792 (N_21792,N_19634,N_20166);
nor U21793 (N_21793,N_20730,N_20882);
and U21794 (N_21794,N_20375,N_20026);
or U21795 (N_21795,N_20255,N_20644);
or U21796 (N_21796,N_19822,N_19961);
or U21797 (N_21797,N_20988,N_20171);
nor U21798 (N_21798,N_19961,N_20863);
nand U21799 (N_21799,N_20125,N_20648);
nor U21800 (N_21800,N_20198,N_20300);
and U21801 (N_21801,N_20290,N_19880);
xnor U21802 (N_21802,N_19906,N_20072);
or U21803 (N_21803,N_20755,N_20901);
and U21804 (N_21804,N_19946,N_19901);
nand U21805 (N_21805,N_19544,N_19589);
xnor U21806 (N_21806,N_20432,N_20930);
xor U21807 (N_21807,N_20034,N_20730);
nor U21808 (N_21808,N_20652,N_19843);
xnor U21809 (N_21809,N_20811,N_19507);
nor U21810 (N_21810,N_20843,N_20884);
or U21811 (N_21811,N_19935,N_20430);
nand U21812 (N_21812,N_20554,N_20336);
and U21813 (N_21813,N_19749,N_19707);
or U21814 (N_21814,N_20359,N_19661);
nand U21815 (N_21815,N_20799,N_20877);
or U21816 (N_21816,N_20211,N_19823);
xor U21817 (N_21817,N_20664,N_20657);
xor U21818 (N_21818,N_20419,N_19592);
xor U21819 (N_21819,N_20756,N_19656);
and U21820 (N_21820,N_20511,N_19584);
xnor U21821 (N_21821,N_20279,N_20049);
nand U21822 (N_21822,N_20758,N_19568);
nor U21823 (N_21823,N_19646,N_20850);
nand U21824 (N_21824,N_20986,N_20088);
and U21825 (N_21825,N_19939,N_20744);
xor U21826 (N_21826,N_19579,N_20245);
and U21827 (N_21827,N_20211,N_19959);
nor U21828 (N_21828,N_19953,N_19783);
or U21829 (N_21829,N_20049,N_20857);
nand U21830 (N_21830,N_19512,N_20392);
or U21831 (N_21831,N_20679,N_20328);
xor U21832 (N_21832,N_20676,N_20416);
nand U21833 (N_21833,N_19578,N_20961);
or U21834 (N_21834,N_20667,N_19861);
nand U21835 (N_21835,N_20811,N_20023);
nand U21836 (N_21836,N_20905,N_20346);
and U21837 (N_21837,N_20840,N_19949);
nand U21838 (N_21838,N_19572,N_19624);
nand U21839 (N_21839,N_20332,N_19896);
and U21840 (N_21840,N_20088,N_19909);
or U21841 (N_21841,N_20322,N_20214);
nand U21842 (N_21842,N_19922,N_20938);
or U21843 (N_21843,N_20453,N_20385);
nand U21844 (N_21844,N_20295,N_19724);
nor U21845 (N_21845,N_20631,N_20093);
nand U21846 (N_21846,N_20883,N_20812);
xor U21847 (N_21847,N_20393,N_19572);
or U21848 (N_21848,N_20356,N_19965);
or U21849 (N_21849,N_19797,N_19889);
or U21850 (N_21850,N_20849,N_20305);
xnor U21851 (N_21851,N_20202,N_20827);
nand U21852 (N_21852,N_19665,N_19510);
and U21853 (N_21853,N_20521,N_20132);
xnor U21854 (N_21854,N_19788,N_19769);
nor U21855 (N_21855,N_19960,N_19937);
nor U21856 (N_21856,N_19975,N_20634);
nor U21857 (N_21857,N_19889,N_19842);
or U21858 (N_21858,N_19587,N_20505);
nor U21859 (N_21859,N_19927,N_20946);
or U21860 (N_21860,N_19970,N_20400);
nand U21861 (N_21861,N_19679,N_20397);
and U21862 (N_21862,N_20604,N_20673);
and U21863 (N_21863,N_20766,N_20887);
or U21864 (N_21864,N_20147,N_20159);
nor U21865 (N_21865,N_20141,N_20284);
nor U21866 (N_21866,N_20490,N_19592);
or U21867 (N_21867,N_20235,N_19607);
nand U21868 (N_21868,N_20092,N_20318);
and U21869 (N_21869,N_20819,N_20016);
xor U21870 (N_21870,N_20116,N_20307);
or U21871 (N_21871,N_20577,N_20963);
nand U21872 (N_21872,N_19800,N_19900);
and U21873 (N_21873,N_20217,N_19653);
and U21874 (N_21874,N_20541,N_20443);
nor U21875 (N_21875,N_20348,N_20103);
xor U21876 (N_21876,N_20785,N_19753);
and U21877 (N_21877,N_19755,N_20380);
xor U21878 (N_21878,N_20009,N_20845);
or U21879 (N_21879,N_20413,N_20425);
or U21880 (N_21880,N_19748,N_19742);
or U21881 (N_21881,N_20837,N_20197);
and U21882 (N_21882,N_20819,N_20531);
nand U21883 (N_21883,N_19916,N_20211);
and U21884 (N_21884,N_19597,N_19901);
or U21885 (N_21885,N_19646,N_19514);
xnor U21886 (N_21886,N_20762,N_20820);
xor U21887 (N_21887,N_20386,N_20297);
nand U21888 (N_21888,N_20563,N_19621);
nor U21889 (N_21889,N_20206,N_19698);
nand U21890 (N_21890,N_19892,N_19723);
and U21891 (N_21891,N_20812,N_20424);
and U21892 (N_21892,N_19956,N_20794);
nand U21893 (N_21893,N_20051,N_20186);
nand U21894 (N_21894,N_20569,N_19867);
xor U21895 (N_21895,N_20029,N_20534);
xnor U21896 (N_21896,N_20402,N_19878);
nor U21897 (N_21897,N_20458,N_19586);
nand U21898 (N_21898,N_19557,N_19643);
nor U21899 (N_21899,N_19589,N_20260);
and U21900 (N_21900,N_20710,N_20447);
nand U21901 (N_21901,N_19729,N_19521);
or U21902 (N_21902,N_19909,N_20701);
nor U21903 (N_21903,N_19964,N_20270);
or U21904 (N_21904,N_20899,N_19512);
xor U21905 (N_21905,N_20629,N_20437);
and U21906 (N_21906,N_20786,N_20282);
or U21907 (N_21907,N_20672,N_20263);
nand U21908 (N_21908,N_20734,N_20014);
nor U21909 (N_21909,N_20197,N_20717);
nand U21910 (N_21910,N_19829,N_20023);
or U21911 (N_21911,N_20337,N_20189);
nor U21912 (N_21912,N_20833,N_20454);
or U21913 (N_21913,N_19765,N_20385);
and U21914 (N_21914,N_19815,N_19856);
nor U21915 (N_21915,N_19654,N_20321);
nor U21916 (N_21916,N_20920,N_20270);
nor U21917 (N_21917,N_20207,N_19837);
xor U21918 (N_21918,N_19951,N_20019);
xnor U21919 (N_21919,N_19807,N_20175);
and U21920 (N_21920,N_19836,N_19947);
nand U21921 (N_21921,N_20424,N_20800);
nor U21922 (N_21922,N_20038,N_20924);
or U21923 (N_21923,N_19920,N_19786);
nand U21924 (N_21924,N_20233,N_20658);
nor U21925 (N_21925,N_19530,N_20682);
or U21926 (N_21926,N_19913,N_19506);
and U21927 (N_21927,N_19961,N_20992);
or U21928 (N_21928,N_20264,N_20084);
or U21929 (N_21929,N_20862,N_19601);
or U21930 (N_21930,N_20257,N_20749);
and U21931 (N_21931,N_20325,N_20480);
nand U21932 (N_21932,N_19746,N_20800);
nor U21933 (N_21933,N_20087,N_19993);
nor U21934 (N_21934,N_20532,N_20490);
nand U21935 (N_21935,N_20971,N_20038);
or U21936 (N_21936,N_20147,N_19518);
and U21937 (N_21937,N_20007,N_19696);
nor U21938 (N_21938,N_20821,N_20018);
or U21939 (N_21939,N_20680,N_20545);
or U21940 (N_21940,N_20054,N_19888);
nor U21941 (N_21941,N_20017,N_20400);
and U21942 (N_21942,N_20493,N_20955);
xnor U21943 (N_21943,N_19956,N_19546);
or U21944 (N_21944,N_20544,N_20262);
nand U21945 (N_21945,N_20930,N_19813);
or U21946 (N_21946,N_19897,N_20995);
nor U21947 (N_21947,N_20424,N_19790);
or U21948 (N_21948,N_20884,N_20109);
and U21949 (N_21949,N_20751,N_20273);
and U21950 (N_21950,N_20503,N_20251);
nor U21951 (N_21951,N_20396,N_20374);
nor U21952 (N_21952,N_20634,N_19854);
and U21953 (N_21953,N_19925,N_20749);
and U21954 (N_21954,N_19705,N_20916);
or U21955 (N_21955,N_19750,N_19542);
nor U21956 (N_21956,N_19948,N_19917);
and U21957 (N_21957,N_20626,N_20349);
or U21958 (N_21958,N_20694,N_19669);
and U21959 (N_21959,N_19531,N_19957);
nor U21960 (N_21960,N_19912,N_20661);
xor U21961 (N_21961,N_20783,N_20412);
xnor U21962 (N_21962,N_20547,N_19624);
and U21963 (N_21963,N_19720,N_20284);
nor U21964 (N_21964,N_20512,N_20585);
and U21965 (N_21965,N_19502,N_20880);
nor U21966 (N_21966,N_19583,N_20357);
or U21967 (N_21967,N_19788,N_20711);
nor U21968 (N_21968,N_20992,N_19554);
and U21969 (N_21969,N_20634,N_19514);
and U21970 (N_21970,N_20762,N_19969);
nor U21971 (N_21971,N_19526,N_19727);
or U21972 (N_21972,N_20319,N_20387);
and U21973 (N_21973,N_20221,N_20656);
xnor U21974 (N_21974,N_20895,N_20344);
nand U21975 (N_21975,N_20181,N_20050);
and U21976 (N_21976,N_20372,N_20859);
nor U21977 (N_21977,N_20410,N_19702);
and U21978 (N_21978,N_20881,N_19767);
or U21979 (N_21979,N_19909,N_20231);
nand U21980 (N_21980,N_20961,N_20081);
nor U21981 (N_21981,N_20975,N_19768);
nor U21982 (N_21982,N_20285,N_20622);
nor U21983 (N_21983,N_19812,N_19876);
or U21984 (N_21984,N_20532,N_19628);
or U21985 (N_21985,N_20469,N_20681);
nor U21986 (N_21986,N_20589,N_19643);
nand U21987 (N_21987,N_19532,N_20093);
xnor U21988 (N_21988,N_20443,N_20784);
or U21989 (N_21989,N_20800,N_20817);
xor U21990 (N_21990,N_19954,N_19703);
or U21991 (N_21991,N_19671,N_19873);
or U21992 (N_21992,N_20413,N_20442);
nor U21993 (N_21993,N_20136,N_20840);
and U21994 (N_21994,N_20010,N_20573);
xor U21995 (N_21995,N_20299,N_20091);
or U21996 (N_21996,N_20516,N_20524);
nand U21997 (N_21997,N_19534,N_19541);
nand U21998 (N_21998,N_20382,N_19758);
xor U21999 (N_21999,N_19622,N_20548);
or U22000 (N_22000,N_20795,N_20366);
or U22001 (N_22001,N_20518,N_20275);
nor U22002 (N_22002,N_19633,N_19974);
nand U22003 (N_22003,N_19638,N_19853);
nand U22004 (N_22004,N_19979,N_20322);
nor U22005 (N_22005,N_20602,N_20349);
nand U22006 (N_22006,N_20599,N_20999);
nor U22007 (N_22007,N_20229,N_19653);
nor U22008 (N_22008,N_20940,N_20171);
xor U22009 (N_22009,N_19970,N_20363);
nand U22010 (N_22010,N_20594,N_19658);
nor U22011 (N_22011,N_19801,N_20778);
nand U22012 (N_22012,N_19611,N_20278);
or U22013 (N_22013,N_19778,N_20456);
nor U22014 (N_22014,N_19599,N_19728);
nand U22015 (N_22015,N_20308,N_20645);
and U22016 (N_22016,N_20448,N_20239);
xnor U22017 (N_22017,N_20950,N_19998);
and U22018 (N_22018,N_20166,N_20741);
nand U22019 (N_22019,N_19813,N_20272);
or U22020 (N_22020,N_19987,N_19750);
nand U22021 (N_22021,N_20725,N_20014);
or U22022 (N_22022,N_20218,N_20393);
and U22023 (N_22023,N_20149,N_20379);
and U22024 (N_22024,N_20342,N_20762);
nand U22025 (N_22025,N_20870,N_19999);
xor U22026 (N_22026,N_20800,N_20620);
or U22027 (N_22027,N_20673,N_20492);
and U22028 (N_22028,N_19547,N_20628);
xnor U22029 (N_22029,N_19814,N_19766);
xor U22030 (N_22030,N_19557,N_20167);
nand U22031 (N_22031,N_20689,N_19526);
nand U22032 (N_22032,N_19860,N_19741);
or U22033 (N_22033,N_20933,N_20970);
and U22034 (N_22034,N_19879,N_20038);
and U22035 (N_22035,N_19677,N_19713);
nand U22036 (N_22036,N_19604,N_20151);
and U22037 (N_22037,N_20063,N_20310);
and U22038 (N_22038,N_20157,N_20689);
xnor U22039 (N_22039,N_19946,N_19848);
xnor U22040 (N_22040,N_19884,N_20745);
nor U22041 (N_22041,N_19903,N_19829);
or U22042 (N_22042,N_20825,N_20414);
and U22043 (N_22043,N_19835,N_19646);
and U22044 (N_22044,N_20689,N_20694);
nand U22045 (N_22045,N_20027,N_20534);
xnor U22046 (N_22046,N_20566,N_19612);
or U22047 (N_22047,N_19532,N_19777);
xnor U22048 (N_22048,N_20053,N_19947);
and U22049 (N_22049,N_20091,N_20793);
and U22050 (N_22050,N_20284,N_20866);
or U22051 (N_22051,N_19819,N_20357);
or U22052 (N_22052,N_20137,N_19714);
nand U22053 (N_22053,N_19699,N_19723);
nor U22054 (N_22054,N_20161,N_19971);
nor U22055 (N_22055,N_20608,N_20191);
or U22056 (N_22056,N_19906,N_20594);
nand U22057 (N_22057,N_19620,N_20390);
nand U22058 (N_22058,N_19951,N_20562);
and U22059 (N_22059,N_20096,N_19705);
nand U22060 (N_22060,N_20904,N_20608);
nor U22061 (N_22061,N_20404,N_20599);
xor U22062 (N_22062,N_20994,N_19985);
and U22063 (N_22063,N_19771,N_20707);
and U22064 (N_22064,N_20346,N_20940);
xor U22065 (N_22065,N_20043,N_20526);
nand U22066 (N_22066,N_19650,N_20052);
nand U22067 (N_22067,N_20357,N_20729);
and U22068 (N_22068,N_19910,N_20371);
xor U22069 (N_22069,N_20742,N_20541);
nor U22070 (N_22070,N_20949,N_20812);
nor U22071 (N_22071,N_20036,N_20416);
and U22072 (N_22072,N_20377,N_20164);
and U22073 (N_22073,N_20630,N_20529);
xor U22074 (N_22074,N_20815,N_19860);
or U22075 (N_22075,N_20981,N_20066);
or U22076 (N_22076,N_20092,N_20977);
nor U22077 (N_22077,N_20061,N_19791);
nand U22078 (N_22078,N_20396,N_20834);
nor U22079 (N_22079,N_20113,N_20942);
xor U22080 (N_22080,N_20766,N_20625);
or U22081 (N_22081,N_19725,N_20725);
or U22082 (N_22082,N_20827,N_20466);
nor U22083 (N_22083,N_20283,N_20546);
or U22084 (N_22084,N_20043,N_19789);
or U22085 (N_22085,N_19635,N_19957);
and U22086 (N_22086,N_20850,N_19977);
nor U22087 (N_22087,N_20752,N_20476);
nand U22088 (N_22088,N_20313,N_20042);
xnor U22089 (N_22089,N_19758,N_19792);
xor U22090 (N_22090,N_19960,N_20574);
nor U22091 (N_22091,N_19630,N_20712);
xor U22092 (N_22092,N_20071,N_20384);
nand U22093 (N_22093,N_19632,N_19775);
nand U22094 (N_22094,N_19882,N_19733);
nand U22095 (N_22095,N_20044,N_20583);
xnor U22096 (N_22096,N_20898,N_20996);
nand U22097 (N_22097,N_20456,N_19786);
xnor U22098 (N_22098,N_20828,N_20414);
nor U22099 (N_22099,N_20040,N_19659);
nand U22100 (N_22100,N_20096,N_20888);
and U22101 (N_22101,N_19993,N_20765);
nand U22102 (N_22102,N_20440,N_20216);
nand U22103 (N_22103,N_19870,N_19974);
xnor U22104 (N_22104,N_20553,N_19544);
nand U22105 (N_22105,N_20267,N_20487);
and U22106 (N_22106,N_20126,N_19834);
nand U22107 (N_22107,N_20919,N_20033);
and U22108 (N_22108,N_20032,N_20942);
or U22109 (N_22109,N_19996,N_19942);
and U22110 (N_22110,N_20786,N_19762);
nor U22111 (N_22111,N_20806,N_20717);
and U22112 (N_22112,N_20009,N_20188);
nand U22113 (N_22113,N_20723,N_20470);
and U22114 (N_22114,N_19999,N_20924);
nand U22115 (N_22115,N_20482,N_20772);
nand U22116 (N_22116,N_20237,N_20998);
nand U22117 (N_22117,N_20851,N_19792);
and U22118 (N_22118,N_20379,N_20084);
nor U22119 (N_22119,N_20608,N_20398);
xor U22120 (N_22120,N_20203,N_20305);
or U22121 (N_22121,N_19541,N_20095);
nor U22122 (N_22122,N_20460,N_19604);
nor U22123 (N_22123,N_19794,N_20839);
and U22124 (N_22124,N_20241,N_20073);
nor U22125 (N_22125,N_20567,N_19700);
or U22126 (N_22126,N_20308,N_20157);
nand U22127 (N_22127,N_20906,N_19847);
and U22128 (N_22128,N_20560,N_20849);
or U22129 (N_22129,N_20537,N_19538);
nor U22130 (N_22130,N_20752,N_19607);
or U22131 (N_22131,N_20172,N_19752);
or U22132 (N_22132,N_19590,N_20741);
or U22133 (N_22133,N_19635,N_20209);
xor U22134 (N_22134,N_20344,N_20141);
and U22135 (N_22135,N_19998,N_20319);
nand U22136 (N_22136,N_20303,N_19967);
nor U22137 (N_22137,N_19810,N_19929);
xor U22138 (N_22138,N_20647,N_20278);
xor U22139 (N_22139,N_20750,N_20339);
nand U22140 (N_22140,N_20958,N_20646);
nand U22141 (N_22141,N_20960,N_20133);
and U22142 (N_22142,N_20995,N_20525);
or U22143 (N_22143,N_20677,N_20725);
or U22144 (N_22144,N_19764,N_20405);
nand U22145 (N_22145,N_20160,N_20680);
nand U22146 (N_22146,N_19925,N_20603);
and U22147 (N_22147,N_19895,N_19797);
or U22148 (N_22148,N_19615,N_20040);
xnor U22149 (N_22149,N_20231,N_19768);
xnor U22150 (N_22150,N_20815,N_20081);
and U22151 (N_22151,N_19538,N_20367);
and U22152 (N_22152,N_20841,N_20157);
and U22153 (N_22153,N_20592,N_19612);
xor U22154 (N_22154,N_19522,N_20686);
nand U22155 (N_22155,N_19802,N_19889);
nand U22156 (N_22156,N_20105,N_20772);
or U22157 (N_22157,N_20812,N_19683);
nor U22158 (N_22158,N_20340,N_19691);
nor U22159 (N_22159,N_20585,N_20338);
and U22160 (N_22160,N_20118,N_20034);
nor U22161 (N_22161,N_19952,N_20658);
and U22162 (N_22162,N_19700,N_20787);
xnor U22163 (N_22163,N_19672,N_20790);
nor U22164 (N_22164,N_20314,N_20636);
xor U22165 (N_22165,N_19766,N_20159);
nand U22166 (N_22166,N_20327,N_19548);
nand U22167 (N_22167,N_20044,N_20326);
nand U22168 (N_22168,N_20518,N_20349);
or U22169 (N_22169,N_20938,N_20082);
or U22170 (N_22170,N_20840,N_19964);
or U22171 (N_22171,N_20194,N_19891);
or U22172 (N_22172,N_19903,N_20251);
nand U22173 (N_22173,N_20272,N_19654);
nand U22174 (N_22174,N_20912,N_19552);
xor U22175 (N_22175,N_19626,N_20399);
or U22176 (N_22176,N_19848,N_19875);
xor U22177 (N_22177,N_19778,N_19535);
xnor U22178 (N_22178,N_20848,N_20114);
nor U22179 (N_22179,N_20772,N_19611);
xnor U22180 (N_22180,N_20220,N_19853);
or U22181 (N_22181,N_20723,N_20648);
xnor U22182 (N_22182,N_20256,N_20571);
nor U22183 (N_22183,N_20950,N_20685);
nand U22184 (N_22184,N_19800,N_19541);
and U22185 (N_22185,N_20889,N_20237);
and U22186 (N_22186,N_19762,N_19905);
nand U22187 (N_22187,N_20605,N_20428);
nand U22188 (N_22188,N_20912,N_20626);
xor U22189 (N_22189,N_20192,N_20187);
nand U22190 (N_22190,N_20563,N_20697);
nor U22191 (N_22191,N_20497,N_20128);
and U22192 (N_22192,N_19790,N_20252);
and U22193 (N_22193,N_20154,N_20120);
xor U22194 (N_22194,N_20953,N_19798);
xor U22195 (N_22195,N_20304,N_20309);
xnor U22196 (N_22196,N_20143,N_20316);
and U22197 (N_22197,N_20476,N_20787);
xor U22198 (N_22198,N_20164,N_20182);
and U22199 (N_22199,N_20375,N_20633);
nor U22200 (N_22200,N_20750,N_20827);
xnor U22201 (N_22201,N_19771,N_20695);
xnor U22202 (N_22202,N_19725,N_19930);
xor U22203 (N_22203,N_20243,N_19832);
nand U22204 (N_22204,N_20017,N_20963);
xnor U22205 (N_22205,N_20767,N_19722);
xor U22206 (N_22206,N_20103,N_19505);
and U22207 (N_22207,N_20948,N_20531);
or U22208 (N_22208,N_20304,N_20491);
xor U22209 (N_22209,N_20413,N_20006);
and U22210 (N_22210,N_20608,N_20600);
nor U22211 (N_22211,N_20058,N_19622);
nand U22212 (N_22212,N_20990,N_20243);
nor U22213 (N_22213,N_19874,N_20520);
nand U22214 (N_22214,N_20313,N_19588);
and U22215 (N_22215,N_20801,N_19899);
or U22216 (N_22216,N_20731,N_20216);
or U22217 (N_22217,N_20799,N_20899);
and U22218 (N_22218,N_19856,N_19732);
and U22219 (N_22219,N_20165,N_20896);
or U22220 (N_22220,N_19723,N_20123);
and U22221 (N_22221,N_19685,N_19771);
and U22222 (N_22222,N_20379,N_20711);
nor U22223 (N_22223,N_19850,N_19507);
or U22224 (N_22224,N_20897,N_20274);
and U22225 (N_22225,N_20863,N_20660);
xor U22226 (N_22226,N_20984,N_20864);
and U22227 (N_22227,N_20331,N_20187);
and U22228 (N_22228,N_19713,N_20018);
and U22229 (N_22229,N_19965,N_20336);
xnor U22230 (N_22230,N_19504,N_19871);
nand U22231 (N_22231,N_19808,N_20509);
nand U22232 (N_22232,N_20560,N_19616);
and U22233 (N_22233,N_19792,N_20251);
and U22234 (N_22234,N_20849,N_20539);
nand U22235 (N_22235,N_19658,N_20413);
nor U22236 (N_22236,N_20172,N_19522);
and U22237 (N_22237,N_20635,N_20095);
nor U22238 (N_22238,N_20772,N_20330);
or U22239 (N_22239,N_20953,N_20687);
or U22240 (N_22240,N_20659,N_19563);
xnor U22241 (N_22241,N_19507,N_20784);
nand U22242 (N_22242,N_20370,N_19655);
xor U22243 (N_22243,N_20203,N_20548);
nand U22244 (N_22244,N_20480,N_19786);
and U22245 (N_22245,N_20089,N_20201);
or U22246 (N_22246,N_20161,N_20882);
and U22247 (N_22247,N_20873,N_19554);
and U22248 (N_22248,N_19837,N_20375);
nand U22249 (N_22249,N_19571,N_19502);
nor U22250 (N_22250,N_20919,N_20559);
xnor U22251 (N_22251,N_20750,N_19962);
and U22252 (N_22252,N_20267,N_19841);
xnor U22253 (N_22253,N_19769,N_20474);
and U22254 (N_22254,N_19792,N_20390);
xor U22255 (N_22255,N_20320,N_20838);
or U22256 (N_22256,N_20842,N_19908);
and U22257 (N_22257,N_20399,N_20355);
nand U22258 (N_22258,N_20193,N_19728);
nand U22259 (N_22259,N_20928,N_19872);
nand U22260 (N_22260,N_20624,N_19972);
nand U22261 (N_22261,N_20643,N_19529);
nor U22262 (N_22262,N_20561,N_20128);
nor U22263 (N_22263,N_20015,N_19841);
and U22264 (N_22264,N_19705,N_20323);
nand U22265 (N_22265,N_19555,N_20516);
or U22266 (N_22266,N_20703,N_20047);
and U22267 (N_22267,N_19973,N_20163);
xor U22268 (N_22268,N_20711,N_20359);
xnor U22269 (N_22269,N_20358,N_19955);
and U22270 (N_22270,N_20402,N_20704);
xnor U22271 (N_22271,N_20515,N_20036);
and U22272 (N_22272,N_20403,N_20537);
and U22273 (N_22273,N_20522,N_19739);
xnor U22274 (N_22274,N_20584,N_20108);
nand U22275 (N_22275,N_19791,N_19830);
nor U22276 (N_22276,N_20219,N_20631);
and U22277 (N_22277,N_19929,N_19734);
nand U22278 (N_22278,N_20690,N_20912);
nand U22279 (N_22279,N_19851,N_19738);
or U22280 (N_22280,N_20555,N_20699);
and U22281 (N_22281,N_19576,N_20445);
xnor U22282 (N_22282,N_20736,N_20396);
nand U22283 (N_22283,N_20658,N_19717);
or U22284 (N_22284,N_20898,N_20706);
nand U22285 (N_22285,N_20154,N_19514);
and U22286 (N_22286,N_19551,N_19638);
nand U22287 (N_22287,N_19920,N_20739);
nand U22288 (N_22288,N_20658,N_20904);
or U22289 (N_22289,N_20680,N_19519);
or U22290 (N_22290,N_20852,N_19724);
nand U22291 (N_22291,N_20512,N_19728);
and U22292 (N_22292,N_20077,N_20955);
xnor U22293 (N_22293,N_20706,N_19860);
and U22294 (N_22294,N_20284,N_19973);
nor U22295 (N_22295,N_20690,N_19603);
xor U22296 (N_22296,N_20505,N_20994);
nor U22297 (N_22297,N_19713,N_20977);
xor U22298 (N_22298,N_19607,N_19737);
nor U22299 (N_22299,N_20575,N_19526);
nand U22300 (N_22300,N_20089,N_20746);
or U22301 (N_22301,N_19546,N_19895);
or U22302 (N_22302,N_20903,N_19698);
or U22303 (N_22303,N_20844,N_20167);
nand U22304 (N_22304,N_20489,N_20960);
nand U22305 (N_22305,N_19585,N_20474);
and U22306 (N_22306,N_20296,N_20128);
nor U22307 (N_22307,N_20200,N_20250);
or U22308 (N_22308,N_20702,N_20634);
xor U22309 (N_22309,N_20739,N_20861);
nand U22310 (N_22310,N_20998,N_20299);
or U22311 (N_22311,N_19716,N_20397);
and U22312 (N_22312,N_20275,N_20403);
nor U22313 (N_22313,N_19842,N_19964);
nor U22314 (N_22314,N_20064,N_19653);
xnor U22315 (N_22315,N_20435,N_20889);
and U22316 (N_22316,N_20026,N_20309);
or U22317 (N_22317,N_20635,N_19670);
nand U22318 (N_22318,N_20853,N_20913);
xnor U22319 (N_22319,N_20007,N_20153);
xor U22320 (N_22320,N_20508,N_20657);
nor U22321 (N_22321,N_20590,N_19917);
xnor U22322 (N_22322,N_19721,N_20531);
nor U22323 (N_22323,N_20968,N_19569);
nor U22324 (N_22324,N_20043,N_19731);
nand U22325 (N_22325,N_19571,N_20762);
and U22326 (N_22326,N_19987,N_20335);
xor U22327 (N_22327,N_19873,N_20366);
or U22328 (N_22328,N_20198,N_20882);
and U22329 (N_22329,N_19654,N_20716);
nor U22330 (N_22330,N_20228,N_19796);
nand U22331 (N_22331,N_20494,N_19844);
and U22332 (N_22332,N_19726,N_20949);
and U22333 (N_22333,N_19744,N_20765);
xor U22334 (N_22334,N_20735,N_20784);
xor U22335 (N_22335,N_20812,N_19536);
and U22336 (N_22336,N_20468,N_20901);
xor U22337 (N_22337,N_19963,N_19821);
nor U22338 (N_22338,N_20361,N_20114);
or U22339 (N_22339,N_20312,N_20239);
and U22340 (N_22340,N_19549,N_19901);
nor U22341 (N_22341,N_19810,N_20582);
and U22342 (N_22342,N_20398,N_19635);
xnor U22343 (N_22343,N_20615,N_20570);
or U22344 (N_22344,N_20894,N_20591);
nand U22345 (N_22345,N_20392,N_19920);
nand U22346 (N_22346,N_20588,N_20931);
or U22347 (N_22347,N_19856,N_20974);
and U22348 (N_22348,N_20317,N_20863);
and U22349 (N_22349,N_19534,N_20224);
and U22350 (N_22350,N_19713,N_19621);
or U22351 (N_22351,N_19837,N_19601);
nor U22352 (N_22352,N_20717,N_20833);
or U22353 (N_22353,N_19835,N_19714);
or U22354 (N_22354,N_19792,N_20642);
or U22355 (N_22355,N_20335,N_20894);
nor U22356 (N_22356,N_20002,N_19808);
xor U22357 (N_22357,N_20336,N_20827);
and U22358 (N_22358,N_19897,N_20356);
and U22359 (N_22359,N_20966,N_20749);
nand U22360 (N_22360,N_19872,N_20397);
nor U22361 (N_22361,N_20691,N_20738);
nor U22362 (N_22362,N_20610,N_19968);
or U22363 (N_22363,N_20938,N_19626);
xnor U22364 (N_22364,N_20573,N_19738);
and U22365 (N_22365,N_20192,N_20528);
nor U22366 (N_22366,N_20921,N_20564);
and U22367 (N_22367,N_19614,N_19603);
nor U22368 (N_22368,N_20628,N_19964);
xnor U22369 (N_22369,N_20153,N_20885);
xnor U22370 (N_22370,N_20395,N_19851);
and U22371 (N_22371,N_20533,N_20835);
and U22372 (N_22372,N_19740,N_20820);
nand U22373 (N_22373,N_19506,N_20086);
and U22374 (N_22374,N_20529,N_20168);
xnor U22375 (N_22375,N_20894,N_20554);
or U22376 (N_22376,N_20739,N_20830);
or U22377 (N_22377,N_20677,N_20574);
nor U22378 (N_22378,N_19818,N_19784);
xnor U22379 (N_22379,N_20654,N_20828);
nor U22380 (N_22380,N_19880,N_20561);
xnor U22381 (N_22381,N_19591,N_19848);
or U22382 (N_22382,N_20108,N_19877);
and U22383 (N_22383,N_19689,N_20526);
nor U22384 (N_22384,N_20118,N_20572);
xnor U22385 (N_22385,N_20122,N_20144);
or U22386 (N_22386,N_19752,N_19811);
nor U22387 (N_22387,N_19568,N_19948);
nand U22388 (N_22388,N_20877,N_20633);
nand U22389 (N_22389,N_19978,N_20216);
or U22390 (N_22390,N_19627,N_20061);
and U22391 (N_22391,N_20095,N_20269);
or U22392 (N_22392,N_19716,N_19903);
and U22393 (N_22393,N_20681,N_20863);
xnor U22394 (N_22394,N_19968,N_20355);
xor U22395 (N_22395,N_19807,N_20984);
nor U22396 (N_22396,N_19553,N_19641);
nor U22397 (N_22397,N_20773,N_19817);
and U22398 (N_22398,N_20912,N_19682);
nor U22399 (N_22399,N_19627,N_20269);
or U22400 (N_22400,N_20122,N_20532);
nor U22401 (N_22401,N_20414,N_20204);
nor U22402 (N_22402,N_19931,N_20283);
or U22403 (N_22403,N_19953,N_19848);
nand U22404 (N_22404,N_20962,N_20195);
and U22405 (N_22405,N_20454,N_20914);
xnor U22406 (N_22406,N_20354,N_19892);
nor U22407 (N_22407,N_19638,N_20609);
nor U22408 (N_22408,N_20207,N_20422);
xnor U22409 (N_22409,N_20077,N_20186);
nor U22410 (N_22410,N_20291,N_19687);
or U22411 (N_22411,N_20749,N_20723);
or U22412 (N_22412,N_20659,N_19990);
nor U22413 (N_22413,N_20145,N_19604);
or U22414 (N_22414,N_19937,N_20852);
xnor U22415 (N_22415,N_20475,N_20794);
or U22416 (N_22416,N_20757,N_20216);
nor U22417 (N_22417,N_19767,N_19563);
nand U22418 (N_22418,N_20015,N_19752);
xnor U22419 (N_22419,N_20767,N_20433);
or U22420 (N_22420,N_20570,N_20883);
and U22421 (N_22421,N_19799,N_20709);
nand U22422 (N_22422,N_20287,N_19845);
or U22423 (N_22423,N_20612,N_19809);
and U22424 (N_22424,N_20087,N_20630);
nor U22425 (N_22425,N_20925,N_19766);
nor U22426 (N_22426,N_20552,N_19871);
or U22427 (N_22427,N_19900,N_20177);
nor U22428 (N_22428,N_19671,N_19660);
nand U22429 (N_22429,N_20143,N_20043);
and U22430 (N_22430,N_20770,N_19883);
xor U22431 (N_22431,N_20860,N_20528);
or U22432 (N_22432,N_20778,N_20558);
nor U22433 (N_22433,N_20884,N_20465);
or U22434 (N_22434,N_20228,N_20551);
nor U22435 (N_22435,N_19598,N_20310);
nand U22436 (N_22436,N_20391,N_20585);
nand U22437 (N_22437,N_19868,N_20388);
or U22438 (N_22438,N_20822,N_20084);
nor U22439 (N_22439,N_20362,N_20587);
or U22440 (N_22440,N_20955,N_19669);
xnor U22441 (N_22441,N_20044,N_20036);
nor U22442 (N_22442,N_19927,N_20468);
or U22443 (N_22443,N_19653,N_20930);
and U22444 (N_22444,N_19622,N_19963);
nor U22445 (N_22445,N_20320,N_20302);
xor U22446 (N_22446,N_20134,N_19716);
nor U22447 (N_22447,N_20014,N_19643);
and U22448 (N_22448,N_20489,N_19510);
and U22449 (N_22449,N_20292,N_20912);
or U22450 (N_22450,N_20641,N_20751);
nand U22451 (N_22451,N_20637,N_20174);
nor U22452 (N_22452,N_20293,N_20932);
nor U22453 (N_22453,N_20769,N_19606);
or U22454 (N_22454,N_20592,N_20677);
and U22455 (N_22455,N_19981,N_19670);
nand U22456 (N_22456,N_20164,N_20819);
and U22457 (N_22457,N_20018,N_20111);
nor U22458 (N_22458,N_20838,N_20386);
nand U22459 (N_22459,N_20365,N_20919);
nand U22460 (N_22460,N_19591,N_20679);
or U22461 (N_22461,N_19768,N_19616);
nand U22462 (N_22462,N_20105,N_20180);
and U22463 (N_22463,N_20300,N_20428);
nand U22464 (N_22464,N_20676,N_20684);
xnor U22465 (N_22465,N_19758,N_20354);
nor U22466 (N_22466,N_19977,N_20657);
nor U22467 (N_22467,N_20536,N_20451);
xnor U22468 (N_22468,N_19611,N_20118);
or U22469 (N_22469,N_19885,N_19974);
nor U22470 (N_22470,N_20191,N_19631);
xor U22471 (N_22471,N_20546,N_20839);
or U22472 (N_22472,N_19671,N_19559);
nand U22473 (N_22473,N_20480,N_20217);
nor U22474 (N_22474,N_20661,N_19949);
xor U22475 (N_22475,N_19857,N_20527);
nor U22476 (N_22476,N_19915,N_19660);
or U22477 (N_22477,N_19807,N_20462);
or U22478 (N_22478,N_20894,N_20713);
xnor U22479 (N_22479,N_20661,N_19677);
nand U22480 (N_22480,N_20084,N_20326);
and U22481 (N_22481,N_20307,N_20421);
xor U22482 (N_22482,N_19979,N_20205);
nor U22483 (N_22483,N_19851,N_19908);
nor U22484 (N_22484,N_19886,N_20023);
nand U22485 (N_22485,N_20023,N_20247);
or U22486 (N_22486,N_19521,N_20114);
and U22487 (N_22487,N_20286,N_19810);
or U22488 (N_22488,N_20931,N_20532);
nor U22489 (N_22489,N_20262,N_20699);
nand U22490 (N_22490,N_19828,N_19841);
nand U22491 (N_22491,N_19649,N_20909);
or U22492 (N_22492,N_19976,N_19750);
nor U22493 (N_22493,N_20879,N_19865);
nor U22494 (N_22494,N_19778,N_20357);
and U22495 (N_22495,N_20563,N_20603);
or U22496 (N_22496,N_20880,N_20673);
and U22497 (N_22497,N_19873,N_20081);
and U22498 (N_22498,N_20903,N_20734);
nand U22499 (N_22499,N_20742,N_20084);
xnor U22500 (N_22500,N_21976,N_21561);
nor U22501 (N_22501,N_21802,N_22394);
xor U22502 (N_22502,N_22144,N_22322);
xor U22503 (N_22503,N_21155,N_22486);
nor U22504 (N_22504,N_22065,N_21182);
xor U22505 (N_22505,N_22362,N_21456);
or U22506 (N_22506,N_22066,N_21143);
nor U22507 (N_22507,N_21839,N_21744);
nor U22508 (N_22508,N_21825,N_21911);
nand U22509 (N_22509,N_21464,N_21851);
or U22510 (N_22510,N_22437,N_22414);
xor U22511 (N_22511,N_22349,N_21909);
nor U22512 (N_22512,N_21245,N_21517);
and U22513 (N_22513,N_22265,N_22418);
or U22514 (N_22514,N_21715,N_21486);
nor U22515 (N_22515,N_21000,N_21535);
and U22516 (N_22516,N_22170,N_21208);
and U22517 (N_22517,N_22267,N_21429);
nor U22518 (N_22518,N_22431,N_21760);
and U22519 (N_22519,N_21427,N_21592);
nand U22520 (N_22520,N_22421,N_22413);
and U22521 (N_22521,N_21354,N_22270);
nand U22522 (N_22522,N_22031,N_21179);
nand U22523 (N_22523,N_22197,N_21952);
or U22524 (N_22524,N_22404,N_21366);
nor U22525 (N_22525,N_21930,N_21985);
or U22526 (N_22526,N_21250,N_22311);
nor U22527 (N_22527,N_22440,N_21872);
nor U22528 (N_22528,N_21448,N_22142);
nor U22529 (N_22529,N_21620,N_21521);
xor U22530 (N_22530,N_22117,N_21948);
or U22531 (N_22531,N_22386,N_21653);
or U22532 (N_22532,N_21614,N_21959);
or U22533 (N_22533,N_21165,N_21576);
nand U22534 (N_22534,N_21216,N_21738);
and U22535 (N_22535,N_21616,N_21575);
or U22536 (N_22536,N_22303,N_21044);
xor U22537 (N_22537,N_21322,N_22347);
and U22538 (N_22538,N_21281,N_22032);
and U22539 (N_22539,N_21038,N_21488);
and U22540 (N_22540,N_21794,N_21907);
nor U22541 (N_22541,N_22381,N_21944);
nor U22542 (N_22542,N_21654,N_21185);
and U22543 (N_22543,N_21373,N_21060);
or U22544 (N_22544,N_21124,N_22175);
nor U22545 (N_22545,N_21070,N_22183);
nor U22546 (N_22546,N_22126,N_21618);
nand U22547 (N_22547,N_21916,N_22106);
xor U22548 (N_22548,N_21398,N_22441);
or U22549 (N_22549,N_22121,N_21048);
nor U22550 (N_22550,N_21351,N_21924);
nand U22551 (N_22551,N_22056,N_21381);
nand U22552 (N_22552,N_21796,N_22368);
and U22553 (N_22553,N_22094,N_21438);
nand U22554 (N_22554,N_21742,N_22044);
xnor U22555 (N_22555,N_21819,N_21568);
nand U22556 (N_22556,N_21040,N_21200);
or U22557 (N_22557,N_22447,N_21183);
xnor U22558 (N_22558,N_21960,N_22231);
and U22559 (N_22559,N_21640,N_22184);
nand U22560 (N_22560,N_21021,N_21673);
nor U22561 (N_22561,N_22237,N_21626);
and U22562 (N_22562,N_21705,N_21524);
nand U22563 (N_22563,N_21827,N_22423);
xor U22564 (N_22564,N_21396,N_21873);
xor U22565 (N_22565,N_22340,N_21732);
or U22566 (N_22566,N_22427,N_22490);
xor U22567 (N_22567,N_21731,N_21162);
nor U22568 (N_22568,N_22107,N_22098);
nor U22569 (N_22569,N_21076,N_21718);
or U22570 (N_22570,N_22057,N_21706);
or U22571 (N_22571,N_21061,N_21422);
xor U22572 (N_22572,N_21650,N_22282);
nand U22573 (N_22573,N_21052,N_21018);
nand U22574 (N_22574,N_21262,N_21225);
or U22575 (N_22575,N_21558,N_21447);
nand U22576 (N_22576,N_21587,N_21619);
nor U22577 (N_22577,N_21666,N_22108);
nor U22578 (N_22578,N_21986,N_22238);
nor U22579 (N_22579,N_21067,N_22475);
and U22580 (N_22580,N_21158,N_21542);
nand U22581 (N_22581,N_22114,N_21609);
nand U22582 (N_22582,N_21117,N_22393);
nand U22583 (N_22583,N_21736,N_21147);
and U22584 (N_22584,N_21831,N_22015);
or U22585 (N_22585,N_22339,N_22296);
and U22586 (N_22586,N_22161,N_21865);
and U22587 (N_22587,N_21605,N_21292);
and U22588 (N_22588,N_21659,N_21947);
nand U22589 (N_22589,N_22116,N_22430);
and U22590 (N_22590,N_22239,N_21621);
xnor U22591 (N_22591,N_21334,N_21739);
or U22592 (N_22592,N_22172,N_22304);
and U22593 (N_22593,N_21312,N_21679);
or U22594 (N_22594,N_21353,N_21638);
xor U22595 (N_22595,N_21298,N_21681);
or U22596 (N_22596,N_21336,N_22289);
nor U22597 (N_22597,N_21215,N_21214);
xor U22598 (N_22598,N_21303,N_21707);
nor U22599 (N_22599,N_21552,N_21202);
and U22600 (N_22600,N_22030,N_21857);
nand U22601 (N_22601,N_22424,N_22467);
nand U22602 (N_22602,N_21495,N_21371);
xnor U22603 (N_22603,N_22281,N_21066);
nor U22604 (N_22604,N_21263,N_21917);
or U22605 (N_22605,N_21932,N_21601);
or U22606 (N_22606,N_21426,N_22152);
and U22607 (N_22607,N_21234,N_22016);
or U22608 (N_22608,N_21759,N_21982);
or U22609 (N_22609,N_21809,N_22343);
nand U22610 (N_22610,N_21277,N_21045);
xnor U22611 (N_22611,N_21166,N_21109);
and U22612 (N_22612,N_22089,N_21551);
nor U22613 (N_22613,N_22211,N_21062);
or U22614 (N_22614,N_22228,N_21583);
xor U22615 (N_22615,N_22224,N_21695);
or U22616 (N_22616,N_22253,N_21193);
and U22617 (N_22617,N_21218,N_21275);
nor U22618 (N_22618,N_21136,N_21417);
and U22619 (N_22619,N_21467,N_22489);
or U22620 (N_22620,N_21037,N_21461);
xor U22621 (N_22621,N_22190,N_21082);
and U22622 (N_22622,N_22261,N_22111);
and U22623 (N_22623,N_21305,N_22419);
and U22624 (N_22624,N_21380,N_22302);
or U22625 (N_22625,N_21157,N_21786);
nand U22626 (N_22626,N_22130,N_21129);
nor U22627 (N_22627,N_22492,N_22271);
and U22628 (N_22628,N_21163,N_21811);
nand U22629 (N_22629,N_21728,N_21748);
xor U22630 (N_22630,N_22084,N_21765);
or U22631 (N_22631,N_21132,N_21206);
and U22632 (N_22632,N_21964,N_22488);
nor U22633 (N_22633,N_22314,N_21347);
nand U22634 (N_22634,N_21570,N_21513);
nor U22635 (N_22635,N_21970,N_21005);
xor U22636 (N_22636,N_21957,N_21125);
or U22637 (N_22637,N_22319,N_22398);
nor U22638 (N_22638,N_21013,N_22298);
or U22639 (N_22639,N_22235,N_21041);
nand U22640 (N_22640,N_22064,N_22451);
and U22641 (N_22641,N_22179,N_21307);
xnor U22642 (N_22642,N_22168,N_22200);
or U22643 (N_22643,N_21914,N_21074);
nor U22644 (N_22644,N_22038,N_21936);
and U22645 (N_22645,N_21859,N_22443);
nor U22646 (N_22646,N_21400,N_22342);
nand U22647 (N_22647,N_21596,N_21327);
nor U22648 (N_22648,N_21606,N_22257);
nor U22649 (N_22649,N_21242,N_21012);
nand U22650 (N_22650,N_22025,N_22407);
nor U22651 (N_22651,N_21492,N_22035);
nand U22652 (N_22652,N_21801,N_21758);
nor U22653 (N_22653,N_22189,N_22405);
xnor U22654 (N_22654,N_22223,N_21671);
nor U22655 (N_22655,N_21852,N_22354);
nor U22656 (N_22656,N_21190,N_21780);
and U22657 (N_22657,N_22410,N_22273);
or U22658 (N_22658,N_21774,N_22350);
or U22659 (N_22659,N_21498,N_21409);
and U22660 (N_22660,N_21874,N_21266);
and U22661 (N_22661,N_21514,N_22454);
and U22662 (N_22662,N_22082,N_21823);
nor U22663 (N_22663,N_21686,N_22290);
xor U22664 (N_22664,N_22258,N_21485);
and U22665 (N_22665,N_21806,N_21028);
nor U22666 (N_22666,N_21634,N_21591);
nand U22667 (N_22667,N_21203,N_22051);
xor U22668 (N_22668,N_21384,N_21518);
or U22669 (N_22669,N_21478,N_21454);
nor U22670 (N_22670,N_21110,N_21466);
or U22671 (N_22671,N_21432,N_21978);
xnor U22672 (N_22672,N_21221,N_22165);
and U22673 (N_22673,N_21661,N_22387);
nor U22674 (N_22674,N_21435,N_22497);
and U22675 (N_22675,N_22462,N_21861);
and U22676 (N_22676,N_21308,N_21593);
nor U22677 (N_22677,N_22491,N_21364);
or U22678 (N_22678,N_22369,N_21643);
nor U22679 (N_22679,N_22213,N_21933);
or U22680 (N_22680,N_22070,N_21159);
nor U22681 (N_22681,N_22245,N_21608);
nand U22682 (N_22682,N_22146,N_22241);
nand U22683 (N_22683,N_21237,N_21582);
or U22684 (N_22684,N_21368,N_21047);
nand U22685 (N_22685,N_21553,N_22498);
nor U22686 (N_22686,N_21820,N_21459);
nand U22687 (N_22687,N_22396,N_22143);
nand U22688 (N_22688,N_21394,N_21385);
nor U22689 (N_22689,N_21479,N_22138);
xor U22690 (N_22690,N_21259,N_22352);
nand U22691 (N_22691,N_21154,N_21229);
or U22692 (N_22692,N_22049,N_21546);
xnor U22693 (N_22693,N_21311,N_21224);
and U22694 (N_22694,N_22156,N_21134);
nand U22695 (N_22695,N_21170,N_21764);
or U22696 (N_22696,N_21296,N_22206);
and U22697 (N_22697,N_21027,N_21714);
nor U22698 (N_22698,N_22356,N_22234);
nand U22699 (N_22699,N_21194,N_22359);
and U22700 (N_22700,N_22483,N_21902);
and U22701 (N_22701,N_21031,N_21137);
nand U22702 (N_22702,N_21847,N_21812);
xnor U22703 (N_22703,N_22309,N_22277);
nand U22704 (N_22704,N_21813,N_21104);
xor U22705 (N_22705,N_21330,N_22134);
nand U22706 (N_22706,N_22177,N_21362);
xnor U22707 (N_22707,N_21670,N_21176);
xnor U22708 (N_22708,N_21750,N_22099);
xor U22709 (N_22709,N_21449,N_21688);
nand U22710 (N_22710,N_21785,N_21669);
or U22711 (N_22711,N_22002,N_22353);
xnor U22712 (N_22712,N_22217,N_21006);
xor U22713 (N_22713,N_21273,N_21337);
xnor U22714 (N_22714,N_21854,N_22360);
or U22715 (N_22715,N_22220,N_21469);
xor U22716 (N_22716,N_22390,N_22422);
nand U22717 (N_22717,N_22485,N_22163);
or U22718 (N_22718,N_22214,N_21173);
or U22719 (N_22719,N_21710,N_21271);
xor U22720 (N_22720,N_21949,N_21174);
or U22721 (N_22721,N_21212,N_21822);
or U22722 (N_22722,N_21472,N_21642);
nor U22723 (N_22723,N_22375,N_21428);
and U22724 (N_22724,N_22230,N_22113);
nand U22725 (N_22725,N_21913,N_22433);
or U22726 (N_22726,N_22236,N_21268);
and U22727 (N_22727,N_22124,N_21776);
or U22728 (N_22728,N_22058,N_22254);
nor U22729 (N_22729,N_21995,N_21286);
or U22730 (N_22730,N_21629,N_21100);
or U22731 (N_22731,N_21545,N_21320);
nand U22732 (N_22732,N_22092,N_21101);
and U22733 (N_22733,N_21633,N_21589);
or U22734 (N_22734,N_22022,N_21317);
and U22735 (N_22735,N_21855,N_21664);
nor U22736 (N_22736,N_21191,N_22248);
and U22737 (N_22737,N_21232,N_21280);
and U22738 (N_22738,N_21999,N_21955);
and U22739 (N_22739,N_21815,N_22274);
or U22740 (N_22740,N_22009,N_21968);
and U22741 (N_22741,N_22147,N_21534);
nand U22742 (N_22742,N_21676,N_21934);
or U22743 (N_22743,N_22005,N_22305);
nor U22744 (N_22744,N_22425,N_21803);
xor U22745 (N_22745,N_21980,N_21572);
nand U22746 (N_22746,N_21723,N_22406);
nand U22747 (N_22747,N_21304,N_21578);
nand U22748 (N_22748,N_22382,N_21318);
nor U22749 (N_22749,N_21249,N_21029);
or U22750 (N_22750,N_22145,N_21864);
or U22751 (N_22751,N_22140,N_21075);
and U22752 (N_22752,N_22180,N_21489);
and U22753 (N_22753,N_21712,N_21397);
nand U22754 (N_22754,N_21319,N_21927);
nor U22755 (N_22755,N_21413,N_21630);
or U22756 (N_22756,N_21945,N_21555);
nand U22757 (N_22757,N_21243,N_21894);
or U22758 (N_22758,N_21525,N_21550);
nand U22759 (N_22759,N_21935,N_21260);
nor U22760 (N_22760,N_21443,N_22346);
or U22761 (N_22761,N_21512,N_21869);
nor U22762 (N_22762,N_21153,N_22389);
nand U22763 (N_22763,N_21356,N_22399);
nor U22764 (N_22764,N_21440,N_21265);
xor U22765 (N_22765,N_21554,N_21641);
nand U22766 (N_22766,N_22329,N_21991);
and U22767 (N_22767,N_21151,N_22203);
and U22768 (N_22768,N_21726,N_21925);
xnor U22769 (N_22769,N_21808,N_21341);
nand U22770 (N_22770,N_21846,N_21713);
nand U22771 (N_22771,N_21365,N_22090);
and U22772 (N_22772,N_21374,N_21310);
nand U22773 (N_22773,N_22464,N_21565);
nand U22774 (N_22774,N_21022,N_21150);
nand U22775 (N_22775,N_22208,N_21775);
nand U22776 (N_22776,N_21994,N_22370);
nor U22777 (N_22777,N_21848,N_22327);
nand U22778 (N_22778,N_22218,N_21223);
and U22779 (N_22779,N_21814,N_21735);
and U22780 (N_22780,N_21391,N_21657);
and U22781 (N_22781,N_22043,N_21187);
nand U22782 (N_22782,N_21511,N_21383);
or U22783 (N_22783,N_22045,N_21862);
xor U22784 (N_22784,N_21437,N_22028);
nand U22785 (N_22785,N_21821,N_21597);
or U22786 (N_22786,N_21624,N_22103);
nand U22787 (N_22787,N_21979,N_21975);
nor U22788 (N_22788,N_22412,N_22279);
nand U22789 (N_22789,N_21496,N_21425);
nor U22790 (N_22790,N_22076,N_22182);
or U22791 (N_22791,N_21007,N_21323);
and U22792 (N_22792,N_21720,N_21463);
or U22793 (N_22793,N_21008,N_21452);
or U22794 (N_22794,N_21126,N_21077);
and U22795 (N_22795,N_22000,N_21491);
or U22796 (N_22796,N_21983,N_21743);
nand U22797 (N_22797,N_21010,N_21559);
or U22798 (N_22798,N_21097,N_21787);
and U22799 (N_22799,N_22306,N_22215);
and U22800 (N_22800,N_21696,N_22008);
and U22801 (N_22801,N_21962,N_21315);
xnor U22802 (N_22802,N_21276,N_22104);
or U22803 (N_22803,N_21966,N_21886);
xor U22804 (N_22804,N_22465,N_21071);
nand U22805 (N_22805,N_21804,N_21716);
xor U22806 (N_22806,N_22122,N_22320);
and U22807 (N_22807,N_22243,N_22307);
nor U22808 (N_22808,N_21526,N_21091);
nor U22809 (N_22809,N_21717,N_21595);
and U22810 (N_22810,N_21344,N_21003);
xnor U22811 (N_22811,N_21210,N_21078);
xnor U22812 (N_22812,N_21516,N_21080);
and U22813 (N_22813,N_21784,N_22110);
and U22814 (N_22814,N_22039,N_21833);
nand U22815 (N_22815,N_22449,N_21842);
nor U22816 (N_22816,N_21046,N_21988);
nand U22817 (N_22817,N_21014,N_21256);
or U22818 (N_22818,N_21617,N_21974);
or U22819 (N_22819,N_21668,N_22366);
nand U22820 (N_22820,N_22242,N_21788);
and U22821 (N_22821,N_21015,N_21025);
xor U22822 (N_22822,N_22364,N_21520);
xor U22823 (N_22823,N_21761,N_21625);
nor U22824 (N_22824,N_21415,N_21849);
and U22825 (N_22825,N_21387,N_21339);
and U22826 (N_22826,N_22021,N_21049);
or U22827 (N_22827,N_21594,N_21752);
and U22828 (N_22828,N_22335,N_21628);
or U22829 (N_22829,N_22194,N_22264);
and U22830 (N_22830,N_22154,N_22232);
nand U22831 (N_22831,N_21611,N_22119);
nor U22832 (N_22832,N_21441,N_21252);
and U22833 (N_22833,N_21908,N_22434);
or U22834 (N_22834,N_21378,N_22326);
nand U22835 (N_22835,N_21832,N_22363);
or U22836 (N_22836,N_22365,N_21816);
nor U22837 (N_22837,N_21471,N_21416);
nor U22838 (N_22838,N_22063,N_22033);
nor U22839 (N_22839,N_22409,N_21433);
nor U22840 (N_22840,N_22436,N_21270);
or U22841 (N_22841,N_21161,N_21401);
nand U22842 (N_22842,N_22323,N_21128);
xor U22843 (N_22843,N_21928,N_21093);
nor U22844 (N_22844,N_21209,N_21294);
xnor U22845 (N_22845,N_21211,N_21922);
nor U22846 (N_22846,N_21703,N_21584);
nor U22847 (N_22847,N_21531,N_21557);
and U22848 (N_22848,N_21325,N_21051);
nor U22849 (N_22849,N_21897,N_21663);
or U22850 (N_22850,N_22459,N_21904);
nand U22851 (N_22851,N_22071,N_21658);
xnor U22852 (N_22852,N_21749,N_21637);
or U22853 (N_22853,N_21369,N_21141);
xnor U22854 (N_22854,N_21411,N_21901);
xor U22855 (N_22855,N_22037,N_21420);
xor U22856 (N_22856,N_21783,N_21042);
nand U22857 (N_22857,N_21841,N_21453);
nand U22858 (N_22858,N_21410,N_22061);
nor U22859 (N_22859,N_21768,N_22402);
and U22860 (N_22860,N_21474,N_21455);
xor U22861 (N_22861,N_22164,N_22374);
nand U22862 (N_22862,N_22087,N_21434);
xnor U22863 (N_22863,N_22479,N_22463);
and U22864 (N_22864,N_21138,N_21996);
and U22865 (N_22865,N_22026,N_21306);
and U22866 (N_22866,N_22275,N_21607);
nor U22867 (N_22867,N_21790,N_21233);
nand U22868 (N_22868,N_21506,N_21896);
xor U22869 (N_22869,N_21840,N_21900);
nand U22870 (N_22870,N_22024,N_21571);
and U22871 (N_22871,N_21830,N_22455);
or U22872 (N_22872,N_21687,N_21274);
xnor U22873 (N_22873,N_21656,N_21184);
and U22874 (N_22874,N_22196,N_21499);
and U22875 (N_22875,N_22095,N_22046);
nand U22876 (N_22876,N_22379,N_21990);
and U22877 (N_22877,N_21358,N_21724);
and U22878 (N_22878,N_21254,N_21675);
and U22879 (N_22879,N_21971,N_21098);
nor U22880 (N_22880,N_22069,N_22293);
nor U22881 (N_22881,N_21326,N_22426);
nor U22882 (N_22882,N_21598,N_22476);
or U22883 (N_22883,N_21540,N_22312);
and U22884 (N_22884,N_22266,N_22195);
or U22885 (N_22885,N_22109,N_21799);
or U22886 (N_22886,N_22417,N_21834);
xor U22887 (N_22887,N_21685,N_22341);
nor U22888 (N_22888,N_22155,N_21198);
or U22889 (N_22889,N_22131,N_21602);
xor U22890 (N_22890,N_21079,N_21148);
nor U22891 (N_22891,N_22445,N_21560);
nor U22892 (N_22892,N_22132,N_21247);
and U22893 (N_22893,N_21192,N_22317);
nor U22894 (N_22894,N_22367,N_21824);
xnor U22895 (N_22895,N_21919,N_21408);
and U22896 (N_22896,N_21073,N_22294);
and U22897 (N_22897,N_21747,N_21282);
nor U22898 (N_22898,N_21860,N_21772);
and U22899 (N_22899,N_22202,N_21054);
xor U22900 (N_22900,N_21941,N_21704);
nand U22901 (N_22901,N_21346,N_22205);
and U22902 (N_22902,N_21639,N_21123);
nand U22903 (N_22903,N_21484,N_21899);
or U22904 (N_22904,N_22227,N_21412);
xor U22905 (N_22905,N_21746,N_21291);
or U22906 (N_22906,N_22286,N_22077);
nand U22907 (N_22907,N_21439,N_22244);
nor U22908 (N_22908,N_21700,N_22252);
and U22909 (N_22909,N_21241,N_21257);
and U22910 (N_22910,N_22469,N_21205);
and U22911 (N_22911,N_21196,N_22384);
xnor U22912 (N_22912,N_21623,N_21998);
or U22913 (N_22913,N_21357,N_21972);
and U22914 (N_22914,N_22011,N_22023);
or U22915 (N_22915,N_21386,N_22251);
xnor U22916 (N_22916,N_21445,N_22338);
nor U22917 (N_22917,N_21235,N_21477);
and U22918 (N_22918,N_21923,N_21251);
and U22919 (N_22919,N_21530,N_22204);
nor U22920 (N_22920,N_22185,N_21992);
nor U22921 (N_22921,N_21329,N_22186);
nor U22922 (N_22922,N_22260,N_22017);
and U22923 (N_22923,N_21355,N_22416);
xnor U22924 (N_22924,N_22181,N_21817);
or U22925 (N_22925,N_22053,N_21088);
xor U22926 (N_22926,N_22229,N_21431);
xor U22927 (N_22927,N_22047,N_21017);
nor U22928 (N_22928,N_21444,N_22357);
nor U22929 (N_22929,N_21946,N_22415);
and U22930 (N_22930,N_21350,N_21652);
xor U22931 (N_22931,N_22333,N_21745);
or U22932 (N_22932,N_22435,N_21680);
and U22933 (N_22933,N_22246,N_22301);
nor U22934 (N_22934,N_22495,N_21016);
nand U22935 (N_22935,N_21677,N_21299);
and U22936 (N_22936,N_22018,N_22036);
nor U22937 (N_22937,N_21239,N_21610);
xnor U22938 (N_22938,N_22118,N_21547);
or U22939 (N_22939,N_21709,N_21068);
and U22940 (N_22940,N_21837,N_21152);
and U22941 (N_22941,N_22129,N_21085);
xnor U22942 (N_22942,N_22403,N_21953);
nand U22943 (N_22943,N_21204,N_22432);
nand U22944 (N_22944,N_21053,N_22392);
nand U22945 (N_22945,N_21244,N_21011);
nor U22946 (N_22946,N_21721,N_22125);
and U22947 (N_22947,N_22153,N_21494);
or U22948 (N_22948,N_21926,N_22300);
and U22949 (N_22949,N_22268,N_21402);
or U22950 (N_22950,N_22219,N_21002);
or U22951 (N_22951,N_22207,N_22158);
nand U22952 (N_22952,N_21906,N_21762);
and U22953 (N_22953,N_21324,N_21149);
or U22954 (N_22954,N_21644,N_21169);
or U22955 (N_22955,N_21580,N_21674);
or U22956 (N_22956,N_21984,N_21267);
or U22957 (N_22957,N_21083,N_21367);
and U22958 (N_22958,N_22233,N_21767);
xnor U22959 (N_22959,N_21197,N_22013);
xor U22960 (N_22960,N_21288,N_21507);
or U22961 (N_22961,N_21564,N_22442);
xor U22962 (N_22962,N_21683,N_22019);
nor U22963 (N_22963,N_21293,N_21056);
and U22964 (N_22964,N_21920,N_22067);
xnor U22965 (N_22965,N_21708,N_21871);
and U22966 (N_22966,N_21751,N_22332);
and U22967 (N_22967,N_22401,N_21084);
nor U22968 (N_22968,N_21487,N_21112);
nor U22969 (N_22969,N_21549,N_21131);
and U22970 (N_22970,N_21423,N_22162);
xnor U22971 (N_22971,N_21095,N_22149);
nand U22972 (N_22972,N_21890,N_21087);
nor U22973 (N_22973,N_21333,N_21631);
and U22974 (N_22974,N_21246,N_22288);
and U22975 (N_22975,N_21436,N_21057);
and U22976 (N_22976,N_21678,N_21177);
xnor U22977 (N_22977,N_22297,N_22086);
xnor U22978 (N_22978,N_21442,N_21562);
nand U22979 (N_22979,N_21912,N_21770);
or U22980 (N_22980,N_21004,N_22383);
nand U22981 (N_22981,N_21573,N_21050);
xnor U22982 (N_22982,N_22083,N_21335);
nand U22983 (N_22983,N_21220,N_22428);
xnor U22984 (N_22984,N_22041,N_22101);
nor U22985 (N_22985,N_22216,N_21782);
nand U22986 (N_22986,N_21284,N_22003);
nand U22987 (N_22987,N_22093,N_22377);
or U22988 (N_22988,N_22188,N_21539);
nand U22989 (N_22989,N_21388,N_21910);
and U22990 (N_22990,N_21810,N_22358);
xnor U22991 (N_22991,N_21236,N_21940);
xor U22992 (N_22992,N_21086,N_21725);
and U22993 (N_22993,N_21156,N_22201);
xnor U22994 (N_22994,N_22001,N_22478);
xor U22995 (N_22995,N_21836,N_22388);
or U22996 (N_22996,N_21430,N_21065);
or U22997 (N_22997,N_21264,N_21997);
or U22998 (N_22998,N_21199,N_21853);
nor U22999 (N_22999,N_21103,N_22336);
or U23000 (N_23000,N_22292,N_22278);
nand U23001 (N_23001,N_22123,N_21682);
nor U23002 (N_23002,N_21145,N_22173);
nor U23003 (N_23003,N_22240,N_21261);
nor U23004 (N_23004,N_22299,N_22088);
nor U23005 (N_23005,N_22285,N_22176);
xnor U23006 (N_23006,N_21043,N_21844);
nor U23007 (N_23007,N_21140,N_21160);
and U23008 (N_23008,N_21905,N_21632);
nor U23009 (N_23009,N_21885,N_21227);
nor U23010 (N_23010,N_21963,N_21189);
or U23011 (N_23011,N_22141,N_21505);
nand U23012 (N_23012,N_21504,N_21240);
or U23013 (N_23013,N_21877,N_21379);
nand U23014 (N_23014,N_22075,N_21195);
nor U23015 (N_23015,N_21989,N_21295);
or U23016 (N_23016,N_21567,N_21349);
or U23017 (N_23017,N_22128,N_21858);
nand U23018 (N_23018,N_21828,N_21393);
nand U23019 (N_23019,N_21102,N_22226);
nor U23020 (N_23020,N_22380,N_22014);
nand U23021 (N_23021,N_21797,N_21302);
nand U23022 (N_23022,N_21702,N_22450);
or U23023 (N_23023,N_21805,N_21771);
xnor U23024 (N_23024,N_21818,N_21961);
xor U23025 (N_23025,N_21272,N_21792);
xnor U23026 (N_23026,N_22198,N_21142);
nand U23027 (N_23027,N_21727,N_21537);
nor U23028 (N_23028,N_22480,N_21921);
nand U23029 (N_23029,N_21701,N_21889);
or U23030 (N_23030,N_22429,N_21144);
nand U23031 (N_23031,N_22085,N_22493);
xor U23032 (N_23032,N_21497,N_21563);
nor U23033 (N_23033,N_22136,N_21672);
nand U23034 (N_23034,N_22477,N_21898);
xnor U23035 (N_23035,N_21689,N_21476);
nor U23036 (N_23036,N_21579,N_22192);
and U23037 (N_23037,N_21577,N_21800);
or U23038 (N_23038,N_21019,N_21590);
nand U23039 (N_23039,N_22269,N_21458);
nand U23040 (N_23040,N_21698,N_21722);
xnor U23041 (N_23041,N_22397,N_21755);
or U23042 (N_23042,N_22328,N_22315);
xnor U23043 (N_23043,N_21058,N_22439);
or U23044 (N_23044,N_22280,N_22096);
xnor U23045 (N_23045,N_22395,N_21331);
nor U23046 (N_23046,N_22178,N_22351);
nand U23047 (N_23047,N_21880,N_21965);
or U23048 (N_23048,N_21791,N_21665);
xor U23049 (N_23049,N_22330,N_21345);
nand U23050 (N_23050,N_21470,N_21360);
nor U23051 (N_23051,N_21217,N_22247);
nand U23052 (N_23052,N_22209,N_21171);
xor U23053 (N_23053,N_21352,N_21509);
and U23054 (N_23054,N_21168,N_22458);
or U23055 (N_23055,N_21481,N_21309);
or U23056 (N_23056,N_22468,N_22007);
nor U23057 (N_23057,N_21033,N_21390);
nor U23058 (N_23058,N_21879,N_21475);
or U23059 (N_23059,N_21691,N_21646);
xor U23060 (N_23060,N_21649,N_21777);
nor U23061 (N_23061,N_21069,N_22334);
nor U23062 (N_23062,N_21807,N_22199);
xnor U23063 (N_23063,N_22484,N_22210);
xor U23064 (N_23064,N_21116,N_21502);
xor U23065 (N_23065,N_22400,N_21023);
and U23066 (N_23066,N_21622,N_21180);
xnor U23067 (N_23067,N_22060,N_21468);
xor U23068 (N_23068,N_21363,N_21756);
or U23069 (N_23069,N_21316,N_21719);
nand U23070 (N_23070,N_21376,N_22284);
and U23071 (N_23071,N_21482,N_21843);
nor U23072 (N_23072,N_21030,N_22408);
nand U23073 (N_23073,N_21581,N_21541);
nor U23074 (N_23074,N_22471,N_21693);
xnor U23075 (N_23075,N_21951,N_21863);
nor U23076 (N_23076,N_22091,N_22004);
or U23077 (N_23077,N_22344,N_21856);
nor U23078 (N_23078,N_21301,N_21793);
or U23079 (N_23079,N_21059,N_21729);
xor U23080 (N_23080,N_22345,N_21175);
or U23081 (N_23081,N_22316,N_21490);
or U23082 (N_23082,N_21887,N_21121);
and U23083 (N_23083,N_21269,N_21122);
xor U23084 (N_23084,N_22159,N_21977);
nor U23085 (N_23085,N_22139,N_21035);
nand U23086 (N_23086,N_22115,N_21107);
nand U23087 (N_23087,N_22081,N_21255);
and U23088 (N_23088,N_21937,N_21009);
nor U23089 (N_23089,N_22100,N_22308);
and U23090 (N_23090,N_22448,N_22287);
xnor U23091 (N_23091,N_22473,N_22112);
nand U23092 (N_23092,N_21939,N_22276);
or U23093 (N_23093,N_21556,N_22105);
nand U23094 (N_23094,N_21627,N_21850);
and U23095 (N_23095,N_21389,N_21648);
xor U23096 (N_23096,N_21884,N_22499);
nor U23097 (N_23097,N_21096,N_21987);
nand U23098 (N_23098,N_21133,N_21248);
and U23099 (N_23099,N_21588,N_21231);
nor U23100 (N_23100,N_22291,N_21789);
xnor U23101 (N_23101,N_21480,N_21950);
and U23102 (N_23102,N_21024,N_21699);
or U23103 (N_23103,N_22355,N_22166);
nor U23104 (N_23104,N_21740,N_22411);
or U23105 (N_23105,N_22385,N_21105);
and U23106 (N_23106,N_21781,N_22496);
xor U23107 (N_23107,N_21285,N_21875);
xnor U23108 (N_23108,N_21929,N_21219);
xor U23109 (N_23109,N_21532,N_21343);
nand U23110 (N_23110,N_21424,N_21026);
nor U23111 (N_23111,N_22054,N_21473);
and U23112 (N_23112,N_22150,N_21892);
nor U23113 (N_23113,N_22027,N_21773);
and U23114 (N_23114,N_21405,N_21446);
nand U23115 (N_23115,N_22078,N_21332);
and U23116 (N_23116,N_21036,N_22474);
nor U23117 (N_23117,N_21938,N_22325);
xor U23118 (N_23118,N_21586,N_22457);
and U23119 (N_23119,N_21651,N_21039);
and U23120 (N_23120,N_21297,N_21943);
and U23121 (N_23121,N_21118,N_21001);
nand U23122 (N_23122,N_21515,N_21450);
xnor U23123 (N_23123,N_21063,N_21451);
nand U23124 (N_23124,N_21766,N_21348);
nor U23125 (N_23125,N_21207,N_21615);
xnor U23126 (N_23126,N_21829,N_21835);
nor U23127 (N_23127,N_21072,N_21845);
nor U23128 (N_23128,N_21600,N_21891);
or U23129 (N_23129,N_22460,N_22048);
nand U23130 (N_23130,N_22102,N_21094);
and U23131 (N_23131,N_21372,N_21645);
or U23132 (N_23132,N_21528,N_21300);
or U23133 (N_23133,N_21692,N_22262);
xor U23134 (N_23134,N_21313,N_22148);
or U23135 (N_23135,N_22494,N_21527);
nand U23136 (N_23136,N_22371,N_21226);
and U23137 (N_23137,N_21993,N_22080);
or U23138 (N_23138,N_21111,N_21838);
and U23139 (N_23139,N_22373,N_22137);
and U23140 (N_23140,N_21893,N_21340);
nand U23141 (N_23141,N_22487,N_21636);
and U23142 (N_23142,N_22127,N_21483);
and U23143 (N_23143,N_22318,N_22391);
or U23144 (N_23144,N_21763,N_21956);
and U23145 (N_23145,N_22456,N_21585);
or U23146 (N_23146,N_22249,N_21569);
and U23147 (N_23147,N_21418,N_22324);
nor U23148 (N_23148,N_21289,N_21711);
nor U23149 (N_23149,N_22250,N_21201);
nand U23150 (N_23150,N_21870,N_21895);
and U23151 (N_23151,N_21876,N_22073);
nor U23152 (N_23152,N_21407,N_22372);
or U23153 (N_23153,N_21279,N_21127);
nor U23154 (N_23154,N_21064,N_22348);
xor U23155 (N_23155,N_22420,N_21613);
nor U23156 (N_23156,N_21228,N_21566);
and U23157 (N_23157,N_21881,N_21278);
or U23158 (N_23158,N_22295,N_22481);
nand U23159 (N_23159,N_21403,N_22470);
nor U23160 (N_23160,N_21090,N_21522);
nand U23161 (N_23161,N_21392,N_21164);
and U23162 (N_23162,N_22040,N_21055);
and U23163 (N_23163,N_22029,N_21798);
nand U23164 (N_23164,N_21108,N_21730);
nand U23165 (N_23165,N_22034,N_21283);
and U23166 (N_23166,N_21868,N_21981);
nor U23167 (N_23167,N_22283,N_22074);
xnor U23168 (N_23168,N_21130,N_21465);
nand U23169 (N_23169,N_21888,N_21328);
and U23170 (N_23170,N_22361,N_22438);
and U23171 (N_23171,N_21778,N_21882);
xor U23172 (N_23172,N_22212,N_21178);
xnor U23173 (N_23173,N_21878,N_21106);
nand U23174 (N_23174,N_21493,N_22376);
and U23175 (N_23175,N_21866,N_22310);
xor U23176 (N_23176,N_22272,N_22068);
xnor U23177 (N_23177,N_21186,N_21697);
nor U23178 (N_23178,N_21883,N_22321);
or U23179 (N_23179,N_22167,N_21503);
xnor U23180 (N_23180,N_22052,N_22059);
or U23181 (N_23181,N_21399,N_21375);
nand U23182 (N_23182,N_21089,N_21114);
nor U23183 (N_23183,N_21604,N_21753);
nand U23184 (N_23184,N_21342,N_21222);
nor U23185 (N_23185,N_21321,N_21635);
nor U23186 (N_23186,N_21181,N_21533);
xnor U23187 (N_23187,N_21135,N_22174);
nor U23188 (N_23188,N_21741,N_21460);
nor U23189 (N_23189,N_21419,N_21574);
or U23190 (N_23190,N_22062,N_21529);
xnor U23191 (N_23191,N_21958,N_21942);
xor U23192 (N_23192,N_21826,N_21523);
xnor U23193 (N_23193,N_22472,N_21667);
nor U23194 (N_23194,N_21359,N_21092);
or U23195 (N_23195,N_21967,N_21032);
and U23196 (N_23196,N_21172,N_22446);
nor U23197 (N_23197,N_21253,N_22010);
and U23198 (N_23198,N_22191,N_21404);
xnor U23199 (N_23199,N_22169,N_21769);
or U23200 (N_23200,N_21238,N_21139);
xnor U23201 (N_23201,N_22120,N_21421);
and U23202 (N_23202,N_22135,N_21020);
nor U23203 (N_23203,N_21734,N_21099);
and U23204 (N_23204,N_22453,N_21382);
xor U23205 (N_23205,N_21501,N_21903);
nor U23206 (N_23206,N_21538,N_21230);
or U23207 (N_23207,N_22461,N_21457);
or U23208 (N_23208,N_21779,N_21213);
or U23209 (N_23209,N_21918,N_22482);
or U23210 (N_23210,N_21548,N_21314);
nor U23211 (N_23211,N_21361,N_22097);
nand U23212 (N_23212,N_21599,N_21660);
and U23213 (N_23213,N_22222,N_21167);
xnor U23214 (N_23214,N_22006,N_22255);
xor U23215 (N_23215,N_22055,N_22020);
and U23216 (N_23216,N_21954,N_21508);
nor U23217 (N_23217,N_22466,N_21510);
nand U23218 (N_23218,N_21370,N_21338);
or U23219 (N_23219,N_22331,N_21377);
nor U23220 (N_23220,N_21258,N_22444);
nor U23221 (N_23221,N_21034,N_21290);
and U23222 (N_23222,N_22313,N_22221);
nand U23223 (N_23223,N_21754,N_21737);
and U23224 (N_23224,N_21612,N_21406);
nor U23225 (N_23225,N_22157,N_22452);
and U23226 (N_23226,N_21973,N_22079);
nor U23227 (N_23227,N_21519,N_22259);
or U23228 (N_23228,N_21146,N_21662);
or U23229 (N_23229,N_21115,N_21120);
nand U23230 (N_23230,N_22187,N_22171);
or U23231 (N_23231,N_22378,N_21543);
nand U23232 (N_23232,N_22050,N_21684);
nand U23233 (N_23233,N_21119,N_21395);
or U23234 (N_23234,N_21462,N_22160);
and U23235 (N_23235,N_21795,N_21931);
nand U23236 (N_23236,N_21500,N_21544);
and U23237 (N_23237,N_21690,N_22263);
xor U23238 (N_23238,N_22337,N_21867);
or U23239 (N_23239,N_21655,N_21287);
or U23240 (N_23240,N_21603,N_22012);
and U23241 (N_23241,N_21188,N_22256);
xnor U23242 (N_23242,N_21694,N_22151);
nand U23243 (N_23243,N_22042,N_22072);
nor U23244 (N_23244,N_21733,N_21536);
or U23245 (N_23245,N_21969,N_21915);
and U23246 (N_23246,N_21647,N_22133);
nand U23247 (N_23247,N_22225,N_21113);
nand U23248 (N_23248,N_21081,N_21414);
and U23249 (N_23249,N_22193,N_21757);
nand U23250 (N_23250,N_21040,N_21270);
nand U23251 (N_23251,N_21240,N_21395);
nand U23252 (N_23252,N_21484,N_21493);
and U23253 (N_23253,N_22144,N_22455);
xnor U23254 (N_23254,N_22349,N_22465);
or U23255 (N_23255,N_21211,N_21029);
nor U23256 (N_23256,N_21731,N_21657);
or U23257 (N_23257,N_21307,N_21885);
xor U23258 (N_23258,N_22189,N_21534);
xnor U23259 (N_23259,N_21870,N_22416);
or U23260 (N_23260,N_21072,N_21029);
nor U23261 (N_23261,N_21469,N_22195);
and U23262 (N_23262,N_22134,N_22322);
xnor U23263 (N_23263,N_21275,N_22496);
or U23264 (N_23264,N_22041,N_21105);
and U23265 (N_23265,N_21783,N_21466);
xor U23266 (N_23266,N_21183,N_22038);
nor U23267 (N_23267,N_21496,N_21942);
or U23268 (N_23268,N_22382,N_21365);
and U23269 (N_23269,N_22244,N_22336);
and U23270 (N_23270,N_22085,N_22428);
and U23271 (N_23271,N_22240,N_22305);
nor U23272 (N_23272,N_21849,N_21961);
and U23273 (N_23273,N_22076,N_21030);
nor U23274 (N_23274,N_21229,N_21380);
xor U23275 (N_23275,N_22281,N_21243);
xor U23276 (N_23276,N_21347,N_21703);
or U23277 (N_23277,N_22036,N_22298);
nand U23278 (N_23278,N_21768,N_21272);
or U23279 (N_23279,N_22112,N_22433);
and U23280 (N_23280,N_21768,N_21444);
or U23281 (N_23281,N_21893,N_21587);
nor U23282 (N_23282,N_21732,N_21002);
xnor U23283 (N_23283,N_22034,N_22018);
nand U23284 (N_23284,N_21146,N_22221);
nand U23285 (N_23285,N_21539,N_21209);
or U23286 (N_23286,N_22110,N_21477);
xnor U23287 (N_23287,N_22243,N_22018);
and U23288 (N_23288,N_21007,N_21381);
nor U23289 (N_23289,N_22418,N_21641);
nand U23290 (N_23290,N_22378,N_21103);
nor U23291 (N_23291,N_22027,N_22048);
or U23292 (N_23292,N_21902,N_22238);
nor U23293 (N_23293,N_21612,N_21038);
nand U23294 (N_23294,N_21081,N_21483);
and U23295 (N_23295,N_21494,N_21204);
nand U23296 (N_23296,N_21122,N_22485);
and U23297 (N_23297,N_21104,N_21057);
nand U23298 (N_23298,N_21519,N_21718);
xnor U23299 (N_23299,N_21202,N_22435);
xor U23300 (N_23300,N_22314,N_21879);
nor U23301 (N_23301,N_21046,N_21507);
nand U23302 (N_23302,N_22246,N_21341);
or U23303 (N_23303,N_22480,N_21061);
or U23304 (N_23304,N_21059,N_21164);
xnor U23305 (N_23305,N_21641,N_21579);
nor U23306 (N_23306,N_21522,N_21886);
and U23307 (N_23307,N_21993,N_21898);
xor U23308 (N_23308,N_21472,N_21309);
nor U23309 (N_23309,N_22302,N_21157);
and U23310 (N_23310,N_22063,N_21554);
or U23311 (N_23311,N_21149,N_21045);
nand U23312 (N_23312,N_21833,N_21615);
nand U23313 (N_23313,N_22412,N_22400);
nand U23314 (N_23314,N_21066,N_21354);
xnor U23315 (N_23315,N_21304,N_22271);
nor U23316 (N_23316,N_22324,N_21946);
nand U23317 (N_23317,N_21572,N_22427);
nand U23318 (N_23318,N_22087,N_22361);
or U23319 (N_23319,N_22320,N_21034);
nand U23320 (N_23320,N_22150,N_22173);
and U23321 (N_23321,N_21967,N_21045);
or U23322 (N_23322,N_21905,N_21138);
nand U23323 (N_23323,N_22288,N_21276);
and U23324 (N_23324,N_22172,N_21042);
and U23325 (N_23325,N_21579,N_21508);
xnor U23326 (N_23326,N_21185,N_22444);
xor U23327 (N_23327,N_21475,N_22025);
xor U23328 (N_23328,N_21607,N_21528);
nor U23329 (N_23329,N_22080,N_22356);
nand U23330 (N_23330,N_21841,N_21790);
xnor U23331 (N_23331,N_22349,N_21311);
xnor U23332 (N_23332,N_21894,N_21521);
or U23333 (N_23333,N_22410,N_21309);
nand U23334 (N_23334,N_22386,N_22150);
nor U23335 (N_23335,N_22235,N_21321);
nand U23336 (N_23336,N_21195,N_21106);
xor U23337 (N_23337,N_22401,N_22154);
nor U23338 (N_23338,N_21239,N_22017);
nor U23339 (N_23339,N_21105,N_22194);
xor U23340 (N_23340,N_21315,N_21780);
or U23341 (N_23341,N_21630,N_21997);
xor U23342 (N_23342,N_21940,N_22425);
or U23343 (N_23343,N_22461,N_21574);
or U23344 (N_23344,N_21690,N_21556);
xnor U23345 (N_23345,N_21987,N_22281);
and U23346 (N_23346,N_22043,N_21882);
xor U23347 (N_23347,N_22488,N_22018);
and U23348 (N_23348,N_22385,N_22468);
and U23349 (N_23349,N_22227,N_21044);
nand U23350 (N_23350,N_22035,N_21632);
and U23351 (N_23351,N_21018,N_21991);
and U23352 (N_23352,N_22467,N_21116);
or U23353 (N_23353,N_22062,N_21434);
nor U23354 (N_23354,N_21077,N_21321);
or U23355 (N_23355,N_21531,N_21985);
nand U23356 (N_23356,N_22001,N_21826);
xor U23357 (N_23357,N_22490,N_21706);
nand U23358 (N_23358,N_21733,N_22000);
or U23359 (N_23359,N_22160,N_21701);
nand U23360 (N_23360,N_21986,N_21065);
nor U23361 (N_23361,N_21985,N_21300);
or U23362 (N_23362,N_21463,N_21692);
nor U23363 (N_23363,N_22388,N_21453);
nor U23364 (N_23364,N_21314,N_21475);
xor U23365 (N_23365,N_22444,N_21953);
and U23366 (N_23366,N_21249,N_21278);
nand U23367 (N_23367,N_21358,N_21528);
and U23368 (N_23368,N_22022,N_21841);
xor U23369 (N_23369,N_22221,N_21997);
nand U23370 (N_23370,N_21751,N_21318);
nand U23371 (N_23371,N_22158,N_21632);
xnor U23372 (N_23372,N_22343,N_22230);
nand U23373 (N_23373,N_21717,N_22250);
nand U23374 (N_23374,N_22385,N_22384);
nand U23375 (N_23375,N_21739,N_21052);
or U23376 (N_23376,N_21397,N_21279);
and U23377 (N_23377,N_22087,N_21130);
or U23378 (N_23378,N_22370,N_21218);
nor U23379 (N_23379,N_21707,N_21206);
nor U23380 (N_23380,N_21410,N_21511);
nand U23381 (N_23381,N_21743,N_21227);
xnor U23382 (N_23382,N_22303,N_21723);
xnor U23383 (N_23383,N_21122,N_22125);
nor U23384 (N_23384,N_21013,N_21143);
nand U23385 (N_23385,N_22082,N_21670);
xnor U23386 (N_23386,N_21769,N_21980);
nor U23387 (N_23387,N_21619,N_22138);
nor U23388 (N_23388,N_21685,N_21501);
nand U23389 (N_23389,N_22279,N_21034);
xor U23390 (N_23390,N_22188,N_21670);
xnor U23391 (N_23391,N_21864,N_21763);
or U23392 (N_23392,N_21863,N_21269);
nand U23393 (N_23393,N_21880,N_21998);
nor U23394 (N_23394,N_21555,N_21287);
xor U23395 (N_23395,N_22156,N_21476);
nand U23396 (N_23396,N_21816,N_21199);
nor U23397 (N_23397,N_21107,N_21932);
nor U23398 (N_23398,N_21108,N_21408);
or U23399 (N_23399,N_21399,N_22362);
xnor U23400 (N_23400,N_21036,N_21246);
xor U23401 (N_23401,N_22211,N_21414);
xnor U23402 (N_23402,N_22462,N_21788);
nor U23403 (N_23403,N_21628,N_21558);
nand U23404 (N_23404,N_21707,N_21660);
nor U23405 (N_23405,N_22131,N_21860);
nor U23406 (N_23406,N_21070,N_22237);
nor U23407 (N_23407,N_21647,N_22000);
and U23408 (N_23408,N_21092,N_21669);
nor U23409 (N_23409,N_21227,N_21613);
xnor U23410 (N_23410,N_21294,N_21157);
and U23411 (N_23411,N_21346,N_21937);
xor U23412 (N_23412,N_21454,N_21351);
nor U23413 (N_23413,N_22489,N_21450);
xnor U23414 (N_23414,N_21163,N_21113);
xor U23415 (N_23415,N_21630,N_21096);
and U23416 (N_23416,N_21323,N_21907);
nor U23417 (N_23417,N_22474,N_22011);
nand U23418 (N_23418,N_21014,N_21806);
and U23419 (N_23419,N_21471,N_21381);
nor U23420 (N_23420,N_21997,N_21624);
and U23421 (N_23421,N_21540,N_21402);
or U23422 (N_23422,N_21477,N_21654);
or U23423 (N_23423,N_22007,N_22016);
or U23424 (N_23424,N_21543,N_21912);
or U23425 (N_23425,N_21466,N_21074);
xor U23426 (N_23426,N_22344,N_21535);
or U23427 (N_23427,N_21880,N_22257);
nand U23428 (N_23428,N_21468,N_21264);
nor U23429 (N_23429,N_21733,N_21715);
or U23430 (N_23430,N_21629,N_21267);
or U23431 (N_23431,N_21336,N_21075);
xor U23432 (N_23432,N_22042,N_21436);
or U23433 (N_23433,N_22030,N_22096);
or U23434 (N_23434,N_21220,N_21285);
nand U23435 (N_23435,N_21355,N_21837);
nor U23436 (N_23436,N_21436,N_21877);
xor U23437 (N_23437,N_21766,N_22491);
or U23438 (N_23438,N_22397,N_21042);
xor U23439 (N_23439,N_21811,N_21090);
and U23440 (N_23440,N_22235,N_21258);
or U23441 (N_23441,N_22331,N_21236);
or U23442 (N_23442,N_21964,N_21750);
and U23443 (N_23443,N_21366,N_21377);
or U23444 (N_23444,N_21400,N_21316);
nand U23445 (N_23445,N_21073,N_22237);
and U23446 (N_23446,N_21236,N_21135);
nor U23447 (N_23447,N_22330,N_22064);
nor U23448 (N_23448,N_22465,N_21512);
nand U23449 (N_23449,N_21872,N_21589);
nor U23450 (N_23450,N_21186,N_22044);
nand U23451 (N_23451,N_21673,N_21496);
nand U23452 (N_23452,N_21506,N_22200);
nor U23453 (N_23453,N_21031,N_21183);
and U23454 (N_23454,N_22004,N_21545);
nor U23455 (N_23455,N_21975,N_22138);
nand U23456 (N_23456,N_21602,N_21698);
or U23457 (N_23457,N_21757,N_21244);
xor U23458 (N_23458,N_21534,N_21864);
nor U23459 (N_23459,N_21718,N_21724);
xnor U23460 (N_23460,N_22117,N_21748);
nand U23461 (N_23461,N_21391,N_22409);
or U23462 (N_23462,N_21127,N_21851);
xnor U23463 (N_23463,N_22359,N_22426);
nor U23464 (N_23464,N_21346,N_22293);
xnor U23465 (N_23465,N_21839,N_21431);
nor U23466 (N_23466,N_22049,N_22145);
nor U23467 (N_23467,N_21910,N_22048);
xnor U23468 (N_23468,N_21594,N_22328);
nor U23469 (N_23469,N_21522,N_21195);
nand U23470 (N_23470,N_22333,N_21255);
and U23471 (N_23471,N_21118,N_21627);
or U23472 (N_23472,N_22003,N_21566);
nand U23473 (N_23473,N_21815,N_21417);
or U23474 (N_23474,N_22296,N_21598);
nor U23475 (N_23475,N_22089,N_21802);
xnor U23476 (N_23476,N_22131,N_22027);
nand U23477 (N_23477,N_21129,N_21948);
and U23478 (N_23478,N_21216,N_21573);
or U23479 (N_23479,N_22046,N_21039);
and U23480 (N_23480,N_22008,N_21612);
or U23481 (N_23481,N_21908,N_21550);
nand U23482 (N_23482,N_22230,N_21319);
xor U23483 (N_23483,N_21073,N_21053);
xnor U23484 (N_23484,N_21121,N_22297);
nor U23485 (N_23485,N_21105,N_21656);
nor U23486 (N_23486,N_21837,N_21448);
or U23487 (N_23487,N_21790,N_21186);
nor U23488 (N_23488,N_21687,N_22450);
nor U23489 (N_23489,N_21595,N_21531);
nand U23490 (N_23490,N_21102,N_21087);
and U23491 (N_23491,N_22425,N_22046);
or U23492 (N_23492,N_21809,N_21924);
or U23493 (N_23493,N_22133,N_21173);
and U23494 (N_23494,N_21069,N_22110);
and U23495 (N_23495,N_22161,N_21924);
and U23496 (N_23496,N_22243,N_21513);
and U23497 (N_23497,N_21541,N_22046);
nand U23498 (N_23498,N_21838,N_21986);
or U23499 (N_23499,N_21153,N_21899);
and U23500 (N_23500,N_21203,N_21326);
xnor U23501 (N_23501,N_21420,N_21221);
nand U23502 (N_23502,N_21411,N_21907);
nand U23503 (N_23503,N_22427,N_22320);
xnor U23504 (N_23504,N_22038,N_22348);
xor U23505 (N_23505,N_22213,N_21666);
xnor U23506 (N_23506,N_21832,N_22364);
or U23507 (N_23507,N_21884,N_22410);
or U23508 (N_23508,N_22279,N_22361);
nand U23509 (N_23509,N_21728,N_22427);
nand U23510 (N_23510,N_22415,N_21576);
xor U23511 (N_23511,N_21235,N_22344);
or U23512 (N_23512,N_21818,N_21556);
nand U23513 (N_23513,N_21988,N_21269);
nor U23514 (N_23514,N_22133,N_22493);
xor U23515 (N_23515,N_21113,N_21839);
nand U23516 (N_23516,N_22170,N_22214);
nor U23517 (N_23517,N_21615,N_21093);
and U23518 (N_23518,N_21671,N_21988);
nand U23519 (N_23519,N_21410,N_22179);
xor U23520 (N_23520,N_21248,N_22154);
nand U23521 (N_23521,N_21428,N_22007);
nand U23522 (N_23522,N_22211,N_21505);
and U23523 (N_23523,N_21251,N_22097);
and U23524 (N_23524,N_21665,N_22108);
nand U23525 (N_23525,N_22112,N_22368);
nor U23526 (N_23526,N_21991,N_21460);
xor U23527 (N_23527,N_21733,N_21356);
nand U23528 (N_23528,N_21766,N_22428);
xor U23529 (N_23529,N_21568,N_22245);
nor U23530 (N_23530,N_21802,N_22391);
nor U23531 (N_23531,N_21747,N_22094);
nor U23532 (N_23532,N_21799,N_21198);
or U23533 (N_23533,N_21853,N_22222);
xor U23534 (N_23534,N_22128,N_21538);
or U23535 (N_23535,N_21902,N_21570);
nor U23536 (N_23536,N_21358,N_21367);
nor U23537 (N_23537,N_21683,N_21270);
xnor U23538 (N_23538,N_21088,N_21003);
nand U23539 (N_23539,N_22103,N_21281);
and U23540 (N_23540,N_21894,N_21517);
or U23541 (N_23541,N_21150,N_21850);
or U23542 (N_23542,N_21185,N_21971);
xor U23543 (N_23543,N_21566,N_21710);
or U23544 (N_23544,N_21647,N_21499);
xnor U23545 (N_23545,N_21809,N_21050);
or U23546 (N_23546,N_21233,N_21641);
or U23547 (N_23547,N_21894,N_22170);
nand U23548 (N_23548,N_22305,N_21578);
xor U23549 (N_23549,N_21068,N_22494);
or U23550 (N_23550,N_21924,N_22472);
nand U23551 (N_23551,N_21425,N_21342);
or U23552 (N_23552,N_21500,N_21704);
nand U23553 (N_23553,N_21822,N_21755);
or U23554 (N_23554,N_22221,N_21999);
nand U23555 (N_23555,N_21022,N_22381);
or U23556 (N_23556,N_21157,N_21054);
nor U23557 (N_23557,N_22394,N_22193);
nor U23558 (N_23558,N_22285,N_22164);
nand U23559 (N_23559,N_21769,N_21880);
nor U23560 (N_23560,N_21749,N_21503);
or U23561 (N_23561,N_22293,N_21629);
or U23562 (N_23562,N_21875,N_22019);
and U23563 (N_23563,N_21103,N_22048);
or U23564 (N_23564,N_21944,N_22020);
nand U23565 (N_23565,N_21319,N_21587);
nand U23566 (N_23566,N_21281,N_21185);
xor U23567 (N_23567,N_22319,N_21202);
xnor U23568 (N_23568,N_21899,N_21546);
xnor U23569 (N_23569,N_21824,N_21207);
nor U23570 (N_23570,N_21642,N_21043);
nor U23571 (N_23571,N_21595,N_21382);
and U23572 (N_23572,N_21681,N_21881);
nor U23573 (N_23573,N_21532,N_22062);
or U23574 (N_23574,N_21242,N_21865);
xnor U23575 (N_23575,N_22436,N_22467);
nand U23576 (N_23576,N_22035,N_21498);
nor U23577 (N_23577,N_22411,N_21388);
and U23578 (N_23578,N_21528,N_21753);
and U23579 (N_23579,N_21681,N_21445);
xor U23580 (N_23580,N_21093,N_21225);
or U23581 (N_23581,N_21761,N_22016);
nand U23582 (N_23582,N_21069,N_21536);
or U23583 (N_23583,N_22298,N_21017);
nand U23584 (N_23584,N_21343,N_21692);
nand U23585 (N_23585,N_21838,N_22021);
or U23586 (N_23586,N_21605,N_22207);
or U23587 (N_23587,N_21459,N_21561);
and U23588 (N_23588,N_21575,N_21853);
nor U23589 (N_23589,N_21774,N_22234);
nand U23590 (N_23590,N_21381,N_21445);
nor U23591 (N_23591,N_21886,N_21492);
and U23592 (N_23592,N_21593,N_21863);
nand U23593 (N_23593,N_22163,N_21298);
and U23594 (N_23594,N_21535,N_22392);
nor U23595 (N_23595,N_22159,N_22098);
nand U23596 (N_23596,N_22298,N_21510);
nand U23597 (N_23597,N_22174,N_21805);
nand U23598 (N_23598,N_22218,N_21703);
or U23599 (N_23599,N_22302,N_21834);
nand U23600 (N_23600,N_21694,N_21828);
or U23601 (N_23601,N_21580,N_21513);
nor U23602 (N_23602,N_22099,N_21387);
nor U23603 (N_23603,N_21495,N_22043);
nand U23604 (N_23604,N_21928,N_21748);
xnor U23605 (N_23605,N_21578,N_21696);
xnor U23606 (N_23606,N_21443,N_22069);
nor U23607 (N_23607,N_21672,N_22309);
or U23608 (N_23608,N_22339,N_22474);
xor U23609 (N_23609,N_22480,N_21747);
nor U23610 (N_23610,N_22026,N_22185);
and U23611 (N_23611,N_22177,N_21350);
and U23612 (N_23612,N_21306,N_21143);
or U23613 (N_23613,N_21094,N_22452);
nand U23614 (N_23614,N_22068,N_21423);
xor U23615 (N_23615,N_22153,N_21705);
xnor U23616 (N_23616,N_22232,N_21620);
nor U23617 (N_23617,N_21262,N_22182);
nand U23618 (N_23618,N_21211,N_22445);
nor U23619 (N_23619,N_21469,N_22388);
xor U23620 (N_23620,N_21661,N_21142);
xnor U23621 (N_23621,N_21998,N_21323);
nand U23622 (N_23622,N_21796,N_21795);
and U23623 (N_23623,N_21929,N_22382);
nor U23624 (N_23624,N_21529,N_21094);
xnor U23625 (N_23625,N_22003,N_22284);
xor U23626 (N_23626,N_22381,N_21286);
nand U23627 (N_23627,N_21757,N_22123);
xor U23628 (N_23628,N_22446,N_21489);
nor U23629 (N_23629,N_21305,N_21130);
nor U23630 (N_23630,N_21143,N_21759);
nand U23631 (N_23631,N_21814,N_22405);
or U23632 (N_23632,N_21777,N_22452);
nor U23633 (N_23633,N_21306,N_21976);
nand U23634 (N_23634,N_22297,N_21170);
nor U23635 (N_23635,N_21386,N_21897);
xor U23636 (N_23636,N_21515,N_22396);
nand U23637 (N_23637,N_22048,N_21168);
xor U23638 (N_23638,N_22416,N_21126);
nand U23639 (N_23639,N_21004,N_22153);
nor U23640 (N_23640,N_22118,N_21974);
and U23641 (N_23641,N_21345,N_21937);
or U23642 (N_23642,N_22327,N_22383);
xnor U23643 (N_23643,N_21752,N_21262);
nand U23644 (N_23644,N_21553,N_21926);
and U23645 (N_23645,N_21450,N_21042);
or U23646 (N_23646,N_22004,N_21199);
and U23647 (N_23647,N_22093,N_22073);
and U23648 (N_23648,N_22421,N_22014);
or U23649 (N_23649,N_22369,N_21082);
nor U23650 (N_23650,N_21806,N_21350);
nand U23651 (N_23651,N_21982,N_21101);
nand U23652 (N_23652,N_22318,N_22207);
or U23653 (N_23653,N_22452,N_22071);
xnor U23654 (N_23654,N_21374,N_21837);
and U23655 (N_23655,N_22246,N_21318);
nor U23656 (N_23656,N_21176,N_21786);
and U23657 (N_23657,N_21406,N_21506);
or U23658 (N_23658,N_21021,N_21607);
and U23659 (N_23659,N_21019,N_21612);
nor U23660 (N_23660,N_21993,N_21195);
nand U23661 (N_23661,N_22050,N_21767);
nor U23662 (N_23662,N_21029,N_22149);
or U23663 (N_23663,N_21646,N_21628);
nand U23664 (N_23664,N_22408,N_22320);
nor U23665 (N_23665,N_21898,N_22003);
nand U23666 (N_23666,N_22342,N_21668);
nor U23667 (N_23667,N_22061,N_21347);
nor U23668 (N_23668,N_22356,N_21483);
nand U23669 (N_23669,N_22066,N_22465);
or U23670 (N_23670,N_22464,N_21637);
nand U23671 (N_23671,N_21297,N_22469);
or U23672 (N_23672,N_21687,N_22247);
or U23673 (N_23673,N_22121,N_22177);
and U23674 (N_23674,N_21609,N_21091);
xor U23675 (N_23675,N_22049,N_21677);
and U23676 (N_23676,N_21590,N_21094);
nand U23677 (N_23677,N_22029,N_21943);
nor U23678 (N_23678,N_22276,N_21582);
xnor U23679 (N_23679,N_22449,N_21401);
nand U23680 (N_23680,N_21743,N_21408);
or U23681 (N_23681,N_21157,N_22265);
nand U23682 (N_23682,N_21828,N_21961);
nand U23683 (N_23683,N_22247,N_21163);
and U23684 (N_23684,N_21009,N_22230);
and U23685 (N_23685,N_22020,N_22181);
and U23686 (N_23686,N_22044,N_21547);
and U23687 (N_23687,N_22117,N_22445);
or U23688 (N_23688,N_21707,N_21491);
nand U23689 (N_23689,N_22392,N_21643);
nor U23690 (N_23690,N_21520,N_21186);
xor U23691 (N_23691,N_22308,N_22201);
nor U23692 (N_23692,N_21647,N_21769);
nand U23693 (N_23693,N_22276,N_21197);
nor U23694 (N_23694,N_21988,N_21207);
and U23695 (N_23695,N_21009,N_22163);
nand U23696 (N_23696,N_21800,N_21121);
nand U23697 (N_23697,N_21485,N_21916);
nand U23698 (N_23698,N_21871,N_22205);
nor U23699 (N_23699,N_22383,N_21574);
xor U23700 (N_23700,N_21040,N_22331);
and U23701 (N_23701,N_21842,N_21664);
nor U23702 (N_23702,N_22383,N_21964);
nand U23703 (N_23703,N_22119,N_21129);
and U23704 (N_23704,N_21643,N_21807);
nand U23705 (N_23705,N_21546,N_22251);
nor U23706 (N_23706,N_22036,N_21776);
nand U23707 (N_23707,N_21020,N_21076);
nor U23708 (N_23708,N_21488,N_22438);
nor U23709 (N_23709,N_21413,N_21503);
nand U23710 (N_23710,N_21932,N_21047);
or U23711 (N_23711,N_21916,N_21816);
or U23712 (N_23712,N_21295,N_21410);
nor U23713 (N_23713,N_21448,N_21172);
and U23714 (N_23714,N_22395,N_22465);
and U23715 (N_23715,N_21253,N_22279);
nand U23716 (N_23716,N_21715,N_21063);
and U23717 (N_23717,N_22367,N_21085);
nand U23718 (N_23718,N_22300,N_21467);
or U23719 (N_23719,N_22355,N_21184);
xnor U23720 (N_23720,N_21414,N_22042);
xnor U23721 (N_23721,N_21408,N_21274);
nor U23722 (N_23722,N_21480,N_21032);
and U23723 (N_23723,N_21165,N_22220);
nor U23724 (N_23724,N_21145,N_21944);
nand U23725 (N_23725,N_22498,N_21024);
and U23726 (N_23726,N_21222,N_21605);
nand U23727 (N_23727,N_21290,N_22260);
or U23728 (N_23728,N_22231,N_21847);
or U23729 (N_23729,N_21373,N_21901);
nor U23730 (N_23730,N_21469,N_21386);
or U23731 (N_23731,N_22442,N_22493);
xnor U23732 (N_23732,N_22494,N_21726);
and U23733 (N_23733,N_22457,N_21364);
and U23734 (N_23734,N_22360,N_21974);
nor U23735 (N_23735,N_21282,N_22483);
xor U23736 (N_23736,N_22152,N_21814);
nand U23737 (N_23737,N_21729,N_21868);
nand U23738 (N_23738,N_21557,N_22369);
nand U23739 (N_23739,N_21068,N_21381);
nor U23740 (N_23740,N_21857,N_21328);
or U23741 (N_23741,N_21417,N_22018);
or U23742 (N_23742,N_21557,N_21295);
and U23743 (N_23743,N_21426,N_21683);
or U23744 (N_23744,N_22494,N_21165);
or U23745 (N_23745,N_21907,N_21240);
and U23746 (N_23746,N_21363,N_21442);
nor U23747 (N_23747,N_21961,N_21888);
or U23748 (N_23748,N_22374,N_21016);
nor U23749 (N_23749,N_21466,N_21846);
xnor U23750 (N_23750,N_21109,N_21771);
nand U23751 (N_23751,N_21974,N_21548);
and U23752 (N_23752,N_22032,N_21943);
or U23753 (N_23753,N_21590,N_22404);
and U23754 (N_23754,N_21730,N_21467);
or U23755 (N_23755,N_21327,N_22434);
nor U23756 (N_23756,N_22139,N_22439);
xor U23757 (N_23757,N_21937,N_21614);
and U23758 (N_23758,N_21752,N_21969);
nor U23759 (N_23759,N_21248,N_21443);
or U23760 (N_23760,N_22017,N_21351);
nor U23761 (N_23761,N_21803,N_21847);
nor U23762 (N_23762,N_22213,N_21038);
or U23763 (N_23763,N_22404,N_21270);
xnor U23764 (N_23764,N_22034,N_21579);
nor U23765 (N_23765,N_21518,N_21774);
nor U23766 (N_23766,N_21890,N_21582);
xnor U23767 (N_23767,N_21033,N_22020);
or U23768 (N_23768,N_21036,N_21206);
nand U23769 (N_23769,N_21896,N_22328);
xnor U23770 (N_23770,N_21975,N_22000);
nor U23771 (N_23771,N_22363,N_21129);
nor U23772 (N_23772,N_21152,N_21106);
nor U23773 (N_23773,N_21733,N_21811);
xnor U23774 (N_23774,N_22016,N_21117);
nand U23775 (N_23775,N_21586,N_22269);
and U23776 (N_23776,N_21666,N_21801);
nor U23777 (N_23777,N_21576,N_21890);
nand U23778 (N_23778,N_22330,N_22414);
xor U23779 (N_23779,N_22425,N_21792);
nand U23780 (N_23780,N_21283,N_21064);
and U23781 (N_23781,N_22232,N_21186);
nor U23782 (N_23782,N_21162,N_22070);
or U23783 (N_23783,N_22020,N_21079);
xor U23784 (N_23784,N_21444,N_21067);
xor U23785 (N_23785,N_22415,N_21710);
nand U23786 (N_23786,N_21087,N_21757);
nor U23787 (N_23787,N_21214,N_21101);
nor U23788 (N_23788,N_22104,N_21393);
nand U23789 (N_23789,N_21894,N_21021);
and U23790 (N_23790,N_22047,N_21424);
or U23791 (N_23791,N_21813,N_21500);
nor U23792 (N_23792,N_21916,N_21635);
and U23793 (N_23793,N_22027,N_21350);
nand U23794 (N_23794,N_21567,N_22058);
and U23795 (N_23795,N_21946,N_21378);
nand U23796 (N_23796,N_21099,N_21161);
and U23797 (N_23797,N_21906,N_21646);
nor U23798 (N_23798,N_21192,N_21223);
xor U23799 (N_23799,N_22030,N_21327);
nor U23800 (N_23800,N_21723,N_21424);
or U23801 (N_23801,N_21815,N_22105);
nor U23802 (N_23802,N_21707,N_21451);
xor U23803 (N_23803,N_22057,N_21674);
and U23804 (N_23804,N_21969,N_22433);
xor U23805 (N_23805,N_22264,N_21763);
and U23806 (N_23806,N_22484,N_22357);
xnor U23807 (N_23807,N_21569,N_21904);
or U23808 (N_23808,N_21725,N_21716);
and U23809 (N_23809,N_21177,N_21164);
xnor U23810 (N_23810,N_21816,N_21590);
xor U23811 (N_23811,N_21493,N_21910);
nor U23812 (N_23812,N_21735,N_22337);
nand U23813 (N_23813,N_22205,N_21310);
or U23814 (N_23814,N_21695,N_21315);
and U23815 (N_23815,N_21257,N_22111);
xor U23816 (N_23816,N_21540,N_21388);
and U23817 (N_23817,N_22476,N_21757);
and U23818 (N_23818,N_22323,N_22399);
nor U23819 (N_23819,N_21666,N_22163);
and U23820 (N_23820,N_21308,N_21754);
xnor U23821 (N_23821,N_22268,N_22150);
and U23822 (N_23822,N_21826,N_22488);
xnor U23823 (N_23823,N_21202,N_21131);
xor U23824 (N_23824,N_21195,N_21399);
nand U23825 (N_23825,N_22327,N_22098);
nor U23826 (N_23826,N_21881,N_21541);
or U23827 (N_23827,N_21936,N_22313);
xor U23828 (N_23828,N_22150,N_21600);
nand U23829 (N_23829,N_22240,N_22355);
nand U23830 (N_23830,N_22266,N_21438);
xor U23831 (N_23831,N_21771,N_21947);
and U23832 (N_23832,N_21234,N_22125);
and U23833 (N_23833,N_21869,N_22300);
xor U23834 (N_23834,N_22315,N_22305);
and U23835 (N_23835,N_21688,N_21377);
xor U23836 (N_23836,N_21700,N_21532);
nor U23837 (N_23837,N_21469,N_22450);
and U23838 (N_23838,N_21647,N_21434);
or U23839 (N_23839,N_22146,N_21662);
and U23840 (N_23840,N_21098,N_21603);
xor U23841 (N_23841,N_22311,N_21193);
nand U23842 (N_23842,N_21808,N_21909);
nand U23843 (N_23843,N_21553,N_21658);
and U23844 (N_23844,N_21812,N_21925);
nand U23845 (N_23845,N_22463,N_22339);
nor U23846 (N_23846,N_21710,N_22280);
and U23847 (N_23847,N_22245,N_21331);
and U23848 (N_23848,N_21354,N_22207);
nor U23849 (N_23849,N_21974,N_21214);
nand U23850 (N_23850,N_21436,N_22197);
xor U23851 (N_23851,N_22209,N_21406);
nor U23852 (N_23852,N_21818,N_21206);
xor U23853 (N_23853,N_21525,N_21668);
xor U23854 (N_23854,N_21471,N_21629);
nor U23855 (N_23855,N_21726,N_21733);
nor U23856 (N_23856,N_21571,N_21509);
and U23857 (N_23857,N_21618,N_22060);
or U23858 (N_23858,N_21578,N_22454);
nor U23859 (N_23859,N_22444,N_21163);
nand U23860 (N_23860,N_21376,N_22282);
xor U23861 (N_23861,N_21479,N_22407);
xnor U23862 (N_23862,N_21713,N_22176);
and U23863 (N_23863,N_21022,N_21720);
and U23864 (N_23864,N_22221,N_21116);
or U23865 (N_23865,N_22101,N_21290);
nand U23866 (N_23866,N_21207,N_22330);
xnor U23867 (N_23867,N_22118,N_21069);
xnor U23868 (N_23868,N_21477,N_21992);
or U23869 (N_23869,N_21344,N_21372);
or U23870 (N_23870,N_22415,N_22356);
nor U23871 (N_23871,N_21555,N_22264);
xor U23872 (N_23872,N_22227,N_22263);
xnor U23873 (N_23873,N_22117,N_21152);
nor U23874 (N_23874,N_21647,N_22059);
or U23875 (N_23875,N_21113,N_22078);
xor U23876 (N_23876,N_21990,N_21036);
and U23877 (N_23877,N_21805,N_22153);
nor U23878 (N_23878,N_22212,N_21195);
xor U23879 (N_23879,N_22410,N_22071);
xor U23880 (N_23880,N_22105,N_22363);
xnor U23881 (N_23881,N_21913,N_21970);
nor U23882 (N_23882,N_21829,N_21963);
or U23883 (N_23883,N_21580,N_21088);
xnor U23884 (N_23884,N_21207,N_22021);
and U23885 (N_23885,N_21567,N_21800);
nand U23886 (N_23886,N_21067,N_21874);
or U23887 (N_23887,N_22448,N_21884);
xor U23888 (N_23888,N_21471,N_21318);
and U23889 (N_23889,N_21878,N_21483);
and U23890 (N_23890,N_22414,N_21628);
nor U23891 (N_23891,N_21149,N_21054);
and U23892 (N_23892,N_21196,N_21454);
nand U23893 (N_23893,N_21654,N_22070);
or U23894 (N_23894,N_21401,N_21545);
nand U23895 (N_23895,N_21625,N_21379);
xnor U23896 (N_23896,N_21793,N_21085);
nand U23897 (N_23897,N_21950,N_21160);
and U23898 (N_23898,N_21153,N_21493);
nor U23899 (N_23899,N_21603,N_22468);
or U23900 (N_23900,N_21419,N_21679);
nand U23901 (N_23901,N_21250,N_22231);
or U23902 (N_23902,N_21770,N_22081);
or U23903 (N_23903,N_22083,N_22151);
nor U23904 (N_23904,N_21623,N_21650);
xor U23905 (N_23905,N_21232,N_21482);
nor U23906 (N_23906,N_22015,N_22372);
nor U23907 (N_23907,N_22022,N_21584);
or U23908 (N_23908,N_22467,N_22124);
xor U23909 (N_23909,N_22482,N_22468);
and U23910 (N_23910,N_21101,N_21944);
nand U23911 (N_23911,N_21075,N_22115);
or U23912 (N_23912,N_21001,N_22382);
and U23913 (N_23913,N_21949,N_21691);
nand U23914 (N_23914,N_21299,N_21738);
nand U23915 (N_23915,N_21305,N_21056);
or U23916 (N_23916,N_21682,N_21723);
and U23917 (N_23917,N_21387,N_21219);
nor U23918 (N_23918,N_21321,N_21683);
nor U23919 (N_23919,N_22000,N_22443);
or U23920 (N_23920,N_22348,N_21486);
nand U23921 (N_23921,N_22455,N_21431);
and U23922 (N_23922,N_21327,N_21697);
nand U23923 (N_23923,N_21754,N_21388);
nor U23924 (N_23924,N_21828,N_21991);
and U23925 (N_23925,N_22455,N_22268);
and U23926 (N_23926,N_21445,N_22415);
nand U23927 (N_23927,N_22380,N_21487);
and U23928 (N_23928,N_22255,N_21652);
nand U23929 (N_23929,N_21853,N_22470);
and U23930 (N_23930,N_21812,N_22086);
nand U23931 (N_23931,N_21599,N_21240);
or U23932 (N_23932,N_22012,N_21849);
xnor U23933 (N_23933,N_22054,N_21357);
and U23934 (N_23934,N_22034,N_22017);
xor U23935 (N_23935,N_21243,N_21259);
and U23936 (N_23936,N_21708,N_22418);
nand U23937 (N_23937,N_21357,N_21781);
xor U23938 (N_23938,N_21993,N_21733);
nand U23939 (N_23939,N_21929,N_21469);
xor U23940 (N_23940,N_22346,N_21066);
or U23941 (N_23941,N_22154,N_21162);
xor U23942 (N_23942,N_21946,N_21302);
or U23943 (N_23943,N_21810,N_21410);
nor U23944 (N_23944,N_21015,N_21416);
xnor U23945 (N_23945,N_21571,N_21425);
or U23946 (N_23946,N_21885,N_22439);
and U23947 (N_23947,N_21460,N_22170);
nand U23948 (N_23948,N_22065,N_21325);
or U23949 (N_23949,N_21156,N_22424);
or U23950 (N_23950,N_21921,N_21779);
xnor U23951 (N_23951,N_22157,N_22336);
nand U23952 (N_23952,N_21308,N_21334);
and U23953 (N_23953,N_22200,N_21430);
xnor U23954 (N_23954,N_21135,N_21558);
xor U23955 (N_23955,N_21097,N_21950);
nor U23956 (N_23956,N_21989,N_21123);
nor U23957 (N_23957,N_21770,N_21027);
xnor U23958 (N_23958,N_22363,N_21074);
nor U23959 (N_23959,N_22280,N_21463);
or U23960 (N_23960,N_21277,N_21132);
nand U23961 (N_23961,N_21187,N_21919);
or U23962 (N_23962,N_21878,N_22004);
nand U23963 (N_23963,N_21717,N_21761);
and U23964 (N_23964,N_21446,N_21485);
and U23965 (N_23965,N_21665,N_21905);
or U23966 (N_23966,N_21132,N_21003);
nor U23967 (N_23967,N_21443,N_21815);
and U23968 (N_23968,N_21503,N_21399);
or U23969 (N_23969,N_22450,N_21429);
nor U23970 (N_23970,N_21297,N_21651);
nor U23971 (N_23971,N_22376,N_21197);
and U23972 (N_23972,N_22372,N_21180);
nor U23973 (N_23973,N_22477,N_22431);
or U23974 (N_23974,N_22248,N_21984);
nor U23975 (N_23975,N_22432,N_21774);
nand U23976 (N_23976,N_22295,N_21906);
nor U23977 (N_23977,N_22234,N_22496);
xnor U23978 (N_23978,N_22319,N_21472);
xor U23979 (N_23979,N_21018,N_21733);
or U23980 (N_23980,N_22372,N_21007);
or U23981 (N_23981,N_21574,N_22449);
nand U23982 (N_23982,N_21056,N_22252);
and U23983 (N_23983,N_21344,N_22426);
and U23984 (N_23984,N_21369,N_21416);
nor U23985 (N_23985,N_22033,N_21170);
xnor U23986 (N_23986,N_22163,N_21510);
or U23987 (N_23987,N_21504,N_21345);
nand U23988 (N_23988,N_21149,N_22266);
nor U23989 (N_23989,N_21778,N_21595);
nor U23990 (N_23990,N_21210,N_22036);
nor U23991 (N_23991,N_22386,N_21212);
or U23992 (N_23992,N_22139,N_21956);
nor U23993 (N_23993,N_22256,N_21618);
and U23994 (N_23994,N_21702,N_22248);
xnor U23995 (N_23995,N_21893,N_22080);
and U23996 (N_23996,N_21702,N_22113);
or U23997 (N_23997,N_21328,N_21807);
and U23998 (N_23998,N_21844,N_22403);
xnor U23999 (N_23999,N_21039,N_21262);
xor U24000 (N_24000,N_23852,N_22940);
nor U24001 (N_24001,N_23396,N_23600);
xor U24002 (N_24002,N_23978,N_23029);
nor U24003 (N_24003,N_23089,N_22644);
nand U24004 (N_24004,N_23502,N_23905);
nor U24005 (N_24005,N_23283,N_23373);
and U24006 (N_24006,N_23950,N_22942);
nand U24007 (N_24007,N_22690,N_23639);
nor U24008 (N_24008,N_22965,N_23590);
xor U24009 (N_24009,N_22646,N_23793);
nor U24010 (N_24010,N_23969,N_23770);
and U24011 (N_24011,N_23232,N_23967);
and U24012 (N_24012,N_23321,N_22887);
xnor U24013 (N_24013,N_23399,N_22811);
and U24014 (N_24014,N_23709,N_23182);
or U24015 (N_24015,N_22615,N_23382);
nor U24016 (N_24016,N_23522,N_22805);
nand U24017 (N_24017,N_23983,N_23724);
or U24018 (N_24018,N_22713,N_23612);
and U24019 (N_24019,N_22996,N_23159);
nand U24020 (N_24020,N_22674,N_23879);
nor U24021 (N_24021,N_23298,N_23333);
nor U24022 (N_24022,N_23164,N_23789);
nor U24023 (N_24023,N_22832,N_23765);
or U24024 (N_24024,N_22914,N_22726);
and U24025 (N_24025,N_22896,N_22558);
nor U24026 (N_24026,N_23657,N_23360);
and U24027 (N_24027,N_23307,N_22560);
and U24028 (N_24028,N_23908,N_23822);
nor U24029 (N_24029,N_23990,N_22852);
nor U24030 (N_24030,N_22592,N_23666);
xor U24031 (N_24031,N_23994,N_23486);
and U24032 (N_24032,N_23376,N_23514);
or U24033 (N_24033,N_23845,N_23915);
xor U24034 (N_24034,N_23052,N_23183);
or U24035 (N_24035,N_23788,N_23912);
xor U24036 (N_24036,N_22841,N_23741);
and U24037 (N_24037,N_23117,N_22597);
or U24038 (N_24038,N_22704,N_22599);
and U24039 (N_24039,N_22532,N_22835);
and U24040 (N_24040,N_22759,N_23478);
or U24041 (N_24041,N_23131,N_22845);
or U24042 (N_24042,N_22997,N_23380);
nand U24043 (N_24043,N_23019,N_22680);
and U24044 (N_24044,N_23447,N_23464);
nor U24045 (N_24045,N_22621,N_22990);
or U24046 (N_24046,N_22717,N_23934);
or U24047 (N_24047,N_23030,N_22628);
xor U24048 (N_24048,N_23489,N_22641);
nand U24049 (N_24049,N_23900,N_23509);
nor U24050 (N_24050,N_23554,N_23677);
xor U24051 (N_24051,N_23103,N_23193);
nand U24052 (N_24052,N_23000,N_23394);
xnor U24053 (N_24053,N_22854,N_23952);
nand U24054 (N_24054,N_23366,N_22760);
nor U24055 (N_24055,N_22744,N_22850);
or U24056 (N_24056,N_23991,N_23093);
and U24057 (N_24057,N_22855,N_23520);
nand U24058 (N_24058,N_22998,N_22693);
or U24059 (N_24059,N_23120,N_23866);
and U24060 (N_24060,N_23722,N_23339);
nor U24061 (N_24061,N_23004,N_22962);
nor U24062 (N_24062,N_22814,N_23169);
nand U24063 (N_24063,N_23986,N_23115);
nor U24064 (N_24064,N_22944,N_22518);
or U24065 (N_24065,N_23242,N_23811);
nand U24066 (N_24066,N_23558,N_22584);
nor U24067 (N_24067,N_23151,N_23303);
nand U24068 (N_24068,N_23816,N_22724);
and U24069 (N_24069,N_23451,N_22889);
and U24070 (N_24070,N_23008,N_23041);
and U24071 (N_24071,N_23174,N_22860);
nor U24072 (N_24072,N_22627,N_23226);
nor U24073 (N_24073,N_23281,N_23252);
or U24074 (N_24074,N_23132,N_22812);
or U24075 (N_24075,N_23446,N_22883);
xor U24076 (N_24076,N_23413,N_23538);
nand U24077 (N_24077,N_23310,N_23818);
nor U24078 (N_24078,N_22777,N_22920);
or U24079 (N_24079,N_22730,N_23608);
xnor U24080 (N_24080,N_23942,N_23425);
nor U24081 (N_24081,N_22506,N_22586);
xnor U24082 (N_24082,N_22712,N_23682);
xnor U24083 (N_24083,N_23481,N_23883);
xnor U24084 (N_24084,N_23302,N_23553);
or U24085 (N_24085,N_22650,N_23492);
nand U24086 (N_24086,N_23686,N_23049);
nor U24087 (N_24087,N_23245,N_22735);
nor U24088 (N_24088,N_23291,N_22977);
xnor U24089 (N_24089,N_23316,N_23614);
xnor U24090 (N_24090,N_22963,N_23441);
xnor U24091 (N_24091,N_23742,N_22587);
xor U24092 (N_24092,N_23386,N_23641);
or U24093 (N_24093,N_22549,N_23306);
nor U24094 (N_24094,N_23733,N_23269);
xnor U24095 (N_24095,N_22636,N_23850);
xnor U24096 (N_24096,N_23582,N_23995);
nor U24097 (N_24097,N_22736,N_23138);
nand U24098 (N_24098,N_23116,N_23749);
or U24099 (N_24099,N_23898,N_23695);
nor U24100 (N_24100,N_23703,N_22995);
and U24101 (N_24101,N_23593,N_22752);
or U24102 (N_24102,N_22754,N_23694);
xnor U24103 (N_24103,N_23985,N_23349);
or U24104 (N_24104,N_22706,N_23456);
and U24105 (N_24105,N_23356,N_23081);
or U24106 (N_24106,N_22799,N_23964);
nor U24107 (N_24107,N_23494,N_23691);
or U24108 (N_24108,N_23145,N_23603);
nor U24109 (N_24109,N_22992,N_22932);
xor U24110 (N_24110,N_22567,N_23851);
and U24111 (N_24111,N_23217,N_23951);
nand U24112 (N_24112,N_23336,N_23053);
and U24113 (N_24113,N_23890,N_23060);
and U24114 (N_24114,N_22741,N_23981);
nor U24115 (N_24115,N_23911,N_22525);
xnor U24116 (N_24116,N_22844,N_22594);
nor U24117 (N_24117,N_23769,N_22661);
or U24118 (N_24118,N_23240,N_23537);
nand U24119 (N_24119,N_22916,N_23491);
nand U24120 (N_24120,N_23244,N_22915);
xor U24121 (N_24121,N_23057,N_22978);
nor U24122 (N_24122,N_22521,N_23391);
nor U24123 (N_24123,N_22865,N_23253);
nand U24124 (N_24124,N_22536,N_23427);
nor U24125 (N_24125,N_22755,N_23927);
nor U24126 (N_24126,N_22642,N_22649);
and U24127 (N_24127,N_22828,N_23877);
or U24128 (N_24128,N_22764,N_22746);
nor U24129 (N_24129,N_23521,N_22512);
nand U24130 (N_24130,N_23073,N_22610);
xnor U24131 (N_24131,N_22581,N_23577);
or U24132 (N_24132,N_22598,N_23676);
or U24133 (N_24133,N_23243,N_23009);
nand U24134 (N_24134,N_22529,N_23842);
nor U24135 (N_24135,N_23598,N_23498);
nor U24136 (N_24136,N_23320,N_23058);
xor U24137 (N_24137,N_23267,N_23723);
and U24138 (N_24138,N_23384,N_23797);
and U24139 (N_24139,N_22602,N_22611);
xor U24140 (N_24140,N_23402,N_23328);
nor U24141 (N_24141,N_23322,N_23566);
and U24142 (N_24142,N_23458,N_23567);
nor U24143 (N_24143,N_23511,N_23337);
or U24144 (N_24144,N_23801,N_23438);
and U24145 (N_24145,N_23664,N_22657);
or U24146 (N_24146,N_23261,N_22546);
or U24147 (N_24147,N_22585,N_23987);
nand U24148 (N_24148,N_22504,N_23312);
and U24149 (N_24149,N_23398,N_23297);
nor U24150 (N_24150,N_22563,N_23585);
nand U24151 (N_24151,N_22846,N_23706);
and U24152 (N_24152,N_22766,N_22705);
or U24153 (N_24153,N_23711,N_23255);
xor U24154 (N_24154,N_23299,N_23815);
nand U24155 (N_24155,N_23365,N_23712);
or U24156 (N_24156,N_22681,N_23370);
nand U24157 (N_24157,N_22534,N_23065);
or U24158 (N_24158,N_23929,N_22707);
xnor U24159 (N_24159,N_22984,N_23238);
or U24160 (N_24160,N_23175,N_22790);
xor U24161 (N_24161,N_23615,N_23841);
xor U24162 (N_24162,N_23048,N_23529);
nand U24163 (N_24163,N_22878,N_23668);
nand U24164 (N_24164,N_22742,N_23550);
and U24165 (N_24165,N_23294,N_22667);
nand U24166 (N_24166,N_23050,N_23410);
nor U24167 (N_24167,N_23139,N_22936);
or U24168 (N_24168,N_23958,N_23836);
nor U24169 (N_24169,N_23647,N_22542);
or U24170 (N_24170,N_23201,N_22502);
xor U24171 (N_24171,N_22588,N_23062);
nor U24172 (N_24172,N_22873,N_23437);
and U24173 (N_24173,N_22576,N_23867);
nand U24174 (N_24174,N_22785,N_22806);
or U24175 (N_24175,N_23070,N_23110);
and U24176 (N_24176,N_23571,N_23804);
or U24177 (N_24177,N_23405,N_22538);
and U24178 (N_24178,N_23018,N_22696);
nor U24179 (N_24179,N_23028,N_23893);
nor U24180 (N_24180,N_23095,N_23725);
or U24181 (N_24181,N_23158,N_23595);
or U24182 (N_24182,N_22810,N_23275);
xor U24183 (N_24183,N_22537,N_22847);
xor U24184 (N_24184,N_23351,N_23228);
and U24185 (N_24185,N_22858,N_22976);
and U24186 (N_24186,N_23189,N_23375);
or U24187 (N_24187,N_23564,N_22901);
nand U24188 (N_24188,N_22609,N_22565);
nor U24189 (N_24189,N_23273,N_23869);
nand U24190 (N_24190,N_23936,N_23693);
nand U24191 (N_24191,N_23806,N_23460);
nor U24192 (N_24192,N_22793,N_22758);
nor U24193 (N_24193,N_23996,N_23221);
nand U24194 (N_24194,N_23755,N_23620);
nor U24195 (N_24195,N_23962,N_23001);
or U24196 (N_24196,N_23493,N_23516);
nand U24197 (N_24197,N_23914,N_23013);
or U24198 (N_24198,N_23670,N_23805);
nor U24199 (N_24199,N_22813,N_22624);
xor U24200 (N_24200,N_23335,N_23718);
xor U24201 (N_24201,N_22983,N_23989);
or U24202 (N_24202,N_23618,N_23527);
nor U24203 (N_24203,N_22662,N_23400);
nor U24204 (N_24204,N_23016,N_23782);
nand U24205 (N_24205,N_22876,N_23417);
and U24206 (N_24206,N_23462,N_22787);
nor U24207 (N_24207,N_22570,N_23681);
nor U24208 (N_24208,N_22648,N_22550);
nand U24209 (N_24209,N_23999,N_23917);
nor U24210 (N_24210,N_23581,N_23717);
nor U24211 (N_24211,N_22678,N_23823);
nor U24212 (N_24212,N_23837,N_22921);
xnor U24213 (N_24213,N_23086,N_23102);
xor U24214 (N_24214,N_23626,N_23781);
and U24215 (N_24215,N_23173,N_23715);
nor U24216 (N_24216,N_23023,N_23621);
nand U24217 (N_24217,N_23326,N_23206);
or U24218 (N_24218,N_23470,N_23500);
or U24219 (N_24219,N_23318,N_23324);
xor U24220 (N_24220,N_23125,N_22899);
or U24221 (N_24221,N_22508,N_23011);
xor U24222 (N_24222,N_23963,N_23141);
xnor U24223 (N_24223,N_22864,N_23531);
nand U24224 (N_24224,N_23534,N_23449);
xnor U24225 (N_24225,N_23416,N_23658);
nor U24226 (N_24226,N_22985,N_22692);
xnor U24227 (N_24227,N_23467,N_23916);
nand U24228 (N_24228,N_23039,N_23076);
nor U24229 (N_24229,N_22653,N_23428);
nand U24230 (N_24230,N_23508,N_22710);
nor U24231 (N_24231,N_22619,N_23932);
nand U24232 (N_24232,N_23469,N_23663);
xor U24233 (N_24233,N_23015,N_23465);
xor U24234 (N_24234,N_22957,N_22722);
xor U24235 (N_24235,N_23036,N_23378);
or U24236 (N_24236,N_23381,N_23955);
and U24237 (N_24237,N_23184,N_23532);
xnor U24238 (N_24238,N_23636,N_23109);
nand U24239 (N_24239,N_22753,N_23007);
or U24240 (N_24240,N_23975,N_23551);
nand U24241 (N_24241,N_23921,N_23640);
xor U24242 (N_24242,N_23388,N_23808);
or U24243 (N_24243,N_22798,N_23803);
or U24244 (N_24244,N_23440,N_22679);
or U24245 (N_24245,N_22817,N_23780);
xor U24246 (N_24246,N_23678,N_23194);
nand U24247 (N_24247,N_22971,N_22723);
or U24248 (N_24248,N_23080,N_22980);
nor U24249 (N_24249,N_23578,N_23988);
nand U24250 (N_24250,N_23107,N_22925);
nand U24251 (N_24251,N_23645,N_23289);
or U24252 (N_24252,N_22573,N_23099);
nor U24253 (N_24253,N_23215,N_23418);
nor U24254 (N_24254,N_23225,N_23147);
xor U24255 (N_24255,N_23431,N_22836);
and U24256 (N_24256,N_23072,N_22756);
nand U24257 (N_24257,N_23022,N_23231);
nor U24258 (N_24258,N_23475,N_22803);
nor U24259 (N_24259,N_22737,N_22800);
nand U24260 (N_24260,N_23843,N_23630);
or U24261 (N_24261,N_23341,N_22590);
nor U24262 (N_24262,N_23933,N_22711);
or U24263 (N_24263,N_23947,N_23497);
nand U24264 (N_24264,N_22913,N_22780);
xnor U24265 (N_24265,N_22929,N_23580);
and U24266 (N_24266,N_23387,N_23587);
and U24267 (N_24267,N_23176,N_22682);
nand U24268 (N_24268,N_23546,N_23859);
nand U24269 (N_24269,N_23482,N_23181);
nand U24270 (N_24270,N_23434,N_22931);
or U24271 (N_24271,N_23419,N_23807);
nand U24272 (N_24272,N_23619,N_23105);
nand U24273 (N_24273,N_22559,N_23443);
nor U24274 (N_24274,N_22986,N_23848);
nor U24275 (N_24275,N_23507,N_22630);
and U24276 (N_24276,N_23777,N_22886);
and U24277 (N_24277,N_23055,N_22954);
nand U24278 (N_24278,N_23730,N_23251);
xor U24279 (N_24279,N_22652,N_23455);
nor U24280 (N_24280,N_22870,N_23834);
or U24281 (N_24281,N_22687,N_23266);
or U24282 (N_24282,N_23922,N_23607);
nor U24283 (N_24283,N_23835,N_23857);
and U24284 (N_24284,N_23756,N_22975);
nor U24285 (N_24285,N_22688,N_23573);
nand U24286 (N_24286,N_22514,N_23894);
nor U24287 (N_24287,N_23510,N_22556);
or U24288 (N_24288,N_23536,N_22769);
or U24289 (N_24289,N_23533,N_23188);
xnor U24290 (N_24290,N_23282,N_23343);
nand U24291 (N_24291,N_23543,N_22815);
and U24292 (N_24292,N_23609,N_23920);
or U24293 (N_24293,N_23684,N_22659);
and U24294 (N_24294,N_22947,N_22909);
or U24295 (N_24295,N_23648,N_23436);
or U24296 (N_24296,N_22786,N_22767);
xor U24297 (N_24297,N_23170,N_23599);
and U24298 (N_24298,N_23892,N_22531);
or U24299 (N_24299,N_22721,N_22733);
xnor U24300 (N_24300,N_23372,N_23487);
and U24301 (N_24301,N_23887,N_22578);
nor U24302 (N_24302,N_23122,N_23068);
and U24303 (N_24303,N_22685,N_23003);
nand U24304 (N_24304,N_23937,N_23045);
xor U24305 (N_24305,N_23746,N_23833);
nor U24306 (N_24306,N_23421,N_23589);
xor U24307 (N_24307,N_23946,N_22981);
or U24308 (N_24308,N_23542,N_23787);
or U24309 (N_24309,N_23944,N_22524);
or U24310 (N_24310,N_23235,N_23526);
xnor U24311 (N_24311,N_23017,N_23878);
and U24312 (N_24312,N_23873,N_23838);
nand U24313 (N_24313,N_22796,N_23463);
or U24314 (N_24314,N_23790,N_23935);
nand U24315 (N_24315,N_23104,N_23424);
xor U24316 (N_24316,N_22684,N_23629);
nand U24317 (N_24317,N_23361,N_23171);
xor U24318 (N_24318,N_23627,N_23984);
nand U24319 (N_24319,N_22604,N_23814);
nand U24320 (N_24320,N_23512,N_22639);
xor U24321 (N_24321,N_23821,N_22867);
or U24322 (N_24322,N_22613,N_22625);
nand U24323 (N_24323,N_22727,N_23847);
nor U24324 (N_24324,N_22930,N_23098);
or U24325 (N_24325,N_23423,N_23972);
nand U24326 (N_24326,N_22953,N_23826);
nor U24327 (N_24327,N_23067,N_22819);
nor U24328 (N_24328,N_23290,N_23819);
xnor U24329 (N_24329,N_22956,N_23503);
nand U24330 (N_24330,N_22999,N_23259);
nor U24331 (N_24331,N_22664,N_23071);
or U24332 (N_24332,N_23404,N_23293);
xnor U24333 (N_24333,N_23654,N_23572);
nor U24334 (N_24334,N_23056,N_22884);
nand U24335 (N_24335,N_23471,N_23027);
nand U24336 (N_24336,N_23268,N_22905);
and U24337 (N_24337,N_22631,N_22959);
or U24338 (N_24338,N_23162,N_23100);
xor U24339 (N_24339,N_22928,N_23897);
and U24340 (N_24340,N_22789,N_22708);
or U24341 (N_24341,N_23993,N_22589);
and U24342 (N_24342,N_23575,N_22862);
nand U24343 (N_24343,N_23800,N_23347);
or U24344 (N_24344,N_23199,N_23736);
nor U24345 (N_24345,N_23344,N_22795);
and U24346 (N_24346,N_23006,N_23314);
or U24347 (N_24347,N_22871,N_23506);
nor U24348 (N_24348,N_23881,N_23832);
and U24349 (N_24349,N_23688,N_23948);
nand U24350 (N_24350,N_23655,N_23762);
and U24351 (N_24351,N_23026,N_22501);
nor U24352 (N_24352,N_23305,N_23864);
and U24353 (N_24353,N_23633,N_23237);
nand U24354 (N_24354,N_23700,N_23625);
nor U24355 (N_24355,N_23635,N_23234);
nand U24356 (N_24356,N_22516,N_23002);
nand U24357 (N_24357,N_22774,N_23278);
nor U24358 (N_24358,N_23524,N_23518);
nor U24359 (N_24359,N_23124,N_23118);
xor U24360 (N_24360,N_23123,N_23477);
or U24361 (N_24361,N_22683,N_23817);
xor U24362 (N_24362,N_23144,N_22991);
or U24363 (N_24363,N_23432,N_22771);
or U24364 (N_24364,N_23576,N_23544);
nor U24365 (N_24365,N_23250,N_23523);
nand U24366 (N_24366,N_23634,N_22666);
nand U24367 (N_24367,N_23484,N_23828);
nor U24368 (N_24368,N_22818,N_22993);
nor U24369 (N_24369,N_23998,N_23876);
nand U24370 (N_24370,N_23236,N_23295);
nand U24371 (N_24371,N_22715,N_23783);
xnor U24372 (N_24372,N_23659,N_23313);
nor U24373 (N_24373,N_23813,N_22903);
or U24374 (N_24374,N_23624,N_22555);
nor U24375 (N_24375,N_23042,N_23389);
nor U24376 (N_24376,N_23622,N_22842);
or U24377 (N_24377,N_23743,N_22988);
nor U24378 (N_24378,N_23172,N_23773);
xor U24379 (N_24379,N_23679,N_23683);
or U24380 (N_24380,N_23092,N_22961);
or U24381 (N_24381,N_23714,N_23829);
and U24382 (N_24382,N_23119,N_23687);
or U24383 (N_24383,N_22545,N_22824);
nand U24384 (N_24384,N_23383,N_22861);
and U24385 (N_24385,N_23101,N_23753);
and U24386 (N_24386,N_23216,N_23980);
nand U24387 (N_24387,N_23160,N_23870);
nand U24388 (N_24388,N_23795,N_23660);
nand U24389 (N_24389,N_23204,N_23439);
and U24390 (N_24390,N_22709,N_22548);
or U24391 (N_24391,N_23561,N_22779);
and U24392 (N_24392,N_23839,N_23457);
nand U24393 (N_24393,N_22513,N_23896);
and U24394 (N_24394,N_22517,N_22562);
or U24395 (N_24395,N_22640,N_23909);
and U24396 (N_24396,N_23161,N_23274);
nor U24397 (N_24397,N_23928,N_23501);
or U24398 (N_24398,N_22698,N_22772);
nand U24399 (N_24399,N_22579,N_23084);
xnor U24400 (N_24400,N_23971,N_23902);
xnor U24401 (N_24401,N_23959,N_23899);
xnor U24402 (N_24402,N_23149,N_22750);
nor U24403 (N_24403,N_23525,N_22637);
nor U24404 (N_24404,N_23309,N_22945);
or U24405 (N_24405,N_23632,N_22571);
and U24406 (N_24406,N_22658,N_22729);
xnor U24407 (N_24407,N_22857,N_22720);
nor U24408 (N_24408,N_23761,N_23854);
nor U24409 (N_24409,N_22569,N_23697);
nor U24410 (N_24410,N_23954,N_23930);
or U24411 (N_24411,N_23708,N_23696);
nor U24412 (N_24412,N_23570,N_23263);
or U24413 (N_24413,N_23209,N_22830);
xnor U24414 (N_24414,N_22601,N_23059);
xnor U24415 (N_24415,N_22906,N_23352);
and U24416 (N_24416,N_22703,N_22552);
nor U24417 (N_24417,N_23358,N_23367);
or U24418 (N_24418,N_22918,N_22701);
or U24419 (N_24419,N_22622,N_23163);
nand U24420 (N_24420,N_23032,N_23220);
nand U24421 (N_24421,N_23111,N_22544);
nand U24422 (N_24422,N_22510,N_23586);
xnor U24423 (N_24423,N_22673,N_23087);
or U24424 (N_24424,N_23637,N_23719);
xor U24425 (N_24425,N_23547,N_22561);
and U24426 (N_24426,N_23563,N_23392);
nand U24427 (N_24427,N_23304,N_22910);
nor U24428 (N_24428,N_23613,N_22574);
or U24429 (N_24429,N_23760,N_22989);
xnor U24430 (N_24430,N_23764,N_23364);
nand U24431 (N_24431,N_22895,N_23051);
xor U24432 (N_24432,N_23541,N_22738);
and U24433 (N_24433,N_22668,N_22827);
nor U24434 (N_24434,N_23338,N_22840);
nand U24435 (N_24435,N_23809,N_23014);
nand U24436 (N_24436,N_23090,N_23568);
or U24437 (N_24437,N_23710,N_22702);
and U24438 (N_24438,N_23415,N_22719);
or U24439 (N_24439,N_23445,N_23628);
and U24440 (N_24440,N_23738,N_23957);
nand U24441 (N_24441,N_23005,N_23129);
xnor U24442 (N_24442,N_23450,N_22645);
xnor U24443 (N_24443,N_22770,N_22872);
nor U24444 (N_24444,N_23043,N_23230);
or U24445 (N_24445,N_23222,N_23812);
nor U24446 (N_24446,N_23831,N_23943);
nand U24447 (N_24447,N_23114,N_23863);
nand U24448 (N_24448,N_23594,N_23794);
xor U24449 (N_24449,N_23368,N_23323);
xor U24450 (N_24450,N_23180,N_22881);
xnor U24451 (N_24451,N_22851,N_23020);
nand U24452 (N_24452,N_23130,N_23113);
and U24453 (N_24453,N_23860,N_23038);
or U24454 (N_24454,N_22922,N_23454);
xor U24455 (N_24455,N_23707,N_22955);
nand U24456 (N_24456,N_23148,N_23519);
nor U24457 (N_24457,N_23606,N_23374);
or U24458 (N_24458,N_23219,N_23342);
or U24459 (N_24459,N_22890,N_23472);
nor U24460 (N_24460,N_23938,N_23285);
nor U24461 (N_24461,N_22877,N_23168);
xnor U24462 (N_24462,N_23403,N_22583);
nor U24463 (N_24463,N_22911,N_23611);
nand U24464 (N_24464,N_23861,N_22775);
xnor U24465 (N_24465,N_23584,N_22926);
nand U24466 (N_24466,N_23406,N_23390);
and U24467 (N_24467,N_23698,N_23094);
or U24468 (N_24468,N_23751,N_23200);
nand U24469 (N_24469,N_22530,N_23750);
xnor U24470 (N_24470,N_23317,N_23940);
or U24471 (N_24471,N_23884,N_22933);
and U24472 (N_24472,N_23840,N_22964);
and U24473 (N_24473,N_23212,N_23674);
or U24474 (N_24474,N_23886,N_23941);
nand U24475 (N_24475,N_23401,N_22638);
xnor U24476 (N_24476,N_23820,N_23505);
nor U24477 (N_24477,N_22671,N_22654);
and U24478 (N_24478,N_23483,N_23397);
nor U24479 (N_24479,N_23588,N_23218);
nor U24480 (N_24480,N_23731,N_22831);
and U24481 (N_24481,N_22807,N_23974);
xnor U24482 (N_24482,N_23137,N_22633);
nand U24483 (N_24483,N_23106,N_22714);
and U24484 (N_24484,N_23150,N_22606);
or U24485 (N_24485,N_22938,N_23889);
and U24486 (N_24486,N_23667,N_22691);
xor U24487 (N_24487,N_23704,N_23191);
nor U24488 (N_24488,N_22617,N_22892);
and U24489 (N_24489,N_23966,N_22825);
and U24490 (N_24490,N_23748,N_23407);
nor U24491 (N_24491,N_22739,N_23379);
and U24492 (N_24492,N_23233,N_23208);
or U24493 (N_24493,N_23882,N_22820);
xor U24494 (N_24494,N_22541,N_22987);
and U24495 (N_24495,N_23047,N_22891);
nor U24496 (N_24496,N_23960,N_22821);
and U24497 (N_24497,N_22700,N_23720);
xor U24498 (N_24498,N_22694,N_23134);
nand U24499 (N_24499,N_23097,N_23798);
nand U24500 (N_24500,N_23597,N_23229);
and U24501 (N_24501,N_23596,N_23740);
xor U24502 (N_24502,N_22937,N_23452);
xor U24503 (N_24503,N_23223,N_23108);
nor U24504 (N_24504,N_23772,N_23775);
nand U24505 (N_24505,N_22672,N_23923);
or U24506 (N_24506,N_23956,N_22982);
xor U24507 (N_24507,N_22522,N_22731);
and U24508 (N_24508,N_23426,N_23369);
nand U24509 (N_24509,N_22600,N_23154);
or U24510 (N_24510,N_23286,N_23965);
nand U24511 (N_24511,N_22695,N_22551);
or U24512 (N_24512,N_22797,N_22826);
nor U24513 (N_24513,N_23555,N_23739);
xnor U24514 (N_24514,N_22970,N_23271);
or U24515 (N_24515,N_23246,N_23735);
xnor U24516 (N_24516,N_23758,N_23414);
xnor U24517 (N_24517,N_22608,N_23669);
nand U24518 (N_24518,N_23925,N_23583);
and U24519 (N_24519,N_23142,N_23385);
or U24520 (N_24520,N_22575,N_23203);
xnor U24521 (N_24521,N_22535,N_22794);
nor U24522 (N_24522,N_22949,N_22859);
nor U24523 (N_24523,N_23112,N_23517);
nand U24524 (N_24524,N_22699,N_23256);
nand U24525 (N_24525,N_22966,N_23734);
and U24526 (N_24526,N_23855,N_23513);
and U24527 (N_24527,N_22950,N_22503);
nor U24528 (N_24528,N_22943,N_22874);
or U24529 (N_24529,N_22591,N_22879);
and U24530 (N_24530,N_22743,N_23552);
nand U24531 (N_24531,N_23824,N_23545);
nand U24532 (N_24532,N_23888,N_23970);
xor U24533 (N_24533,N_22647,N_23673);
and U24534 (N_24534,N_23140,N_22823);
nor U24535 (N_24535,N_23579,N_22623);
or U24536 (N_24536,N_23591,N_22749);
and U24537 (N_24537,N_23918,N_23239);
and U24538 (N_24538,N_23354,N_23187);
nand U24539 (N_24539,N_23891,N_23759);
xnor U24540 (N_24540,N_23644,N_22540);
nand U24541 (N_24541,N_23270,N_22519);
xor U24542 (N_24542,N_22734,N_23178);
nor U24543 (N_24543,N_23862,N_23796);
nand U24544 (N_24544,N_23377,N_22868);
nor U24545 (N_24545,N_23907,N_23319);
nor U24546 (N_24546,N_23973,N_23393);
nor U24547 (N_24547,N_23858,N_23540);
and U24548 (N_24548,N_22686,N_22788);
xor U24549 (N_24549,N_23631,N_23021);
and U24550 (N_24550,N_22747,N_23198);
or U24551 (N_24551,N_23247,N_22596);
nor U24552 (N_24552,N_23224,N_23904);
or U24553 (N_24553,N_23953,N_22568);
nand U24554 (N_24554,N_23747,N_22716);
xnor U24555 (N_24555,N_23348,N_23033);
and U24556 (N_24556,N_23992,N_22935);
xnor U24557 (N_24557,N_22768,N_23190);
nor U24558 (N_24558,N_22566,N_23121);
and U24559 (N_24559,N_23779,N_22665);
or U24560 (N_24560,N_23827,N_23136);
xnor U24561 (N_24561,N_22757,N_23165);
xor U24562 (N_24562,N_23528,N_23474);
nor U24563 (N_24563,N_23325,N_23279);
nand U24564 (N_24564,N_23444,N_23292);
nor U24565 (N_24565,N_23549,N_23646);
or U24566 (N_24566,N_23926,N_22582);
or U24567 (N_24567,N_23311,N_23559);
xnor U24568 (N_24568,N_23331,N_23776);
or U24569 (N_24569,N_23284,N_23650);
or U24570 (N_24570,N_22888,N_22635);
xor U24571 (N_24571,N_23504,N_23288);
and U24572 (N_24572,N_22848,N_23355);
and U24573 (N_24573,N_23146,N_22782);
or U24574 (N_24574,N_23716,N_23262);
nor U24575 (N_24575,N_23064,N_22968);
and U24576 (N_24576,N_23671,N_22547);
nor U24577 (N_24577,N_22923,N_22773);
nand U24578 (N_24578,N_23063,N_22751);
xor U24579 (N_24579,N_23949,N_23466);
xnor U24580 (N_24580,N_23156,N_22974);
xor U24581 (N_24581,N_22880,N_22612);
or U24582 (N_24582,N_22778,N_23496);
or U24583 (N_24583,N_23665,N_22553);
nand U24584 (N_24584,N_23025,N_22934);
nand U24585 (N_24585,N_23562,N_22564);
xnor U24586 (N_24586,N_23079,N_22958);
nor U24587 (N_24587,N_23713,N_22897);
nor U24588 (N_24588,N_23468,N_23872);
xor U24589 (N_24589,N_23539,N_23257);
and U24590 (N_24590,N_22500,N_22669);
xor U24591 (N_24591,N_22802,N_23656);
xnor U24592 (N_24592,N_22792,N_23473);
or U24593 (N_24593,N_23557,N_22539);
or U24594 (N_24594,N_23945,N_22967);
or U24595 (N_24595,N_22675,N_23901);
and U24596 (N_24596,N_23638,N_23903);
nand U24597 (N_24597,N_23556,N_23874);
and U24598 (N_24598,N_23913,N_23091);
or U24599 (N_24599,N_23791,N_23702);
nor U24600 (N_24600,N_23069,N_22919);
xor U24601 (N_24601,N_22969,N_22725);
xor U24602 (N_24602,N_23672,N_22941);
nor U24603 (N_24603,N_23721,N_22626);
nor U24604 (N_24604,N_22776,N_23802);
and U24605 (N_24605,N_23301,N_23085);
or U24606 (N_24606,N_23430,N_22781);
xor U24607 (N_24607,N_23096,N_23906);
and U24608 (N_24608,N_23997,N_23675);
xor U24609 (N_24609,N_23411,N_22924);
xnor U24610 (N_24610,N_22973,N_22783);
or U24611 (N_24611,N_23592,N_23353);
and U24612 (N_24612,N_23083,N_23345);
xnor U24613 (N_24613,N_23034,N_22620);
and U24614 (N_24614,N_23155,N_22939);
and U24615 (N_24615,N_22839,N_22894);
and U24616 (N_24616,N_22801,N_22603);
xnor U24617 (N_24617,N_22904,N_22595);
or U24618 (N_24618,N_22605,N_22528);
and U24619 (N_24619,N_23729,N_22557);
and U24620 (N_24620,N_23442,N_23340);
and U24621 (N_24621,N_23535,N_22614);
nor U24622 (N_24622,N_23433,N_23185);
and U24623 (N_24623,N_23260,N_22520);
nand U24624 (N_24624,N_23362,N_22822);
and U24625 (N_24625,N_23651,N_23153);
nand U24626 (N_24626,N_23334,N_23810);
and U24627 (N_24627,N_22697,N_22740);
and U24628 (N_24628,N_22927,N_22527);
or U24629 (N_24629,N_23490,N_23037);
or U24630 (N_24630,N_23485,N_23329);
and U24631 (N_24631,N_22618,N_23300);
nand U24632 (N_24632,N_23705,N_23830);
nor U24633 (N_24633,N_23254,N_22885);
nand U24634 (N_24634,N_23601,N_23825);
and U24635 (N_24635,N_23359,N_23895);
or U24636 (N_24636,N_23024,N_23602);
nand U24637 (N_24637,N_22663,N_23196);
or U24638 (N_24638,N_22809,N_23249);
nand U24639 (N_24639,N_23258,N_23128);
xor U24640 (N_24640,N_22632,N_22960);
xnor U24641 (N_24641,N_23885,N_23692);
nor U24642 (N_24642,N_23357,N_23412);
or U24643 (N_24643,N_23409,N_22634);
nand U24644 (N_24644,N_23135,N_23177);
and U24645 (N_24645,N_22863,N_23610);
nand U24646 (N_24646,N_23616,N_23371);
or U24647 (N_24647,N_23910,N_23074);
or U24648 (N_24648,N_23784,N_23287);
xor U24649 (N_24649,N_22670,N_22656);
nor U24650 (N_24650,N_23799,N_23979);
xor U24651 (N_24651,N_22728,N_23774);
and U24652 (N_24652,N_22946,N_22948);
or U24653 (N_24653,N_23574,N_22543);
nand U24654 (N_24654,N_23661,N_23846);
and U24655 (N_24655,N_23210,N_22875);
nor U24656 (N_24656,N_22660,N_22689);
and U24657 (N_24657,N_23875,N_23363);
or U24658 (N_24658,N_22515,N_22834);
or U24659 (N_24659,N_23786,N_23332);
or U24660 (N_24660,N_22765,N_22748);
nand U24661 (N_24661,N_23479,N_22912);
xnor U24662 (N_24662,N_23088,N_23737);
xnor U24663 (N_24663,N_22763,N_22853);
nand U24664 (N_24664,N_23308,N_23977);
nor U24665 (N_24665,N_22676,N_22629);
and U24666 (N_24666,N_23754,N_23488);
nor U24667 (N_24667,N_22593,N_23054);
nand U24668 (N_24668,N_22837,N_23690);
and U24669 (N_24669,N_22507,N_23924);
or U24670 (N_24670,N_22866,N_22856);
nor U24671 (N_24671,N_22972,N_22833);
nor U24672 (N_24672,N_23939,N_23241);
xnor U24673 (N_24673,N_23197,N_23642);
nor U24674 (N_24674,N_23728,N_23012);
nand U24675 (N_24675,N_22523,N_22761);
or U24676 (N_24676,N_23968,N_23767);
or U24677 (N_24677,N_23315,N_23689);
nor U24678 (N_24678,N_22791,N_23082);
nand U24679 (N_24679,N_23530,N_22732);
nor U24680 (N_24680,N_22509,N_23652);
nand U24681 (N_24681,N_23649,N_22577);
nand U24682 (N_24682,N_22902,N_22917);
or U24683 (N_24683,N_23330,N_23849);
or U24684 (N_24684,N_23227,N_22808);
and U24685 (N_24685,N_23179,N_23515);
nand U24686 (N_24686,N_23276,N_23976);
nor U24687 (N_24687,N_23346,N_22951);
xor U24688 (N_24688,N_23046,N_23685);
and U24689 (N_24689,N_22898,N_22952);
xnor U24690 (N_24690,N_23031,N_22843);
and U24691 (N_24691,N_23395,N_23560);
nand U24692 (N_24692,N_23213,N_23662);
and U24693 (N_24693,N_22869,N_23066);
and U24694 (N_24694,N_23919,N_22655);
nand U24695 (N_24695,N_23569,N_23186);
and U24696 (N_24696,N_22505,N_23192);
or U24697 (N_24697,N_23277,N_23766);
and U24698 (N_24698,N_23844,N_23296);
nor U24699 (N_24699,N_23461,N_22816);
nand U24700 (N_24700,N_23133,N_23771);
xnor U24701 (N_24701,N_22572,N_23459);
and U24702 (N_24702,N_23763,N_23078);
nand U24703 (N_24703,N_23680,N_23726);
and U24704 (N_24704,N_23166,N_23195);
nor U24705 (N_24705,N_23422,N_23853);
or U24706 (N_24706,N_23499,N_23420);
nand U24707 (N_24707,N_23768,N_23868);
and U24708 (N_24708,N_23408,N_23126);
or U24709 (N_24709,N_23010,N_23453);
nor U24710 (N_24710,N_23605,N_22554);
nor U24711 (N_24711,N_22616,N_23152);
or U24712 (N_24712,N_22607,N_22718);
or U24713 (N_24713,N_23075,N_23061);
nor U24714 (N_24714,N_23350,N_23643);
and U24715 (N_24715,N_23265,N_23077);
nor U24716 (N_24716,N_23727,N_23264);
nor U24717 (N_24717,N_23880,N_23205);
or U24718 (N_24718,N_23040,N_23653);
nand U24719 (N_24719,N_23272,N_23931);
nand U24720 (N_24720,N_22979,N_23604);
nand U24721 (N_24721,N_22849,N_23476);
xor U24722 (N_24722,N_23961,N_23745);
or U24723 (N_24723,N_23143,N_22643);
and U24724 (N_24724,N_23871,N_23744);
nor U24725 (N_24725,N_23214,N_23701);
nand U24726 (N_24726,N_23327,N_23035);
xor U24727 (N_24727,N_22677,N_23856);
and U24728 (N_24728,N_23435,N_23548);
or U24729 (N_24729,N_22580,N_23865);
xor U24730 (N_24730,N_22893,N_23495);
nand U24731 (N_24731,N_22882,N_23699);
or U24732 (N_24732,N_22907,N_23429);
xor U24733 (N_24733,N_23207,N_23044);
and U24734 (N_24734,N_23211,N_23127);
and U24735 (N_24735,N_23785,N_22908);
nor U24736 (N_24736,N_23757,N_23778);
nand U24737 (N_24737,N_22784,N_23982);
and U24738 (N_24738,N_22511,N_23167);
nand U24739 (N_24739,N_22829,N_23448);
nor U24740 (N_24740,N_23202,N_23157);
and U24741 (N_24741,N_22651,N_22745);
xnor U24742 (N_24742,N_22900,N_23732);
xor U24743 (N_24743,N_23752,N_23623);
xor U24744 (N_24744,N_22533,N_23565);
nor U24745 (N_24745,N_23617,N_23248);
xnor U24746 (N_24746,N_23792,N_23480);
or U24747 (N_24747,N_22762,N_23280);
and U24748 (N_24748,N_22804,N_22838);
or U24749 (N_24749,N_22994,N_22526);
and U24750 (N_24750,N_23142,N_22510);
and U24751 (N_24751,N_23036,N_23159);
nor U24752 (N_24752,N_23356,N_23058);
and U24753 (N_24753,N_23141,N_23084);
and U24754 (N_24754,N_23309,N_23455);
and U24755 (N_24755,N_22697,N_23992);
nand U24756 (N_24756,N_22757,N_23861);
and U24757 (N_24757,N_23052,N_22510);
and U24758 (N_24758,N_23222,N_22974);
or U24759 (N_24759,N_23214,N_22910);
nor U24760 (N_24760,N_22846,N_22679);
nand U24761 (N_24761,N_23331,N_23285);
xor U24762 (N_24762,N_23176,N_22543);
and U24763 (N_24763,N_23733,N_23270);
or U24764 (N_24764,N_23523,N_23705);
or U24765 (N_24765,N_23281,N_23654);
or U24766 (N_24766,N_22977,N_23875);
or U24767 (N_24767,N_23286,N_23853);
nand U24768 (N_24768,N_23279,N_23602);
nand U24769 (N_24769,N_22580,N_22875);
nand U24770 (N_24770,N_23313,N_23101);
nand U24771 (N_24771,N_23147,N_22582);
and U24772 (N_24772,N_23381,N_23199);
or U24773 (N_24773,N_23185,N_23770);
nand U24774 (N_24774,N_22908,N_22785);
nor U24775 (N_24775,N_23389,N_23776);
or U24776 (N_24776,N_23684,N_23898);
nor U24777 (N_24777,N_22564,N_23395);
nor U24778 (N_24778,N_23460,N_23467);
or U24779 (N_24779,N_23325,N_23822);
and U24780 (N_24780,N_23062,N_22975);
nor U24781 (N_24781,N_22657,N_23452);
or U24782 (N_24782,N_23207,N_23040);
nand U24783 (N_24783,N_22910,N_23241);
nand U24784 (N_24784,N_23879,N_22758);
or U24785 (N_24785,N_23826,N_23072);
and U24786 (N_24786,N_23440,N_23466);
xor U24787 (N_24787,N_23454,N_23243);
xor U24788 (N_24788,N_23261,N_23124);
nand U24789 (N_24789,N_23118,N_22999);
and U24790 (N_24790,N_23844,N_23316);
xor U24791 (N_24791,N_23914,N_23767);
and U24792 (N_24792,N_22790,N_23161);
xnor U24793 (N_24793,N_23551,N_22511);
nor U24794 (N_24794,N_22702,N_23219);
xor U24795 (N_24795,N_23858,N_23264);
xor U24796 (N_24796,N_23370,N_23951);
and U24797 (N_24797,N_23908,N_23003);
nor U24798 (N_24798,N_23671,N_23346);
nand U24799 (N_24799,N_22783,N_23118);
xnor U24800 (N_24800,N_23693,N_22892);
and U24801 (N_24801,N_22640,N_23922);
xor U24802 (N_24802,N_22971,N_23654);
or U24803 (N_24803,N_23021,N_22743);
xor U24804 (N_24804,N_23509,N_22703);
xor U24805 (N_24805,N_23694,N_23268);
nor U24806 (N_24806,N_23932,N_23527);
or U24807 (N_24807,N_22634,N_22557);
nor U24808 (N_24808,N_22887,N_23296);
and U24809 (N_24809,N_23671,N_23505);
xor U24810 (N_24810,N_22615,N_23461);
or U24811 (N_24811,N_22989,N_23055);
xor U24812 (N_24812,N_22897,N_22914);
nand U24813 (N_24813,N_23132,N_22737);
or U24814 (N_24814,N_23950,N_22934);
or U24815 (N_24815,N_22747,N_22975);
or U24816 (N_24816,N_23486,N_23513);
or U24817 (N_24817,N_23447,N_23833);
or U24818 (N_24818,N_23217,N_23824);
and U24819 (N_24819,N_22849,N_23504);
xor U24820 (N_24820,N_22787,N_22729);
xor U24821 (N_24821,N_23798,N_23473);
or U24822 (N_24822,N_23774,N_22663);
xor U24823 (N_24823,N_23348,N_22692);
xor U24824 (N_24824,N_22722,N_23464);
xnor U24825 (N_24825,N_23787,N_22712);
or U24826 (N_24826,N_23488,N_23926);
or U24827 (N_24827,N_23476,N_23230);
or U24828 (N_24828,N_23845,N_23746);
and U24829 (N_24829,N_22700,N_23208);
nand U24830 (N_24830,N_22884,N_22823);
nor U24831 (N_24831,N_23993,N_22766);
or U24832 (N_24832,N_22820,N_22548);
xnor U24833 (N_24833,N_23150,N_23388);
nand U24834 (N_24834,N_23647,N_23862);
xor U24835 (N_24835,N_23077,N_22864);
or U24836 (N_24836,N_23165,N_22821);
nand U24837 (N_24837,N_23836,N_22952);
nor U24838 (N_24838,N_22616,N_22960);
nand U24839 (N_24839,N_23731,N_22942);
nand U24840 (N_24840,N_23505,N_22904);
nand U24841 (N_24841,N_23767,N_23475);
or U24842 (N_24842,N_22915,N_23286);
nand U24843 (N_24843,N_23862,N_23247);
nand U24844 (N_24844,N_22522,N_23602);
or U24845 (N_24845,N_23886,N_23958);
or U24846 (N_24846,N_23464,N_23271);
xnor U24847 (N_24847,N_22857,N_23711);
or U24848 (N_24848,N_23328,N_22927);
nor U24849 (N_24849,N_23267,N_23672);
or U24850 (N_24850,N_23975,N_23713);
and U24851 (N_24851,N_23292,N_23745);
and U24852 (N_24852,N_23137,N_23619);
xor U24853 (N_24853,N_23522,N_22753);
or U24854 (N_24854,N_22610,N_23756);
nor U24855 (N_24855,N_23412,N_23666);
nor U24856 (N_24856,N_23326,N_23420);
or U24857 (N_24857,N_23864,N_23336);
nand U24858 (N_24858,N_23016,N_23429);
or U24859 (N_24859,N_22565,N_23405);
nand U24860 (N_24860,N_23399,N_23503);
or U24861 (N_24861,N_23695,N_22516);
xnor U24862 (N_24862,N_22758,N_23893);
xor U24863 (N_24863,N_22889,N_23057);
nand U24864 (N_24864,N_23109,N_23385);
and U24865 (N_24865,N_22830,N_23131);
nand U24866 (N_24866,N_23816,N_22890);
nor U24867 (N_24867,N_23897,N_23665);
nor U24868 (N_24868,N_22797,N_23624);
or U24869 (N_24869,N_23982,N_22924);
nor U24870 (N_24870,N_22529,N_23241);
nand U24871 (N_24871,N_22970,N_23688);
or U24872 (N_24872,N_23372,N_23071);
and U24873 (N_24873,N_22799,N_23280);
or U24874 (N_24874,N_23769,N_22721);
nor U24875 (N_24875,N_22654,N_23413);
nand U24876 (N_24876,N_22934,N_23389);
and U24877 (N_24877,N_22746,N_23018);
nand U24878 (N_24878,N_23395,N_23732);
nand U24879 (N_24879,N_23480,N_23177);
nand U24880 (N_24880,N_23415,N_23325);
xor U24881 (N_24881,N_22745,N_22694);
xor U24882 (N_24882,N_22735,N_22696);
xor U24883 (N_24883,N_23478,N_23262);
or U24884 (N_24884,N_23776,N_23076);
xnor U24885 (N_24885,N_23013,N_23852);
nand U24886 (N_24886,N_23027,N_23747);
and U24887 (N_24887,N_22930,N_23659);
xor U24888 (N_24888,N_22512,N_23165);
nand U24889 (N_24889,N_22753,N_23387);
or U24890 (N_24890,N_23537,N_22622);
and U24891 (N_24891,N_23792,N_23862);
or U24892 (N_24892,N_23723,N_22834);
or U24893 (N_24893,N_22809,N_23815);
xnor U24894 (N_24894,N_23012,N_23456);
nor U24895 (N_24895,N_23271,N_23534);
nand U24896 (N_24896,N_23321,N_22943);
xor U24897 (N_24897,N_22981,N_23479);
nand U24898 (N_24898,N_23459,N_23997);
nor U24899 (N_24899,N_23162,N_23105);
and U24900 (N_24900,N_23317,N_23835);
xor U24901 (N_24901,N_22675,N_23919);
or U24902 (N_24902,N_23802,N_22690);
nand U24903 (N_24903,N_22701,N_23174);
xor U24904 (N_24904,N_23412,N_23452);
nand U24905 (N_24905,N_23907,N_22526);
xor U24906 (N_24906,N_23888,N_23805);
nand U24907 (N_24907,N_23264,N_23090);
nor U24908 (N_24908,N_22540,N_23868);
xnor U24909 (N_24909,N_23011,N_23093);
nand U24910 (N_24910,N_23753,N_23621);
and U24911 (N_24911,N_23208,N_22970);
nor U24912 (N_24912,N_22959,N_22540);
nand U24913 (N_24913,N_23159,N_23543);
nor U24914 (N_24914,N_22557,N_23139);
or U24915 (N_24915,N_23853,N_23708);
and U24916 (N_24916,N_23274,N_23065);
xor U24917 (N_24917,N_22668,N_22873);
nand U24918 (N_24918,N_23977,N_23540);
or U24919 (N_24919,N_23173,N_23057);
and U24920 (N_24920,N_22510,N_23546);
or U24921 (N_24921,N_22862,N_22950);
xor U24922 (N_24922,N_23553,N_23645);
or U24923 (N_24923,N_22557,N_23662);
or U24924 (N_24924,N_23006,N_22935);
xor U24925 (N_24925,N_22501,N_23180);
xor U24926 (N_24926,N_22634,N_23008);
xor U24927 (N_24927,N_23437,N_22577);
xnor U24928 (N_24928,N_22837,N_23992);
nand U24929 (N_24929,N_23313,N_23455);
or U24930 (N_24930,N_23129,N_23647);
nand U24931 (N_24931,N_22586,N_23337);
or U24932 (N_24932,N_22921,N_23055);
nand U24933 (N_24933,N_23110,N_23001);
xor U24934 (N_24934,N_22712,N_23894);
nand U24935 (N_24935,N_23861,N_23466);
xnor U24936 (N_24936,N_22665,N_23241);
or U24937 (N_24937,N_23507,N_22995);
or U24938 (N_24938,N_23517,N_22948);
and U24939 (N_24939,N_23974,N_23094);
nor U24940 (N_24940,N_22962,N_23133);
nor U24941 (N_24941,N_23045,N_23652);
nand U24942 (N_24942,N_23763,N_23868);
xor U24943 (N_24943,N_23220,N_22925);
or U24944 (N_24944,N_23913,N_22719);
xor U24945 (N_24945,N_23090,N_23598);
xor U24946 (N_24946,N_22651,N_23765);
nand U24947 (N_24947,N_22943,N_23599);
nor U24948 (N_24948,N_23545,N_22935);
and U24949 (N_24949,N_23957,N_22597);
nor U24950 (N_24950,N_23893,N_22537);
nor U24951 (N_24951,N_22695,N_22576);
and U24952 (N_24952,N_22937,N_22858);
and U24953 (N_24953,N_23579,N_23580);
nor U24954 (N_24954,N_23698,N_22870);
nor U24955 (N_24955,N_23166,N_23276);
nand U24956 (N_24956,N_22896,N_23751);
nand U24957 (N_24957,N_23864,N_23121);
or U24958 (N_24958,N_23859,N_23969);
and U24959 (N_24959,N_23991,N_23529);
nand U24960 (N_24960,N_22910,N_23195);
xnor U24961 (N_24961,N_22617,N_23651);
nand U24962 (N_24962,N_22616,N_22699);
xor U24963 (N_24963,N_23161,N_23152);
xnor U24964 (N_24964,N_23706,N_22782);
nor U24965 (N_24965,N_22691,N_22690);
nor U24966 (N_24966,N_23061,N_23693);
nand U24967 (N_24967,N_23549,N_23495);
xor U24968 (N_24968,N_23269,N_23334);
nand U24969 (N_24969,N_23982,N_23347);
nand U24970 (N_24970,N_22946,N_23983);
or U24971 (N_24971,N_23542,N_23577);
xor U24972 (N_24972,N_23166,N_23900);
or U24973 (N_24973,N_23025,N_23689);
or U24974 (N_24974,N_22669,N_23289);
and U24975 (N_24975,N_23692,N_22506);
or U24976 (N_24976,N_23362,N_22863);
or U24977 (N_24977,N_22883,N_23127);
xor U24978 (N_24978,N_23682,N_23749);
or U24979 (N_24979,N_22504,N_23418);
or U24980 (N_24980,N_23371,N_22943);
or U24981 (N_24981,N_22943,N_23126);
xnor U24982 (N_24982,N_23963,N_22514);
nand U24983 (N_24983,N_23060,N_22819);
nor U24984 (N_24984,N_22601,N_22518);
xor U24985 (N_24985,N_22903,N_23999);
or U24986 (N_24986,N_22740,N_22967);
xnor U24987 (N_24987,N_23458,N_22694);
nand U24988 (N_24988,N_22655,N_22758);
nand U24989 (N_24989,N_23237,N_23724);
nor U24990 (N_24990,N_23568,N_22804);
xnor U24991 (N_24991,N_22703,N_22618);
nor U24992 (N_24992,N_22675,N_23896);
nand U24993 (N_24993,N_23099,N_23408);
and U24994 (N_24994,N_22881,N_23785);
nand U24995 (N_24995,N_22515,N_23489);
and U24996 (N_24996,N_22936,N_23878);
or U24997 (N_24997,N_22979,N_22818);
or U24998 (N_24998,N_22733,N_23498);
nand U24999 (N_24999,N_23517,N_23045);
nand U25000 (N_25000,N_23202,N_23353);
or U25001 (N_25001,N_23122,N_23406);
nand U25002 (N_25002,N_22984,N_23865);
nand U25003 (N_25003,N_22535,N_23199);
nand U25004 (N_25004,N_23569,N_23309);
or U25005 (N_25005,N_22818,N_22556);
nor U25006 (N_25006,N_22923,N_23118);
and U25007 (N_25007,N_23575,N_23855);
nand U25008 (N_25008,N_23622,N_23487);
or U25009 (N_25009,N_23409,N_22507);
nor U25010 (N_25010,N_22788,N_23239);
xnor U25011 (N_25011,N_22772,N_23561);
nor U25012 (N_25012,N_22789,N_23451);
xnor U25013 (N_25013,N_22538,N_23436);
nand U25014 (N_25014,N_23595,N_22587);
or U25015 (N_25015,N_22970,N_23588);
nand U25016 (N_25016,N_23779,N_23344);
xnor U25017 (N_25017,N_23183,N_23909);
nand U25018 (N_25018,N_22583,N_23755);
nand U25019 (N_25019,N_23129,N_22901);
nand U25020 (N_25020,N_23532,N_22532);
or U25021 (N_25021,N_23012,N_23892);
and U25022 (N_25022,N_22606,N_23959);
xnor U25023 (N_25023,N_23341,N_23010);
or U25024 (N_25024,N_23735,N_23112);
nor U25025 (N_25025,N_23677,N_23571);
nor U25026 (N_25026,N_23600,N_23473);
nor U25027 (N_25027,N_23808,N_22747);
or U25028 (N_25028,N_23035,N_23178);
nor U25029 (N_25029,N_23640,N_22593);
and U25030 (N_25030,N_23828,N_22957);
or U25031 (N_25031,N_23196,N_23699);
xor U25032 (N_25032,N_23209,N_23555);
xor U25033 (N_25033,N_22597,N_23265);
and U25034 (N_25034,N_23084,N_22553);
nand U25035 (N_25035,N_22732,N_23747);
nand U25036 (N_25036,N_22682,N_23955);
xnor U25037 (N_25037,N_23393,N_23429);
nor U25038 (N_25038,N_23160,N_23448);
or U25039 (N_25039,N_23441,N_22769);
and U25040 (N_25040,N_23250,N_22636);
or U25041 (N_25041,N_22672,N_22950);
nor U25042 (N_25042,N_22810,N_23035);
nor U25043 (N_25043,N_22797,N_23684);
nor U25044 (N_25044,N_22507,N_22838);
or U25045 (N_25045,N_22507,N_22891);
or U25046 (N_25046,N_22960,N_23969);
and U25047 (N_25047,N_22914,N_23457);
xor U25048 (N_25048,N_23723,N_23570);
or U25049 (N_25049,N_23590,N_23096);
and U25050 (N_25050,N_23447,N_23608);
and U25051 (N_25051,N_23386,N_23042);
or U25052 (N_25052,N_23506,N_22914);
and U25053 (N_25053,N_22646,N_23455);
nor U25054 (N_25054,N_23442,N_23246);
and U25055 (N_25055,N_22976,N_23127);
nor U25056 (N_25056,N_23105,N_22855);
or U25057 (N_25057,N_23353,N_23386);
nand U25058 (N_25058,N_23557,N_23535);
nor U25059 (N_25059,N_23642,N_22835);
and U25060 (N_25060,N_23615,N_22998);
or U25061 (N_25061,N_23462,N_23388);
and U25062 (N_25062,N_23144,N_23707);
xnor U25063 (N_25063,N_23738,N_23510);
xor U25064 (N_25064,N_23178,N_23953);
and U25065 (N_25065,N_23305,N_22543);
and U25066 (N_25066,N_23049,N_23698);
nand U25067 (N_25067,N_23499,N_22859);
or U25068 (N_25068,N_23876,N_23596);
and U25069 (N_25069,N_23388,N_23335);
nand U25070 (N_25070,N_23285,N_23714);
nand U25071 (N_25071,N_23956,N_22574);
nand U25072 (N_25072,N_22523,N_22611);
or U25073 (N_25073,N_23921,N_23329);
and U25074 (N_25074,N_23979,N_22539);
and U25075 (N_25075,N_23682,N_23802);
nand U25076 (N_25076,N_23680,N_22900);
nor U25077 (N_25077,N_23529,N_23820);
nand U25078 (N_25078,N_22655,N_23695);
and U25079 (N_25079,N_23561,N_23626);
nand U25080 (N_25080,N_23196,N_23393);
and U25081 (N_25081,N_23176,N_23657);
xor U25082 (N_25082,N_23928,N_23090);
and U25083 (N_25083,N_23484,N_23066);
nor U25084 (N_25084,N_23548,N_22746);
and U25085 (N_25085,N_23377,N_23503);
xor U25086 (N_25086,N_22756,N_23588);
and U25087 (N_25087,N_22925,N_23649);
or U25088 (N_25088,N_23104,N_22950);
or U25089 (N_25089,N_23388,N_23555);
or U25090 (N_25090,N_23593,N_23361);
xnor U25091 (N_25091,N_22713,N_22710);
nor U25092 (N_25092,N_23481,N_23354);
nor U25093 (N_25093,N_23810,N_23561);
and U25094 (N_25094,N_22853,N_22786);
nand U25095 (N_25095,N_23225,N_23848);
xnor U25096 (N_25096,N_22832,N_23907);
and U25097 (N_25097,N_23661,N_23273);
or U25098 (N_25098,N_23799,N_22951);
or U25099 (N_25099,N_22854,N_23188);
and U25100 (N_25100,N_23377,N_23118);
or U25101 (N_25101,N_23771,N_23798);
or U25102 (N_25102,N_23720,N_22664);
nor U25103 (N_25103,N_22879,N_22848);
nor U25104 (N_25104,N_23246,N_23270);
nand U25105 (N_25105,N_22793,N_23728);
nor U25106 (N_25106,N_23259,N_23542);
nand U25107 (N_25107,N_23958,N_23138);
or U25108 (N_25108,N_22561,N_23793);
xor U25109 (N_25109,N_23844,N_22566);
nor U25110 (N_25110,N_23076,N_23981);
and U25111 (N_25111,N_23281,N_22991);
and U25112 (N_25112,N_22634,N_23720);
nand U25113 (N_25113,N_22614,N_23605);
xnor U25114 (N_25114,N_23151,N_23457);
nand U25115 (N_25115,N_23371,N_23696);
nand U25116 (N_25116,N_23665,N_22890);
nor U25117 (N_25117,N_23235,N_23606);
nand U25118 (N_25118,N_23510,N_23443);
nor U25119 (N_25119,N_22999,N_22707);
nand U25120 (N_25120,N_23080,N_22800);
or U25121 (N_25121,N_22890,N_23390);
or U25122 (N_25122,N_23444,N_23967);
nand U25123 (N_25123,N_23307,N_22657);
xnor U25124 (N_25124,N_23974,N_23507);
or U25125 (N_25125,N_23531,N_23467);
or U25126 (N_25126,N_23846,N_22890);
xor U25127 (N_25127,N_23904,N_23289);
nor U25128 (N_25128,N_23426,N_22562);
nand U25129 (N_25129,N_22517,N_23592);
xor U25130 (N_25130,N_23105,N_23449);
nand U25131 (N_25131,N_23458,N_22916);
xnor U25132 (N_25132,N_23598,N_23939);
or U25133 (N_25133,N_23339,N_23775);
xnor U25134 (N_25134,N_22662,N_23230);
and U25135 (N_25135,N_23702,N_22918);
xor U25136 (N_25136,N_23204,N_23434);
nor U25137 (N_25137,N_23892,N_23668);
and U25138 (N_25138,N_22890,N_22900);
nand U25139 (N_25139,N_23486,N_23913);
and U25140 (N_25140,N_22999,N_22529);
xnor U25141 (N_25141,N_22571,N_23414);
or U25142 (N_25142,N_22597,N_23135);
or U25143 (N_25143,N_22997,N_23690);
or U25144 (N_25144,N_22558,N_23520);
xor U25145 (N_25145,N_23287,N_23140);
nand U25146 (N_25146,N_23242,N_23932);
nor U25147 (N_25147,N_23175,N_23384);
xnor U25148 (N_25148,N_22908,N_22750);
xnor U25149 (N_25149,N_22831,N_23861);
nand U25150 (N_25150,N_22649,N_23141);
nand U25151 (N_25151,N_23303,N_23625);
nor U25152 (N_25152,N_23194,N_22994);
and U25153 (N_25153,N_23984,N_22805);
and U25154 (N_25154,N_23913,N_23071);
or U25155 (N_25155,N_23153,N_23199);
nor U25156 (N_25156,N_23658,N_23883);
nand U25157 (N_25157,N_23775,N_23172);
nand U25158 (N_25158,N_23438,N_23605);
nand U25159 (N_25159,N_22828,N_23637);
and U25160 (N_25160,N_22779,N_23447);
or U25161 (N_25161,N_23877,N_22993);
and U25162 (N_25162,N_22529,N_22642);
and U25163 (N_25163,N_22905,N_23768);
xnor U25164 (N_25164,N_23850,N_22712);
and U25165 (N_25165,N_23594,N_23829);
xnor U25166 (N_25166,N_23483,N_23369);
or U25167 (N_25167,N_23615,N_23510);
nand U25168 (N_25168,N_22675,N_23476);
or U25169 (N_25169,N_22596,N_23548);
and U25170 (N_25170,N_22882,N_23623);
or U25171 (N_25171,N_23893,N_23683);
nor U25172 (N_25172,N_22673,N_22761);
or U25173 (N_25173,N_23434,N_23470);
xnor U25174 (N_25174,N_22737,N_23550);
and U25175 (N_25175,N_23086,N_23453);
nor U25176 (N_25176,N_22557,N_22619);
nand U25177 (N_25177,N_23283,N_23899);
and U25178 (N_25178,N_23395,N_23791);
nor U25179 (N_25179,N_22641,N_23081);
nand U25180 (N_25180,N_23381,N_23546);
nor U25181 (N_25181,N_23456,N_23679);
xnor U25182 (N_25182,N_23939,N_22824);
xnor U25183 (N_25183,N_23473,N_22723);
nor U25184 (N_25184,N_23680,N_23325);
nand U25185 (N_25185,N_23908,N_23756);
and U25186 (N_25186,N_22872,N_22780);
xor U25187 (N_25187,N_23868,N_23329);
nand U25188 (N_25188,N_23136,N_23049);
and U25189 (N_25189,N_23970,N_23765);
or U25190 (N_25190,N_23392,N_22957);
or U25191 (N_25191,N_22759,N_23965);
and U25192 (N_25192,N_23483,N_22502);
and U25193 (N_25193,N_23198,N_22551);
xnor U25194 (N_25194,N_23462,N_22537);
nor U25195 (N_25195,N_23294,N_22544);
nand U25196 (N_25196,N_23105,N_23142);
and U25197 (N_25197,N_22569,N_22693);
xnor U25198 (N_25198,N_23728,N_23721);
and U25199 (N_25199,N_22544,N_23645);
and U25200 (N_25200,N_22508,N_22876);
nand U25201 (N_25201,N_22558,N_23575);
xor U25202 (N_25202,N_23787,N_23096);
nand U25203 (N_25203,N_23167,N_22652);
and U25204 (N_25204,N_23627,N_23922);
and U25205 (N_25205,N_23884,N_23991);
nand U25206 (N_25206,N_22614,N_23786);
nor U25207 (N_25207,N_23865,N_23300);
nand U25208 (N_25208,N_23330,N_22550);
and U25209 (N_25209,N_23432,N_23655);
and U25210 (N_25210,N_23600,N_22636);
and U25211 (N_25211,N_23053,N_23873);
nand U25212 (N_25212,N_23464,N_23834);
xnor U25213 (N_25213,N_23943,N_23186);
nand U25214 (N_25214,N_23928,N_23115);
or U25215 (N_25215,N_22763,N_23935);
xor U25216 (N_25216,N_23433,N_23006);
nor U25217 (N_25217,N_22757,N_23634);
or U25218 (N_25218,N_22538,N_23398);
xor U25219 (N_25219,N_23672,N_22533);
nor U25220 (N_25220,N_22825,N_23495);
xnor U25221 (N_25221,N_23658,N_23769);
xnor U25222 (N_25222,N_23211,N_23357);
nor U25223 (N_25223,N_23459,N_23687);
nand U25224 (N_25224,N_23880,N_23489);
nor U25225 (N_25225,N_22690,N_22566);
xor U25226 (N_25226,N_23067,N_22649);
xor U25227 (N_25227,N_22860,N_22843);
or U25228 (N_25228,N_23483,N_22689);
and U25229 (N_25229,N_22585,N_23037);
nor U25230 (N_25230,N_22633,N_22727);
or U25231 (N_25231,N_23367,N_22572);
nand U25232 (N_25232,N_23055,N_23221);
and U25233 (N_25233,N_23820,N_23254);
xnor U25234 (N_25234,N_23892,N_22782);
nand U25235 (N_25235,N_23473,N_22615);
or U25236 (N_25236,N_23566,N_22557);
and U25237 (N_25237,N_23279,N_22832);
or U25238 (N_25238,N_23266,N_23061);
xor U25239 (N_25239,N_23003,N_22531);
and U25240 (N_25240,N_22883,N_23032);
nand U25241 (N_25241,N_23411,N_22962);
xnor U25242 (N_25242,N_22857,N_22599);
nand U25243 (N_25243,N_23757,N_23785);
and U25244 (N_25244,N_23865,N_22957);
or U25245 (N_25245,N_22958,N_22590);
nand U25246 (N_25246,N_23328,N_22887);
xor U25247 (N_25247,N_22687,N_23932);
or U25248 (N_25248,N_22868,N_22746);
or U25249 (N_25249,N_22857,N_23527);
or U25250 (N_25250,N_23837,N_23598);
xor U25251 (N_25251,N_22994,N_23728);
xnor U25252 (N_25252,N_23460,N_23678);
or U25253 (N_25253,N_22960,N_22916);
or U25254 (N_25254,N_22555,N_23168);
nor U25255 (N_25255,N_22705,N_23479);
xor U25256 (N_25256,N_23391,N_23344);
and U25257 (N_25257,N_22829,N_22643);
and U25258 (N_25258,N_23613,N_23880);
xnor U25259 (N_25259,N_23679,N_22963);
xor U25260 (N_25260,N_23856,N_22752);
nand U25261 (N_25261,N_23015,N_22946);
or U25262 (N_25262,N_22783,N_23772);
or U25263 (N_25263,N_23969,N_23869);
nand U25264 (N_25264,N_23854,N_23258);
nand U25265 (N_25265,N_23273,N_23112);
nor U25266 (N_25266,N_23774,N_23563);
xor U25267 (N_25267,N_23885,N_23557);
nor U25268 (N_25268,N_23997,N_23632);
or U25269 (N_25269,N_23000,N_22664);
xnor U25270 (N_25270,N_22735,N_23764);
nand U25271 (N_25271,N_23713,N_23608);
and U25272 (N_25272,N_23991,N_23626);
nand U25273 (N_25273,N_22766,N_23951);
nor U25274 (N_25274,N_23056,N_23490);
or U25275 (N_25275,N_22695,N_23977);
nor U25276 (N_25276,N_23226,N_22918);
nand U25277 (N_25277,N_23931,N_23810);
nor U25278 (N_25278,N_22748,N_22941);
xnor U25279 (N_25279,N_22728,N_23992);
and U25280 (N_25280,N_23264,N_22971);
and U25281 (N_25281,N_23146,N_23526);
and U25282 (N_25282,N_22547,N_23346);
nand U25283 (N_25283,N_23981,N_23519);
xnor U25284 (N_25284,N_23821,N_23133);
nand U25285 (N_25285,N_22963,N_22821);
nand U25286 (N_25286,N_23438,N_23659);
nand U25287 (N_25287,N_23054,N_23243);
nor U25288 (N_25288,N_23532,N_23666);
xor U25289 (N_25289,N_22610,N_23170);
and U25290 (N_25290,N_22596,N_22578);
nand U25291 (N_25291,N_23688,N_23565);
or U25292 (N_25292,N_23770,N_22624);
xnor U25293 (N_25293,N_23070,N_23235);
xnor U25294 (N_25294,N_23763,N_23487);
xor U25295 (N_25295,N_23750,N_23228);
or U25296 (N_25296,N_22590,N_23814);
or U25297 (N_25297,N_23451,N_22852);
xor U25298 (N_25298,N_23171,N_23327);
or U25299 (N_25299,N_23522,N_23773);
and U25300 (N_25300,N_23436,N_23403);
or U25301 (N_25301,N_22926,N_23016);
nor U25302 (N_25302,N_23349,N_22920);
nor U25303 (N_25303,N_23569,N_22735);
or U25304 (N_25304,N_22934,N_22818);
nand U25305 (N_25305,N_23305,N_23015);
or U25306 (N_25306,N_23907,N_23736);
and U25307 (N_25307,N_22988,N_23836);
nand U25308 (N_25308,N_23740,N_22858);
nand U25309 (N_25309,N_22806,N_23480);
xnor U25310 (N_25310,N_23955,N_23916);
nor U25311 (N_25311,N_23725,N_23074);
nor U25312 (N_25312,N_22780,N_23338);
nor U25313 (N_25313,N_22842,N_23117);
or U25314 (N_25314,N_22661,N_23960);
xnor U25315 (N_25315,N_23186,N_23313);
nor U25316 (N_25316,N_23830,N_23843);
and U25317 (N_25317,N_22934,N_23496);
nand U25318 (N_25318,N_23952,N_23358);
xor U25319 (N_25319,N_23662,N_23543);
or U25320 (N_25320,N_22969,N_22590);
nand U25321 (N_25321,N_23823,N_22700);
xor U25322 (N_25322,N_23371,N_23340);
xnor U25323 (N_25323,N_22782,N_23583);
nor U25324 (N_25324,N_23780,N_22741);
nand U25325 (N_25325,N_23048,N_23039);
nor U25326 (N_25326,N_23207,N_22648);
or U25327 (N_25327,N_23575,N_23696);
nor U25328 (N_25328,N_23386,N_23809);
and U25329 (N_25329,N_22628,N_23445);
or U25330 (N_25330,N_23575,N_23229);
and U25331 (N_25331,N_23671,N_23619);
nor U25332 (N_25332,N_23989,N_23728);
or U25333 (N_25333,N_23019,N_22965);
nor U25334 (N_25334,N_23034,N_22905);
or U25335 (N_25335,N_23550,N_22782);
or U25336 (N_25336,N_23915,N_22623);
and U25337 (N_25337,N_23304,N_23934);
nand U25338 (N_25338,N_23643,N_23740);
xor U25339 (N_25339,N_23927,N_22909);
and U25340 (N_25340,N_22800,N_23629);
nor U25341 (N_25341,N_23837,N_22520);
xor U25342 (N_25342,N_23452,N_23598);
or U25343 (N_25343,N_23179,N_23125);
nor U25344 (N_25344,N_22549,N_23760);
nor U25345 (N_25345,N_22677,N_22809);
and U25346 (N_25346,N_23252,N_23457);
nand U25347 (N_25347,N_23024,N_23387);
or U25348 (N_25348,N_22610,N_23975);
or U25349 (N_25349,N_22722,N_23064);
nand U25350 (N_25350,N_23483,N_23480);
nand U25351 (N_25351,N_22867,N_23143);
nand U25352 (N_25352,N_23830,N_22531);
or U25353 (N_25353,N_22543,N_23898);
xnor U25354 (N_25354,N_23179,N_23424);
and U25355 (N_25355,N_23339,N_22641);
nor U25356 (N_25356,N_22703,N_23641);
nor U25357 (N_25357,N_23832,N_23954);
and U25358 (N_25358,N_22532,N_22589);
xnor U25359 (N_25359,N_23579,N_22889);
nand U25360 (N_25360,N_23415,N_23974);
nor U25361 (N_25361,N_22918,N_22971);
and U25362 (N_25362,N_22787,N_23931);
xor U25363 (N_25363,N_23680,N_23739);
nor U25364 (N_25364,N_22771,N_23503);
or U25365 (N_25365,N_23330,N_22590);
nor U25366 (N_25366,N_22971,N_23150);
and U25367 (N_25367,N_23508,N_23779);
nor U25368 (N_25368,N_22968,N_23802);
nand U25369 (N_25369,N_23259,N_22546);
nand U25370 (N_25370,N_22547,N_23951);
nor U25371 (N_25371,N_23489,N_23054);
nand U25372 (N_25372,N_23693,N_23383);
xor U25373 (N_25373,N_22715,N_22801);
xnor U25374 (N_25374,N_23219,N_23236);
xnor U25375 (N_25375,N_22948,N_22903);
nand U25376 (N_25376,N_22573,N_23809);
or U25377 (N_25377,N_23724,N_23083);
or U25378 (N_25378,N_23640,N_23134);
xor U25379 (N_25379,N_22987,N_23936);
nor U25380 (N_25380,N_22688,N_22796);
xnor U25381 (N_25381,N_22896,N_23333);
and U25382 (N_25382,N_22790,N_23699);
xor U25383 (N_25383,N_23754,N_23356);
nand U25384 (N_25384,N_23160,N_22688);
or U25385 (N_25385,N_23646,N_23291);
or U25386 (N_25386,N_22917,N_23610);
or U25387 (N_25387,N_23751,N_22998);
nand U25388 (N_25388,N_23288,N_23175);
nor U25389 (N_25389,N_23263,N_22887);
nand U25390 (N_25390,N_22672,N_22675);
xor U25391 (N_25391,N_23592,N_22582);
nand U25392 (N_25392,N_23250,N_23718);
nor U25393 (N_25393,N_23353,N_22596);
or U25394 (N_25394,N_23566,N_22934);
and U25395 (N_25395,N_23457,N_23610);
and U25396 (N_25396,N_23426,N_22731);
xor U25397 (N_25397,N_23694,N_23132);
or U25398 (N_25398,N_23322,N_23469);
nor U25399 (N_25399,N_23196,N_22853);
nor U25400 (N_25400,N_23314,N_22508);
nor U25401 (N_25401,N_23219,N_23624);
nor U25402 (N_25402,N_23013,N_23370);
nor U25403 (N_25403,N_23518,N_22706);
nand U25404 (N_25404,N_23180,N_23952);
xnor U25405 (N_25405,N_22717,N_22897);
nor U25406 (N_25406,N_22882,N_23279);
xor U25407 (N_25407,N_22814,N_23561);
and U25408 (N_25408,N_23899,N_22644);
nor U25409 (N_25409,N_22733,N_23230);
nand U25410 (N_25410,N_23450,N_23022);
xor U25411 (N_25411,N_22651,N_23779);
and U25412 (N_25412,N_22526,N_22877);
nor U25413 (N_25413,N_23352,N_23852);
nand U25414 (N_25414,N_23882,N_23189);
nand U25415 (N_25415,N_23904,N_23825);
and U25416 (N_25416,N_22992,N_23185);
nor U25417 (N_25417,N_23903,N_23006);
xnor U25418 (N_25418,N_23086,N_23399);
and U25419 (N_25419,N_23695,N_23791);
and U25420 (N_25420,N_23133,N_22993);
xnor U25421 (N_25421,N_23044,N_22631);
nor U25422 (N_25422,N_23503,N_23061);
and U25423 (N_25423,N_23288,N_22780);
and U25424 (N_25424,N_23789,N_23331);
or U25425 (N_25425,N_23382,N_23097);
and U25426 (N_25426,N_23843,N_23334);
or U25427 (N_25427,N_23425,N_23463);
nor U25428 (N_25428,N_22825,N_23693);
nand U25429 (N_25429,N_23543,N_23031);
xnor U25430 (N_25430,N_22774,N_22812);
nand U25431 (N_25431,N_23042,N_23260);
xnor U25432 (N_25432,N_23745,N_23952);
xor U25433 (N_25433,N_23034,N_23103);
nor U25434 (N_25434,N_23893,N_23590);
nor U25435 (N_25435,N_23295,N_22753);
nor U25436 (N_25436,N_23408,N_23260);
nor U25437 (N_25437,N_22942,N_23990);
and U25438 (N_25438,N_23748,N_23545);
nand U25439 (N_25439,N_22909,N_22867);
xor U25440 (N_25440,N_22884,N_23272);
xnor U25441 (N_25441,N_22950,N_22884);
and U25442 (N_25442,N_23930,N_23194);
or U25443 (N_25443,N_22940,N_23116);
nand U25444 (N_25444,N_23241,N_23090);
nand U25445 (N_25445,N_23661,N_23249);
or U25446 (N_25446,N_23864,N_23873);
nor U25447 (N_25447,N_22671,N_22614);
nand U25448 (N_25448,N_22826,N_22651);
nor U25449 (N_25449,N_23084,N_22620);
or U25450 (N_25450,N_23723,N_23549);
xnor U25451 (N_25451,N_22935,N_23943);
and U25452 (N_25452,N_22749,N_23516);
or U25453 (N_25453,N_22888,N_23914);
xnor U25454 (N_25454,N_23138,N_23637);
and U25455 (N_25455,N_23407,N_23881);
and U25456 (N_25456,N_23247,N_22737);
nand U25457 (N_25457,N_23576,N_23711);
and U25458 (N_25458,N_22639,N_22637);
xor U25459 (N_25459,N_22548,N_23045);
nor U25460 (N_25460,N_23665,N_22733);
and U25461 (N_25461,N_23042,N_22610);
and U25462 (N_25462,N_23526,N_22629);
xor U25463 (N_25463,N_23476,N_22734);
and U25464 (N_25464,N_23668,N_23370);
and U25465 (N_25465,N_23690,N_23689);
nand U25466 (N_25466,N_23357,N_23246);
and U25467 (N_25467,N_23177,N_23291);
and U25468 (N_25468,N_22954,N_23700);
and U25469 (N_25469,N_23631,N_22778);
xor U25470 (N_25470,N_23197,N_23367);
or U25471 (N_25471,N_22910,N_22817);
or U25472 (N_25472,N_23474,N_23894);
nor U25473 (N_25473,N_23289,N_23563);
xnor U25474 (N_25474,N_22635,N_22604);
nand U25475 (N_25475,N_23261,N_23861);
xor U25476 (N_25476,N_23018,N_23278);
and U25477 (N_25477,N_23106,N_23446);
or U25478 (N_25478,N_23191,N_23033);
nor U25479 (N_25479,N_23276,N_23354);
xnor U25480 (N_25480,N_23078,N_23536);
xnor U25481 (N_25481,N_22957,N_23369);
nor U25482 (N_25482,N_23095,N_23186);
or U25483 (N_25483,N_23389,N_23073);
and U25484 (N_25484,N_23490,N_23731);
nand U25485 (N_25485,N_22863,N_23219);
or U25486 (N_25486,N_23618,N_22945);
xnor U25487 (N_25487,N_23291,N_22946);
or U25488 (N_25488,N_23610,N_22617);
xor U25489 (N_25489,N_23460,N_22807);
nor U25490 (N_25490,N_23280,N_22597);
or U25491 (N_25491,N_23576,N_23984);
nand U25492 (N_25492,N_23567,N_23694);
or U25493 (N_25493,N_23481,N_23100);
or U25494 (N_25494,N_23493,N_23080);
xor U25495 (N_25495,N_23192,N_23252);
and U25496 (N_25496,N_22595,N_23152);
or U25497 (N_25497,N_23492,N_23834);
nor U25498 (N_25498,N_22984,N_23794);
nand U25499 (N_25499,N_23033,N_23530);
xor U25500 (N_25500,N_24083,N_24699);
xnor U25501 (N_25501,N_25205,N_24755);
nand U25502 (N_25502,N_24730,N_24163);
nor U25503 (N_25503,N_24238,N_24891);
and U25504 (N_25504,N_24579,N_25450);
nand U25505 (N_25505,N_24265,N_24071);
xnor U25506 (N_25506,N_24952,N_24229);
nor U25507 (N_25507,N_24501,N_24742);
nor U25508 (N_25508,N_24748,N_24478);
and U25509 (N_25509,N_24523,N_24351);
xnor U25510 (N_25510,N_24459,N_24322);
nand U25511 (N_25511,N_24987,N_24414);
nand U25512 (N_25512,N_24837,N_24195);
or U25513 (N_25513,N_25323,N_25135);
and U25514 (N_25514,N_24946,N_24740);
xnor U25515 (N_25515,N_24108,N_24037);
and U25516 (N_25516,N_24081,N_25038);
nor U25517 (N_25517,N_24209,N_25181);
nand U25518 (N_25518,N_25453,N_24471);
nor U25519 (N_25519,N_24529,N_24665);
or U25520 (N_25520,N_25271,N_24403);
nor U25521 (N_25521,N_24479,N_24863);
xor U25522 (N_25522,N_24741,N_25253);
xor U25523 (N_25523,N_24261,N_24972);
xnor U25524 (N_25524,N_24399,N_24527);
or U25525 (N_25525,N_24213,N_25367);
or U25526 (N_25526,N_24556,N_24519);
and U25527 (N_25527,N_25020,N_24206);
nand U25528 (N_25528,N_24067,N_24207);
and U25529 (N_25529,N_25082,N_25345);
nand U25530 (N_25530,N_24744,N_24180);
and U25531 (N_25531,N_24375,N_24049);
xor U25532 (N_25532,N_24227,N_25073);
nand U25533 (N_25533,N_24088,N_24043);
xor U25534 (N_25534,N_24161,N_24805);
nor U25535 (N_25535,N_24457,N_25241);
and U25536 (N_25536,N_25454,N_24600);
and U25537 (N_25537,N_25190,N_24378);
or U25538 (N_25538,N_24691,N_24650);
or U25539 (N_25539,N_25342,N_24311);
xnor U25540 (N_25540,N_24924,N_25457);
or U25541 (N_25541,N_24709,N_24361);
nand U25542 (N_25542,N_24566,N_24135);
or U25543 (N_25543,N_24706,N_25145);
xor U25544 (N_25544,N_24446,N_24063);
nor U25545 (N_25545,N_25121,N_25123);
nand U25546 (N_25546,N_24156,N_24644);
and U25547 (N_25547,N_24336,N_25156);
or U25548 (N_25548,N_24241,N_24096);
nand U25549 (N_25549,N_24027,N_24050);
or U25550 (N_25550,N_24326,N_25305);
xnor U25551 (N_25551,N_24452,N_24392);
and U25552 (N_25552,N_24642,N_24723);
xnor U25553 (N_25553,N_25136,N_24567);
or U25554 (N_25554,N_25297,N_25062);
xor U25555 (N_25555,N_24331,N_25105);
or U25556 (N_25556,N_25255,N_24362);
xor U25557 (N_25557,N_24258,N_24493);
nor U25558 (N_25558,N_24211,N_24692);
nand U25559 (N_25559,N_24761,N_24445);
nor U25560 (N_25560,N_25442,N_25462);
nand U25561 (N_25561,N_24455,N_24500);
nand U25562 (N_25562,N_24118,N_25460);
nand U25563 (N_25563,N_25226,N_24803);
xor U25564 (N_25564,N_24450,N_25258);
xnor U25565 (N_25565,N_25292,N_24386);
nand U25566 (N_25566,N_24492,N_24041);
xnor U25567 (N_25567,N_24094,N_24400);
and U25568 (N_25568,N_24340,N_24460);
nand U25569 (N_25569,N_24697,N_24150);
nand U25570 (N_25570,N_25419,N_24530);
and U25571 (N_25571,N_24465,N_24447);
or U25572 (N_25572,N_25482,N_24107);
and U25573 (N_25573,N_24698,N_24965);
or U25574 (N_25574,N_24069,N_24239);
or U25575 (N_25575,N_24578,N_24806);
or U25576 (N_25576,N_25393,N_25054);
nor U25577 (N_25577,N_24836,N_25083);
and U25578 (N_25578,N_25163,N_25494);
nor U25579 (N_25579,N_24275,N_24616);
and U25580 (N_25580,N_24320,N_24487);
and U25581 (N_25581,N_24055,N_24352);
or U25582 (N_25582,N_25473,N_24504);
nand U25583 (N_25583,N_25228,N_25227);
and U25584 (N_25584,N_25458,N_24330);
or U25585 (N_25585,N_24164,N_24750);
nor U25586 (N_25586,N_25491,N_24090);
nand U25587 (N_25587,N_24700,N_24169);
xor U25588 (N_25588,N_24569,N_25027);
xnor U25589 (N_25589,N_24285,N_25065);
xor U25590 (N_25590,N_24598,N_24084);
and U25591 (N_25591,N_25213,N_24917);
nand U25592 (N_25592,N_25488,N_24677);
nand U25593 (N_25593,N_24724,N_25268);
xor U25594 (N_25594,N_24483,N_24068);
and U25595 (N_25595,N_24981,N_24571);
xor U25596 (N_25596,N_24266,N_24781);
or U25597 (N_25597,N_24589,N_24097);
and U25598 (N_25598,N_25189,N_24271);
nand U25599 (N_25599,N_25372,N_24606);
nor U25600 (N_25600,N_24839,N_24797);
or U25601 (N_25601,N_24407,N_24299);
or U25602 (N_25602,N_25196,N_24536);
nand U25603 (N_25603,N_24018,N_24484);
nand U25604 (N_25604,N_25273,N_24248);
or U25605 (N_25605,N_24601,N_25310);
and U25606 (N_25606,N_24053,N_24890);
nand U25607 (N_25607,N_25395,N_25006);
nor U25608 (N_25608,N_24105,N_25120);
nand U25609 (N_25609,N_25328,N_24634);
nand U25610 (N_25610,N_24720,N_24327);
nor U25611 (N_25611,N_24651,N_25053);
or U25612 (N_25612,N_24413,N_25324);
nor U25613 (N_25613,N_24418,N_24905);
and U25614 (N_25614,N_25425,N_25366);
or U25615 (N_25615,N_25118,N_24898);
nand U25616 (N_25616,N_24522,N_24762);
xnor U25617 (N_25617,N_25103,N_25363);
xnor U25618 (N_25618,N_24660,N_24872);
nand U25619 (N_25619,N_25111,N_25249);
nand U25620 (N_25620,N_24707,N_24387);
xnor U25621 (N_25621,N_24035,N_24807);
and U25622 (N_25622,N_24737,N_24818);
and U25623 (N_25623,N_24974,N_25362);
xor U25624 (N_25624,N_25252,N_24103);
or U25625 (N_25625,N_25451,N_24678);
and U25626 (N_25626,N_24732,N_24743);
nand U25627 (N_25627,N_24372,N_24419);
and U25628 (N_25628,N_24931,N_24325);
or U25629 (N_25629,N_24555,N_24516);
xor U25630 (N_25630,N_24810,N_24782);
nor U25631 (N_25631,N_24428,N_25140);
nand U25632 (N_25632,N_24437,N_24553);
or U25633 (N_25633,N_24186,N_24683);
nand U25634 (N_25634,N_25339,N_24996);
xor U25635 (N_25635,N_24199,N_25476);
and U25636 (N_25636,N_24177,N_25160);
and U25637 (N_25637,N_24901,N_25202);
nor U25638 (N_25638,N_24409,N_25315);
and U25639 (N_25639,N_24545,N_25229);
xnor U25640 (N_25640,N_24052,N_25282);
or U25641 (N_25641,N_24552,N_25427);
or U25642 (N_25642,N_24429,N_25321);
nand U25643 (N_25643,N_24039,N_25257);
xor U25644 (N_25644,N_24194,N_25404);
and U25645 (N_25645,N_25192,N_25433);
xnor U25646 (N_25646,N_25167,N_24726);
nand U25647 (N_25647,N_24800,N_25304);
xor U25648 (N_25648,N_24232,N_24592);
xnor U25649 (N_25649,N_24219,N_25264);
and U25650 (N_25650,N_25398,N_24851);
nand U25651 (N_25651,N_24764,N_24821);
nor U25652 (N_25652,N_24597,N_25408);
or U25653 (N_25653,N_25231,N_24915);
nand U25654 (N_25654,N_24703,N_24846);
xnor U25655 (N_25655,N_24612,N_24621);
xor U25656 (N_25656,N_25267,N_25432);
or U25657 (N_25657,N_25183,N_25005);
nand U25658 (N_25658,N_25104,N_24481);
nand U25659 (N_25659,N_24937,N_25341);
or U25660 (N_25660,N_24510,N_24899);
and U25661 (N_25661,N_24801,N_25025);
nor U25662 (N_25662,N_25349,N_25287);
or U25663 (N_25663,N_25336,N_24142);
xor U25664 (N_25664,N_24633,N_25001);
or U25665 (N_25665,N_24879,N_24645);
xnor U25666 (N_25666,N_24104,N_25221);
or U25667 (N_25667,N_25012,N_24319);
nor U25668 (N_25668,N_24300,N_24792);
nor U25669 (N_25669,N_25275,N_24431);
xor U25670 (N_25670,N_24815,N_24283);
xor U25671 (N_25671,N_24985,N_25477);
xnor U25672 (N_25672,N_24903,N_24860);
or U25673 (N_25673,N_24246,N_25334);
nor U25674 (N_25674,N_25331,N_24923);
or U25675 (N_25675,N_24512,N_24282);
and U25676 (N_25676,N_25391,N_24046);
xnor U25677 (N_25677,N_24524,N_25172);
nor U25678 (N_25678,N_25217,N_25385);
and U25679 (N_25679,N_24005,N_25098);
or U25680 (N_25680,N_25470,N_24630);
or U25681 (N_25681,N_24448,N_24121);
xor U25682 (N_25682,N_24247,N_25165);
nor U25683 (N_25683,N_24943,N_24395);
or U25684 (N_25684,N_24874,N_24377);
nor U25685 (N_25685,N_25444,N_24091);
and U25686 (N_25686,N_25070,N_25148);
and U25687 (N_25687,N_24405,N_24042);
or U25688 (N_25688,N_24876,N_25000);
or U25689 (N_25689,N_24205,N_24930);
or U25690 (N_25690,N_25466,N_24973);
or U25691 (N_25691,N_24058,N_24131);
xor U25692 (N_25692,N_25194,N_24988);
xnor U25693 (N_25693,N_25492,N_25302);
xor U25694 (N_25694,N_25050,N_25371);
nor U25695 (N_25695,N_24780,N_24065);
and U25696 (N_25696,N_24430,N_24040);
nand U25697 (N_25697,N_25233,N_24031);
xnor U25698 (N_25698,N_25319,N_24296);
xor U25699 (N_25699,N_24680,N_24820);
or U25700 (N_25700,N_24619,N_25277);
xnor U25701 (N_25701,N_25344,N_24226);
nand U25702 (N_25702,N_24017,N_24470);
xnor U25703 (N_25703,N_25019,N_24986);
or U25704 (N_25704,N_24558,N_24926);
nor U25705 (N_25705,N_25298,N_25312);
nor U25706 (N_25706,N_24751,N_24662);
and U25707 (N_25707,N_24286,N_24659);
and U25708 (N_25708,N_25177,N_25060);
nand U25709 (N_25709,N_25224,N_24664);
nor U25710 (N_25710,N_24568,N_25126);
nand U25711 (N_25711,N_24280,N_25033);
or U25712 (N_25712,N_24440,N_24365);
or U25713 (N_25713,N_24577,N_24812);
or U25714 (N_25714,N_24904,N_24363);
xor U25715 (N_25715,N_25346,N_25097);
and U25716 (N_25716,N_25379,N_25072);
nand U25717 (N_25717,N_25130,N_24835);
and U25718 (N_25718,N_25011,N_25184);
nor U25719 (N_25719,N_24026,N_24747);
and U25720 (N_25720,N_24292,N_24441);
or U25721 (N_25721,N_24914,N_24396);
and U25722 (N_25722,N_24626,N_24822);
xnor U25723 (N_25723,N_24305,N_24770);
or U25724 (N_25724,N_24845,N_25320);
nor U25725 (N_25725,N_25499,N_25317);
nor U25726 (N_25726,N_25447,N_24971);
or U25727 (N_25727,N_25124,N_24938);
nand U25728 (N_25728,N_25422,N_24402);
or U25729 (N_25729,N_24294,N_25159);
nor U25730 (N_25730,N_24162,N_24954);
or U25731 (N_25731,N_24323,N_24989);
nand U25732 (N_25732,N_25057,N_25311);
or U25733 (N_25733,N_25101,N_24346);
or U25734 (N_25734,N_24334,N_24604);
xnor U25735 (N_25735,N_24314,N_24394);
nor U25736 (N_25736,N_24153,N_24383);
xnor U25737 (N_25737,N_25359,N_25368);
or U25738 (N_25738,N_24370,N_24853);
or U25739 (N_25739,N_24649,N_25479);
nor U25740 (N_25740,N_24913,N_25112);
and U25741 (N_25741,N_24992,N_24540);
nor U25742 (N_25742,N_25230,N_24588);
or U25743 (N_25743,N_24980,N_24712);
xor U25744 (N_25744,N_25348,N_24875);
xor U25745 (N_25745,N_24798,N_24663);
or U25746 (N_25746,N_24843,N_24841);
or U25747 (N_25747,N_24288,N_25200);
and U25748 (N_25748,N_24324,N_24412);
nor U25749 (N_25749,N_24811,N_24969);
or U25750 (N_25750,N_24574,N_25399);
or U25751 (N_25751,N_24379,N_24714);
nand U25752 (N_25752,N_24968,N_25193);
nand U25753 (N_25753,N_24886,N_25037);
and U25754 (N_25754,N_24201,N_24696);
nand U25755 (N_25755,N_25007,N_25113);
xor U25756 (N_25756,N_24033,N_24725);
nand U25757 (N_25757,N_24823,N_24754);
nor U25758 (N_25758,N_25219,N_24273);
nand U25759 (N_25759,N_24611,N_24263);
and U25760 (N_25760,N_25276,N_25131);
nand U25761 (N_25761,N_24038,N_24353);
xnor U25762 (N_25762,N_24185,N_25467);
or U25763 (N_25763,N_24244,N_25188);
or U25764 (N_25764,N_25443,N_24496);
and U25765 (N_25765,N_25360,N_25474);
nor U25766 (N_25766,N_24878,N_25023);
or U25767 (N_25767,N_24842,N_25223);
or U25768 (N_25768,N_24715,N_24546);
xor U25769 (N_25769,N_25141,N_25114);
nand U25770 (N_25770,N_24561,N_24434);
xor U25771 (N_25771,N_24307,N_24264);
xor U25772 (N_25772,N_25309,N_24997);
xnor U25773 (N_25773,N_25409,N_24358);
nand U25774 (N_25774,N_24464,N_24652);
and U25775 (N_25775,N_24735,N_25370);
xnor U25776 (N_25776,N_24242,N_24117);
nand U25777 (N_25777,N_24149,N_24354);
xnor U25778 (N_25778,N_24147,N_25220);
xor U25779 (N_25779,N_24250,N_25441);
or U25780 (N_25780,N_24559,N_24062);
nor U25781 (N_25781,N_24749,N_24667);
or U25782 (N_25782,N_25388,N_25461);
nor U25783 (N_25783,N_24738,N_25495);
and U25784 (N_25784,N_25102,N_24298);
and U25785 (N_25785,N_24635,N_24548);
and U25786 (N_25786,N_24858,N_24137);
or U25787 (N_25787,N_24710,N_24290);
or U25788 (N_25788,N_24245,N_24277);
xor U25789 (N_25789,N_25475,N_24593);
and U25790 (N_25790,N_25410,N_24256);
nor U25791 (N_25791,N_24936,N_24584);
nor U25792 (N_25792,N_25353,N_24349);
xor U25793 (N_25793,N_25178,N_25058);
or U25794 (N_25794,N_25150,N_24356);
nand U25795 (N_25795,N_25356,N_24002);
nand U25796 (N_25796,N_24883,N_24927);
xor U25797 (N_25797,N_25081,N_24894);
and U25798 (N_25798,N_24560,N_24140);
xnor U25799 (N_25799,N_24773,N_24767);
or U25800 (N_25800,N_25326,N_24861);
nand U25801 (N_25801,N_24838,N_24393);
nor U25802 (N_25802,N_25246,N_24585);
or U25803 (N_25803,N_25248,N_24032);
xnor U25804 (N_25804,N_25280,N_25208);
xor U25805 (N_25805,N_25047,N_25168);
and U25806 (N_25806,N_24507,N_24006);
and U25807 (N_25807,N_24774,N_25293);
nand U25808 (N_25808,N_24557,N_25179);
nand U25809 (N_25809,N_24231,N_24688);
xor U25810 (N_25810,N_24882,N_24908);
nor U25811 (N_25811,N_24126,N_24857);
or U25812 (N_25812,N_25009,N_24073);
nand U25813 (N_25813,N_24979,N_25024);
nor U25814 (N_25814,N_25236,N_25066);
xnor U25815 (N_25815,N_24884,N_24112);
nand U25816 (N_25816,N_24200,N_25465);
nand U25817 (N_25817,N_24581,N_24854);
or U25818 (N_25818,N_24935,N_24036);
and U25819 (N_25819,N_24243,N_24912);
nand U25820 (N_25820,N_25376,N_24255);
and U25821 (N_25821,N_24813,N_24144);
nor U25822 (N_25822,N_24109,N_25064);
or U25823 (N_25823,N_24061,N_24456);
nor U25824 (N_25824,N_25086,N_24364);
or U25825 (N_25825,N_25459,N_25307);
nand U25826 (N_25826,N_24054,N_24515);
nand U25827 (N_25827,N_25191,N_25242);
or U25828 (N_25828,N_24538,N_24982);
and U25829 (N_25829,N_24176,N_24834);
or U25830 (N_25830,N_25373,N_24490);
nor U25831 (N_25831,N_25127,N_25288);
and U25832 (N_25832,N_24763,N_24454);
or U25833 (N_25833,N_25115,N_24066);
xnor U25834 (N_25834,N_24423,N_24350);
and U25835 (N_25835,N_24308,N_24933);
nand U25836 (N_25836,N_24825,N_25034);
xnor U25837 (N_25837,N_25182,N_24388);
nor U25838 (N_25838,N_24814,N_25496);
or U25839 (N_25839,N_24315,N_25284);
xor U25840 (N_25840,N_24681,N_24718);
xnor U25841 (N_25841,N_24525,N_25158);
nor U25842 (N_25842,N_24535,N_24020);
and U25843 (N_25843,N_24833,N_25424);
nor U25844 (N_25844,N_24449,N_24444);
and U25845 (N_25845,N_24721,N_25416);
xor U25846 (N_25846,N_24141,N_24092);
nand U25847 (N_25847,N_25418,N_24847);
nor U25848 (N_25848,N_24095,N_24008);
or U25849 (N_25849,N_25122,N_25303);
or U25850 (N_25850,N_24316,N_24087);
and U25851 (N_25851,N_24178,N_25269);
nand U25852 (N_25852,N_24304,N_24328);
nand U25853 (N_25853,N_24840,N_24240);
or U25854 (N_25854,N_25008,N_24949);
and U25855 (N_25855,N_24376,N_24306);
nor U25856 (N_25856,N_24279,N_24003);
or U25857 (N_25857,N_24406,N_24499);
nor U25858 (N_25858,N_24295,N_25212);
or U25859 (N_25859,N_25274,N_24978);
and U25860 (N_25860,N_25116,N_25110);
nand U25861 (N_25861,N_24016,N_24809);
nand U25862 (N_25862,N_24785,N_24671);
and U25863 (N_25863,N_25014,N_24110);
nor U25864 (N_25864,N_24397,N_24249);
or U25865 (N_25865,N_25243,N_24371);
nand U25866 (N_25866,N_24543,N_24733);
or U25867 (N_25867,N_25092,N_25489);
nand U25868 (N_25868,N_25405,N_24015);
nand U25869 (N_25869,N_24260,N_24958);
xnor U25870 (N_25870,N_24472,N_24717);
or U25871 (N_25871,N_24582,N_24534);
nand U25872 (N_25872,N_24064,N_24369);
nor U25873 (N_25873,N_25089,N_24966);
and U25874 (N_25874,N_24831,N_24181);
and U25875 (N_25875,N_24918,N_24716);
and U25876 (N_25876,N_24676,N_24477);
xnor U25877 (N_25877,N_24786,N_24480);
nand U25878 (N_25878,N_25109,N_24237);
xnor U25879 (N_25879,N_24998,N_24702);
xnor U25880 (N_25880,N_24640,N_25365);
xor U25881 (N_25881,N_24114,N_25031);
xor U25882 (N_25882,N_24768,N_25045);
nor U25883 (N_25883,N_24673,N_24228);
or U25884 (N_25884,N_24059,N_24906);
or U25885 (N_25885,N_24120,N_24101);
nor U25886 (N_25886,N_25361,N_24160);
or U25887 (N_25887,N_25308,N_24432);
nor U25888 (N_25888,N_25445,N_24159);
xnor U25889 (N_25889,N_24942,N_24870);
nand U25890 (N_25890,N_25335,N_25439);
or U25891 (N_25891,N_24485,N_24007);
or U25892 (N_25892,N_24495,N_24230);
and U25893 (N_25893,N_25080,N_25322);
or U25894 (N_25894,N_24367,N_25375);
or U25895 (N_25895,N_24647,N_24654);
or U25896 (N_25896,N_24505,N_24796);
or U25897 (N_25897,N_24010,N_24617);
nor U25898 (N_25898,N_25210,N_24580);
and U25899 (N_25899,N_24922,N_25497);
xnor U25900 (N_25900,N_24850,N_24877);
nand U25901 (N_25901,N_25093,N_24832);
xnor U25902 (N_25902,N_24517,N_25134);
xor U25903 (N_25903,N_25046,N_25382);
xor U25904 (N_25904,N_24408,N_25199);
or U25905 (N_25905,N_24045,N_24089);
xnor U25906 (N_25906,N_25107,N_24024);
nor U25907 (N_25907,N_25314,N_24541);
and U25908 (N_25908,N_24636,N_25330);
and U25909 (N_25909,N_24234,N_25383);
or U25910 (N_25910,N_25266,N_25117);
and U25911 (N_25911,N_24424,N_24900);
nor U25912 (N_25912,N_24453,N_24928);
and U25913 (N_25913,N_24728,N_24210);
nor U25914 (N_25914,N_24047,N_24236);
nor U25915 (N_25915,N_25487,N_25449);
nor U25916 (N_25916,N_24920,N_24547);
xnor U25917 (N_25917,N_25187,N_24675);
nand U25918 (N_25918,N_24272,N_24284);
nand U25919 (N_25919,N_24518,N_24888);
or U25920 (N_25920,N_24102,N_24520);
xnor U25921 (N_25921,N_24766,N_24991);
or U25922 (N_25922,N_25251,N_25206);
nand U25923 (N_25923,N_25438,N_24791);
nand U25924 (N_25924,N_24215,N_25095);
nor U25925 (N_25925,N_24187,N_24021);
nor U25926 (N_25926,N_24214,N_25214);
nand U25927 (N_25927,N_24175,N_25392);
or U25928 (N_25928,N_24293,N_24804);
nand U25929 (N_25929,N_25333,N_24939);
nor U25930 (N_25930,N_24948,N_25401);
or U25931 (N_25931,N_24777,N_24193);
or U25932 (N_25932,N_24701,N_25316);
nand U25933 (N_25933,N_24357,N_24070);
xnor U25934 (N_25934,N_24208,N_24669);
or U25935 (N_25935,N_25042,N_24648);
xor U25936 (N_25936,N_24222,N_24224);
nand U25937 (N_25937,N_24956,N_24827);
and U25938 (N_25938,N_24544,N_24503);
and U25939 (N_25939,N_24416,N_25068);
xor U25940 (N_25940,N_24990,N_24333);
nand U25941 (N_25941,N_25256,N_24380);
or U25942 (N_25942,N_24329,N_24360);
nor U25943 (N_25943,N_24573,N_25094);
nand U25944 (N_25944,N_24550,N_24190);
or U25945 (N_25945,N_24653,N_24173);
nand U25946 (N_25946,N_24301,N_25318);
xnor U25947 (N_25947,N_24950,N_25380);
xnor U25948 (N_25948,N_25225,N_25394);
xnor U25949 (N_25949,N_24607,N_24257);
and U25950 (N_25950,N_24591,N_25436);
or U25951 (N_25951,N_24599,N_24960);
or U25952 (N_25952,N_25381,N_25142);
nor U25953 (N_25953,N_24947,N_24753);
xor U25954 (N_25954,N_24184,N_24482);
xor U25955 (N_25955,N_25018,N_24022);
nand U25956 (N_25956,N_24586,N_24911);
nor U25957 (N_25957,N_24034,N_24984);
nand U25958 (N_25958,N_24051,N_24204);
nor U25959 (N_25959,N_25203,N_24303);
and U25960 (N_25960,N_25010,N_24784);
xor U25961 (N_25961,N_25435,N_25234);
nor U25962 (N_25962,N_24174,N_24494);
nand U25963 (N_25963,N_24562,N_24614);
nor U25964 (N_25964,N_25239,N_24892);
nor U25965 (N_25965,N_25270,N_25036);
or U25966 (N_25966,N_24844,N_24613);
xnor U25967 (N_25967,N_24687,N_24044);
nor U25968 (N_25968,N_24521,N_24401);
and U25969 (N_25969,N_25201,N_24463);
nor U25970 (N_25970,N_24790,N_24759);
nand U25971 (N_25971,N_24713,N_25291);
or U25972 (N_25972,N_25468,N_24216);
or U25973 (N_25973,N_25285,N_25162);
nor U25974 (N_25974,N_25283,N_24443);
nor U25975 (N_25975,N_24233,N_25071);
nand U25976 (N_25976,N_24916,N_24461);
or U25977 (N_25977,N_24011,N_24977);
nor U25978 (N_25978,N_25481,N_24919);
or U25979 (N_25979,N_25166,N_25055);
or U25980 (N_25980,N_24398,N_25149);
nand U25981 (N_25981,N_24502,N_24620);
nand U25982 (N_25982,N_25232,N_25133);
or U25983 (N_25983,N_24695,N_24218);
and U25984 (N_25984,N_24077,N_24615);
nand U25985 (N_25985,N_24605,N_25456);
or U25986 (N_25986,N_25056,N_24475);
xor U25987 (N_25987,N_24253,N_25138);
nand U25988 (N_25988,N_24945,N_25247);
or U25989 (N_25989,N_24631,N_24570);
xor U25990 (N_25990,N_25088,N_24632);
nor U25991 (N_25991,N_24993,N_24139);
nand U25992 (N_25992,N_24909,N_25369);
nand U25993 (N_25993,N_24955,N_24417);
and U25994 (N_25994,N_24188,N_24385);
and U25995 (N_25995,N_24953,N_25125);
nand U25996 (N_25996,N_24995,N_24563);
and U25997 (N_25997,N_24148,N_25087);
nor U25998 (N_25998,N_25396,N_25452);
nor U25999 (N_25999,N_24123,N_25143);
or U26000 (N_26000,N_24335,N_25407);
and U26001 (N_26001,N_25137,N_24321);
nand U26002 (N_26002,N_24030,N_24929);
nor U26003 (N_26003,N_24771,N_25079);
nor U26004 (N_26004,N_25096,N_24212);
nor U26005 (N_26005,N_25169,N_24468);
nor U26006 (N_26006,N_24341,N_25176);
or U26007 (N_26007,N_24276,N_25286);
or U26008 (N_26008,N_24235,N_24896);
and U26009 (N_26009,N_25157,N_25483);
nor U26010 (N_26010,N_24668,N_24093);
or U26011 (N_26011,N_24381,N_24289);
nor U26012 (N_26012,N_25170,N_24309);
and U26013 (N_26013,N_24004,N_25250);
xor U26014 (N_26014,N_24136,N_24347);
and U26015 (N_26015,N_25197,N_24439);
nand U26016 (N_26016,N_25099,N_24013);
nand U26017 (N_26017,N_25440,N_24157);
xnor U26018 (N_26018,N_24679,N_25175);
nand U26019 (N_26019,N_24532,N_24138);
nand U26020 (N_26020,N_24154,N_24146);
and U26021 (N_26021,N_24012,N_24817);
or U26022 (N_26022,N_25430,N_24368);
xnor U26023 (N_26023,N_24684,N_25090);
nand U26024 (N_26024,N_24921,N_24506);
nor U26025 (N_26025,N_24115,N_25464);
and U26026 (N_26026,N_24694,N_25329);
or U26027 (N_26027,N_24191,N_25244);
nor U26028 (N_26028,N_24602,N_24745);
nand U26029 (N_26029,N_24610,N_24145);
or U26030 (N_26030,N_25044,N_25076);
nand U26031 (N_26031,N_24192,N_25455);
and U26032 (N_26032,N_24511,N_25364);
nand U26033 (N_26033,N_24783,N_24513);
and U26034 (N_26034,N_24072,N_24098);
and U26035 (N_26035,N_24436,N_24317);
xnor U26036 (N_26036,N_24488,N_24348);
nand U26037 (N_26037,N_24152,N_24658);
nor U26038 (N_26038,N_24217,N_24787);
nand U26039 (N_26039,N_24869,N_24171);
nor U26040 (N_26040,N_25198,N_25313);
or U26041 (N_26041,N_24458,N_24902);
nor U26042 (N_26042,N_25043,N_24539);
xor U26043 (N_26043,N_25003,N_25352);
nor U26044 (N_26044,N_25245,N_25414);
nor U26045 (N_26045,N_24338,N_24421);
and U26046 (N_26046,N_24462,N_25423);
or U26047 (N_26047,N_25147,N_24125);
nor U26048 (N_26048,N_25144,N_24172);
nor U26049 (N_26049,N_24183,N_25139);
nand U26050 (N_26050,N_25486,N_24128);
nor U26051 (N_26051,N_24772,N_24789);
nor U26052 (N_26052,N_24343,N_24583);
and U26053 (N_26053,N_24198,N_25263);
nor U26054 (N_26054,N_24885,N_24389);
and U26055 (N_26055,N_25084,N_24816);
xor U26056 (N_26056,N_24332,N_24451);
nand U26057 (N_26057,N_25161,N_25069);
and U26058 (N_26058,N_25480,N_25209);
nor U26059 (N_26059,N_24442,N_25237);
nor U26060 (N_26060,N_24666,N_24639);
xnor U26061 (N_26061,N_24862,N_24438);
xnor U26062 (N_26062,N_24078,N_25406);
nand U26063 (N_26063,N_24491,N_24951);
nand U26064 (N_26064,N_24151,N_25420);
nor U26065 (N_26065,N_25185,N_24819);
nand U26066 (N_26066,N_24656,N_24704);
xor U26067 (N_26067,N_25289,N_24690);
and U26068 (N_26068,N_25049,N_24057);
nor U26069 (N_26069,N_25343,N_25485);
nand U26070 (N_26070,N_25278,N_24856);
xor U26071 (N_26071,N_24025,N_25294);
nand U26072 (N_26072,N_24124,N_24934);
or U26073 (N_26073,N_24983,N_25254);
and U26074 (N_26074,N_25281,N_24624);
or U26075 (N_26075,N_25164,N_25195);
nor U26076 (N_26076,N_25351,N_24080);
nand U26077 (N_26077,N_24337,N_24291);
nand U26078 (N_26078,N_24056,N_24608);
and U26079 (N_26079,N_24278,N_25048);
nor U26080 (N_26080,N_25015,N_24776);
nand U26081 (N_26081,N_25355,N_24655);
nor U26082 (N_26082,N_25028,N_24179);
nand U26083 (N_26083,N_24893,N_24719);
nor U26084 (N_26084,N_24100,N_25129);
nand U26085 (N_26085,N_24533,N_25059);
nor U26086 (N_26086,N_24734,N_25354);
nand U26087 (N_26087,N_25207,N_25063);
or U26088 (N_26088,N_24779,N_25215);
xnor U26089 (N_26089,N_24359,N_24384);
nand U26090 (N_26090,N_25421,N_24168);
and U26091 (N_26091,N_24476,N_25358);
and U26092 (N_26092,N_25490,N_25347);
nor U26093 (N_26093,N_24760,N_24082);
and U26094 (N_26094,N_25067,N_24079);
and U26095 (N_26095,N_24202,N_25106);
nor U26096 (N_26096,N_24752,N_24964);
nand U26097 (N_26097,N_24603,N_25146);
xor U26098 (N_26098,N_25016,N_25377);
and U26099 (N_26099,N_24674,N_24404);
nand U26100 (N_26100,N_25128,N_24318);
and U26101 (N_26101,N_24940,N_24134);
and U26102 (N_26102,N_24824,N_24758);
and U26103 (N_26103,N_24765,N_25415);
nor U26104 (N_26104,N_24203,N_25428);
or U26105 (N_26105,N_24587,N_25074);
nand U26106 (N_26106,N_24287,N_24514);
nand U26107 (N_26107,N_25426,N_24970);
or U26108 (N_26108,N_24312,N_24994);
xor U26109 (N_26109,N_24269,N_24672);
nor U26110 (N_26110,N_24474,N_24623);
or U26111 (N_26111,N_24722,N_24143);
nand U26112 (N_26112,N_25032,N_24618);
or U26113 (N_26113,N_25261,N_24076);
or U26114 (N_26114,N_24411,N_24575);
nor U26115 (N_26115,N_25327,N_25030);
nor U26116 (N_26116,N_24155,N_24802);
nor U26117 (N_26117,N_24382,N_25389);
and U26118 (N_26118,N_24641,N_25040);
xnor U26119 (N_26119,N_25350,N_24873);
and U26120 (N_26120,N_24963,N_24373);
nor U26121 (N_26121,N_25337,N_25417);
and U26122 (N_26122,N_24910,N_25472);
nor U26123 (N_26123,N_24526,N_24009);
and U26124 (N_26124,N_24967,N_24158);
or U26125 (N_26125,N_25021,N_24473);
nor U26126 (N_26126,N_24711,N_24111);
nor U26127 (N_26127,N_25029,N_24793);
nand U26128 (N_26128,N_24795,N_25386);
nor U26129 (N_26129,N_25387,N_25338);
xnor U26130 (N_26130,N_24975,N_24390);
nor U26131 (N_26131,N_25265,N_24374);
or U26132 (N_26132,N_25357,N_25153);
nor U26133 (N_26133,N_24881,N_24961);
or U26134 (N_26134,N_24689,N_25400);
xor U26135 (N_26135,N_24957,N_25119);
or U26136 (N_26136,N_24182,N_24422);
nand U26137 (N_26137,N_24859,N_24262);
xnor U26138 (N_26138,N_24576,N_25211);
or U26139 (N_26139,N_24661,N_24014);
and U26140 (N_26140,N_25173,N_25378);
or U26141 (N_26141,N_24941,N_25411);
nor U26142 (N_26142,N_24867,N_24622);
xor U26143 (N_26143,N_24225,N_25051);
xor U26144 (N_26144,N_25204,N_24756);
nand U26145 (N_26145,N_24799,N_25402);
nor U26146 (N_26146,N_24628,N_24705);
or U26147 (N_26147,N_24999,N_24627);
xor U26148 (N_26148,N_24252,N_24196);
nor U26149 (N_26149,N_25446,N_24739);
or U26150 (N_26150,N_25171,N_24849);
xor U26151 (N_26151,N_24537,N_24119);
xnor U26152 (N_26152,N_24757,N_24420);
or U26153 (N_26153,N_24729,N_24609);
or U26154 (N_26154,N_24489,N_24880);
nor U26155 (N_26155,N_24682,N_25085);
or U26156 (N_26156,N_25384,N_25240);
or U26157 (N_26157,N_24746,N_24197);
and U26158 (N_26158,N_24727,N_24976);
xor U26159 (N_26159,N_24638,N_24251);
and U26160 (N_26160,N_24132,N_25013);
and U26161 (N_26161,N_24085,N_24427);
nand U26162 (N_26162,N_25478,N_25108);
and U26163 (N_26163,N_24433,N_24564);
nand U26164 (N_26164,N_25295,N_25152);
or U26165 (N_26165,N_24466,N_24129);
xnor U26166 (N_26166,N_24415,N_24528);
nor U26167 (N_26167,N_25272,N_24932);
and U26168 (N_26168,N_25431,N_24855);
nand U26169 (N_26169,N_25035,N_24270);
and U26170 (N_26170,N_24469,N_25180);
and U26171 (N_26171,N_25151,N_24133);
xnor U26172 (N_26172,N_24596,N_25279);
xor U26173 (N_26173,N_25077,N_24345);
nand U26174 (N_26174,N_25300,N_24113);
nor U26175 (N_26175,N_24028,N_24775);
and U26176 (N_26176,N_24788,N_24259);
or U26177 (N_26177,N_24708,N_24852);
nand U26178 (N_26178,N_24267,N_24830);
and U26179 (N_26179,N_25259,N_25100);
nand U26180 (N_26180,N_24731,N_25429);
and U26181 (N_26181,N_24542,N_24274);
and U26182 (N_26182,N_24075,N_24625);
nand U26183 (N_26183,N_25469,N_24355);
nor U26184 (N_26184,N_24572,N_24590);
nand U26185 (N_26185,N_24736,N_25002);
and U26186 (N_26186,N_24106,N_24116);
or U26187 (N_26187,N_24907,N_24944);
xnor U26188 (N_26188,N_24167,N_24829);
nor U26189 (N_26189,N_24344,N_25403);
xnor U26190 (N_26190,N_24865,N_24048);
and U26191 (N_26191,N_25325,N_24099);
nand U26192 (N_26192,N_24670,N_24122);
nand U26193 (N_26193,N_25238,N_24467);
and U26194 (N_26194,N_24594,N_24887);
or U26195 (N_26195,N_24508,N_24029);
nand U26196 (N_26196,N_25075,N_24268);
xor U26197 (N_26197,N_24866,N_24629);
nor U26198 (N_26198,N_24127,N_25004);
and U26199 (N_26199,N_24693,N_25299);
nor U26200 (N_26200,N_25306,N_25413);
xor U26201 (N_26201,N_25434,N_24166);
nand U26202 (N_26202,N_24685,N_25026);
and U26203 (N_26203,N_24646,N_24828);
nor U26204 (N_26204,N_24897,N_25290);
nor U26205 (N_26205,N_24808,N_25186);
or U26206 (N_26206,N_25296,N_24871);
or U26207 (N_26207,N_24643,N_24220);
nor U26208 (N_26208,N_24000,N_24657);
xor U26209 (N_26209,N_24130,N_25222);
and U26210 (N_26210,N_24551,N_25017);
nand U26211 (N_26211,N_24595,N_25091);
xor U26212 (N_26212,N_25390,N_25260);
and U26213 (N_26213,N_24864,N_24281);
nand U26214 (N_26214,N_25216,N_24794);
nand U26215 (N_26215,N_24848,N_24410);
or U26216 (N_26216,N_24425,N_24223);
nor U26217 (N_26217,N_24426,N_24165);
xnor U26218 (N_26218,N_25374,N_24019);
xnor U26219 (N_26219,N_24060,N_25498);
nor U26220 (N_26220,N_24435,N_25463);
nor U26221 (N_26221,N_24959,N_25235);
nor U26222 (N_26222,N_25174,N_24925);
and U26223 (N_26223,N_24637,N_24391);
and U26224 (N_26224,N_25132,N_24509);
nor U26225 (N_26225,N_25484,N_24302);
nor U26226 (N_26226,N_24778,N_24366);
or U26227 (N_26227,N_25340,N_25022);
xnor U26228 (N_26228,N_25262,N_25448);
or U26229 (N_26229,N_25471,N_25218);
or U26230 (N_26230,N_24086,N_24023);
nand U26231 (N_26231,N_25412,N_24074);
and U26232 (N_26232,N_24221,N_24549);
xor U26233 (N_26233,N_24486,N_24895);
or U26234 (N_26234,N_24339,N_24554);
and U26235 (N_26235,N_24254,N_24313);
nor U26236 (N_26236,N_24769,N_25078);
xor U26237 (N_26237,N_25039,N_24498);
xor U26238 (N_26238,N_24310,N_24531);
and U26239 (N_26239,N_25155,N_25041);
and U26240 (N_26240,N_24497,N_24686);
nand U26241 (N_26241,N_24962,N_24868);
and U26242 (N_26242,N_24826,N_25301);
xor U26243 (N_26243,N_24565,N_25061);
or U26244 (N_26244,N_24342,N_25397);
nand U26245 (N_26245,N_25332,N_25493);
nand U26246 (N_26246,N_25154,N_25437);
nand U26247 (N_26247,N_24889,N_24170);
and U26248 (N_26248,N_25052,N_24189);
nand U26249 (N_26249,N_24297,N_24001);
nand U26250 (N_26250,N_24197,N_25090);
nor U26251 (N_26251,N_25433,N_25418);
xor U26252 (N_26252,N_25036,N_25104);
nor U26253 (N_26253,N_24138,N_24174);
nand U26254 (N_26254,N_24285,N_24546);
and U26255 (N_26255,N_24900,N_24982);
nand U26256 (N_26256,N_25025,N_24444);
nor U26257 (N_26257,N_24262,N_24724);
xor U26258 (N_26258,N_24840,N_25213);
and U26259 (N_26259,N_25138,N_25121);
nor U26260 (N_26260,N_24701,N_24301);
and U26261 (N_26261,N_25310,N_24909);
xnor U26262 (N_26262,N_24290,N_24087);
or U26263 (N_26263,N_24851,N_24266);
and U26264 (N_26264,N_24110,N_24861);
or U26265 (N_26265,N_24772,N_24599);
or U26266 (N_26266,N_24372,N_24898);
nand U26267 (N_26267,N_24456,N_24320);
or U26268 (N_26268,N_25126,N_24386);
nand U26269 (N_26269,N_24607,N_24998);
xor U26270 (N_26270,N_24114,N_25216);
nor U26271 (N_26271,N_25148,N_24605);
or U26272 (N_26272,N_24555,N_25407);
nand U26273 (N_26273,N_25133,N_25462);
and U26274 (N_26274,N_25076,N_24379);
nand U26275 (N_26275,N_25085,N_25451);
xnor U26276 (N_26276,N_24334,N_24998);
xnor U26277 (N_26277,N_24192,N_24505);
or U26278 (N_26278,N_24092,N_24377);
xor U26279 (N_26279,N_24153,N_24026);
nor U26280 (N_26280,N_24481,N_25283);
nand U26281 (N_26281,N_25112,N_24498);
or U26282 (N_26282,N_24193,N_24993);
nand U26283 (N_26283,N_24755,N_24691);
or U26284 (N_26284,N_24091,N_24077);
xnor U26285 (N_26285,N_24120,N_24029);
nand U26286 (N_26286,N_24364,N_24522);
and U26287 (N_26287,N_25222,N_24171);
nor U26288 (N_26288,N_24461,N_24661);
and U26289 (N_26289,N_24327,N_24560);
or U26290 (N_26290,N_24650,N_25153);
xor U26291 (N_26291,N_24697,N_25221);
and U26292 (N_26292,N_24445,N_24472);
nand U26293 (N_26293,N_24498,N_24639);
nand U26294 (N_26294,N_25336,N_25109);
nor U26295 (N_26295,N_24519,N_24488);
or U26296 (N_26296,N_25065,N_24725);
and U26297 (N_26297,N_25400,N_24908);
xnor U26298 (N_26298,N_25347,N_24722);
nand U26299 (N_26299,N_24495,N_25037);
or U26300 (N_26300,N_24164,N_24444);
nor U26301 (N_26301,N_24199,N_25469);
or U26302 (N_26302,N_24845,N_24164);
or U26303 (N_26303,N_24297,N_24547);
nand U26304 (N_26304,N_25153,N_24192);
and U26305 (N_26305,N_24051,N_25279);
and U26306 (N_26306,N_24131,N_25345);
nor U26307 (N_26307,N_24181,N_24142);
xor U26308 (N_26308,N_24945,N_24561);
and U26309 (N_26309,N_25266,N_24149);
or U26310 (N_26310,N_24700,N_24495);
nand U26311 (N_26311,N_24746,N_24610);
xnor U26312 (N_26312,N_25469,N_25006);
nand U26313 (N_26313,N_24220,N_25380);
nor U26314 (N_26314,N_24808,N_25280);
and U26315 (N_26315,N_24111,N_24496);
nand U26316 (N_26316,N_24507,N_24555);
nand U26317 (N_26317,N_24810,N_24605);
or U26318 (N_26318,N_24764,N_25392);
nand U26319 (N_26319,N_25053,N_24272);
or U26320 (N_26320,N_24534,N_24732);
or U26321 (N_26321,N_24588,N_24825);
nor U26322 (N_26322,N_25364,N_25312);
nor U26323 (N_26323,N_24095,N_25098);
or U26324 (N_26324,N_25191,N_25117);
xor U26325 (N_26325,N_25146,N_24349);
xnor U26326 (N_26326,N_24886,N_24277);
nand U26327 (N_26327,N_24753,N_24459);
nor U26328 (N_26328,N_25449,N_24322);
nand U26329 (N_26329,N_25447,N_24834);
nor U26330 (N_26330,N_24261,N_24831);
or U26331 (N_26331,N_25399,N_25440);
or U26332 (N_26332,N_24405,N_25200);
and U26333 (N_26333,N_24642,N_24399);
xnor U26334 (N_26334,N_24675,N_24571);
or U26335 (N_26335,N_24145,N_25288);
xnor U26336 (N_26336,N_24078,N_25173);
or U26337 (N_26337,N_24648,N_24547);
and U26338 (N_26338,N_25367,N_24651);
or U26339 (N_26339,N_25212,N_24522);
xor U26340 (N_26340,N_24720,N_24731);
nor U26341 (N_26341,N_25022,N_24389);
or U26342 (N_26342,N_25481,N_25320);
nand U26343 (N_26343,N_24737,N_24085);
xnor U26344 (N_26344,N_24273,N_25106);
or U26345 (N_26345,N_25446,N_25437);
nor U26346 (N_26346,N_24414,N_25017);
nor U26347 (N_26347,N_24824,N_24774);
and U26348 (N_26348,N_24511,N_25092);
nand U26349 (N_26349,N_24589,N_24829);
nor U26350 (N_26350,N_24939,N_25218);
xnor U26351 (N_26351,N_24577,N_24802);
nor U26352 (N_26352,N_24414,N_25242);
xnor U26353 (N_26353,N_24324,N_25336);
or U26354 (N_26354,N_24721,N_25122);
nor U26355 (N_26355,N_25028,N_24275);
or U26356 (N_26356,N_24700,N_25484);
nor U26357 (N_26357,N_25239,N_24696);
and U26358 (N_26358,N_24338,N_24968);
nor U26359 (N_26359,N_24416,N_24666);
or U26360 (N_26360,N_24988,N_24490);
and U26361 (N_26361,N_24231,N_24519);
nand U26362 (N_26362,N_24388,N_25456);
or U26363 (N_26363,N_25486,N_25152);
nand U26364 (N_26364,N_24462,N_24966);
nand U26365 (N_26365,N_25360,N_25361);
nand U26366 (N_26366,N_24699,N_24632);
xnor U26367 (N_26367,N_25184,N_24069);
nor U26368 (N_26368,N_25369,N_24578);
nand U26369 (N_26369,N_24827,N_24724);
or U26370 (N_26370,N_25442,N_25319);
nand U26371 (N_26371,N_25401,N_25173);
xnor U26372 (N_26372,N_24199,N_24761);
nand U26373 (N_26373,N_25122,N_24447);
nor U26374 (N_26374,N_25367,N_24391);
nor U26375 (N_26375,N_24249,N_25416);
and U26376 (N_26376,N_24871,N_25453);
or U26377 (N_26377,N_24819,N_24553);
nand U26378 (N_26378,N_24616,N_24967);
nand U26379 (N_26379,N_24114,N_24580);
nor U26380 (N_26380,N_24267,N_25049);
nor U26381 (N_26381,N_24638,N_25364);
nand U26382 (N_26382,N_24361,N_24619);
nand U26383 (N_26383,N_24348,N_25080);
or U26384 (N_26384,N_24845,N_24000);
nand U26385 (N_26385,N_25395,N_24712);
or U26386 (N_26386,N_25469,N_24928);
nand U26387 (N_26387,N_25044,N_24150);
xor U26388 (N_26388,N_24993,N_24744);
nand U26389 (N_26389,N_24760,N_24522);
nor U26390 (N_26390,N_24896,N_24603);
and U26391 (N_26391,N_24871,N_24139);
nand U26392 (N_26392,N_24078,N_24555);
or U26393 (N_26393,N_25171,N_25479);
xor U26394 (N_26394,N_24320,N_25419);
xnor U26395 (N_26395,N_25002,N_24817);
or U26396 (N_26396,N_25281,N_25180);
or U26397 (N_26397,N_24418,N_25268);
or U26398 (N_26398,N_24348,N_24841);
nor U26399 (N_26399,N_24252,N_25289);
or U26400 (N_26400,N_24012,N_25174);
xnor U26401 (N_26401,N_24894,N_24579);
or U26402 (N_26402,N_25346,N_25190);
nor U26403 (N_26403,N_24699,N_24965);
nor U26404 (N_26404,N_24710,N_25083);
nand U26405 (N_26405,N_24352,N_24981);
nor U26406 (N_26406,N_24657,N_24598);
or U26407 (N_26407,N_25003,N_24797);
or U26408 (N_26408,N_24197,N_24176);
xor U26409 (N_26409,N_24115,N_24760);
xnor U26410 (N_26410,N_25096,N_25367);
nor U26411 (N_26411,N_24269,N_25112);
and U26412 (N_26412,N_25308,N_24321);
nand U26413 (N_26413,N_24858,N_25486);
nor U26414 (N_26414,N_24235,N_24762);
and U26415 (N_26415,N_25241,N_24349);
and U26416 (N_26416,N_24366,N_24789);
or U26417 (N_26417,N_25027,N_25224);
nor U26418 (N_26418,N_24680,N_24903);
nor U26419 (N_26419,N_25115,N_24798);
nor U26420 (N_26420,N_24225,N_24727);
and U26421 (N_26421,N_24616,N_24426);
nand U26422 (N_26422,N_24406,N_24144);
and U26423 (N_26423,N_24600,N_25417);
nor U26424 (N_26424,N_24298,N_24887);
or U26425 (N_26425,N_25009,N_25124);
nand U26426 (N_26426,N_24708,N_24040);
nor U26427 (N_26427,N_25430,N_25266);
nand U26428 (N_26428,N_24366,N_24384);
or U26429 (N_26429,N_24382,N_24629);
nor U26430 (N_26430,N_25079,N_24174);
and U26431 (N_26431,N_24883,N_25465);
xor U26432 (N_26432,N_25167,N_24507);
or U26433 (N_26433,N_24725,N_24834);
xnor U26434 (N_26434,N_25242,N_25218);
xnor U26435 (N_26435,N_24801,N_25178);
nand U26436 (N_26436,N_24791,N_24188);
xnor U26437 (N_26437,N_24422,N_24058);
nand U26438 (N_26438,N_25235,N_24944);
and U26439 (N_26439,N_24119,N_25489);
xor U26440 (N_26440,N_25241,N_25389);
and U26441 (N_26441,N_24014,N_25452);
or U26442 (N_26442,N_24120,N_24758);
or U26443 (N_26443,N_25200,N_25272);
nor U26444 (N_26444,N_24606,N_25140);
and U26445 (N_26445,N_24545,N_24986);
and U26446 (N_26446,N_24993,N_24290);
or U26447 (N_26447,N_24329,N_24162);
nand U26448 (N_26448,N_24038,N_25292);
xor U26449 (N_26449,N_24142,N_24138);
and U26450 (N_26450,N_25078,N_24551);
nor U26451 (N_26451,N_24803,N_24860);
nand U26452 (N_26452,N_24049,N_25382);
and U26453 (N_26453,N_24371,N_24886);
xnor U26454 (N_26454,N_25074,N_24127);
nor U26455 (N_26455,N_24560,N_24486);
and U26456 (N_26456,N_24104,N_24636);
nand U26457 (N_26457,N_25178,N_25342);
and U26458 (N_26458,N_24239,N_25313);
nor U26459 (N_26459,N_24122,N_25098);
or U26460 (N_26460,N_24031,N_24056);
nand U26461 (N_26461,N_24003,N_24835);
or U26462 (N_26462,N_25455,N_24968);
xnor U26463 (N_26463,N_24616,N_25451);
nand U26464 (N_26464,N_24073,N_25385);
or U26465 (N_26465,N_24741,N_25436);
nor U26466 (N_26466,N_24144,N_25207);
nand U26467 (N_26467,N_24248,N_25223);
xnor U26468 (N_26468,N_24068,N_24333);
and U26469 (N_26469,N_24417,N_25144);
nor U26470 (N_26470,N_24091,N_25110);
or U26471 (N_26471,N_24820,N_24182);
nor U26472 (N_26472,N_24095,N_25029);
nand U26473 (N_26473,N_25200,N_24971);
and U26474 (N_26474,N_25400,N_25227);
or U26475 (N_26475,N_24912,N_24388);
or U26476 (N_26476,N_24910,N_24468);
or U26477 (N_26477,N_24146,N_24636);
xnor U26478 (N_26478,N_24352,N_24757);
nor U26479 (N_26479,N_24794,N_24625);
nor U26480 (N_26480,N_24045,N_25118);
and U26481 (N_26481,N_24455,N_25125);
nand U26482 (N_26482,N_24998,N_25494);
or U26483 (N_26483,N_24882,N_24252);
nor U26484 (N_26484,N_24803,N_25232);
and U26485 (N_26485,N_25162,N_24863);
and U26486 (N_26486,N_25395,N_25382);
xnor U26487 (N_26487,N_24871,N_25318);
nand U26488 (N_26488,N_25299,N_24011);
and U26489 (N_26489,N_24292,N_24670);
nor U26490 (N_26490,N_24508,N_24428);
nor U26491 (N_26491,N_25441,N_25427);
or U26492 (N_26492,N_25338,N_24113);
and U26493 (N_26493,N_25420,N_25441);
or U26494 (N_26494,N_25250,N_25107);
and U26495 (N_26495,N_24752,N_24845);
nor U26496 (N_26496,N_25440,N_24862);
nand U26497 (N_26497,N_24700,N_24976);
or U26498 (N_26498,N_25450,N_25277);
xor U26499 (N_26499,N_24102,N_24361);
xor U26500 (N_26500,N_25104,N_25432);
nor U26501 (N_26501,N_24121,N_24210);
nor U26502 (N_26502,N_24902,N_24601);
and U26503 (N_26503,N_24828,N_25206);
nand U26504 (N_26504,N_24436,N_24773);
nand U26505 (N_26505,N_24001,N_25040);
nand U26506 (N_26506,N_25068,N_25411);
nand U26507 (N_26507,N_24633,N_24294);
nor U26508 (N_26508,N_24940,N_25289);
nor U26509 (N_26509,N_24658,N_24714);
xnor U26510 (N_26510,N_25332,N_24812);
nand U26511 (N_26511,N_24846,N_25168);
and U26512 (N_26512,N_24865,N_24428);
nand U26513 (N_26513,N_24509,N_24981);
nor U26514 (N_26514,N_24340,N_25238);
nand U26515 (N_26515,N_25121,N_24797);
nor U26516 (N_26516,N_24073,N_24558);
and U26517 (N_26517,N_25411,N_25132);
and U26518 (N_26518,N_24647,N_24678);
xor U26519 (N_26519,N_24184,N_24843);
nor U26520 (N_26520,N_25295,N_25433);
nor U26521 (N_26521,N_25281,N_25481);
nor U26522 (N_26522,N_24898,N_24180);
nand U26523 (N_26523,N_25446,N_25383);
or U26524 (N_26524,N_25206,N_24384);
xor U26525 (N_26525,N_24757,N_24543);
nor U26526 (N_26526,N_25284,N_24295);
nor U26527 (N_26527,N_24005,N_24699);
and U26528 (N_26528,N_24648,N_24541);
xor U26529 (N_26529,N_24853,N_24931);
and U26530 (N_26530,N_24898,N_24919);
nor U26531 (N_26531,N_25057,N_25393);
nor U26532 (N_26532,N_24952,N_24377);
xor U26533 (N_26533,N_24632,N_25292);
nand U26534 (N_26534,N_24486,N_25348);
and U26535 (N_26535,N_25338,N_24305);
xnor U26536 (N_26536,N_24470,N_24010);
nand U26537 (N_26537,N_24649,N_24571);
xor U26538 (N_26538,N_25264,N_24333);
xnor U26539 (N_26539,N_24420,N_24440);
xor U26540 (N_26540,N_24054,N_24108);
xnor U26541 (N_26541,N_25208,N_25201);
nand U26542 (N_26542,N_24155,N_25177);
or U26543 (N_26543,N_25387,N_24375);
nor U26544 (N_26544,N_24550,N_25002);
nand U26545 (N_26545,N_25455,N_25052);
nor U26546 (N_26546,N_24702,N_24920);
and U26547 (N_26547,N_25088,N_24194);
or U26548 (N_26548,N_25218,N_24139);
and U26549 (N_26549,N_25010,N_24259);
nand U26550 (N_26550,N_25287,N_24006);
and U26551 (N_26551,N_24952,N_25226);
or U26552 (N_26552,N_25125,N_25178);
nor U26553 (N_26553,N_24503,N_24456);
and U26554 (N_26554,N_24920,N_24792);
xnor U26555 (N_26555,N_24519,N_25254);
or U26556 (N_26556,N_24128,N_24156);
and U26557 (N_26557,N_24305,N_24673);
or U26558 (N_26558,N_24015,N_25474);
xnor U26559 (N_26559,N_24939,N_24457);
xor U26560 (N_26560,N_24884,N_24498);
xnor U26561 (N_26561,N_24781,N_24375);
and U26562 (N_26562,N_25340,N_25304);
xnor U26563 (N_26563,N_25432,N_24724);
or U26564 (N_26564,N_24430,N_24545);
nand U26565 (N_26565,N_24072,N_24114);
nand U26566 (N_26566,N_25268,N_24232);
xor U26567 (N_26567,N_24187,N_24142);
or U26568 (N_26568,N_24231,N_24673);
nand U26569 (N_26569,N_24136,N_24295);
nor U26570 (N_26570,N_24064,N_24761);
or U26571 (N_26571,N_25230,N_25294);
nor U26572 (N_26572,N_24341,N_24092);
nor U26573 (N_26573,N_25263,N_24489);
nor U26574 (N_26574,N_24489,N_24472);
or U26575 (N_26575,N_24750,N_25230);
and U26576 (N_26576,N_24021,N_24119);
xor U26577 (N_26577,N_24684,N_24925);
and U26578 (N_26578,N_24949,N_24405);
or U26579 (N_26579,N_24395,N_25451);
and U26580 (N_26580,N_24430,N_24477);
or U26581 (N_26581,N_25365,N_24620);
nor U26582 (N_26582,N_24966,N_24539);
and U26583 (N_26583,N_25144,N_24085);
and U26584 (N_26584,N_25279,N_25214);
and U26585 (N_26585,N_24274,N_24331);
or U26586 (N_26586,N_24658,N_24721);
or U26587 (N_26587,N_24029,N_24965);
xnor U26588 (N_26588,N_24735,N_24357);
nand U26589 (N_26589,N_25387,N_25374);
nand U26590 (N_26590,N_24362,N_25263);
or U26591 (N_26591,N_24222,N_24694);
or U26592 (N_26592,N_25408,N_24197);
and U26593 (N_26593,N_25270,N_25304);
xor U26594 (N_26594,N_25170,N_24312);
xor U26595 (N_26595,N_24575,N_24228);
nand U26596 (N_26596,N_24938,N_24940);
nand U26597 (N_26597,N_24438,N_24127);
or U26598 (N_26598,N_25467,N_24737);
and U26599 (N_26599,N_24995,N_24762);
or U26600 (N_26600,N_24347,N_24927);
xor U26601 (N_26601,N_24679,N_24215);
nor U26602 (N_26602,N_24297,N_24720);
nand U26603 (N_26603,N_25182,N_24828);
or U26604 (N_26604,N_24087,N_24030);
xor U26605 (N_26605,N_24719,N_24206);
nand U26606 (N_26606,N_24964,N_25259);
xnor U26607 (N_26607,N_25024,N_25430);
or U26608 (N_26608,N_25129,N_25088);
or U26609 (N_26609,N_24131,N_24602);
or U26610 (N_26610,N_25471,N_24424);
xnor U26611 (N_26611,N_24065,N_24391);
nand U26612 (N_26612,N_24634,N_25264);
xor U26613 (N_26613,N_24185,N_24313);
xnor U26614 (N_26614,N_24269,N_24242);
or U26615 (N_26615,N_24704,N_24069);
and U26616 (N_26616,N_24259,N_24337);
xnor U26617 (N_26617,N_25324,N_25117);
and U26618 (N_26618,N_25359,N_24087);
nand U26619 (N_26619,N_24135,N_24212);
nand U26620 (N_26620,N_24975,N_25218);
and U26621 (N_26621,N_24041,N_24029);
or U26622 (N_26622,N_25213,N_24843);
nand U26623 (N_26623,N_24113,N_24551);
nor U26624 (N_26624,N_25240,N_24638);
and U26625 (N_26625,N_24231,N_25453);
nor U26626 (N_26626,N_25284,N_25341);
or U26627 (N_26627,N_24086,N_24414);
or U26628 (N_26628,N_24195,N_25472);
nor U26629 (N_26629,N_24917,N_24178);
nor U26630 (N_26630,N_24974,N_24440);
nor U26631 (N_26631,N_24433,N_25101);
nor U26632 (N_26632,N_24937,N_24706);
and U26633 (N_26633,N_24991,N_25321);
nand U26634 (N_26634,N_25330,N_25059);
nand U26635 (N_26635,N_24065,N_25462);
and U26636 (N_26636,N_25452,N_24745);
nand U26637 (N_26637,N_24369,N_24204);
nand U26638 (N_26638,N_24474,N_25333);
and U26639 (N_26639,N_24075,N_24645);
or U26640 (N_26640,N_24295,N_24876);
and U26641 (N_26641,N_25252,N_24998);
nor U26642 (N_26642,N_24623,N_24015);
xnor U26643 (N_26643,N_25112,N_24583);
nor U26644 (N_26644,N_24323,N_24531);
or U26645 (N_26645,N_24170,N_25025);
and U26646 (N_26646,N_25019,N_24906);
and U26647 (N_26647,N_24550,N_25478);
nand U26648 (N_26648,N_25350,N_24131);
or U26649 (N_26649,N_25170,N_25209);
and U26650 (N_26650,N_24963,N_24513);
and U26651 (N_26651,N_25147,N_24398);
nor U26652 (N_26652,N_24787,N_24335);
or U26653 (N_26653,N_24747,N_24431);
nor U26654 (N_26654,N_24330,N_24564);
nand U26655 (N_26655,N_24510,N_24497);
or U26656 (N_26656,N_25175,N_24629);
nand U26657 (N_26657,N_24416,N_24084);
xnor U26658 (N_26658,N_25070,N_25194);
nand U26659 (N_26659,N_24055,N_25352);
nor U26660 (N_26660,N_24684,N_24381);
nor U26661 (N_26661,N_25064,N_24852);
nor U26662 (N_26662,N_24681,N_25151);
nand U26663 (N_26663,N_24291,N_24609);
nor U26664 (N_26664,N_24235,N_24891);
or U26665 (N_26665,N_25259,N_25004);
nor U26666 (N_26666,N_25399,N_24097);
or U26667 (N_26667,N_25137,N_25299);
nand U26668 (N_26668,N_25297,N_24606);
nand U26669 (N_26669,N_24638,N_24585);
or U26670 (N_26670,N_24140,N_25020);
and U26671 (N_26671,N_24520,N_24926);
xnor U26672 (N_26672,N_25397,N_25420);
nand U26673 (N_26673,N_24669,N_25036);
nand U26674 (N_26674,N_24539,N_24010);
xor U26675 (N_26675,N_25328,N_24524);
xnor U26676 (N_26676,N_24069,N_24091);
xor U26677 (N_26677,N_25279,N_25347);
or U26678 (N_26678,N_24961,N_24312);
xnor U26679 (N_26679,N_24198,N_24539);
xnor U26680 (N_26680,N_25297,N_24429);
or U26681 (N_26681,N_24105,N_24541);
nand U26682 (N_26682,N_25229,N_25439);
nor U26683 (N_26683,N_24679,N_24496);
nor U26684 (N_26684,N_24625,N_24460);
or U26685 (N_26685,N_24510,N_25035);
or U26686 (N_26686,N_24368,N_25345);
nor U26687 (N_26687,N_25000,N_25214);
nor U26688 (N_26688,N_24376,N_25024);
nand U26689 (N_26689,N_24179,N_25099);
or U26690 (N_26690,N_24000,N_25381);
and U26691 (N_26691,N_25448,N_24490);
xnor U26692 (N_26692,N_25185,N_25324);
or U26693 (N_26693,N_24845,N_24271);
nand U26694 (N_26694,N_24652,N_25235);
xnor U26695 (N_26695,N_25065,N_25226);
nor U26696 (N_26696,N_24022,N_24567);
nor U26697 (N_26697,N_24532,N_24296);
nor U26698 (N_26698,N_24640,N_25233);
or U26699 (N_26699,N_24106,N_24630);
nor U26700 (N_26700,N_24919,N_24441);
or U26701 (N_26701,N_24577,N_24254);
nand U26702 (N_26702,N_25381,N_24386);
and U26703 (N_26703,N_24090,N_25158);
or U26704 (N_26704,N_24308,N_24648);
nand U26705 (N_26705,N_24220,N_24346);
xor U26706 (N_26706,N_24887,N_25474);
xor U26707 (N_26707,N_24895,N_25180);
and U26708 (N_26708,N_25439,N_24980);
nor U26709 (N_26709,N_25076,N_24260);
nand U26710 (N_26710,N_24990,N_24583);
and U26711 (N_26711,N_24598,N_24854);
nor U26712 (N_26712,N_25108,N_25361);
xnor U26713 (N_26713,N_24099,N_25283);
nand U26714 (N_26714,N_24840,N_25059);
nor U26715 (N_26715,N_24169,N_24479);
xor U26716 (N_26716,N_24543,N_25294);
nor U26717 (N_26717,N_24399,N_24336);
xor U26718 (N_26718,N_24036,N_24275);
xor U26719 (N_26719,N_25055,N_24095);
and U26720 (N_26720,N_25354,N_25466);
and U26721 (N_26721,N_25012,N_24047);
and U26722 (N_26722,N_24382,N_25316);
and U26723 (N_26723,N_25310,N_24798);
or U26724 (N_26724,N_24238,N_24300);
and U26725 (N_26725,N_24872,N_24683);
xnor U26726 (N_26726,N_25415,N_24447);
nor U26727 (N_26727,N_24522,N_24268);
nand U26728 (N_26728,N_24298,N_24056);
and U26729 (N_26729,N_24873,N_24546);
or U26730 (N_26730,N_24149,N_24536);
nand U26731 (N_26731,N_25291,N_25062);
nand U26732 (N_26732,N_24607,N_24997);
xor U26733 (N_26733,N_24388,N_24767);
xnor U26734 (N_26734,N_24484,N_24824);
and U26735 (N_26735,N_25086,N_24968);
or U26736 (N_26736,N_24257,N_25382);
and U26737 (N_26737,N_24102,N_24367);
and U26738 (N_26738,N_24513,N_24510);
nand U26739 (N_26739,N_24479,N_25157);
and U26740 (N_26740,N_25354,N_24980);
or U26741 (N_26741,N_25289,N_24484);
or U26742 (N_26742,N_24079,N_24981);
and U26743 (N_26743,N_25244,N_25135);
nand U26744 (N_26744,N_24091,N_24912);
or U26745 (N_26745,N_24678,N_25196);
xor U26746 (N_26746,N_25395,N_25252);
and U26747 (N_26747,N_24907,N_24515);
or U26748 (N_26748,N_25315,N_25341);
nor U26749 (N_26749,N_24150,N_24026);
xnor U26750 (N_26750,N_25256,N_24404);
nor U26751 (N_26751,N_25001,N_24356);
nor U26752 (N_26752,N_24127,N_25455);
xnor U26753 (N_26753,N_24435,N_24226);
and U26754 (N_26754,N_25135,N_24800);
and U26755 (N_26755,N_24354,N_24761);
or U26756 (N_26756,N_24790,N_24348);
or U26757 (N_26757,N_25358,N_24420);
or U26758 (N_26758,N_25400,N_25411);
and U26759 (N_26759,N_24735,N_25106);
and U26760 (N_26760,N_24761,N_25013);
and U26761 (N_26761,N_24566,N_24842);
or U26762 (N_26762,N_25398,N_24903);
or U26763 (N_26763,N_25456,N_25139);
xor U26764 (N_26764,N_24071,N_24413);
and U26765 (N_26765,N_24170,N_25323);
xnor U26766 (N_26766,N_24477,N_24697);
nand U26767 (N_26767,N_25443,N_24096);
and U26768 (N_26768,N_24876,N_24065);
and U26769 (N_26769,N_24147,N_25246);
nand U26770 (N_26770,N_24963,N_25446);
and U26771 (N_26771,N_24010,N_24261);
nand U26772 (N_26772,N_24159,N_24031);
and U26773 (N_26773,N_24578,N_24920);
nor U26774 (N_26774,N_24204,N_24563);
and U26775 (N_26775,N_24445,N_24580);
and U26776 (N_26776,N_24799,N_24082);
or U26777 (N_26777,N_24462,N_24839);
nor U26778 (N_26778,N_25424,N_25075);
nand U26779 (N_26779,N_25008,N_25218);
or U26780 (N_26780,N_24392,N_24600);
xor U26781 (N_26781,N_25374,N_24794);
nand U26782 (N_26782,N_24555,N_24148);
and U26783 (N_26783,N_25082,N_24353);
xor U26784 (N_26784,N_24440,N_25281);
nand U26785 (N_26785,N_24576,N_24938);
nor U26786 (N_26786,N_24796,N_24524);
nor U26787 (N_26787,N_25451,N_24634);
and U26788 (N_26788,N_24011,N_24517);
nand U26789 (N_26789,N_25432,N_24705);
nor U26790 (N_26790,N_25275,N_24565);
nand U26791 (N_26791,N_24169,N_24739);
or U26792 (N_26792,N_24320,N_24361);
or U26793 (N_26793,N_24414,N_24534);
and U26794 (N_26794,N_24238,N_24464);
xnor U26795 (N_26795,N_24514,N_24765);
nor U26796 (N_26796,N_24648,N_25158);
nand U26797 (N_26797,N_24792,N_24789);
nand U26798 (N_26798,N_24476,N_25448);
or U26799 (N_26799,N_25232,N_24447);
xnor U26800 (N_26800,N_24749,N_24128);
nand U26801 (N_26801,N_24638,N_24144);
xnor U26802 (N_26802,N_25094,N_24839);
nand U26803 (N_26803,N_24570,N_24955);
nand U26804 (N_26804,N_24889,N_24762);
or U26805 (N_26805,N_24623,N_24882);
xnor U26806 (N_26806,N_24458,N_25459);
or U26807 (N_26807,N_24813,N_24938);
and U26808 (N_26808,N_24039,N_24684);
xnor U26809 (N_26809,N_25078,N_24194);
nor U26810 (N_26810,N_24998,N_25100);
and U26811 (N_26811,N_24519,N_25439);
and U26812 (N_26812,N_24539,N_25451);
xor U26813 (N_26813,N_24094,N_25402);
nand U26814 (N_26814,N_24946,N_24191);
and U26815 (N_26815,N_24328,N_24141);
and U26816 (N_26816,N_24102,N_24196);
xnor U26817 (N_26817,N_24672,N_25182);
nor U26818 (N_26818,N_24138,N_25373);
and U26819 (N_26819,N_24228,N_25164);
and U26820 (N_26820,N_24226,N_24746);
or U26821 (N_26821,N_24585,N_24981);
and U26822 (N_26822,N_24973,N_25268);
and U26823 (N_26823,N_24741,N_24623);
and U26824 (N_26824,N_25035,N_24641);
or U26825 (N_26825,N_24624,N_24897);
or U26826 (N_26826,N_24384,N_24248);
and U26827 (N_26827,N_24017,N_24846);
and U26828 (N_26828,N_24143,N_24342);
xnor U26829 (N_26829,N_25422,N_25116);
nor U26830 (N_26830,N_25114,N_25431);
or U26831 (N_26831,N_24328,N_24807);
xnor U26832 (N_26832,N_25084,N_24789);
nand U26833 (N_26833,N_25150,N_24912);
xnor U26834 (N_26834,N_24380,N_24582);
nor U26835 (N_26835,N_24029,N_25477);
or U26836 (N_26836,N_25000,N_25397);
xnor U26837 (N_26837,N_24592,N_24543);
and U26838 (N_26838,N_25452,N_24571);
xnor U26839 (N_26839,N_25106,N_24229);
nand U26840 (N_26840,N_24737,N_24138);
nor U26841 (N_26841,N_24226,N_25406);
nand U26842 (N_26842,N_25104,N_24435);
or U26843 (N_26843,N_24947,N_24164);
and U26844 (N_26844,N_24042,N_24881);
xor U26845 (N_26845,N_25036,N_24537);
nor U26846 (N_26846,N_24668,N_25042);
and U26847 (N_26847,N_24644,N_24719);
nand U26848 (N_26848,N_24650,N_24669);
or U26849 (N_26849,N_24108,N_25319);
nand U26850 (N_26850,N_24308,N_24695);
xnor U26851 (N_26851,N_24594,N_24822);
and U26852 (N_26852,N_24584,N_25242);
xnor U26853 (N_26853,N_24153,N_24039);
nor U26854 (N_26854,N_24916,N_24319);
and U26855 (N_26855,N_24487,N_24469);
xnor U26856 (N_26856,N_24963,N_24381);
nor U26857 (N_26857,N_24745,N_25331);
and U26858 (N_26858,N_24767,N_24029);
nor U26859 (N_26859,N_24716,N_24663);
and U26860 (N_26860,N_25466,N_24232);
xor U26861 (N_26861,N_24352,N_24272);
or U26862 (N_26862,N_24897,N_25009);
xor U26863 (N_26863,N_24027,N_25449);
xor U26864 (N_26864,N_24257,N_24858);
xnor U26865 (N_26865,N_24996,N_24491);
xor U26866 (N_26866,N_24799,N_24948);
xnor U26867 (N_26867,N_24623,N_25158);
xor U26868 (N_26868,N_25254,N_24268);
and U26869 (N_26869,N_25141,N_24752);
xor U26870 (N_26870,N_25081,N_24532);
and U26871 (N_26871,N_24470,N_24526);
and U26872 (N_26872,N_24833,N_24201);
nor U26873 (N_26873,N_25324,N_24113);
nand U26874 (N_26874,N_24666,N_24815);
or U26875 (N_26875,N_24339,N_25385);
nand U26876 (N_26876,N_24804,N_25263);
or U26877 (N_26877,N_25063,N_25480);
nand U26878 (N_26878,N_25441,N_25033);
nand U26879 (N_26879,N_24034,N_25473);
nor U26880 (N_26880,N_25422,N_24607);
nand U26881 (N_26881,N_24838,N_24014);
nor U26882 (N_26882,N_24387,N_24543);
or U26883 (N_26883,N_24572,N_24345);
nor U26884 (N_26884,N_25367,N_24756);
xnor U26885 (N_26885,N_25027,N_24695);
xor U26886 (N_26886,N_24723,N_25123);
nand U26887 (N_26887,N_24907,N_25336);
nor U26888 (N_26888,N_24231,N_24429);
nand U26889 (N_26889,N_24031,N_24020);
nor U26890 (N_26890,N_24730,N_24250);
xor U26891 (N_26891,N_24211,N_25053);
or U26892 (N_26892,N_25020,N_24434);
nand U26893 (N_26893,N_24291,N_25093);
nand U26894 (N_26894,N_24978,N_25096);
xor U26895 (N_26895,N_24889,N_24143);
or U26896 (N_26896,N_24950,N_25219);
or U26897 (N_26897,N_24423,N_24539);
nor U26898 (N_26898,N_25034,N_25386);
nor U26899 (N_26899,N_25240,N_24577);
or U26900 (N_26900,N_24408,N_25405);
xnor U26901 (N_26901,N_24897,N_24455);
and U26902 (N_26902,N_24393,N_24356);
xnor U26903 (N_26903,N_24674,N_25481);
or U26904 (N_26904,N_24840,N_25093);
nand U26905 (N_26905,N_24548,N_24971);
and U26906 (N_26906,N_24552,N_24969);
xor U26907 (N_26907,N_24665,N_24896);
xnor U26908 (N_26908,N_24149,N_24400);
xor U26909 (N_26909,N_25207,N_25194);
nor U26910 (N_26910,N_25414,N_24725);
nor U26911 (N_26911,N_25348,N_25024);
nor U26912 (N_26912,N_24910,N_25489);
nor U26913 (N_26913,N_24869,N_24360);
and U26914 (N_26914,N_25317,N_24488);
xnor U26915 (N_26915,N_24415,N_24395);
nand U26916 (N_26916,N_24435,N_24108);
or U26917 (N_26917,N_25226,N_24815);
and U26918 (N_26918,N_24525,N_25023);
xnor U26919 (N_26919,N_25335,N_25067);
xnor U26920 (N_26920,N_25104,N_24381);
nor U26921 (N_26921,N_25226,N_25306);
or U26922 (N_26922,N_25358,N_24671);
nor U26923 (N_26923,N_24919,N_24750);
and U26924 (N_26924,N_24303,N_25243);
nand U26925 (N_26925,N_24910,N_24041);
nor U26926 (N_26926,N_24847,N_24242);
and U26927 (N_26927,N_24477,N_24257);
xnor U26928 (N_26928,N_24859,N_24620);
xnor U26929 (N_26929,N_25332,N_24813);
nand U26930 (N_26930,N_24782,N_24772);
nand U26931 (N_26931,N_24790,N_24394);
nand U26932 (N_26932,N_25139,N_25305);
and U26933 (N_26933,N_24670,N_24557);
xor U26934 (N_26934,N_25233,N_25303);
or U26935 (N_26935,N_24551,N_24281);
and U26936 (N_26936,N_25102,N_24094);
nand U26937 (N_26937,N_25139,N_24655);
or U26938 (N_26938,N_25451,N_24792);
and U26939 (N_26939,N_25449,N_24730);
or U26940 (N_26940,N_25453,N_24322);
nor U26941 (N_26941,N_24786,N_25458);
nor U26942 (N_26942,N_24696,N_24744);
and U26943 (N_26943,N_24523,N_24568);
or U26944 (N_26944,N_25231,N_24015);
nor U26945 (N_26945,N_24688,N_24973);
or U26946 (N_26946,N_25052,N_24572);
or U26947 (N_26947,N_24332,N_24724);
xor U26948 (N_26948,N_24416,N_25309);
xnor U26949 (N_26949,N_24168,N_24003);
xor U26950 (N_26950,N_24388,N_24874);
nor U26951 (N_26951,N_24863,N_25222);
nor U26952 (N_26952,N_25425,N_25480);
nand U26953 (N_26953,N_24542,N_25423);
nand U26954 (N_26954,N_25200,N_24621);
nand U26955 (N_26955,N_25235,N_24370);
and U26956 (N_26956,N_25161,N_24848);
nand U26957 (N_26957,N_24593,N_25476);
nand U26958 (N_26958,N_24223,N_24326);
nor U26959 (N_26959,N_24143,N_24715);
xnor U26960 (N_26960,N_24406,N_24452);
xnor U26961 (N_26961,N_25372,N_24020);
and U26962 (N_26962,N_24851,N_25448);
xor U26963 (N_26963,N_25418,N_24210);
and U26964 (N_26964,N_25328,N_24402);
xor U26965 (N_26965,N_24988,N_24690);
or U26966 (N_26966,N_25445,N_24530);
or U26967 (N_26967,N_24824,N_24561);
or U26968 (N_26968,N_24568,N_25070);
nor U26969 (N_26969,N_24352,N_25404);
or U26970 (N_26970,N_24936,N_24792);
nand U26971 (N_26971,N_24891,N_25215);
xnor U26972 (N_26972,N_25123,N_25080);
nand U26973 (N_26973,N_25303,N_24503);
nand U26974 (N_26974,N_25308,N_24710);
nor U26975 (N_26975,N_24583,N_25486);
xnor U26976 (N_26976,N_25065,N_25133);
or U26977 (N_26977,N_24572,N_24847);
or U26978 (N_26978,N_25396,N_24500);
nor U26979 (N_26979,N_24194,N_24978);
and U26980 (N_26980,N_25381,N_24871);
xnor U26981 (N_26981,N_25039,N_24674);
xnor U26982 (N_26982,N_25213,N_24813);
xor U26983 (N_26983,N_24715,N_25057);
and U26984 (N_26984,N_24101,N_25381);
and U26985 (N_26985,N_24107,N_24011);
nand U26986 (N_26986,N_24521,N_24832);
nor U26987 (N_26987,N_24257,N_24384);
or U26988 (N_26988,N_25065,N_24458);
and U26989 (N_26989,N_25187,N_24678);
or U26990 (N_26990,N_25263,N_24853);
nor U26991 (N_26991,N_25088,N_24620);
and U26992 (N_26992,N_24096,N_24317);
nor U26993 (N_26993,N_24741,N_24891);
or U26994 (N_26994,N_24562,N_24764);
and U26995 (N_26995,N_24851,N_24342);
xnor U26996 (N_26996,N_25213,N_24345);
or U26997 (N_26997,N_25128,N_24759);
xor U26998 (N_26998,N_25098,N_25049);
and U26999 (N_26999,N_24412,N_24616);
xnor U27000 (N_27000,N_25765,N_25722);
and U27001 (N_27001,N_25952,N_26066);
nor U27002 (N_27002,N_26379,N_26905);
or U27003 (N_27003,N_26097,N_26179);
or U27004 (N_27004,N_26679,N_26747);
xnor U27005 (N_27005,N_25978,N_26552);
nor U27006 (N_27006,N_26983,N_26248);
and U27007 (N_27007,N_25552,N_26559);
nor U27008 (N_27008,N_26616,N_26249);
or U27009 (N_27009,N_25850,N_25922);
and U27010 (N_27010,N_26499,N_26801);
xor U27011 (N_27011,N_25646,N_26807);
or U27012 (N_27012,N_26207,N_26105);
nand U27013 (N_27013,N_26196,N_25670);
nor U27014 (N_27014,N_26129,N_25890);
and U27015 (N_27015,N_26203,N_25676);
xor U27016 (N_27016,N_26871,N_26660);
xnor U27017 (N_27017,N_26082,N_25840);
and U27018 (N_27018,N_26416,N_26316);
nor U27019 (N_27019,N_25699,N_25925);
and U27020 (N_27020,N_26624,N_26091);
xnor U27021 (N_27021,N_25883,N_26818);
and U27022 (N_27022,N_26995,N_25508);
and U27023 (N_27023,N_26694,N_26543);
or U27024 (N_27024,N_26682,N_26511);
or U27025 (N_27025,N_26822,N_26956);
or U27026 (N_27026,N_26057,N_26572);
nand U27027 (N_27027,N_26787,N_26570);
nand U27028 (N_27028,N_26607,N_25982);
nand U27029 (N_27029,N_26696,N_26889);
nor U27030 (N_27030,N_26672,N_26406);
xor U27031 (N_27031,N_26929,N_26612);
nor U27032 (N_27032,N_26111,N_25521);
xor U27033 (N_27033,N_26400,N_25798);
or U27034 (N_27034,N_25664,N_26859);
nand U27035 (N_27035,N_26226,N_25872);
nand U27036 (N_27036,N_26709,N_25945);
nand U27037 (N_27037,N_26974,N_25632);
nor U27038 (N_27038,N_25962,N_25677);
and U27039 (N_27039,N_25750,N_26356);
nand U27040 (N_27040,N_26518,N_26069);
nand U27041 (N_27041,N_25690,N_26132);
nand U27042 (N_27042,N_26899,N_26122);
nand U27043 (N_27043,N_26538,N_26913);
xor U27044 (N_27044,N_25910,N_25814);
nand U27045 (N_27045,N_26458,N_26760);
nand U27046 (N_27046,N_26286,N_26701);
xnor U27047 (N_27047,N_25902,N_26390);
or U27048 (N_27048,N_26233,N_26331);
xnor U27049 (N_27049,N_26988,N_26200);
xnor U27050 (N_27050,N_25913,N_26049);
xnor U27051 (N_27051,N_25635,N_26103);
xnor U27052 (N_27052,N_26231,N_26131);
or U27053 (N_27053,N_25625,N_26460);
and U27054 (N_27054,N_26710,N_26523);
nand U27055 (N_27055,N_25783,N_26445);
xor U27056 (N_27056,N_26405,N_25748);
nor U27057 (N_27057,N_26618,N_26961);
and U27058 (N_27058,N_25611,N_26408);
xor U27059 (N_27059,N_26973,N_26350);
nand U27060 (N_27060,N_26072,N_25874);
nand U27061 (N_27061,N_25881,N_26483);
nor U27062 (N_27062,N_26415,N_26649);
nor U27063 (N_27063,N_25615,N_25606);
xnor U27064 (N_27064,N_26969,N_26150);
or U27065 (N_27065,N_26833,N_26761);
or U27066 (N_27066,N_26068,N_25599);
xnor U27067 (N_27067,N_26904,N_26875);
or U27068 (N_27068,N_26396,N_26100);
or U27069 (N_27069,N_26579,N_26500);
nand U27070 (N_27070,N_25863,N_25667);
nand U27071 (N_27071,N_26133,N_26005);
xor U27072 (N_27072,N_26026,N_25880);
xor U27073 (N_27073,N_26770,N_25973);
or U27074 (N_27074,N_26653,N_26638);
or U27075 (N_27075,N_25708,N_26520);
or U27076 (N_27076,N_26703,N_25774);
or U27077 (N_27077,N_25688,N_26325);
and U27078 (N_27078,N_26490,N_26942);
and U27079 (N_27079,N_26903,N_26213);
nor U27080 (N_27080,N_26711,N_26492);
xor U27081 (N_27081,N_26312,N_26369);
or U27082 (N_27082,N_25551,N_26881);
nor U27083 (N_27083,N_25549,N_25693);
nor U27084 (N_27084,N_26420,N_25991);
nor U27085 (N_27085,N_26724,N_25530);
and U27086 (N_27086,N_25939,N_26853);
and U27087 (N_27087,N_26870,N_25598);
xnor U27088 (N_27088,N_26955,N_26303);
xnor U27089 (N_27089,N_25741,N_26972);
and U27090 (N_27090,N_25852,N_26962);
or U27091 (N_27091,N_26437,N_26298);
xnor U27092 (N_27092,N_26188,N_26240);
xor U27093 (N_27093,N_25640,N_26885);
xnor U27094 (N_27094,N_25532,N_26705);
and U27095 (N_27095,N_25586,N_26773);
xnor U27096 (N_27096,N_26750,N_26832);
xnor U27097 (N_27097,N_26937,N_26178);
nand U27098 (N_27098,N_25697,N_26952);
xor U27099 (N_27099,N_25957,N_25777);
or U27100 (N_27100,N_26181,N_25847);
or U27101 (N_27101,N_25614,N_26451);
nor U27102 (N_27102,N_26510,N_25828);
xnor U27103 (N_27103,N_25658,N_25869);
nand U27104 (N_27104,N_26976,N_26245);
and U27105 (N_27105,N_26153,N_25865);
and U27106 (N_27106,N_26023,N_26975);
or U27107 (N_27107,N_26836,N_26693);
nor U27108 (N_27108,N_26798,N_26762);
and U27109 (N_27109,N_26247,N_26565);
and U27110 (N_27110,N_26002,N_26474);
or U27111 (N_27111,N_26968,N_26439);
xnor U27112 (N_27112,N_25579,N_26235);
and U27113 (N_27113,N_26916,N_26751);
nand U27114 (N_27114,N_26699,N_26868);
nor U27115 (N_27115,N_26075,N_26174);
and U27116 (N_27116,N_26238,N_26222);
nor U27117 (N_27117,N_26475,N_26692);
xnor U27118 (N_27118,N_26009,N_26085);
nor U27119 (N_27119,N_26627,N_26344);
nor U27120 (N_27120,N_26494,N_26923);
nor U27121 (N_27121,N_25637,N_25897);
or U27122 (N_27122,N_26255,N_26504);
or U27123 (N_27123,N_26934,N_26555);
and U27124 (N_27124,N_26834,N_25833);
and U27125 (N_27125,N_26289,N_26996);
and U27126 (N_27126,N_26993,N_25636);
or U27127 (N_27127,N_26927,N_26404);
xor U27128 (N_27128,N_26635,N_25948);
nor U27129 (N_27129,N_26159,N_26733);
nor U27130 (N_27130,N_26382,N_26394);
xor U27131 (N_27131,N_25516,N_26526);
and U27132 (N_27132,N_26381,N_26387);
nor U27133 (N_27133,N_26160,N_25547);
nor U27134 (N_27134,N_26809,N_25590);
and U27135 (N_27135,N_26139,N_25812);
nand U27136 (N_27136,N_26986,N_26880);
nand U27137 (N_27137,N_25935,N_26096);
nand U27138 (N_27138,N_26625,N_25903);
and U27139 (N_27139,N_26055,N_25749);
nand U27140 (N_27140,N_26343,N_25582);
nor U27141 (N_27141,N_25862,N_25984);
or U27142 (N_27142,N_25622,N_26270);
and U27143 (N_27143,N_26623,N_26330);
nand U27144 (N_27144,N_25909,N_26514);
nand U27145 (N_27145,N_25805,N_26723);
and U27146 (N_27146,N_26077,N_25896);
or U27147 (N_27147,N_25976,N_26323);
and U27148 (N_27148,N_26121,N_25643);
and U27149 (N_27149,N_26999,N_25953);
xor U27150 (N_27150,N_26535,N_25936);
nor U27151 (N_27151,N_26357,N_26290);
nand U27152 (N_27152,N_26041,N_25678);
nand U27153 (N_27153,N_26366,N_26363);
nor U27154 (N_27154,N_26315,N_26815);
or U27155 (N_27155,N_25930,N_26496);
nor U27156 (N_27156,N_26658,N_26489);
or U27157 (N_27157,N_26378,N_26027);
nand U27158 (N_27158,N_25796,N_26887);
or U27159 (N_27159,N_26509,N_26865);
and U27160 (N_27160,N_25811,N_25575);
xnor U27161 (N_27161,N_26283,N_26634);
nand U27162 (N_27162,N_26578,N_26680);
nand U27163 (N_27163,N_26182,N_26124);
xnor U27164 (N_27164,N_25761,N_26948);
or U27165 (N_27165,N_26980,N_25555);
xnor U27166 (N_27166,N_26301,N_26838);
or U27167 (N_27167,N_25832,N_25920);
and U27168 (N_27168,N_26257,N_25884);
or U27169 (N_27169,N_26151,N_26361);
and U27170 (N_27170,N_26007,N_26449);
xor U27171 (N_27171,N_25723,N_25797);
nor U27172 (N_27172,N_25639,N_25546);
or U27173 (N_27173,N_25806,N_26730);
nor U27174 (N_27174,N_25914,N_26412);
xnor U27175 (N_27175,N_26950,N_26052);
or U27176 (N_27176,N_26697,N_26383);
xnor U27177 (N_27177,N_26893,N_25698);
or U27178 (N_27178,N_26202,N_26120);
xor U27179 (N_27179,N_25506,N_26757);
and U27180 (N_27180,N_25951,N_25657);
xor U27181 (N_27181,N_26610,N_25556);
or U27182 (N_27182,N_25710,N_26718);
xor U27183 (N_27183,N_26924,N_26266);
xor U27184 (N_27184,N_26668,N_26583);
nor U27185 (N_27185,N_26713,N_26640);
nand U27186 (N_27186,N_26939,N_25545);
xnor U27187 (N_27187,N_26117,N_26531);
or U27188 (N_27188,N_25608,N_26358);
nor U27189 (N_27189,N_25602,N_26154);
nand U27190 (N_27190,N_25908,N_26424);
and U27191 (N_27191,N_25500,N_26090);
xor U27192 (N_27192,N_26727,N_25958);
nand U27193 (N_27193,N_26690,N_25992);
nor U27194 (N_27194,N_26902,N_26519);
nor U27195 (N_27195,N_26130,N_25858);
and U27196 (N_27196,N_25591,N_26210);
or U27197 (N_27197,N_25857,N_26554);
and U27198 (N_27198,N_25648,N_26593);
xnor U27199 (N_27199,N_25975,N_26287);
nor U27200 (N_27200,N_26731,N_26142);
nand U27201 (N_27201,N_25706,N_26843);
xnor U27202 (N_27202,N_26944,N_25911);
nand U27203 (N_27203,N_25559,N_25649);
nor U27204 (N_27204,N_25916,N_26192);
xnor U27205 (N_27205,N_26018,N_26167);
or U27206 (N_27206,N_26146,N_25673);
and U27207 (N_27207,N_26790,N_25770);
xor U27208 (N_27208,N_26766,N_25929);
or U27209 (N_27209,N_26183,N_26528);
xor U27210 (N_27210,N_26646,N_26276);
xor U27211 (N_27211,N_26004,N_26295);
or U27212 (N_27212,N_26087,N_26571);
or U27213 (N_27213,N_25612,N_25986);
and U27214 (N_27214,N_25966,N_26918);
or U27215 (N_27215,N_25877,N_26076);
or U27216 (N_27216,N_25644,N_26294);
and U27217 (N_27217,N_26098,N_26340);
or U27218 (N_27218,N_26687,N_25983);
or U27219 (N_27219,N_25548,N_25729);
and U27220 (N_27220,N_26686,N_26012);
and U27221 (N_27221,N_26503,N_26456);
nor U27222 (N_27222,N_26165,N_26959);
or U27223 (N_27223,N_26862,N_26958);
nor U27224 (N_27224,N_26855,N_26803);
xnor U27225 (N_27225,N_26780,N_25790);
nor U27226 (N_27226,N_25887,N_26546);
or U27227 (N_27227,N_25617,N_26155);
nor U27228 (N_27228,N_25918,N_25701);
or U27229 (N_27229,N_26198,N_26211);
and U27230 (N_27230,N_26926,N_26373);
nor U27231 (N_27231,N_26814,N_26191);
xor U27232 (N_27232,N_26220,N_25836);
nand U27233 (N_27233,N_26837,N_26675);
xnor U27234 (N_27234,N_25515,N_25789);
and U27235 (N_27235,N_26655,N_26367);
and U27236 (N_27236,N_26670,N_25566);
nor U27237 (N_27237,N_26613,N_25999);
and U27238 (N_27238,N_26236,N_26921);
xnor U27239 (N_27239,N_26112,N_26250);
nand U27240 (N_27240,N_26407,N_25653);
and U27241 (N_27241,N_25845,N_26915);
or U27242 (N_27242,N_25569,N_26252);
xor U27243 (N_27243,N_26953,N_26943);
or U27244 (N_27244,N_25771,N_25985);
xnor U27245 (N_27245,N_25853,N_26793);
nand U27246 (N_27246,N_26168,N_25736);
and U27247 (N_27247,N_26830,N_26438);
xor U27248 (N_27248,N_26561,N_26947);
or U27249 (N_27249,N_26669,N_26264);
xnor U27250 (N_27250,N_26397,N_25692);
or U27251 (N_27251,N_25624,N_26332);
xnor U27252 (N_27252,N_26984,N_26059);
nand U27253 (N_27253,N_26721,N_26019);
nor U27254 (N_27254,N_25573,N_25672);
nor U27255 (N_27255,N_26774,N_26548);
nand U27256 (N_27256,N_26001,N_26997);
nor U27257 (N_27257,N_26989,N_26030);
nand U27258 (N_27258,N_26978,N_26472);
or U27259 (N_27259,N_26603,N_26898);
nor U27260 (N_27260,N_26930,N_26597);
nand U27261 (N_27261,N_26386,N_26678);
nor U27262 (N_27262,N_26455,N_26223);
nand U27263 (N_27263,N_25820,N_26043);
nand U27264 (N_27264,N_25600,N_26324);
xnor U27265 (N_27265,N_25921,N_26345);
xnor U27266 (N_27266,N_26015,N_26608);
nand U27267 (N_27267,N_26448,N_26785);
nand U27268 (N_27268,N_26810,N_26204);
xor U27269 (N_27269,N_25915,N_26588);
or U27270 (N_27270,N_26058,N_26278);
and U27271 (N_27271,N_26138,N_25571);
nor U27272 (N_27272,N_26611,N_26062);
nand U27273 (N_27273,N_25661,N_26308);
nor U27274 (N_27274,N_26906,N_25861);
or U27275 (N_27275,N_26605,N_25864);
nand U27276 (N_27276,N_26313,N_25679);
nand U27277 (N_27277,N_26657,N_26190);
xor U27278 (N_27278,N_26089,N_25859);
xnor U27279 (N_27279,N_26883,N_26365);
and U27280 (N_27280,N_26602,N_25717);
and U27281 (N_27281,N_25860,N_26576);
or U27282 (N_27282,N_26740,N_26981);
xnor U27283 (N_27283,N_26544,N_26706);
nand U27284 (N_27284,N_25821,N_26851);
and U27285 (N_27285,N_25627,N_26194);
nor U27286 (N_27286,N_25619,N_26094);
nor U27287 (N_27287,N_26767,N_26073);
or U27288 (N_27288,N_26229,N_25987);
nand U27289 (N_27289,N_26482,N_26212);
and U27290 (N_27290,N_25731,N_26752);
and U27291 (N_27291,N_26877,N_26963);
nor U27292 (N_27292,N_26991,N_26031);
xnor U27293 (N_27293,N_26804,N_25971);
nand U27294 (N_27294,N_26484,N_26466);
and U27295 (N_27295,N_26342,N_25629);
or U27296 (N_27296,N_26435,N_25905);
or U27297 (N_27297,N_26088,N_25507);
and U27298 (N_27298,N_26800,N_25901);
nand U27299 (N_27299,N_26429,N_26442);
or U27300 (N_27300,N_25509,N_25809);
xnor U27301 (N_27301,N_26254,N_25768);
xnor U27302 (N_27302,N_26127,N_26376);
xnor U27303 (N_27303,N_25567,N_26065);
nand U27304 (N_27304,N_26550,N_26674);
or U27305 (N_27305,N_25596,N_26008);
nand U27306 (N_27306,N_26197,N_26487);
nor U27307 (N_27307,N_26932,N_25737);
nand U27308 (N_27308,N_26353,N_25756);
and U27309 (N_27309,N_26779,N_26447);
nor U27310 (N_27310,N_25685,N_26292);
or U27311 (N_27311,N_26631,N_26563);
nand U27312 (N_27312,N_25711,N_26452);
nor U27313 (N_27313,N_26600,N_25659);
nand U27314 (N_27314,N_26081,N_25876);
or U27315 (N_27315,N_26218,N_25968);
and U27316 (N_27316,N_25724,N_25526);
nand U27317 (N_27317,N_26615,N_26735);
xnor U27318 (N_27318,N_25808,N_26113);
or U27319 (N_27319,N_26695,N_26428);
or U27320 (N_27320,N_25965,N_25570);
nor U27321 (N_27321,N_26173,N_26025);
and U27322 (N_27322,N_26951,N_26060);
or U27323 (N_27323,N_25531,N_26849);
xnor U27324 (N_27324,N_26691,N_25686);
or U27325 (N_27325,N_26046,N_26101);
nand U27326 (N_27326,N_26099,N_26527);
and U27327 (N_27327,N_26582,N_26553);
nand U27328 (N_27328,N_25815,N_26243);
and U27329 (N_27329,N_26147,N_26145);
or U27330 (N_27330,N_26890,N_25926);
xor U27331 (N_27331,N_26427,N_25932);
and U27332 (N_27332,N_25666,N_26253);
nor U27333 (N_27333,N_25959,N_26949);
nand U27334 (N_27334,N_26558,N_26063);
or U27335 (N_27335,N_25631,N_26792);
nand U27336 (N_27336,N_26549,N_26219);
or U27337 (N_27337,N_26529,N_26650);
xor U27338 (N_27338,N_25759,N_26891);
or U27339 (N_27339,N_26728,N_26737);
or U27340 (N_27340,N_25517,N_26551);
xnor U27341 (N_27341,N_25684,N_26258);
xnor U27342 (N_27342,N_26388,N_25763);
nand U27343 (N_27343,N_26114,N_26359);
and U27344 (N_27344,N_25618,N_25871);
and U27345 (N_27345,N_25709,N_26506);
or U27346 (N_27346,N_26874,N_25504);
or U27347 (N_27347,N_26601,N_26193);
nand U27348 (N_27348,N_26645,N_25848);
nor U27349 (N_27349,N_26093,N_26022);
xor U27350 (N_27350,N_26216,N_26663);
nor U27351 (N_27351,N_26560,N_25753);
or U27352 (N_27352,N_26311,N_26931);
xor U27353 (N_27353,N_26722,N_25889);
and U27354 (N_27354,N_26628,N_26592);
or U27355 (N_27355,N_25954,N_25824);
and U27356 (N_27356,N_26897,N_26444);
nor U27357 (N_27357,N_26162,N_26187);
or U27358 (N_27358,N_26741,N_26493);
or U27359 (N_27359,N_25947,N_26432);
or U27360 (N_27360,N_26430,N_26346);
xnor U27361 (N_27361,N_26532,N_25937);
xnor U27362 (N_27362,N_26771,N_25513);
and U27363 (N_27363,N_26816,N_25819);
and U27364 (N_27364,N_26821,N_26826);
nand U27365 (N_27365,N_25536,N_26446);
nand U27366 (N_27366,N_25795,N_26010);
nand U27367 (N_27367,N_26037,N_26758);
or U27368 (N_27368,N_25616,N_26199);
or U27369 (N_27369,N_26636,N_26481);
nor U27370 (N_27370,N_26497,N_26857);
or U27371 (N_27371,N_25785,N_25665);
xnor U27372 (N_27372,N_25621,N_26907);
and U27373 (N_27373,N_26643,N_25503);
or U27374 (N_27374,N_26119,N_25511);
and U27375 (N_27375,N_26933,N_26542);
and U27376 (N_27376,N_26884,N_26620);
xor U27377 (N_27377,N_25528,N_26209);
and U27378 (N_27378,N_26300,N_26954);
nand U27379 (N_27379,N_26297,N_26642);
or U27380 (N_27380,N_26080,N_26912);
nor U27381 (N_27381,N_26436,N_25671);
xor U27382 (N_27382,N_26016,N_26647);
nand U27383 (N_27383,N_25813,N_25838);
and U27384 (N_27384,N_26648,N_26321);
or U27385 (N_27385,N_26491,N_26845);
nand U27386 (N_27386,N_26314,N_26423);
and U27387 (N_27387,N_26116,N_26654);
or U27388 (N_27388,N_25620,N_26777);
xnor U27389 (N_27389,N_25518,N_25519);
nand U27390 (N_27390,N_26054,N_25727);
nor U27391 (N_27391,N_25703,N_26661);
nor U27392 (N_27392,N_26143,N_25822);
or U27393 (N_27393,N_26273,N_25660);
nor U27394 (N_27394,N_25593,N_26744);
and U27395 (N_27395,N_26714,N_26239);
and U27396 (N_27396,N_26769,N_26461);
xnor U27397 (N_27397,N_25743,N_26765);
and U27398 (N_27398,N_26854,N_25681);
and U27399 (N_27399,N_26337,N_26683);
nor U27400 (N_27400,N_26587,N_25581);
or U27401 (N_27401,N_25738,N_26749);
or U27402 (N_27402,N_26320,N_25527);
or U27403 (N_27403,N_26374,N_26126);
xor U27404 (N_27404,N_26502,N_26265);
and U27405 (N_27405,N_26074,N_26860);
and U27406 (N_27406,N_26288,N_26403);
nor U27407 (N_27407,N_26707,N_26900);
or U27408 (N_27408,N_26928,N_25735);
nor U27409 (N_27409,N_26095,N_26775);
and U27410 (N_27410,N_26486,N_26419);
or U27411 (N_27411,N_25875,N_26161);
and U27412 (N_27412,N_26633,N_26465);
nor U27413 (N_27413,N_25565,N_25779);
nand U27414 (N_27414,N_25514,N_26115);
or U27415 (N_27415,N_26227,N_26042);
nand U27416 (N_27416,N_26585,N_25733);
and U27417 (N_27417,N_26977,N_26477);
or U27418 (N_27418,N_26047,N_26318);
nor U27419 (N_27419,N_26568,N_25584);
xnor U27420 (N_27420,N_26205,N_25597);
or U27421 (N_27421,N_25972,N_26401);
nor U27422 (N_27422,N_26957,N_26739);
nand U27423 (N_27423,N_26802,N_25651);
or U27424 (N_27424,N_26584,N_26433);
xor U27425 (N_27425,N_25906,N_26776);
nand U27426 (N_27426,N_25782,N_26869);
xnor U27427 (N_27427,N_25645,N_25792);
nor U27428 (N_27428,N_26979,N_26317);
and U27429 (N_27429,N_25534,N_25944);
nand U27430 (N_27430,N_26755,N_25940);
or U27431 (N_27431,N_25719,N_25818);
and U27432 (N_27432,N_26569,N_26684);
xor U27433 (N_27433,N_26327,N_25787);
xor U27434 (N_27434,N_26328,N_26794);
or U27435 (N_27435,N_25993,N_26786);
or U27436 (N_27436,N_26322,N_26524);
xor U27437 (N_27437,N_26917,N_26338);
nor U27438 (N_27438,N_26846,N_26453);
nor U27439 (N_27439,N_26992,N_26268);
or U27440 (N_27440,N_25757,N_26418);
xnor U27441 (N_27441,N_26866,N_26319);
or U27442 (N_27442,N_25970,N_26632);
xnor U27443 (N_27443,N_25802,N_26743);
or U27444 (N_27444,N_26044,N_25980);
nor U27445 (N_27445,N_26371,N_26108);
and U27446 (N_27446,N_26333,N_25835);
xnor U27447 (N_27447,N_25907,N_26967);
xor U27448 (N_27448,N_25543,N_26895);
xor U27449 (N_27449,N_26596,N_25823);
or U27450 (N_27450,N_26941,N_25715);
or U27451 (N_27451,N_25766,N_26351);
or U27452 (N_27452,N_26440,N_26470);
nor U27453 (N_27453,N_26329,N_25873);
nand U27454 (N_27454,N_26036,N_26277);
nor U27455 (N_27455,N_26156,N_25899);
nor U27456 (N_27456,N_26982,N_26285);
xor U27457 (N_27457,N_25674,N_25781);
xnor U27458 (N_27458,N_26228,N_26513);
nor U27459 (N_27459,N_25745,N_25794);
xnor U27460 (N_27460,N_26756,N_25946);
and U27461 (N_27461,N_26035,N_25900);
and U27462 (N_27462,N_25767,N_25726);
nor U27463 (N_27463,N_26864,N_26184);
and U27464 (N_27464,N_26000,N_26349);
nor U27465 (N_27465,N_26720,N_26341);
xor U27466 (N_27466,N_26517,N_25758);
and U27467 (N_27467,N_26157,N_26392);
nand U27468 (N_27468,N_26828,N_26421);
nor U27469 (N_27469,N_25610,N_26516);
and U27470 (N_27470,N_25641,N_25760);
nand U27471 (N_27471,N_26457,N_26753);
nand U27472 (N_27472,N_26736,N_26852);
nor U27473 (N_27473,N_25963,N_26665);
and U27474 (N_27474,N_26411,N_26732);
nand U27475 (N_27475,N_25843,N_25541);
and U27476 (N_27476,N_26867,N_26604);
xor U27477 (N_27477,N_25524,N_26861);
xor U27478 (N_27478,N_26965,N_26163);
and U27479 (N_27479,N_26462,N_25817);
nor U27480 (N_27480,N_26398,N_26464);
nand U27481 (N_27481,N_25577,N_26454);
and U27482 (N_27482,N_25594,N_25834);
xnor U27483 (N_27483,N_26033,N_25694);
or U27484 (N_27484,N_26848,N_26971);
xor U27485 (N_27485,N_25669,N_26911);
xnor U27486 (N_27486,N_25583,N_25841);
xor U27487 (N_27487,N_26629,N_26825);
nand U27488 (N_27488,N_26135,N_26310);
and U27489 (N_27489,N_26987,N_25996);
nand U27490 (N_27490,N_26799,N_26764);
nor U27491 (N_27491,N_26246,N_26637);
nor U27492 (N_27492,N_26215,N_26123);
xnor U27493 (N_27493,N_26206,N_26562);
xor U27494 (N_27494,N_26788,N_25683);
nor U27495 (N_27495,N_26677,N_26856);
nor U27496 (N_27496,N_26508,N_26556);
or U27497 (N_27497,N_25854,N_25941);
or U27498 (N_27498,N_26053,N_25775);
xnor U27499 (N_27499,N_25751,N_25553);
xnor U27500 (N_27500,N_26813,N_26940);
nor U27501 (N_27501,N_26639,N_26106);
nand U27502 (N_27502,N_25537,N_26589);
nand U27503 (N_27503,N_26014,N_25592);
nor U27504 (N_27504,N_26476,N_25851);
and U27505 (N_27505,N_26414,N_26360);
nand U27506 (N_27506,N_26488,N_26621);
nor U27507 (N_27507,N_26305,N_26362);
or U27508 (N_27508,N_26778,N_25997);
nor U27509 (N_27509,N_25713,N_25687);
nor U27510 (N_27510,N_25846,N_25680);
xnor U27511 (N_27511,N_26347,N_25867);
nor U27512 (N_27512,N_26662,N_26795);
nor U27513 (N_27513,N_26039,N_26048);
or U27514 (N_27514,N_25560,N_26208);
xor U27515 (N_27515,N_25604,N_25977);
and U27516 (N_27516,N_26545,N_25585);
and U27517 (N_27517,N_26805,N_26013);
nand U27518 (N_27518,N_25855,N_26279);
xnor U27519 (N_27519,N_26434,N_26512);
or U27520 (N_27520,N_25827,N_26914);
or U27521 (N_27521,N_26689,N_26034);
nand U27522 (N_27522,N_26990,N_26185);
xnor U27523 (N_27523,N_26812,N_26772);
and U27524 (N_27524,N_25718,N_25525);
nand U27525 (N_27525,N_25689,N_26726);
and U27526 (N_27526,N_26079,N_25655);
nor U27527 (N_27527,N_26269,N_26501);
and U27528 (N_27528,N_26051,N_26617);
or U27529 (N_27529,N_25974,N_25825);
or U27530 (N_27530,N_26463,N_25998);
nand U27531 (N_27531,N_26450,N_26431);
or U27532 (N_27532,N_26232,N_25712);
nand U27533 (N_27533,N_26140,N_26355);
nor U27534 (N_27534,N_26873,N_25501);
and U27535 (N_27535,N_26032,N_26557);
nor U27536 (N_27536,N_26540,N_25788);
or U27537 (N_27537,N_25964,N_26479);
nand U27538 (N_27538,N_25704,N_26384);
and U27539 (N_27539,N_25675,N_25634);
and U27540 (N_27540,N_26970,N_26468);
nor U27541 (N_27541,N_25576,N_26306);
xnor U27542 (N_27542,N_25923,N_26791);
xor U27543 (N_27543,N_26537,N_26067);
nor U27544 (N_27544,N_25885,N_26781);
and U27545 (N_27545,N_26644,N_26811);
nand U27546 (N_27546,N_26136,N_25603);
and U27547 (N_27547,N_26110,N_26888);
or U27548 (N_27548,N_26507,N_25772);
and U27549 (N_27549,N_26425,N_26656);
and U27550 (N_27550,N_25754,N_25943);
xnor U27551 (N_27551,N_25879,N_25831);
xor U27552 (N_27552,N_25520,N_26498);
nor U27553 (N_27553,N_25844,N_26024);
xor U27554 (N_27554,N_26417,N_26372);
nand U27555 (N_27555,N_25563,N_26175);
nand U27556 (N_27556,N_26244,N_26831);
nand U27557 (N_27557,N_26704,N_26230);
xor U27558 (N_27558,N_26823,N_25691);
xor U27559 (N_27559,N_26716,N_26495);
nor U27560 (N_27560,N_26681,N_26935);
xnor U27561 (N_27561,N_25642,N_26152);
xnor U27562 (N_27562,N_26274,N_25512);
xnor U27563 (N_27563,N_26021,N_26370);
and U27564 (N_27564,N_25842,N_26170);
nor U27565 (N_27565,N_26134,N_26104);
xnor U27566 (N_27566,N_26820,N_26599);
or U27567 (N_27567,N_26485,N_25605);
nor U27568 (N_27568,N_26824,N_26158);
nor U27569 (N_27569,N_26595,N_26784);
or U27570 (N_27570,N_25917,N_26186);
or U27571 (N_27571,N_25564,N_25742);
nor U27572 (N_27572,N_26729,N_25934);
or U27573 (N_27573,N_26242,N_26946);
or U27574 (N_27574,N_26667,N_25588);
nor U27575 (N_27575,N_26876,N_25568);
xnor U27576 (N_27576,N_25924,N_26473);
nand U27577 (N_27577,N_26748,N_25540);
or U27578 (N_27578,N_26195,N_26630);
nand U27579 (N_27579,N_25849,N_26896);
xor U27580 (N_27580,N_26029,N_26092);
xor U27581 (N_27581,N_25786,N_25979);
and U27582 (N_27582,N_26070,N_26960);
xor U27583 (N_27583,N_25702,N_26177);
nand U27584 (N_27584,N_26061,N_26754);
nor U27585 (N_27585,N_26441,N_25626);
or U27586 (N_27586,N_26234,N_25894);
and U27587 (N_27587,N_26377,N_25990);
nor U27588 (N_27588,N_26006,N_25888);
nand U27589 (N_27589,N_26309,N_25572);
nor U27590 (N_27590,N_26064,N_26702);
nor U27591 (N_27591,N_25956,N_26863);
xnor U27592 (N_27592,N_26541,N_26598);
or U27593 (N_27593,N_25942,N_26505);
and U27594 (N_27594,N_25928,N_25744);
or U27595 (N_27595,N_26410,N_25969);
and U27596 (N_27596,N_26872,N_25740);
nor U27597 (N_27597,N_25695,N_26263);
nand U27598 (N_27598,N_26581,N_26180);
nand U27599 (N_27599,N_26609,N_26149);
or U27600 (N_27600,N_26829,N_25539);
xnor U27601 (N_27601,N_26380,N_25700);
or U27602 (N_27602,N_26922,N_26938);
nor U27603 (N_27603,N_26471,N_25801);
and U27604 (N_27604,N_25557,N_26385);
and U27605 (N_27605,N_25663,N_26045);
xor U27606 (N_27606,N_25510,N_26573);
nor U27607 (N_27607,N_25960,N_26844);
or U27608 (N_27608,N_26606,N_25607);
xor U27609 (N_27609,N_25830,N_25762);
nand U27610 (N_27610,N_26348,N_26789);
xor U27611 (N_27611,N_25967,N_26413);
and U27612 (N_27612,N_26391,N_26574);
and U27613 (N_27613,N_26260,N_25989);
xnor U27614 (N_27614,N_26368,N_25799);
or U27615 (N_27615,N_26272,N_26050);
or U27616 (N_27616,N_26858,N_26925);
nand U27617 (N_27617,N_25898,N_26144);
or U27618 (N_27618,N_25949,N_25562);
nor U27619 (N_27619,N_25720,N_26577);
and U27620 (N_27620,N_26827,N_25601);
nor U27621 (N_27621,N_26354,N_26291);
and U27622 (N_27622,N_26304,N_25776);
xnor U27623 (N_27623,N_26522,N_26275);
xnor U27624 (N_27624,N_26326,N_26302);
xor U27625 (N_27625,N_26251,N_25550);
and U27626 (N_27626,N_26746,N_26171);
and U27627 (N_27627,N_26125,N_26894);
nor U27628 (N_27628,N_25950,N_26671);
or U27629 (N_27629,N_26256,N_25868);
or U27630 (N_27630,N_25931,N_26622);
or U27631 (N_27631,N_25662,N_26796);
and U27632 (N_27632,N_26530,N_26782);
nand U27633 (N_27633,N_26241,N_26738);
nor U27634 (N_27634,N_26017,N_26352);
and U27635 (N_27635,N_26817,N_25633);
or U27636 (N_27636,N_26614,N_26539);
nand U27637 (N_27637,N_25609,N_26745);
nand U27638 (N_27638,N_26426,N_26651);
xnor U27639 (N_27639,N_25716,N_26841);
and U27640 (N_27640,N_26763,N_25994);
xnor U27641 (N_27641,N_25529,N_26919);
xor U27642 (N_27642,N_26201,N_26020);
nand U27643 (N_27643,N_26128,N_26259);
nand U27644 (N_27644,N_25542,N_26725);
xor U27645 (N_27645,N_26664,N_25933);
or U27646 (N_27646,N_26892,N_26071);
and U27647 (N_27647,N_25988,N_26708);
nand U27648 (N_27648,N_26567,N_25891);
or U27649 (N_27649,N_26712,N_26580);
nor U27650 (N_27650,N_25725,N_26118);
xor U27651 (N_27651,N_26698,N_26882);
or U27652 (N_27652,N_25714,N_26217);
xnor U27653 (N_27653,N_25791,N_25780);
and U27654 (N_27654,N_26399,N_26237);
nor U27655 (N_27655,N_25580,N_26284);
nand U27656 (N_27656,N_25856,N_25574);
or U27657 (N_27657,N_25502,N_26536);
and U27658 (N_27658,N_25535,N_26469);
nor U27659 (N_27659,N_25628,N_26307);
xnor U27660 (N_27660,N_26221,N_25747);
or U27661 (N_27661,N_25728,N_26534);
or U27662 (N_27662,N_26945,N_26847);
and U27663 (N_27663,N_26840,N_26626);
nand U27664 (N_27664,N_26083,N_26028);
and U27665 (N_27665,N_25837,N_25882);
and U27666 (N_27666,N_25638,N_26107);
nand U27667 (N_27667,N_26566,N_26586);
and U27668 (N_27668,N_26334,N_26715);
nor U27669 (N_27669,N_26920,N_26364);
xnor U27670 (N_27670,N_25826,N_25839);
and U27671 (N_27671,N_25755,N_26806);
nand U27672 (N_27672,N_26393,N_25505);
xor U27673 (N_27673,N_26443,N_25652);
xnor U27674 (N_27674,N_25533,N_25810);
nor U27675 (N_27675,N_26459,N_26293);
nand U27676 (N_27676,N_26966,N_26214);
or U27677 (N_27677,N_25893,N_26389);
xor U27678 (N_27678,N_26688,N_26478);
and U27679 (N_27679,N_25554,N_25734);
nand U27680 (N_27680,N_26594,N_25981);
nand U27681 (N_27681,N_26086,N_26985);
nand U27682 (N_27682,N_25892,N_25919);
and U27683 (N_27683,N_26964,N_25752);
nor U27684 (N_27684,N_26547,N_25656);
nor U27685 (N_27685,N_25784,N_25804);
nand U27686 (N_27686,N_26591,N_25587);
xnor U27687 (N_27687,N_25650,N_26335);
nand U27688 (N_27688,N_25878,N_25904);
and U27689 (N_27689,N_25630,N_25895);
and U27690 (N_27690,N_26003,N_25793);
nand U27691 (N_27691,N_26225,N_26619);
and U27692 (N_27692,N_26102,N_25739);
nand U27693 (N_27693,N_26908,N_26189);
nor U27694 (N_27694,N_26685,N_25773);
nor U27695 (N_27695,N_26422,N_25961);
or U27696 (N_27696,N_26533,N_25732);
xnor U27697 (N_27697,N_25589,N_25707);
nor U27698 (N_27698,N_26267,N_25705);
xnor U27699 (N_27699,N_26467,N_25613);
or U27700 (N_27700,N_26282,N_25696);
nor U27701 (N_27701,N_25595,N_26850);
nor U27702 (N_27702,N_26998,N_26719);
nand U27703 (N_27703,N_26480,N_25668);
xnor U27704 (N_27704,N_26652,N_26521);
xor U27705 (N_27705,N_26909,N_25623);
xnor U27706 (N_27706,N_26078,N_26717);
xor U27707 (N_27707,N_26375,N_26666);
and U27708 (N_27708,N_26176,N_26299);
or U27709 (N_27709,N_26525,N_25764);
xor U27710 (N_27710,N_26395,N_25544);
or U27711 (N_27711,N_26768,N_26835);
and U27712 (N_27712,N_25803,N_26936);
or U27713 (N_27713,N_26673,N_26109);
xor U27714 (N_27714,N_26564,N_25886);
nor U27715 (N_27715,N_26141,N_25778);
nand U27716 (N_27716,N_25769,N_26901);
nor U27717 (N_27717,N_25927,N_26084);
xor U27718 (N_27718,N_26839,N_26148);
nand U27719 (N_27719,N_26137,N_26339);
and U27720 (N_27720,N_26878,N_25721);
and U27721 (N_27721,N_26575,N_26336);
and U27722 (N_27722,N_26797,N_26819);
or U27723 (N_27723,N_26402,N_26886);
and U27724 (N_27724,N_25807,N_26910);
xor U27725 (N_27725,N_25995,N_26842);
and U27726 (N_27726,N_25682,N_26224);
or U27727 (N_27727,N_25870,N_26994);
and U27728 (N_27728,N_26676,N_25538);
nand U27729 (N_27729,N_26759,N_25800);
and U27730 (N_27730,N_26261,N_26734);
and U27731 (N_27731,N_26166,N_25578);
nor U27732 (N_27732,N_26808,N_25938);
and U27733 (N_27733,N_25561,N_26172);
and U27734 (N_27734,N_26040,N_26271);
and U27735 (N_27735,N_25912,N_26281);
nand U27736 (N_27736,N_26164,N_25730);
or U27737 (N_27737,N_26262,N_26296);
and U27738 (N_27738,N_25746,N_25866);
nand U27739 (N_27739,N_26700,N_26056);
xor U27740 (N_27740,N_25829,N_26280);
nor U27741 (N_27741,N_25558,N_25522);
nor U27742 (N_27742,N_26879,N_26641);
nor U27743 (N_27743,N_26659,N_26742);
nor U27744 (N_27744,N_26011,N_26783);
or U27745 (N_27745,N_26169,N_25816);
or U27746 (N_27746,N_26409,N_26038);
or U27747 (N_27747,N_26590,N_25955);
xor U27748 (N_27748,N_25523,N_25654);
and U27749 (N_27749,N_26515,N_25647);
nor U27750 (N_27750,N_26505,N_25701);
xnor U27751 (N_27751,N_25760,N_26193);
or U27752 (N_27752,N_25744,N_25808);
xor U27753 (N_27753,N_26908,N_25787);
xnor U27754 (N_27754,N_26003,N_25898);
and U27755 (N_27755,N_26072,N_25861);
nor U27756 (N_27756,N_26817,N_26153);
and U27757 (N_27757,N_26219,N_25726);
xor U27758 (N_27758,N_26016,N_25848);
xnor U27759 (N_27759,N_26491,N_26945);
nor U27760 (N_27760,N_25646,N_25591);
or U27761 (N_27761,N_26099,N_25710);
nor U27762 (N_27762,N_25548,N_26671);
and U27763 (N_27763,N_26933,N_26848);
nand U27764 (N_27764,N_26643,N_26971);
nor U27765 (N_27765,N_25624,N_26812);
nor U27766 (N_27766,N_26009,N_26239);
and U27767 (N_27767,N_26944,N_25629);
xnor U27768 (N_27768,N_26915,N_26504);
and U27769 (N_27769,N_26839,N_26084);
xnor U27770 (N_27770,N_26889,N_25997);
or U27771 (N_27771,N_25924,N_25845);
nand U27772 (N_27772,N_26412,N_26479);
and U27773 (N_27773,N_26139,N_26622);
or U27774 (N_27774,N_26970,N_26650);
and U27775 (N_27775,N_26934,N_26253);
nand U27776 (N_27776,N_26749,N_26411);
nor U27777 (N_27777,N_26976,N_26938);
nand U27778 (N_27778,N_26125,N_25716);
or U27779 (N_27779,N_25718,N_26132);
and U27780 (N_27780,N_26905,N_26616);
and U27781 (N_27781,N_26031,N_26760);
nor U27782 (N_27782,N_25711,N_25796);
nand U27783 (N_27783,N_25738,N_25714);
and U27784 (N_27784,N_26276,N_26903);
nor U27785 (N_27785,N_25522,N_26407);
or U27786 (N_27786,N_26610,N_26775);
or U27787 (N_27787,N_26831,N_25811);
and U27788 (N_27788,N_26577,N_26075);
xor U27789 (N_27789,N_25549,N_25942);
nor U27790 (N_27790,N_25986,N_25780);
nand U27791 (N_27791,N_26606,N_26436);
or U27792 (N_27792,N_25746,N_26305);
nor U27793 (N_27793,N_26447,N_26491);
xor U27794 (N_27794,N_26115,N_25812);
nor U27795 (N_27795,N_26655,N_26523);
and U27796 (N_27796,N_26943,N_26098);
and U27797 (N_27797,N_25588,N_25615);
or U27798 (N_27798,N_25681,N_26455);
and U27799 (N_27799,N_26573,N_26413);
xor U27800 (N_27800,N_26543,N_26366);
xnor U27801 (N_27801,N_26826,N_26434);
or U27802 (N_27802,N_26236,N_26829);
nand U27803 (N_27803,N_25728,N_26980);
or U27804 (N_27804,N_26453,N_26620);
xor U27805 (N_27805,N_25642,N_26180);
and U27806 (N_27806,N_26771,N_26611);
or U27807 (N_27807,N_25701,N_26160);
nand U27808 (N_27808,N_26353,N_26267);
xnor U27809 (N_27809,N_25923,N_25507);
nand U27810 (N_27810,N_26389,N_26162);
and U27811 (N_27811,N_25774,N_25691);
xnor U27812 (N_27812,N_26861,N_26209);
xor U27813 (N_27813,N_26493,N_25715);
xor U27814 (N_27814,N_25708,N_25787);
nor U27815 (N_27815,N_26290,N_25978);
xnor U27816 (N_27816,N_26100,N_26339);
or U27817 (N_27817,N_26431,N_26713);
nand U27818 (N_27818,N_25551,N_26456);
and U27819 (N_27819,N_26447,N_26831);
nor U27820 (N_27820,N_25585,N_26747);
and U27821 (N_27821,N_26968,N_26853);
xnor U27822 (N_27822,N_26311,N_25570);
or U27823 (N_27823,N_25628,N_26975);
xor U27824 (N_27824,N_26235,N_26367);
or U27825 (N_27825,N_26003,N_26185);
or U27826 (N_27826,N_26170,N_26952);
or U27827 (N_27827,N_26640,N_26495);
or U27828 (N_27828,N_25806,N_26932);
xnor U27829 (N_27829,N_25911,N_25800);
nor U27830 (N_27830,N_26428,N_26731);
nor U27831 (N_27831,N_26397,N_26185);
nor U27832 (N_27832,N_26068,N_26911);
and U27833 (N_27833,N_25564,N_26216);
xor U27834 (N_27834,N_26349,N_25967);
nor U27835 (N_27835,N_26055,N_26635);
nand U27836 (N_27836,N_26301,N_25532);
nor U27837 (N_27837,N_25689,N_25799);
xnor U27838 (N_27838,N_26809,N_26707);
nor U27839 (N_27839,N_26646,N_26628);
nand U27840 (N_27840,N_26208,N_26333);
nand U27841 (N_27841,N_26229,N_25763);
or U27842 (N_27842,N_26062,N_25963);
xnor U27843 (N_27843,N_25781,N_26405);
nand U27844 (N_27844,N_25653,N_25503);
nand U27845 (N_27845,N_26173,N_25502);
and U27846 (N_27846,N_25957,N_26600);
nor U27847 (N_27847,N_25724,N_25599);
xnor U27848 (N_27848,N_25765,N_25869);
nor U27849 (N_27849,N_25696,N_25930);
xor U27850 (N_27850,N_26405,N_26461);
nor U27851 (N_27851,N_26412,N_26106);
and U27852 (N_27852,N_26468,N_26718);
nand U27853 (N_27853,N_26775,N_26969);
nand U27854 (N_27854,N_25834,N_26744);
or U27855 (N_27855,N_26989,N_26591);
nand U27856 (N_27856,N_26746,N_26884);
nor U27857 (N_27857,N_25889,N_26759);
nand U27858 (N_27858,N_26330,N_26545);
and U27859 (N_27859,N_25876,N_25734);
nor U27860 (N_27860,N_26876,N_26218);
nand U27861 (N_27861,N_26682,N_26236);
and U27862 (N_27862,N_25809,N_26138);
nor U27863 (N_27863,N_25572,N_25767);
xor U27864 (N_27864,N_26952,N_26241);
xor U27865 (N_27865,N_26431,N_25800);
or U27866 (N_27866,N_26457,N_25848);
xnor U27867 (N_27867,N_25989,N_26181);
or U27868 (N_27868,N_26354,N_25727);
and U27869 (N_27869,N_25535,N_26697);
xnor U27870 (N_27870,N_25863,N_25518);
or U27871 (N_27871,N_26022,N_25532);
nor U27872 (N_27872,N_26642,N_26380);
or U27873 (N_27873,N_25639,N_26348);
xnor U27874 (N_27874,N_25773,N_26509);
or U27875 (N_27875,N_26287,N_25728);
nor U27876 (N_27876,N_26515,N_26070);
nand U27877 (N_27877,N_26665,N_25604);
nor U27878 (N_27878,N_26593,N_26898);
nand U27879 (N_27879,N_26034,N_26332);
nor U27880 (N_27880,N_26391,N_25866);
and U27881 (N_27881,N_26404,N_26330);
xnor U27882 (N_27882,N_26299,N_25511);
xor U27883 (N_27883,N_25501,N_25843);
xnor U27884 (N_27884,N_26429,N_26582);
and U27885 (N_27885,N_26697,N_26532);
xnor U27886 (N_27886,N_26792,N_26208);
or U27887 (N_27887,N_26176,N_26283);
nand U27888 (N_27888,N_26270,N_26762);
nand U27889 (N_27889,N_25976,N_25716);
xor U27890 (N_27890,N_25535,N_26625);
nand U27891 (N_27891,N_26468,N_25755);
or U27892 (N_27892,N_26630,N_25731);
nand U27893 (N_27893,N_25592,N_25743);
or U27894 (N_27894,N_26493,N_26269);
and U27895 (N_27895,N_25720,N_26298);
or U27896 (N_27896,N_26070,N_25925);
and U27897 (N_27897,N_26260,N_26041);
xnor U27898 (N_27898,N_26259,N_26795);
and U27899 (N_27899,N_26658,N_26627);
nor U27900 (N_27900,N_26874,N_26705);
or U27901 (N_27901,N_26106,N_26710);
xor U27902 (N_27902,N_26318,N_26526);
or U27903 (N_27903,N_26248,N_25514);
or U27904 (N_27904,N_26220,N_26485);
or U27905 (N_27905,N_25927,N_26594);
nor U27906 (N_27906,N_25841,N_25721);
and U27907 (N_27907,N_26305,N_26871);
nor U27908 (N_27908,N_26159,N_26327);
or U27909 (N_27909,N_25904,N_25608);
or U27910 (N_27910,N_25762,N_25563);
or U27911 (N_27911,N_26241,N_26985);
nand U27912 (N_27912,N_25695,N_25646);
and U27913 (N_27913,N_26539,N_25926);
xnor U27914 (N_27914,N_25687,N_26610);
and U27915 (N_27915,N_25986,N_26603);
nand U27916 (N_27916,N_26654,N_26569);
and U27917 (N_27917,N_25659,N_26500);
xnor U27918 (N_27918,N_25615,N_25772);
nor U27919 (N_27919,N_26411,N_26628);
nand U27920 (N_27920,N_26185,N_25726);
or U27921 (N_27921,N_25786,N_26777);
xnor U27922 (N_27922,N_26572,N_26010);
nor U27923 (N_27923,N_26199,N_25686);
nand U27924 (N_27924,N_26212,N_25865);
or U27925 (N_27925,N_26592,N_25953);
and U27926 (N_27926,N_25949,N_26339);
nor U27927 (N_27927,N_26187,N_26817);
and U27928 (N_27928,N_26595,N_26989);
and U27929 (N_27929,N_26176,N_26545);
nand U27930 (N_27930,N_26900,N_25545);
xor U27931 (N_27931,N_26982,N_26739);
and U27932 (N_27932,N_26846,N_26700);
or U27933 (N_27933,N_26548,N_25527);
nand U27934 (N_27934,N_26391,N_25920);
nand U27935 (N_27935,N_26350,N_26233);
nor U27936 (N_27936,N_25792,N_26424);
or U27937 (N_27937,N_26487,N_26927);
or U27938 (N_27938,N_26954,N_26620);
or U27939 (N_27939,N_26235,N_25569);
xor U27940 (N_27940,N_25976,N_26246);
nor U27941 (N_27941,N_26187,N_25656);
or U27942 (N_27942,N_26461,N_25696);
and U27943 (N_27943,N_26737,N_26180);
nor U27944 (N_27944,N_26344,N_26304);
nor U27945 (N_27945,N_26818,N_26691);
or U27946 (N_27946,N_26312,N_25997);
nand U27947 (N_27947,N_26605,N_25520);
nand U27948 (N_27948,N_25925,N_25971);
xor U27949 (N_27949,N_26223,N_26851);
or U27950 (N_27950,N_26803,N_26400);
nor U27951 (N_27951,N_25701,N_26434);
xor U27952 (N_27952,N_26222,N_26025);
nand U27953 (N_27953,N_25592,N_26844);
nand U27954 (N_27954,N_25559,N_26465);
nand U27955 (N_27955,N_26522,N_25842);
or U27956 (N_27956,N_26866,N_26448);
nor U27957 (N_27957,N_26445,N_26926);
nor U27958 (N_27958,N_25874,N_25821);
nor U27959 (N_27959,N_26990,N_25765);
xor U27960 (N_27960,N_26375,N_26685);
nand U27961 (N_27961,N_26040,N_26385);
nand U27962 (N_27962,N_26827,N_26768);
or U27963 (N_27963,N_26967,N_25965);
and U27964 (N_27964,N_26669,N_26301);
nand U27965 (N_27965,N_26687,N_25847);
or U27966 (N_27966,N_26625,N_26569);
nor U27967 (N_27967,N_25587,N_25988);
or U27968 (N_27968,N_25503,N_26642);
xnor U27969 (N_27969,N_26465,N_26258);
nor U27970 (N_27970,N_26293,N_26774);
xor U27971 (N_27971,N_25527,N_26985);
xnor U27972 (N_27972,N_26716,N_25967);
xnor U27973 (N_27973,N_26814,N_25944);
nor U27974 (N_27974,N_26068,N_25752);
nand U27975 (N_27975,N_26144,N_26599);
and U27976 (N_27976,N_26949,N_25824);
or U27977 (N_27977,N_26943,N_26857);
xnor U27978 (N_27978,N_26586,N_26820);
or U27979 (N_27979,N_26696,N_25509);
nor U27980 (N_27980,N_26336,N_26020);
nor U27981 (N_27981,N_26693,N_26964);
nor U27982 (N_27982,N_26955,N_25674);
nand U27983 (N_27983,N_26301,N_26582);
and U27984 (N_27984,N_25582,N_26695);
xor U27985 (N_27985,N_26711,N_26414);
nor U27986 (N_27986,N_26511,N_26071);
and U27987 (N_27987,N_26562,N_26061);
or U27988 (N_27988,N_26514,N_26619);
and U27989 (N_27989,N_25702,N_26296);
nand U27990 (N_27990,N_25540,N_26603);
nand U27991 (N_27991,N_26268,N_26223);
or U27992 (N_27992,N_26287,N_26122);
nor U27993 (N_27993,N_25882,N_26819);
xnor U27994 (N_27994,N_26341,N_26206);
or U27995 (N_27995,N_26328,N_25867);
or U27996 (N_27996,N_26430,N_26275);
xnor U27997 (N_27997,N_26974,N_26433);
nor U27998 (N_27998,N_26665,N_26894);
nand U27999 (N_27999,N_26203,N_26259);
xor U28000 (N_28000,N_26373,N_26711);
nand U28001 (N_28001,N_25879,N_26883);
or U28002 (N_28002,N_26190,N_26278);
or U28003 (N_28003,N_26440,N_26723);
nor U28004 (N_28004,N_26171,N_26106);
xnor U28005 (N_28005,N_26322,N_26351);
nand U28006 (N_28006,N_25552,N_25929);
and U28007 (N_28007,N_26984,N_25817);
nor U28008 (N_28008,N_26777,N_25680);
xor U28009 (N_28009,N_25917,N_26235);
xor U28010 (N_28010,N_26964,N_26477);
and U28011 (N_28011,N_26382,N_26208);
and U28012 (N_28012,N_25980,N_25967);
or U28013 (N_28013,N_26905,N_26877);
nand U28014 (N_28014,N_26260,N_25664);
nor U28015 (N_28015,N_26414,N_26386);
xor U28016 (N_28016,N_26024,N_26284);
and U28017 (N_28017,N_26004,N_26665);
and U28018 (N_28018,N_25709,N_25592);
xor U28019 (N_28019,N_26893,N_26505);
or U28020 (N_28020,N_26498,N_26652);
and U28021 (N_28021,N_25739,N_26252);
xor U28022 (N_28022,N_26708,N_26502);
and U28023 (N_28023,N_26107,N_26052);
or U28024 (N_28024,N_25978,N_25660);
and U28025 (N_28025,N_26265,N_25932);
and U28026 (N_28026,N_26288,N_26967);
or U28027 (N_28027,N_25875,N_25686);
and U28028 (N_28028,N_26441,N_26814);
or U28029 (N_28029,N_26348,N_26801);
or U28030 (N_28030,N_26584,N_26650);
nand U28031 (N_28031,N_26769,N_25558);
and U28032 (N_28032,N_25653,N_25778);
xor U28033 (N_28033,N_26972,N_26961);
nand U28034 (N_28034,N_26690,N_26496);
nand U28035 (N_28035,N_26709,N_25556);
nand U28036 (N_28036,N_26077,N_25880);
or U28037 (N_28037,N_26007,N_25990);
xor U28038 (N_28038,N_25537,N_26634);
nand U28039 (N_28039,N_26975,N_26346);
xor U28040 (N_28040,N_26603,N_26218);
nor U28041 (N_28041,N_25533,N_26567);
nor U28042 (N_28042,N_26906,N_26352);
nand U28043 (N_28043,N_25703,N_26728);
and U28044 (N_28044,N_25529,N_25762);
and U28045 (N_28045,N_26143,N_25596);
nor U28046 (N_28046,N_26391,N_25646);
nand U28047 (N_28047,N_26594,N_26902);
xor U28048 (N_28048,N_26343,N_26898);
nand U28049 (N_28049,N_25668,N_26349);
nand U28050 (N_28050,N_26665,N_26488);
nor U28051 (N_28051,N_25731,N_26974);
or U28052 (N_28052,N_26504,N_26913);
nand U28053 (N_28053,N_25797,N_25623);
nor U28054 (N_28054,N_25926,N_26457);
nand U28055 (N_28055,N_26608,N_25682);
or U28056 (N_28056,N_25636,N_26127);
nor U28057 (N_28057,N_25699,N_25882);
nand U28058 (N_28058,N_25812,N_26040);
nand U28059 (N_28059,N_26410,N_25906);
and U28060 (N_28060,N_26685,N_26757);
nor U28061 (N_28061,N_25884,N_26102);
xor U28062 (N_28062,N_26870,N_26196);
or U28063 (N_28063,N_26839,N_26176);
nor U28064 (N_28064,N_26875,N_26545);
or U28065 (N_28065,N_26340,N_26408);
or U28066 (N_28066,N_25528,N_25818);
nand U28067 (N_28067,N_25534,N_26026);
xor U28068 (N_28068,N_26356,N_26063);
nand U28069 (N_28069,N_25773,N_25691);
nand U28070 (N_28070,N_26495,N_25687);
xor U28071 (N_28071,N_25962,N_26937);
nor U28072 (N_28072,N_25848,N_26973);
or U28073 (N_28073,N_26529,N_26924);
nor U28074 (N_28074,N_25649,N_25892);
xnor U28075 (N_28075,N_26858,N_25568);
nor U28076 (N_28076,N_26250,N_26501);
xnor U28077 (N_28077,N_26623,N_26723);
xor U28078 (N_28078,N_25829,N_26952);
nand U28079 (N_28079,N_26076,N_26970);
or U28080 (N_28080,N_25731,N_25645);
or U28081 (N_28081,N_25700,N_25603);
nand U28082 (N_28082,N_26695,N_26544);
and U28083 (N_28083,N_26476,N_26207);
and U28084 (N_28084,N_25626,N_26882);
or U28085 (N_28085,N_26204,N_26825);
and U28086 (N_28086,N_25683,N_26579);
or U28087 (N_28087,N_26729,N_26213);
nand U28088 (N_28088,N_26942,N_26136);
and U28089 (N_28089,N_25944,N_25916);
xnor U28090 (N_28090,N_26589,N_26166);
xnor U28091 (N_28091,N_26790,N_25813);
xor U28092 (N_28092,N_26547,N_26280);
xnor U28093 (N_28093,N_26629,N_26836);
nand U28094 (N_28094,N_26806,N_26574);
or U28095 (N_28095,N_26659,N_26995);
nor U28096 (N_28096,N_25842,N_25911);
xor U28097 (N_28097,N_26873,N_26916);
nand U28098 (N_28098,N_26231,N_25821);
and U28099 (N_28099,N_25823,N_26969);
nor U28100 (N_28100,N_26102,N_26109);
nand U28101 (N_28101,N_26474,N_26409);
or U28102 (N_28102,N_26615,N_26981);
nand U28103 (N_28103,N_26130,N_26581);
or U28104 (N_28104,N_25916,N_26234);
nor U28105 (N_28105,N_26290,N_26929);
and U28106 (N_28106,N_25549,N_26113);
nor U28107 (N_28107,N_26305,N_26850);
and U28108 (N_28108,N_26080,N_25918);
or U28109 (N_28109,N_26517,N_26144);
xnor U28110 (N_28110,N_26436,N_25693);
or U28111 (N_28111,N_26174,N_25863);
or U28112 (N_28112,N_26626,N_25938);
xnor U28113 (N_28113,N_25972,N_26589);
xor U28114 (N_28114,N_26211,N_26786);
and U28115 (N_28115,N_25597,N_25518);
or U28116 (N_28116,N_26827,N_26589);
and U28117 (N_28117,N_25769,N_25873);
xor U28118 (N_28118,N_26624,N_26471);
nor U28119 (N_28119,N_25892,N_25512);
nand U28120 (N_28120,N_25757,N_26710);
xnor U28121 (N_28121,N_26334,N_26469);
nor U28122 (N_28122,N_25599,N_25896);
xnor U28123 (N_28123,N_26201,N_26788);
nor U28124 (N_28124,N_25725,N_25629);
nand U28125 (N_28125,N_26828,N_26424);
xor U28126 (N_28126,N_25847,N_26194);
xor U28127 (N_28127,N_26358,N_25828);
xor U28128 (N_28128,N_26775,N_25974);
and U28129 (N_28129,N_26579,N_25872);
xnor U28130 (N_28130,N_26921,N_25662);
xnor U28131 (N_28131,N_26608,N_25871);
and U28132 (N_28132,N_26967,N_26954);
or U28133 (N_28133,N_26785,N_26704);
xnor U28134 (N_28134,N_26657,N_25991);
or U28135 (N_28135,N_25972,N_26044);
nand U28136 (N_28136,N_25810,N_26718);
nand U28137 (N_28137,N_25962,N_26716);
xnor U28138 (N_28138,N_26055,N_25925);
xnor U28139 (N_28139,N_26206,N_26094);
nand U28140 (N_28140,N_26351,N_26224);
nor U28141 (N_28141,N_26708,N_26106);
nor U28142 (N_28142,N_26514,N_26006);
nand U28143 (N_28143,N_26924,N_26438);
and U28144 (N_28144,N_26134,N_26519);
or U28145 (N_28145,N_25647,N_25510);
and U28146 (N_28146,N_25517,N_25741);
or U28147 (N_28147,N_26136,N_25821);
and U28148 (N_28148,N_26523,N_26546);
or U28149 (N_28149,N_26269,N_26970);
nand U28150 (N_28150,N_26989,N_26888);
nor U28151 (N_28151,N_25766,N_25514);
and U28152 (N_28152,N_26079,N_26936);
or U28153 (N_28153,N_25958,N_26061);
nor U28154 (N_28154,N_26534,N_25662);
or U28155 (N_28155,N_26617,N_25971);
and U28156 (N_28156,N_26179,N_26382);
and U28157 (N_28157,N_26608,N_26694);
nand U28158 (N_28158,N_26618,N_26283);
xnor U28159 (N_28159,N_26545,N_26094);
or U28160 (N_28160,N_26023,N_26123);
nor U28161 (N_28161,N_26258,N_26598);
nand U28162 (N_28162,N_25671,N_26485);
xnor U28163 (N_28163,N_26588,N_25541);
nor U28164 (N_28164,N_26681,N_25756);
and U28165 (N_28165,N_26244,N_26194);
and U28166 (N_28166,N_26726,N_25719);
or U28167 (N_28167,N_25799,N_26743);
xor U28168 (N_28168,N_26408,N_26506);
nand U28169 (N_28169,N_25977,N_26095);
xnor U28170 (N_28170,N_25920,N_26584);
or U28171 (N_28171,N_25631,N_26460);
nand U28172 (N_28172,N_26000,N_26539);
nand U28173 (N_28173,N_26799,N_26627);
and U28174 (N_28174,N_26813,N_25982);
or U28175 (N_28175,N_26788,N_26052);
or U28176 (N_28176,N_25835,N_26537);
nor U28177 (N_28177,N_26603,N_26876);
and U28178 (N_28178,N_25637,N_26868);
nand U28179 (N_28179,N_25699,N_25737);
or U28180 (N_28180,N_26367,N_26968);
or U28181 (N_28181,N_26026,N_25517);
nand U28182 (N_28182,N_26463,N_26260);
nor U28183 (N_28183,N_26057,N_25624);
and U28184 (N_28184,N_25654,N_25653);
nand U28185 (N_28185,N_25739,N_26977);
and U28186 (N_28186,N_26081,N_25870);
xnor U28187 (N_28187,N_26370,N_26362);
xnor U28188 (N_28188,N_26728,N_25643);
xnor U28189 (N_28189,N_26716,N_26348);
or U28190 (N_28190,N_26007,N_25988);
or U28191 (N_28191,N_26524,N_26362);
xnor U28192 (N_28192,N_26048,N_26736);
nor U28193 (N_28193,N_26066,N_26907);
xor U28194 (N_28194,N_26401,N_26947);
and U28195 (N_28195,N_26162,N_26704);
nand U28196 (N_28196,N_25842,N_26639);
nand U28197 (N_28197,N_26351,N_25807);
and U28198 (N_28198,N_26270,N_26925);
xor U28199 (N_28199,N_26924,N_26074);
nand U28200 (N_28200,N_26655,N_26882);
xor U28201 (N_28201,N_25564,N_25846);
nor U28202 (N_28202,N_25505,N_26863);
nand U28203 (N_28203,N_26687,N_26902);
nand U28204 (N_28204,N_26128,N_26075);
and U28205 (N_28205,N_26601,N_25924);
xor U28206 (N_28206,N_26683,N_25651);
and U28207 (N_28207,N_26709,N_26446);
nand U28208 (N_28208,N_25956,N_26393);
nand U28209 (N_28209,N_26071,N_25903);
nor U28210 (N_28210,N_26722,N_25688);
nor U28211 (N_28211,N_25992,N_26105);
and U28212 (N_28212,N_25727,N_26832);
nor U28213 (N_28213,N_26696,N_25836);
nor U28214 (N_28214,N_25743,N_26776);
nand U28215 (N_28215,N_26031,N_26114);
xor U28216 (N_28216,N_25779,N_26070);
xnor U28217 (N_28217,N_25543,N_26611);
nor U28218 (N_28218,N_26522,N_26663);
and U28219 (N_28219,N_25601,N_26709);
nand U28220 (N_28220,N_25813,N_25904);
xor U28221 (N_28221,N_25684,N_25590);
and U28222 (N_28222,N_25880,N_26430);
or U28223 (N_28223,N_25921,N_26366);
nor U28224 (N_28224,N_25605,N_26102);
or U28225 (N_28225,N_25838,N_25979);
nand U28226 (N_28226,N_26080,N_25683);
nor U28227 (N_28227,N_25537,N_26712);
xnor U28228 (N_28228,N_26455,N_25575);
xnor U28229 (N_28229,N_25616,N_25570);
and U28230 (N_28230,N_25975,N_25939);
nor U28231 (N_28231,N_26018,N_26952);
nand U28232 (N_28232,N_26954,N_26154);
xor U28233 (N_28233,N_25605,N_26462);
xor U28234 (N_28234,N_26586,N_26778);
and U28235 (N_28235,N_26129,N_26430);
xnor U28236 (N_28236,N_26082,N_25813);
nand U28237 (N_28237,N_25812,N_26187);
nor U28238 (N_28238,N_25817,N_26271);
nor U28239 (N_28239,N_26117,N_26960);
nand U28240 (N_28240,N_26607,N_26681);
or U28241 (N_28241,N_25828,N_26765);
and U28242 (N_28242,N_25698,N_26000);
nor U28243 (N_28243,N_25665,N_26701);
or U28244 (N_28244,N_25743,N_25508);
nor U28245 (N_28245,N_26989,N_25724);
xnor U28246 (N_28246,N_26132,N_26054);
and U28247 (N_28247,N_26866,N_26246);
and U28248 (N_28248,N_26386,N_26131);
nand U28249 (N_28249,N_26218,N_26746);
xnor U28250 (N_28250,N_26598,N_26375);
or U28251 (N_28251,N_26489,N_26078);
or U28252 (N_28252,N_26273,N_26507);
xor U28253 (N_28253,N_26810,N_25849);
and U28254 (N_28254,N_26464,N_26107);
nor U28255 (N_28255,N_26033,N_26189);
or U28256 (N_28256,N_25675,N_26600);
nand U28257 (N_28257,N_26274,N_26106);
xnor U28258 (N_28258,N_26606,N_25659);
and U28259 (N_28259,N_26534,N_25797);
or U28260 (N_28260,N_26499,N_26318);
and U28261 (N_28261,N_25697,N_26241);
and U28262 (N_28262,N_25942,N_26957);
or U28263 (N_28263,N_25701,N_26295);
nand U28264 (N_28264,N_25565,N_26813);
xor U28265 (N_28265,N_26194,N_26054);
xnor U28266 (N_28266,N_25711,N_25841);
nor U28267 (N_28267,N_26261,N_26334);
xnor U28268 (N_28268,N_26660,N_26844);
and U28269 (N_28269,N_25985,N_26843);
and U28270 (N_28270,N_26240,N_25950);
xor U28271 (N_28271,N_26757,N_26017);
xor U28272 (N_28272,N_26714,N_26340);
nor U28273 (N_28273,N_25919,N_26329);
nand U28274 (N_28274,N_26730,N_26734);
xnor U28275 (N_28275,N_26822,N_25964);
or U28276 (N_28276,N_26380,N_26439);
nor U28277 (N_28277,N_26314,N_26248);
nand U28278 (N_28278,N_26180,N_26990);
xnor U28279 (N_28279,N_26248,N_25980);
nor U28280 (N_28280,N_26575,N_26393);
or U28281 (N_28281,N_26798,N_26310);
nand U28282 (N_28282,N_26462,N_25636);
or U28283 (N_28283,N_26113,N_26691);
and U28284 (N_28284,N_26277,N_26395);
nor U28285 (N_28285,N_26323,N_26952);
or U28286 (N_28286,N_26540,N_26085);
nor U28287 (N_28287,N_25642,N_26615);
nor U28288 (N_28288,N_26246,N_26964);
xor U28289 (N_28289,N_25619,N_26652);
or U28290 (N_28290,N_26638,N_25640);
nand U28291 (N_28291,N_25792,N_25994);
or U28292 (N_28292,N_26236,N_26445);
xnor U28293 (N_28293,N_26527,N_25747);
nor U28294 (N_28294,N_25539,N_26266);
nand U28295 (N_28295,N_26474,N_26576);
nand U28296 (N_28296,N_26318,N_26517);
or U28297 (N_28297,N_26658,N_25526);
and U28298 (N_28298,N_26975,N_26377);
or U28299 (N_28299,N_25796,N_25534);
nand U28300 (N_28300,N_26968,N_26783);
and U28301 (N_28301,N_25920,N_26842);
nand U28302 (N_28302,N_26139,N_25797);
nor U28303 (N_28303,N_26829,N_26170);
and U28304 (N_28304,N_26682,N_26683);
or U28305 (N_28305,N_25895,N_25891);
and U28306 (N_28306,N_26478,N_26547);
nor U28307 (N_28307,N_26792,N_25899);
or U28308 (N_28308,N_25767,N_26339);
nor U28309 (N_28309,N_25748,N_26052);
nand U28310 (N_28310,N_25927,N_26003);
nor U28311 (N_28311,N_26853,N_26050);
and U28312 (N_28312,N_26783,N_26622);
xor U28313 (N_28313,N_26774,N_26147);
and U28314 (N_28314,N_26946,N_26377);
nand U28315 (N_28315,N_26957,N_26762);
nor U28316 (N_28316,N_26587,N_26950);
nor U28317 (N_28317,N_25991,N_26291);
nand U28318 (N_28318,N_26598,N_26102);
xnor U28319 (N_28319,N_26804,N_25582);
and U28320 (N_28320,N_26390,N_26847);
nand U28321 (N_28321,N_26157,N_26918);
nand U28322 (N_28322,N_25668,N_26873);
xor U28323 (N_28323,N_25525,N_26513);
or U28324 (N_28324,N_25937,N_25673);
nor U28325 (N_28325,N_26971,N_25713);
nor U28326 (N_28326,N_26105,N_26777);
nand U28327 (N_28327,N_26341,N_26316);
nor U28328 (N_28328,N_25617,N_25710);
and U28329 (N_28329,N_26598,N_26487);
xnor U28330 (N_28330,N_25752,N_26719);
nor U28331 (N_28331,N_26674,N_25993);
nand U28332 (N_28332,N_26047,N_25546);
and U28333 (N_28333,N_25829,N_26730);
or U28334 (N_28334,N_25674,N_25876);
or U28335 (N_28335,N_26632,N_26965);
xor U28336 (N_28336,N_26861,N_26172);
nand U28337 (N_28337,N_25823,N_26801);
nor U28338 (N_28338,N_26163,N_26640);
or U28339 (N_28339,N_26072,N_25713);
or U28340 (N_28340,N_26774,N_25971);
nand U28341 (N_28341,N_26957,N_26267);
or U28342 (N_28342,N_26539,N_26408);
xnor U28343 (N_28343,N_25744,N_25876);
nor U28344 (N_28344,N_25780,N_26298);
nand U28345 (N_28345,N_26532,N_26900);
or U28346 (N_28346,N_26438,N_26774);
xnor U28347 (N_28347,N_26359,N_25914);
or U28348 (N_28348,N_26798,N_25926);
nor U28349 (N_28349,N_26403,N_26600);
or U28350 (N_28350,N_25854,N_26185);
or U28351 (N_28351,N_26678,N_26357);
or U28352 (N_28352,N_26038,N_25946);
or U28353 (N_28353,N_25772,N_26064);
nor U28354 (N_28354,N_26192,N_26720);
xor U28355 (N_28355,N_25727,N_25930);
and U28356 (N_28356,N_25719,N_26704);
or U28357 (N_28357,N_26312,N_26154);
nor U28358 (N_28358,N_25617,N_26923);
xor U28359 (N_28359,N_26468,N_26061);
nor U28360 (N_28360,N_25931,N_26593);
and U28361 (N_28361,N_26025,N_25758);
xor U28362 (N_28362,N_26892,N_25855);
nand U28363 (N_28363,N_25551,N_26443);
xnor U28364 (N_28364,N_26917,N_26972);
nand U28365 (N_28365,N_26580,N_25516);
xor U28366 (N_28366,N_26571,N_26584);
xor U28367 (N_28367,N_26169,N_25922);
nor U28368 (N_28368,N_26476,N_26618);
and U28369 (N_28369,N_26876,N_26007);
or U28370 (N_28370,N_25866,N_25735);
nor U28371 (N_28371,N_26464,N_26629);
xor U28372 (N_28372,N_25665,N_25606);
nand U28373 (N_28373,N_26547,N_26796);
or U28374 (N_28374,N_26670,N_26363);
xnor U28375 (N_28375,N_25854,N_25572);
nor U28376 (N_28376,N_25995,N_25938);
or U28377 (N_28377,N_26258,N_25526);
xor U28378 (N_28378,N_26615,N_25855);
nand U28379 (N_28379,N_26735,N_26801);
nor U28380 (N_28380,N_26948,N_26435);
or U28381 (N_28381,N_26337,N_26966);
nand U28382 (N_28382,N_26179,N_26146);
and U28383 (N_28383,N_26430,N_26972);
nand U28384 (N_28384,N_26509,N_26462);
and U28385 (N_28385,N_25972,N_26498);
and U28386 (N_28386,N_25830,N_26622);
and U28387 (N_28387,N_26015,N_26161);
and U28388 (N_28388,N_25772,N_25791);
and U28389 (N_28389,N_25791,N_26669);
and U28390 (N_28390,N_25748,N_25808);
or U28391 (N_28391,N_25632,N_26822);
or U28392 (N_28392,N_25793,N_25930);
xnor U28393 (N_28393,N_25626,N_26179);
xnor U28394 (N_28394,N_26192,N_26583);
xnor U28395 (N_28395,N_25985,N_25691);
nand U28396 (N_28396,N_26627,N_25750);
and U28397 (N_28397,N_25614,N_26132);
xnor U28398 (N_28398,N_26937,N_26457);
xnor U28399 (N_28399,N_26502,N_26445);
and U28400 (N_28400,N_25884,N_26330);
nor U28401 (N_28401,N_25950,N_25931);
nand U28402 (N_28402,N_25997,N_26055);
nand U28403 (N_28403,N_26828,N_25886);
or U28404 (N_28404,N_26414,N_26855);
nand U28405 (N_28405,N_25620,N_26272);
and U28406 (N_28406,N_26381,N_25573);
or U28407 (N_28407,N_25625,N_25503);
or U28408 (N_28408,N_26842,N_26777);
and U28409 (N_28409,N_26515,N_26604);
nor U28410 (N_28410,N_26263,N_25977);
nor U28411 (N_28411,N_26806,N_26956);
nand U28412 (N_28412,N_26705,N_25972);
or U28413 (N_28413,N_26512,N_26620);
and U28414 (N_28414,N_25755,N_25769);
or U28415 (N_28415,N_25651,N_26010);
and U28416 (N_28416,N_26799,N_26790);
and U28417 (N_28417,N_25806,N_26841);
xnor U28418 (N_28418,N_25656,N_26284);
or U28419 (N_28419,N_26669,N_26410);
or U28420 (N_28420,N_26255,N_26098);
nand U28421 (N_28421,N_25847,N_25638);
or U28422 (N_28422,N_26972,N_26750);
nor U28423 (N_28423,N_25673,N_26839);
nor U28424 (N_28424,N_26560,N_26011);
xor U28425 (N_28425,N_25822,N_26078);
nor U28426 (N_28426,N_26977,N_26991);
nor U28427 (N_28427,N_25780,N_26811);
nor U28428 (N_28428,N_25927,N_26374);
xor U28429 (N_28429,N_26225,N_26089);
nand U28430 (N_28430,N_25827,N_26848);
nor U28431 (N_28431,N_26224,N_25754);
or U28432 (N_28432,N_25533,N_25735);
xnor U28433 (N_28433,N_26796,N_26838);
xnor U28434 (N_28434,N_25941,N_25814);
and U28435 (N_28435,N_26017,N_25576);
and U28436 (N_28436,N_26195,N_25947);
or U28437 (N_28437,N_25907,N_26829);
and U28438 (N_28438,N_26700,N_25765);
nand U28439 (N_28439,N_26770,N_26168);
and U28440 (N_28440,N_26940,N_26014);
or U28441 (N_28441,N_26383,N_26303);
and U28442 (N_28442,N_25609,N_26773);
nor U28443 (N_28443,N_26772,N_26407);
or U28444 (N_28444,N_26259,N_26112);
nand U28445 (N_28445,N_26426,N_25817);
or U28446 (N_28446,N_25789,N_26776);
xnor U28447 (N_28447,N_26001,N_26682);
xnor U28448 (N_28448,N_26855,N_25704);
or U28449 (N_28449,N_26954,N_25584);
nand U28450 (N_28450,N_26900,N_25925);
nor U28451 (N_28451,N_26671,N_26013);
and U28452 (N_28452,N_26131,N_26958);
xnor U28453 (N_28453,N_25912,N_26022);
or U28454 (N_28454,N_26456,N_26055);
nor U28455 (N_28455,N_25553,N_26327);
nand U28456 (N_28456,N_26858,N_25955);
and U28457 (N_28457,N_26088,N_26774);
nand U28458 (N_28458,N_26029,N_25648);
nor U28459 (N_28459,N_26939,N_26644);
nor U28460 (N_28460,N_25524,N_25753);
or U28461 (N_28461,N_25655,N_26781);
xnor U28462 (N_28462,N_25848,N_26070);
nand U28463 (N_28463,N_26622,N_26208);
and U28464 (N_28464,N_26579,N_26326);
nand U28465 (N_28465,N_26161,N_26219);
xor U28466 (N_28466,N_26390,N_26246);
nand U28467 (N_28467,N_26950,N_26700);
and U28468 (N_28468,N_26773,N_26862);
and U28469 (N_28469,N_25661,N_25643);
nor U28470 (N_28470,N_26042,N_25696);
nor U28471 (N_28471,N_26796,N_26575);
nor U28472 (N_28472,N_26734,N_25879);
nor U28473 (N_28473,N_26246,N_25898);
and U28474 (N_28474,N_26852,N_26374);
nand U28475 (N_28475,N_25652,N_26224);
and U28476 (N_28476,N_26418,N_26056);
nor U28477 (N_28477,N_26650,N_25704);
and U28478 (N_28478,N_26292,N_26736);
or U28479 (N_28479,N_25890,N_26318);
nand U28480 (N_28480,N_26320,N_25593);
or U28481 (N_28481,N_25597,N_26468);
xor U28482 (N_28482,N_26655,N_25998);
and U28483 (N_28483,N_26285,N_25813);
or U28484 (N_28484,N_26368,N_26611);
nand U28485 (N_28485,N_26640,N_26110);
nand U28486 (N_28486,N_26438,N_26958);
and U28487 (N_28487,N_26068,N_26201);
or U28488 (N_28488,N_26010,N_25623);
nand U28489 (N_28489,N_26068,N_26459);
and U28490 (N_28490,N_26349,N_25645);
xor U28491 (N_28491,N_26785,N_26252);
xnor U28492 (N_28492,N_26912,N_26084);
and U28493 (N_28493,N_26101,N_25973);
nor U28494 (N_28494,N_25928,N_25866);
nor U28495 (N_28495,N_25569,N_26000);
xor U28496 (N_28496,N_26534,N_26844);
nand U28497 (N_28497,N_25901,N_25714);
nor U28498 (N_28498,N_25974,N_25946);
nand U28499 (N_28499,N_25922,N_26435);
nor U28500 (N_28500,N_27132,N_28233);
xor U28501 (N_28501,N_27075,N_27598);
nand U28502 (N_28502,N_27767,N_27231);
nor U28503 (N_28503,N_27530,N_28326);
and U28504 (N_28504,N_28410,N_27082);
nor U28505 (N_28505,N_27574,N_28393);
or U28506 (N_28506,N_28034,N_27243);
xor U28507 (N_28507,N_28386,N_27868);
nand U28508 (N_28508,N_27623,N_27663);
and U28509 (N_28509,N_27269,N_28276);
nor U28510 (N_28510,N_27485,N_27312);
and U28511 (N_28511,N_27510,N_28292);
xnor U28512 (N_28512,N_27923,N_27008);
xnor U28513 (N_28513,N_28044,N_27771);
nand U28514 (N_28514,N_28452,N_27221);
xnor U28515 (N_28515,N_28318,N_27464);
nor U28516 (N_28516,N_27539,N_27276);
nor U28517 (N_28517,N_27810,N_27885);
and U28518 (N_28518,N_27319,N_27053);
xnor U28519 (N_28519,N_28475,N_27209);
and U28520 (N_28520,N_28270,N_28461);
nand U28521 (N_28521,N_28399,N_27861);
and U28522 (N_28522,N_27650,N_27831);
xor U28523 (N_28523,N_28086,N_27138);
xor U28524 (N_28524,N_28129,N_27415);
and U28525 (N_28525,N_28430,N_27707);
or U28526 (N_28526,N_28235,N_27286);
xnor U28527 (N_28527,N_27896,N_28496);
or U28528 (N_28528,N_28466,N_27747);
or U28529 (N_28529,N_28001,N_28269);
and U28530 (N_28530,N_27103,N_27427);
nor U28531 (N_28531,N_27121,N_28405);
nor U28532 (N_28532,N_28415,N_27124);
or U28533 (N_28533,N_27993,N_28121);
nand U28534 (N_28534,N_28319,N_28073);
xnor U28535 (N_28535,N_27755,N_28230);
or U28536 (N_28536,N_27324,N_27323);
nor U28537 (N_28537,N_28147,N_27791);
or U28538 (N_28538,N_27382,N_27271);
nor U28539 (N_28539,N_27632,N_28289);
or U28540 (N_28540,N_27070,N_27552);
and U28541 (N_28541,N_27912,N_27529);
xor U28542 (N_28542,N_27190,N_27919);
xor U28543 (N_28543,N_28153,N_27633);
nor U28544 (N_28544,N_27402,N_28371);
xor U28545 (N_28545,N_28241,N_28188);
or U28546 (N_28546,N_27524,N_28332);
nand U28547 (N_28547,N_28013,N_28493);
and U28548 (N_28548,N_28464,N_27975);
and U28549 (N_28549,N_27191,N_27836);
or U28550 (N_28550,N_27676,N_27715);
or U28551 (N_28551,N_27911,N_28412);
and U28552 (N_28552,N_28113,N_28271);
xnor U28553 (N_28553,N_27514,N_27216);
xnor U28554 (N_28554,N_27520,N_27815);
nand U28555 (N_28555,N_28028,N_27828);
and U28556 (N_28556,N_28005,N_28402);
xor U28557 (N_28557,N_28211,N_28221);
or U28558 (N_28558,N_27400,N_27389);
nand U28559 (N_28559,N_27294,N_28063);
or U28560 (N_28560,N_28354,N_27056);
and U28561 (N_28561,N_27973,N_27928);
xor U28562 (N_28562,N_28409,N_28240);
or U28563 (N_28563,N_27962,N_28075);
nor U28564 (N_28564,N_27852,N_27983);
and U28565 (N_28565,N_27732,N_27544);
xor U28566 (N_28566,N_27410,N_27097);
xnor U28567 (N_28567,N_27435,N_27335);
nand U28568 (N_28568,N_27417,N_27526);
or U28569 (N_28569,N_27274,N_27307);
xor U28570 (N_28570,N_27576,N_27541);
or U28571 (N_28571,N_27786,N_27395);
nand U28572 (N_28572,N_27292,N_27545);
nand U28573 (N_28573,N_27062,N_27260);
and U28574 (N_28574,N_27645,N_27575);
and U28575 (N_28575,N_28408,N_27193);
xor U28576 (N_28576,N_27423,N_27291);
nor U28577 (N_28577,N_28307,N_28268);
or U28578 (N_28578,N_28096,N_28195);
xnor U28579 (N_28579,N_28352,N_27431);
nor U28580 (N_28580,N_28131,N_27929);
nor U28581 (N_28581,N_27931,N_27807);
or U28582 (N_28582,N_27522,N_27957);
nand U28583 (N_28583,N_27573,N_27240);
nand U28584 (N_28584,N_27586,N_27613);
nand U28585 (N_28585,N_28051,N_27763);
and U28586 (N_28586,N_28469,N_27135);
and U28587 (N_28587,N_27250,N_28202);
xor U28588 (N_28588,N_28298,N_27501);
or U28589 (N_28589,N_27607,N_27184);
and U28590 (N_28590,N_28036,N_27015);
xnor U28591 (N_28591,N_28128,N_28181);
nor U28592 (N_28592,N_27453,N_27067);
and U28593 (N_28593,N_27314,N_28377);
xor U28594 (N_28594,N_27662,N_28481);
and U28595 (N_28595,N_27517,N_28209);
or U28596 (N_28596,N_28116,N_28480);
xnor U28597 (N_28597,N_27420,N_27803);
and U28598 (N_28598,N_28123,N_27069);
nand U28599 (N_28599,N_28262,N_27030);
xor U28600 (N_28600,N_27330,N_27599);
nand U28601 (N_28601,N_28168,N_27328);
or U28602 (N_28602,N_27867,N_28379);
xor U28603 (N_28603,N_27927,N_27716);
or U28604 (N_28604,N_27381,N_27512);
nand U28605 (N_28605,N_27338,N_28249);
or U28606 (N_28606,N_27034,N_27013);
nor U28607 (N_28607,N_27155,N_27845);
and U28608 (N_28608,N_28474,N_28068);
nand U28609 (N_28609,N_28117,N_27835);
nand U28610 (N_28610,N_28070,N_28085);
or U28611 (N_28611,N_28038,N_27438);
or U28612 (N_28612,N_28421,N_27612);
xor U28613 (N_28613,N_27806,N_28373);
xor U28614 (N_28614,N_27717,N_27698);
and U28615 (N_28615,N_27805,N_27089);
nor U28616 (N_28616,N_27133,N_27948);
nand U28617 (N_28617,N_27683,N_28312);
nand U28618 (N_28618,N_28056,N_27985);
and U28619 (N_28619,N_28033,N_27907);
and U28620 (N_28620,N_28148,N_27478);
and U28621 (N_28621,N_27699,N_27119);
and U28622 (N_28622,N_27198,N_27331);
or U28623 (N_28623,N_27793,N_27101);
xor U28624 (N_28624,N_28215,N_27939);
nor U28625 (N_28625,N_27293,N_27935);
or U28626 (N_28626,N_28093,N_27998);
nor U28627 (N_28627,N_27022,N_27201);
and U28628 (N_28628,N_27005,N_28160);
and U28629 (N_28629,N_27149,N_27516);
or U28630 (N_28630,N_27126,N_27403);
and U28631 (N_28631,N_27629,N_27457);
nor U28632 (N_28632,N_27981,N_28426);
nand U28633 (N_28633,N_27146,N_27021);
nor U28634 (N_28634,N_27970,N_27233);
xor U28635 (N_28635,N_27525,N_27822);
and U28636 (N_28636,N_27002,N_28010);
and U28637 (N_28637,N_27688,N_27383);
xnor U28638 (N_28638,N_28463,N_27606);
and U28639 (N_28639,N_27242,N_27665);
xor U28640 (N_28640,N_27009,N_27055);
nand U28641 (N_28641,N_28169,N_27932);
xnor U28642 (N_28642,N_27901,N_28105);
nor U28643 (N_28643,N_27262,N_27057);
nor U28644 (N_28644,N_27470,N_27642);
or U28645 (N_28645,N_27533,N_27549);
xor U28646 (N_28646,N_27279,N_27950);
xor U28647 (N_28647,N_27284,N_27441);
nor U28648 (N_28648,N_27466,N_27397);
or U28649 (N_28649,N_27780,N_27891);
nand U28650 (N_28650,N_27345,N_27820);
or U28651 (N_28651,N_28002,N_28444);
xnor U28652 (N_28652,N_28356,N_27158);
nand U28653 (N_28653,N_27167,N_27433);
nor U28654 (N_28654,N_27289,N_27694);
nor U28655 (N_28655,N_27313,N_27701);
nand U28656 (N_28656,N_28017,N_27593);
and U28657 (N_28657,N_27963,N_27727);
nor U28658 (N_28658,N_27961,N_27166);
or U28659 (N_28659,N_27120,N_27559);
nor U28660 (N_28660,N_28037,N_27589);
or U28661 (N_28661,N_27334,N_27494);
and U28662 (N_28662,N_27326,N_27143);
xnor U28663 (N_28663,N_27875,N_27239);
nor U28664 (N_28664,N_27758,N_28264);
and U28665 (N_28665,N_27404,N_27863);
xnor U28666 (N_28666,N_28341,N_28114);
nor U28667 (N_28667,N_27208,N_27624);
xor U28668 (N_28668,N_27904,N_27964);
nand U28669 (N_28669,N_27686,N_27257);
and U28670 (N_28670,N_27086,N_27267);
nand U28671 (N_28671,N_27064,N_28431);
and U28672 (N_28672,N_28258,N_27342);
or U28673 (N_28673,N_28171,N_27367);
xor U28674 (N_28674,N_27557,N_27532);
or U28675 (N_28675,N_27600,N_27995);
nor U28676 (N_28676,N_27712,N_27482);
xor U28677 (N_28677,N_27789,N_27808);
or U28678 (N_28678,N_27169,N_27817);
xor U28679 (N_28679,N_28369,N_27211);
nor U28680 (N_28680,N_27737,N_28316);
nor U28681 (N_28681,N_27503,N_27653);
and U28682 (N_28682,N_27361,N_27247);
and U28683 (N_28683,N_28484,N_27369);
nor U28684 (N_28684,N_27540,N_27459);
nand U28685 (N_28685,N_27677,N_28035);
or U28686 (N_28686,N_27892,N_27204);
nor U28687 (N_28687,N_28178,N_28237);
nor U28688 (N_28688,N_27638,N_27227);
and U28689 (N_28689,N_27496,N_27620);
or U28690 (N_28690,N_27074,N_27451);
nor U28691 (N_28691,N_28045,N_27012);
or U28692 (N_28692,N_27764,N_27223);
or U28693 (N_28693,N_27684,N_28203);
xnor U28694 (N_28694,N_28141,N_27579);
or U28695 (N_28695,N_27136,N_27432);
nor U28696 (N_28696,N_28004,N_27956);
or U28697 (N_28697,N_27477,N_28227);
and U28698 (N_28698,N_27192,N_27238);
and U28699 (N_28699,N_27736,N_28065);
nor U28700 (N_28700,N_28222,N_27938);
or U28701 (N_28701,N_27813,N_27194);
nand U28702 (N_28702,N_27263,N_27385);
and U28703 (N_28703,N_27253,N_27856);
nand U28704 (N_28704,N_28259,N_27029);
xnor U28705 (N_28705,N_27832,N_28254);
xor U28706 (N_28706,N_27475,N_27602);
xnor U28707 (N_28707,N_27615,N_27387);
or U28708 (N_28708,N_27375,N_27173);
xor U28709 (N_28709,N_27456,N_27798);
and U28710 (N_28710,N_28427,N_27418);
nand U28711 (N_28711,N_27337,N_27827);
xnor U28712 (N_28712,N_27654,N_28458);
xor U28713 (N_28713,N_28353,N_27960);
and U28714 (N_28714,N_27226,N_27171);
nor U28715 (N_28715,N_27316,N_27241);
xnor U28716 (N_28716,N_28455,N_27587);
or U28717 (N_28717,N_27864,N_28328);
and U28718 (N_28718,N_27799,N_27042);
or U28719 (N_28719,N_27430,N_28360);
or U28720 (N_28720,N_28363,N_28150);
nand U28721 (N_28721,N_28416,N_28253);
and U28722 (N_28722,N_27584,N_28300);
nor U28723 (N_28723,N_27842,N_27185);
nand U28724 (N_28724,N_28494,N_27333);
or U28725 (N_28725,N_28392,N_27290);
and U28726 (N_28726,N_27673,N_28087);
nand U28727 (N_28727,N_28330,N_27087);
or U28728 (N_28728,N_27353,N_27726);
xnor U28729 (N_28729,N_27505,N_28336);
nand U28730 (N_28730,N_27183,N_27486);
nand U28731 (N_28731,N_28216,N_27643);
nor U28732 (N_28732,N_27866,N_27405);
xor U28733 (N_28733,N_27644,N_27481);
nor U28734 (N_28734,N_28283,N_27657);
nand U28735 (N_28735,N_27844,N_27955);
or U28736 (N_28736,N_27007,N_27770);
or U28737 (N_28737,N_27422,N_28201);
nand U28738 (N_28738,N_28378,N_28314);
and U28739 (N_28739,N_27743,N_27161);
xnor U28740 (N_28740,N_28324,N_27660);
or U28741 (N_28741,N_27959,N_27838);
and U28742 (N_28742,N_27092,N_27601);
xnor U28743 (N_28743,N_27641,N_27611);
and U28744 (N_28744,N_27018,N_27968);
xnor U28745 (N_28745,N_28000,N_27869);
or U28746 (N_28746,N_27926,N_27272);
nor U28747 (N_28747,N_27814,N_27592);
xnor U28748 (N_28748,N_27152,N_27084);
nor U28749 (N_28749,N_27947,N_28208);
xor U28750 (N_28750,N_27548,N_27256);
and U28751 (N_28751,N_27218,N_27350);
nor U28752 (N_28752,N_27249,N_28471);
nand U28753 (N_28753,N_27298,N_27823);
nor U28754 (N_28754,N_27225,N_28048);
nor U28755 (N_28755,N_27873,N_27401);
or U28756 (N_28756,N_27098,N_27168);
and U28757 (N_28757,N_28125,N_28435);
xnor U28758 (N_28758,N_27199,N_28008);
nand U28759 (N_28759,N_28217,N_27693);
xor U28760 (N_28760,N_27027,N_28091);
or U28761 (N_28761,N_28295,N_27761);
and U28762 (N_28762,N_27941,N_28489);
xnor U28763 (N_28763,N_28055,N_27877);
and U28764 (N_28764,N_27329,N_27762);
nand U28765 (N_28765,N_27170,N_27031);
nand U28766 (N_28766,N_27449,N_27523);
xnor U28767 (N_28767,N_27380,N_27635);
nand U28768 (N_28768,N_27426,N_27550);
nor U28769 (N_28769,N_28453,N_27851);
nand U28770 (N_28770,N_28454,N_27910);
nand U28771 (N_28771,N_27346,N_27439);
xor U28772 (N_28772,N_28343,N_27492);
xnor U28773 (N_28773,N_27140,N_27206);
nor U28774 (N_28774,N_27854,N_27547);
xor U28775 (N_28775,N_27434,N_27407);
nand U28776 (N_28776,N_27718,N_27855);
and U28777 (N_28777,N_27145,N_27872);
xnor U28778 (N_28778,N_27376,N_28012);
xnor U28779 (N_28779,N_27108,N_27966);
or U28780 (N_28780,N_27936,N_27930);
and U28781 (N_28781,N_27871,N_28071);
or U28782 (N_28782,N_27977,N_28257);
xor U28783 (N_28783,N_28383,N_27571);
nand U28784 (N_28784,N_27413,N_27659);
nand U28785 (N_28785,N_27390,N_28438);
xor U28786 (N_28786,N_28149,N_27651);
xnor U28787 (N_28787,N_28401,N_27270);
nand U28788 (N_28788,N_27436,N_27819);
xor U28789 (N_28789,N_27618,N_28288);
and U28790 (N_28790,N_27965,N_28250);
nand U28791 (N_28791,N_27588,N_28029);
or U28792 (N_28792,N_28205,N_27740);
nor U28793 (N_28793,N_28337,N_27924);
nand U28794 (N_28794,N_28166,N_27577);
nand U28795 (N_28795,N_28122,N_28433);
and U28796 (N_28796,N_27640,N_27255);
xnor U28797 (N_28797,N_27462,N_28425);
or U28798 (N_28798,N_28245,N_28076);
nor U28799 (N_28799,N_27542,N_27165);
nor U28800 (N_28800,N_27306,N_28236);
nor U28801 (N_28801,N_27655,N_28311);
nand U28802 (N_28802,N_27339,N_27036);
xnor U28803 (N_28803,N_27077,N_27578);
xnor U28804 (N_28804,N_27646,N_28439);
and U28805 (N_28805,N_28339,N_27045);
nand U28806 (N_28806,N_28473,N_27969);
nor U28807 (N_28807,N_27038,N_28424);
nor U28808 (N_28808,N_28140,N_27858);
nand U28809 (N_28809,N_27213,N_28238);
or U28810 (N_28810,N_28303,N_27252);
and U28811 (N_28811,N_28476,N_27258);
and U28812 (N_28812,N_28462,N_28478);
nand U28813 (N_28813,N_28305,N_27795);
nand U28814 (N_28814,N_28152,N_27776);
xnor U28815 (N_28815,N_27078,N_28003);
and U28816 (N_28816,N_27399,N_27428);
xnor U28817 (N_28817,N_28403,N_28491);
nand U28818 (N_28818,N_27489,N_27849);
nor U28819 (N_28819,N_27090,N_28170);
xnor U28820 (N_28820,N_27754,N_28180);
and U28821 (N_28821,N_27172,N_27044);
or U28822 (N_28822,N_27102,N_28186);
xor U28823 (N_28823,N_27534,N_28077);
nand U28824 (N_28824,N_27862,N_27859);
nand U28825 (N_28825,N_27610,N_28313);
and U28826 (N_28826,N_27130,N_27105);
nor U28827 (N_28827,N_28165,N_27236);
or U28828 (N_28828,N_27359,N_28135);
nor U28829 (N_28829,N_27784,N_27502);
or U28830 (N_28830,N_28119,N_28362);
nor U28831 (N_28831,N_27181,N_28176);
or U28832 (N_28832,N_28483,N_27468);
and U28833 (N_28833,N_27551,N_27695);
and U28834 (N_28834,N_27412,N_27095);
xor U28835 (N_28835,N_28375,N_27893);
nor U28836 (N_28836,N_27750,N_27508);
or U28837 (N_28837,N_27971,N_28025);
nand U28838 (N_28838,N_28499,N_27809);
and U28839 (N_28839,N_27200,N_28239);
and U28840 (N_28840,N_27178,N_27702);
or U28841 (N_28841,N_28108,N_27365);
or U28842 (N_28842,N_28225,N_27648);
nor U28843 (N_28843,N_27488,N_27521);
or U28844 (N_28844,N_27019,N_27847);
and U28845 (N_28845,N_27691,N_27821);
or U28846 (N_28846,N_28118,N_28218);
and U28847 (N_28847,N_27134,N_27409);
xnor U28848 (N_28848,N_27982,N_27748);
xor U28849 (N_28849,N_28043,N_27281);
or U28850 (N_28850,N_27555,N_28023);
xor U28851 (N_28851,N_27017,N_28187);
or U28852 (N_28852,N_27709,N_28272);
xor U28853 (N_28853,N_28112,N_28376);
and U28854 (N_28854,N_28136,N_27467);
xnor U28855 (N_28855,N_27921,N_28364);
nand U28856 (N_28856,N_27116,N_28109);
or U28857 (N_28857,N_27972,N_28232);
nor U28858 (N_28858,N_28206,N_28185);
or U28859 (N_28859,N_27379,N_27558);
or U28860 (N_28860,N_28107,N_27952);
nand U28861 (N_28861,N_28223,N_28139);
xnor U28862 (N_28862,N_28275,N_27065);
or U28863 (N_28863,N_27091,N_27857);
and U28864 (N_28864,N_28164,N_27890);
nand U28865 (N_28865,N_27127,N_27583);
xor U28866 (N_28866,N_27215,N_27051);
or U28867 (N_28867,N_27829,N_28340);
nand U28868 (N_28868,N_27352,N_27107);
and U28869 (N_28869,N_27280,N_27419);
or U28870 (N_28870,N_28212,N_27561);
nand U28871 (N_28871,N_27656,N_27690);
and U28872 (N_28872,N_28361,N_27093);
or U28873 (N_28873,N_27604,N_27878);
and U28874 (N_28874,N_27913,N_28022);
and U28875 (N_28875,N_27569,N_27949);
or U28876 (N_28876,N_27408,N_28226);
and U28877 (N_28877,N_27917,N_27028);
nand U28878 (N_28878,N_27499,N_28006);
nand U28879 (N_28879,N_27565,N_27368);
or U28880 (N_28880,N_27076,N_28050);
nand U28881 (N_28881,N_27850,N_28310);
nand U28882 (N_28882,N_28159,N_28460);
xnor U28883 (N_28883,N_27630,N_27264);
xnor U28884 (N_28884,N_27287,N_28320);
and U28885 (N_28885,N_27111,N_27830);
nor U28886 (N_28886,N_27765,N_27528);
or U28887 (N_28887,N_27392,N_27465);
nand U28888 (N_28888,N_27493,N_28059);
and U28889 (N_28889,N_27224,N_27682);
and U28890 (N_28890,N_27870,N_27942);
and U28891 (N_28891,N_27685,N_27112);
xnor U28892 (N_28892,N_27636,N_28154);
xor U28893 (N_28893,N_27853,N_27637);
or U28894 (N_28894,N_28115,N_28143);
and U28895 (N_28895,N_28231,N_27538);
and U28896 (N_28896,N_27908,N_27816);
nor U28897 (N_28897,N_27440,N_27273);
nand U28898 (N_28898,N_27667,N_27824);
nand U28899 (N_28899,N_27980,N_28284);
xnor U28900 (N_28900,N_27788,N_28089);
xnor U28901 (N_28901,N_27720,N_27511);
or U28902 (N_28902,N_27536,N_27356);
nand U28903 (N_28903,N_27234,N_28391);
nand U28904 (N_28904,N_27518,N_27837);
xnor U28905 (N_28905,N_27778,N_27495);
or U28906 (N_28906,N_27487,N_28083);
or U28907 (N_28907,N_28306,N_28014);
xor U28908 (N_28908,N_28368,N_27230);
nand U28909 (N_28909,N_28447,N_27474);
nand U28910 (N_28910,N_28039,N_27443);
or U28911 (N_28911,N_28220,N_28101);
nor U28912 (N_28912,N_28331,N_27394);
and U28913 (N_28913,N_27189,N_28219);
nor U28914 (N_28914,N_28321,N_28302);
xor U28915 (N_28915,N_27745,N_27933);
nand U28916 (N_28916,N_27631,N_27976);
and U28917 (N_28917,N_27661,N_27760);
and U28918 (N_28918,N_27148,N_27840);
nand U28919 (N_28919,N_27905,N_27621);
and U28920 (N_28920,N_28229,N_27724);
nand U28921 (N_28921,N_27043,N_27498);
nand U28922 (N_28922,N_27781,N_27251);
nand U28923 (N_28923,N_27527,N_27647);
or U28924 (N_28924,N_27777,N_27915);
and U28925 (N_28925,N_27902,N_28103);
nor U28926 (N_28926,N_27164,N_28459);
nand U28927 (N_28927,N_27050,N_28026);
and U28928 (N_28928,N_27446,N_27071);
nand U28929 (N_28929,N_28440,N_27425);
nand U28930 (N_28930,N_27773,N_27100);
or U28931 (N_28931,N_27129,N_28327);
and U28932 (N_28932,N_27713,N_28088);
and U28933 (N_28933,N_27792,N_28266);
xnor U28934 (N_28934,N_27160,N_27708);
nand U28935 (N_28935,N_28106,N_27480);
nand U28936 (N_28936,N_28120,N_28432);
nor U28937 (N_28937,N_28009,N_27244);
nand U28938 (N_28938,N_28296,N_27914);
nor U28939 (N_28939,N_27305,N_28423);
or U28940 (N_28940,N_27336,N_28351);
or U28941 (N_28941,N_28054,N_28064);
and U28942 (N_28942,N_28132,N_28381);
and U28943 (N_28943,N_27176,N_27219);
nand U28944 (N_28944,N_28420,N_27603);
or U28945 (N_28945,N_28246,N_27311);
or U28946 (N_28946,N_28315,N_27010);
nor U28947 (N_28947,N_27590,N_27634);
or U28948 (N_28948,N_27207,N_27396);
or U28949 (N_28949,N_27714,N_27944);
xor U28950 (N_28950,N_27174,N_28485);
and U28951 (N_28951,N_28357,N_27594);
nor U28952 (N_28952,N_28082,N_27014);
nand U28953 (N_28953,N_27039,N_28058);
nand U28954 (N_28954,N_27888,N_28344);
xnor U28955 (N_28955,N_28414,N_27741);
xnor U28956 (N_28956,N_27188,N_27566);
and U28957 (N_28957,N_27066,N_27288);
and U28958 (N_28958,N_28488,N_27609);
nand U28959 (N_28959,N_27114,N_28052);
nor U28960 (N_28960,N_28286,N_27490);
nor U28961 (N_28961,N_27406,N_28278);
and U28962 (N_28962,N_27729,N_27327);
and U28963 (N_28963,N_27779,N_27063);
and U28964 (N_28964,N_27001,N_28124);
or U28965 (N_28965,N_27026,N_27903);
or U28966 (N_28966,N_27774,N_27687);
xor U28967 (N_28967,N_27783,N_27749);
nor U28968 (N_28968,N_28495,N_27974);
and U28969 (N_28969,N_28347,N_27384);
and U28970 (N_28970,N_28279,N_28338);
and U28971 (N_28971,N_27568,N_27833);
or U28972 (N_28972,N_27483,N_27627);
xor U28973 (N_28973,N_28090,N_28290);
and U28974 (N_28974,N_27372,N_28387);
nand U28975 (N_28975,N_27343,N_27790);
xor U28976 (N_28976,N_27000,N_28384);
xor U28977 (N_28977,N_28449,N_27308);
nor U28978 (N_28978,N_27060,N_27731);
xnor U28979 (N_28979,N_28281,N_28406);
and U28980 (N_28980,N_27801,N_28365);
xor U28981 (N_28981,N_28104,N_27535);
xnor U28982 (N_28982,N_28027,N_27989);
nand U28983 (N_28983,N_28134,N_27374);
or U28984 (N_28984,N_27506,N_28057);
and U28985 (N_28985,N_28099,N_27591);
and U28986 (N_28986,N_28299,N_28042);
and U28987 (N_28987,N_27616,N_28062);
nand U28988 (N_28988,N_27797,N_27068);
and U28989 (N_28989,N_27259,N_28097);
nor U28990 (N_28990,N_27572,N_28446);
nor U28991 (N_28991,N_28251,N_27706);
nor U28992 (N_28992,N_27117,N_27710);
or U28993 (N_28993,N_27567,N_27297);
nor U28994 (N_28994,N_27079,N_28252);
or U28995 (N_28995,N_27006,N_27237);
nor U28996 (N_28996,N_27414,N_28385);
nand U28997 (N_28997,N_27934,N_28265);
nand U28998 (N_28998,N_27622,N_27059);
nand U28999 (N_28999,N_27388,N_27865);
xnor U29000 (N_29000,N_27049,N_28400);
nand U29001 (N_29001,N_27652,N_28078);
nor U29002 (N_29002,N_27442,N_28244);
nor U29003 (N_29003,N_28182,N_28192);
nor U29004 (N_29004,N_27922,N_27639);
xor U29005 (N_29005,N_27154,N_27347);
and U29006 (N_29006,N_27879,N_27246);
nand U29007 (N_29007,N_28172,N_27671);
nor U29008 (N_29008,N_28418,N_28293);
nand U29009 (N_29009,N_27826,N_27794);
nor U29010 (N_29010,N_27672,N_28015);
nand U29011 (N_29011,N_27800,N_28323);
xnor U29012 (N_29012,N_27378,N_28177);
xor U29013 (N_29013,N_28100,N_27450);
xor U29014 (N_29014,N_27841,N_28157);
nor U29015 (N_29015,N_27448,N_27469);
and U29016 (N_29016,N_28467,N_27220);
or U29017 (N_29017,N_28443,N_28079);
or U29018 (N_29018,N_27563,N_27564);
or U29019 (N_29019,N_28228,N_27898);
nor U29020 (N_29020,N_27197,N_28450);
nand U29021 (N_29021,N_28191,N_27811);
and U29022 (N_29022,N_28308,N_28407);
or U29023 (N_29023,N_28273,N_27366);
nor U29024 (N_29024,N_28031,N_28448);
xnor U29025 (N_29025,N_28094,N_27580);
nand U29026 (N_29026,N_27984,N_27674);
nand U29027 (N_29027,N_28456,N_27649);
nor U29028 (N_29028,N_28477,N_27889);
xnor U29029 (N_29029,N_27048,N_27282);
and U29030 (N_29030,N_27785,N_27759);
and U29031 (N_29031,N_28146,N_27245);
and U29032 (N_29032,N_27109,N_28282);
nand U29033 (N_29033,N_27473,N_28144);
xor U29034 (N_29034,N_28248,N_27562);
nand U29035 (N_29035,N_27883,N_27757);
nand U29036 (N_29036,N_27072,N_28374);
xor U29037 (N_29037,N_28173,N_27115);
nor U29038 (N_29038,N_28189,N_28417);
and U29039 (N_29039,N_27680,N_27137);
nor U29040 (N_29040,N_27011,N_27210);
nor U29041 (N_29041,N_28081,N_28445);
nand U29042 (N_29042,N_27177,N_28479);
xor U29043 (N_29043,N_28145,N_28267);
nor U29044 (N_29044,N_28335,N_27354);
and U29045 (N_29045,N_27187,N_27131);
nor U29046 (N_29046,N_28179,N_27118);
or U29047 (N_29047,N_27222,N_27304);
or U29048 (N_29048,N_27424,N_27991);
and U29049 (N_29049,N_27196,N_28021);
nand U29050 (N_29050,N_27476,N_27585);
nand U29051 (N_29051,N_28397,N_28472);
nor U29052 (N_29052,N_27205,N_28138);
nor U29053 (N_29053,N_28429,N_27159);
or U29054 (N_29054,N_28317,N_28053);
xor U29055 (N_29055,N_28102,N_28199);
and U29056 (N_29056,N_27628,N_27248);
and U29057 (N_29057,N_28277,N_28370);
or U29058 (N_29058,N_28007,N_27004);
nor U29059 (N_29059,N_27543,N_27775);
or U29060 (N_29060,N_28047,N_27461);
and U29061 (N_29061,N_27228,N_27739);
and U29062 (N_29062,N_27491,N_27229);
or U29063 (N_29063,N_28256,N_28127);
nand U29064 (N_29064,N_27625,N_27605);
nand U29065 (N_29065,N_27519,N_27348);
nor U29066 (N_29066,N_27768,N_28074);
nand U29067 (N_29067,N_27681,N_28492);
or U29068 (N_29068,N_27320,N_27212);
and U29069 (N_29069,N_27554,N_27033);
and U29070 (N_29070,N_28126,N_27581);
xor U29071 (N_29071,N_27825,N_27735);
and U29072 (N_29072,N_28247,N_28260);
or U29073 (N_29073,N_27391,N_27678);
and U29074 (N_29074,N_27742,N_27035);
or U29075 (N_29075,N_27283,N_27099);
and U29076 (N_29076,N_27300,N_27846);
nand U29077 (N_29077,N_27513,N_28255);
xnor U29078 (N_29078,N_28175,N_28190);
nor U29079 (N_29079,N_28436,N_28200);
xor U29080 (N_29080,N_28049,N_28297);
nand U29081 (N_29081,N_27988,N_27711);
nand U29082 (N_29082,N_28301,N_28437);
nor U29083 (N_29083,N_27696,N_27373);
or U29084 (N_29084,N_27411,N_27679);
and U29085 (N_29085,N_28390,N_27357);
xnor U29086 (N_29086,N_28018,N_27992);
xnor U29087 (N_29087,N_27725,N_28294);
nand U29088 (N_29088,N_27182,N_27332);
or U29089 (N_29089,N_28198,N_27179);
or U29090 (N_29090,N_27703,N_27344);
xnor U29091 (N_29091,N_28183,N_27582);
nor U29092 (N_29092,N_28263,N_28046);
or U29093 (N_29093,N_27860,N_27309);
xor U29094 (N_29094,N_28358,N_28024);
or U29095 (N_29095,N_28213,N_27722);
and U29096 (N_29096,N_27455,N_27953);
and U29097 (N_29097,N_27358,N_27734);
nor U29098 (N_29098,N_27900,N_27445);
nand U29099 (N_29099,N_27032,N_28309);
or U29100 (N_29100,N_28156,N_27839);
or U29101 (N_29101,N_27556,N_27484);
nor U29102 (N_29102,N_27986,N_28355);
xor U29103 (N_29103,N_28348,N_27416);
or U29104 (N_29104,N_27531,N_27322);
nor U29105 (N_29105,N_28304,N_28349);
nor U29106 (N_29106,N_28411,N_28224);
nand U29107 (N_29107,N_28490,N_27744);
or U29108 (N_29108,N_27507,N_28291);
and U29109 (N_29109,N_27472,N_27364);
xor U29110 (N_29110,N_27876,N_28468);
nor U29111 (N_29111,N_27509,N_27106);
or U29112 (N_29112,N_27738,N_28396);
nor U29113 (N_29113,N_27088,N_27772);
nor U29114 (N_29114,N_28133,N_27360);
and U29115 (N_29115,N_27125,N_28367);
or U29116 (N_29116,N_28388,N_27925);
and U29117 (N_29117,N_27546,N_28080);
nand U29118 (N_29118,N_27997,N_28174);
nor U29119 (N_29119,N_28151,N_27692);
xnor U29120 (N_29120,N_27139,N_28382);
and U29121 (N_29121,N_27214,N_27421);
and U29122 (N_29122,N_28016,N_27769);
or U29123 (N_29123,N_27967,N_27265);
nand U29124 (N_29124,N_27664,N_27954);
nor U29125 (N_29125,N_27945,N_27882);
and U29126 (N_29126,N_28366,N_28389);
or U29127 (N_29127,N_27398,N_27818);
nor U29128 (N_29128,N_27370,N_27894);
and U29129 (N_29129,N_28451,N_28197);
nand U29130 (N_29130,N_27751,N_27321);
nand U29131 (N_29131,N_27728,N_27147);
nand U29132 (N_29132,N_27073,N_27595);
nand U29133 (N_29133,N_27151,N_27317);
and U29134 (N_29134,N_27393,N_28486);
nor U29135 (N_29135,N_28342,N_27377);
and U29136 (N_29136,N_28441,N_28497);
and U29137 (N_29137,N_27315,N_27515);
nor U29138 (N_29138,N_27340,N_27150);
xnor U29139 (N_29139,N_27083,N_28040);
xor U29140 (N_29140,N_27041,N_27040);
or U29141 (N_29141,N_28465,N_27874);
xor U29142 (N_29142,N_27025,N_27597);
xnor U29143 (N_29143,N_28457,N_27937);
nand U29144 (N_29144,N_27386,N_27016);
xor U29145 (N_29145,N_28072,N_28142);
nor U29146 (N_29146,N_27046,N_27429);
nor U29147 (N_29147,N_27619,N_28110);
nand U29148 (N_29148,N_27162,N_28428);
nor U29149 (N_29149,N_27899,N_27085);
and U29150 (N_29150,N_28020,N_27463);
nand U29151 (N_29151,N_28395,N_27113);
nand U29152 (N_29152,N_28011,N_27142);
nor U29153 (N_29153,N_27979,N_28158);
or U29154 (N_29154,N_27918,N_27999);
nand U29155 (N_29155,N_27617,N_27733);
xor U29156 (N_29156,N_27054,N_27700);
or U29157 (N_29157,N_27277,N_28130);
and U29158 (N_29158,N_27987,N_28204);
nand U29159 (N_29159,N_28214,N_28243);
nand U29160 (N_29160,N_28193,N_27895);
or U29161 (N_29161,N_27299,N_28394);
nor U29162 (N_29162,N_28207,N_27202);
nor U29163 (N_29163,N_27812,N_27887);
nor U29164 (N_29164,N_27203,N_27024);
nand U29165 (N_29165,N_27596,N_27668);
nor U29166 (N_29166,N_27752,N_27195);
or U29167 (N_29167,N_27553,N_27047);
nor U29168 (N_29168,N_27094,N_27163);
nor U29169 (N_29169,N_27666,N_27537);
xor U29170 (N_29170,N_28155,N_28334);
or U29171 (N_29171,N_28019,N_28322);
and U29172 (N_29172,N_28069,N_28242);
xnor U29173 (N_29173,N_27848,N_28030);
or U29174 (N_29174,N_28032,N_28163);
xor U29175 (N_29175,N_27834,N_27504);
nand U29176 (N_29176,N_27080,N_27217);
nand U29177 (N_29177,N_27303,N_27122);
nor U29178 (N_29178,N_27940,N_27285);
or U29179 (N_29179,N_27437,N_28350);
and U29180 (N_29180,N_27301,N_27278);
nand U29181 (N_29181,N_27884,N_27447);
and U29182 (N_29182,N_27958,N_28482);
and U29183 (N_29183,N_27052,N_27254);
or U29184 (N_29184,N_27881,N_27802);
nor U29185 (N_29185,N_27906,N_28060);
xnor U29186 (N_29186,N_27951,N_27766);
nor U29187 (N_29187,N_28194,N_27782);
nor U29188 (N_29188,N_27110,N_28346);
or U29189 (N_29189,N_27705,N_27669);
nand U29190 (N_29190,N_27880,N_27670);
nand U29191 (N_29191,N_27123,N_28442);
and U29192 (N_29192,N_28359,N_28196);
and U29193 (N_29193,N_27753,N_27061);
nand U29194 (N_29194,N_28329,N_27626);
or U29195 (N_29195,N_27454,N_27295);
or U29196 (N_29196,N_28167,N_28422);
xnor U29197 (N_29197,N_27341,N_28210);
or U29198 (N_29198,N_27471,N_28470);
nand U29199 (N_29199,N_28487,N_27500);
and U29200 (N_29200,N_28285,N_27362);
and U29201 (N_29201,N_28184,N_28372);
and U29202 (N_29202,N_27232,N_27349);
nor U29203 (N_29203,N_28261,N_28067);
or U29204 (N_29204,N_27897,N_27796);
xnor U29205 (N_29205,N_28413,N_27275);
nand U29206 (N_29206,N_28419,N_27175);
nor U29207 (N_29207,N_27153,N_27675);
or U29208 (N_29208,N_27943,N_27721);
nand U29209 (N_29209,N_27371,N_28398);
or U29210 (N_29210,N_27658,N_27023);
nor U29211 (N_29211,N_27302,N_27037);
and U29212 (N_29212,N_28333,N_28325);
and U29213 (N_29213,N_27996,N_27746);
nand U29214 (N_29214,N_27909,N_27235);
xnor U29215 (N_29215,N_28111,N_27268);
and U29216 (N_29216,N_28061,N_27261);
xnor U29217 (N_29217,N_27128,N_27058);
xnor U29218 (N_29218,N_27104,N_28498);
nand U29219 (N_29219,N_27296,N_27723);
xnor U29220 (N_29220,N_27689,N_27730);
and U29221 (N_29221,N_27614,N_28084);
xor U29222 (N_29222,N_27978,N_27020);
xor U29223 (N_29223,N_28098,N_27156);
xor U29224 (N_29224,N_27608,N_27920);
and U29225 (N_29225,N_27946,N_28434);
xnor U29226 (N_29226,N_27570,N_27916);
or U29227 (N_29227,N_27697,N_27186);
nor U29228 (N_29228,N_27351,N_28280);
or U29229 (N_29229,N_27458,N_28287);
and U29230 (N_29230,N_27325,N_27560);
xnor U29231 (N_29231,N_27310,N_27719);
and U29232 (N_29232,N_28162,N_28095);
nor U29233 (N_29233,N_27452,N_27157);
xnor U29234 (N_29234,N_27704,N_27096);
nor U29235 (N_29235,N_27990,N_28137);
nor U29236 (N_29236,N_27994,N_28161);
and U29237 (N_29237,N_27318,N_27804);
xor U29238 (N_29238,N_27479,N_27756);
nand U29239 (N_29239,N_28345,N_28092);
nor U29240 (N_29240,N_27363,N_27355);
or U29241 (N_29241,N_28066,N_28404);
and U29242 (N_29242,N_27144,N_27886);
and U29243 (N_29243,N_27497,N_28274);
nand U29244 (N_29244,N_27266,N_27843);
and U29245 (N_29245,N_27003,N_27081);
xnor U29246 (N_29246,N_28041,N_28234);
nand U29247 (N_29247,N_27141,N_28380);
nand U29248 (N_29248,N_27787,N_27460);
nor U29249 (N_29249,N_27444,N_27180);
nand U29250 (N_29250,N_28391,N_27266);
and U29251 (N_29251,N_27790,N_27322);
nor U29252 (N_29252,N_27113,N_27561);
nand U29253 (N_29253,N_27986,N_27608);
nor U29254 (N_29254,N_27528,N_27654);
or U29255 (N_29255,N_27766,N_27271);
nand U29256 (N_29256,N_27485,N_27558);
nand U29257 (N_29257,N_27973,N_27744);
nor U29258 (N_29258,N_27295,N_27122);
or U29259 (N_29259,N_28197,N_27255);
nand U29260 (N_29260,N_27928,N_27034);
and U29261 (N_29261,N_28260,N_27347);
nor U29262 (N_29262,N_28286,N_27624);
and U29263 (N_29263,N_27739,N_27658);
or U29264 (N_29264,N_27522,N_27139);
and U29265 (N_29265,N_28295,N_27795);
or U29266 (N_29266,N_27318,N_28404);
nand U29267 (N_29267,N_27049,N_28072);
nor U29268 (N_29268,N_27811,N_27407);
nor U29269 (N_29269,N_28446,N_27243);
nor U29270 (N_29270,N_28226,N_27136);
and U29271 (N_29271,N_28052,N_27492);
nor U29272 (N_29272,N_27623,N_27096);
xnor U29273 (N_29273,N_28393,N_28122);
nand U29274 (N_29274,N_27563,N_27067);
or U29275 (N_29275,N_27699,N_27503);
or U29276 (N_29276,N_28241,N_28216);
or U29277 (N_29277,N_28414,N_28251);
and U29278 (N_29278,N_28173,N_27625);
nor U29279 (N_29279,N_28386,N_28473);
nand U29280 (N_29280,N_27325,N_28248);
nand U29281 (N_29281,N_27495,N_28048);
or U29282 (N_29282,N_28018,N_27944);
nor U29283 (N_29283,N_27297,N_28496);
nand U29284 (N_29284,N_27292,N_28475);
xor U29285 (N_29285,N_27595,N_27894);
and U29286 (N_29286,N_28471,N_28371);
or U29287 (N_29287,N_27810,N_27414);
nor U29288 (N_29288,N_28082,N_28494);
xnor U29289 (N_29289,N_28499,N_28394);
xor U29290 (N_29290,N_27962,N_27552);
or U29291 (N_29291,N_28136,N_27019);
or U29292 (N_29292,N_27747,N_27594);
or U29293 (N_29293,N_27826,N_27267);
and U29294 (N_29294,N_27896,N_28115);
nand U29295 (N_29295,N_27440,N_28137);
xor U29296 (N_29296,N_28388,N_27617);
or U29297 (N_29297,N_28479,N_27689);
and U29298 (N_29298,N_28308,N_27709);
and U29299 (N_29299,N_28119,N_27812);
xor U29300 (N_29300,N_28375,N_27006);
nor U29301 (N_29301,N_27339,N_28453);
or U29302 (N_29302,N_28009,N_27044);
xnor U29303 (N_29303,N_28082,N_27096);
nand U29304 (N_29304,N_28401,N_27275);
and U29305 (N_29305,N_27821,N_27082);
and U29306 (N_29306,N_27016,N_27772);
and U29307 (N_29307,N_27591,N_28004);
nor U29308 (N_29308,N_27477,N_27899);
xor U29309 (N_29309,N_28347,N_28054);
xnor U29310 (N_29310,N_27510,N_27440);
and U29311 (N_29311,N_28134,N_28102);
or U29312 (N_29312,N_27368,N_27521);
or U29313 (N_29313,N_27140,N_28222);
nor U29314 (N_29314,N_27984,N_27639);
and U29315 (N_29315,N_27588,N_27927);
and U29316 (N_29316,N_27217,N_27303);
xor U29317 (N_29317,N_27680,N_27812);
xor U29318 (N_29318,N_27237,N_28345);
nor U29319 (N_29319,N_27523,N_28310);
or U29320 (N_29320,N_27245,N_28211);
or U29321 (N_29321,N_28449,N_28014);
nor U29322 (N_29322,N_28245,N_28455);
nor U29323 (N_29323,N_28206,N_27202);
and U29324 (N_29324,N_28326,N_27459);
and U29325 (N_29325,N_27256,N_27434);
and U29326 (N_29326,N_27648,N_27109);
nor U29327 (N_29327,N_28006,N_28240);
xor U29328 (N_29328,N_27582,N_27912);
xor U29329 (N_29329,N_28099,N_28266);
nor U29330 (N_29330,N_27326,N_28309);
and U29331 (N_29331,N_27185,N_27959);
nor U29332 (N_29332,N_28205,N_27801);
nor U29333 (N_29333,N_27088,N_27918);
nand U29334 (N_29334,N_27642,N_28097);
xor U29335 (N_29335,N_28158,N_28428);
or U29336 (N_29336,N_27257,N_27839);
or U29337 (N_29337,N_27897,N_27056);
xnor U29338 (N_29338,N_27429,N_27251);
or U29339 (N_29339,N_27604,N_27356);
or U29340 (N_29340,N_27575,N_28134);
nor U29341 (N_29341,N_27232,N_28381);
and U29342 (N_29342,N_27012,N_27352);
nand U29343 (N_29343,N_27402,N_27401);
nor U29344 (N_29344,N_27166,N_27904);
nor U29345 (N_29345,N_27692,N_27634);
nor U29346 (N_29346,N_28460,N_27923);
nand U29347 (N_29347,N_27229,N_27818);
and U29348 (N_29348,N_27682,N_27272);
nor U29349 (N_29349,N_27617,N_27378);
nand U29350 (N_29350,N_28084,N_27723);
or U29351 (N_29351,N_28475,N_28255);
nand U29352 (N_29352,N_28131,N_27085);
nor U29353 (N_29353,N_27153,N_28304);
or U29354 (N_29354,N_27641,N_27823);
or U29355 (N_29355,N_27115,N_27027);
and U29356 (N_29356,N_28458,N_27719);
or U29357 (N_29357,N_27100,N_27086);
or U29358 (N_29358,N_28393,N_27754);
or U29359 (N_29359,N_28382,N_28400);
nor U29360 (N_29360,N_27504,N_28159);
and U29361 (N_29361,N_27265,N_27026);
nand U29362 (N_29362,N_28191,N_27243);
nand U29363 (N_29363,N_27685,N_28367);
nand U29364 (N_29364,N_27917,N_27764);
nand U29365 (N_29365,N_28409,N_27875);
or U29366 (N_29366,N_27719,N_28365);
or U29367 (N_29367,N_28363,N_27529);
xnor U29368 (N_29368,N_27053,N_27125);
nand U29369 (N_29369,N_28298,N_27877);
xnor U29370 (N_29370,N_27271,N_27917);
nor U29371 (N_29371,N_27513,N_28486);
and U29372 (N_29372,N_27289,N_28423);
nor U29373 (N_29373,N_28227,N_28438);
nor U29374 (N_29374,N_27685,N_27369);
xor U29375 (N_29375,N_27219,N_28231);
and U29376 (N_29376,N_27744,N_27505);
and U29377 (N_29377,N_27390,N_28372);
and U29378 (N_29378,N_27315,N_28330);
xnor U29379 (N_29379,N_28071,N_28404);
or U29380 (N_29380,N_27528,N_27894);
or U29381 (N_29381,N_28366,N_27952);
and U29382 (N_29382,N_27964,N_27657);
nand U29383 (N_29383,N_27363,N_28387);
or U29384 (N_29384,N_27990,N_27303);
or U29385 (N_29385,N_27222,N_27625);
or U29386 (N_29386,N_27180,N_28025);
and U29387 (N_29387,N_27159,N_27586);
or U29388 (N_29388,N_27641,N_28119);
and U29389 (N_29389,N_27566,N_27848);
nor U29390 (N_29390,N_28468,N_28341);
or U29391 (N_29391,N_27815,N_27934);
nand U29392 (N_29392,N_27854,N_28168);
and U29393 (N_29393,N_28074,N_27674);
xnor U29394 (N_29394,N_28342,N_28209);
nand U29395 (N_29395,N_27421,N_27877);
nand U29396 (N_29396,N_28422,N_27796);
nor U29397 (N_29397,N_28319,N_27093);
xnor U29398 (N_29398,N_27722,N_27303);
and U29399 (N_29399,N_27331,N_27867);
xor U29400 (N_29400,N_28302,N_27865);
xnor U29401 (N_29401,N_27449,N_27395);
nand U29402 (N_29402,N_27942,N_28241);
nor U29403 (N_29403,N_27933,N_27873);
nor U29404 (N_29404,N_28214,N_27633);
xor U29405 (N_29405,N_28148,N_27554);
or U29406 (N_29406,N_27538,N_27631);
xnor U29407 (N_29407,N_27576,N_28365);
nand U29408 (N_29408,N_27888,N_27010);
or U29409 (N_29409,N_27574,N_27476);
nor U29410 (N_29410,N_27136,N_27903);
nand U29411 (N_29411,N_27446,N_27024);
xor U29412 (N_29412,N_27759,N_27863);
or U29413 (N_29413,N_27938,N_28018);
or U29414 (N_29414,N_27597,N_27203);
and U29415 (N_29415,N_27922,N_27710);
xnor U29416 (N_29416,N_27298,N_28307);
nand U29417 (N_29417,N_27806,N_28252);
nand U29418 (N_29418,N_27965,N_27249);
nand U29419 (N_29419,N_27970,N_27307);
xnor U29420 (N_29420,N_27797,N_28341);
and U29421 (N_29421,N_28130,N_27948);
nand U29422 (N_29422,N_27200,N_27203);
or U29423 (N_29423,N_27192,N_27054);
and U29424 (N_29424,N_28316,N_28341);
or U29425 (N_29425,N_28228,N_27581);
or U29426 (N_29426,N_27119,N_27628);
xnor U29427 (N_29427,N_28269,N_27011);
and U29428 (N_29428,N_27344,N_27534);
or U29429 (N_29429,N_28372,N_27443);
xnor U29430 (N_29430,N_27068,N_27589);
and U29431 (N_29431,N_28047,N_28193);
nor U29432 (N_29432,N_27422,N_27545);
and U29433 (N_29433,N_28250,N_27895);
or U29434 (N_29434,N_27381,N_28231);
xor U29435 (N_29435,N_28195,N_28315);
and U29436 (N_29436,N_28220,N_27813);
and U29437 (N_29437,N_27955,N_27923);
nor U29438 (N_29438,N_27927,N_28238);
nand U29439 (N_29439,N_27591,N_27378);
nand U29440 (N_29440,N_27715,N_28402);
and U29441 (N_29441,N_28207,N_27840);
nand U29442 (N_29442,N_28280,N_27442);
or U29443 (N_29443,N_28452,N_27907);
nor U29444 (N_29444,N_28064,N_28148);
nor U29445 (N_29445,N_28283,N_28065);
or U29446 (N_29446,N_28352,N_27540);
nand U29447 (N_29447,N_28334,N_27275);
nor U29448 (N_29448,N_27765,N_27939);
nor U29449 (N_29449,N_27208,N_27642);
nand U29450 (N_29450,N_27324,N_27327);
xor U29451 (N_29451,N_28281,N_27685);
or U29452 (N_29452,N_27574,N_27970);
nor U29453 (N_29453,N_28052,N_27686);
nor U29454 (N_29454,N_28373,N_27388);
nor U29455 (N_29455,N_27734,N_27949);
or U29456 (N_29456,N_27965,N_27138);
nor U29457 (N_29457,N_27770,N_27017);
nor U29458 (N_29458,N_27326,N_27917);
nand U29459 (N_29459,N_27649,N_28289);
nand U29460 (N_29460,N_28335,N_28318);
nand U29461 (N_29461,N_28359,N_27895);
and U29462 (N_29462,N_27140,N_27543);
xor U29463 (N_29463,N_28113,N_27275);
or U29464 (N_29464,N_28270,N_27455);
or U29465 (N_29465,N_27068,N_27442);
nor U29466 (N_29466,N_27771,N_27496);
or U29467 (N_29467,N_28210,N_27658);
xnor U29468 (N_29468,N_28341,N_27070);
and U29469 (N_29469,N_28174,N_27248);
and U29470 (N_29470,N_28428,N_27652);
xnor U29471 (N_29471,N_27880,N_27404);
nor U29472 (N_29472,N_27157,N_27352);
xor U29473 (N_29473,N_27783,N_27631);
nor U29474 (N_29474,N_27017,N_27368);
or U29475 (N_29475,N_28401,N_28497);
nand U29476 (N_29476,N_27492,N_28180);
and U29477 (N_29477,N_27094,N_27622);
nand U29478 (N_29478,N_28203,N_27585);
or U29479 (N_29479,N_27225,N_27768);
nor U29480 (N_29480,N_27320,N_27674);
and U29481 (N_29481,N_27002,N_27381);
xnor U29482 (N_29482,N_28054,N_27708);
and U29483 (N_29483,N_28273,N_27702);
nor U29484 (N_29484,N_27766,N_28349);
and U29485 (N_29485,N_27024,N_27206);
nand U29486 (N_29486,N_27971,N_27134);
or U29487 (N_29487,N_27191,N_28095);
and U29488 (N_29488,N_28467,N_27231);
or U29489 (N_29489,N_27459,N_28303);
nor U29490 (N_29490,N_27583,N_27793);
xor U29491 (N_29491,N_27703,N_27935);
xnor U29492 (N_29492,N_27987,N_27195);
or U29493 (N_29493,N_27354,N_27300);
and U29494 (N_29494,N_27336,N_28001);
or U29495 (N_29495,N_28454,N_27271);
xor U29496 (N_29496,N_27177,N_27071);
xor U29497 (N_29497,N_28375,N_27004);
xor U29498 (N_29498,N_27637,N_27576);
nor U29499 (N_29499,N_27866,N_28202);
and U29500 (N_29500,N_28065,N_28189);
or U29501 (N_29501,N_28114,N_27923);
nor U29502 (N_29502,N_27356,N_28064);
and U29503 (N_29503,N_28320,N_27550);
and U29504 (N_29504,N_27014,N_28099);
nor U29505 (N_29505,N_28272,N_27169);
or U29506 (N_29506,N_27147,N_27172);
or U29507 (N_29507,N_27709,N_27472);
xnor U29508 (N_29508,N_27457,N_27521);
or U29509 (N_29509,N_27067,N_28192);
or U29510 (N_29510,N_27085,N_27259);
or U29511 (N_29511,N_28185,N_27526);
nand U29512 (N_29512,N_28186,N_28409);
or U29513 (N_29513,N_27476,N_27457);
and U29514 (N_29514,N_27561,N_28410);
nand U29515 (N_29515,N_28192,N_28311);
nand U29516 (N_29516,N_27773,N_27249);
nand U29517 (N_29517,N_27729,N_27196);
nand U29518 (N_29518,N_28145,N_27484);
nor U29519 (N_29519,N_28139,N_28030);
or U29520 (N_29520,N_27473,N_28391);
nor U29521 (N_29521,N_27363,N_27151);
and U29522 (N_29522,N_27464,N_27494);
or U29523 (N_29523,N_28468,N_27634);
and U29524 (N_29524,N_28070,N_27069);
and U29525 (N_29525,N_27018,N_28312);
nor U29526 (N_29526,N_27081,N_27833);
and U29527 (N_29527,N_27547,N_27566);
or U29528 (N_29528,N_27373,N_27052);
or U29529 (N_29529,N_27114,N_27798);
xor U29530 (N_29530,N_27669,N_27004);
and U29531 (N_29531,N_27744,N_27861);
nand U29532 (N_29532,N_27004,N_27245);
xor U29533 (N_29533,N_28436,N_28360);
nand U29534 (N_29534,N_27196,N_27998);
nor U29535 (N_29535,N_27625,N_27062);
and U29536 (N_29536,N_28120,N_27379);
and U29537 (N_29537,N_28312,N_27497);
nor U29538 (N_29538,N_28353,N_28498);
nor U29539 (N_29539,N_27651,N_28237);
xor U29540 (N_29540,N_27255,N_27601);
nor U29541 (N_29541,N_27519,N_27833);
nor U29542 (N_29542,N_28272,N_28016);
xor U29543 (N_29543,N_27316,N_28150);
or U29544 (N_29544,N_27941,N_27480);
or U29545 (N_29545,N_27586,N_27918);
xnor U29546 (N_29546,N_27768,N_28447);
nand U29547 (N_29547,N_28428,N_27383);
and U29548 (N_29548,N_28194,N_28220);
nand U29549 (N_29549,N_27208,N_28126);
and U29550 (N_29550,N_28075,N_28448);
xor U29551 (N_29551,N_27930,N_27887);
xnor U29552 (N_29552,N_28471,N_28381);
and U29553 (N_29553,N_27600,N_27673);
or U29554 (N_29554,N_27584,N_27214);
or U29555 (N_29555,N_27719,N_27269);
nand U29556 (N_29556,N_28000,N_28055);
nor U29557 (N_29557,N_27118,N_27177);
nor U29558 (N_29558,N_27200,N_27618);
or U29559 (N_29559,N_28025,N_27601);
nand U29560 (N_29560,N_27761,N_27154);
or U29561 (N_29561,N_27678,N_27224);
or U29562 (N_29562,N_27463,N_28248);
nand U29563 (N_29563,N_27229,N_28199);
nor U29564 (N_29564,N_27630,N_28196);
or U29565 (N_29565,N_28461,N_27104);
nand U29566 (N_29566,N_27548,N_28196);
nand U29567 (N_29567,N_27357,N_27716);
or U29568 (N_29568,N_28317,N_28055);
nand U29569 (N_29569,N_27184,N_28459);
or U29570 (N_29570,N_27964,N_27092);
nor U29571 (N_29571,N_27245,N_27749);
and U29572 (N_29572,N_28287,N_28345);
or U29573 (N_29573,N_27904,N_28422);
xnor U29574 (N_29574,N_28222,N_28050);
xor U29575 (N_29575,N_27101,N_27260);
nor U29576 (N_29576,N_27550,N_27933);
nor U29577 (N_29577,N_27579,N_27304);
xor U29578 (N_29578,N_27071,N_28305);
nand U29579 (N_29579,N_27441,N_27180);
and U29580 (N_29580,N_28279,N_27851);
nand U29581 (N_29581,N_27293,N_27589);
nor U29582 (N_29582,N_27608,N_28024);
xor U29583 (N_29583,N_27569,N_27252);
nand U29584 (N_29584,N_28050,N_27872);
and U29585 (N_29585,N_27297,N_27493);
or U29586 (N_29586,N_27184,N_27097);
and U29587 (N_29587,N_28296,N_27233);
nor U29588 (N_29588,N_27851,N_28206);
or U29589 (N_29589,N_27880,N_27467);
and U29590 (N_29590,N_27476,N_27400);
nand U29591 (N_29591,N_27289,N_27243);
nand U29592 (N_29592,N_27409,N_27146);
and U29593 (N_29593,N_27881,N_27282);
nand U29594 (N_29594,N_27177,N_27633);
nand U29595 (N_29595,N_27950,N_27107);
nor U29596 (N_29596,N_27156,N_27146);
xnor U29597 (N_29597,N_27156,N_28467);
and U29598 (N_29598,N_27712,N_27910);
nand U29599 (N_29599,N_27715,N_28173);
nor U29600 (N_29600,N_27563,N_27648);
and U29601 (N_29601,N_28078,N_28019);
and U29602 (N_29602,N_27998,N_27008);
and U29603 (N_29603,N_27853,N_27494);
and U29604 (N_29604,N_27304,N_28351);
or U29605 (N_29605,N_27173,N_27175);
nand U29606 (N_29606,N_27518,N_28191);
and U29607 (N_29607,N_27302,N_28128);
or U29608 (N_29608,N_27443,N_27052);
nand U29609 (N_29609,N_27542,N_27518);
nand U29610 (N_29610,N_27958,N_27850);
nor U29611 (N_29611,N_27113,N_27655);
nand U29612 (N_29612,N_27349,N_27279);
or U29613 (N_29613,N_27916,N_27769);
or U29614 (N_29614,N_27466,N_28083);
nand U29615 (N_29615,N_27546,N_27421);
xor U29616 (N_29616,N_27421,N_27805);
and U29617 (N_29617,N_27755,N_27783);
and U29618 (N_29618,N_27382,N_27362);
nand U29619 (N_29619,N_28050,N_27142);
nand U29620 (N_29620,N_27187,N_27417);
xnor U29621 (N_29621,N_28334,N_27999);
and U29622 (N_29622,N_27932,N_28000);
nand U29623 (N_29623,N_28101,N_27720);
and U29624 (N_29624,N_27455,N_27840);
nor U29625 (N_29625,N_27812,N_27545);
nor U29626 (N_29626,N_27205,N_27572);
or U29627 (N_29627,N_28358,N_27282);
nand U29628 (N_29628,N_27549,N_27220);
nand U29629 (N_29629,N_28179,N_27915);
nand U29630 (N_29630,N_27458,N_28134);
and U29631 (N_29631,N_27497,N_27652);
and U29632 (N_29632,N_27081,N_27921);
nor U29633 (N_29633,N_27283,N_28312);
nor U29634 (N_29634,N_27125,N_27520);
xnor U29635 (N_29635,N_27986,N_27287);
nand U29636 (N_29636,N_27064,N_27944);
or U29637 (N_29637,N_27216,N_27761);
nor U29638 (N_29638,N_27511,N_27228);
or U29639 (N_29639,N_27424,N_27514);
xnor U29640 (N_29640,N_27444,N_27884);
nor U29641 (N_29641,N_27817,N_28204);
nor U29642 (N_29642,N_28016,N_27316);
nor U29643 (N_29643,N_27528,N_27822);
nand U29644 (N_29644,N_28265,N_27965);
nor U29645 (N_29645,N_27082,N_27125);
or U29646 (N_29646,N_27483,N_28129);
or U29647 (N_29647,N_27523,N_28130);
or U29648 (N_29648,N_27677,N_27102);
nor U29649 (N_29649,N_27749,N_27041);
nand U29650 (N_29650,N_27186,N_27964);
nor U29651 (N_29651,N_27179,N_27147);
xnor U29652 (N_29652,N_28059,N_28104);
nor U29653 (N_29653,N_27316,N_27730);
nor U29654 (N_29654,N_28133,N_28290);
and U29655 (N_29655,N_28407,N_27157);
xor U29656 (N_29656,N_28256,N_27869);
nor U29657 (N_29657,N_27804,N_28299);
xnor U29658 (N_29658,N_27275,N_27794);
or U29659 (N_29659,N_27697,N_27766);
xnor U29660 (N_29660,N_28028,N_27567);
or U29661 (N_29661,N_27523,N_27455);
nand U29662 (N_29662,N_28472,N_27812);
nand U29663 (N_29663,N_28215,N_27751);
and U29664 (N_29664,N_28351,N_27655);
nor U29665 (N_29665,N_27594,N_28202);
xor U29666 (N_29666,N_27572,N_28486);
nor U29667 (N_29667,N_28030,N_28302);
nor U29668 (N_29668,N_28446,N_28487);
nor U29669 (N_29669,N_27157,N_28455);
nor U29670 (N_29670,N_27299,N_28284);
or U29671 (N_29671,N_27192,N_27198);
nand U29672 (N_29672,N_28209,N_27352);
or U29673 (N_29673,N_28064,N_28203);
xnor U29674 (N_29674,N_27379,N_27457);
nand U29675 (N_29675,N_27922,N_27171);
nand U29676 (N_29676,N_27324,N_27865);
or U29677 (N_29677,N_27854,N_27744);
xor U29678 (N_29678,N_27146,N_27802);
nor U29679 (N_29679,N_28051,N_27333);
nand U29680 (N_29680,N_27219,N_27690);
and U29681 (N_29681,N_27023,N_27004);
or U29682 (N_29682,N_27496,N_27301);
xor U29683 (N_29683,N_28409,N_28469);
and U29684 (N_29684,N_27725,N_28319);
and U29685 (N_29685,N_27399,N_27455);
nand U29686 (N_29686,N_27800,N_27217);
nand U29687 (N_29687,N_27328,N_28464);
nor U29688 (N_29688,N_27436,N_28417);
xnor U29689 (N_29689,N_28482,N_27356);
nand U29690 (N_29690,N_27392,N_27292);
and U29691 (N_29691,N_27558,N_27919);
xor U29692 (N_29692,N_28419,N_27308);
nand U29693 (N_29693,N_27780,N_27034);
nor U29694 (N_29694,N_27840,N_27333);
or U29695 (N_29695,N_27380,N_27323);
or U29696 (N_29696,N_28458,N_27339);
or U29697 (N_29697,N_27573,N_27237);
and U29698 (N_29698,N_27630,N_27084);
nand U29699 (N_29699,N_28022,N_27917);
xnor U29700 (N_29700,N_27036,N_27202);
nor U29701 (N_29701,N_28068,N_27686);
and U29702 (N_29702,N_27298,N_28322);
or U29703 (N_29703,N_28356,N_27626);
and U29704 (N_29704,N_27890,N_27393);
xor U29705 (N_29705,N_27942,N_27083);
xnor U29706 (N_29706,N_27813,N_27967);
and U29707 (N_29707,N_27433,N_27055);
xnor U29708 (N_29708,N_28279,N_28391);
nand U29709 (N_29709,N_28433,N_28365);
xnor U29710 (N_29710,N_28280,N_27548);
nor U29711 (N_29711,N_27988,N_28337);
nor U29712 (N_29712,N_28317,N_27222);
nor U29713 (N_29713,N_27107,N_27041);
nor U29714 (N_29714,N_28154,N_27593);
or U29715 (N_29715,N_28037,N_27563);
nor U29716 (N_29716,N_27325,N_27391);
and U29717 (N_29717,N_27042,N_28391);
and U29718 (N_29718,N_27934,N_27701);
and U29719 (N_29719,N_27295,N_28353);
or U29720 (N_29720,N_27403,N_27019);
and U29721 (N_29721,N_27193,N_27067);
nand U29722 (N_29722,N_27431,N_27748);
or U29723 (N_29723,N_27036,N_27775);
xnor U29724 (N_29724,N_27444,N_28270);
and U29725 (N_29725,N_28171,N_28044);
nand U29726 (N_29726,N_27978,N_27065);
or U29727 (N_29727,N_27579,N_27039);
nand U29728 (N_29728,N_27228,N_27585);
nand U29729 (N_29729,N_27117,N_27164);
and U29730 (N_29730,N_27219,N_27207);
and U29731 (N_29731,N_27500,N_28283);
and U29732 (N_29732,N_27936,N_27929);
and U29733 (N_29733,N_27922,N_28244);
or U29734 (N_29734,N_27217,N_27824);
nor U29735 (N_29735,N_27894,N_27935);
nand U29736 (N_29736,N_27430,N_27187);
or U29737 (N_29737,N_28237,N_28186);
nor U29738 (N_29738,N_28326,N_27298);
or U29739 (N_29739,N_28077,N_28091);
nor U29740 (N_29740,N_27958,N_28144);
or U29741 (N_29741,N_27628,N_27346);
and U29742 (N_29742,N_27698,N_27453);
xnor U29743 (N_29743,N_27595,N_27925);
or U29744 (N_29744,N_28230,N_27420);
and U29745 (N_29745,N_28427,N_27715);
or U29746 (N_29746,N_28451,N_27903);
nor U29747 (N_29747,N_28181,N_27206);
and U29748 (N_29748,N_28131,N_27151);
nand U29749 (N_29749,N_28456,N_27016);
xnor U29750 (N_29750,N_27471,N_27252);
and U29751 (N_29751,N_27756,N_27504);
and U29752 (N_29752,N_27873,N_27073);
and U29753 (N_29753,N_28067,N_28372);
or U29754 (N_29754,N_27771,N_28428);
or U29755 (N_29755,N_27891,N_27135);
and U29756 (N_29756,N_27730,N_27583);
or U29757 (N_29757,N_28409,N_27406);
or U29758 (N_29758,N_27174,N_27129);
and U29759 (N_29759,N_28065,N_27076);
and U29760 (N_29760,N_28407,N_28367);
and U29761 (N_29761,N_27963,N_27978);
xor U29762 (N_29762,N_28021,N_27429);
or U29763 (N_29763,N_27794,N_27499);
nor U29764 (N_29764,N_27267,N_27137);
nand U29765 (N_29765,N_27606,N_28376);
nor U29766 (N_29766,N_27929,N_28267);
or U29767 (N_29767,N_27291,N_27508);
or U29768 (N_29768,N_27119,N_27335);
and U29769 (N_29769,N_27538,N_27710);
xnor U29770 (N_29770,N_27991,N_27267);
xor U29771 (N_29771,N_28210,N_27788);
and U29772 (N_29772,N_27217,N_27209);
and U29773 (N_29773,N_27438,N_27304);
or U29774 (N_29774,N_28329,N_28450);
nand U29775 (N_29775,N_27323,N_27322);
xnor U29776 (N_29776,N_27403,N_27343);
and U29777 (N_29777,N_27751,N_28154);
nand U29778 (N_29778,N_27072,N_27646);
or U29779 (N_29779,N_27599,N_28162);
nor U29780 (N_29780,N_28455,N_28110);
and U29781 (N_29781,N_27087,N_27678);
nor U29782 (N_29782,N_27968,N_28461);
nand U29783 (N_29783,N_28253,N_28093);
nor U29784 (N_29784,N_28291,N_27851);
nor U29785 (N_29785,N_27343,N_27398);
xnor U29786 (N_29786,N_27491,N_27021);
nand U29787 (N_29787,N_27458,N_27345);
nand U29788 (N_29788,N_28354,N_28433);
xor U29789 (N_29789,N_27245,N_27863);
nand U29790 (N_29790,N_28238,N_27215);
nor U29791 (N_29791,N_27012,N_27753);
nand U29792 (N_29792,N_27993,N_27277);
and U29793 (N_29793,N_27689,N_28446);
nand U29794 (N_29794,N_27316,N_27642);
nand U29795 (N_29795,N_27674,N_28145);
and U29796 (N_29796,N_28249,N_28345);
or U29797 (N_29797,N_28444,N_27439);
and U29798 (N_29798,N_27178,N_27866);
or U29799 (N_29799,N_27605,N_28216);
nor U29800 (N_29800,N_27722,N_27279);
nor U29801 (N_29801,N_27021,N_27078);
nor U29802 (N_29802,N_27310,N_27729);
nand U29803 (N_29803,N_27553,N_27121);
xnor U29804 (N_29804,N_28304,N_27669);
or U29805 (N_29805,N_27664,N_27934);
and U29806 (N_29806,N_27952,N_28106);
nor U29807 (N_29807,N_28332,N_28129);
nand U29808 (N_29808,N_27347,N_27541);
and U29809 (N_29809,N_27160,N_27961);
or U29810 (N_29810,N_27223,N_27756);
or U29811 (N_29811,N_27201,N_27036);
nand U29812 (N_29812,N_27931,N_27922);
and U29813 (N_29813,N_28209,N_27546);
nor U29814 (N_29814,N_28344,N_27921);
and U29815 (N_29815,N_27858,N_27769);
and U29816 (N_29816,N_27164,N_27826);
xor U29817 (N_29817,N_28451,N_28493);
and U29818 (N_29818,N_28380,N_27639);
nand U29819 (N_29819,N_28198,N_27034);
nor U29820 (N_29820,N_27655,N_27937);
and U29821 (N_29821,N_27932,N_27908);
or U29822 (N_29822,N_27419,N_28470);
nor U29823 (N_29823,N_27215,N_27908);
nor U29824 (N_29824,N_27512,N_28121);
and U29825 (N_29825,N_27460,N_28483);
xnor U29826 (N_29826,N_27473,N_27311);
xor U29827 (N_29827,N_28004,N_27125);
nor U29828 (N_29828,N_28358,N_27740);
and U29829 (N_29829,N_27846,N_28483);
nor U29830 (N_29830,N_27227,N_27514);
xnor U29831 (N_29831,N_27733,N_27321);
xnor U29832 (N_29832,N_27114,N_27773);
or U29833 (N_29833,N_28406,N_27403);
and U29834 (N_29834,N_27701,N_27718);
or U29835 (N_29835,N_27316,N_27282);
xor U29836 (N_29836,N_27657,N_27521);
nand U29837 (N_29837,N_27379,N_27401);
or U29838 (N_29838,N_27292,N_27441);
nand U29839 (N_29839,N_27716,N_28171);
nand U29840 (N_29840,N_27821,N_28281);
and U29841 (N_29841,N_28444,N_27946);
xnor U29842 (N_29842,N_27922,N_27968);
and U29843 (N_29843,N_28046,N_28246);
nand U29844 (N_29844,N_28435,N_27423);
xnor U29845 (N_29845,N_27428,N_28209);
nand U29846 (N_29846,N_27951,N_27669);
xor U29847 (N_29847,N_28258,N_27969);
xor U29848 (N_29848,N_28283,N_28270);
xnor U29849 (N_29849,N_27202,N_28201);
xnor U29850 (N_29850,N_28480,N_27362);
nor U29851 (N_29851,N_27291,N_27795);
nand U29852 (N_29852,N_27747,N_28074);
and U29853 (N_29853,N_27976,N_28397);
and U29854 (N_29854,N_28078,N_27489);
xnor U29855 (N_29855,N_27543,N_28134);
nand U29856 (N_29856,N_27114,N_28392);
nor U29857 (N_29857,N_27859,N_27036);
nor U29858 (N_29858,N_27740,N_28000);
xor U29859 (N_29859,N_27461,N_27980);
xor U29860 (N_29860,N_27762,N_27730);
xor U29861 (N_29861,N_28132,N_27870);
or U29862 (N_29862,N_27037,N_28425);
nand U29863 (N_29863,N_27383,N_27471);
nor U29864 (N_29864,N_27957,N_27341);
and U29865 (N_29865,N_27024,N_27751);
or U29866 (N_29866,N_27522,N_27025);
xor U29867 (N_29867,N_27535,N_27295);
or U29868 (N_29868,N_28432,N_28126);
nor U29869 (N_29869,N_27332,N_27809);
nand U29870 (N_29870,N_27712,N_28481);
nand U29871 (N_29871,N_28221,N_27045);
and U29872 (N_29872,N_27545,N_28230);
nand U29873 (N_29873,N_27038,N_27751);
nor U29874 (N_29874,N_27178,N_28287);
and U29875 (N_29875,N_27973,N_27643);
xnor U29876 (N_29876,N_27671,N_28365);
and U29877 (N_29877,N_28375,N_27766);
nand U29878 (N_29878,N_28398,N_27045);
and U29879 (N_29879,N_27932,N_27968);
nor U29880 (N_29880,N_27509,N_28489);
xnor U29881 (N_29881,N_28253,N_28215);
nor U29882 (N_29882,N_27859,N_27682);
or U29883 (N_29883,N_27774,N_27090);
nand U29884 (N_29884,N_28241,N_27866);
xnor U29885 (N_29885,N_28246,N_27889);
nand U29886 (N_29886,N_28229,N_27873);
nor U29887 (N_29887,N_27823,N_28060);
xor U29888 (N_29888,N_27070,N_27236);
nor U29889 (N_29889,N_28024,N_28204);
or U29890 (N_29890,N_27677,N_27064);
xor U29891 (N_29891,N_27853,N_27192);
nand U29892 (N_29892,N_27445,N_27942);
xnor U29893 (N_29893,N_28163,N_28001);
or U29894 (N_29894,N_27521,N_27526);
or U29895 (N_29895,N_28404,N_27775);
xnor U29896 (N_29896,N_28128,N_28355);
xor U29897 (N_29897,N_27273,N_28064);
xor U29898 (N_29898,N_28412,N_27198);
and U29899 (N_29899,N_27020,N_27030);
xnor U29900 (N_29900,N_27229,N_27548);
nor U29901 (N_29901,N_27865,N_28227);
nor U29902 (N_29902,N_27870,N_27229);
or U29903 (N_29903,N_27083,N_27385);
xnor U29904 (N_29904,N_27378,N_27546);
or U29905 (N_29905,N_27644,N_28121);
or U29906 (N_29906,N_27890,N_27226);
xnor U29907 (N_29907,N_28027,N_27293);
xor U29908 (N_29908,N_27173,N_27751);
xor U29909 (N_29909,N_27856,N_28461);
nand U29910 (N_29910,N_28134,N_27422);
and U29911 (N_29911,N_28194,N_27707);
xnor U29912 (N_29912,N_27821,N_28276);
nand U29913 (N_29913,N_28220,N_28478);
and U29914 (N_29914,N_27972,N_27844);
xnor U29915 (N_29915,N_27270,N_27923);
xor U29916 (N_29916,N_27551,N_27033);
or U29917 (N_29917,N_27901,N_28116);
nor U29918 (N_29918,N_27574,N_28074);
nand U29919 (N_29919,N_27994,N_27257);
or U29920 (N_29920,N_28032,N_27002);
nand U29921 (N_29921,N_27651,N_28265);
and U29922 (N_29922,N_28425,N_27080);
and U29923 (N_29923,N_27146,N_28371);
nand U29924 (N_29924,N_28166,N_27469);
xnor U29925 (N_29925,N_28295,N_27176);
nor U29926 (N_29926,N_27867,N_27971);
or U29927 (N_29927,N_27845,N_27620);
and U29928 (N_29928,N_27232,N_28494);
nand U29929 (N_29929,N_27714,N_28365);
or U29930 (N_29930,N_28410,N_27693);
nor U29931 (N_29931,N_27654,N_28312);
and U29932 (N_29932,N_28393,N_27781);
nand U29933 (N_29933,N_28316,N_27461);
nor U29934 (N_29934,N_28305,N_28276);
nand U29935 (N_29935,N_28457,N_28490);
xnor U29936 (N_29936,N_27420,N_28269);
or U29937 (N_29937,N_27778,N_27540);
nor U29938 (N_29938,N_27175,N_27092);
xnor U29939 (N_29939,N_27863,N_28180);
or U29940 (N_29940,N_27386,N_27037);
and U29941 (N_29941,N_27894,N_27859);
and U29942 (N_29942,N_27051,N_27675);
xor U29943 (N_29943,N_27670,N_27841);
xnor U29944 (N_29944,N_27189,N_28359);
nand U29945 (N_29945,N_27553,N_27522);
nand U29946 (N_29946,N_27693,N_27292);
nand U29947 (N_29947,N_27604,N_28320);
nor U29948 (N_29948,N_28180,N_27009);
and U29949 (N_29949,N_27247,N_27285);
and U29950 (N_29950,N_28057,N_27778);
xnor U29951 (N_29951,N_27050,N_27613);
xnor U29952 (N_29952,N_27131,N_28030);
or U29953 (N_29953,N_28349,N_27263);
xor U29954 (N_29954,N_27201,N_27845);
xor U29955 (N_29955,N_27768,N_28153);
or U29956 (N_29956,N_28393,N_27865);
and U29957 (N_29957,N_27275,N_27429);
nor U29958 (N_29958,N_28487,N_28496);
or U29959 (N_29959,N_28176,N_28451);
xnor U29960 (N_29960,N_28429,N_27488);
nor U29961 (N_29961,N_27430,N_27571);
or U29962 (N_29962,N_27999,N_27627);
xor U29963 (N_29963,N_27697,N_27006);
xnor U29964 (N_29964,N_28056,N_27738);
xor U29965 (N_29965,N_27641,N_28399);
and U29966 (N_29966,N_27722,N_27431);
xor U29967 (N_29967,N_28495,N_27278);
or U29968 (N_29968,N_28182,N_27927);
or U29969 (N_29969,N_27193,N_28330);
nand U29970 (N_29970,N_27366,N_28360);
nand U29971 (N_29971,N_28276,N_27162);
and U29972 (N_29972,N_27346,N_28012);
or U29973 (N_29973,N_27990,N_27191);
xnor U29974 (N_29974,N_27111,N_27914);
and U29975 (N_29975,N_27949,N_27899);
xor U29976 (N_29976,N_28210,N_28390);
nand U29977 (N_29977,N_27845,N_27162);
and U29978 (N_29978,N_28380,N_28222);
xnor U29979 (N_29979,N_28252,N_27871);
nor U29980 (N_29980,N_28157,N_28455);
nor U29981 (N_29981,N_27292,N_27349);
and U29982 (N_29982,N_28360,N_28024);
nor U29983 (N_29983,N_27586,N_28435);
nor U29984 (N_29984,N_27490,N_27079);
nand U29985 (N_29985,N_27513,N_27447);
nor U29986 (N_29986,N_28245,N_27612);
nand U29987 (N_29987,N_27682,N_28253);
and U29988 (N_29988,N_28414,N_28434);
or U29989 (N_29989,N_27279,N_27835);
xnor U29990 (N_29990,N_27556,N_27910);
xor U29991 (N_29991,N_27883,N_27419);
and U29992 (N_29992,N_27016,N_28383);
or U29993 (N_29993,N_27351,N_27459);
nand U29994 (N_29994,N_27056,N_27516);
or U29995 (N_29995,N_27169,N_27540);
and U29996 (N_29996,N_28151,N_27630);
or U29997 (N_29997,N_27444,N_27751);
nor U29998 (N_29998,N_27881,N_27640);
xor U29999 (N_29999,N_27158,N_28438);
and UO_0 (O_0,N_28960,N_29018);
and UO_1 (O_1,N_28934,N_28644);
nor UO_2 (O_2,N_29714,N_28942);
nor UO_3 (O_3,N_29751,N_29229);
and UO_4 (O_4,N_29896,N_29130);
and UO_5 (O_5,N_29556,N_29511);
nand UO_6 (O_6,N_29155,N_28936);
nor UO_7 (O_7,N_28522,N_29030);
nor UO_8 (O_8,N_29231,N_28704);
nor UO_9 (O_9,N_29547,N_29303);
xor UO_10 (O_10,N_28844,N_29581);
nand UO_11 (O_11,N_29418,N_28684);
or UO_12 (O_12,N_29446,N_29333);
or UO_13 (O_13,N_28915,N_29572);
xor UO_14 (O_14,N_28845,N_29631);
and UO_15 (O_15,N_28618,N_29692);
nand UO_16 (O_16,N_29490,N_29072);
or UO_17 (O_17,N_29459,N_29887);
nand UO_18 (O_18,N_28948,N_29538);
or UO_19 (O_19,N_29386,N_29242);
nor UO_20 (O_20,N_28977,N_29080);
or UO_21 (O_21,N_28952,N_29010);
xor UO_22 (O_22,N_29008,N_28968);
or UO_23 (O_23,N_29148,N_29188);
nand UO_24 (O_24,N_28842,N_28790);
nand UO_25 (O_25,N_29644,N_28892);
and UO_26 (O_26,N_29639,N_28713);
nor UO_27 (O_27,N_29709,N_29756);
xor UO_28 (O_28,N_28871,N_29701);
or UO_29 (O_29,N_28819,N_29736);
nor UO_30 (O_30,N_29895,N_29795);
nand UO_31 (O_31,N_28873,N_28654);
and UO_32 (O_32,N_28885,N_28856);
or UO_33 (O_33,N_29510,N_29994);
nor UO_34 (O_34,N_28808,N_28578);
nand UO_35 (O_35,N_28610,N_29608);
xnor UO_36 (O_36,N_29611,N_29002);
xnor UO_37 (O_37,N_29554,N_29814);
nor UO_38 (O_38,N_29761,N_29367);
nor UO_39 (O_39,N_29657,N_29758);
or UO_40 (O_40,N_28553,N_29577);
nor UO_41 (O_41,N_28816,N_29175);
nor UO_42 (O_42,N_29413,N_28523);
and UO_43 (O_43,N_29810,N_28696);
or UO_44 (O_44,N_29889,N_29100);
or UO_45 (O_45,N_28539,N_29196);
nand UO_46 (O_46,N_29868,N_29444);
nand UO_47 (O_47,N_28920,N_28671);
xor UO_48 (O_48,N_29423,N_28529);
nor UO_49 (O_49,N_28812,N_29506);
and UO_50 (O_50,N_28966,N_29183);
or UO_51 (O_51,N_29278,N_29335);
and UO_52 (O_52,N_28983,N_28877);
or UO_53 (O_53,N_29304,N_28769);
nand UO_54 (O_54,N_28503,N_28643);
or UO_55 (O_55,N_28849,N_29266);
and UO_56 (O_56,N_28957,N_29001);
nor UO_57 (O_57,N_29797,N_28992);
or UO_58 (O_58,N_29660,N_29258);
and UO_59 (O_59,N_28917,N_29700);
and UO_60 (O_60,N_28520,N_28614);
nand UO_61 (O_61,N_28994,N_29762);
or UO_62 (O_62,N_29443,N_28758);
nand UO_63 (O_63,N_29450,N_29629);
and UO_64 (O_64,N_28649,N_28792);
nor UO_65 (O_65,N_28891,N_29414);
or UO_66 (O_66,N_28680,N_29673);
and UO_67 (O_67,N_28787,N_29993);
xor UO_68 (O_68,N_29293,N_29527);
nand UO_69 (O_69,N_29697,N_29056);
and UO_70 (O_70,N_28878,N_29964);
xor UO_71 (O_71,N_29533,N_29383);
xnor UO_72 (O_72,N_29058,N_29416);
and UO_73 (O_73,N_29238,N_28552);
or UO_74 (O_74,N_28574,N_28551);
or UO_75 (O_75,N_29967,N_29374);
and UO_76 (O_76,N_29234,N_29957);
nor UO_77 (O_77,N_29358,N_29310);
xor UO_78 (O_78,N_29366,N_29775);
and UO_79 (O_79,N_29865,N_28987);
and UO_80 (O_80,N_29060,N_29405);
and UO_81 (O_81,N_29212,N_29388);
nor UO_82 (O_82,N_28733,N_29997);
nand UO_83 (O_83,N_28521,N_29634);
nor UO_84 (O_84,N_29926,N_29636);
xnor UO_85 (O_85,N_29479,N_28586);
nand UO_86 (O_86,N_28558,N_28918);
nor UO_87 (O_87,N_29544,N_28827);
nor UO_88 (O_88,N_29771,N_29850);
nand UO_89 (O_89,N_29866,N_29815);
nand UO_90 (O_90,N_28867,N_29355);
or UO_91 (O_91,N_29471,N_29017);
nor UO_92 (O_92,N_29228,N_29842);
nor UO_93 (O_93,N_29772,N_29539);
xor UO_94 (O_94,N_29792,N_28774);
and UO_95 (O_95,N_29821,N_29637);
nor UO_96 (O_96,N_29859,N_29050);
or UO_97 (O_97,N_28836,N_29504);
nand UO_98 (O_98,N_29723,N_28533);
nor UO_99 (O_99,N_29667,N_29354);
nand UO_100 (O_100,N_29939,N_28985);
nand UO_101 (O_101,N_29064,N_29166);
and UO_102 (O_102,N_29400,N_29919);
and UO_103 (O_103,N_28795,N_28595);
nand UO_104 (O_104,N_29077,N_29147);
nand UO_105 (O_105,N_29104,N_29257);
xor UO_106 (O_106,N_28548,N_29301);
and UO_107 (O_107,N_28638,N_29208);
nand UO_108 (O_108,N_28879,N_29733);
nor UO_109 (O_109,N_29852,N_29916);
nor UO_110 (O_110,N_28720,N_29051);
or UO_111 (O_111,N_28530,N_28932);
xnor UO_112 (O_112,N_29747,N_29805);
and UO_113 (O_113,N_29809,N_28993);
xnor UO_114 (O_114,N_29171,N_29528);
xnor UO_115 (O_115,N_28974,N_29913);
or UO_116 (O_116,N_28516,N_29774);
and UO_117 (O_117,N_28597,N_28954);
nand UO_118 (O_118,N_29296,N_29728);
or UO_119 (O_119,N_28799,N_29676);
and UO_120 (O_120,N_28658,N_29904);
nor UO_121 (O_121,N_29176,N_29543);
xor UO_122 (O_122,N_28837,N_29849);
and UO_123 (O_123,N_28961,N_29575);
nor UO_124 (O_124,N_29128,N_29055);
and UO_125 (O_125,N_29584,N_28901);
nand UO_126 (O_126,N_29937,N_28701);
nor UO_127 (O_127,N_29131,N_29947);
nand UO_128 (O_128,N_29347,N_28681);
or UO_129 (O_129,N_29189,N_29067);
xnor UO_130 (O_130,N_28576,N_29779);
nand UO_131 (O_131,N_28645,N_28828);
or UO_132 (O_132,N_29605,N_29826);
or UO_133 (O_133,N_28880,N_28661);
xnor UO_134 (O_134,N_29541,N_29401);
and UO_135 (O_135,N_29698,N_29380);
nand UO_136 (O_136,N_29163,N_29844);
or UO_137 (O_137,N_29760,N_28545);
xor UO_138 (O_138,N_28870,N_28935);
and UO_139 (O_139,N_28674,N_29499);
and UO_140 (O_140,N_28986,N_28855);
xor UO_141 (O_141,N_29284,N_28949);
and UO_142 (O_142,N_29206,N_29936);
xor UO_143 (O_143,N_29759,N_28707);
xnor UO_144 (O_144,N_29734,N_29118);
nand UO_145 (O_145,N_28928,N_29226);
or UO_146 (O_146,N_28746,N_29306);
xor UO_147 (O_147,N_28741,N_29819);
xor UO_148 (O_148,N_28969,N_29940);
and UO_149 (O_149,N_29315,N_28889);
and UO_150 (O_150,N_29363,N_29594);
xor UO_151 (O_151,N_29856,N_28923);
xnor UO_152 (O_152,N_29573,N_28927);
nand UO_153 (O_153,N_29591,N_29551);
or UO_154 (O_154,N_28629,N_28862);
nand UO_155 (O_155,N_29465,N_29861);
xnor UO_156 (O_156,N_28998,N_29715);
and UO_157 (O_157,N_28738,N_29890);
nand UO_158 (O_158,N_28921,N_29767);
nand UO_159 (O_159,N_28951,N_28822);
xor UO_160 (O_160,N_29616,N_29717);
nor UO_161 (O_161,N_29683,N_29390);
and UO_162 (O_162,N_28639,N_28538);
xnor UO_163 (O_163,N_28834,N_29567);
nand UO_164 (O_164,N_28564,N_29518);
and UO_165 (O_165,N_29879,N_28874);
xor UO_166 (O_166,N_28515,N_28630);
and UO_167 (O_167,N_28734,N_29839);
nor UO_168 (O_168,N_29144,N_29827);
or UO_169 (O_169,N_29409,N_29113);
nand UO_170 (O_170,N_29508,N_28710);
and UO_171 (O_171,N_28956,N_28668);
nand UO_172 (O_172,N_29691,N_29903);
and UO_173 (O_173,N_28852,N_29353);
xor UO_174 (O_174,N_29763,N_29449);
nand UO_175 (O_175,N_29312,N_29180);
and UO_176 (O_176,N_29738,N_29812);
nor UO_177 (O_177,N_29299,N_28579);
nor UO_178 (O_178,N_29534,N_29387);
and UO_179 (O_179,N_29106,N_29251);
xnor UO_180 (O_180,N_29600,N_28762);
nor UO_181 (O_181,N_29513,N_28943);
xor UO_182 (O_182,N_29433,N_29472);
nor UO_183 (O_183,N_29599,N_29192);
or UO_184 (O_184,N_29469,N_29702);
nor UO_185 (O_185,N_29794,N_28781);
xor UO_186 (O_186,N_29870,N_29776);
nand UO_187 (O_187,N_28692,N_29824);
or UO_188 (O_188,N_29960,N_29976);
and UO_189 (O_189,N_28785,N_28544);
xor UO_190 (O_190,N_28648,N_29352);
xor UO_191 (O_191,N_29005,N_29341);
nor UO_192 (O_192,N_29343,N_28970);
nand UO_193 (O_193,N_28640,N_29796);
nor UO_194 (O_194,N_29754,N_29090);
or UO_195 (O_195,N_29791,N_29329);
nand UO_196 (O_196,N_28688,N_29091);
and UO_197 (O_197,N_28670,N_29901);
nor UO_198 (O_198,N_29378,N_29029);
or UO_199 (O_199,N_28978,N_29381);
xor UO_200 (O_200,N_29984,N_29831);
nand UO_201 (O_201,N_28624,N_28582);
nand UO_202 (O_202,N_29942,N_29597);
nor UO_203 (O_203,N_29781,N_29127);
xnor UO_204 (O_204,N_29991,N_29954);
nand UO_205 (O_205,N_29654,N_28612);
nand UO_206 (O_206,N_29068,N_28659);
xnor UO_207 (O_207,N_29019,N_29275);
xnor UO_208 (O_208,N_28991,N_28646);
and UO_209 (O_209,N_29421,N_28601);
nand UO_210 (O_210,N_29169,N_28726);
xor UO_211 (O_211,N_29439,N_29497);
nand UO_212 (O_212,N_28611,N_28673);
nand UO_213 (O_213,N_29972,N_29834);
or UO_214 (O_214,N_28633,N_29495);
nand UO_215 (O_215,N_29862,N_28851);
nor UO_216 (O_216,N_29998,N_28818);
xnor UO_217 (O_217,N_28771,N_28814);
and UO_218 (O_218,N_29888,N_28660);
or UO_219 (O_219,N_29272,N_29959);
nand UO_220 (O_220,N_29620,N_29004);
nor UO_221 (O_221,N_29243,N_29607);
nand UO_222 (O_222,N_29201,N_29992);
nand UO_223 (O_223,N_29370,N_28759);
and UO_224 (O_224,N_29951,N_28667);
nor UO_225 (O_225,N_29837,N_29097);
or UO_226 (O_226,N_29209,N_28541);
and UO_227 (O_227,N_28984,N_28950);
xnor UO_228 (O_228,N_28619,N_29489);
nor UO_229 (O_229,N_29109,N_28575);
nand UO_230 (O_230,N_28568,N_29222);
xor UO_231 (O_231,N_29034,N_28797);
nand UO_232 (O_232,N_29143,N_29501);
nand UO_233 (O_233,N_28534,N_28693);
or UO_234 (O_234,N_29033,N_29777);
xor UO_235 (O_235,N_28922,N_29220);
nand UO_236 (O_236,N_28897,N_29214);
nor UO_237 (O_237,N_28859,N_29855);
or UO_238 (O_238,N_29811,N_29339);
nor UO_239 (O_239,N_29632,N_29485);
nor UO_240 (O_240,N_29788,N_29987);
and UO_241 (O_241,N_29360,N_29535);
xnor UO_242 (O_242,N_28846,N_29086);
and UO_243 (O_243,N_29053,N_29571);
nor UO_244 (O_244,N_28823,N_28953);
and UO_245 (O_245,N_29117,N_28603);
xor UO_246 (O_246,N_29142,N_29289);
or UO_247 (O_247,N_28714,N_29872);
nand UO_248 (O_248,N_28702,N_29045);
and UO_249 (O_249,N_29021,N_28898);
or UO_250 (O_250,N_29248,N_29198);
xnor UO_251 (O_251,N_29379,N_29741);
nand UO_252 (O_252,N_29269,N_29912);
nand UO_253 (O_253,N_28802,N_28571);
and UO_254 (O_254,N_29268,N_29059);
xor UO_255 (O_255,N_29087,N_29375);
and UO_256 (O_256,N_29442,N_29566);
or UO_257 (O_257,N_28708,N_28860);
or UO_258 (O_258,N_29372,N_29704);
and UO_259 (O_259,N_28524,N_29665);
or UO_260 (O_260,N_29563,N_28941);
or UO_261 (O_261,N_29292,N_29536);
xor UO_262 (O_262,N_29769,N_29641);
or UO_263 (O_263,N_29349,N_29822);
nor UO_264 (O_264,N_29848,N_28752);
nor UO_265 (O_265,N_29402,N_29316);
nor UO_266 (O_266,N_28596,N_28755);
or UO_267 (O_267,N_29786,N_29156);
xor UO_268 (O_268,N_28532,N_28697);
xor UO_269 (O_269,N_29914,N_28606);
nand UO_270 (O_270,N_28770,N_29902);
and UO_271 (O_271,N_29807,N_29419);
nand UO_272 (O_272,N_29340,N_29748);
nor UO_273 (O_273,N_28685,N_28763);
nand UO_274 (O_274,N_28919,N_29863);
nor UO_275 (O_275,N_28735,N_29677);
nand UO_276 (O_276,N_29832,N_29925);
nand UO_277 (O_277,N_29186,N_29217);
nor UO_278 (O_278,N_29125,N_29049);
and UO_279 (O_279,N_29598,N_29294);
xor UO_280 (O_280,N_29435,N_28662);
nand UO_281 (O_281,N_29491,N_29083);
nand UO_282 (O_282,N_29194,N_29860);
nand UO_283 (O_283,N_29445,N_29035);
nand UO_284 (O_284,N_29514,N_29195);
or UO_285 (O_285,N_28514,N_29966);
nor UO_286 (O_286,N_29393,N_29494);
nor UO_287 (O_287,N_28937,N_28536);
and UO_288 (O_288,N_29202,N_29927);
nand UO_289 (O_289,N_29219,N_28925);
xnor UO_290 (O_290,N_29773,N_28890);
nand UO_291 (O_291,N_29197,N_29725);
and UO_292 (O_292,N_28519,N_29894);
nor UO_293 (O_293,N_29505,N_29564);
and UO_294 (O_294,N_29530,N_29980);
or UO_295 (O_295,N_29922,N_28604);
xor UO_296 (O_296,N_29448,N_29643);
nor UO_297 (O_297,N_29264,N_28929);
nor UO_298 (O_298,N_28881,N_29282);
xnor UO_299 (O_299,N_29707,N_29230);
and UO_300 (O_300,N_28700,N_28506);
xor UO_301 (O_301,N_28945,N_28587);
or UO_302 (O_302,N_29580,N_28768);
xnor UO_303 (O_303,N_29256,N_28793);
nor UO_304 (O_304,N_28843,N_29813);
nor UO_305 (O_305,N_29119,N_29182);
nand UO_306 (O_306,N_29502,N_29766);
and UO_307 (O_307,N_29377,N_29908);
nand UO_308 (O_308,N_28636,N_29975);
nor UO_309 (O_309,N_29199,N_29949);
xnor UO_310 (O_310,N_29311,N_29675);
xor UO_311 (O_311,N_29108,N_28613);
nand UO_312 (O_312,N_29968,N_28589);
nor UO_313 (O_313,N_28902,N_29417);
xor UO_314 (O_314,N_28504,N_29604);
nand UO_315 (O_315,N_28971,N_29606);
and UO_316 (O_316,N_29524,N_29503);
or UO_317 (O_317,N_29924,N_29619);
or UO_318 (O_318,N_29670,N_29568);
nand UO_319 (O_319,N_29962,N_28806);
or UO_320 (O_320,N_29693,N_29730);
nor UO_321 (O_321,N_29999,N_28657);
nor UO_322 (O_322,N_28537,N_29874);
xor UO_323 (O_323,N_29955,N_29732);
and UO_324 (O_324,N_29408,N_29820);
and UO_325 (O_325,N_28989,N_29941);
nor UO_326 (O_326,N_29240,N_29977);
nor UO_327 (O_327,N_28801,N_28866);
and UO_328 (O_328,N_28800,N_29261);
xnor UO_329 (O_329,N_28690,N_28794);
and UO_330 (O_330,N_29337,N_29368);
nand UO_331 (O_331,N_28562,N_29618);
and UO_332 (O_332,N_28655,N_28711);
and UO_333 (O_333,N_29254,N_29274);
and UO_334 (O_334,N_29162,N_29878);
nor UO_335 (O_335,N_29037,N_28543);
nand UO_336 (O_336,N_29237,N_29043);
xnor UO_337 (O_337,N_28507,N_29559);
and UO_338 (O_338,N_29244,N_29308);
and UO_339 (O_339,N_29114,N_29875);
xnor UO_340 (O_340,N_29120,N_29746);
nor UO_341 (O_341,N_29094,N_28815);
or UO_342 (O_342,N_28678,N_29473);
nand UO_343 (O_343,N_29046,N_28577);
and UO_344 (O_344,N_28739,N_29453);
nand UO_345 (O_345,N_29107,N_29138);
and UO_346 (O_346,N_29345,N_29829);
and UO_347 (O_347,N_28566,N_29519);
nand UO_348 (O_348,N_28627,N_29079);
nand UO_349 (O_349,N_29398,N_28924);
or UO_350 (O_350,N_29688,N_29552);
xnor UO_351 (O_351,N_28740,N_29057);
and UO_352 (O_352,N_29731,N_29253);
nor UO_353 (O_353,N_29415,N_28729);
and UO_354 (O_354,N_29578,N_29458);
and UO_355 (O_355,N_29656,N_29307);
nand UO_356 (O_356,N_29655,N_28912);
or UO_357 (O_357,N_29481,N_29394);
xor UO_358 (O_358,N_28620,N_28930);
or UO_359 (O_359,N_28505,N_29235);
nor UO_360 (O_360,N_28663,N_28683);
xor UO_361 (O_361,N_29883,N_29135);
nor UO_362 (O_362,N_29215,N_29540);
xor UO_363 (O_363,N_29082,N_29323);
and UO_364 (O_364,N_29102,N_29074);
and UO_365 (O_365,N_28625,N_29392);
or UO_366 (O_366,N_28725,N_29297);
nand UO_367 (O_367,N_29800,N_29515);
or UO_368 (O_368,N_29396,N_29092);
xnor UO_369 (O_369,N_29140,N_29406);
nand UO_370 (O_370,N_29854,N_29262);
nor UO_371 (O_371,N_28580,N_29016);
xor UO_372 (O_372,N_28753,N_29790);
nor UO_373 (O_373,N_28996,N_29252);
and UO_374 (O_374,N_28841,N_29298);
or UO_375 (O_375,N_29684,N_29950);
xor UO_376 (O_376,N_29526,N_29451);
xnor UO_377 (O_377,N_29151,N_28803);
nor UO_378 (O_378,N_29179,N_29174);
xnor UO_379 (O_379,N_29752,N_29646);
xnor UO_380 (O_380,N_28776,N_29134);
nand UO_381 (O_381,N_29793,N_29427);
nand UO_382 (O_382,N_28981,N_28900);
nand UO_383 (O_383,N_29545,N_29084);
and UO_384 (O_384,N_29601,N_28672);
nor UO_385 (O_385,N_29522,N_29953);
nor UO_386 (O_386,N_28807,N_28896);
nand UO_387 (O_387,N_29468,N_29236);
or UO_388 (O_388,N_28581,N_28590);
or UO_389 (O_389,N_29757,N_28913);
xnor UO_390 (O_390,N_29893,N_28691);
xnor UO_391 (O_391,N_29012,N_28825);
xnor UO_392 (O_392,N_29085,N_28557);
xnor UO_393 (O_393,N_29132,N_28591);
and UO_394 (O_394,N_29466,N_29098);
or UO_395 (O_395,N_29024,N_28911);
xor UO_396 (O_396,N_29934,N_29227);
nand UO_397 (O_397,N_29020,N_29452);
and UO_398 (O_398,N_28742,N_29753);
nand UO_399 (O_399,N_29054,N_29270);
and UO_400 (O_400,N_29165,N_28748);
nor UO_401 (O_401,N_29322,N_28997);
and UO_402 (O_402,N_28546,N_29283);
nor UO_403 (O_403,N_28567,N_28958);
nand UO_404 (O_404,N_29350,N_29042);
nand UO_405 (O_405,N_28865,N_29721);
nand UO_406 (O_406,N_28626,N_28869);
and UO_407 (O_407,N_28829,N_28513);
or UO_408 (O_408,N_28549,N_29477);
nor UO_409 (O_409,N_29787,N_28926);
or UO_410 (O_410,N_29898,N_29317);
nor UO_411 (O_411,N_28973,N_28511);
nand UO_412 (O_412,N_28631,N_28868);
nand UO_413 (O_413,N_29007,N_29213);
xor UO_414 (O_414,N_29089,N_29716);
and UO_415 (O_415,N_29770,N_29447);
and UO_416 (O_416,N_29205,N_29133);
xnor UO_417 (O_417,N_29300,N_29560);
xnor UO_418 (O_418,N_28585,N_29263);
nor UO_419 (O_419,N_29804,N_28717);
nor UO_420 (O_420,N_29152,N_29403);
or UO_421 (O_421,N_29146,N_29886);
nand UO_422 (O_422,N_29687,N_28850);
and UO_423 (O_423,N_29330,N_29410);
xnor UO_424 (O_424,N_29871,N_29935);
or UO_425 (O_425,N_29441,N_29905);
nor UO_426 (O_426,N_28811,N_29595);
nor UO_427 (O_427,N_28675,N_29036);
and UO_428 (O_428,N_29173,N_28838);
nand UO_429 (O_429,N_28709,N_28602);
xnor UO_430 (O_430,N_29614,N_29295);
and UO_431 (O_431,N_29621,N_28666);
xor UO_432 (O_432,N_28689,N_29642);
nor UO_433 (O_433,N_29562,N_29153);
and UO_434 (O_434,N_28599,N_29718);
nor UO_435 (O_435,N_29255,N_29429);
and UO_436 (O_436,N_28664,N_29145);
xnor UO_437 (O_437,N_28605,N_29267);
and UO_438 (O_438,N_28723,N_28583);
or UO_439 (O_439,N_29320,N_29063);
or UO_440 (O_440,N_29764,N_28528);
xnor UO_441 (O_441,N_29755,N_29588);
xnor UO_442 (O_442,N_29995,N_29900);
or UO_443 (O_443,N_28903,N_29799);
nor UO_444 (O_444,N_28616,N_28854);
nor UO_445 (O_445,N_28750,N_29585);
nand UO_446 (O_446,N_29626,N_28999);
and UO_447 (O_447,N_29187,N_28563);
or UO_448 (O_448,N_29498,N_28731);
or UO_449 (O_449,N_29703,N_29101);
xnor UO_450 (O_450,N_29280,N_28550);
xnor UO_451 (O_451,N_29455,N_29603);
and UO_452 (O_452,N_28547,N_29464);
xnor UO_453 (O_453,N_29635,N_28712);
nor UO_454 (O_454,N_29440,N_29407);
nand UO_455 (O_455,N_29332,N_28847);
nor UO_456 (O_456,N_29149,N_29897);
or UO_457 (O_457,N_29137,N_28882);
or UO_458 (O_458,N_29110,N_29789);
xnor UO_459 (O_459,N_29369,N_29589);
or UO_460 (O_460,N_29853,N_28510);
xnor UO_461 (O_461,N_29742,N_29425);
and UO_462 (O_462,N_29570,N_29930);
nor UO_463 (O_463,N_28560,N_29389);
and UO_464 (O_464,N_28526,N_29052);
nor UO_465 (O_465,N_29743,N_29663);
nor UO_466 (O_466,N_29287,N_29139);
xor UO_467 (O_467,N_29361,N_28780);
xnor UO_468 (O_468,N_29348,N_29136);
nand UO_469 (O_469,N_29129,N_29044);
and UO_470 (O_470,N_29487,N_28863);
xor UO_471 (O_471,N_28905,N_29432);
nand UO_472 (O_472,N_29249,N_29633);
nand UO_473 (O_473,N_29971,N_29845);
and UO_474 (O_474,N_29190,N_29918);
and UO_475 (O_475,N_29668,N_28652);
xnor UO_476 (O_476,N_29482,N_29729);
or UO_477 (O_477,N_28588,N_29899);
nand UO_478 (O_478,N_29986,N_29362);
nor UO_479 (O_479,N_28721,N_29661);
nand UO_480 (O_480,N_29509,N_28669);
and UO_481 (O_481,N_29672,N_28884);
and UO_482 (O_482,N_29877,N_29630);
nor UO_483 (O_483,N_29193,N_29088);
and UO_484 (O_484,N_29719,N_29241);
xor UO_485 (O_485,N_29027,N_28817);
xnor UO_486 (O_486,N_29828,N_29923);
and UO_487 (O_487,N_29989,N_29111);
and UO_488 (O_488,N_28724,N_28910);
or UO_489 (O_489,N_29325,N_29569);
nand UO_490 (O_490,N_29124,N_28955);
xor UO_491 (O_491,N_29346,N_29404);
and UO_492 (O_492,N_29365,N_29537);
and UO_493 (O_493,N_28858,N_28760);
and UO_494 (O_494,N_29679,N_29070);
nand UO_495 (O_495,N_29517,N_28650);
nand UO_496 (O_496,N_29061,N_28786);
xnor UO_497 (O_497,N_29483,N_29265);
xor UO_498 (O_498,N_29973,N_29022);
or UO_499 (O_499,N_29470,N_28569);
and UO_500 (O_500,N_29833,N_28775);
and UO_501 (O_501,N_28699,N_28635);
or UO_502 (O_502,N_28833,N_28593);
nand UO_503 (O_503,N_28682,N_29671);
xnor UO_504 (O_504,N_29579,N_29737);
and UO_505 (O_505,N_28964,N_29069);
or UO_506 (O_506,N_29945,N_29529);
and UO_507 (O_507,N_29512,N_29424);
nand UO_508 (O_508,N_29028,N_28933);
nand UO_509 (O_509,N_28764,N_29210);
xor UO_510 (O_510,N_28535,N_29159);
and UO_511 (O_511,N_28813,N_29553);
nand UO_512 (O_512,N_29768,N_29956);
or UO_513 (O_513,N_29288,N_29115);
nand UO_514 (O_514,N_28540,N_28939);
and UO_515 (O_515,N_29457,N_29395);
nor UO_516 (O_516,N_29938,N_28899);
or UO_517 (O_517,N_28600,N_28784);
or UO_518 (O_518,N_28779,N_28963);
or UO_519 (O_519,N_28820,N_28778);
nor UO_520 (O_520,N_28621,N_28694);
and UO_521 (O_521,N_28853,N_28908);
nand UO_522 (O_522,N_28608,N_29801);
xnor UO_523 (O_523,N_29961,N_28687);
or UO_524 (O_524,N_28722,N_29203);
or UO_525 (O_525,N_29281,N_28745);
xnor UO_526 (O_526,N_28570,N_29694);
nor UO_527 (O_527,N_29682,N_28531);
xnor UO_528 (O_528,N_29931,N_29873);
nor UO_529 (O_529,N_28502,N_29981);
nand UO_530 (O_530,N_29699,N_29123);
and UO_531 (O_531,N_28517,N_29817);
xnor UO_532 (O_532,N_29548,N_28525);
and UO_533 (O_533,N_28761,N_29958);
xnor UO_534 (O_534,N_29532,N_28572);
and UO_535 (O_535,N_28573,N_29071);
nand UO_536 (O_536,N_29836,N_28556);
xnor UO_537 (O_537,N_29891,N_29011);
or UO_538 (O_538,N_29461,N_29590);
or UO_539 (O_539,N_28959,N_29550);
and UO_540 (O_540,N_29041,N_29014);
nand UO_541 (O_541,N_29200,N_28665);
nand UO_542 (O_542,N_29625,N_29397);
or UO_543 (O_543,N_29979,N_28904);
nor UO_544 (O_544,N_29239,N_28783);
xor UO_545 (O_545,N_28861,N_29917);
xor UO_546 (O_546,N_28979,N_28864);
nor UO_547 (O_547,N_29969,N_28821);
nand UO_548 (O_548,N_29876,N_28757);
or UO_549 (O_549,N_29765,N_28743);
nor UO_550 (O_550,N_29224,N_28791);
nor UO_551 (O_551,N_29066,N_29841);
and UO_552 (O_552,N_29710,N_28512);
and UO_553 (O_553,N_29778,N_29420);
nor UO_554 (O_554,N_29467,N_29664);
nand UO_555 (O_555,N_28848,N_28632);
nor UO_556 (O_556,N_29290,N_29546);
xor UO_557 (O_557,N_28893,N_29009);
nand UO_558 (O_558,N_29640,N_28796);
nand UO_559 (O_559,N_29689,N_29740);
and UO_560 (O_560,N_28831,N_29627);
and UO_561 (O_561,N_29726,N_29434);
and UO_562 (O_562,N_29150,N_28767);
nor UO_563 (O_563,N_29520,N_29326);
or UO_564 (O_564,N_28906,N_29218);
nand UO_565 (O_565,N_29232,N_28886);
xnor UO_566 (O_566,N_29516,N_29484);
xnor UO_567 (O_567,N_28501,N_28876);
and UO_568 (O_568,N_29031,N_29624);
nand UO_569 (O_569,N_28565,N_29185);
xor UO_570 (O_570,N_29909,N_29221);
nor UO_571 (O_571,N_28940,N_29475);
nor UO_572 (O_572,N_28653,N_29920);
nor UO_573 (O_573,N_29065,N_29858);
or UO_574 (O_574,N_29096,N_28705);
or UO_575 (O_575,N_28615,N_28656);
nor UO_576 (O_576,N_29696,N_28500);
xnor UO_577 (O_577,N_29040,N_29602);
or UO_578 (O_578,N_28598,N_29026);
and UO_579 (O_579,N_28609,N_29076);
and UO_580 (O_580,N_29160,N_29430);
or UO_581 (O_581,N_29158,N_29233);
nand UO_582 (O_582,N_29384,N_29492);
or UO_583 (O_583,N_28766,N_29783);
nor UO_584 (O_584,N_29674,N_29869);
and UO_585 (O_585,N_28698,N_29431);
or UO_586 (O_586,N_29780,N_29613);
xor UO_587 (O_587,N_29932,N_29121);
xor UO_588 (O_588,N_29302,N_28832);
nand UO_589 (O_589,N_29460,N_29686);
xor UO_590 (O_590,N_28839,N_29259);
or UO_591 (O_591,N_28727,N_29816);
or UO_592 (O_592,N_29116,N_28810);
or UO_593 (O_593,N_28875,N_29474);
or UO_594 (O_594,N_29105,N_29685);
nor UO_595 (O_595,N_29652,N_29648);
nor UO_596 (O_596,N_28982,N_29610);
nand UO_597 (O_597,N_28895,N_29892);
or UO_598 (O_598,N_28990,N_29750);
nand UO_599 (O_599,N_29708,N_29593);
xor UO_600 (O_600,N_28772,N_29319);
nand UO_601 (O_601,N_29279,N_29542);
and UO_602 (O_602,N_28972,N_28527);
and UO_603 (O_603,N_29921,N_29411);
and UO_604 (O_604,N_29802,N_29982);
and UO_605 (O_605,N_28555,N_29880);
or UO_606 (O_606,N_29713,N_29662);
xnor UO_607 (O_607,N_29929,N_28988);
nor UO_608 (O_608,N_29612,N_29706);
and UO_609 (O_609,N_28715,N_29285);
and UO_610 (O_610,N_29276,N_28686);
and UO_611 (O_611,N_28773,N_28508);
nor UO_612 (O_612,N_29745,N_29669);
or UO_613 (O_613,N_29985,N_29628);
nand UO_614 (O_614,N_29565,N_29587);
nand UO_615 (O_615,N_29586,N_29032);
or UO_616 (O_616,N_29735,N_28830);
or UO_617 (O_617,N_29617,N_29561);
or UO_618 (O_618,N_29651,N_28938);
nand UO_619 (O_619,N_29507,N_29609);
or UO_620 (O_620,N_29006,N_29364);
xnor UO_621 (O_621,N_29583,N_28518);
xnor UO_622 (O_622,N_28736,N_28931);
xnor UO_623 (O_623,N_28679,N_29681);
xnor UO_624 (O_624,N_29531,N_28909);
nor UO_625 (O_625,N_29313,N_29650);
or UO_626 (O_626,N_28634,N_29486);
or UO_627 (O_627,N_28995,N_29965);
or UO_628 (O_628,N_29328,N_28751);
xnor UO_629 (O_629,N_29023,N_28914);
nand UO_630 (O_630,N_28676,N_28789);
or UO_631 (O_631,N_29334,N_29371);
or UO_632 (O_632,N_29557,N_29373);
nor UO_633 (O_633,N_28809,N_29164);
nand UO_634 (O_634,N_28840,N_28980);
and UO_635 (O_635,N_28622,N_29141);
nand UO_636 (O_636,N_29331,N_29178);
and UO_637 (O_637,N_29952,N_29412);
nor UO_638 (O_638,N_28732,N_29666);
and UO_639 (O_639,N_29399,N_29454);
nand UO_640 (O_640,N_28916,N_29013);
nand UO_641 (O_641,N_29247,N_29885);
nand UO_642 (O_642,N_29428,N_29273);
nor UO_643 (O_643,N_29351,N_29093);
nand UO_644 (O_644,N_29025,N_29911);
nor UO_645 (O_645,N_28907,N_29216);
nor UO_646 (O_646,N_28888,N_29808);
nand UO_647 (O_647,N_29038,N_29456);
nand UO_648 (O_648,N_29944,N_29463);
and UO_649 (O_649,N_28947,N_29928);
nand UO_650 (O_650,N_28706,N_29978);
and UO_651 (O_651,N_29376,N_29974);
or UO_652 (O_652,N_29356,N_28617);
xor UO_653 (O_653,N_29422,N_29623);
nor UO_654 (O_654,N_28594,N_29948);
or UO_655 (O_655,N_29112,N_29720);
or UO_656 (O_656,N_28749,N_28509);
and UO_657 (O_657,N_28695,N_29309);
and UO_658 (O_658,N_29154,N_29823);
or UO_659 (O_659,N_29615,N_29695);
and UO_660 (O_660,N_29983,N_29705);
or UO_661 (O_661,N_28542,N_29385);
nor UO_662 (O_662,N_29803,N_29592);
and UO_663 (O_663,N_29500,N_29881);
xor UO_664 (O_664,N_29582,N_29277);
and UO_665 (O_665,N_29649,N_29382);
nand UO_666 (O_666,N_29867,N_29437);
nor UO_667 (O_667,N_29291,N_28647);
and UO_668 (O_668,N_29739,N_29818);
nor UO_669 (O_669,N_29048,N_28894);
or UO_670 (O_670,N_28824,N_29181);
or UO_671 (O_671,N_29157,N_28944);
nor UO_672 (O_672,N_29426,N_28805);
or UO_673 (O_673,N_29882,N_29207);
xor UO_674 (O_674,N_29884,N_29191);
or UO_675 (O_675,N_29963,N_29525);
or UO_676 (O_676,N_29324,N_29555);
or UO_677 (O_677,N_29910,N_29305);
and UO_678 (O_678,N_29843,N_28777);
xnor UO_679 (O_679,N_28962,N_29680);
or UO_680 (O_680,N_28835,N_28883);
nand UO_681 (O_681,N_29168,N_29521);
and UO_682 (O_682,N_28967,N_29488);
xnor UO_683 (O_683,N_29095,N_29493);
or UO_684 (O_684,N_28788,N_29073);
and UO_685 (O_685,N_29223,N_29359);
or UO_686 (O_686,N_29172,N_28730);
xor UO_687 (O_687,N_29081,N_29907);
nor UO_688 (O_688,N_29647,N_29177);
and UO_689 (O_689,N_29047,N_29622);
nand UO_690 (O_690,N_29204,N_28765);
nor UO_691 (O_691,N_29835,N_28637);
nand UO_692 (O_692,N_28756,N_28623);
nand UO_693 (O_693,N_29170,N_28965);
nand UO_694 (O_694,N_29075,N_29711);
nor UO_695 (O_695,N_28826,N_29840);
nand UO_696 (O_696,N_29318,N_29336);
or UO_697 (O_697,N_28592,N_29915);
xnor UO_698 (O_698,N_28857,N_29436);
nand UO_699 (O_699,N_29039,N_28651);
xnor UO_700 (O_700,N_29184,N_28607);
nor UO_701 (O_701,N_29250,N_29825);
or UO_702 (O_702,N_29785,N_29000);
nor UO_703 (O_703,N_28561,N_29806);
or UO_704 (O_704,N_29321,N_29712);
nand UO_705 (O_705,N_29744,N_29838);
xnor UO_706 (O_706,N_28703,N_29596);
and UO_707 (O_707,N_29357,N_28628);
xnor UO_708 (O_708,N_29943,N_29327);
nand UO_709 (O_709,N_29690,N_29271);
nand UO_710 (O_710,N_29523,N_29211);
xor UO_711 (O_711,N_29798,N_29344);
and UO_712 (O_712,N_29658,N_29782);
and UO_713 (O_713,N_28716,N_28754);
nand UO_714 (O_714,N_29438,N_29003);
or UO_715 (O_715,N_29161,N_28804);
nand UO_716 (O_716,N_28946,N_29099);
and UO_717 (O_717,N_29906,N_29314);
xnor UO_718 (O_718,N_29857,N_28719);
or UO_719 (O_719,N_28677,N_28641);
or UO_720 (O_720,N_28554,N_28728);
and UO_721 (O_721,N_29286,N_29576);
or UO_722 (O_722,N_28872,N_29476);
or UO_723 (O_723,N_28747,N_29260);
nand UO_724 (O_724,N_29462,N_28782);
nor UO_725 (O_725,N_28975,N_29722);
xnor UO_726 (O_726,N_29480,N_28798);
xor UO_727 (O_727,N_29574,N_29851);
xor UO_728 (O_728,N_29246,N_29864);
or UO_729 (O_729,N_29638,N_29558);
and UO_730 (O_730,N_29749,N_29933);
nand UO_731 (O_731,N_29996,N_28737);
xor UO_732 (O_732,N_29645,N_29338);
and UO_733 (O_733,N_29078,N_29126);
nand UO_734 (O_734,N_29245,N_28559);
nand UO_735 (O_735,N_29659,N_29724);
xnor UO_736 (O_736,N_29062,N_28976);
nor UO_737 (O_737,N_29103,N_28642);
and UO_738 (O_738,N_28718,N_29496);
xnor UO_739 (O_739,N_29167,N_29678);
nor UO_740 (O_740,N_29122,N_29225);
and UO_741 (O_741,N_29549,N_29391);
or UO_742 (O_742,N_29015,N_29970);
and UO_743 (O_743,N_28744,N_29830);
and UO_744 (O_744,N_28887,N_29946);
nor UO_745 (O_745,N_29342,N_29988);
xor UO_746 (O_746,N_29653,N_29784);
xor UO_747 (O_747,N_29727,N_29478);
and UO_748 (O_748,N_29990,N_28584);
and UO_749 (O_749,N_29847,N_29846);
and UO_750 (O_750,N_29802,N_29852);
nor UO_751 (O_751,N_28597,N_29674);
xor UO_752 (O_752,N_29952,N_28860);
nor UO_753 (O_753,N_28648,N_29585);
or UO_754 (O_754,N_29262,N_28712);
xor UO_755 (O_755,N_28547,N_29113);
or UO_756 (O_756,N_29196,N_29675);
nor UO_757 (O_757,N_29947,N_29577);
nor UO_758 (O_758,N_28611,N_28727);
or UO_759 (O_759,N_29618,N_28719);
nor UO_760 (O_760,N_28971,N_28505);
or UO_761 (O_761,N_29797,N_28839);
xnor UO_762 (O_762,N_29556,N_28735);
or UO_763 (O_763,N_29062,N_28836);
and UO_764 (O_764,N_29248,N_29257);
xnor UO_765 (O_765,N_28937,N_29729);
and UO_766 (O_766,N_28754,N_29260);
xor UO_767 (O_767,N_28715,N_29237);
and UO_768 (O_768,N_29123,N_28500);
or UO_769 (O_769,N_29650,N_28740);
nand UO_770 (O_770,N_29791,N_28937);
nand UO_771 (O_771,N_28921,N_29438);
and UO_772 (O_772,N_29417,N_29754);
nor UO_773 (O_773,N_29534,N_29606);
or UO_774 (O_774,N_29312,N_29897);
nor UO_775 (O_775,N_29023,N_29661);
or UO_776 (O_776,N_29520,N_29695);
nor UO_777 (O_777,N_28939,N_28635);
xor UO_778 (O_778,N_29808,N_28985);
nor UO_779 (O_779,N_29820,N_28572);
or UO_780 (O_780,N_29310,N_28812);
nand UO_781 (O_781,N_29233,N_29872);
nand UO_782 (O_782,N_29009,N_28736);
and UO_783 (O_783,N_28664,N_29273);
or UO_784 (O_784,N_29268,N_29256);
or UO_785 (O_785,N_29459,N_29903);
nand UO_786 (O_786,N_29429,N_28849);
xor UO_787 (O_787,N_29020,N_29768);
and UO_788 (O_788,N_29820,N_29978);
and UO_789 (O_789,N_29273,N_29805);
and UO_790 (O_790,N_28709,N_29897);
nand UO_791 (O_791,N_28779,N_29272);
xor UO_792 (O_792,N_29103,N_29329);
nand UO_793 (O_793,N_28575,N_29803);
or UO_794 (O_794,N_29657,N_28937);
xor UO_795 (O_795,N_28756,N_29673);
xnor UO_796 (O_796,N_29700,N_29409);
xnor UO_797 (O_797,N_29579,N_29192);
xnor UO_798 (O_798,N_29094,N_29546);
nor UO_799 (O_799,N_29036,N_29506);
nand UO_800 (O_800,N_29978,N_28665);
xor UO_801 (O_801,N_29540,N_28749);
xnor UO_802 (O_802,N_29281,N_28779);
nor UO_803 (O_803,N_28708,N_29304);
nand UO_804 (O_804,N_29497,N_28907);
or UO_805 (O_805,N_29691,N_29185);
and UO_806 (O_806,N_28960,N_28565);
nor UO_807 (O_807,N_29272,N_29152);
xor UO_808 (O_808,N_29351,N_29857);
or UO_809 (O_809,N_28657,N_29809);
or UO_810 (O_810,N_29005,N_29638);
or UO_811 (O_811,N_28646,N_28928);
or UO_812 (O_812,N_28682,N_29382);
nor UO_813 (O_813,N_28782,N_28583);
or UO_814 (O_814,N_29453,N_29206);
nand UO_815 (O_815,N_29603,N_28578);
nor UO_816 (O_816,N_29206,N_29128);
nand UO_817 (O_817,N_28587,N_29579);
xor UO_818 (O_818,N_29206,N_29614);
nand UO_819 (O_819,N_29611,N_28946);
nand UO_820 (O_820,N_29841,N_29560);
nor UO_821 (O_821,N_28608,N_29025);
nand UO_822 (O_822,N_29400,N_28621);
xnor UO_823 (O_823,N_29076,N_29347);
nand UO_824 (O_824,N_28819,N_29661);
and UO_825 (O_825,N_29227,N_28944);
xor UO_826 (O_826,N_28628,N_29618);
nand UO_827 (O_827,N_29004,N_28640);
nor UO_828 (O_828,N_29889,N_29198);
or UO_829 (O_829,N_29260,N_29794);
xor UO_830 (O_830,N_28798,N_28641);
xnor UO_831 (O_831,N_29361,N_29529);
nand UO_832 (O_832,N_29337,N_29796);
or UO_833 (O_833,N_28595,N_28659);
or UO_834 (O_834,N_28658,N_29033);
nor UO_835 (O_835,N_28855,N_29001);
or UO_836 (O_836,N_29468,N_29811);
and UO_837 (O_837,N_28557,N_29014);
nand UO_838 (O_838,N_29699,N_28836);
and UO_839 (O_839,N_29547,N_29293);
or UO_840 (O_840,N_29922,N_28750);
nor UO_841 (O_841,N_29065,N_28951);
or UO_842 (O_842,N_29115,N_29226);
or UO_843 (O_843,N_29195,N_29175);
and UO_844 (O_844,N_28980,N_28606);
and UO_845 (O_845,N_28653,N_28536);
and UO_846 (O_846,N_28889,N_29093);
nor UO_847 (O_847,N_28744,N_29082);
and UO_848 (O_848,N_29480,N_29481);
or UO_849 (O_849,N_29432,N_29159);
or UO_850 (O_850,N_29561,N_29632);
nor UO_851 (O_851,N_29013,N_29037);
nand UO_852 (O_852,N_29769,N_29173);
or UO_853 (O_853,N_29698,N_28891);
nor UO_854 (O_854,N_29006,N_29651);
or UO_855 (O_855,N_29312,N_28953);
or UO_856 (O_856,N_28653,N_29272);
nand UO_857 (O_857,N_29194,N_29580);
and UO_858 (O_858,N_29213,N_29365);
nand UO_859 (O_859,N_29967,N_28642);
and UO_860 (O_860,N_29872,N_29881);
nor UO_861 (O_861,N_29154,N_29196);
nor UO_862 (O_862,N_28649,N_29391);
xor UO_863 (O_863,N_29416,N_29968);
nor UO_864 (O_864,N_29752,N_28517);
and UO_865 (O_865,N_29457,N_29301);
nand UO_866 (O_866,N_29128,N_28579);
or UO_867 (O_867,N_29670,N_28752);
and UO_868 (O_868,N_29763,N_29121);
nand UO_869 (O_869,N_28711,N_28722);
nand UO_870 (O_870,N_29923,N_28629);
or UO_871 (O_871,N_29648,N_29887);
nor UO_872 (O_872,N_28578,N_28970);
xnor UO_873 (O_873,N_29360,N_28720);
nand UO_874 (O_874,N_29067,N_29178);
and UO_875 (O_875,N_29824,N_29505);
nand UO_876 (O_876,N_28927,N_29854);
and UO_877 (O_877,N_29486,N_28685);
xor UO_878 (O_878,N_29959,N_28610);
and UO_879 (O_879,N_29014,N_28591);
xor UO_880 (O_880,N_28951,N_29823);
nor UO_881 (O_881,N_28732,N_29392);
nand UO_882 (O_882,N_29026,N_29987);
nor UO_883 (O_883,N_29955,N_29117);
nor UO_884 (O_884,N_28587,N_29790);
nand UO_885 (O_885,N_29835,N_28519);
or UO_886 (O_886,N_28692,N_29772);
or UO_887 (O_887,N_28934,N_29580);
nor UO_888 (O_888,N_29084,N_28881);
nor UO_889 (O_889,N_29018,N_28928);
xor UO_890 (O_890,N_28521,N_29723);
nor UO_891 (O_891,N_29711,N_29727);
and UO_892 (O_892,N_29685,N_28542);
or UO_893 (O_893,N_29613,N_29088);
xor UO_894 (O_894,N_29505,N_28910);
nor UO_895 (O_895,N_29719,N_29687);
and UO_896 (O_896,N_28890,N_28796);
xor UO_897 (O_897,N_28588,N_29919);
nand UO_898 (O_898,N_29699,N_29555);
nand UO_899 (O_899,N_29181,N_29945);
nor UO_900 (O_900,N_28697,N_29888);
nor UO_901 (O_901,N_29158,N_29613);
nand UO_902 (O_902,N_29988,N_29105);
xnor UO_903 (O_903,N_29106,N_28515);
nor UO_904 (O_904,N_29521,N_29811);
xnor UO_905 (O_905,N_29009,N_28685);
xnor UO_906 (O_906,N_29969,N_28596);
nor UO_907 (O_907,N_29085,N_28631);
and UO_908 (O_908,N_28894,N_29288);
nand UO_909 (O_909,N_29721,N_28535);
xor UO_910 (O_910,N_29423,N_28783);
nand UO_911 (O_911,N_29388,N_29901);
or UO_912 (O_912,N_28665,N_29958);
or UO_913 (O_913,N_29030,N_28941);
and UO_914 (O_914,N_29948,N_29392);
and UO_915 (O_915,N_29211,N_29673);
xnor UO_916 (O_916,N_29933,N_29889);
or UO_917 (O_917,N_29837,N_28546);
and UO_918 (O_918,N_29755,N_29248);
xor UO_919 (O_919,N_29816,N_29576);
nand UO_920 (O_920,N_28662,N_29747);
and UO_921 (O_921,N_29917,N_29194);
nor UO_922 (O_922,N_29206,N_29138);
xor UO_923 (O_923,N_29641,N_29863);
xnor UO_924 (O_924,N_28686,N_29105);
nand UO_925 (O_925,N_29947,N_29919);
or UO_926 (O_926,N_28768,N_29969);
and UO_927 (O_927,N_29669,N_29395);
or UO_928 (O_928,N_28590,N_29623);
xor UO_929 (O_929,N_29894,N_29978);
or UO_930 (O_930,N_29531,N_29957);
nand UO_931 (O_931,N_29589,N_29539);
nand UO_932 (O_932,N_29310,N_29309);
xnor UO_933 (O_933,N_29959,N_28968);
or UO_934 (O_934,N_28640,N_29735);
or UO_935 (O_935,N_28935,N_29098);
nor UO_936 (O_936,N_28594,N_29035);
nor UO_937 (O_937,N_28633,N_29442);
or UO_938 (O_938,N_28708,N_29053);
nand UO_939 (O_939,N_29760,N_28798);
xnor UO_940 (O_940,N_28745,N_29559);
or UO_941 (O_941,N_28675,N_28798);
or UO_942 (O_942,N_29862,N_29834);
or UO_943 (O_943,N_29260,N_28920);
nor UO_944 (O_944,N_29051,N_29631);
and UO_945 (O_945,N_29094,N_29436);
nand UO_946 (O_946,N_29798,N_28933);
xnor UO_947 (O_947,N_29637,N_29152);
xor UO_948 (O_948,N_29952,N_28572);
nor UO_949 (O_949,N_29369,N_29575);
and UO_950 (O_950,N_28771,N_29318);
or UO_951 (O_951,N_28579,N_29389);
xor UO_952 (O_952,N_29272,N_29579);
or UO_953 (O_953,N_29434,N_29452);
and UO_954 (O_954,N_28617,N_29947);
nor UO_955 (O_955,N_28763,N_29539);
or UO_956 (O_956,N_28976,N_29513);
and UO_957 (O_957,N_29261,N_29441);
xnor UO_958 (O_958,N_29618,N_29705);
nand UO_959 (O_959,N_29524,N_28871);
xor UO_960 (O_960,N_28717,N_28926);
xor UO_961 (O_961,N_29993,N_29522);
nor UO_962 (O_962,N_29355,N_28995);
xnor UO_963 (O_963,N_29544,N_29670);
nand UO_964 (O_964,N_29150,N_29981);
nand UO_965 (O_965,N_29246,N_29908);
xor UO_966 (O_966,N_29966,N_28849);
or UO_967 (O_967,N_28901,N_28570);
or UO_968 (O_968,N_29015,N_28766);
and UO_969 (O_969,N_29718,N_29790);
and UO_970 (O_970,N_28506,N_28929);
nor UO_971 (O_971,N_29795,N_28822);
xor UO_972 (O_972,N_29052,N_29668);
or UO_973 (O_973,N_28574,N_29377);
nor UO_974 (O_974,N_29800,N_29963);
nand UO_975 (O_975,N_29984,N_29895);
nor UO_976 (O_976,N_28624,N_29635);
xnor UO_977 (O_977,N_29486,N_29503);
nand UO_978 (O_978,N_29292,N_29206);
or UO_979 (O_979,N_28952,N_29459);
and UO_980 (O_980,N_29769,N_29213);
xnor UO_981 (O_981,N_29625,N_29820);
or UO_982 (O_982,N_28864,N_29914);
xnor UO_983 (O_983,N_29177,N_29315);
xnor UO_984 (O_984,N_29992,N_28686);
or UO_985 (O_985,N_29500,N_29628);
nand UO_986 (O_986,N_29170,N_28650);
and UO_987 (O_987,N_29925,N_29373);
xor UO_988 (O_988,N_28898,N_29966);
nand UO_989 (O_989,N_29822,N_28983);
nor UO_990 (O_990,N_29392,N_29146);
xnor UO_991 (O_991,N_29728,N_29827);
xnor UO_992 (O_992,N_29674,N_29594);
xnor UO_993 (O_993,N_29094,N_29122);
nand UO_994 (O_994,N_29748,N_29784);
nand UO_995 (O_995,N_29039,N_28671);
xnor UO_996 (O_996,N_29861,N_29568);
nand UO_997 (O_997,N_29845,N_28906);
xnor UO_998 (O_998,N_29529,N_29585);
nand UO_999 (O_999,N_29438,N_29425);
xor UO_1000 (O_1000,N_29584,N_29924);
or UO_1001 (O_1001,N_28609,N_29502);
nor UO_1002 (O_1002,N_29762,N_29214);
or UO_1003 (O_1003,N_29813,N_29108);
xor UO_1004 (O_1004,N_29445,N_28532);
nor UO_1005 (O_1005,N_28997,N_28826);
xor UO_1006 (O_1006,N_28996,N_28559);
or UO_1007 (O_1007,N_28823,N_29061);
or UO_1008 (O_1008,N_29185,N_29521);
and UO_1009 (O_1009,N_29545,N_28942);
or UO_1010 (O_1010,N_28533,N_29025);
xnor UO_1011 (O_1011,N_29925,N_28669);
nor UO_1012 (O_1012,N_28783,N_28564);
nand UO_1013 (O_1013,N_28759,N_28751);
or UO_1014 (O_1014,N_28651,N_28721);
and UO_1015 (O_1015,N_29174,N_29593);
nor UO_1016 (O_1016,N_29925,N_29883);
xor UO_1017 (O_1017,N_29778,N_28581);
and UO_1018 (O_1018,N_29209,N_29480);
nor UO_1019 (O_1019,N_29635,N_28708);
nand UO_1020 (O_1020,N_29333,N_29079);
nand UO_1021 (O_1021,N_29252,N_29917);
or UO_1022 (O_1022,N_29700,N_28663);
and UO_1023 (O_1023,N_29932,N_29230);
and UO_1024 (O_1024,N_29160,N_28766);
nand UO_1025 (O_1025,N_29276,N_28749);
nor UO_1026 (O_1026,N_29815,N_28713);
xor UO_1027 (O_1027,N_28621,N_28951);
and UO_1028 (O_1028,N_29886,N_28782);
and UO_1029 (O_1029,N_28855,N_29995);
nand UO_1030 (O_1030,N_28512,N_29953);
xnor UO_1031 (O_1031,N_29293,N_28516);
or UO_1032 (O_1032,N_28646,N_28946);
xor UO_1033 (O_1033,N_28895,N_28744);
or UO_1034 (O_1034,N_29971,N_29178);
nor UO_1035 (O_1035,N_28743,N_28767);
or UO_1036 (O_1036,N_28893,N_28664);
or UO_1037 (O_1037,N_28816,N_28534);
nand UO_1038 (O_1038,N_28914,N_29829);
xor UO_1039 (O_1039,N_28776,N_29861);
xnor UO_1040 (O_1040,N_28680,N_29325);
nor UO_1041 (O_1041,N_28785,N_29081);
xnor UO_1042 (O_1042,N_29989,N_29686);
or UO_1043 (O_1043,N_29881,N_29372);
nand UO_1044 (O_1044,N_29833,N_28641);
nor UO_1045 (O_1045,N_29301,N_29293);
or UO_1046 (O_1046,N_29058,N_29291);
and UO_1047 (O_1047,N_28947,N_29880);
nand UO_1048 (O_1048,N_29255,N_29367);
or UO_1049 (O_1049,N_29909,N_29338);
xor UO_1050 (O_1050,N_29854,N_29997);
nand UO_1051 (O_1051,N_29328,N_29814);
xor UO_1052 (O_1052,N_28830,N_29269);
and UO_1053 (O_1053,N_28880,N_29893);
and UO_1054 (O_1054,N_29503,N_28540);
xor UO_1055 (O_1055,N_29064,N_29774);
nor UO_1056 (O_1056,N_29528,N_28654);
nand UO_1057 (O_1057,N_29419,N_29834);
and UO_1058 (O_1058,N_29767,N_28549);
nand UO_1059 (O_1059,N_29709,N_28713);
nand UO_1060 (O_1060,N_29662,N_29086);
and UO_1061 (O_1061,N_29457,N_29545);
nor UO_1062 (O_1062,N_29563,N_29730);
and UO_1063 (O_1063,N_29657,N_28701);
xnor UO_1064 (O_1064,N_29769,N_28625);
nand UO_1065 (O_1065,N_28895,N_28524);
and UO_1066 (O_1066,N_28613,N_29037);
and UO_1067 (O_1067,N_29171,N_28866);
nor UO_1068 (O_1068,N_28508,N_29106);
or UO_1069 (O_1069,N_29905,N_29413);
or UO_1070 (O_1070,N_28638,N_28959);
and UO_1071 (O_1071,N_29233,N_29407);
and UO_1072 (O_1072,N_29773,N_29627);
nor UO_1073 (O_1073,N_28588,N_29879);
or UO_1074 (O_1074,N_29456,N_29079);
and UO_1075 (O_1075,N_29910,N_28579);
or UO_1076 (O_1076,N_29935,N_28859);
or UO_1077 (O_1077,N_29727,N_29521);
or UO_1078 (O_1078,N_28762,N_28512);
nand UO_1079 (O_1079,N_28827,N_29586);
xor UO_1080 (O_1080,N_29732,N_29087);
or UO_1081 (O_1081,N_29660,N_29755);
nand UO_1082 (O_1082,N_29003,N_28791);
nand UO_1083 (O_1083,N_28711,N_29968);
nand UO_1084 (O_1084,N_29628,N_29134);
or UO_1085 (O_1085,N_28741,N_29301);
and UO_1086 (O_1086,N_29477,N_29196);
and UO_1087 (O_1087,N_29898,N_29015);
nand UO_1088 (O_1088,N_28769,N_29006);
xor UO_1089 (O_1089,N_29645,N_29254);
and UO_1090 (O_1090,N_29126,N_29149);
xnor UO_1091 (O_1091,N_29953,N_28851);
xor UO_1092 (O_1092,N_28607,N_29454);
nor UO_1093 (O_1093,N_28530,N_29202);
nand UO_1094 (O_1094,N_29097,N_29824);
or UO_1095 (O_1095,N_29609,N_29174);
or UO_1096 (O_1096,N_29326,N_28852);
xnor UO_1097 (O_1097,N_29696,N_29402);
and UO_1098 (O_1098,N_28551,N_28901);
nor UO_1099 (O_1099,N_29082,N_29349);
or UO_1100 (O_1100,N_28822,N_29176);
and UO_1101 (O_1101,N_29965,N_29958);
and UO_1102 (O_1102,N_29433,N_29625);
and UO_1103 (O_1103,N_29645,N_28706);
and UO_1104 (O_1104,N_28903,N_29923);
xor UO_1105 (O_1105,N_28657,N_29657);
or UO_1106 (O_1106,N_29958,N_29756);
nor UO_1107 (O_1107,N_28726,N_29407);
nor UO_1108 (O_1108,N_29739,N_29284);
or UO_1109 (O_1109,N_28660,N_28518);
and UO_1110 (O_1110,N_29510,N_29907);
xnor UO_1111 (O_1111,N_29473,N_29619);
xnor UO_1112 (O_1112,N_28785,N_29157);
nor UO_1113 (O_1113,N_28723,N_29702);
xnor UO_1114 (O_1114,N_29506,N_29633);
and UO_1115 (O_1115,N_29598,N_29924);
or UO_1116 (O_1116,N_29682,N_28826);
nor UO_1117 (O_1117,N_29143,N_29455);
and UO_1118 (O_1118,N_29370,N_29055);
nor UO_1119 (O_1119,N_29719,N_29991);
or UO_1120 (O_1120,N_29996,N_28572);
nand UO_1121 (O_1121,N_29091,N_29099);
nor UO_1122 (O_1122,N_29945,N_29094);
nor UO_1123 (O_1123,N_28681,N_29199);
nand UO_1124 (O_1124,N_28582,N_29122);
and UO_1125 (O_1125,N_28952,N_29758);
xnor UO_1126 (O_1126,N_29183,N_29382);
and UO_1127 (O_1127,N_29644,N_28587);
nor UO_1128 (O_1128,N_28896,N_28713);
nand UO_1129 (O_1129,N_29446,N_28755);
nand UO_1130 (O_1130,N_29978,N_29592);
xor UO_1131 (O_1131,N_29118,N_29210);
nand UO_1132 (O_1132,N_29151,N_28500);
xor UO_1133 (O_1133,N_29993,N_28655);
nand UO_1134 (O_1134,N_29009,N_28656);
nor UO_1135 (O_1135,N_29785,N_29399);
and UO_1136 (O_1136,N_29616,N_29880);
xnor UO_1137 (O_1137,N_28832,N_28762);
and UO_1138 (O_1138,N_29218,N_28669);
nand UO_1139 (O_1139,N_29420,N_29025);
and UO_1140 (O_1140,N_28753,N_29413);
xnor UO_1141 (O_1141,N_28837,N_29930);
nor UO_1142 (O_1142,N_29298,N_29775);
nor UO_1143 (O_1143,N_29301,N_29879);
or UO_1144 (O_1144,N_29958,N_29952);
and UO_1145 (O_1145,N_28532,N_28751);
or UO_1146 (O_1146,N_29244,N_29404);
nor UO_1147 (O_1147,N_28651,N_29285);
or UO_1148 (O_1148,N_29712,N_29694);
nor UO_1149 (O_1149,N_29146,N_29835);
and UO_1150 (O_1150,N_28723,N_29413);
xnor UO_1151 (O_1151,N_29199,N_28579);
and UO_1152 (O_1152,N_28907,N_28889);
xor UO_1153 (O_1153,N_28902,N_29355);
nor UO_1154 (O_1154,N_29120,N_28550);
nor UO_1155 (O_1155,N_28987,N_28830);
xnor UO_1156 (O_1156,N_29039,N_28528);
nor UO_1157 (O_1157,N_28719,N_29919);
nand UO_1158 (O_1158,N_29112,N_29009);
and UO_1159 (O_1159,N_29566,N_29987);
nor UO_1160 (O_1160,N_28706,N_29310);
nand UO_1161 (O_1161,N_28902,N_29443);
xnor UO_1162 (O_1162,N_28845,N_29617);
and UO_1163 (O_1163,N_28651,N_28504);
and UO_1164 (O_1164,N_29442,N_29499);
nor UO_1165 (O_1165,N_29197,N_29564);
xnor UO_1166 (O_1166,N_29587,N_29385);
and UO_1167 (O_1167,N_29194,N_29695);
xnor UO_1168 (O_1168,N_29917,N_28735);
nand UO_1169 (O_1169,N_29237,N_29493);
and UO_1170 (O_1170,N_29823,N_29543);
or UO_1171 (O_1171,N_29643,N_28920);
and UO_1172 (O_1172,N_28833,N_29053);
or UO_1173 (O_1173,N_29669,N_29796);
nor UO_1174 (O_1174,N_29996,N_28754);
nor UO_1175 (O_1175,N_28650,N_29088);
nor UO_1176 (O_1176,N_29667,N_29095);
xor UO_1177 (O_1177,N_29786,N_29491);
nand UO_1178 (O_1178,N_28565,N_29016);
or UO_1179 (O_1179,N_29823,N_29015);
and UO_1180 (O_1180,N_29703,N_29406);
and UO_1181 (O_1181,N_29937,N_29291);
nand UO_1182 (O_1182,N_28571,N_29208);
nor UO_1183 (O_1183,N_29428,N_29452);
or UO_1184 (O_1184,N_29893,N_29847);
nand UO_1185 (O_1185,N_29127,N_29920);
and UO_1186 (O_1186,N_28896,N_29368);
nor UO_1187 (O_1187,N_29999,N_29222);
and UO_1188 (O_1188,N_29193,N_29870);
nand UO_1189 (O_1189,N_28695,N_29281);
nand UO_1190 (O_1190,N_29871,N_29207);
nand UO_1191 (O_1191,N_29397,N_29506);
xnor UO_1192 (O_1192,N_29131,N_29944);
nand UO_1193 (O_1193,N_29246,N_29642);
nand UO_1194 (O_1194,N_28956,N_29070);
nand UO_1195 (O_1195,N_28765,N_29398);
nor UO_1196 (O_1196,N_29407,N_29369);
nand UO_1197 (O_1197,N_29234,N_29852);
xor UO_1198 (O_1198,N_28623,N_28511);
nor UO_1199 (O_1199,N_29422,N_29848);
nand UO_1200 (O_1200,N_29462,N_29688);
xor UO_1201 (O_1201,N_29031,N_29606);
xnor UO_1202 (O_1202,N_29692,N_29941);
xnor UO_1203 (O_1203,N_29894,N_28802);
xor UO_1204 (O_1204,N_29222,N_29233);
or UO_1205 (O_1205,N_28777,N_29447);
nor UO_1206 (O_1206,N_28744,N_28514);
and UO_1207 (O_1207,N_29488,N_29423);
nand UO_1208 (O_1208,N_29500,N_29233);
nand UO_1209 (O_1209,N_29216,N_29348);
and UO_1210 (O_1210,N_28523,N_29859);
xor UO_1211 (O_1211,N_28955,N_29330);
and UO_1212 (O_1212,N_29107,N_28853);
nor UO_1213 (O_1213,N_29059,N_29027);
nand UO_1214 (O_1214,N_29154,N_28827);
nand UO_1215 (O_1215,N_28853,N_29085);
or UO_1216 (O_1216,N_29236,N_28970);
nor UO_1217 (O_1217,N_29956,N_28577);
or UO_1218 (O_1218,N_29271,N_29783);
or UO_1219 (O_1219,N_28588,N_29645);
nor UO_1220 (O_1220,N_29339,N_29840);
xor UO_1221 (O_1221,N_28589,N_28652);
nor UO_1222 (O_1222,N_29661,N_29740);
nor UO_1223 (O_1223,N_28596,N_29006);
xnor UO_1224 (O_1224,N_29976,N_28565);
nor UO_1225 (O_1225,N_28837,N_29274);
or UO_1226 (O_1226,N_28925,N_28610);
xor UO_1227 (O_1227,N_29589,N_29677);
and UO_1228 (O_1228,N_29252,N_29396);
nand UO_1229 (O_1229,N_28636,N_29073);
nor UO_1230 (O_1230,N_29514,N_28629);
and UO_1231 (O_1231,N_29176,N_29109);
or UO_1232 (O_1232,N_29604,N_29529);
nor UO_1233 (O_1233,N_29580,N_28704);
and UO_1234 (O_1234,N_28675,N_29553);
and UO_1235 (O_1235,N_29719,N_29256);
xnor UO_1236 (O_1236,N_29899,N_29063);
and UO_1237 (O_1237,N_29950,N_28500);
nor UO_1238 (O_1238,N_29531,N_28551);
and UO_1239 (O_1239,N_29836,N_29991);
and UO_1240 (O_1240,N_28605,N_28542);
xnor UO_1241 (O_1241,N_29653,N_29726);
nand UO_1242 (O_1242,N_29705,N_28608);
nand UO_1243 (O_1243,N_28585,N_28844);
nor UO_1244 (O_1244,N_29190,N_28682);
or UO_1245 (O_1245,N_29068,N_28627);
and UO_1246 (O_1246,N_29651,N_29344);
xor UO_1247 (O_1247,N_29714,N_29306);
and UO_1248 (O_1248,N_29901,N_28956);
or UO_1249 (O_1249,N_28551,N_29902);
xnor UO_1250 (O_1250,N_28612,N_29442);
nor UO_1251 (O_1251,N_28679,N_29740);
or UO_1252 (O_1252,N_28702,N_29588);
nor UO_1253 (O_1253,N_29727,N_29286);
nand UO_1254 (O_1254,N_29661,N_29273);
or UO_1255 (O_1255,N_28925,N_29038);
xnor UO_1256 (O_1256,N_29923,N_29065);
and UO_1257 (O_1257,N_29511,N_28727);
or UO_1258 (O_1258,N_29138,N_28655);
and UO_1259 (O_1259,N_28955,N_29065);
xnor UO_1260 (O_1260,N_28937,N_29738);
or UO_1261 (O_1261,N_28746,N_29614);
or UO_1262 (O_1262,N_29669,N_29474);
nand UO_1263 (O_1263,N_29998,N_28711);
nor UO_1264 (O_1264,N_29824,N_29455);
and UO_1265 (O_1265,N_29228,N_29526);
nand UO_1266 (O_1266,N_29671,N_29672);
nand UO_1267 (O_1267,N_29057,N_29110);
and UO_1268 (O_1268,N_28776,N_29656);
and UO_1269 (O_1269,N_29455,N_29919);
nand UO_1270 (O_1270,N_29755,N_29849);
nor UO_1271 (O_1271,N_29820,N_28582);
or UO_1272 (O_1272,N_28862,N_28642);
or UO_1273 (O_1273,N_29710,N_29959);
nand UO_1274 (O_1274,N_28915,N_29574);
nor UO_1275 (O_1275,N_29933,N_28898);
nand UO_1276 (O_1276,N_29195,N_28822);
or UO_1277 (O_1277,N_29802,N_29422);
nand UO_1278 (O_1278,N_28509,N_29024);
xnor UO_1279 (O_1279,N_28922,N_28703);
nor UO_1280 (O_1280,N_29546,N_28637);
nand UO_1281 (O_1281,N_28963,N_29503);
nor UO_1282 (O_1282,N_29952,N_29230);
and UO_1283 (O_1283,N_29971,N_28537);
or UO_1284 (O_1284,N_29863,N_29279);
xnor UO_1285 (O_1285,N_28560,N_28619);
or UO_1286 (O_1286,N_29052,N_29191);
xor UO_1287 (O_1287,N_29891,N_29475);
and UO_1288 (O_1288,N_29423,N_29394);
xnor UO_1289 (O_1289,N_29836,N_28859);
or UO_1290 (O_1290,N_29965,N_28517);
nand UO_1291 (O_1291,N_29568,N_29162);
xor UO_1292 (O_1292,N_29114,N_28604);
or UO_1293 (O_1293,N_29261,N_29942);
nand UO_1294 (O_1294,N_29575,N_29872);
xnor UO_1295 (O_1295,N_29781,N_29715);
and UO_1296 (O_1296,N_28926,N_29055);
or UO_1297 (O_1297,N_29763,N_28984);
xnor UO_1298 (O_1298,N_29076,N_29723);
xnor UO_1299 (O_1299,N_28801,N_29563);
nor UO_1300 (O_1300,N_29963,N_29237);
nor UO_1301 (O_1301,N_29944,N_28558);
nor UO_1302 (O_1302,N_29832,N_29434);
xor UO_1303 (O_1303,N_29105,N_29486);
nor UO_1304 (O_1304,N_29662,N_29312);
xor UO_1305 (O_1305,N_28623,N_28523);
nand UO_1306 (O_1306,N_28924,N_28839);
and UO_1307 (O_1307,N_29425,N_29348);
and UO_1308 (O_1308,N_29706,N_29596);
and UO_1309 (O_1309,N_29099,N_29371);
and UO_1310 (O_1310,N_29921,N_29172);
or UO_1311 (O_1311,N_29941,N_28753);
nand UO_1312 (O_1312,N_29849,N_29072);
or UO_1313 (O_1313,N_28755,N_29247);
or UO_1314 (O_1314,N_29597,N_28811);
and UO_1315 (O_1315,N_29023,N_29387);
nor UO_1316 (O_1316,N_29105,N_29861);
and UO_1317 (O_1317,N_29167,N_28889);
or UO_1318 (O_1318,N_29881,N_28600);
nand UO_1319 (O_1319,N_29100,N_28676);
or UO_1320 (O_1320,N_29656,N_29425);
nor UO_1321 (O_1321,N_29241,N_29833);
nand UO_1322 (O_1322,N_28931,N_29847);
nand UO_1323 (O_1323,N_29167,N_29410);
nand UO_1324 (O_1324,N_29506,N_29289);
and UO_1325 (O_1325,N_29727,N_29264);
nand UO_1326 (O_1326,N_28838,N_28713);
or UO_1327 (O_1327,N_29854,N_29794);
nand UO_1328 (O_1328,N_28973,N_28640);
and UO_1329 (O_1329,N_28911,N_29245);
or UO_1330 (O_1330,N_29825,N_28663);
and UO_1331 (O_1331,N_28708,N_29548);
or UO_1332 (O_1332,N_29446,N_29220);
and UO_1333 (O_1333,N_28944,N_29706);
xor UO_1334 (O_1334,N_29845,N_28758);
nand UO_1335 (O_1335,N_28697,N_29034);
and UO_1336 (O_1336,N_28785,N_29393);
nor UO_1337 (O_1337,N_29261,N_28619);
or UO_1338 (O_1338,N_29216,N_29025);
xor UO_1339 (O_1339,N_28866,N_28681);
nor UO_1340 (O_1340,N_29523,N_29757);
nand UO_1341 (O_1341,N_29727,N_29664);
nand UO_1342 (O_1342,N_29602,N_28997);
nor UO_1343 (O_1343,N_29246,N_29654);
nor UO_1344 (O_1344,N_28510,N_28715);
or UO_1345 (O_1345,N_28845,N_29611);
or UO_1346 (O_1346,N_28832,N_28848);
and UO_1347 (O_1347,N_29421,N_29144);
xnor UO_1348 (O_1348,N_29911,N_28729);
or UO_1349 (O_1349,N_28548,N_28925);
or UO_1350 (O_1350,N_28615,N_28884);
or UO_1351 (O_1351,N_28817,N_29487);
and UO_1352 (O_1352,N_28982,N_29038);
and UO_1353 (O_1353,N_29542,N_29124);
and UO_1354 (O_1354,N_29487,N_29527);
and UO_1355 (O_1355,N_29005,N_28730);
or UO_1356 (O_1356,N_29557,N_28827);
nor UO_1357 (O_1357,N_29304,N_29459);
or UO_1358 (O_1358,N_28678,N_29906);
nor UO_1359 (O_1359,N_29924,N_29553);
nand UO_1360 (O_1360,N_29537,N_28589);
or UO_1361 (O_1361,N_29813,N_28709);
or UO_1362 (O_1362,N_29650,N_29618);
xnor UO_1363 (O_1363,N_29124,N_29223);
or UO_1364 (O_1364,N_29964,N_28974);
or UO_1365 (O_1365,N_29779,N_28753);
xor UO_1366 (O_1366,N_29728,N_28848);
or UO_1367 (O_1367,N_28943,N_28817);
nand UO_1368 (O_1368,N_29468,N_29880);
or UO_1369 (O_1369,N_29358,N_29237);
and UO_1370 (O_1370,N_29169,N_29688);
and UO_1371 (O_1371,N_29133,N_29554);
nand UO_1372 (O_1372,N_29090,N_29294);
and UO_1373 (O_1373,N_29064,N_29559);
xnor UO_1374 (O_1374,N_28966,N_28664);
nor UO_1375 (O_1375,N_28604,N_29565);
and UO_1376 (O_1376,N_28938,N_29187);
xnor UO_1377 (O_1377,N_28590,N_28944);
and UO_1378 (O_1378,N_28989,N_29040);
nor UO_1379 (O_1379,N_28544,N_29950);
nand UO_1380 (O_1380,N_29382,N_29426);
xor UO_1381 (O_1381,N_28538,N_28736);
or UO_1382 (O_1382,N_28741,N_28636);
nor UO_1383 (O_1383,N_29812,N_29366);
xor UO_1384 (O_1384,N_29459,N_29336);
and UO_1385 (O_1385,N_29496,N_28781);
and UO_1386 (O_1386,N_28696,N_28861);
or UO_1387 (O_1387,N_29111,N_29906);
nand UO_1388 (O_1388,N_29421,N_29560);
nor UO_1389 (O_1389,N_29945,N_29066);
nor UO_1390 (O_1390,N_28926,N_28959);
xnor UO_1391 (O_1391,N_28622,N_28824);
and UO_1392 (O_1392,N_28913,N_28982);
or UO_1393 (O_1393,N_29353,N_29815);
xor UO_1394 (O_1394,N_29549,N_29159);
nand UO_1395 (O_1395,N_28642,N_28841);
and UO_1396 (O_1396,N_28808,N_28540);
xor UO_1397 (O_1397,N_28993,N_29325);
xnor UO_1398 (O_1398,N_28730,N_28893);
nor UO_1399 (O_1399,N_29967,N_28897);
and UO_1400 (O_1400,N_28935,N_29109);
or UO_1401 (O_1401,N_29525,N_29691);
xor UO_1402 (O_1402,N_29645,N_28988);
xnor UO_1403 (O_1403,N_29010,N_29487);
nand UO_1404 (O_1404,N_29523,N_28873);
xnor UO_1405 (O_1405,N_29639,N_28882);
or UO_1406 (O_1406,N_29898,N_29903);
and UO_1407 (O_1407,N_28515,N_28982);
nand UO_1408 (O_1408,N_29559,N_29312);
nor UO_1409 (O_1409,N_29495,N_29713);
or UO_1410 (O_1410,N_28969,N_29383);
nor UO_1411 (O_1411,N_29529,N_29917);
xor UO_1412 (O_1412,N_29947,N_29598);
or UO_1413 (O_1413,N_29317,N_29655);
and UO_1414 (O_1414,N_28539,N_28597);
nor UO_1415 (O_1415,N_29503,N_28874);
nand UO_1416 (O_1416,N_28922,N_29591);
xor UO_1417 (O_1417,N_28684,N_29109);
nor UO_1418 (O_1418,N_28622,N_29887);
nand UO_1419 (O_1419,N_28817,N_29951);
xor UO_1420 (O_1420,N_29760,N_28720);
xnor UO_1421 (O_1421,N_29499,N_28860);
and UO_1422 (O_1422,N_29243,N_28786);
nand UO_1423 (O_1423,N_29056,N_28885);
nand UO_1424 (O_1424,N_29532,N_28768);
and UO_1425 (O_1425,N_29590,N_29084);
xor UO_1426 (O_1426,N_28660,N_28696);
and UO_1427 (O_1427,N_29632,N_29783);
nor UO_1428 (O_1428,N_28876,N_29370);
nor UO_1429 (O_1429,N_28580,N_29341);
or UO_1430 (O_1430,N_29022,N_28747);
nand UO_1431 (O_1431,N_29819,N_29599);
nand UO_1432 (O_1432,N_29505,N_29332);
nand UO_1433 (O_1433,N_29095,N_28542);
and UO_1434 (O_1434,N_29387,N_29609);
nand UO_1435 (O_1435,N_29459,N_29939);
nand UO_1436 (O_1436,N_29460,N_28509);
nor UO_1437 (O_1437,N_29595,N_29548);
or UO_1438 (O_1438,N_29509,N_28649);
and UO_1439 (O_1439,N_29248,N_28770);
nand UO_1440 (O_1440,N_29404,N_29302);
and UO_1441 (O_1441,N_29716,N_29408);
xor UO_1442 (O_1442,N_29534,N_29869);
and UO_1443 (O_1443,N_29413,N_28598);
nor UO_1444 (O_1444,N_28883,N_29497);
or UO_1445 (O_1445,N_29502,N_29311);
or UO_1446 (O_1446,N_28990,N_29571);
xor UO_1447 (O_1447,N_29563,N_29013);
nand UO_1448 (O_1448,N_29678,N_29696);
nand UO_1449 (O_1449,N_29137,N_29851);
nand UO_1450 (O_1450,N_29319,N_29337);
or UO_1451 (O_1451,N_29424,N_29903);
xnor UO_1452 (O_1452,N_29685,N_29605);
and UO_1453 (O_1453,N_29078,N_29005);
or UO_1454 (O_1454,N_29346,N_29170);
or UO_1455 (O_1455,N_28545,N_28758);
xor UO_1456 (O_1456,N_29531,N_29719);
xnor UO_1457 (O_1457,N_28843,N_29349);
and UO_1458 (O_1458,N_29268,N_28580);
and UO_1459 (O_1459,N_29978,N_29625);
nand UO_1460 (O_1460,N_29009,N_29592);
xor UO_1461 (O_1461,N_29095,N_28906);
nor UO_1462 (O_1462,N_29341,N_28787);
and UO_1463 (O_1463,N_29140,N_29292);
nand UO_1464 (O_1464,N_29844,N_28817);
or UO_1465 (O_1465,N_29009,N_28973);
and UO_1466 (O_1466,N_29926,N_29444);
nor UO_1467 (O_1467,N_28560,N_28967);
nand UO_1468 (O_1468,N_28828,N_28601);
nor UO_1469 (O_1469,N_29171,N_29861);
nand UO_1470 (O_1470,N_29147,N_29447);
xnor UO_1471 (O_1471,N_28620,N_28983);
xor UO_1472 (O_1472,N_29670,N_29366);
xnor UO_1473 (O_1473,N_29102,N_29031);
xnor UO_1474 (O_1474,N_28554,N_28598);
and UO_1475 (O_1475,N_29436,N_29069);
xnor UO_1476 (O_1476,N_29802,N_29781);
xnor UO_1477 (O_1477,N_28890,N_28671);
or UO_1478 (O_1478,N_28569,N_29674);
xnor UO_1479 (O_1479,N_29246,N_29097);
nor UO_1480 (O_1480,N_28564,N_29218);
nor UO_1481 (O_1481,N_29424,N_28864);
nand UO_1482 (O_1482,N_29064,N_29303);
and UO_1483 (O_1483,N_29522,N_29562);
and UO_1484 (O_1484,N_28772,N_29734);
or UO_1485 (O_1485,N_28916,N_28635);
nand UO_1486 (O_1486,N_28759,N_29149);
and UO_1487 (O_1487,N_29605,N_28986);
or UO_1488 (O_1488,N_28999,N_29801);
nor UO_1489 (O_1489,N_29674,N_28904);
and UO_1490 (O_1490,N_29821,N_29155);
and UO_1491 (O_1491,N_28895,N_28559);
or UO_1492 (O_1492,N_28992,N_29149);
xnor UO_1493 (O_1493,N_28926,N_29802);
or UO_1494 (O_1494,N_28676,N_29742);
or UO_1495 (O_1495,N_29115,N_28527);
nand UO_1496 (O_1496,N_29888,N_29523);
nand UO_1497 (O_1497,N_29376,N_29200);
nand UO_1498 (O_1498,N_28678,N_29956);
nor UO_1499 (O_1499,N_28952,N_29429);
nor UO_1500 (O_1500,N_28594,N_29842);
or UO_1501 (O_1501,N_29769,N_28674);
nand UO_1502 (O_1502,N_28511,N_28822);
nand UO_1503 (O_1503,N_28633,N_29223);
nand UO_1504 (O_1504,N_29001,N_28857);
and UO_1505 (O_1505,N_29583,N_28665);
xnor UO_1506 (O_1506,N_28872,N_29335);
xnor UO_1507 (O_1507,N_29683,N_29803);
or UO_1508 (O_1508,N_28952,N_29175);
nor UO_1509 (O_1509,N_29729,N_28825);
or UO_1510 (O_1510,N_29988,N_28748);
nand UO_1511 (O_1511,N_29768,N_29525);
nor UO_1512 (O_1512,N_28603,N_29209);
or UO_1513 (O_1513,N_28942,N_29338);
or UO_1514 (O_1514,N_28540,N_29052);
or UO_1515 (O_1515,N_29971,N_29262);
nand UO_1516 (O_1516,N_29117,N_28795);
nand UO_1517 (O_1517,N_29470,N_28577);
nand UO_1518 (O_1518,N_29587,N_29327);
or UO_1519 (O_1519,N_29678,N_29857);
nand UO_1520 (O_1520,N_29683,N_28603);
nand UO_1521 (O_1521,N_28831,N_29691);
nand UO_1522 (O_1522,N_29461,N_28875);
or UO_1523 (O_1523,N_29974,N_29727);
xor UO_1524 (O_1524,N_29138,N_29664);
nand UO_1525 (O_1525,N_29168,N_28609);
or UO_1526 (O_1526,N_29540,N_29693);
or UO_1527 (O_1527,N_29836,N_29564);
and UO_1528 (O_1528,N_29090,N_28881);
or UO_1529 (O_1529,N_29812,N_29399);
xor UO_1530 (O_1530,N_29588,N_29242);
xor UO_1531 (O_1531,N_29778,N_29483);
nand UO_1532 (O_1532,N_28966,N_29739);
xor UO_1533 (O_1533,N_29752,N_29809);
and UO_1534 (O_1534,N_29592,N_29211);
and UO_1535 (O_1535,N_29655,N_28916);
and UO_1536 (O_1536,N_29827,N_29872);
xor UO_1537 (O_1537,N_29706,N_29366);
xnor UO_1538 (O_1538,N_29494,N_28500);
or UO_1539 (O_1539,N_28819,N_29847);
xor UO_1540 (O_1540,N_28765,N_29490);
nor UO_1541 (O_1541,N_29350,N_29296);
and UO_1542 (O_1542,N_28862,N_29789);
nand UO_1543 (O_1543,N_29821,N_28797);
or UO_1544 (O_1544,N_28999,N_28749);
xor UO_1545 (O_1545,N_29007,N_29246);
nand UO_1546 (O_1546,N_29077,N_29315);
or UO_1547 (O_1547,N_29786,N_28989);
nand UO_1548 (O_1548,N_28934,N_28643);
and UO_1549 (O_1549,N_29175,N_28988);
and UO_1550 (O_1550,N_28904,N_29122);
nand UO_1551 (O_1551,N_28852,N_29460);
xnor UO_1552 (O_1552,N_29306,N_28574);
or UO_1553 (O_1553,N_29737,N_28931);
or UO_1554 (O_1554,N_29970,N_29988);
nand UO_1555 (O_1555,N_29599,N_29313);
or UO_1556 (O_1556,N_28961,N_29229);
nand UO_1557 (O_1557,N_29686,N_29850);
nand UO_1558 (O_1558,N_29008,N_28661);
and UO_1559 (O_1559,N_29234,N_28648);
xnor UO_1560 (O_1560,N_28561,N_29917);
xor UO_1561 (O_1561,N_29513,N_28512);
or UO_1562 (O_1562,N_28912,N_29865);
nor UO_1563 (O_1563,N_29844,N_29193);
nor UO_1564 (O_1564,N_29636,N_29289);
nor UO_1565 (O_1565,N_29685,N_29065);
xnor UO_1566 (O_1566,N_28953,N_29191);
xor UO_1567 (O_1567,N_29483,N_29245);
nand UO_1568 (O_1568,N_29618,N_28518);
xor UO_1569 (O_1569,N_28546,N_29850);
and UO_1570 (O_1570,N_29917,N_29405);
nor UO_1571 (O_1571,N_29573,N_28691);
nand UO_1572 (O_1572,N_29013,N_28704);
and UO_1573 (O_1573,N_29722,N_28517);
or UO_1574 (O_1574,N_29465,N_28722);
or UO_1575 (O_1575,N_29704,N_29037);
nand UO_1576 (O_1576,N_29015,N_28515);
and UO_1577 (O_1577,N_29218,N_28992);
xnor UO_1578 (O_1578,N_29335,N_29409);
and UO_1579 (O_1579,N_29067,N_29882);
or UO_1580 (O_1580,N_29980,N_29248);
nor UO_1581 (O_1581,N_29286,N_28604);
nor UO_1582 (O_1582,N_29618,N_28992);
nor UO_1583 (O_1583,N_28902,N_29291);
nor UO_1584 (O_1584,N_28697,N_29306);
nor UO_1585 (O_1585,N_29005,N_28737);
nand UO_1586 (O_1586,N_28726,N_28564);
xor UO_1587 (O_1587,N_29514,N_28883);
xor UO_1588 (O_1588,N_29519,N_29993);
xor UO_1589 (O_1589,N_28518,N_28791);
or UO_1590 (O_1590,N_28903,N_29751);
nand UO_1591 (O_1591,N_28920,N_29210);
xor UO_1592 (O_1592,N_29541,N_28854);
or UO_1593 (O_1593,N_29013,N_28644);
or UO_1594 (O_1594,N_28928,N_28785);
or UO_1595 (O_1595,N_29374,N_29104);
or UO_1596 (O_1596,N_29035,N_29462);
and UO_1597 (O_1597,N_28533,N_29860);
and UO_1598 (O_1598,N_28723,N_29203);
xnor UO_1599 (O_1599,N_29323,N_28580);
and UO_1600 (O_1600,N_28753,N_29934);
or UO_1601 (O_1601,N_29100,N_29126);
or UO_1602 (O_1602,N_28716,N_29697);
nor UO_1603 (O_1603,N_28802,N_29518);
nand UO_1604 (O_1604,N_28511,N_28542);
xor UO_1605 (O_1605,N_29447,N_28629);
xnor UO_1606 (O_1606,N_28529,N_28764);
xnor UO_1607 (O_1607,N_29521,N_29455);
or UO_1608 (O_1608,N_29077,N_29078);
nand UO_1609 (O_1609,N_29074,N_29744);
and UO_1610 (O_1610,N_29007,N_29053);
xor UO_1611 (O_1611,N_29148,N_29749);
xnor UO_1612 (O_1612,N_29553,N_29029);
and UO_1613 (O_1613,N_29442,N_28508);
nor UO_1614 (O_1614,N_29704,N_29546);
xnor UO_1615 (O_1615,N_29442,N_29168);
and UO_1616 (O_1616,N_29105,N_29572);
nand UO_1617 (O_1617,N_29876,N_28884);
or UO_1618 (O_1618,N_28729,N_29384);
and UO_1619 (O_1619,N_29013,N_28811);
xor UO_1620 (O_1620,N_29655,N_28787);
or UO_1621 (O_1621,N_29987,N_28682);
nor UO_1622 (O_1622,N_29598,N_28593);
xor UO_1623 (O_1623,N_29385,N_29459);
and UO_1624 (O_1624,N_29249,N_28551);
or UO_1625 (O_1625,N_28586,N_28588);
xor UO_1626 (O_1626,N_29420,N_29349);
nor UO_1627 (O_1627,N_29966,N_28897);
nand UO_1628 (O_1628,N_29349,N_29099);
nor UO_1629 (O_1629,N_29429,N_28755);
and UO_1630 (O_1630,N_29966,N_28895);
xor UO_1631 (O_1631,N_29020,N_29236);
nor UO_1632 (O_1632,N_29177,N_28682);
and UO_1633 (O_1633,N_28977,N_28626);
or UO_1634 (O_1634,N_28710,N_29275);
and UO_1635 (O_1635,N_28553,N_29179);
xnor UO_1636 (O_1636,N_29269,N_28994);
xnor UO_1637 (O_1637,N_29476,N_29489);
xor UO_1638 (O_1638,N_29086,N_29496);
xor UO_1639 (O_1639,N_29795,N_29812);
xor UO_1640 (O_1640,N_28567,N_29144);
xor UO_1641 (O_1641,N_29367,N_28980);
xor UO_1642 (O_1642,N_28704,N_29179);
or UO_1643 (O_1643,N_28669,N_29773);
and UO_1644 (O_1644,N_28780,N_28688);
or UO_1645 (O_1645,N_28778,N_29262);
xnor UO_1646 (O_1646,N_29631,N_29320);
xnor UO_1647 (O_1647,N_29322,N_29768);
and UO_1648 (O_1648,N_29889,N_29662);
xnor UO_1649 (O_1649,N_29862,N_29472);
nand UO_1650 (O_1650,N_29336,N_29752);
or UO_1651 (O_1651,N_29917,N_28528);
and UO_1652 (O_1652,N_29169,N_28626);
or UO_1653 (O_1653,N_28616,N_29095);
nor UO_1654 (O_1654,N_28810,N_29988);
and UO_1655 (O_1655,N_29827,N_29012);
or UO_1656 (O_1656,N_28955,N_28715);
or UO_1657 (O_1657,N_28569,N_28912);
and UO_1658 (O_1658,N_29528,N_29372);
nor UO_1659 (O_1659,N_28645,N_28721);
or UO_1660 (O_1660,N_29774,N_29186);
nand UO_1661 (O_1661,N_29000,N_28649);
nor UO_1662 (O_1662,N_29178,N_29009);
and UO_1663 (O_1663,N_29124,N_29503);
nand UO_1664 (O_1664,N_29822,N_29874);
or UO_1665 (O_1665,N_29662,N_29989);
or UO_1666 (O_1666,N_28867,N_29123);
nand UO_1667 (O_1667,N_28673,N_28633);
and UO_1668 (O_1668,N_28530,N_29317);
nor UO_1669 (O_1669,N_29597,N_29295);
nor UO_1670 (O_1670,N_29023,N_29789);
nand UO_1671 (O_1671,N_28867,N_29722);
nor UO_1672 (O_1672,N_29801,N_29236);
and UO_1673 (O_1673,N_29699,N_29588);
xnor UO_1674 (O_1674,N_28737,N_29359);
xnor UO_1675 (O_1675,N_29786,N_29046);
and UO_1676 (O_1676,N_28825,N_28636);
and UO_1677 (O_1677,N_29357,N_28614);
or UO_1678 (O_1678,N_29260,N_29635);
nor UO_1679 (O_1679,N_28764,N_29683);
nor UO_1680 (O_1680,N_29584,N_29548);
and UO_1681 (O_1681,N_29185,N_28776);
and UO_1682 (O_1682,N_29639,N_29225);
nand UO_1683 (O_1683,N_29601,N_29826);
nand UO_1684 (O_1684,N_29057,N_29803);
or UO_1685 (O_1685,N_28561,N_29573);
and UO_1686 (O_1686,N_29875,N_29544);
and UO_1687 (O_1687,N_29380,N_29745);
nand UO_1688 (O_1688,N_29824,N_28549);
nor UO_1689 (O_1689,N_28785,N_29513);
nand UO_1690 (O_1690,N_29360,N_28925);
xnor UO_1691 (O_1691,N_29146,N_29454);
nand UO_1692 (O_1692,N_29709,N_29066);
nand UO_1693 (O_1693,N_29215,N_29859);
nor UO_1694 (O_1694,N_29788,N_28625);
and UO_1695 (O_1695,N_29603,N_28702);
nand UO_1696 (O_1696,N_29054,N_28634);
nand UO_1697 (O_1697,N_28534,N_28984);
nor UO_1698 (O_1698,N_29057,N_29461);
and UO_1699 (O_1699,N_29662,N_29148);
and UO_1700 (O_1700,N_29205,N_28686);
or UO_1701 (O_1701,N_29177,N_29801);
nor UO_1702 (O_1702,N_28570,N_29466);
and UO_1703 (O_1703,N_28636,N_29621);
nand UO_1704 (O_1704,N_29256,N_29072);
nand UO_1705 (O_1705,N_28689,N_28505);
or UO_1706 (O_1706,N_28916,N_28792);
or UO_1707 (O_1707,N_28817,N_28646);
nand UO_1708 (O_1708,N_28660,N_28639);
nand UO_1709 (O_1709,N_28929,N_29121);
xor UO_1710 (O_1710,N_28550,N_29484);
nor UO_1711 (O_1711,N_29935,N_29371);
xor UO_1712 (O_1712,N_29109,N_29998);
and UO_1713 (O_1713,N_29641,N_29834);
xor UO_1714 (O_1714,N_28878,N_29047);
nor UO_1715 (O_1715,N_29225,N_29873);
or UO_1716 (O_1716,N_29078,N_29477);
or UO_1717 (O_1717,N_28979,N_28774);
nor UO_1718 (O_1718,N_28859,N_28614);
and UO_1719 (O_1719,N_29109,N_29054);
xnor UO_1720 (O_1720,N_29484,N_28741);
or UO_1721 (O_1721,N_29625,N_29905);
and UO_1722 (O_1722,N_29231,N_29002);
xor UO_1723 (O_1723,N_28683,N_29193);
nor UO_1724 (O_1724,N_29200,N_29540);
nand UO_1725 (O_1725,N_28610,N_29746);
nand UO_1726 (O_1726,N_29604,N_29536);
xnor UO_1727 (O_1727,N_29785,N_29827);
nand UO_1728 (O_1728,N_29302,N_29531);
nand UO_1729 (O_1729,N_28534,N_28702);
xnor UO_1730 (O_1730,N_29996,N_28696);
xnor UO_1731 (O_1731,N_28928,N_28818);
nor UO_1732 (O_1732,N_29072,N_29543);
or UO_1733 (O_1733,N_29770,N_29793);
or UO_1734 (O_1734,N_28842,N_28866);
and UO_1735 (O_1735,N_28721,N_29313);
nand UO_1736 (O_1736,N_29524,N_29315);
nor UO_1737 (O_1737,N_29131,N_29050);
or UO_1738 (O_1738,N_29365,N_28679);
nand UO_1739 (O_1739,N_28965,N_28540);
nand UO_1740 (O_1740,N_28688,N_28580);
and UO_1741 (O_1741,N_28989,N_28927);
and UO_1742 (O_1742,N_29612,N_28555);
or UO_1743 (O_1743,N_28658,N_29632);
or UO_1744 (O_1744,N_29782,N_29757);
or UO_1745 (O_1745,N_29925,N_28696);
and UO_1746 (O_1746,N_29375,N_29852);
xor UO_1747 (O_1747,N_28934,N_29622);
xor UO_1748 (O_1748,N_29079,N_29162);
nor UO_1749 (O_1749,N_28737,N_29851);
or UO_1750 (O_1750,N_29674,N_29772);
or UO_1751 (O_1751,N_29101,N_29035);
or UO_1752 (O_1752,N_29490,N_29998);
nand UO_1753 (O_1753,N_29475,N_29248);
xnor UO_1754 (O_1754,N_28733,N_28813);
nand UO_1755 (O_1755,N_29030,N_28977);
nand UO_1756 (O_1756,N_29271,N_29104);
nor UO_1757 (O_1757,N_28924,N_29362);
or UO_1758 (O_1758,N_29707,N_29109);
nor UO_1759 (O_1759,N_29587,N_28684);
xor UO_1760 (O_1760,N_29843,N_29065);
and UO_1761 (O_1761,N_28996,N_29367);
and UO_1762 (O_1762,N_28985,N_29369);
xor UO_1763 (O_1763,N_28617,N_29741);
nor UO_1764 (O_1764,N_29653,N_28613);
nand UO_1765 (O_1765,N_28618,N_28950);
xor UO_1766 (O_1766,N_29693,N_29253);
xnor UO_1767 (O_1767,N_29848,N_28802);
or UO_1768 (O_1768,N_28859,N_28590);
nor UO_1769 (O_1769,N_28657,N_29775);
xor UO_1770 (O_1770,N_29621,N_29433);
nand UO_1771 (O_1771,N_29882,N_29943);
nand UO_1772 (O_1772,N_29771,N_28641);
nor UO_1773 (O_1773,N_29270,N_28924);
nand UO_1774 (O_1774,N_29197,N_29271);
xnor UO_1775 (O_1775,N_29115,N_29043);
or UO_1776 (O_1776,N_28528,N_28732);
or UO_1777 (O_1777,N_28814,N_29469);
xnor UO_1778 (O_1778,N_29333,N_28664);
or UO_1779 (O_1779,N_29683,N_29664);
nand UO_1780 (O_1780,N_28875,N_29652);
or UO_1781 (O_1781,N_29376,N_29490);
nor UO_1782 (O_1782,N_29740,N_29860);
xor UO_1783 (O_1783,N_29101,N_29919);
and UO_1784 (O_1784,N_29498,N_28520);
nor UO_1785 (O_1785,N_28839,N_29881);
and UO_1786 (O_1786,N_29603,N_28843);
or UO_1787 (O_1787,N_29622,N_28557);
and UO_1788 (O_1788,N_29153,N_29439);
xnor UO_1789 (O_1789,N_29520,N_29628);
nor UO_1790 (O_1790,N_29294,N_29520);
xnor UO_1791 (O_1791,N_29378,N_29339);
and UO_1792 (O_1792,N_29554,N_29031);
nor UO_1793 (O_1793,N_29831,N_29944);
nor UO_1794 (O_1794,N_28676,N_29853);
or UO_1795 (O_1795,N_29553,N_28780);
xor UO_1796 (O_1796,N_29822,N_29574);
or UO_1797 (O_1797,N_28840,N_29090);
and UO_1798 (O_1798,N_28898,N_29005);
and UO_1799 (O_1799,N_28525,N_28970);
and UO_1800 (O_1800,N_29953,N_29565);
or UO_1801 (O_1801,N_29553,N_29745);
or UO_1802 (O_1802,N_29254,N_28802);
xor UO_1803 (O_1803,N_29291,N_29805);
or UO_1804 (O_1804,N_29647,N_28811);
nand UO_1805 (O_1805,N_29029,N_29883);
or UO_1806 (O_1806,N_29057,N_29574);
xor UO_1807 (O_1807,N_28895,N_28513);
nor UO_1808 (O_1808,N_29382,N_28783);
xnor UO_1809 (O_1809,N_28830,N_28784);
or UO_1810 (O_1810,N_29506,N_29453);
and UO_1811 (O_1811,N_29106,N_29243);
xnor UO_1812 (O_1812,N_29768,N_29302);
nand UO_1813 (O_1813,N_29265,N_29262);
xnor UO_1814 (O_1814,N_29175,N_29045);
and UO_1815 (O_1815,N_29175,N_29962);
or UO_1816 (O_1816,N_29284,N_28599);
and UO_1817 (O_1817,N_28961,N_28739);
xnor UO_1818 (O_1818,N_28595,N_29718);
nand UO_1819 (O_1819,N_29439,N_28895);
nand UO_1820 (O_1820,N_28910,N_28935);
or UO_1821 (O_1821,N_29616,N_29063);
nand UO_1822 (O_1822,N_29759,N_29713);
and UO_1823 (O_1823,N_29864,N_28558);
nand UO_1824 (O_1824,N_29487,N_29294);
and UO_1825 (O_1825,N_29735,N_28980);
or UO_1826 (O_1826,N_29387,N_28985);
nor UO_1827 (O_1827,N_28828,N_29879);
nor UO_1828 (O_1828,N_28619,N_28993);
nand UO_1829 (O_1829,N_29815,N_29591);
or UO_1830 (O_1830,N_28598,N_28613);
nand UO_1831 (O_1831,N_29602,N_28788);
and UO_1832 (O_1832,N_28930,N_29990);
xor UO_1833 (O_1833,N_29787,N_29239);
or UO_1834 (O_1834,N_29566,N_29388);
nand UO_1835 (O_1835,N_28770,N_29838);
and UO_1836 (O_1836,N_28762,N_29581);
and UO_1837 (O_1837,N_29357,N_29503);
or UO_1838 (O_1838,N_29342,N_29597);
xnor UO_1839 (O_1839,N_29034,N_29164);
nand UO_1840 (O_1840,N_28976,N_28565);
or UO_1841 (O_1841,N_28922,N_29920);
xor UO_1842 (O_1842,N_29135,N_28886);
or UO_1843 (O_1843,N_29351,N_28650);
nand UO_1844 (O_1844,N_28994,N_28753);
nand UO_1845 (O_1845,N_29911,N_28608);
or UO_1846 (O_1846,N_29820,N_28733);
nor UO_1847 (O_1847,N_29742,N_28727);
xnor UO_1848 (O_1848,N_28613,N_29352);
and UO_1849 (O_1849,N_29122,N_29746);
nor UO_1850 (O_1850,N_29423,N_29114);
nor UO_1851 (O_1851,N_29813,N_29401);
or UO_1852 (O_1852,N_28944,N_28842);
xor UO_1853 (O_1853,N_29235,N_29000);
nor UO_1854 (O_1854,N_29383,N_28841);
xnor UO_1855 (O_1855,N_29627,N_28724);
or UO_1856 (O_1856,N_29199,N_29098);
nand UO_1857 (O_1857,N_29236,N_29515);
nand UO_1858 (O_1858,N_29371,N_28908);
xnor UO_1859 (O_1859,N_28710,N_29990);
nand UO_1860 (O_1860,N_29738,N_29832);
nor UO_1861 (O_1861,N_29365,N_28871);
nand UO_1862 (O_1862,N_29181,N_29811);
nand UO_1863 (O_1863,N_29873,N_28566);
nor UO_1864 (O_1864,N_28700,N_28990);
nor UO_1865 (O_1865,N_29036,N_29777);
nand UO_1866 (O_1866,N_28743,N_28533);
or UO_1867 (O_1867,N_28738,N_29088);
nor UO_1868 (O_1868,N_28529,N_29081);
nor UO_1869 (O_1869,N_29290,N_28918);
and UO_1870 (O_1870,N_28921,N_28902);
nand UO_1871 (O_1871,N_29586,N_28852);
nor UO_1872 (O_1872,N_29995,N_28795);
nand UO_1873 (O_1873,N_29322,N_28705);
xor UO_1874 (O_1874,N_29179,N_29071);
and UO_1875 (O_1875,N_28648,N_28805);
nand UO_1876 (O_1876,N_29563,N_29222);
and UO_1877 (O_1877,N_29177,N_28571);
and UO_1878 (O_1878,N_29305,N_28709);
or UO_1879 (O_1879,N_28974,N_29419);
and UO_1880 (O_1880,N_29897,N_29953);
and UO_1881 (O_1881,N_28624,N_29728);
nor UO_1882 (O_1882,N_29579,N_29227);
xnor UO_1883 (O_1883,N_29115,N_29234);
nand UO_1884 (O_1884,N_29476,N_29117);
and UO_1885 (O_1885,N_28792,N_28748);
nor UO_1886 (O_1886,N_28940,N_29588);
and UO_1887 (O_1887,N_29131,N_29942);
nand UO_1888 (O_1888,N_29331,N_29017);
or UO_1889 (O_1889,N_29371,N_28878);
and UO_1890 (O_1890,N_28704,N_28705);
and UO_1891 (O_1891,N_29003,N_29099);
or UO_1892 (O_1892,N_29382,N_29844);
xnor UO_1893 (O_1893,N_29141,N_29867);
and UO_1894 (O_1894,N_29205,N_29650);
nand UO_1895 (O_1895,N_28679,N_28991);
or UO_1896 (O_1896,N_28557,N_28584);
nor UO_1897 (O_1897,N_29119,N_29660);
nor UO_1898 (O_1898,N_28941,N_29983);
nand UO_1899 (O_1899,N_28722,N_29413);
xor UO_1900 (O_1900,N_29036,N_29161);
or UO_1901 (O_1901,N_28535,N_29106);
and UO_1902 (O_1902,N_29839,N_29009);
or UO_1903 (O_1903,N_29788,N_28941);
nand UO_1904 (O_1904,N_29603,N_29506);
or UO_1905 (O_1905,N_28846,N_29390);
and UO_1906 (O_1906,N_28796,N_29727);
nand UO_1907 (O_1907,N_29519,N_28770);
xor UO_1908 (O_1908,N_29100,N_28715);
or UO_1909 (O_1909,N_29535,N_29838);
xnor UO_1910 (O_1910,N_29571,N_29384);
xor UO_1911 (O_1911,N_29788,N_29271);
nor UO_1912 (O_1912,N_28575,N_29003);
nand UO_1913 (O_1913,N_29929,N_29490);
nor UO_1914 (O_1914,N_29992,N_29675);
xnor UO_1915 (O_1915,N_29548,N_29856);
or UO_1916 (O_1916,N_29763,N_29130);
nor UO_1917 (O_1917,N_28671,N_28698);
nand UO_1918 (O_1918,N_29294,N_29560);
nand UO_1919 (O_1919,N_28604,N_29069);
or UO_1920 (O_1920,N_28651,N_29882);
nand UO_1921 (O_1921,N_29966,N_29089);
xor UO_1922 (O_1922,N_29618,N_29955);
or UO_1923 (O_1923,N_29630,N_29466);
xnor UO_1924 (O_1924,N_29670,N_29042);
or UO_1925 (O_1925,N_29920,N_28764);
or UO_1926 (O_1926,N_29109,N_29641);
nor UO_1927 (O_1927,N_28541,N_29818);
nand UO_1928 (O_1928,N_29783,N_29755);
xnor UO_1929 (O_1929,N_29777,N_28604);
or UO_1930 (O_1930,N_28543,N_29960);
or UO_1931 (O_1931,N_29646,N_29154);
nor UO_1932 (O_1932,N_28687,N_29965);
nor UO_1933 (O_1933,N_29107,N_28952);
xor UO_1934 (O_1934,N_29112,N_28576);
nand UO_1935 (O_1935,N_28611,N_29729);
and UO_1936 (O_1936,N_29337,N_29784);
xor UO_1937 (O_1937,N_28561,N_29501);
nor UO_1938 (O_1938,N_29265,N_29506);
and UO_1939 (O_1939,N_29891,N_29767);
nor UO_1940 (O_1940,N_29172,N_28901);
xor UO_1941 (O_1941,N_29828,N_29132);
xor UO_1942 (O_1942,N_28732,N_29413);
xnor UO_1943 (O_1943,N_29249,N_28921);
or UO_1944 (O_1944,N_29795,N_28619);
xor UO_1945 (O_1945,N_29815,N_29304);
nor UO_1946 (O_1946,N_29757,N_29491);
and UO_1947 (O_1947,N_28811,N_29402);
xor UO_1948 (O_1948,N_28714,N_29353);
nand UO_1949 (O_1949,N_29857,N_28532);
nor UO_1950 (O_1950,N_29272,N_29737);
and UO_1951 (O_1951,N_28662,N_28758);
or UO_1952 (O_1952,N_29504,N_29970);
xor UO_1953 (O_1953,N_29161,N_29422);
nor UO_1954 (O_1954,N_28870,N_29649);
or UO_1955 (O_1955,N_28945,N_28641);
and UO_1956 (O_1956,N_29305,N_29264);
nand UO_1957 (O_1957,N_29492,N_29807);
and UO_1958 (O_1958,N_29869,N_29207);
nand UO_1959 (O_1959,N_29658,N_29426);
nand UO_1960 (O_1960,N_29187,N_29776);
xor UO_1961 (O_1961,N_28801,N_29639);
or UO_1962 (O_1962,N_28670,N_29511);
xnor UO_1963 (O_1963,N_29352,N_29140);
and UO_1964 (O_1964,N_29404,N_29904);
or UO_1965 (O_1965,N_29898,N_29743);
and UO_1966 (O_1966,N_29104,N_28537);
and UO_1967 (O_1967,N_28758,N_28920);
or UO_1968 (O_1968,N_29969,N_29280);
xnor UO_1969 (O_1969,N_29749,N_29705);
nor UO_1970 (O_1970,N_29060,N_29109);
nand UO_1971 (O_1971,N_28713,N_28655);
xor UO_1972 (O_1972,N_28832,N_29812);
or UO_1973 (O_1973,N_28781,N_28974);
and UO_1974 (O_1974,N_29568,N_28902);
xor UO_1975 (O_1975,N_28625,N_29924);
or UO_1976 (O_1976,N_29360,N_29614);
or UO_1977 (O_1977,N_29952,N_29727);
nor UO_1978 (O_1978,N_29791,N_29771);
or UO_1979 (O_1979,N_28760,N_28516);
xnor UO_1980 (O_1980,N_28576,N_29730);
and UO_1981 (O_1981,N_29466,N_29526);
xnor UO_1982 (O_1982,N_28647,N_28889);
nor UO_1983 (O_1983,N_28536,N_29669);
nor UO_1984 (O_1984,N_28676,N_29860);
nand UO_1985 (O_1985,N_28784,N_28838);
and UO_1986 (O_1986,N_29231,N_29091);
nand UO_1987 (O_1987,N_28807,N_29908);
xnor UO_1988 (O_1988,N_29069,N_29336);
nand UO_1989 (O_1989,N_29603,N_29687);
and UO_1990 (O_1990,N_29701,N_29574);
and UO_1991 (O_1991,N_28925,N_29151);
nand UO_1992 (O_1992,N_29018,N_28531);
xnor UO_1993 (O_1993,N_29123,N_28982);
nor UO_1994 (O_1994,N_29774,N_29948);
nor UO_1995 (O_1995,N_29004,N_29777);
nor UO_1996 (O_1996,N_28575,N_28909);
xor UO_1997 (O_1997,N_29002,N_29890);
or UO_1998 (O_1998,N_29318,N_29630);
nor UO_1999 (O_1999,N_28620,N_29991);
or UO_2000 (O_2000,N_29630,N_29756);
nor UO_2001 (O_2001,N_28846,N_29951);
nor UO_2002 (O_2002,N_28629,N_29546);
or UO_2003 (O_2003,N_29297,N_29408);
xor UO_2004 (O_2004,N_29730,N_29190);
or UO_2005 (O_2005,N_29847,N_28690);
nor UO_2006 (O_2006,N_29071,N_29579);
nand UO_2007 (O_2007,N_28748,N_29570);
nand UO_2008 (O_2008,N_29867,N_28541);
and UO_2009 (O_2009,N_28787,N_29587);
and UO_2010 (O_2010,N_29861,N_29370);
or UO_2011 (O_2011,N_28817,N_29633);
nand UO_2012 (O_2012,N_28568,N_29616);
nor UO_2013 (O_2013,N_29976,N_28506);
xnor UO_2014 (O_2014,N_29008,N_29521);
nand UO_2015 (O_2015,N_28510,N_29474);
and UO_2016 (O_2016,N_28952,N_29901);
and UO_2017 (O_2017,N_29140,N_29939);
xor UO_2018 (O_2018,N_29269,N_29537);
or UO_2019 (O_2019,N_28523,N_29094);
nand UO_2020 (O_2020,N_29306,N_29843);
xnor UO_2021 (O_2021,N_29276,N_29083);
xnor UO_2022 (O_2022,N_28730,N_28504);
xor UO_2023 (O_2023,N_28631,N_29222);
and UO_2024 (O_2024,N_29159,N_28895);
nand UO_2025 (O_2025,N_29703,N_29462);
nand UO_2026 (O_2026,N_29991,N_29498);
or UO_2027 (O_2027,N_29195,N_29239);
xnor UO_2028 (O_2028,N_29051,N_29630);
xor UO_2029 (O_2029,N_29739,N_29099);
nor UO_2030 (O_2030,N_29820,N_29867);
nor UO_2031 (O_2031,N_29407,N_28520);
xor UO_2032 (O_2032,N_28803,N_28733);
nor UO_2033 (O_2033,N_28697,N_29991);
or UO_2034 (O_2034,N_29710,N_29321);
nand UO_2035 (O_2035,N_28644,N_29638);
xor UO_2036 (O_2036,N_29039,N_29728);
nand UO_2037 (O_2037,N_28563,N_29254);
xor UO_2038 (O_2038,N_29172,N_29481);
and UO_2039 (O_2039,N_29870,N_29520);
or UO_2040 (O_2040,N_29696,N_29076);
nor UO_2041 (O_2041,N_29278,N_28711);
or UO_2042 (O_2042,N_29483,N_29756);
xor UO_2043 (O_2043,N_29069,N_29678);
nor UO_2044 (O_2044,N_29282,N_29465);
or UO_2045 (O_2045,N_28581,N_29683);
and UO_2046 (O_2046,N_29538,N_28987);
nand UO_2047 (O_2047,N_29900,N_29367);
or UO_2048 (O_2048,N_29347,N_29597);
and UO_2049 (O_2049,N_28776,N_28977);
or UO_2050 (O_2050,N_28531,N_28606);
xnor UO_2051 (O_2051,N_29759,N_29950);
nor UO_2052 (O_2052,N_28602,N_29822);
and UO_2053 (O_2053,N_29886,N_28779);
and UO_2054 (O_2054,N_29777,N_29020);
nand UO_2055 (O_2055,N_28871,N_29563);
nand UO_2056 (O_2056,N_29977,N_29899);
nand UO_2057 (O_2057,N_29297,N_29156);
nand UO_2058 (O_2058,N_29418,N_29489);
xor UO_2059 (O_2059,N_29872,N_29360);
and UO_2060 (O_2060,N_28565,N_28985);
nand UO_2061 (O_2061,N_29154,N_29009);
and UO_2062 (O_2062,N_29495,N_29611);
nor UO_2063 (O_2063,N_29807,N_28588);
nand UO_2064 (O_2064,N_28937,N_29327);
nand UO_2065 (O_2065,N_29016,N_29362);
xor UO_2066 (O_2066,N_29650,N_29469);
xor UO_2067 (O_2067,N_29307,N_29619);
nand UO_2068 (O_2068,N_29170,N_28500);
nor UO_2069 (O_2069,N_28513,N_29798);
or UO_2070 (O_2070,N_29687,N_29331);
or UO_2071 (O_2071,N_29364,N_29803);
or UO_2072 (O_2072,N_29539,N_29005);
nor UO_2073 (O_2073,N_28778,N_29998);
xor UO_2074 (O_2074,N_29547,N_29481);
nand UO_2075 (O_2075,N_29212,N_29476);
or UO_2076 (O_2076,N_29071,N_29254);
or UO_2077 (O_2077,N_29771,N_28803);
xor UO_2078 (O_2078,N_29586,N_28833);
or UO_2079 (O_2079,N_29679,N_29728);
nand UO_2080 (O_2080,N_28584,N_29920);
and UO_2081 (O_2081,N_29186,N_28950);
nor UO_2082 (O_2082,N_28868,N_28578);
or UO_2083 (O_2083,N_29996,N_29513);
or UO_2084 (O_2084,N_29176,N_28893);
xnor UO_2085 (O_2085,N_28988,N_29418);
or UO_2086 (O_2086,N_28628,N_29630);
and UO_2087 (O_2087,N_28704,N_29096);
and UO_2088 (O_2088,N_29025,N_29874);
xnor UO_2089 (O_2089,N_29310,N_29731);
nor UO_2090 (O_2090,N_28693,N_29251);
xor UO_2091 (O_2091,N_29999,N_29590);
nor UO_2092 (O_2092,N_29335,N_28752);
or UO_2093 (O_2093,N_29501,N_28633);
and UO_2094 (O_2094,N_29158,N_28905);
nand UO_2095 (O_2095,N_29133,N_29012);
nand UO_2096 (O_2096,N_28662,N_29256);
and UO_2097 (O_2097,N_29210,N_29906);
and UO_2098 (O_2098,N_29725,N_29017);
xor UO_2099 (O_2099,N_29084,N_28903);
xor UO_2100 (O_2100,N_29892,N_28695);
nor UO_2101 (O_2101,N_29577,N_29918);
and UO_2102 (O_2102,N_29991,N_29857);
xnor UO_2103 (O_2103,N_29107,N_29228);
xor UO_2104 (O_2104,N_29068,N_29990);
xnor UO_2105 (O_2105,N_28557,N_28849);
nand UO_2106 (O_2106,N_29545,N_29017);
and UO_2107 (O_2107,N_28731,N_29809);
xor UO_2108 (O_2108,N_29282,N_28884);
and UO_2109 (O_2109,N_28537,N_29805);
nor UO_2110 (O_2110,N_29425,N_29559);
nor UO_2111 (O_2111,N_28532,N_29983);
and UO_2112 (O_2112,N_29386,N_28816);
or UO_2113 (O_2113,N_29399,N_28822);
and UO_2114 (O_2114,N_29046,N_29575);
nand UO_2115 (O_2115,N_28618,N_29487);
or UO_2116 (O_2116,N_29679,N_29641);
nand UO_2117 (O_2117,N_29884,N_28977);
and UO_2118 (O_2118,N_28582,N_28917);
and UO_2119 (O_2119,N_29993,N_28996);
nand UO_2120 (O_2120,N_28627,N_29327);
or UO_2121 (O_2121,N_28671,N_29114);
and UO_2122 (O_2122,N_29033,N_29909);
or UO_2123 (O_2123,N_28603,N_29930);
nand UO_2124 (O_2124,N_29797,N_29105);
and UO_2125 (O_2125,N_28805,N_29880);
nor UO_2126 (O_2126,N_29909,N_29639);
or UO_2127 (O_2127,N_28523,N_29111);
and UO_2128 (O_2128,N_28991,N_28623);
xor UO_2129 (O_2129,N_29724,N_29318);
nand UO_2130 (O_2130,N_28818,N_28772);
nor UO_2131 (O_2131,N_29691,N_29007);
or UO_2132 (O_2132,N_28961,N_29996);
or UO_2133 (O_2133,N_29456,N_29235);
or UO_2134 (O_2134,N_29426,N_29906);
xnor UO_2135 (O_2135,N_29142,N_29757);
nand UO_2136 (O_2136,N_28588,N_28836);
nand UO_2137 (O_2137,N_29490,N_29657);
nor UO_2138 (O_2138,N_29271,N_29907);
or UO_2139 (O_2139,N_29039,N_29969);
nand UO_2140 (O_2140,N_28686,N_28924);
or UO_2141 (O_2141,N_28881,N_29376);
nand UO_2142 (O_2142,N_28628,N_29954);
nand UO_2143 (O_2143,N_29926,N_28595);
nor UO_2144 (O_2144,N_29539,N_29671);
or UO_2145 (O_2145,N_29816,N_28953);
nand UO_2146 (O_2146,N_29843,N_29378);
nand UO_2147 (O_2147,N_28655,N_29367);
nand UO_2148 (O_2148,N_29264,N_28864);
nor UO_2149 (O_2149,N_28916,N_29927);
xor UO_2150 (O_2150,N_29732,N_28945);
nand UO_2151 (O_2151,N_29602,N_28676);
xnor UO_2152 (O_2152,N_29752,N_29597);
or UO_2153 (O_2153,N_29668,N_28550);
and UO_2154 (O_2154,N_28891,N_29373);
xor UO_2155 (O_2155,N_29846,N_29280);
or UO_2156 (O_2156,N_28948,N_29612);
or UO_2157 (O_2157,N_29108,N_28985);
and UO_2158 (O_2158,N_29026,N_29284);
and UO_2159 (O_2159,N_28710,N_29431);
xnor UO_2160 (O_2160,N_28656,N_29217);
nor UO_2161 (O_2161,N_29185,N_29077);
nand UO_2162 (O_2162,N_28583,N_29163);
nor UO_2163 (O_2163,N_28997,N_28729);
nor UO_2164 (O_2164,N_29473,N_28634);
nand UO_2165 (O_2165,N_29710,N_28532);
xnor UO_2166 (O_2166,N_29578,N_28864);
xor UO_2167 (O_2167,N_28805,N_29193);
xnor UO_2168 (O_2168,N_29633,N_29565);
or UO_2169 (O_2169,N_29002,N_29203);
xor UO_2170 (O_2170,N_29949,N_29850);
and UO_2171 (O_2171,N_29716,N_29761);
or UO_2172 (O_2172,N_28933,N_28779);
or UO_2173 (O_2173,N_28751,N_29911);
xnor UO_2174 (O_2174,N_29824,N_28763);
xnor UO_2175 (O_2175,N_28757,N_28823);
nor UO_2176 (O_2176,N_29932,N_29609);
nor UO_2177 (O_2177,N_29750,N_29473);
or UO_2178 (O_2178,N_29006,N_29060);
xor UO_2179 (O_2179,N_29508,N_28629);
nand UO_2180 (O_2180,N_29161,N_29100);
nor UO_2181 (O_2181,N_29326,N_29339);
nand UO_2182 (O_2182,N_29274,N_29094);
xor UO_2183 (O_2183,N_28591,N_28581);
or UO_2184 (O_2184,N_28886,N_28681);
nand UO_2185 (O_2185,N_29062,N_29292);
nand UO_2186 (O_2186,N_29551,N_28789);
and UO_2187 (O_2187,N_29743,N_28987);
nor UO_2188 (O_2188,N_29358,N_29788);
nor UO_2189 (O_2189,N_29801,N_28896);
nor UO_2190 (O_2190,N_28673,N_29320);
nand UO_2191 (O_2191,N_29083,N_29665);
and UO_2192 (O_2192,N_29873,N_29480);
nand UO_2193 (O_2193,N_28878,N_29281);
nand UO_2194 (O_2194,N_28910,N_28534);
or UO_2195 (O_2195,N_29145,N_28655);
and UO_2196 (O_2196,N_28671,N_29986);
xnor UO_2197 (O_2197,N_29898,N_29920);
xnor UO_2198 (O_2198,N_29465,N_29952);
or UO_2199 (O_2199,N_29614,N_29671);
xor UO_2200 (O_2200,N_29270,N_29150);
nand UO_2201 (O_2201,N_29944,N_29598);
nor UO_2202 (O_2202,N_29546,N_28966);
xnor UO_2203 (O_2203,N_29995,N_29328);
or UO_2204 (O_2204,N_29747,N_28975);
and UO_2205 (O_2205,N_28676,N_29454);
nor UO_2206 (O_2206,N_29733,N_29275);
or UO_2207 (O_2207,N_29589,N_29568);
nand UO_2208 (O_2208,N_28599,N_28902);
nor UO_2209 (O_2209,N_29923,N_28717);
nor UO_2210 (O_2210,N_29903,N_29807);
nor UO_2211 (O_2211,N_29601,N_29240);
nand UO_2212 (O_2212,N_29623,N_29980);
nor UO_2213 (O_2213,N_29741,N_28720);
nor UO_2214 (O_2214,N_28574,N_29028);
or UO_2215 (O_2215,N_28544,N_29331);
nand UO_2216 (O_2216,N_29872,N_29247);
or UO_2217 (O_2217,N_28746,N_28866);
nand UO_2218 (O_2218,N_29161,N_29152);
or UO_2219 (O_2219,N_28737,N_28592);
nor UO_2220 (O_2220,N_29521,N_29778);
and UO_2221 (O_2221,N_28773,N_28519);
and UO_2222 (O_2222,N_29586,N_29455);
xnor UO_2223 (O_2223,N_28526,N_28896);
xor UO_2224 (O_2224,N_29731,N_28874);
or UO_2225 (O_2225,N_28742,N_29412);
nand UO_2226 (O_2226,N_28760,N_29396);
nor UO_2227 (O_2227,N_28700,N_29700);
nand UO_2228 (O_2228,N_29067,N_29809);
and UO_2229 (O_2229,N_29681,N_29469);
nand UO_2230 (O_2230,N_29976,N_29958);
nor UO_2231 (O_2231,N_29061,N_29660);
and UO_2232 (O_2232,N_29012,N_28873);
nand UO_2233 (O_2233,N_29954,N_29527);
nand UO_2234 (O_2234,N_29694,N_29962);
nand UO_2235 (O_2235,N_29572,N_29672);
xor UO_2236 (O_2236,N_29742,N_28907);
xnor UO_2237 (O_2237,N_29396,N_29264);
and UO_2238 (O_2238,N_29263,N_28988);
and UO_2239 (O_2239,N_28923,N_29093);
xor UO_2240 (O_2240,N_28711,N_29158);
xnor UO_2241 (O_2241,N_28741,N_29651);
and UO_2242 (O_2242,N_28701,N_29464);
and UO_2243 (O_2243,N_29956,N_29311);
xnor UO_2244 (O_2244,N_28592,N_29791);
xor UO_2245 (O_2245,N_29897,N_29610);
and UO_2246 (O_2246,N_29727,N_29609);
and UO_2247 (O_2247,N_28908,N_29585);
nand UO_2248 (O_2248,N_29377,N_29260);
and UO_2249 (O_2249,N_28520,N_28724);
and UO_2250 (O_2250,N_29515,N_29932);
and UO_2251 (O_2251,N_28939,N_29088);
or UO_2252 (O_2252,N_29111,N_29079);
nor UO_2253 (O_2253,N_29901,N_29917);
nand UO_2254 (O_2254,N_29532,N_29821);
or UO_2255 (O_2255,N_29272,N_29642);
or UO_2256 (O_2256,N_29288,N_28811);
nand UO_2257 (O_2257,N_29570,N_29689);
or UO_2258 (O_2258,N_29243,N_28776);
nand UO_2259 (O_2259,N_28891,N_28764);
or UO_2260 (O_2260,N_29545,N_29927);
xnor UO_2261 (O_2261,N_29196,N_29127);
xor UO_2262 (O_2262,N_29955,N_28611);
nand UO_2263 (O_2263,N_29927,N_28870);
nand UO_2264 (O_2264,N_29775,N_29022);
nand UO_2265 (O_2265,N_29677,N_28765);
nand UO_2266 (O_2266,N_29487,N_28975);
and UO_2267 (O_2267,N_28848,N_29514);
xor UO_2268 (O_2268,N_29382,N_29945);
nor UO_2269 (O_2269,N_28983,N_28982);
or UO_2270 (O_2270,N_29220,N_29192);
or UO_2271 (O_2271,N_29180,N_29490);
or UO_2272 (O_2272,N_29234,N_28943);
and UO_2273 (O_2273,N_29261,N_28773);
xor UO_2274 (O_2274,N_28957,N_29043);
nor UO_2275 (O_2275,N_29452,N_29002);
or UO_2276 (O_2276,N_29325,N_29000);
or UO_2277 (O_2277,N_29812,N_28947);
xor UO_2278 (O_2278,N_29377,N_28795);
nand UO_2279 (O_2279,N_29603,N_28789);
or UO_2280 (O_2280,N_29744,N_29700);
and UO_2281 (O_2281,N_29380,N_28637);
or UO_2282 (O_2282,N_28930,N_29730);
and UO_2283 (O_2283,N_29283,N_28894);
nor UO_2284 (O_2284,N_29023,N_29311);
nand UO_2285 (O_2285,N_29268,N_29809);
nand UO_2286 (O_2286,N_29227,N_29534);
xor UO_2287 (O_2287,N_28641,N_28784);
nand UO_2288 (O_2288,N_29230,N_28736);
nor UO_2289 (O_2289,N_29739,N_29358);
nor UO_2290 (O_2290,N_29008,N_28980);
nand UO_2291 (O_2291,N_28703,N_28511);
or UO_2292 (O_2292,N_29704,N_28717);
xor UO_2293 (O_2293,N_28773,N_29777);
xnor UO_2294 (O_2294,N_29690,N_29309);
nor UO_2295 (O_2295,N_29443,N_29954);
nand UO_2296 (O_2296,N_28572,N_29081);
and UO_2297 (O_2297,N_29285,N_28720);
nand UO_2298 (O_2298,N_29253,N_28669);
xnor UO_2299 (O_2299,N_29390,N_29062);
nor UO_2300 (O_2300,N_28946,N_29519);
nand UO_2301 (O_2301,N_29481,N_29092);
and UO_2302 (O_2302,N_28870,N_29223);
or UO_2303 (O_2303,N_29932,N_29257);
or UO_2304 (O_2304,N_29306,N_29783);
xor UO_2305 (O_2305,N_29375,N_29981);
or UO_2306 (O_2306,N_29975,N_28653);
nor UO_2307 (O_2307,N_29560,N_29969);
or UO_2308 (O_2308,N_28953,N_29240);
nand UO_2309 (O_2309,N_29223,N_29024);
nor UO_2310 (O_2310,N_28777,N_29231);
xnor UO_2311 (O_2311,N_29593,N_29337);
xnor UO_2312 (O_2312,N_29482,N_28574);
xor UO_2313 (O_2313,N_28895,N_28812);
nand UO_2314 (O_2314,N_29302,N_29627);
xnor UO_2315 (O_2315,N_29791,N_29870);
nor UO_2316 (O_2316,N_29888,N_29636);
xnor UO_2317 (O_2317,N_29038,N_28847);
and UO_2318 (O_2318,N_28682,N_29940);
nor UO_2319 (O_2319,N_29709,N_28812);
xor UO_2320 (O_2320,N_28992,N_28670);
xor UO_2321 (O_2321,N_29830,N_28869);
and UO_2322 (O_2322,N_28778,N_29661);
and UO_2323 (O_2323,N_29820,N_29034);
nor UO_2324 (O_2324,N_29682,N_28566);
xor UO_2325 (O_2325,N_29291,N_29779);
nor UO_2326 (O_2326,N_29160,N_29865);
and UO_2327 (O_2327,N_29382,N_29808);
or UO_2328 (O_2328,N_28981,N_28877);
xnor UO_2329 (O_2329,N_29390,N_29722);
nand UO_2330 (O_2330,N_28846,N_29582);
and UO_2331 (O_2331,N_28865,N_29466);
or UO_2332 (O_2332,N_28580,N_29055);
and UO_2333 (O_2333,N_28775,N_28712);
nand UO_2334 (O_2334,N_29114,N_29869);
or UO_2335 (O_2335,N_29717,N_29318);
nor UO_2336 (O_2336,N_29791,N_29952);
and UO_2337 (O_2337,N_29655,N_29974);
or UO_2338 (O_2338,N_29189,N_28745);
nor UO_2339 (O_2339,N_29363,N_29510);
or UO_2340 (O_2340,N_29076,N_28777);
and UO_2341 (O_2341,N_29018,N_29528);
xnor UO_2342 (O_2342,N_28698,N_29497);
and UO_2343 (O_2343,N_29161,N_28612);
xor UO_2344 (O_2344,N_29229,N_28700);
and UO_2345 (O_2345,N_29512,N_29902);
xnor UO_2346 (O_2346,N_29347,N_28817);
or UO_2347 (O_2347,N_29033,N_29246);
or UO_2348 (O_2348,N_29609,N_28507);
nor UO_2349 (O_2349,N_29533,N_28753);
xor UO_2350 (O_2350,N_29498,N_29077);
nand UO_2351 (O_2351,N_29104,N_28613);
or UO_2352 (O_2352,N_28732,N_28645);
or UO_2353 (O_2353,N_28845,N_29295);
or UO_2354 (O_2354,N_29237,N_28849);
xor UO_2355 (O_2355,N_29318,N_28673);
nand UO_2356 (O_2356,N_28705,N_29023);
nand UO_2357 (O_2357,N_28876,N_28652);
or UO_2358 (O_2358,N_29224,N_28864);
and UO_2359 (O_2359,N_29946,N_29867);
and UO_2360 (O_2360,N_29303,N_29631);
nand UO_2361 (O_2361,N_28525,N_28564);
nor UO_2362 (O_2362,N_28709,N_29203);
xor UO_2363 (O_2363,N_28734,N_28758);
xnor UO_2364 (O_2364,N_29885,N_28791);
nor UO_2365 (O_2365,N_28842,N_29884);
nand UO_2366 (O_2366,N_28843,N_29067);
nor UO_2367 (O_2367,N_29090,N_28973);
or UO_2368 (O_2368,N_29015,N_28755);
xnor UO_2369 (O_2369,N_29842,N_28509);
or UO_2370 (O_2370,N_29075,N_29482);
nand UO_2371 (O_2371,N_29667,N_28516);
xor UO_2372 (O_2372,N_29484,N_29833);
and UO_2373 (O_2373,N_28756,N_28664);
nand UO_2374 (O_2374,N_29701,N_28543);
nand UO_2375 (O_2375,N_28851,N_29025);
nand UO_2376 (O_2376,N_29998,N_29951);
or UO_2377 (O_2377,N_28942,N_28588);
nand UO_2378 (O_2378,N_29652,N_29227);
nor UO_2379 (O_2379,N_28576,N_29857);
or UO_2380 (O_2380,N_29901,N_29990);
nor UO_2381 (O_2381,N_29226,N_28638);
nor UO_2382 (O_2382,N_28756,N_29766);
nor UO_2383 (O_2383,N_29900,N_28632);
or UO_2384 (O_2384,N_29410,N_28824);
xnor UO_2385 (O_2385,N_29772,N_28890);
and UO_2386 (O_2386,N_29354,N_29435);
and UO_2387 (O_2387,N_28712,N_29628);
or UO_2388 (O_2388,N_29007,N_28670);
and UO_2389 (O_2389,N_29342,N_28822);
xor UO_2390 (O_2390,N_29538,N_29119);
nor UO_2391 (O_2391,N_29156,N_29314);
nor UO_2392 (O_2392,N_29294,N_29046);
or UO_2393 (O_2393,N_28812,N_28769);
nor UO_2394 (O_2394,N_29932,N_29013);
nand UO_2395 (O_2395,N_29792,N_28710);
or UO_2396 (O_2396,N_28841,N_28695);
xor UO_2397 (O_2397,N_29106,N_29017);
nand UO_2398 (O_2398,N_28894,N_28896);
nor UO_2399 (O_2399,N_28517,N_29176);
xor UO_2400 (O_2400,N_29672,N_29022);
or UO_2401 (O_2401,N_29040,N_28815);
nand UO_2402 (O_2402,N_29721,N_29475);
or UO_2403 (O_2403,N_29706,N_28760);
and UO_2404 (O_2404,N_29577,N_29704);
nand UO_2405 (O_2405,N_29272,N_29255);
or UO_2406 (O_2406,N_29953,N_29519);
or UO_2407 (O_2407,N_29730,N_28799);
xnor UO_2408 (O_2408,N_29334,N_29547);
nand UO_2409 (O_2409,N_29401,N_28644);
nor UO_2410 (O_2410,N_29033,N_29208);
nor UO_2411 (O_2411,N_28649,N_29577);
nor UO_2412 (O_2412,N_29097,N_28940);
or UO_2413 (O_2413,N_29965,N_29636);
and UO_2414 (O_2414,N_29288,N_29146);
nand UO_2415 (O_2415,N_28789,N_29306);
xnor UO_2416 (O_2416,N_28961,N_28879);
and UO_2417 (O_2417,N_29998,N_29404);
nor UO_2418 (O_2418,N_28644,N_29979);
or UO_2419 (O_2419,N_28722,N_29613);
and UO_2420 (O_2420,N_29060,N_28883);
nand UO_2421 (O_2421,N_28914,N_29378);
and UO_2422 (O_2422,N_28990,N_29812);
nor UO_2423 (O_2423,N_29827,N_28715);
and UO_2424 (O_2424,N_29353,N_29634);
or UO_2425 (O_2425,N_28764,N_29867);
and UO_2426 (O_2426,N_28722,N_29511);
nand UO_2427 (O_2427,N_29100,N_28938);
xnor UO_2428 (O_2428,N_28913,N_28509);
or UO_2429 (O_2429,N_29199,N_29322);
nand UO_2430 (O_2430,N_29675,N_29805);
and UO_2431 (O_2431,N_29915,N_28937);
xor UO_2432 (O_2432,N_28812,N_29885);
nand UO_2433 (O_2433,N_28691,N_29654);
nand UO_2434 (O_2434,N_28781,N_29787);
or UO_2435 (O_2435,N_28966,N_29509);
nand UO_2436 (O_2436,N_29426,N_29378);
nand UO_2437 (O_2437,N_29478,N_29194);
or UO_2438 (O_2438,N_29039,N_29807);
or UO_2439 (O_2439,N_29200,N_28703);
nor UO_2440 (O_2440,N_29059,N_29020);
or UO_2441 (O_2441,N_29162,N_29807);
or UO_2442 (O_2442,N_29034,N_28585);
nand UO_2443 (O_2443,N_29079,N_28751);
or UO_2444 (O_2444,N_29784,N_29199);
nor UO_2445 (O_2445,N_29813,N_29722);
and UO_2446 (O_2446,N_29433,N_29185);
nand UO_2447 (O_2447,N_29888,N_28515);
or UO_2448 (O_2448,N_29357,N_29416);
and UO_2449 (O_2449,N_29612,N_29595);
xnor UO_2450 (O_2450,N_29416,N_28758);
nand UO_2451 (O_2451,N_28859,N_29857);
nand UO_2452 (O_2452,N_28770,N_29766);
nand UO_2453 (O_2453,N_29993,N_29439);
nand UO_2454 (O_2454,N_29769,N_29363);
nand UO_2455 (O_2455,N_28909,N_28698);
xnor UO_2456 (O_2456,N_28714,N_28615);
nand UO_2457 (O_2457,N_29204,N_28701);
and UO_2458 (O_2458,N_29000,N_29776);
and UO_2459 (O_2459,N_29962,N_29975);
or UO_2460 (O_2460,N_29526,N_28964);
or UO_2461 (O_2461,N_29207,N_28685);
nand UO_2462 (O_2462,N_28799,N_29204);
nand UO_2463 (O_2463,N_29397,N_28711);
or UO_2464 (O_2464,N_29936,N_29738);
nand UO_2465 (O_2465,N_28515,N_29505);
xor UO_2466 (O_2466,N_29159,N_29057);
nand UO_2467 (O_2467,N_29652,N_29249);
or UO_2468 (O_2468,N_29521,N_29884);
nor UO_2469 (O_2469,N_28753,N_29198);
nor UO_2470 (O_2470,N_29998,N_29952);
nor UO_2471 (O_2471,N_29348,N_29624);
xnor UO_2472 (O_2472,N_29547,N_29173);
or UO_2473 (O_2473,N_28524,N_29897);
or UO_2474 (O_2474,N_28594,N_29984);
nor UO_2475 (O_2475,N_28516,N_29441);
nor UO_2476 (O_2476,N_28854,N_29537);
nor UO_2477 (O_2477,N_28931,N_28614);
and UO_2478 (O_2478,N_29900,N_28996);
xnor UO_2479 (O_2479,N_28818,N_29994);
or UO_2480 (O_2480,N_29048,N_29194);
and UO_2481 (O_2481,N_29701,N_29440);
or UO_2482 (O_2482,N_28982,N_29948);
and UO_2483 (O_2483,N_29721,N_29875);
or UO_2484 (O_2484,N_28951,N_29729);
nand UO_2485 (O_2485,N_29797,N_28772);
and UO_2486 (O_2486,N_29037,N_29021);
xnor UO_2487 (O_2487,N_29971,N_29001);
nand UO_2488 (O_2488,N_28567,N_28786);
nand UO_2489 (O_2489,N_28909,N_29468);
nand UO_2490 (O_2490,N_29990,N_29734);
xnor UO_2491 (O_2491,N_29273,N_29580);
nor UO_2492 (O_2492,N_28977,N_28571);
and UO_2493 (O_2493,N_28655,N_29435);
xnor UO_2494 (O_2494,N_28979,N_28996);
nand UO_2495 (O_2495,N_29381,N_29151);
or UO_2496 (O_2496,N_29451,N_28518);
or UO_2497 (O_2497,N_29447,N_29293);
nor UO_2498 (O_2498,N_28585,N_29568);
nand UO_2499 (O_2499,N_29183,N_29915);
nand UO_2500 (O_2500,N_29121,N_29469);
and UO_2501 (O_2501,N_29570,N_28664);
and UO_2502 (O_2502,N_29950,N_29640);
or UO_2503 (O_2503,N_29081,N_29113);
xnor UO_2504 (O_2504,N_29058,N_29111);
xor UO_2505 (O_2505,N_29494,N_28682);
or UO_2506 (O_2506,N_28524,N_28641);
and UO_2507 (O_2507,N_29131,N_28594);
nand UO_2508 (O_2508,N_29593,N_28937);
nand UO_2509 (O_2509,N_28558,N_29590);
nor UO_2510 (O_2510,N_28904,N_29007);
or UO_2511 (O_2511,N_29072,N_29353);
xor UO_2512 (O_2512,N_29665,N_29654);
nand UO_2513 (O_2513,N_28658,N_28891);
and UO_2514 (O_2514,N_29841,N_29789);
xnor UO_2515 (O_2515,N_29519,N_29629);
or UO_2516 (O_2516,N_28527,N_29931);
or UO_2517 (O_2517,N_29274,N_29605);
nor UO_2518 (O_2518,N_29504,N_28663);
or UO_2519 (O_2519,N_29071,N_29114);
nor UO_2520 (O_2520,N_28786,N_28774);
and UO_2521 (O_2521,N_29039,N_29224);
and UO_2522 (O_2522,N_29560,N_29920);
or UO_2523 (O_2523,N_28594,N_29574);
xnor UO_2524 (O_2524,N_29787,N_28522);
or UO_2525 (O_2525,N_29302,N_29746);
xor UO_2526 (O_2526,N_28749,N_28868);
xor UO_2527 (O_2527,N_29930,N_29747);
nor UO_2528 (O_2528,N_29147,N_29506);
or UO_2529 (O_2529,N_29406,N_29567);
or UO_2530 (O_2530,N_29173,N_29289);
or UO_2531 (O_2531,N_29529,N_29649);
xor UO_2532 (O_2532,N_28609,N_29877);
nand UO_2533 (O_2533,N_28711,N_29202);
xnor UO_2534 (O_2534,N_28774,N_29599);
nor UO_2535 (O_2535,N_29726,N_29178);
nor UO_2536 (O_2536,N_29440,N_28700);
or UO_2537 (O_2537,N_29429,N_29656);
xnor UO_2538 (O_2538,N_28876,N_28653);
xnor UO_2539 (O_2539,N_28885,N_29975);
or UO_2540 (O_2540,N_29146,N_29948);
or UO_2541 (O_2541,N_29309,N_29269);
or UO_2542 (O_2542,N_29743,N_29208);
or UO_2543 (O_2543,N_28577,N_29672);
nor UO_2544 (O_2544,N_29320,N_29512);
nor UO_2545 (O_2545,N_29332,N_29363);
nand UO_2546 (O_2546,N_28725,N_28739);
or UO_2547 (O_2547,N_29354,N_29796);
nand UO_2548 (O_2548,N_29516,N_29564);
and UO_2549 (O_2549,N_29922,N_29258);
nor UO_2550 (O_2550,N_29818,N_29859);
and UO_2551 (O_2551,N_29924,N_29527);
xor UO_2552 (O_2552,N_28616,N_28908);
nand UO_2553 (O_2553,N_29229,N_28809);
xnor UO_2554 (O_2554,N_28747,N_28874);
nand UO_2555 (O_2555,N_29539,N_28637);
xnor UO_2556 (O_2556,N_29370,N_28750);
nand UO_2557 (O_2557,N_29833,N_29823);
nand UO_2558 (O_2558,N_28701,N_29422);
xnor UO_2559 (O_2559,N_29786,N_29713);
xnor UO_2560 (O_2560,N_29040,N_29767);
or UO_2561 (O_2561,N_28684,N_29633);
xor UO_2562 (O_2562,N_29057,N_29261);
or UO_2563 (O_2563,N_29111,N_29406);
or UO_2564 (O_2564,N_29739,N_28756);
xnor UO_2565 (O_2565,N_28962,N_29440);
xnor UO_2566 (O_2566,N_29306,N_29289);
xnor UO_2567 (O_2567,N_28871,N_29345);
nor UO_2568 (O_2568,N_28852,N_29165);
nor UO_2569 (O_2569,N_29461,N_28600);
and UO_2570 (O_2570,N_29138,N_28958);
xnor UO_2571 (O_2571,N_29414,N_28965);
or UO_2572 (O_2572,N_29038,N_29229);
nand UO_2573 (O_2573,N_29223,N_29386);
and UO_2574 (O_2574,N_28939,N_29556);
or UO_2575 (O_2575,N_29528,N_29290);
xnor UO_2576 (O_2576,N_29859,N_29847);
nand UO_2577 (O_2577,N_29809,N_28809);
nor UO_2578 (O_2578,N_29937,N_29720);
xor UO_2579 (O_2579,N_29611,N_29319);
or UO_2580 (O_2580,N_28823,N_29939);
and UO_2581 (O_2581,N_28901,N_29515);
nand UO_2582 (O_2582,N_28518,N_28753);
and UO_2583 (O_2583,N_29337,N_28947);
or UO_2584 (O_2584,N_29908,N_29064);
xnor UO_2585 (O_2585,N_29795,N_29454);
or UO_2586 (O_2586,N_29606,N_28955);
or UO_2587 (O_2587,N_29471,N_29446);
xnor UO_2588 (O_2588,N_29537,N_29428);
xor UO_2589 (O_2589,N_29996,N_29439);
nor UO_2590 (O_2590,N_28542,N_29870);
xor UO_2591 (O_2591,N_28501,N_29819);
nor UO_2592 (O_2592,N_28535,N_29932);
nor UO_2593 (O_2593,N_29939,N_28664);
nand UO_2594 (O_2594,N_28695,N_29465);
nor UO_2595 (O_2595,N_29186,N_29369);
xnor UO_2596 (O_2596,N_29525,N_29103);
and UO_2597 (O_2597,N_29952,N_29237);
nor UO_2598 (O_2598,N_29155,N_29531);
xor UO_2599 (O_2599,N_29342,N_29679);
or UO_2600 (O_2600,N_28723,N_29948);
and UO_2601 (O_2601,N_29185,N_28652);
nand UO_2602 (O_2602,N_29803,N_28518);
or UO_2603 (O_2603,N_29476,N_28761);
and UO_2604 (O_2604,N_28852,N_29061);
or UO_2605 (O_2605,N_29739,N_29803);
nand UO_2606 (O_2606,N_28547,N_29408);
xor UO_2607 (O_2607,N_29516,N_29659);
nor UO_2608 (O_2608,N_29496,N_29146);
and UO_2609 (O_2609,N_29408,N_29110);
xor UO_2610 (O_2610,N_29170,N_29660);
or UO_2611 (O_2611,N_29582,N_29800);
nand UO_2612 (O_2612,N_29692,N_29828);
nor UO_2613 (O_2613,N_29248,N_28672);
nor UO_2614 (O_2614,N_28886,N_29375);
and UO_2615 (O_2615,N_28874,N_29985);
and UO_2616 (O_2616,N_29521,N_29244);
nor UO_2617 (O_2617,N_29169,N_28972);
and UO_2618 (O_2618,N_29779,N_29967);
and UO_2619 (O_2619,N_28860,N_29192);
or UO_2620 (O_2620,N_29331,N_29035);
or UO_2621 (O_2621,N_29122,N_29532);
and UO_2622 (O_2622,N_28516,N_29500);
nor UO_2623 (O_2623,N_29027,N_29246);
xnor UO_2624 (O_2624,N_29375,N_29957);
and UO_2625 (O_2625,N_28651,N_29825);
xor UO_2626 (O_2626,N_29473,N_28887);
and UO_2627 (O_2627,N_29080,N_29932);
and UO_2628 (O_2628,N_28509,N_29792);
nor UO_2629 (O_2629,N_29246,N_28571);
nor UO_2630 (O_2630,N_28748,N_29784);
xnor UO_2631 (O_2631,N_29481,N_28650);
nor UO_2632 (O_2632,N_29155,N_29757);
and UO_2633 (O_2633,N_29307,N_29398);
and UO_2634 (O_2634,N_29516,N_28505);
or UO_2635 (O_2635,N_29493,N_29926);
nor UO_2636 (O_2636,N_29190,N_28966);
nand UO_2637 (O_2637,N_28875,N_28781);
nand UO_2638 (O_2638,N_29310,N_28553);
nand UO_2639 (O_2639,N_28565,N_29877);
xnor UO_2640 (O_2640,N_29733,N_28967);
nor UO_2641 (O_2641,N_28803,N_29072);
and UO_2642 (O_2642,N_28980,N_29668);
nand UO_2643 (O_2643,N_29793,N_28682);
or UO_2644 (O_2644,N_29299,N_28606);
or UO_2645 (O_2645,N_29555,N_28776);
nor UO_2646 (O_2646,N_29283,N_28681);
or UO_2647 (O_2647,N_28972,N_28646);
nand UO_2648 (O_2648,N_29821,N_29250);
or UO_2649 (O_2649,N_29045,N_28693);
and UO_2650 (O_2650,N_29736,N_29527);
nor UO_2651 (O_2651,N_29910,N_29366);
xor UO_2652 (O_2652,N_29339,N_29946);
nor UO_2653 (O_2653,N_29335,N_28543);
nand UO_2654 (O_2654,N_29338,N_29180);
or UO_2655 (O_2655,N_29587,N_29543);
nor UO_2656 (O_2656,N_29663,N_29562);
nand UO_2657 (O_2657,N_29271,N_29113);
nand UO_2658 (O_2658,N_29075,N_28889);
or UO_2659 (O_2659,N_29681,N_29428);
nand UO_2660 (O_2660,N_29937,N_29438);
and UO_2661 (O_2661,N_29807,N_28580);
xor UO_2662 (O_2662,N_29840,N_29114);
and UO_2663 (O_2663,N_29715,N_29954);
nand UO_2664 (O_2664,N_29214,N_28951);
nor UO_2665 (O_2665,N_29482,N_29541);
nor UO_2666 (O_2666,N_29608,N_28572);
nor UO_2667 (O_2667,N_28848,N_29223);
and UO_2668 (O_2668,N_29322,N_29790);
and UO_2669 (O_2669,N_28511,N_28907);
or UO_2670 (O_2670,N_29502,N_29930);
and UO_2671 (O_2671,N_29980,N_29549);
xor UO_2672 (O_2672,N_29286,N_29366);
xnor UO_2673 (O_2673,N_29178,N_28758);
nor UO_2674 (O_2674,N_28592,N_28992);
and UO_2675 (O_2675,N_29602,N_29343);
xnor UO_2676 (O_2676,N_28804,N_28681);
xor UO_2677 (O_2677,N_29247,N_29600);
and UO_2678 (O_2678,N_28638,N_29381);
nor UO_2679 (O_2679,N_28536,N_29117);
nor UO_2680 (O_2680,N_29926,N_29733);
nor UO_2681 (O_2681,N_29681,N_29583);
nand UO_2682 (O_2682,N_29745,N_29248);
nor UO_2683 (O_2683,N_29795,N_28576);
or UO_2684 (O_2684,N_28574,N_29384);
nor UO_2685 (O_2685,N_28881,N_28698);
xnor UO_2686 (O_2686,N_29456,N_29156);
or UO_2687 (O_2687,N_29556,N_28543);
and UO_2688 (O_2688,N_28771,N_28616);
nand UO_2689 (O_2689,N_29509,N_29122);
xor UO_2690 (O_2690,N_29279,N_29425);
and UO_2691 (O_2691,N_29759,N_29399);
or UO_2692 (O_2692,N_28507,N_29240);
xor UO_2693 (O_2693,N_29933,N_29932);
and UO_2694 (O_2694,N_29163,N_28722);
nor UO_2695 (O_2695,N_28774,N_28969);
or UO_2696 (O_2696,N_28950,N_29009);
or UO_2697 (O_2697,N_29504,N_29788);
and UO_2698 (O_2698,N_28739,N_29459);
nor UO_2699 (O_2699,N_29016,N_29165);
nor UO_2700 (O_2700,N_29152,N_28730);
nor UO_2701 (O_2701,N_29105,N_28837);
nor UO_2702 (O_2702,N_29879,N_29462);
or UO_2703 (O_2703,N_28989,N_29578);
nor UO_2704 (O_2704,N_29373,N_28978);
nand UO_2705 (O_2705,N_29620,N_29075);
or UO_2706 (O_2706,N_29809,N_29338);
or UO_2707 (O_2707,N_29342,N_28884);
and UO_2708 (O_2708,N_28665,N_29572);
and UO_2709 (O_2709,N_28820,N_29189);
nor UO_2710 (O_2710,N_29392,N_29154);
nor UO_2711 (O_2711,N_28851,N_29106);
or UO_2712 (O_2712,N_29309,N_28896);
nor UO_2713 (O_2713,N_29448,N_29911);
and UO_2714 (O_2714,N_29924,N_28916);
xnor UO_2715 (O_2715,N_28549,N_29123);
or UO_2716 (O_2716,N_28574,N_29477);
nand UO_2717 (O_2717,N_29454,N_29487);
xor UO_2718 (O_2718,N_29492,N_29397);
and UO_2719 (O_2719,N_29375,N_29840);
nor UO_2720 (O_2720,N_29163,N_29510);
and UO_2721 (O_2721,N_29964,N_29020);
nor UO_2722 (O_2722,N_29723,N_29979);
and UO_2723 (O_2723,N_29914,N_29629);
and UO_2724 (O_2724,N_29869,N_28802);
or UO_2725 (O_2725,N_29320,N_28869);
and UO_2726 (O_2726,N_29099,N_28702);
or UO_2727 (O_2727,N_28834,N_28643);
nor UO_2728 (O_2728,N_29635,N_28769);
xnor UO_2729 (O_2729,N_28667,N_29401);
nor UO_2730 (O_2730,N_29832,N_28944);
nand UO_2731 (O_2731,N_29961,N_29124);
nor UO_2732 (O_2732,N_29661,N_29834);
nand UO_2733 (O_2733,N_29303,N_28708);
and UO_2734 (O_2734,N_28695,N_29742);
or UO_2735 (O_2735,N_28652,N_28734);
or UO_2736 (O_2736,N_29775,N_29830);
or UO_2737 (O_2737,N_29766,N_29032);
and UO_2738 (O_2738,N_28647,N_29332);
nor UO_2739 (O_2739,N_28668,N_28540);
xor UO_2740 (O_2740,N_29389,N_29473);
xor UO_2741 (O_2741,N_28959,N_28591);
xor UO_2742 (O_2742,N_29551,N_29863);
nor UO_2743 (O_2743,N_29831,N_28754);
nor UO_2744 (O_2744,N_29620,N_28740);
nor UO_2745 (O_2745,N_29594,N_28500);
nand UO_2746 (O_2746,N_29556,N_29434);
or UO_2747 (O_2747,N_29387,N_29891);
or UO_2748 (O_2748,N_29021,N_29171);
nand UO_2749 (O_2749,N_29587,N_29502);
or UO_2750 (O_2750,N_28837,N_29224);
xor UO_2751 (O_2751,N_29400,N_28708);
xnor UO_2752 (O_2752,N_28980,N_29247);
xor UO_2753 (O_2753,N_28654,N_29440);
nand UO_2754 (O_2754,N_29417,N_28944);
and UO_2755 (O_2755,N_28921,N_29745);
nor UO_2756 (O_2756,N_29699,N_28779);
xor UO_2757 (O_2757,N_29368,N_29776);
and UO_2758 (O_2758,N_28755,N_29529);
and UO_2759 (O_2759,N_29464,N_29317);
nor UO_2760 (O_2760,N_29192,N_29476);
nor UO_2761 (O_2761,N_29111,N_28907);
and UO_2762 (O_2762,N_29412,N_29878);
or UO_2763 (O_2763,N_28880,N_29005);
nor UO_2764 (O_2764,N_28520,N_28843);
nor UO_2765 (O_2765,N_29206,N_29533);
and UO_2766 (O_2766,N_29036,N_28974);
xnor UO_2767 (O_2767,N_28883,N_29839);
nor UO_2768 (O_2768,N_29555,N_29734);
nor UO_2769 (O_2769,N_29583,N_28863);
or UO_2770 (O_2770,N_28770,N_28718);
or UO_2771 (O_2771,N_29547,N_29992);
nor UO_2772 (O_2772,N_29243,N_29025);
or UO_2773 (O_2773,N_29163,N_28628);
or UO_2774 (O_2774,N_29399,N_29623);
nor UO_2775 (O_2775,N_29907,N_28924);
and UO_2776 (O_2776,N_28882,N_29153);
nand UO_2777 (O_2777,N_29712,N_28780);
and UO_2778 (O_2778,N_28845,N_28690);
nor UO_2779 (O_2779,N_28860,N_29389);
nor UO_2780 (O_2780,N_29853,N_29995);
or UO_2781 (O_2781,N_28581,N_29716);
nor UO_2782 (O_2782,N_29003,N_29382);
nor UO_2783 (O_2783,N_28700,N_29892);
nand UO_2784 (O_2784,N_29054,N_29782);
nor UO_2785 (O_2785,N_29672,N_29383);
xnor UO_2786 (O_2786,N_29955,N_28766);
xnor UO_2787 (O_2787,N_29848,N_29226);
or UO_2788 (O_2788,N_29812,N_28773);
nor UO_2789 (O_2789,N_29428,N_28666);
nand UO_2790 (O_2790,N_29020,N_28942);
or UO_2791 (O_2791,N_28933,N_29143);
and UO_2792 (O_2792,N_29461,N_29190);
nand UO_2793 (O_2793,N_28816,N_29892);
xnor UO_2794 (O_2794,N_28677,N_29449);
nand UO_2795 (O_2795,N_29346,N_28827);
nor UO_2796 (O_2796,N_29700,N_29990);
xor UO_2797 (O_2797,N_28816,N_28694);
and UO_2798 (O_2798,N_29697,N_28859);
xnor UO_2799 (O_2799,N_29127,N_28552);
and UO_2800 (O_2800,N_28979,N_29070);
or UO_2801 (O_2801,N_29646,N_29742);
xnor UO_2802 (O_2802,N_29810,N_29750);
or UO_2803 (O_2803,N_28797,N_29619);
xnor UO_2804 (O_2804,N_29290,N_28754);
or UO_2805 (O_2805,N_28941,N_29368);
or UO_2806 (O_2806,N_29181,N_29065);
and UO_2807 (O_2807,N_28589,N_29848);
and UO_2808 (O_2808,N_29511,N_28979);
or UO_2809 (O_2809,N_28545,N_29076);
and UO_2810 (O_2810,N_29850,N_29753);
xor UO_2811 (O_2811,N_29378,N_28648);
and UO_2812 (O_2812,N_29853,N_29554);
nor UO_2813 (O_2813,N_29461,N_29004);
nor UO_2814 (O_2814,N_29184,N_28945);
xor UO_2815 (O_2815,N_29573,N_29073);
and UO_2816 (O_2816,N_29512,N_29178);
nand UO_2817 (O_2817,N_28982,N_28570);
and UO_2818 (O_2818,N_29838,N_28855);
nor UO_2819 (O_2819,N_29651,N_28522);
xnor UO_2820 (O_2820,N_29589,N_28610);
nand UO_2821 (O_2821,N_28747,N_29172);
and UO_2822 (O_2822,N_29922,N_28533);
nor UO_2823 (O_2823,N_29878,N_28870);
and UO_2824 (O_2824,N_29480,N_28603);
and UO_2825 (O_2825,N_29163,N_28910);
xnor UO_2826 (O_2826,N_28656,N_28586);
and UO_2827 (O_2827,N_29575,N_29959);
nand UO_2828 (O_2828,N_29400,N_28776);
or UO_2829 (O_2829,N_29560,N_28655);
xor UO_2830 (O_2830,N_29452,N_29824);
and UO_2831 (O_2831,N_29550,N_29422);
or UO_2832 (O_2832,N_29818,N_28898);
or UO_2833 (O_2833,N_28664,N_29277);
and UO_2834 (O_2834,N_28807,N_29084);
nand UO_2835 (O_2835,N_28600,N_29523);
nand UO_2836 (O_2836,N_29643,N_28985);
xnor UO_2837 (O_2837,N_29069,N_28558);
nand UO_2838 (O_2838,N_28783,N_28502);
nor UO_2839 (O_2839,N_29645,N_29793);
or UO_2840 (O_2840,N_29494,N_28585);
nand UO_2841 (O_2841,N_29363,N_28578);
or UO_2842 (O_2842,N_29997,N_29233);
xor UO_2843 (O_2843,N_28651,N_29756);
or UO_2844 (O_2844,N_28520,N_29117);
nand UO_2845 (O_2845,N_29073,N_29820);
nand UO_2846 (O_2846,N_29994,N_29240);
nor UO_2847 (O_2847,N_28552,N_29576);
or UO_2848 (O_2848,N_29206,N_29779);
nand UO_2849 (O_2849,N_28685,N_28525);
xnor UO_2850 (O_2850,N_29408,N_28901);
xor UO_2851 (O_2851,N_28565,N_29609);
and UO_2852 (O_2852,N_29947,N_28812);
xor UO_2853 (O_2853,N_28923,N_29545);
nand UO_2854 (O_2854,N_29161,N_29219);
nand UO_2855 (O_2855,N_29984,N_28956);
nand UO_2856 (O_2856,N_29803,N_28531);
nor UO_2857 (O_2857,N_29801,N_29103);
or UO_2858 (O_2858,N_28801,N_29694);
nand UO_2859 (O_2859,N_29623,N_29034);
nor UO_2860 (O_2860,N_29101,N_29344);
and UO_2861 (O_2861,N_29361,N_29383);
or UO_2862 (O_2862,N_29367,N_28641);
or UO_2863 (O_2863,N_28951,N_29841);
xnor UO_2864 (O_2864,N_28871,N_29907);
nand UO_2865 (O_2865,N_29181,N_29024);
or UO_2866 (O_2866,N_29230,N_29403);
or UO_2867 (O_2867,N_28570,N_29391);
or UO_2868 (O_2868,N_28505,N_28730);
or UO_2869 (O_2869,N_29800,N_28967);
nand UO_2870 (O_2870,N_29347,N_29034);
nand UO_2871 (O_2871,N_29600,N_28945);
and UO_2872 (O_2872,N_29315,N_28999);
and UO_2873 (O_2873,N_28714,N_28798);
and UO_2874 (O_2874,N_29291,N_28857);
nand UO_2875 (O_2875,N_28698,N_29212);
or UO_2876 (O_2876,N_29545,N_29648);
xor UO_2877 (O_2877,N_29922,N_28878);
or UO_2878 (O_2878,N_29799,N_28970);
xnor UO_2879 (O_2879,N_29452,N_29968);
or UO_2880 (O_2880,N_28661,N_29425);
and UO_2881 (O_2881,N_29470,N_29341);
nor UO_2882 (O_2882,N_29959,N_29265);
xnor UO_2883 (O_2883,N_29064,N_28915);
nor UO_2884 (O_2884,N_29907,N_29758);
or UO_2885 (O_2885,N_29568,N_28966);
xor UO_2886 (O_2886,N_29593,N_29809);
xor UO_2887 (O_2887,N_29517,N_28653);
and UO_2888 (O_2888,N_28873,N_29928);
nor UO_2889 (O_2889,N_28831,N_29917);
nand UO_2890 (O_2890,N_29712,N_29005);
nand UO_2891 (O_2891,N_29193,N_28680);
xor UO_2892 (O_2892,N_29313,N_29020);
or UO_2893 (O_2893,N_28793,N_28849);
and UO_2894 (O_2894,N_29516,N_29243);
nand UO_2895 (O_2895,N_29068,N_28753);
nor UO_2896 (O_2896,N_28714,N_29403);
nor UO_2897 (O_2897,N_28876,N_28837);
and UO_2898 (O_2898,N_28650,N_29007);
nor UO_2899 (O_2899,N_29868,N_29244);
or UO_2900 (O_2900,N_29804,N_29765);
and UO_2901 (O_2901,N_29264,N_29717);
nand UO_2902 (O_2902,N_29839,N_28921);
xor UO_2903 (O_2903,N_29629,N_29689);
or UO_2904 (O_2904,N_28752,N_28918);
xor UO_2905 (O_2905,N_29653,N_29015);
or UO_2906 (O_2906,N_28807,N_29485);
and UO_2907 (O_2907,N_28661,N_28891);
nand UO_2908 (O_2908,N_29443,N_29238);
nand UO_2909 (O_2909,N_28524,N_28712);
xnor UO_2910 (O_2910,N_29358,N_29400);
xnor UO_2911 (O_2911,N_29764,N_28504);
and UO_2912 (O_2912,N_29886,N_29154);
or UO_2913 (O_2913,N_29675,N_29784);
or UO_2914 (O_2914,N_29174,N_28897);
xnor UO_2915 (O_2915,N_29137,N_28610);
nor UO_2916 (O_2916,N_29309,N_28940);
and UO_2917 (O_2917,N_29045,N_29988);
or UO_2918 (O_2918,N_29609,N_29555);
nor UO_2919 (O_2919,N_29323,N_29808);
nand UO_2920 (O_2920,N_29778,N_29759);
nand UO_2921 (O_2921,N_29940,N_29088);
or UO_2922 (O_2922,N_28910,N_28925);
xnor UO_2923 (O_2923,N_28911,N_29431);
xor UO_2924 (O_2924,N_28562,N_29508);
nand UO_2925 (O_2925,N_29277,N_28843);
xor UO_2926 (O_2926,N_29451,N_29094);
and UO_2927 (O_2927,N_29039,N_28784);
and UO_2928 (O_2928,N_29295,N_28742);
nor UO_2929 (O_2929,N_29818,N_28884);
xor UO_2930 (O_2930,N_29059,N_28661);
nor UO_2931 (O_2931,N_29880,N_29695);
or UO_2932 (O_2932,N_29603,N_28664);
or UO_2933 (O_2933,N_29265,N_29313);
nand UO_2934 (O_2934,N_28777,N_29140);
or UO_2935 (O_2935,N_29912,N_29613);
xor UO_2936 (O_2936,N_29484,N_28693);
and UO_2937 (O_2937,N_29217,N_29914);
or UO_2938 (O_2938,N_29118,N_29307);
and UO_2939 (O_2939,N_28586,N_29040);
nand UO_2940 (O_2940,N_29380,N_29232);
xnor UO_2941 (O_2941,N_28562,N_29933);
nor UO_2942 (O_2942,N_29021,N_29185);
nand UO_2943 (O_2943,N_29667,N_28740);
or UO_2944 (O_2944,N_29773,N_28959);
nor UO_2945 (O_2945,N_29818,N_29806);
xor UO_2946 (O_2946,N_29854,N_29107);
and UO_2947 (O_2947,N_29527,N_28860);
and UO_2948 (O_2948,N_29459,N_29564);
nor UO_2949 (O_2949,N_29203,N_28975);
nor UO_2950 (O_2950,N_28848,N_28920);
xor UO_2951 (O_2951,N_28823,N_28611);
and UO_2952 (O_2952,N_29860,N_28978);
nor UO_2953 (O_2953,N_29212,N_29161);
or UO_2954 (O_2954,N_29045,N_29544);
xor UO_2955 (O_2955,N_29568,N_29490);
or UO_2956 (O_2956,N_29025,N_28634);
or UO_2957 (O_2957,N_29075,N_29061);
and UO_2958 (O_2958,N_29176,N_29906);
and UO_2959 (O_2959,N_29966,N_28881);
nor UO_2960 (O_2960,N_29595,N_28577);
and UO_2961 (O_2961,N_29438,N_29806);
xnor UO_2962 (O_2962,N_28527,N_29319);
or UO_2963 (O_2963,N_29506,N_29113);
and UO_2964 (O_2964,N_29478,N_28625);
nor UO_2965 (O_2965,N_29797,N_29033);
nor UO_2966 (O_2966,N_29309,N_28857);
and UO_2967 (O_2967,N_29015,N_29287);
or UO_2968 (O_2968,N_29793,N_29106);
nand UO_2969 (O_2969,N_29771,N_29350);
xnor UO_2970 (O_2970,N_29613,N_28995);
and UO_2971 (O_2971,N_28786,N_29153);
or UO_2972 (O_2972,N_29629,N_29733);
xnor UO_2973 (O_2973,N_28921,N_29768);
nor UO_2974 (O_2974,N_29321,N_29021);
nor UO_2975 (O_2975,N_28582,N_29768);
and UO_2976 (O_2976,N_29990,N_29438);
nand UO_2977 (O_2977,N_28753,N_28547);
nand UO_2978 (O_2978,N_29733,N_29491);
or UO_2979 (O_2979,N_29947,N_28515);
nor UO_2980 (O_2980,N_28734,N_28638);
and UO_2981 (O_2981,N_28855,N_29527);
and UO_2982 (O_2982,N_28808,N_29587);
and UO_2983 (O_2983,N_29396,N_29902);
or UO_2984 (O_2984,N_29079,N_29440);
nand UO_2985 (O_2985,N_28545,N_28861);
and UO_2986 (O_2986,N_29160,N_28734);
nand UO_2987 (O_2987,N_28764,N_29840);
and UO_2988 (O_2988,N_29007,N_29739);
or UO_2989 (O_2989,N_29896,N_29613);
nand UO_2990 (O_2990,N_29089,N_29334);
nand UO_2991 (O_2991,N_29546,N_28833);
or UO_2992 (O_2992,N_28916,N_29234);
or UO_2993 (O_2993,N_28601,N_28760);
and UO_2994 (O_2994,N_29835,N_29243);
nor UO_2995 (O_2995,N_29022,N_29890);
nand UO_2996 (O_2996,N_29485,N_29158);
xor UO_2997 (O_2997,N_29901,N_29861);
xor UO_2998 (O_2998,N_29091,N_29013);
or UO_2999 (O_2999,N_29682,N_29241);
or UO_3000 (O_3000,N_29164,N_28996);
or UO_3001 (O_3001,N_29805,N_29711);
and UO_3002 (O_3002,N_29568,N_28997);
and UO_3003 (O_3003,N_29948,N_29619);
nor UO_3004 (O_3004,N_29374,N_29564);
nand UO_3005 (O_3005,N_28560,N_28639);
nor UO_3006 (O_3006,N_28919,N_28627);
xnor UO_3007 (O_3007,N_29322,N_28695);
and UO_3008 (O_3008,N_29454,N_29689);
xnor UO_3009 (O_3009,N_29003,N_29525);
or UO_3010 (O_3010,N_29138,N_28875);
or UO_3011 (O_3011,N_29562,N_29919);
nand UO_3012 (O_3012,N_28527,N_28616);
or UO_3013 (O_3013,N_28803,N_29101);
nor UO_3014 (O_3014,N_28796,N_28799);
or UO_3015 (O_3015,N_28531,N_28911);
xnor UO_3016 (O_3016,N_29003,N_29807);
nor UO_3017 (O_3017,N_29058,N_29704);
or UO_3018 (O_3018,N_29034,N_29065);
and UO_3019 (O_3019,N_29488,N_29235);
nor UO_3020 (O_3020,N_28742,N_28729);
nand UO_3021 (O_3021,N_29082,N_28645);
nor UO_3022 (O_3022,N_29312,N_28521);
and UO_3023 (O_3023,N_29680,N_29879);
and UO_3024 (O_3024,N_29849,N_29917);
nand UO_3025 (O_3025,N_28856,N_28773);
and UO_3026 (O_3026,N_29843,N_29770);
and UO_3027 (O_3027,N_29146,N_29147);
nand UO_3028 (O_3028,N_29588,N_29353);
nor UO_3029 (O_3029,N_28954,N_28655);
nor UO_3030 (O_3030,N_29590,N_29172);
or UO_3031 (O_3031,N_29675,N_28585);
and UO_3032 (O_3032,N_29538,N_28782);
or UO_3033 (O_3033,N_29699,N_29200);
nand UO_3034 (O_3034,N_28602,N_29159);
nor UO_3035 (O_3035,N_29142,N_28774);
nor UO_3036 (O_3036,N_28701,N_28822);
nor UO_3037 (O_3037,N_28557,N_28881);
nand UO_3038 (O_3038,N_28760,N_29315);
nand UO_3039 (O_3039,N_28617,N_28513);
xnor UO_3040 (O_3040,N_29194,N_29848);
nor UO_3041 (O_3041,N_29511,N_29756);
nor UO_3042 (O_3042,N_29845,N_28771);
xor UO_3043 (O_3043,N_29410,N_29877);
or UO_3044 (O_3044,N_28511,N_28847);
or UO_3045 (O_3045,N_29413,N_28997);
nor UO_3046 (O_3046,N_29064,N_28652);
nor UO_3047 (O_3047,N_29909,N_29767);
nand UO_3048 (O_3048,N_29831,N_29574);
xnor UO_3049 (O_3049,N_28849,N_29037);
nand UO_3050 (O_3050,N_29376,N_29781);
or UO_3051 (O_3051,N_28797,N_28796);
nand UO_3052 (O_3052,N_29220,N_29305);
nor UO_3053 (O_3053,N_28690,N_29022);
and UO_3054 (O_3054,N_29048,N_29108);
nor UO_3055 (O_3055,N_29432,N_29728);
nor UO_3056 (O_3056,N_29372,N_29546);
nand UO_3057 (O_3057,N_28547,N_29003);
nand UO_3058 (O_3058,N_29726,N_29088);
and UO_3059 (O_3059,N_29060,N_29896);
and UO_3060 (O_3060,N_28548,N_29078);
and UO_3061 (O_3061,N_29064,N_29435);
nand UO_3062 (O_3062,N_29883,N_29205);
nor UO_3063 (O_3063,N_28817,N_29733);
nor UO_3064 (O_3064,N_29907,N_28948);
nand UO_3065 (O_3065,N_29812,N_28961);
and UO_3066 (O_3066,N_28997,N_29033);
xnor UO_3067 (O_3067,N_29735,N_28896);
and UO_3068 (O_3068,N_29853,N_29584);
and UO_3069 (O_3069,N_29503,N_29869);
nand UO_3070 (O_3070,N_29640,N_29904);
or UO_3071 (O_3071,N_29624,N_29874);
or UO_3072 (O_3072,N_28910,N_28761);
nor UO_3073 (O_3073,N_29685,N_29590);
nor UO_3074 (O_3074,N_29160,N_29769);
xor UO_3075 (O_3075,N_29803,N_28797);
xor UO_3076 (O_3076,N_28625,N_29378);
xnor UO_3077 (O_3077,N_29995,N_29366);
nor UO_3078 (O_3078,N_29171,N_29776);
xor UO_3079 (O_3079,N_29170,N_28798);
xnor UO_3080 (O_3080,N_28579,N_29549);
nor UO_3081 (O_3081,N_29980,N_29355);
nor UO_3082 (O_3082,N_29290,N_29856);
or UO_3083 (O_3083,N_28504,N_29679);
and UO_3084 (O_3084,N_28993,N_29896);
and UO_3085 (O_3085,N_28961,N_29969);
or UO_3086 (O_3086,N_29926,N_28722);
nand UO_3087 (O_3087,N_29153,N_29716);
or UO_3088 (O_3088,N_29541,N_29169);
xnor UO_3089 (O_3089,N_29695,N_28891);
nand UO_3090 (O_3090,N_28572,N_28793);
nand UO_3091 (O_3091,N_28771,N_29695);
nor UO_3092 (O_3092,N_29755,N_29080);
xor UO_3093 (O_3093,N_29266,N_29965);
and UO_3094 (O_3094,N_28549,N_29753);
xnor UO_3095 (O_3095,N_29919,N_29321);
and UO_3096 (O_3096,N_28661,N_28841);
xor UO_3097 (O_3097,N_29213,N_29933);
nand UO_3098 (O_3098,N_29134,N_29292);
or UO_3099 (O_3099,N_28999,N_29850);
or UO_3100 (O_3100,N_29201,N_29263);
nor UO_3101 (O_3101,N_28702,N_29799);
nor UO_3102 (O_3102,N_29332,N_29059);
nor UO_3103 (O_3103,N_29996,N_29579);
nor UO_3104 (O_3104,N_29077,N_29201);
nor UO_3105 (O_3105,N_29900,N_29160);
or UO_3106 (O_3106,N_29769,N_29862);
nor UO_3107 (O_3107,N_29183,N_29113);
and UO_3108 (O_3108,N_29949,N_28900);
nor UO_3109 (O_3109,N_29335,N_29952);
and UO_3110 (O_3110,N_29854,N_28535);
nor UO_3111 (O_3111,N_29751,N_29515);
xnor UO_3112 (O_3112,N_28930,N_29238);
and UO_3113 (O_3113,N_29576,N_29578);
nor UO_3114 (O_3114,N_29448,N_29651);
nand UO_3115 (O_3115,N_28792,N_29536);
or UO_3116 (O_3116,N_29576,N_29348);
nand UO_3117 (O_3117,N_29848,N_29498);
and UO_3118 (O_3118,N_29845,N_29042);
xnor UO_3119 (O_3119,N_28589,N_29963);
nand UO_3120 (O_3120,N_28830,N_29849);
nand UO_3121 (O_3121,N_29872,N_29664);
xor UO_3122 (O_3122,N_29376,N_29142);
nand UO_3123 (O_3123,N_29312,N_29185);
xnor UO_3124 (O_3124,N_28876,N_29532);
or UO_3125 (O_3125,N_28767,N_29054);
xor UO_3126 (O_3126,N_28514,N_28503);
nand UO_3127 (O_3127,N_28518,N_28542);
and UO_3128 (O_3128,N_29696,N_29827);
and UO_3129 (O_3129,N_29554,N_29616);
xor UO_3130 (O_3130,N_29237,N_29473);
xnor UO_3131 (O_3131,N_29824,N_28967);
xor UO_3132 (O_3132,N_28909,N_29607);
nand UO_3133 (O_3133,N_29829,N_29834);
nand UO_3134 (O_3134,N_28658,N_29717);
nor UO_3135 (O_3135,N_29742,N_29542);
xor UO_3136 (O_3136,N_28606,N_29273);
nand UO_3137 (O_3137,N_29923,N_28647);
and UO_3138 (O_3138,N_29019,N_28620);
or UO_3139 (O_3139,N_29367,N_29202);
xor UO_3140 (O_3140,N_28640,N_28596);
or UO_3141 (O_3141,N_29824,N_29772);
or UO_3142 (O_3142,N_28864,N_29120);
and UO_3143 (O_3143,N_28629,N_29593);
nor UO_3144 (O_3144,N_29556,N_29508);
nand UO_3145 (O_3145,N_29051,N_29195);
and UO_3146 (O_3146,N_28793,N_28870);
nor UO_3147 (O_3147,N_29317,N_29078);
nand UO_3148 (O_3148,N_29845,N_29816);
or UO_3149 (O_3149,N_29720,N_29873);
or UO_3150 (O_3150,N_29447,N_29276);
nor UO_3151 (O_3151,N_29780,N_29419);
and UO_3152 (O_3152,N_29046,N_28601);
nor UO_3153 (O_3153,N_29366,N_29308);
nor UO_3154 (O_3154,N_29431,N_29180);
or UO_3155 (O_3155,N_28554,N_29831);
nand UO_3156 (O_3156,N_28755,N_29758);
nand UO_3157 (O_3157,N_29230,N_28682);
nor UO_3158 (O_3158,N_29233,N_29207);
and UO_3159 (O_3159,N_29084,N_28950);
nand UO_3160 (O_3160,N_28595,N_29980);
xor UO_3161 (O_3161,N_29208,N_29552);
or UO_3162 (O_3162,N_29150,N_28610);
xnor UO_3163 (O_3163,N_29977,N_28724);
xor UO_3164 (O_3164,N_29397,N_29422);
nand UO_3165 (O_3165,N_29182,N_29967);
and UO_3166 (O_3166,N_28736,N_28977);
and UO_3167 (O_3167,N_28511,N_28879);
nand UO_3168 (O_3168,N_28580,N_29820);
nor UO_3169 (O_3169,N_29806,N_29187);
xor UO_3170 (O_3170,N_29207,N_29942);
nand UO_3171 (O_3171,N_29586,N_28616);
nor UO_3172 (O_3172,N_28667,N_29232);
nand UO_3173 (O_3173,N_29127,N_29789);
nor UO_3174 (O_3174,N_28617,N_29780);
or UO_3175 (O_3175,N_28776,N_29169);
nor UO_3176 (O_3176,N_29457,N_28921);
nand UO_3177 (O_3177,N_29732,N_28536);
and UO_3178 (O_3178,N_29244,N_29836);
xor UO_3179 (O_3179,N_29593,N_28672);
nand UO_3180 (O_3180,N_28708,N_28598);
or UO_3181 (O_3181,N_28889,N_29884);
and UO_3182 (O_3182,N_29216,N_29263);
and UO_3183 (O_3183,N_29318,N_29904);
and UO_3184 (O_3184,N_29385,N_29422);
or UO_3185 (O_3185,N_29362,N_29649);
and UO_3186 (O_3186,N_29533,N_29870);
xnor UO_3187 (O_3187,N_28604,N_29354);
or UO_3188 (O_3188,N_28659,N_29264);
and UO_3189 (O_3189,N_28653,N_28877);
nor UO_3190 (O_3190,N_29158,N_29063);
or UO_3191 (O_3191,N_29607,N_29469);
or UO_3192 (O_3192,N_29382,N_29027);
nor UO_3193 (O_3193,N_29359,N_29869);
or UO_3194 (O_3194,N_29266,N_29804);
or UO_3195 (O_3195,N_28986,N_29870);
nand UO_3196 (O_3196,N_29980,N_28815);
xor UO_3197 (O_3197,N_29911,N_28880);
and UO_3198 (O_3198,N_29755,N_29877);
xor UO_3199 (O_3199,N_28717,N_28562);
nand UO_3200 (O_3200,N_29309,N_29022);
nand UO_3201 (O_3201,N_28960,N_29948);
or UO_3202 (O_3202,N_29893,N_28723);
xor UO_3203 (O_3203,N_29683,N_28517);
nor UO_3204 (O_3204,N_28863,N_29206);
nor UO_3205 (O_3205,N_29381,N_29069);
xnor UO_3206 (O_3206,N_29094,N_29052);
nor UO_3207 (O_3207,N_29550,N_28984);
and UO_3208 (O_3208,N_29321,N_29744);
nand UO_3209 (O_3209,N_29259,N_28822);
nor UO_3210 (O_3210,N_28551,N_29759);
or UO_3211 (O_3211,N_28817,N_29055);
or UO_3212 (O_3212,N_28599,N_28810);
or UO_3213 (O_3213,N_29467,N_28589);
nor UO_3214 (O_3214,N_29517,N_29118);
nand UO_3215 (O_3215,N_29844,N_29233);
and UO_3216 (O_3216,N_29070,N_29240);
xor UO_3217 (O_3217,N_29573,N_29421);
and UO_3218 (O_3218,N_28593,N_28559);
nand UO_3219 (O_3219,N_29974,N_28853);
nand UO_3220 (O_3220,N_29624,N_29665);
nor UO_3221 (O_3221,N_29973,N_28847);
and UO_3222 (O_3222,N_29849,N_29289);
xnor UO_3223 (O_3223,N_29053,N_29031);
or UO_3224 (O_3224,N_28601,N_28659);
or UO_3225 (O_3225,N_29788,N_29047);
nor UO_3226 (O_3226,N_29080,N_29749);
xnor UO_3227 (O_3227,N_28675,N_28754);
and UO_3228 (O_3228,N_28791,N_29746);
nand UO_3229 (O_3229,N_28575,N_29069);
nand UO_3230 (O_3230,N_29321,N_29237);
xor UO_3231 (O_3231,N_28625,N_29231);
xor UO_3232 (O_3232,N_28884,N_28854);
and UO_3233 (O_3233,N_29536,N_29788);
nor UO_3234 (O_3234,N_28578,N_29357);
xor UO_3235 (O_3235,N_29952,N_28571);
nand UO_3236 (O_3236,N_28591,N_29444);
or UO_3237 (O_3237,N_29081,N_28805);
nor UO_3238 (O_3238,N_28989,N_28916);
nor UO_3239 (O_3239,N_29652,N_29523);
and UO_3240 (O_3240,N_29740,N_28523);
xnor UO_3241 (O_3241,N_28918,N_29058);
and UO_3242 (O_3242,N_29697,N_28878);
or UO_3243 (O_3243,N_29502,N_29824);
nand UO_3244 (O_3244,N_29523,N_29133);
nand UO_3245 (O_3245,N_29986,N_29547);
or UO_3246 (O_3246,N_28862,N_29730);
or UO_3247 (O_3247,N_29919,N_29399);
or UO_3248 (O_3248,N_29832,N_29060);
xnor UO_3249 (O_3249,N_28585,N_29126);
nor UO_3250 (O_3250,N_29458,N_28504);
and UO_3251 (O_3251,N_28756,N_29533);
and UO_3252 (O_3252,N_29085,N_28872);
or UO_3253 (O_3253,N_29316,N_28613);
nand UO_3254 (O_3254,N_29777,N_29143);
and UO_3255 (O_3255,N_29457,N_28506);
nor UO_3256 (O_3256,N_28847,N_29396);
and UO_3257 (O_3257,N_28642,N_28557);
and UO_3258 (O_3258,N_29512,N_29586);
nor UO_3259 (O_3259,N_29281,N_29419);
nor UO_3260 (O_3260,N_29273,N_29614);
nor UO_3261 (O_3261,N_29100,N_28850);
or UO_3262 (O_3262,N_29555,N_29370);
nand UO_3263 (O_3263,N_29807,N_29626);
xnor UO_3264 (O_3264,N_28670,N_28500);
and UO_3265 (O_3265,N_29061,N_29704);
and UO_3266 (O_3266,N_29376,N_28694);
and UO_3267 (O_3267,N_29031,N_29426);
nor UO_3268 (O_3268,N_29615,N_28658);
xor UO_3269 (O_3269,N_29387,N_29572);
and UO_3270 (O_3270,N_28696,N_28767);
xor UO_3271 (O_3271,N_29056,N_28672);
nor UO_3272 (O_3272,N_29305,N_29804);
nand UO_3273 (O_3273,N_28808,N_28855);
and UO_3274 (O_3274,N_28755,N_29878);
and UO_3275 (O_3275,N_29600,N_28525);
or UO_3276 (O_3276,N_29307,N_28778);
nor UO_3277 (O_3277,N_29111,N_29908);
xor UO_3278 (O_3278,N_29864,N_28801);
nor UO_3279 (O_3279,N_28697,N_29164);
and UO_3280 (O_3280,N_29350,N_29470);
nor UO_3281 (O_3281,N_29849,N_29453);
or UO_3282 (O_3282,N_28613,N_29130);
xnor UO_3283 (O_3283,N_28768,N_29413);
xnor UO_3284 (O_3284,N_29488,N_28905);
or UO_3285 (O_3285,N_29533,N_29343);
nor UO_3286 (O_3286,N_29740,N_29253);
and UO_3287 (O_3287,N_29349,N_29374);
xor UO_3288 (O_3288,N_28802,N_29614);
or UO_3289 (O_3289,N_29248,N_29499);
and UO_3290 (O_3290,N_29979,N_28959);
xnor UO_3291 (O_3291,N_29473,N_28744);
nand UO_3292 (O_3292,N_28508,N_28964);
nor UO_3293 (O_3293,N_29514,N_28504);
and UO_3294 (O_3294,N_29604,N_29289);
nand UO_3295 (O_3295,N_28888,N_28529);
nor UO_3296 (O_3296,N_29105,N_29196);
or UO_3297 (O_3297,N_28712,N_29605);
nor UO_3298 (O_3298,N_29454,N_29443);
xor UO_3299 (O_3299,N_29462,N_29689);
nand UO_3300 (O_3300,N_29271,N_29593);
xor UO_3301 (O_3301,N_29056,N_28947);
nor UO_3302 (O_3302,N_29917,N_28588);
nor UO_3303 (O_3303,N_28531,N_29101);
xnor UO_3304 (O_3304,N_29481,N_28979);
and UO_3305 (O_3305,N_29428,N_29594);
or UO_3306 (O_3306,N_29510,N_28822);
xnor UO_3307 (O_3307,N_29583,N_28675);
and UO_3308 (O_3308,N_28982,N_28883);
or UO_3309 (O_3309,N_28630,N_29829);
and UO_3310 (O_3310,N_29142,N_29939);
xnor UO_3311 (O_3311,N_29190,N_29410);
nand UO_3312 (O_3312,N_28539,N_28572);
and UO_3313 (O_3313,N_29143,N_29442);
nor UO_3314 (O_3314,N_29971,N_29708);
xnor UO_3315 (O_3315,N_29060,N_29501);
xor UO_3316 (O_3316,N_29666,N_28602);
nor UO_3317 (O_3317,N_28991,N_29532);
nor UO_3318 (O_3318,N_28744,N_29891);
xnor UO_3319 (O_3319,N_28901,N_29080);
nand UO_3320 (O_3320,N_29119,N_28869);
nand UO_3321 (O_3321,N_29438,N_29631);
or UO_3322 (O_3322,N_29548,N_28803);
xor UO_3323 (O_3323,N_29627,N_29926);
and UO_3324 (O_3324,N_29691,N_29318);
nand UO_3325 (O_3325,N_29464,N_29266);
nor UO_3326 (O_3326,N_28865,N_29883);
and UO_3327 (O_3327,N_28585,N_29881);
nand UO_3328 (O_3328,N_29273,N_29388);
or UO_3329 (O_3329,N_29626,N_28517);
or UO_3330 (O_3330,N_28730,N_28823);
and UO_3331 (O_3331,N_29322,N_28841);
nor UO_3332 (O_3332,N_28817,N_29975);
nand UO_3333 (O_3333,N_28506,N_29943);
nand UO_3334 (O_3334,N_28776,N_29663);
nand UO_3335 (O_3335,N_29512,N_29244);
nor UO_3336 (O_3336,N_29766,N_28589);
xor UO_3337 (O_3337,N_28619,N_29727);
nand UO_3338 (O_3338,N_29912,N_29381);
nor UO_3339 (O_3339,N_29919,N_29876);
nor UO_3340 (O_3340,N_29012,N_29878);
xnor UO_3341 (O_3341,N_29331,N_28766);
or UO_3342 (O_3342,N_29316,N_29116);
or UO_3343 (O_3343,N_29634,N_29227);
xor UO_3344 (O_3344,N_28882,N_29097);
nand UO_3345 (O_3345,N_29604,N_29524);
and UO_3346 (O_3346,N_29104,N_28975);
and UO_3347 (O_3347,N_29444,N_29866);
nor UO_3348 (O_3348,N_29128,N_29801);
nor UO_3349 (O_3349,N_29409,N_29892);
and UO_3350 (O_3350,N_29487,N_29621);
or UO_3351 (O_3351,N_28786,N_28551);
or UO_3352 (O_3352,N_29394,N_28963);
or UO_3353 (O_3353,N_29044,N_29333);
or UO_3354 (O_3354,N_29882,N_28938);
xor UO_3355 (O_3355,N_29006,N_28980);
or UO_3356 (O_3356,N_29118,N_29091);
nand UO_3357 (O_3357,N_29148,N_29059);
or UO_3358 (O_3358,N_29012,N_29915);
nor UO_3359 (O_3359,N_28769,N_29791);
nor UO_3360 (O_3360,N_28876,N_29580);
nor UO_3361 (O_3361,N_28906,N_29838);
nand UO_3362 (O_3362,N_28595,N_28612);
xor UO_3363 (O_3363,N_29666,N_29773);
nand UO_3364 (O_3364,N_28659,N_29498);
xor UO_3365 (O_3365,N_29639,N_29257);
nand UO_3366 (O_3366,N_28726,N_28839);
xor UO_3367 (O_3367,N_29243,N_29129);
nor UO_3368 (O_3368,N_29351,N_29274);
xor UO_3369 (O_3369,N_28530,N_28702);
or UO_3370 (O_3370,N_29497,N_29930);
nor UO_3371 (O_3371,N_29990,N_29228);
xor UO_3372 (O_3372,N_29123,N_29911);
or UO_3373 (O_3373,N_29590,N_28848);
nand UO_3374 (O_3374,N_29097,N_29263);
or UO_3375 (O_3375,N_29758,N_28735);
nor UO_3376 (O_3376,N_29394,N_29239);
or UO_3377 (O_3377,N_29905,N_29722);
nor UO_3378 (O_3378,N_28833,N_29880);
xor UO_3379 (O_3379,N_29323,N_28991);
and UO_3380 (O_3380,N_28645,N_29983);
and UO_3381 (O_3381,N_29183,N_29317);
xor UO_3382 (O_3382,N_29531,N_29310);
nand UO_3383 (O_3383,N_28739,N_28979);
or UO_3384 (O_3384,N_29154,N_29586);
nor UO_3385 (O_3385,N_29469,N_28561);
or UO_3386 (O_3386,N_29597,N_29795);
nand UO_3387 (O_3387,N_29457,N_29161);
and UO_3388 (O_3388,N_29259,N_29792);
and UO_3389 (O_3389,N_28949,N_29442);
and UO_3390 (O_3390,N_29477,N_28690);
xnor UO_3391 (O_3391,N_29542,N_29062);
nand UO_3392 (O_3392,N_29579,N_28838);
xnor UO_3393 (O_3393,N_29524,N_28525);
or UO_3394 (O_3394,N_29038,N_28506);
and UO_3395 (O_3395,N_29692,N_29631);
nand UO_3396 (O_3396,N_29261,N_28885);
nand UO_3397 (O_3397,N_29690,N_29434);
nor UO_3398 (O_3398,N_29226,N_29155);
or UO_3399 (O_3399,N_29364,N_29894);
nand UO_3400 (O_3400,N_29988,N_28642);
nand UO_3401 (O_3401,N_28669,N_29033);
nor UO_3402 (O_3402,N_28738,N_29343);
xnor UO_3403 (O_3403,N_29211,N_29265);
xnor UO_3404 (O_3404,N_29383,N_28907);
nor UO_3405 (O_3405,N_29656,N_28908);
nor UO_3406 (O_3406,N_29160,N_29713);
xnor UO_3407 (O_3407,N_29918,N_29520);
or UO_3408 (O_3408,N_29584,N_28854);
nand UO_3409 (O_3409,N_29763,N_29907);
or UO_3410 (O_3410,N_29668,N_28678);
nor UO_3411 (O_3411,N_29745,N_29274);
and UO_3412 (O_3412,N_29338,N_29178);
nor UO_3413 (O_3413,N_29547,N_29066);
xor UO_3414 (O_3414,N_28711,N_28792);
nor UO_3415 (O_3415,N_28672,N_29069);
xor UO_3416 (O_3416,N_29983,N_29198);
nor UO_3417 (O_3417,N_29861,N_29742);
and UO_3418 (O_3418,N_29483,N_29011);
nand UO_3419 (O_3419,N_29196,N_29499);
and UO_3420 (O_3420,N_29651,N_29783);
and UO_3421 (O_3421,N_28978,N_29571);
or UO_3422 (O_3422,N_28700,N_29492);
xor UO_3423 (O_3423,N_29160,N_28626);
nor UO_3424 (O_3424,N_29766,N_29729);
nor UO_3425 (O_3425,N_29477,N_29704);
xor UO_3426 (O_3426,N_29803,N_28553);
nand UO_3427 (O_3427,N_29185,N_29400);
and UO_3428 (O_3428,N_28988,N_29185);
and UO_3429 (O_3429,N_29374,N_29634);
nor UO_3430 (O_3430,N_29849,N_29880);
or UO_3431 (O_3431,N_28737,N_29414);
xnor UO_3432 (O_3432,N_29013,N_28559);
nor UO_3433 (O_3433,N_28636,N_28769);
and UO_3434 (O_3434,N_29933,N_29195);
nand UO_3435 (O_3435,N_29233,N_28607);
nor UO_3436 (O_3436,N_29659,N_28648);
or UO_3437 (O_3437,N_29530,N_29281);
or UO_3438 (O_3438,N_29848,N_29036);
nor UO_3439 (O_3439,N_29502,N_28635);
xnor UO_3440 (O_3440,N_29608,N_28988);
and UO_3441 (O_3441,N_28854,N_28832);
and UO_3442 (O_3442,N_29525,N_28949);
and UO_3443 (O_3443,N_29678,N_29926);
nand UO_3444 (O_3444,N_29597,N_28758);
xor UO_3445 (O_3445,N_29080,N_28933);
or UO_3446 (O_3446,N_29401,N_28771);
and UO_3447 (O_3447,N_29143,N_29904);
and UO_3448 (O_3448,N_29596,N_28712);
nand UO_3449 (O_3449,N_29539,N_29173);
nand UO_3450 (O_3450,N_29460,N_29336);
nand UO_3451 (O_3451,N_28644,N_28947);
nand UO_3452 (O_3452,N_29740,N_29489);
or UO_3453 (O_3453,N_29067,N_28760);
nand UO_3454 (O_3454,N_29723,N_28597);
and UO_3455 (O_3455,N_28925,N_29695);
xor UO_3456 (O_3456,N_29107,N_29776);
or UO_3457 (O_3457,N_29517,N_29679);
nor UO_3458 (O_3458,N_29196,N_28673);
nand UO_3459 (O_3459,N_28658,N_29553);
nor UO_3460 (O_3460,N_28709,N_29740);
xor UO_3461 (O_3461,N_28829,N_28809);
nand UO_3462 (O_3462,N_29272,N_29296);
or UO_3463 (O_3463,N_29015,N_28735);
nor UO_3464 (O_3464,N_28747,N_28791);
nor UO_3465 (O_3465,N_28975,N_29379);
or UO_3466 (O_3466,N_29681,N_28986);
xor UO_3467 (O_3467,N_29264,N_28602);
xnor UO_3468 (O_3468,N_28835,N_29675);
nor UO_3469 (O_3469,N_28764,N_29652);
nor UO_3470 (O_3470,N_28910,N_28985);
or UO_3471 (O_3471,N_29024,N_29785);
and UO_3472 (O_3472,N_28614,N_29266);
nor UO_3473 (O_3473,N_29426,N_29193);
nand UO_3474 (O_3474,N_29836,N_29780);
or UO_3475 (O_3475,N_29327,N_28725);
nor UO_3476 (O_3476,N_29876,N_29670);
xor UO_3477 (O_3477,N_29512,N_29884);
or UO_3478 (O_3478,N_29658,N_28843);
nand UO_3479 (O_3479,N_29348,N_28956);
or UO_3480 (O_3480,N_29560,N_28511);
nand UO_3481 (O_3481,N_29635,N_29278);
nor UO_3482 (O_3482,N_29835,N_29099);
and UO_3483 (O_3483,N_28969,N_29289);
nor UO_3484 (O_3484,N_28580,N_29144);
nand UO_3485 (O_3485,N_29268,N_29339);
or UO_3486 (O_3486,N_29474,N_29878);
and UO_3487 (O_3487,N_28953,N_29046);
xnor UO_3488 (O_3488,N_29909,N_29285);
nor UO_3489 (O_3489,N_28637,N_28923);
xnor UO_3490 (O_3490,N_28505,N_29134);
nor UO_3491 (O_3491,N_29292,N_28808);
nor UO_3492 (O_3492,N_28923,N_28587);
and UO_3493 (O_3493,N_28814,N_29918);
or UO_3494 (O_3494,N_28933,N_28760);
nor UO_3495 (O_3495,N_29100,N_29149);
xor UO_3496 (O_3496,N_29422,N_29874);
and UO_3497 (O_3497,N_28737,N_29859);
nand UO_3498 (O_3498,N_29607,N_29312);
nand UO_3499 (O_3499,N_29730,N_29323);
endmodule