module basic_500_3000_500_40_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_296,In_415);
xnor U1 (N_1,In_324,In_476);
nand U2 (N_2,In_217,In_27);
xor U3 (N_3,In_123,In_224);
and U4 (N_4,In_312,In_180);
nor U5 (N_5,In_348,In_406);
or U6 (N_6,In_298,In_332);
or U7 (N_7,In_439,In_374);
nor U8 (N_8,In_148,In_239);
nand U9 (N_9,In_183,In_231);
nand U10 (N_10,In_256,In_350);
nor U11 (N_11,In_356,In_252);
nor U12 (N_12,In_15,In_477);
nor U13 (N_13,In_488,In_301);
xor U14 (N_14,In_54,In_216);
or U15 (N_15,In_331,In_293);
nor U16 (N_16,In_174,In_479);
and U17 (N_17,In_189,In_138);
and U18 (N_18,In_264,In_468);
xor U19 (N_19,In_47,In_304);
nor U20 (N_20,In_319,In_421);
nor U21 (N_21,In_462,In_107);
nand U22 (N_22,In_418,In_170);
nor U23 (N_23,In_494,In_102);
or U24 (N_24,In_59,In_105);
xor U25 (N_25,In_288,In_423);
nor U26 (N_26,In_93,In_145);
and U27 (N_27,In_322,In_339);
nor U28 (N_28,In_393,In_355);
xor U29 (N_29,In_318,In_237);
nor U30 (N_30,In_436,In_323);
nand U31 (N_31,In_362,In_291);
and U32 (N_32,In_26,In_354);
nor U33 (N_33,In_390,In_70);
nand U34 (N_34,In_140,In_430);
xnor U35 (N_35,In_413,In_81);
and U36 (N_36,In_317,In_187);
nand U37 (N_37,In_375,In_313);
and U38 (N_38,In_46,In_396);
nor U39 (N_39,In_17,In_496);
and U40 (N_40,In_246,In_410);
and U41 (N_41,In_94,In_340);
and U42 (N_42,In_156,In_35);
nand U43 (N_43,In_172,In_97);
nor U44 (N_44,In_425,In_162);
or U45 (N_45,In_474,In_297);
or U46 (N_46,In_361,In_403);
or U47 (N_47,In_447,In_20);
nor U48 (N_48,In_373,In_25);
and U49 (N_49,In_490,In_167);
or U50 (N_50,In_409,In_249);
or U51 (N_51,In_21,In_111);
nor U52 (N_52,In_214,In_96);
nand U53 (N_53,In_234,In_446);
nand U54 (N_54,In_364,In_404);
nor U55 (N_55,In_248,In_328);
nor U56 (N_56,In_75,In_386);
nor U57 (N_57,In_407,In_0);
and U58 (N_58,In_456,In_347);
and U59 (N_59,In_242,In_114);
and U60 (N_60,In_177,In_441);
and U61 (N_61,In_470,In_427);
or U62 (N_62,In_98,In_487);
and U63 (N_63,In_334,In_371);
nor U64 (N_64,In_58,In_164);
nor U65 (N_65,In_306,In_119);
and U66 (N_66,In_489,In_49);
or U67 (N_67,In_417,In_357);
or U68 (N_68,In_336,In_48);
nor U69 (N_69,In_163,In_268);
nor U70 (N_70,In_335,In_157);
and U71 (N_71,In_220,In_330);
or U72 (N_72,In_181,In_30);
nor U73 (N_73,In_397,In_428);
nor U74 (N_74,In_38,In_192);
or U75 (N_75,In_412,In_86);
and U76 (N_76,In_414,N_66);
and U77 (N_77,In_118,N_35);
and U78 (N_78,In_92,In_314);
nor U79 (N_79,N_72,In_22);
and U80 (N_80,N_20,In_395);
and U81 (N_81,In_131,In_465);
and U82 (N_82,In_139,In_60);
and U83 (N_83,In_154,In_377);
nand U84 (N_84,In_241,In_121);
nand U85 (N_85,In_196,In_55);
and U86 (N_86,In_277,N_41);
or U87 (N_87,In_448,In_169);
or U88 (N_88,In_73,In_50);
nor U89 (N_89,In_345,In_41);
or U90 (N_90,In_278,In_191);
nand U91 (N_91,In_7,N_6);
nand U92 (N_92,In_101,In_302);
nor U93 (N_93,In_360,In_178);
nor U94 (N_94,In_149,In_284);
and U95 (N_95,In_150,In_270);
nor U96 (N_96,In_272,In_303);
nand U97 (N_97,N_32,In_159);
and U98 (N_98,In_218,N_33);
and U99 (N_99,In_28,N_53);
nor U100 (N_100,In_32,In_199);
nor U101 (N_101,N_73,In_385);
nand U102 (N_102,In_308,In_299);
or U103 (N_103,In_112,N_67);
or U104 (N_104,In_126,N_24);
nand U105 (N_105,In_52,N_18);
nor U106 (N_106,In_37,N_13);
and U107 (N_107,In_255,In_85);
and U108 (N_108,In_295,In_491);
nand U109 (N_109,In_51,In_369);
or U110 (N_110,In_440,In_10);
nor U111 (N_111,N_1,In_457);
nor U112 (N_112,In_432,N_49);
and U113 (N_113,N_36,In_84);
nand U114 (N_114,In_168,In_482);
and U115 (N_115,In_435,In_113);
or U116 (N_116,In_144,In_245);
nand U117 (N_117,In_160,In_387);
and U118 (N_118,In_247,In_100);
or U119 (N_119,In_115,In_333);
nor U120 (N_120,In_275,In_405);
and U121 (N_121,In_8,In_53);
nand U122 (N_122,In_290,In_108);
and U123 (N_123,In_327,In_408);
nor U124 (N_124,In_366,In_307);
or U125 (N_125,In_380,In_207);
nand U126 (N_126,In_120,In_473);
or U127 (N_127,In_254,In_212);
nand U128 (N_128,In_244,In_176);
or U129 (N_129,N_59,In_135);
xnor U130 (N_130,In_351,N_68);
nand U131 (N_131,In_469,In_151);
and U132 (N_132,In_5,In_34);
and U133 (N_133,N_63,In_99);
nor U134 (N_134,In_147,N_2);
and U135 (N_135,In_424,In_230);
nand U136 (N_136,In_226,In_341);
or U137 (N_137,N_64,In_376);
nand U138 (N_138,N_7,In_36);
or U139 (N_139,In_219,In_227);
nor U140 (N_140,In_292,In_280);
nand U141 (N_141,In_40,In_240);
or U142 (N_142,In_184,In_14);
nand U143 (N_143,In_250,In_103);
nand U144 (N_144,In_186,In_394);
or U145 (N_145,In_95,In_261);
or U146 (N_146,In_276,In_3);
xnor U147 (N_147,N_15,In_152);
or U148 (N_148,In_200,In_266);
nor U149 (N_149,In_11,In_461);
or U150 (N_150,In_72,N_110);
or U151 (N_151,In_78,In_236);
nand U152 (N_152,N_14,N_5);
and U153 (N_153,In_143,In_420);
or U154 (N_154,N_109,In_451);
or U155 (N_155,In_353,In_197);
nand U156 (N_156,In_453,In_201);
or U157 (N_157,In_315,N_116);
nand U158 (N_158,N_12,In_82);
and U159 (N_159,In_158,In_124);
and U160 (N_160,N_87,N_22);
nor U161 (N_161,In_274,N_62);
or U162 (N_162,In_76,In_251);
or U163 (N_163,N_149,In_179);
nand U164 (N_164,In_223,N_69);
nor U165 (N_165,In_188,In_459);
or U166 (N_166,N_144,In_475);
nor U167 (N_167,In_260,In_210);
or U168 (N_168,In_259,In_358);
nand U169 (N_169,N_78,In_381);
nand U170 (N_170,In_87,In_182);
or U171 (N_171,In_205,In_134);
nand U172 (N_172,In_80,In_311);
nand U173 (N_173,N_0,In_391);
nor U174 (N_174,In_401,In_392);
xnor U175 (N_175,In_44,In_171);
and U176 (N_176,N_141,In_206);
and U177 (N_177,In_438,In_166);
and U178 (N_178,In_283,In_122);
or U179 (N_179,In_43,N_107);
or U180 (N_180,In_463,In_19);
nand U181 (N_181,In_130,In_454);
nand U182 (N_182,In_16,In_363);
and U183 (N_183,N_130,N_95);
nor U184 (N_184,In_471,In_271);
or U185 (N_185,In_128,In_6);
and U186 (N_186,N_44,N_89);
nand U187 (N_187,N_28,In_88);
nor U188 (N_188,N_80,In_63);
nor U189 (N_189,N_47,In_127);
nand U190 (N_190,In_203,In_285);
and U191 (N_191,In_384,In_359);
nand U192 (N_192,N_85,In_225);
or U193 (N_193,In_495,N_88);
xnor U194 (N_194,In_342,In_24);
nor U195 (N_195,In_265,N_11);
and U196 (N_196,In_57,N_9);
nor U197 (N_197,N_92,In_222);
nor U198 (N_198,In_452,N_125);
and U199 (N_199,In_9,In_56);
or U200 (N_200,In_398,In_208);
nor U201 (N_201,In_137,N_51);
and U202 (N_202,In_13,In_258);
and U203 (N_203,N_119,In_287);
nor U204 (N_204,In_337,In_116);
or U205 (N_205,In_77,In_91);
and U206 (N_206,In_343,In_195);
and U207 (N_207,N_118,N_117);
nor U208 (N_208,In_444,In_23);
or U209 (N_209,N_104,N_111);
and U210 (N_210,In_173,N_105);
nor U211 (N_211,In_455,In_243);
nand U212 (N_212,N_131,In_281);
nor U213 (N_213,N_40,N_8);
or U214 (N_214,N_124,In_229);
and U215 (N_215,In_133,In_213);
nand U216 (N_216,N_137,In_29);
nand U217 (N_217,N_34,N_112);
or U218 (N_218,In_309,In_483);
or U219 (N_219,In_419,In_185);
xnor U220 (N_220,N_106,N_93);
or U221 (N_221,N_126,N_143);
xnor U222 (N_222,In_485,In_365);
nor U223 (N_223,In_399,N_122);
nor U224 (N_224,In_190,In_458);
or U225 (N_225,In_62,N_84);
and U226 (N_226,N_193,N_65);
nand U227 (N_227,N_181,In_202);
nand U228 (N_228,In_464,N_4);
nor U229 (N_229,N_102,N_57);
and U230 (N_230,In_132,N_195);
and U231 (N_231,N_101,In_372);
and U232 (N_232,N_170,N_163);
nor U233 (N_233,In_316,In_478);
nor U234 (N_234,N_90,In_39);
or U235 (N_235,In_480,In_45);
nand U236 (N_236,N_153,In_194);
and U237 (N_237,N_145,In_106);
nor U238 (N_238,N_182,N_140);
nor U239 (N_239,N_60,N_76);
xor U240 (N_240,In_71,N_25);
and U241 (N_241,In_33,N_175);
nor U242 (N_242,N_100,In_267);
or U243 (N_243,N_142,In_155);
and U244 (N_244,In_370,In_338);
nor U245 (N_245,In_69,N_211);
or U246 (N_246,In_228,In_310);
nand U247 (N_247,In_257,N_98);
nor U248 (N_248,N_129,In_67);
nand U249 (N_249,N_45,N_91);
nor U250 (N_250,N_192,In_110);
nor U251 (N_251,N_43,N_29);
nand U252 (N_252,N_139,In_389);
and U253 (N_253,N_169,In_273);
or U254 (N_254,N_177,In_198);
or U255 (N_255,N_113,In_129);
nand U256 (N_256,N_152,N_220);
nor U257 (N_257,N_38,N_61);
or U258 (N_258,In_499,N_198);
and U259 (N_259,N_205,In_422);
and U260 (N_260,N_171,N_162);
or U261 (N_261,N_179,N_196);
nand U262 (N_262,N_56,N_223);
nor U263 (N_263,In_329,In_450);
nor U264 (N_264,N_58,N_75);
nor U265 (N_265,N_82,In_294);
nand U266 (N_266,N_99,In_42);
nand U267 (N_267,N_133,N_121);
nor U268 (N_268,In_64,In_1);
nand U269 (N_269,N_127,N_176);
or U270 (N_270,In_141,N_197);
and U271 (N_271,In_445,N_31);
nor U272 (N_272,In_497,N_180);
or U273 (N_273,N_46,In_125);
or U274 (N_274,N_54,N_218);
nand U275 (N_275,In_79,N_108);
or U276 (N_276,In_238,N_39);
nor U277 (N_277,In_175,In_215);
nand U278 (N_278,N_200,In_378);
and U279 (N_279,In_136,In_31);
or U280 (N_280,N_189,N_103);
or U281 (N_281,N_52,N_30);
nor U282 (N_282,N_212,N_132);
nand U283 (N_283,N_120,N_190);
or U284 (N_284,In_18,In_320);
nor U285 (N_285,In_346,N_174);
nor U286 (N_286,N_214,In_4);
nand U287 (N_287,In_65,In_193);
nor U288 (N_288,N_79,N_207);
nand U289 (N_289,In_486,In_382);
and U290 (N_290,N_157,N_26);
and U291 (N_291,N_96,In_305);
nand U292 (N_292,N_213,N_187);
or U293 (N_293,N_202,N_167);
and U294 (N_294,In_279,In_282);
nor U295 (N_295,N_165,N_154);
nor U296 (N_296,In_493,In_300);
nor U297 (N_297,N_210,In_221);
nor U298 (N_298,In_431,N_71);
nand U299 (N_299,In_442,N_222);
or U300 (N_300,N_238,N_270);
nor U301 (N_301,N_263,N_86);
or U302 (N_302,N_81,In_443);
or U303 (N_303,N_243,In_153);
nand U304 (N_304,N_42,In_429);
or U305 (N_305,N_249,In_400);
nand U306 (N_306,N_274,N_50);
nor U307 (N_307,N_159,N_256);
nor U308 (N_308,N_209,In_146);
nand U309 (N_309,In_321,N_183);
and U310 (N_310,N_224,N_156);
nand U311 (N_311,N_269,N_10);
or U312 (N_312,In_388,In_383);
and U313 (N_313,In_68,In_117);
nand U314 (N_314,N_281,N_246);
and U315 (N_315,N_275,N_204);
or U316 (N_316,In_289,N_173);
nand U317 (N_317,N_286,In_83);
nor U318 (N_318,In_498,In_209);
nand U319 (N_319,N_288,N_236);
nor U320 (N_320,N_215,N_294);
nor U321 (N_321,N_16,N_283);
and U322 (N_322,In_433,In_204);
nor U323 (N_323,N_241,N_19);
or U324 (N_324,N_250,N_234);
nand U325 (N_325,N_261,N_248);
and U326 (N_326,In_437,N_295);
and U327 (N_327,N_199,N_146);
nor U328 (N_328,N_221,In_379);
or U329 (N_329,N_55,N_266);
and U330 (N_330,In_262,N_186);
nand U331 (N_331,N_259,In_61);
nand U332 (N_332,N_147,N_237);
or U333 (N_333,In_426,N_226);
xnor U334 (N_334,N_292,N_164);
and U335 (N_335,In_411,N_216);
or U336 (N_336,N_228,N_225);
or U337 (N_337,In_492,In_434);
or U338 (N_338,N_245,N_148);
nand U339 (N_339,In_466,N_252);
or U340 (N_340,In_269,N_206);
nand U341 (N_341,N_285,In_104);
nor U342 (N_342,N_115,N_282);
and U343 (N_343,N_27,In_74);
or U344 (N_344,In_349,N_297);
or U345 (N_345,N_217,N_208);
or U346 (N_346,N_279,In_286);
or U347 (N_347,In_484,N_136);
xnor U348 (N_348,In_211,N_188);
nor U349 (N_349,N_254,In_263);
nor U350 (N_350,In_460,N_227);
and U351 (N_351,N_134,N_97);
nand U352 (N_352,In_165,N_191);
or U353 (N_353,In_2,In_235);
or U354 (N_354,N_155,N_290);
or U355 (N_355,N_150,N_17);
nor U356 (N_356,In_481,N_253);
and U357 (N_357,N_178,In_161);
or U358 (N_358,N_293,In_66);
and U359 (N_359,In_233,N_172);
and U360 (N_360,N_151,N_94);
or U361 (N_361,N_160,N_114);
nor U362 (N_362,N_203,N_185);
or U363 (N_363,N_299,N_158);
nor U364 (N_364,In_142,N_267);
nor U365 (N_365,In_325,N_219);
and U366 (N_366,In_89,In_402);
nand U367 (N_367,In_367,N_255);
nand U368 (N_368,N_272,N_70);
or U369 (N_369,N_289,N_276);
nand U370 (N_370,N_201,N_264);
xnor U371 (N_371,In_467,N_135);
or U372 (N_372,N_287,N_48);
nand U373 (N_373,N_23,N_3);
and U374 (N_374,N_74,In_449);
nor U375 (N_375,N_324,N_359);
and U376 (N_376,N_331,N_332);
and U377 (N_377,N_291,N_361);
nand U378 (N_378,N_262,In_352);
nand U379 (N_379,N_341,N_347);
and U380 (N_380,N_307,In_109);
or U381 (N_381,N_358,N_345);
nand U382 (N_382,N_356,N_330);
nand U383 (N_383,N_138,N_373);
xnor U384 (N_384,N_360,N_369);
or U385 (N_385,N_333,In_253);
or U386 (N_386,N_320,N_364);
and U387 (N_387,N_326,N_317);
nor U388 (N_388,N_350,N_346);
or U389 (N_389,N_239,N_268);
or U390 (N_390,N_368,N_240);
nand U391 (N_391,N_230,N_344);
and U392 (N_392,N_351,N_296);
and U393 (N_393,N_314,In_368);
nor U394 (N_394,N_349,N_371);
nor U395 (N_395,In_326,N_309);
or U396 (N_396,N_325,In_12);
nor U397 (N_397,In_416,N_21);
nand U398 (N_398,N_298,N_319);
nor U399 (N_399,N_302,N_329);
or U400 (N_400,N_322,N_305);
nand U401 (N_401,N_370,N_280);
or U402 (N_402,N_316,N_339);
nand U403 (N_403,In_232,N_271);
and U404 (N_404,N_321,N_355);
or U405 (N_405,N_374,N_323);
or U406 (N_406,N_336,N_278);
or U407 (N_407,N_308,N_306);
or U408 (N_408,N_334,N_363);
nor U409 (N_409,N_343,N_258);
or U410 (N_410,In_472,N_310);
nand U411 (N_411,N_229,N_232);
nand U412 (N_412,N_367,N_168);
nand U413 (N_413,N_335,N_265);
nand U414 (N_414,N_313,N_357);
nand U415 (N_415,N_338,N_247);
xor U416 (N_416,N_37,N_311);
nand U417 (N_417,N_184,N_83);
xor U418 (N_418,N_366,N_312);
nand U419 (N_419,N_327,N_251);
and U420 (N_420,N_194,N_300);
or U421 (N_421,N_123,In_90);
nand U422 (N_422,N_244,N_303);
xor U423 (N_423,N_352,In_344);
or U424 (N_424,N_354,N_242);
nor U425 (N_425,N_166,N_318);
nand U426 (N_426,N_284,N_128);
or U427 (N_427,N_235,N_304);
and U428 (N_428,N_362,N_77);
and U429 (N_429,N_301,N_342);
and U430 (N_430,N_231,N_372);
and U431 (N_431,N_277,N_337);
xor U432 (N_432,N_353,N_257);
and U433 (N_433,N_365,N_328);
nor U434 (N_434,N_233,N_260);
nor U435 (N_435,N_161,N_315);
and U436 (N_436,N_340,N_273);
xor U437 (N_437,N_348,N_364);
nand U438 (N_438,N_325,N_308);
nand U439 (N_439,N_349,N_336);
nor U440 (N_440,N_77,N_333);
nand U441 (N_441,N_334,N_336);
nand U442 (N_442,N_367,In_12);
or U443 (N_443,N_240,N_352);
nand U444 (N_444,N_326,N_339);
or U445 (N_445,N_305,N_229);
and U446 (N_446,N_242,N_83);
nand U447 (N_447,In_368,N_128);
or U448 (N_448,N_336,N_232);
and U449 (N_449,N_306,N_268);
or U450 (N_450,N_386,N_441);
or U451 (N_451,N_396,N_378);
and U452 (N_452,N_379,N_417);
or U453 (N_453,N_411,N_383);
and U454 (N_454,N_399,N_433);
nand U455 (N_455,N_427,N_413);
nor U456 (N_456,N_403,N_415);
and U457 (N_457,N_442,N_430);
nand U458 (N_458,N_416,N_388);
and U459 (N_459,N_406,N_381);
xor U460 (N_460,N_444,N_449);
nor U461 (N_461,N_432,N_409);
nand U462 (N_462,N_407,N_385);
nor U463 (N_463,N_422,N_418);
xor U464 (N_464,N_426,N_446);
nand U465 (N_465,N_448,N_419);
and U466 (N_466,N_437,N_440);
or U467 (N_467,N_424,N_404);
nand U468 (N_468,N_402,N_423);
and U469 (N_469,N_376,N_387);
nand U470 (N_470,N_412,N_429);
or U471 (N_471,N_377,N_375);
and U472 (N_472,N_397,N_414);
nand U473 (N_473,N_436,N_408);
xor U474 (N_474,N_384,N_443);
nand U475 (N_475,N_410,N_401);
or U476 (N_476,N_400,N_421);
xnor U477 (N_477,N_445,N_382);
nand U478 (N_478,N_434,N_380);
nand U479 (N_479,N_439,N_425);
and U480 (N_480,N_398,N_405);
xnor U481 (N_481,N_392,N_447);
and U482 (N_482,N_393,N_390);
nor U483 (N_483,N_389,N_438);
nor U484 (N_484,N_428,N_431);
and U485 (N_485,N_391,N_435);
or U486 (N_486,N_420,N_395);
nand U487 (N_487,N_394,N_378);
or U488 (N_488,N_383,N_445);
and U489 (N_489,N_427,N_404);
or U490 (N_490,N_410,N_406);
nand U491 (N_491,N_394,N_410);
or U492 (N_492,N_418,N_445);
nor U493 (N_493,N_404,N_423);
and U494 (N_494,N_383,N_427);
or U495 (N_495,N_382,N_396);
and U496 (N_496,N_406,N_428);
and U497 (N_497,N_449,N_447);
nand U498 (N_498,N_393,N_433);
and U499 (N_499,N_417,N_424);
and U500 (N_500,N_381,N_385);
nor U501 (N_501,N_401,N_441);
nor U502 (N_502,N_435,N_442);
and U503 (N_503,N_426,N_393);
nand U504 (N_504,N_413,N_433);
nor U505 (N_505,N_431,N_377);
or U506 (N_506,N_415,N_389);
nand U507 (N_507,N_407,N_398);
nand U508 (N_508,N_396,N_419);
and U509 (N_509,N_418,N_432);
nand U510 (N_510,N_416,N_394);
nand U511 (N_511,N_378,N_384);
nand U512 (N_512,N_383,N_402);
or U513 (N_513,N_442,N_416);
nand U514 (N_514,N_378,N_376);
or U515 (N_515,N_379,N_390);
nand U516 (N_516,N_427,N_447);
and U517 (N_517,N_389,N_417);
nor U518 (N_518,N_417,N_421);
and U519 (N_519,N_445,N_424);
nand U520 (N_520,N_412,N_382);
and U521 (N_521,N_405,N_389);
nand U522 (N_522,N_399,N_445);
and U523 (N_523,N_399,N_423);
or U524 (N_524,N_382,N_415);
or U525 (N_525,N_474,N_460);
or U526 (N_526,N_502,N_517);
and U527 (N_527,N_472,N_512);
and U528 (N_528,N_499,N_467);
and U529 (N_529,N_478,N_506);
xnor U530 (N_530,N_484,N_519);
or U531 (N_531,N_490,N_469);
nor U532 (N_532,N_461,N_508);
or U533 (N_533,N_524,N_462);
or U534 (N_534,N_520,N_488);
and U535 (N_535,N_452,N_471);
and U536 (N_536,N_455,N_498);
and U537 (N_537,N_507,N_513);
nand U538 (N_538,N_494,N_465);
nand U539 (N_539,N_493,N_492);
or U540 (N_540,N_489,N_496);
and U541 (N_541,N_509,N_491);
nor U542 (N_542,N_504,N_516);
or U543 (N_543,N_477,N_453);
or U544 (N_544,N_486,N_495);
nor U545 (N_545,N_523,N_505);
and U546 (N_546,N_468,N_473);
or U547 (N_547,N_500,N_487);
nand U548 (N_548,N_464,N_514);
and U549 (N_549,N_456,N_458);
and U550 (N_550,N_457,N_483);
nand U551 (N_551,N_485,N_475);
and U552 (N_552,N_466,N_503);
and U553 (N_553,N_482,N_521);
nand U554 (N_554,N_501,N_511);
nor U555 (N_555,N_451,N_510);
and U556 (N_556,N_459,N_463);
and U557 (N_557,N_515,N_480);
nand U558 (N_558,N_497,N_479);
or U559 (N_559,N_518,N_522);
and U560 (N_560,N_476,N_454);
and U561 (N_561,N_481,N_450);
or U562 (N_562,N_470,N_496);
and U563 (N_563,N_453,N_515);
nand U564 (N_564,N_455,N_495);
nand U565 (N_565,N_460,N_458);
nor U566 (N_566,N_466,N_508);
or U567 (N_567,N_452,N_479);
nor U568 (N_568,N_462,N_492);
or U569 (N_569,N_490,N_473);
nand U570 (N_570,N_457,N_471);
nor U571 (N_571,N_473,N_521);
or U572 (N_572,N_500,N_460);
xor U573 (N_573,N_506,N_520);
nand U574 (N_574,N_495,N_463);
nand U575 (N_575,N_459,N_471);
and U576 (N_576,N_506,N_461);
nor U577 (N_577,N_516,N_495);
or U578 (N_578,N_509,N_463);
and U579 (N_579,N_513,N_492);
and U580 (N_580,N_515,N_452);
and U581 (N_581,N_456,N_503);
nand U582 (N_582,N_517,N_463);
nor U583 (N_583,N_475,N_488);
nand U584 (N_584,N_456,N_499);
nor U585 (N_585,N_458,N_487);
or U586 (N_586,N_472,N_506);
and U587 (N_587,N_450,N_468);
or U588 (N_588,N_491,N_508);
nand U589 (N_589,N_506,N_468);
and U590 (N_590,N_498,N_501);
nand U591 (N_591,N_514,N_477);
nor U592 (N_592,N_473,N_524);
nor U593 (N_593,N_481,N_470);
or U594 (N_594,N_452,N_485);
and U595 (N_595,N_524,N_455);
nor U596 (N_596,N_456,N_488);
nor U597 (N_597,N_455,N_465);
nand U598 (N_598,N_524,N_486);
and U599 (N_599,N_480,N_455);
nor U600 (N_600,N_566,N_576);
nor U601 (N_601,N_577,N_538);
nand U602 (N_602,N_541,N_567);
or U603 (N_603,N_593,N_547);
nor U604 (N_604,N_580,N_544);
nor U605 (N_605,N_579,N_569);
nand U606 (N_606,N_527,N_531);
nor U607 (N_607,N_546,N_586);
nand U608 (N_608,N_591,N_578);
and U609 (N_609,N_525,N_584);
xnor U610 (N_610,N_583,N_570);
nand U611 (N_611,N_588,N_598);
or U612 (N_612,N_581,N_550);
nand U613 (N_613,N_597,N_534);
or U614 (N_614,N_565,N_554);
nand U615 (N_615,N_543,N_542);
nor U616 (N_616,N_568,N_573);
nor U617 (N_617,N_553,N_529);
nor U618 (N_618,N_552,N_587);
xor U619 (N_619,N_599,N_539);
nor U620 (N_620,N_549,N_557);
nor U621 (N_621,N_537,N_571);
or U622 (N_622,N_564,N_556);
and U623 (N_623,N_536,N_560);
nand U624 (N_624,N_551,N_540);
nand U625 (N_625,N_526,N_595);
and U626 (N_626,N_572,N_555);
nor U627 (N_627,N_548,N_562);
and U628 (N_628,N_535,N_596);
and U629 (N_629,N_589,N_532);
and U630 (N_630,N_563,N_558);
nand U631 (N_631,N_528,N_530);
nand U632 (N_632,N_575,N_545);
and U633 (N_633,N_533,N_590);
nor U634 (N_634,N_592,N_594);
xor U635 (N_635,N_585,N_561);
and U636 (N_636,N_574,N_559);
nor U637 (N_637,N_582,N_570);
and U638 (N_638,N_541,N_529);
or U639 (N_639,N_579,N_577);
nor U640 (N_640,N_550,N_549);
or U641 (N_641,N_565,N_543);
and U642 (N_642,N_578,N_534);
nand U643 (N_643,N_556,N_587);
or U644 (N_644,N_562,N_586);
and U645 (N_645,N_577,N_527);
nor U646 (N_646,N_550,N_585);
xnor U647 (N_647,N_560,N_544);
nor U648 (N_648,N_571,N_531);
nor U649 (N_649,N_576,N_578);
or U650 (N_650,N_591,N_542);
or U651 (N_651,N_592,N_529);
xor U652 (N_652,N_543,N_589);
nand U653 (N_653,N_544,N_533);
or U654 (N_654,N_534,N_544);
and U655 (N_655,N_589,N_538);
or U656 (N_656,N_587,N_541);
nor U657 (N_657,N_546,N_548);
and U658 (N_658,N_552,N_597);
or U659 (N_659,N_583,N_549);
and U660 (N_660,N_575,N_549);
nor U661 (N_661,N_568,N_599);
or U662 (N_662,N_573,N_536);
nand U663 (N_663,N_567,N_574);
nor U664 (N_664,N_559,N_588);
and U665 (N_665,N_533,N_553);
and U666 (N_666,N_552,N_599);
nor U667 (N_667,N_575,N_597);
xnor U668 (N_668,N_566,N_555);
and U669 (N_669,N_575,N_525);
xnor U670 (N_670,N_525,N_545);
nand U671 (N_671,N_561,N_571);
nor U672 (N_672,N_568,N_529);
and U673 (N_673,N_534,N_592);
nor U674 (N_674,N_525,N_592);
nand U675 (N_675,N_653,N_644);
nand U676 (N_676,N_612,N_643);
or U677 (N_677,N_632,N_636);
nor U678 (N_678,N_648,N_624);
and U679 (N_679,N_618,N_659);
nor U680 (N_680,N_608,N_656);
nand U681 (N_681,N_664,N_646);
nor U682 (N_682,N_621,N_652);
nand U683 (N_683,N_671,N_665);
nor U684 (N_684,N_606,N_668);
and U685 (N_685,N_601,N_610);
xnor U686 (N_686,N_633,N_672);
nor U687 (N_687,N_640,N_611);
nor U688 (N_688,N_666,N_645);
and U689 (N_689,N_634,N_670);
nor U690 (N_690,N_667,N_649);
or U691 (N_691,N_655,N_658);
and U692 (N_692,N_669,N_663);
nor U693 (N_693,N_625,N_660);
or U694 (N_694,N_674,N_637);
nor U695 (N_695,N_613,N_615);
and U696 (N_696,N_604,N_673);
nor U697 (N_697,N_635,N_616);
nand U698 (N_698,N_657,N_605);
and U699 (N_699,N_647,N_602);
nand U700 (N_700,N_614,N_650);
or U701 (N_701,N_627,N_641);
nand U702 (N_702,N_617,N_622);
or U703 (N_703,N_623,N_661);
or U704 (N_704,N_662,N_609);
or U705 (N_705,N_654,N_600);
and U706 (N_706,N_603,N_607);
nor U707 (N_707,N_628,N_630);
and U708 (N_708,N_626,N_620);
nand U709 (N_709,N_651,N_638);
or U710 (N_710,N_631,N_629);
xor U711 (N_711,N_642,N_639);
and U712 (N_712,N_619,N_647);
or U713 (N_713,N_644,N_629);
nor U714 (N_714,N_639,N_647);
nor U715 (N_715,N_662,N_659);
and U716 (N_716,N_635,N_664);
and U717 (N_717,N_650,N_663);
xnor U718 (N_718,N_619,N_646);
or U719 (N_719,N_627,N_672);
or U720 (N_720,N_656,N_604);
xnor U721 (N_721,N_663,N_619);
or U722 (N_722,N_645,N_658);
nor U723 (N_723,N_610,N_646);
nor U724 (N_724,N_629,N_673);
nor U725 (N_725,N_647,N_642);
nor U726 (N_726,N_667,N_604);
nor U727 (N_727,N_651,N_611);
nor U728 (N_728,N_635,N_646);
and U729 (N_729,N_644,N_643);
and U730 (N_730,N_617,N_673);
or U731 (N_731,N_673,N_650);
and U732 (N_732,N_626,N_647);
nor U733 (N_733,N_600,N_602);
xnor U734 (N_734,N_617,N_656);
nor U735 (N_735,N_624,N_639);
or U736 (N_736,N_610,N_609);
nor U737 (N_737,N_645,N_617);
or U738 (N_738,N_646,N_605);
and U739 (N_739,N_611,N_608);
nor U740 (N_740,N_669,N_602);
or U741 (N_741,N_663,N_622);
nand U742 (N_742,N_631,N_621);
and U743 (N_743,N_671,N_642);
nor U744 (N_744,N_621,N_646);
nand U745 (N_745,N_649,N_615);
nand U746 (N_746,N_622,N_653);
or U747 (N_747,N_635,N_604);
and U748 (N_748,N_613,N_623);
and U749 (N_749,N_630,N_655);
nand U750 (N_750,N_734,N_710);
and U751 (N_751,N_700,N_706);
nand U752 (N_752,N_685,N_748);
or U753 (N_753,N_695,N_686);
nand U754 (N_754,N_737,N_716);
and U755 (N_755,N_677,N_688);
nor U756 (N_756,N_684,N_738);
and U757 (N_757,N_736,N_744);
nand U758 (N_758,N_701,N_742);
nand U759 (N_759,N_683,N_733);
nand U760 (N_760,N_715,N_735);
xor U761 (N_761,N_722,N_709);
nor U762 (N_762,N_718,N_717);
or U763 (N_763,N_681,N_689);
nor U764 (N_764,N_729,N_679);
nand U765 (N_765,N_714,N_699);
nand U766 (N_766,N_678,N_711);
nor U767 (N_767,N_720,N_708);
and U768 (N_768,N_676,N_746);
and U769 (N_769,N_694,N_697);
and U770 (N_770,N_713,N_731);
or U771 (N_771,N_704,N_707);
and U772 (N_772,N_728,N_705);
or U773 (N_773,N_682,N_691);
or U774 (N_774,N_721,N_696);
nand U775 (N_775,N_745,N_743);
nand U776 (N_776,N_712,N_702);
and U777 (N_777,N_740,N_727);
and U778 (N_778,N_724,N_725);
nor U779 (N_779,N_732,N_692);
and U780 (N_780,N_680,N_693);
or U781 (N_781,N_747,N_690);
nor U782 (N_782,N_675,N_719);
or U783 (N_783,N_739,N_698);
or U784 (N_784,N_703,N_687);
nand U785 (N_785,N_726,N_723);
or U786 (N_786,N_749,N_741);
or U787 (N_787,N_730,N_692);
or U788 (N_788,N_706,N_732);
nor U789 (N_789,N_733,N_694);
or U790 (N_790,N_678,N_714);
nor U791 (N_791,N_746,N_725);
or U792 (N_792,N_706,N_679);
nor U793 (N_793,N_730,N_745);
or U794 (N_794,N_685,N_722);
nor U795 (N_795,N_695,N_740);
nor U796 (N_796,N_743,N_725);
or U797 (N_797,N_689,N_715);
and U798 (N_798,N_697,N_706);
or U799 (N_799,N_731,N_741);
and U800 (N_800,N_677,N_724);
nor U801 (N_801,N_714,N_731);
nor U802 (N_802,N_707,N_695);
nand U803 (N_803,N_694,N_735);
xnor U804 (N_804,N_743,N_720);
and U805 (N_805,N_699,N_717);
and U806 (N_806,N_679,N_687);
nor U807 (N_807,N_738,N_683);
and U808 (N_808,N_681,N_744);
nor U809 (N_809,N_722,N_737);
or U810 (N_810,N_701,N_713);
and U811 (N_811,N_726,N_713);
nand U812 (N_812,N_683,N_743);
or U813 (N_813,N_699,N_723);
nor U814 (N_814,N_680,N_719);
nand U815 (N_815,N_729,N_722);
nand U816 (N_816,N_698,N_694);
and U817 (N_817,N_729,N_744);
nand U818 (N_818,N_699,N_688);
nand U819 (N_819,N_748,N_732);
and U820 (N_820,N_695,N_678);
xnor U821 (N_821,N_711,N_717);
nand U822 (N_822,N_701,N_703);
and U823 (N_823,N_749,N_706);
or U824 (N_824,N_736,N_686);
and U825 (N_825,N_754,N_758);
nor U826 (N_826,N_770,N_813);
xor U827 (N_827,N_784,N_816);
nor U828 (N_828,N_802,N_760);
nand U829 (N_829,N_771,N_804);
xnor U830 (N_830,N_791,N_801);
or U831 (N_831,N_785,N_778);
nor U832 (N_832,N_756,N_795);
or U833 (N_833,N_798,N_788);
nor U834 (N_834,N_805,N_768);
nand U835 (N_835,N_777,N_815);
and U836 (N_836,N_794,N_790);
and U837 (N_837,N_774,N_799);
nand U838 (N_838,N_766,N_807);
nand U839 (N_839,N_789,N_757);
and U840 (N_840,N_759,N_765);
nor U841 (N_841,N_773,N_817);
nand U842 (N_842,N_796,N_786);
and U843 (N_843,N_776,N_814);
or U844 (N_844,N_767,N_811);
and U845 (N_845,N_810,N_803);
or U846 (N_846,N_762,N_822);
and U847 (N_847,N_809,N_797);
or U848 (N_848,N_793,N_824);
and U849 (N_849,N_818,N_800);
nor U850 (N_850,N_752,N_769);
and U851 (N_851,N_820,N_780);
and U852 (N_852,N_812,N_763);
and U853 (N_853,N_823,N_751);
nor U854 (N_854,N_819,N_781);
or U855 (N_855,N_750,N_792);
and U856 (N_856,N_821,N_782);
or U857 (N_857,N_761,N_806);
nand U858 (N_858,N_775,N_779);
nor U859 (N_859,N_753,N_772);
and U860 (N_860,N_787,N_783);
nor U861 (N_861,N_764,N_808);
and U862 (N_862,N_755,N_766);
nand U863 (N_863,N_760,N_750);
and U864 (N_864,N_760,N_774);
and U865 (N_865,N_767,N_750);
xnor U866 (N_866,N_820,N_751);
or U867 (N_867,N_816,N_801);
or U868 (N_868,N_790,N_798);
and U869 (N_869,N_766,N_758);
and U870 (N_870,N_796,N_776);
nor U871 (N_871,N_804,N_806);
xnor U872 (N_872,N_771,N_759);
nand U873 (N_873,N_795,N_810);
nor U874 (N_874,N_805,N_793);
nand U875 (N_875,N_792,N_761);
nand U876 (N_876,N_750,N_818);
or U877 (N_877,N_764,N_762);
and U878 (N_878,N_820,N_775);
or U879 (N_879,N_750,N_791);
and U880 (N_880,N_811,N_778);
and U881 (N_881,N_810,N_752);
nand U882 (N_882,N_756,N_761);
xnor U883 (N_883,N_811,N_759);
and U884 (N_884,N_755,N_767);
and U885 (N_885,N_780,N_791);
nand U886 (N_886,N_770,N_750);
nand U887 (N_887,N_811,N_750);
or U888 (N_888,N_823,N_787);
and U889 (N_889,N_794,N_797);
nand U890 (N_890,N_770,N_765);
or U891 (N_891,N_791,N_777);
and U892 (N_892,N_822,N_754);
nor U893 (N_893,N_803,N_765);
and U894 (N_894,N_779,N_798);
or U895 (N_895,N_752,N_764);
xor U896 (N_896,N_778,N_812);
or U897 (N_897,N_762,N_774);
nor U898 (N_898,N_768,N_810);
or U899 (N_899,N_817,N_807);
and U900 (N_900,N_892,N_849);
nand U901 (N_901,N_875,N_825);
or U902 (N_902,N_836,N_827);
and U903 (N_903,N_887,N_898);
nand U904 (N_904,N_869,N_839);
and U905 (N_905,N_840,N_896);
nand U906 (N_906,N_854,N_856);
nor U907 (N_907,N_890,N_837);
and U908 (N_908,N_883,N_845);
nor U909 (N_909,N_880,N_895);
and U910 (N_910,N_860,N_888);
or U911 (N_911,N_865,N_833);
nor U912 (N_912,N_870,N_864);
nor U913 (N_913,N_829,N_866);
or U914 (N_914,N_832,N_847);
or U915 (N_915,N_867,N_861);
or U916 (N_916,N_835,N_873);
nand U917 (N_917,N_826,N_876);
nand U918 (N_918,N_834,N_885);
xnor U919 (N_919,N_882,N_862);
nand U920 (N_920,N_848,N_863);
and U921 (N_921,N_846,N_841);
and U922 (N_922,N_853,N_844);
nor U923 (N_923,N_838,N_828);
or U924 (N_924,N_843,N_881);
nor U925 (N_925,N_852,N_855);
and U926 (N_926,N_874,N_899);
nor U927 (N_927,N_886,N_859);
nand U928 (N_928,N_894,N_842);
and U929 (N_929,N_877,N_893);
or U930 (N_930,N_857,N_831);
or U931 (N_931,N_858,N_878);
or U932 (N_932,N_897,N_871);
nor U933 (N_933,N_830,N_884);
xor U934 (N_934,N_889,N_872);
and U935 (N_935,N_850,N_868);
or U936 (N_936,N_891,N_851);
and U937 (N_937,N_879,N_838);
nor U938 (N_938,N_852,N_836);
or U939 (N_939,N_827,N_852);
nor U940 (N_940,N_884,N_829);
and U941 (N_941,N_897,N_856);
nor U942 (N_942,N_860,N_825);
xor U943 (N_943,N_841,N_827);
and U944 (N_944,N_860,N_867);
nand U945 (N_945,N_869,N_875);
nor U946 (N_946,N_850,N_872);
or U947 (N_947,N_885,N_867);
nand U948 (N_948,N_844,N_866);
nand U949 (N_949,N_828,N_850);
nand U950 (N_950,N_831,N_854);
nand U951 (N_951,N_857,N_867);
and U952 (N_952,N_856,N_862);
nand U953 (N_953,N_834,N_879);
nand U954 (N_954,N_852,N_826);
nand U955 (N_955,N_846,N_891);
nor U956 (N_956,N_831,N_860);
nor U957 (N_957,N_852,N_849);
or U958 (N_958,N_831,N_874);
or U959 (N_959,N_841,N_870);
and U960 (N_960,N_877,N_884);
and U961 (N_961,N_888,N_868);
nand U962 (N_962,N_873,N_880);
or U963 (N_963,N_827,N_846);
and U964 (N_964,N_895,N_835);
and U965 (N_965,N_829,N_891);
nand U966 (N_966,N_861,N_829);
nor U967 (N_967,N_854,N_842);
and U968 (N_968,N_884,N_864);
nand U969 (N_969,N_872,N_888);
nor U970 (N_970,N_894,N_836);
or U971 (N_971,N_886,N_831);
and U972 (N_972,N_863,N_868);
nor U973 (N_973,N_879,N_851);
nand U974 (N_974,N_890,N_861);
nand U975 (N_975,N_911,N_926);
nand U976 (N_976,N_946,N_922);
or U977 (N_977,N_939,N_950);
and U978 (N_978,N_940,N_963);
nor U979 (N_979,N_923,N_912);
nand U980 (N_980,N_945,N_942);
or U981 (N_981,N_902,N_930);
nand U982 (N_982,N_970,N_925);
nor U983 (N_983,N_948,N_944);
and U984 (N_984,N_968,N_924);
or U985 (N_985,N_907,N_933);
nand U986 (N_986,N_938,N_953);
nand U987 (N_987,N_960,N_969);
xor U988 (N_988,N_956,N_931);
and U989 (N_989,N_958,N_949);
and U990 (N_990,N_962,N_967);
nand U991 (N_991,N_959,N_951);
or U992 (N_992,N_919,N_965);
nand U993 (N_993,N_928,N_900);
and U994 (N_994,N_916,N_901);
or U995 (N_995,N_934,N_961);
and U996 (N_996,N_908,N_914);
nand U997 (N_997,N_910,N_905);
and U998 (N_998,N_941,N_909);
and U999 (N_999,N_906,N_937);
and U1000 (N_1000,N_915,N_920);
or U1001 (N_1001,N_932,N_927);
nand U1002 (N_1002,N_964,N_974);
nand U1003 (N_1003,N_936,N_973);
and U1004 (N_1004,N_918,N_972);
or U1005 (N_1005,N_952,N_935);
nand U1006 (N_1006,N_971,N_955);
nor U1007 (N_1007,N_903,N_904);
nand U1008 (N_1008,N_947,N_917);
nand U1009 (N_1009,N_954,N_913);
or U1010 (N_1010,N_929,N_957);
and U1011 (N_1011,N_943,N_966);
and U1012 (N_1012,N_921,N_918);
or U1013 (N_1013,N_955,N_932);
and U1014 (N_1014,N_900,N_971);
nand U1015 (N_1015,N_926,N_913);
or U1016 (N_1016,N_936,N_904);
nand U1017 (N_1017,N_960,N_974);
nand U1018 (N_1018,N_955,N_930);
and U1019 (N_1019,N_961,N_922);
nand U1020 (N_1020,N_968,N_963);
nor U1021 (N_1021,N_939,N_945);
or U1022 (N_1022,N_954,N_968);
xor U1023 (N_1023,N_974,N_946);
or U1024 (N_1024,N_914,N_959);
nand U1025 (N_1025,N_959,N_950);
and U1026 (N_1026,N_971,N_944);
or U1027 (N_1027,N_908,N_939);
and U1028 (N_1028,N_916,N_971);
nor U1029 (N_1029,N_908,N_960);
and U1030 (N_1030,N_955,N_938);
or U1031 (N_1031,N_958,N_973);
nand U1032 (N_1032,N_906,N_968);
nand U1033 (N_1033,N_917,N_916);
and U1034 (N_1034,N_941,N_925);
nor U1035 (N_1035,N_937,N_934);
and U1036 (N_1036,N_901,N_944);
nor U1037 (N_1037,N_958,N_902);
nor U1038 (N_1038,N_913,N_929);
nand U1039 (N_1039,N_942,N_903);
nor U1040 (N_1040,N_906,N_907);
and U1041 (N_1041,N_912,N_971);
and U1042 (N_1042,N_906,N_971);
nand U1043 (N_1043,N_935,N_914);
xor U1044 (N_1044,N_955,N_966);
or U1045 (N_1045,N_932,N_951);
nor U1046 (N_1046,N_949,N_903);
or U1047 (N_1047,N_912,N_947);
xor U1048 (N_1048,N_964,N_973);
or U1049 (N_1049,N_961,N_963);
nand U1050 (N_1050,N_1043,N_1041);
and U1051 (N_1051,N_1029,N_982);
and U1052 (N_1052,N_1003,N_1031);
and U1053 (N_1053,N_1023,N_1010);
nand U1054 (N_1054,N_1048,N_985);
and U1055 (N_1055,N_1024,N_996);
nor U1056 (N_1056,N_990,N_1033);
nand U1057 (N_1057,N_997,N_999);
or U1058 (N_1058,N_1005,N_1047);
nor U1059 (N_1059,N_986,N_1007);
or U1060 (N_1060,N_1019,N_1008);
and U1061 (N_1061,N_1020,N_975);
nand U1062 (N_1062,N_1036,N_1034);
and U1063 (N_1063,N_1017,N_1037);
or U1064 (N_1064,N_1038,N_1045);
xnor U1065 (N_1065,N_991,N_998);
or U1066 (N_1066,N_1049,N_1012);
nor U1067 (N_1067,N_995,N_1044);
nor U1068 (N_1068,N_1039,N_1015);
or U1069 (N_1069,N_1000,N_1013);
nor U1070 (N_1070,N_1006,N_989);
and U1071 (N_1071,N_1025,N_979);
or U1072 (N_1072,N_976,N_1016);
nor U1073 (N_1073,N_987,N_980);
nand U1074 (N_1074,N_1018,N_1032);
nand U1075 (N_1075,N_1004,N_983);
and U1076 (N_1076,N_1042,N_994);
or U1077 (N_1077,N_1001,N_988);
nor U1078 (N_1078,N_978,N_1046);
and U1079 (N_1079,N_1002,N_1014);
nor U1080 (N_1080,N_1011,N_992);
nor U1081 (N_1081,N_1035,N_1021);
and U1082 (N_1082,N_1028,N_1022);
nor U1083 (N_1083,N_981,N_1027);
or U1084 (N_1084,N_993,N_1026);
or U1085 (N_1085,N_977,N_1009);
nor U1086 (N_1086,N_984,N_1040);
nor U1087 (N_1087,N_1030,N_983);
nor U1088 (N_1088,N_1045,N_1010);
and U1089 (N_1089,N_1015,N_976);
and U1090 (N_1090,N_1032,N_1030);
and U1091 (N_1091,N_1035,N_988);
nand U1092 (N_1092,N_990,N_1048);
nor U1093 (N_1093,N_1026,N_1045);
xnor U1094 (N_1094,N_1005,N_992);
and U1095 (N_1095,N_997,N_1039);
and U1096 (N_1096,N_1020,N_1014);
or U1097 (N_1097,N_1025,N_1049);
nor U1098 (N_1098,N_1030,N_1045);
and U1099 (N_1099,N_1006,N_978);
or U1100 (N_1100,N_1037,N_1000);
or U1101 (N_1101,N_1010,N_998);
nor U1102 (N_1102,N_1027,N_988);
and U1103 (N_1103,N_991,N_1037);
nor U1104 (N_1104,N_1049,N_985);
or U1105 (N_1105,N_1042,N_1029);
and U1106 (N_1106,N_1041,N_1011);
nor U1107 (N_1107,N_982,N_1018);
or U1108 (N_1108,N_1019,N_1000);
or U1109 (N_1109,N_1028,N_991);
nor U1110 (N_1110,N_1048,N_979);
nand U1111 (N_1111,N_1039,N_982);
and U1112 (N_1112,N_1000,N_990);
or U1113 (N_1113,N_983,N_1018);
nand U1114 (N_1114,N_1042,N_1001);
nand U1115 (N_1115,N_1010,N_1026);
nor U1116 (N_1116,N_976,N_987);
xor U1117 (N_1117,N_1001,N_1002);
and U1118 (N_1118,N_1040,N_1029);
and U1119 (N_1119,N_1026,N_989);
nand U1120 (N_1120,N_1043,N_1009);
and U1121 (N_1121,N_1006,N_982);
nor U1122 (N_1122,N_1017,N_1016);
and U1123 (N_1123,N_986,N_1043);
nor U1124 (N_1124,N_1027,N_994);
and U1125 (N_1125,N_1100,N_1070);
or U1126 (N_1126,N_1072,N_1092);
nand U1127 (N_1127,N_1071,N_1054);
nor U1128 (N_1128,N_1085,N_1109);
nor U1129 (N_1129,N_1051,N_1050);
nand U1130 (N_1130,N_1115,N_1124);
and U1131 (N_1131,N_1069,N_1056);
nor U1132 (N_1132,N_1113,N_1061);
or U1133 (N_1133,N_1063,N_1053);
or U1134 (N_1134,N_1097,N_1060);
nor U1135 (N_1135,N_1062,N_1108);
or U1136 (N_1136,N_1084,N_1103);
nand U1137 (N_1137,N_1102,N_1078);
and U1138 (N_1138,N_1101,N_1067);
nor U1139 (N_1139,N_1119,N_1118);
and U1140 (N_1140,N_1088,N_1089);
nor U1141 (N_1141,N_1120,N_1095);
or U1142 (N_1142,N_1117,N_1066);
nand U1143 (N_1143,N_1075,N_1091);
or U1144 (N_1144,N_1074,N_1064);
or U1145 (N_1145,N_1082,N_1107);
nand U1146 (N_1146,N_1055,N_1099);
or U1147 (N_1147,N_1110,N_1094);
nor U1148 (N_1148,N_1111,N_1058);
and U1149 (N_1149,N_1093,N_1122);
and U1150 (N_1150,N_1096,N_1080);
nor U1151 (N_1151,N_1098,N_1057);
and U1152 (N_1152,N_1077,N_1104);
or U1153 (N_1153,N_1090,N_1076);
and U1154 (N_1154,N_1083,N_1106);
nor U1155 (N_1155,N_1116,N_1114);
xor U1156 (N_1156,N_1087,N_1073);
and U1157 (N_1157,N_1065,N_1112);
or U1158 (N_1158,N_1052,N_1079);
and U1159 (N_1159,N_1086,N_1123);
or U1160 (N_1160,N_1081,N_1105);
nor U1161 (N_1161,N_1059,N_1121);
or U1162 (N_1162,N_1068,N_1120);
and U1163 (N_1163,N_1093,N_1059);
nand U1164 (N_1164,N_1123,N_1058);
and U1165 (N_1165,N_1110,N_1080);
and U1166 (N_1166,N_1110,N_1101);
nand U1167 (N_1167,N_1073,N_1070);
and U1168 (N_1168,N_1076,N_1087);
or U1169 (N_1169,N_1059,N_1083);
nor U1170 (N_1170,N_1117,N_1120);
nor U1171 (N_1171,N_1053,N_1114);
or U1172 (N_1172,N_1058,N_1122);
or U1173 (N_1173,N_1059,N_1114);
or U1174 (N_1174,N_1076,N_1086);
nor U1175 (N_1175,N_1081,N_1106);
nand U1176 (N_1176,N_1073,N_1100);
and U1177 (N_1177,N_1109,N_1099);
and U1178 (N_1178,N_1074,N_1062);
or U1179 (N_1179,N_1069,N_1050);
and U1180 (N_1180,N_1065,N_1061);
and U1181 (N_1181,N_1074,N_1097);
nand U1182 (N_1182,N_1123,N_1075);
and U1183 (N_1183,N_1095,N_1101);
nand U1184 (N_1184,N_1064,N_1066);
nor U1185 (N_1185,N_1089,N_1069);
nand U1186 (N_1186,N_1121,N_1057);
xor U1187 (N_1187,N_1081,N_1059);
nor U1188 (N_1188,N_1077,N_1115);
nor U1189 (N_1189,N_1052,N_1069);
nand U1190 (N_1190,N_1106,N_1086);
or U1191 (N_1191,N_1106,N_1070);
nor U1192 (N_1192,N_1112,N_1069);
and U1193 (N_1193,N_1052,N_1082);
or U1194 (N_1194,N_1123,N_1068);
or U1195 (N_1195,N_1069,N_1108);
and U1196 (N_1196,N_1069,N_1095);
nand U1197 (N_1197,N_1102,N_1064);
nand U1198 (N_1198,N_1051,N_1052);
nand U1199 (N_1199,N_1097,N_1103);
or U1200 (N_1200,N_1176,N_1141);
nor U1201 (N_1201,N_1171,N_1189);
nand U1202 (N_1202,N_1148,N_1151);
or U1203 (N_1203,N_1193,N_1129);
nor U1204 (N_1204,N_1144,N_1139);
nor U1205 (N_1205,N_1132,N_1172);
nand U1206 (N_1206,N_1184,N_1138);
nor U1207 (N_1207,N_1149,N_1175);
nand U1208 (N_1208,N_1192,N_1170);
and U1209 (N_1209,N_1196,N_1190);
nor U1210 (N_1210,N_1186,N_1197);
and U1211 (N_1211,N_1162,N_1147);
nand U1212 (N_1212,N_1153,N_1167);
and U1213 (N_1213,N_1159,N_1187);
and U1214 (N_1214,N_1150,N_1152);
nand U1215 (N_1215,N_1191,N_1163);
nor U1216 (N_1216,N_1142,N_1194);
nor U1217 (N_1217,N_1181,N_1155);
nand U1218 (N_1218,N_1134,N_1168);
and U1219 (N_1219,N_1140,N_1156);
or U1220 (N_1220,N_1165,N_1195);
nand U1221 (N_1221,N_1157,N_1131);
nor U1222 (N_1222,N_1128,N_1135);
nand U1223 (N_1223,N_1178,N_1161);
nor U1224 (N_1224,N_1164,N_1133);
or U1225 (N_1225,N_1137,N_1160);
or U1226 (N_1226,N_1180,N_1125);
or U1227 (N_1227,N_1174,N_1126);
nor U1228 (N_1228,N_1127,N_1173);
and U1229 (N_1229,N_1130,N_1185);
and U1230 (N_1230,N_1143,N_1154);
and U1231 (N_1231,N_1177,N_1188);
nand U1232 (N_1232,N_1183,N_1146);
xor U1233 (N_1233,N_1158,N_1166);
or U1234 (N_1234,N_1199,N_1169);
nor U1235 (N_1235,N_1145,N_1182);
or U1236 (N_1236,N_1198,N_1136);
xnor U1237 (N_1237,N_1179,N_1178);
and U1238 (N_1238,N_1146,N_1136);
or U1239 (N_1239,N_1164,N_1126);
nand U1240 (N_1240,N_1133,N_1125);
nand U1241 (N_1241,N_1127,N_1147);
nand U1242 (N_1242,N_1128,N_1160);
nor U1243 (N_1243,N_1132,N_1193);
nand U1244 (N_1244,N_1174,N_1155);
and U1245 (N_1245,N_1172,N_1150);
or U1246 (N_1246,N_1182,N_1178);
nor U1247 (N_1247,N_1137,N_1140);
or U1248 (N_1248,N_1136,N_1129);
or U1249 (N_1249,N_1157,N_1137);
nand U1250 (N_1250,N_1164,N_1179);
or U1251 (N_1251,N_1140,N_1129);
and U1252 (N_1252,N_1152,N_1196);
or U1253 (N_1253,N_1184,N_1135);
nor U1254 (N_1254,N_1136,N_1181);
or U1255 (N_1255,N_1132,N_1159);
and U1256 (N_1256,N_1198,N_1137);
nor U1257 (N_1257,N_1151,N_1141);
and U1258 (N_1258,N_1157,N_1175);
nand U1259 (N_1259,N_1198,N_1163);
nor U1260 (N_1260,N_1135,N_1194);
and U1261 (N_1261,N_1166,N_1155);
nand U1262 (N_1262,N_1169,N_1193);
and U1263 (N_1263,N_1163,N_1129);
and U1264 (N_1264,N_1133,N_1185);
and U1265 (N_1265,N_1129,N_1130);
nor U1266 (N_1266,N_1160,N_1154);
nor U1267 (N_1267,N_1192,N_1126);
nor U1268 (N_1268,N_1197,N_1155);
nand U1269 (N_1269,N_1180,N_1127);
or U1270 (N_1270,N_1150,N_1180);
nor U1271 (N_1271,N_1178,N_1196);
nor U1272 (N_1272,N_1158,N_1157);
nor U1273 (N_1273,N_1188,N_1138);
and U1274 (N_1274,N_1177,N_1139);
and U1275 (N_1275,N_1202,N_1236);
or U1276 (N_1276,N_1271,N_1247);
or U1277 (N_1277,N_1246,N_1257);
nand U1278 (N_1278,N_1266,N_1217);
nor U1279 (N_1279,N_1237,N_1212);
and U1280 (N_1280,N_1260,N_1208);
and U1281 (N_1281,N_1225,N_1258);
and U1282 (N_1282,N_1223,N_1262);
or U1283 (N_1283,N_1221,N_1245);
nand U1284 (N_1284,N_1209,N_1235);
or U1285 (N_1285,N_1205,N_1268);
or U1286 (N_1286,N_1244,N_1249);
and U1287 (N_1287,N_1255,N_1252);
nand U1288 (N_1288,N_1238,N_1259);
or U1289 (N_1289,N_1211,N_1233);
or U1290 (N_1290,N_1256,N_1272);
nor U1291 (N_1291,N_1261,N_1269);
or U1292 (N_1292,N_1216,N_1273);
nor U1293 (N_1293,N_1206,N_1253);
or U1294 (N_1294,N_1274,N_1222);
nor U1295 (N_1295,N_1215,N_1239);
or U1296 (N_1296,N_1241,N_1232);
nand U1297 (N_1297,N_1254,N_1220);
nand U1298 (N_1298,N_1219,N_1270);
or U1299 (N_1299,N_1226,N_1200);
and U1300 (N_1300,N_1230,N_1204);
nand U1301 (N_1301,N_1242,N_1207);
and U1302 (N_1302,N_1265,N_1213);
or U1303 (N_1303,N_1229,N_1201);
nor U1304 (N_1304,N_1243,N_1224);
nand U1305 (N_1305,N_1263,N_1248);
nand U1306 (N_1306,N_1267,N_1214);
nor U1307 (N_1307,N_1250,N_1264);
nand U1308 (N_1308,N_1234,N_1210);
nand U1309 (N_1309,N_1203,N_1231);
nand U1310 (N_1310,N_1240,N_1228);
nor U1311 (N_1311,N_1227,N_1218);
nand U1312 (N_1312,N_1251,N_1200);
or U1313 (N_1313,N_1265,N_1271);
and U1314 (N_1314,N_1268,N_1217);
nand U1315 (N_1315,N_1205,N_1207);
nand U1316 (N_1316,N_1265,N_1223);
nand U1317 (N_1317,N_1206,N_1261);
nand U1318 (N_1318,N_1262,N_1204);
nand U1319 (N_1319,N_1231,N_1246);
and U1320 (N_1320,N_1200,N_1259);
nor U1321 (N_1321,N_1251,N_1250);
nand U1322 (N_1322,N_1251,N_1213);
nand U1323 (N_1323,N_1211,N_1201);
and U1324 (N_1324,N_1233,N_1263);
nor U1325 (N_1325,N_1266,N_1226);
nor U1326 (N_1326,N_1223,N_1231);
nor U1327 (N_1327,N_1257,N_1266);
nor U1328 (N_1328,N_1223,N_1242);
nor U1329 (N_1329,N_1209,N_1272);
nor U1330 (N_1330,N_1226,N_1268);
nand U1331 (N_1331,N_1251,N_1240);
and U1332 (N_1332,N_1229,N_1273);
and U1333 (N_1333,N_1213,N_1254);
nand U1334 (N_1334,N_1257,N_1260);
or U1335 (N_1335,N_1235,N_1207);
or U1336 (N_1336,N_1222,N_1242);
and U1337 (N_1337,N_1250,N_1231);
or U1338 (N_1338,N_1264,N_1271);
or U1339 (N_1339,N_1207,N_1216);
and U1340 (N_1340,N_1249,N_1224);
nand U1341 (N_1341,N_1211,N_1229);
nand U1342 (N_1342,N_1258,N_1249);
or U1343 (N_1343,N_1254,N_1203);
and U1344 (N_1344,N_1224,N_1251);
and U1345 (N_1345,N_1241,N_1212);
or U1346 (N_1346,N_1241,N_1273);
or U1347 (N_1347,N_1257,N_1242);
and U1348 (N_1348,N_1248,N_1242);
nand U1349 (N_1349,N_1235,N_1254);
nand U1350 (N_1350,N_1312,N_1310);
nor U1351 (N_1351,N_1342,N_1311);
and U1352 (N_1352,N_1283,N_1331);
nand U1353 (N_1353,N_1302,N_1287);
nor U1354 (N_1354,N_1316,N_1275);
and U1355 (N_1355,N_1319,N_1345);
nor U1356 (N_1356,N_1299,N_1346);
nand U1357 (N_1357,N_1315,N_1300);
or U1358 (N_1358,N_1286,N_1307);
and U1359 (N_1359,N_1320,N_1292);
nand U1360 (N_1360,N_1303,N_1308);
nand U1361 (N_1361,N_1289,N_1340);
nand U1362 (N_1362,N_1278,N_1277);
or U1363 (N_1363,N_1306,N_1334);
nor U1364 (N_1364,N_1317,N_1294);
and U1365 (N_1365,N_1322,N_1276);
and U1366 (N_1366,N_1305,N_1296);
nand U1367 (N_1367,N_1281,N_1328);
or U1368 (N_1368,N_1326,N_1347);
nor U1369 (N_1369,N_1343,N_1309);
nand U1370 (N_1370,N_1332,N_1344);
nand U1371 (N_1371,N_1291,N_1327);
and U1372 (N_1372,N_1293,N_1333);
nor U1373 (N_1373,N_1325,N_1336);
or U1374 (N_1374,N_1297,N_1330);
nor U1375 (N_1375,N_1324,N_1339);
nand U1376 (N_1376,N_1338,N_1335);
nand U1377 (N_1377,N_1304,N_1282);
xor U1378 (N_1378,N_1337,N_1290);
nor U1379 (N_1379,N_1280,N_1285);
or U1380 (N_1380,N_1329,N_1314);
and U1381 (N_1381,N_1301,N_1288);
nand U1382 (N_1382,N_1321,N_1341);
and U1383 (N_1383,N_1295,N_1348);
or U1384 (N_1384,N_1298,N_1313);
and U1385 (N_1385,N_1318,N_1349);
nand U1386 (N_1386,N_1279,N_1284);
nor U1387 (N_1387,N_1323,N_1292);
and U1388 (N_1388,N_1342,N_1326);
or U1389 (N_1389,N_1310,N_1322);
and U1390 (N_1390,N_1340,N_1329);
nand U1391 (N_1391,N_1332,N_1348);
or U1392 (N_1392,N_1284,N_1287);
nor U1393 (N_1393,N_1297,N_1344);
and U1394 (N_1394,N_1287,N_1300);
nor U1395 (N_1395,N_1297,N_1335);
or U1396 (N_1396,N_1341,N_1298);
nand U1397 (N_1397,N_1277,N_1318);
nor U1398 (N_1398,N_1336,N_1324);
or U1399 (N_1399,N_1281,N_1295);
nand U1400 (N_1400,N_1294,N_1285);
or U1401 (N_1401,N_1276,N_1303);
or U1402 (N_1402,N_1336,N_1347);
nor U1403 (N_1403,N_1310,N_1317);
or U1404 (N_1404,N_1292,N_1312);
or U1405 (N_1405,N_1280,N_1334);
nand U1406 (N_1406,N_1285,N_1331);
or U1407 (N_1407,N_1277,N_1283);
nor U1408 (N_1408,N_1279,N_1297);
nand U1409 (N_1409,N_1303,N_1285);
nor U1410 (N_1410,N_1344,N_1296);
nand U1411 (N_1411,N_1286,N_1301);
nor U1412 (N_1412,N_1342,N_1338);
and U1413 (N_1413,N_1342,N_1294);
or U1414 (N_1414,N_1330,N_1333);
nand U1415 (N_1415,N_1331,N_1314);
nand U1416 (N_1416,N_1281,N_1326);
nor U1417 (N_1417,N_1328,N_1345);
nand U1418 (N_1418,N_1296,N_1286);
nand U1419 (N_1419,N_1300,N_1323);
nand U1420 (N_1420,N_1322,N_1314);
or U1421 (N_1421,N_1328,N_1332);
xnor U1422 (N_1422,N_1344,N_1336);
xnor U1423 (N_1423,N_1284,N_1308);
nor U1424 (N_1424,N_1275,N_1277);
or U1425 (N_1425,N_1405,N_1372);
nand U1426 (N_1426,N_1416,N_1421);
and U1427 (N_1427,N_1409,N_1384);
or U1428 (N_1428,N_1406,N_1375);
nor U1429 (N_1429,N_1412,N_1380);
and U1430 (N_1430,N_1420,N_1368);
nor U1431 (N_1431,N_1408,N_1402);
nand U1432 (N_1432,N_1369,N_1355);
nand U1433 (N_1433,N_1371,N_1387);
and U1434 (N_1434,N_1417,N_1389);
and U1435 (N_1435,N_1395,N_1366);
or U1436 (N_1436,N_1400,N_1398);
and U1437 (N_1437,N_1363,N_1364);
and U1438 (N_1438,N_1423,N_1357);
or U1439 (N_1439,N_1388,N_1391);
nor U1440 (N_1440,N_1381,N_1397);
nand U1441 (N_1441,N_1382,N_1404);
or U1442 (N_1442,N_1386,N_1359);
or U1443 (N_1443,N_1358,N_1376);
or U1444 (N_1444,N_1351,N_1352);
nor U1445 (N_1445,N_1403,N_1396);
nor U1446 (N_1446,N_1399,N_1393);
nand U1447 (N_1447,N_1361,N_1401);
nor U1448 (N_1448,N_1362,N_1353);
and U1449 (N_1449,N_1365,N_1374);
nor U1450 (N_1450,N_1415,N_1378);
and U1451 (N_1451,N_1422,N_1419);
nand U1452 (N_1452,N_1385,N_1373);
or U1453 (N_1453,N_1418,N_1392);
nand U1454 (N_1454,N_1354,N_1410);
nand U1455 (N_1455,N_1424,N_1367);
or U1456 (N_1456,N_1411,N_1350);
or U1457 (N_1457,N_1356,N_1407);
nor U1458 (N_1458,N_1360,N_1379);
nand U1459 (N_1459,N_1370,N_1383);
nand U1460 (N_1460,N_1394,N_1390);
nor U1461 (N_1461,N_1377,N_1413);
nand U1462 (N_1462,N_1414,N_1354);
nor U1463 (N_1463,N_1376,N_1405);
nor U1464 (N_1464,N_1410,N_1405);
or U1465 (N_1465,N_1350,N_1404);
or U1466 (N_1466,N_1406,N_1379);
and U1467 (N_1467,N_1385,N_1366);
and U1468 (N_1468,N_1424,N_1393);
and U1469 (N_1469,N_1388,N_1368);
nor U1470 (N_1470,N_1417,N_1358);
nor U1471 (N_1471,N_1384,N_1392);
nand U1472 (N_1472,N_1418,N_1382);
nor U1473 (N_1473,N_1365,N_1421);
nand U1474 (N_1474,N_1350,N_1351);
xor U1475 (N_1475,N_1402,N_1400);
or U1476 (N_1476,N_1366,N_1369);
nand U1477 (N_1477,N_1402,N_1396);
and U1478 (N_1478,N_1374,N_1355);
or U1479 (N_1479,N_1414,N_1406);
xor U1480 (N_1480,N_1392,N_1421);
or U1481 (N_1481,N_1394,N_1410);
nand U1482 (N_1482,N_1423,N_1365);
nand U1483 (N_1483,N_1379,N_1359);
nand U1484 (N_1484,N_1412,N_1378);
nor U1485 (N_1485,N_1377,N_1382);
or U1486 (N_1486,N_1376,N_1401);
nor U1487 (N_1487,N_1384,N_1414);
nor U1488 (N_1488,N_1363,N_1416);
nand U1489 (N_1489,N_1422,N_1408);
nand U1490 (N_1490,N_1355,N_1360);
nor U1491 (N_1491,N_1404,N_1377);
or U1492 (N_1492,N_1385,N_1417);
nor U1493 (N_1493,N_1376,N_1360);
or U1494 (N_1494,N_1385,N_1367);
and U1495 (N_1495,N_1414,N_1362);
nor U1496 (N_1496,N_1384,N_1406);
nand U1497 (N_1497,N_1356,N_1365);
or U1498 (N_1498,N_1417,N_1393);
nand U1499 (N_1499,N_1362,N_1384);
nand U1500 (N_1500,N_1427,N_1449);
nor U1501 (N_1501,N_1465,N_1429);
nor U1502 (N_1502,N_1468,N_1474);
and U1503 (N_1503,N_1483,N_1448);
nor U1504 (N_1504,N_1477,N_1456);
and U1505 (N_1505,N_1473,N_1489);
or U1506 (N_1506,N_1475,N_1433);
or U1507 (N_1507,N_1485,N_1461);
or U1508 (N_1508,N_1454,N_1493);
or U1509 (N_1509,N_1442,N_1492);
nand U1510 (N_1510,N_1484,N_1452);
nor U1511 (N_1511,N_1497,N_1457);
or U1512 (N_1512,N_1495,N_1435);
nor U1513 (N_1513,N_1460,N_1488);
or U1514 (N_1514,N_1446,N_1428);
nand U1515 (N_1515,N_1471,N_1455);
and U1516 (N_1516,N_1466,N_1496);
and U1517 (N_1517,N_1478,N_1470);
and U1518 (N_1518,N_1440,N_1469);
nand U1519 (N_1519,N_1445,N_1444);
or U1520 (N_1520,N_1482,N_1476);
or U1521 (N_1521,N_1491,N_1436);
nand U1522 (N_1522,N_1479,N_1451);
nand U1523 (N_1523,N_1459,N_1481);
and U1524 (N_1524,N_1458,N_1438);
or U1525 (N_1525,N_1490,N_1462);
nor U1526 (N_1526,N_1498,N_1431);
and U1527 (N_1527,N_1426,N_1463);
or U1528 (N_1528,N_1425,N_1480);
and U1529 (N_1529,N_1487,N_1472);
or U1530 (N_1530,N_1447,N_1441);
and U1531 (N_1531,N_1437,N_1439);
nand U1532 (N_1532,N_1453,N_1467);
or U1533 (N_1533,N_1450,N_1494);
and U1534 (N_1534,N_1432,N_1486);
and U1535 (N_1535,N_1430,N_1443);
and U1536 (N_1536,N_1434,N_1499);
or U1537 (N_1537,N_1464,N_1454);
and U1538 (N_1538,N_1489,N_1445);
nor U1539 (N_1539,N_1426,N_1449);
or U1540 (N_1540,N_1468,N_1447);
nand U1541 (N_1541,N_1461,N_1435);
nand U1542 (N_1542,N_1470,N_1459);
or U1543 (N_1543,N_1468,N_1431);
nand U1544 (N_1544,N_1441,N_1439);
or U1545 (N_1545,N_1430,N_1437);
or U1546 (N_1546,N_1425,N_1439);
or U1547 (N_1547,N_1452,N_1434);
nand U1548 (N_1548,N_1461,N_1463);
or U1549 (N_1549,N_1495,N_1449);
nor U1550 (N_1550,N_1435,N_1491);
nand U1551 (N_1551,N_1477,N_1485);
and U1552 (N_1552,N_1456,N_1457);
or U1553 (N_1553,N_1494,N_1451);
nor U1554 (N_1554,N_1482,N_1437);
xnor U1555 (N_1555,N_1436,N_1454);
or U1556 (N_1556,N_1467,N_1441);
nand U1557 (N_1557,N_1469,N_1494);
or U1558 (N_1558,N_1492,N_1485);
nor U1559 (N_1559,N_1432,N_1455);
or U1560 (N_1560,N_1480,N_1436);
nand U1561 (N_1561,N_1445,N_1432);
or U1562 (N_1562,N_1431,N_1457);
and U1563 (N_1563,N_1432,N_1435);
or U1564 (N_1564,N_1494,N_1490);
nor U1565 (N_1565,N_1489,N_1434);
and U1566 (N_1566,N_1448,N_1439);
nor U1567 (N_1567,N_1488,N_1448);
and U1568 (N_1568,N_1488,N_1444);
and U1569 (N_1569,N_1461,N_1464);
and U1570 (N_1570,N_1449,N_1439);
nand U1571 (N_1571,N_1486,N_1458);
nand U1572 (N_1572,N_1490,N_1471);
or U1573 (N_1573,N_1489,N_1479);
and U1574 (N_1574,N_1486,N_1468);
or U1575 (N_1575,N_1506,N_1565);
and U1576 (N_1576,N_1522,N_1549);
or U1577 (N_1577,N_1515,N_1550);
nand U1578 (N_1578,N_1514,N_1542);
and U1579 (N_1579,N_1523,N_1509);
or U1580 (N_1580,N_1546,N_1548);
and U1581 (N_1581,N_1518,N_1529);
or U1582 (N_1582,N_1502,N_1524);
nand U1583 (N_1583,N_1566,N_1525);
nand U1584 (N_1584,N_1530,N_1526);
or U1585 (N_1585,N_1562,N_1553);
or U1586 (N_1586,N_1554,N_1528);
nor U1587 (N_1587,N_1574,N_1521);
and U1588 (N_1588,N_1500,N_1520);
nand U1589 (N_1589,N_1517,N_1507);
nor U1590 (N_1590,N_1551,N_1552);
nor U1591 (N_1591,N_1559,N_1563);
or U1592 (N_1592,N_1508,N_1539);
and U1593 (N_1593,N_1569,N_1560);
nand U1594 (N_1594,N_1501,N_1547);
and U1595 (N_1595,N_1503,N_1556);
nor U1596 (N_1596,N_1564,N_1544);
and U1597 (N_1597,N_1504,N_1532);
and U1598 (N_1598,N_1505,N_1531);
nor U1599 (N_1599,N_1511,N_1541);
nand U1600 (N_1600,N_1527,N_1510);
nand U1601 (N_1601,N_1558,N_1535);
nand U1602 (N_1602,N_1573,N_1545);
and U1603 (N_1603,N_1534,N_1533);
nand U1604 (N_1604,N_1571,N_1570);
and U1605 (N_1605,N_1536,N_1512);
nor U1606 (N_1606,N_1543,N_1516);
nand U1607 (N_1607,N_1567,N_1555);
nand U1608 (N_1608,N_1572,N_1537);
nand U1609 (N_1609,N_1519,N_1557);
and U1610 (N_1610,N_1568,N_1538);
and U1611 (N_1611,N_1513,N_1540);
or U1612 (N_1612,N_1561,N_1562);
or U1613 (N_1613,N_1511,N_1551);
and U1614 (N_1614,N_1515,N_1528);
nor U1615 (N_1615,N_1514,N_1549);
nand U1616 (N_1616,N_1504,N_1531);
nand U1617 (N_1617,N_1556,N_1531);
or U1618 (N_1618,N_1567,N_1558);
or U1619 (N_1619,N_1513,N_1536);
and U1620 (N_1620,N_1528,N_1502);
nand U1621 (N_1621,N_1522,N_1541);
nor U1622 (N_1622,N_1563,N_1552);
or U1623 (N_1623,N_1518,N_1523);
or U1624 (N_1624,N_1512,N_1545);
nor U1625 (N_1625,N_1507,N_1560);
nand U1626 (N_1626,N_1554,N_1563);
nor U1627 (N_1627,N_1566,N_1533);
or U1628 (N_1628,N_1555,N_1568);
or U1629 (N_1629,N_1528,N_1570);
or U1630 (N_1630,N_1509,N_1541);
or U1631 (N_1631,N_1556,N_1560);
or U1632 (N_1632,N_1573,N_1502);
nand U1633 (N_1633,N_1529,N_1515);
nor U1634 (N_1634,N_1543,N_1552);
nand U1635 (N_1635,N_1528,N_1501);
nor U1636 (N_1636,N_1512,N_1528);
or U1637 (N_1637,N_1535,N_1505);
and U1638 (N_1638,N_1513,N_1529);
and U1639 (N_1639,N_1529,N_1538);
xnor U1640 (N_1640,N_1513,N_1517);
nand U1641 (N_1641,N_1570,N_1556);
nor U1642 (N_1642,N_1551,N_1535);
or U1643 (N_1643,N_1544,N_1571);
xnor U1644 (N_1644,N_1520,N_1564);
nor U1645 (N_1645,N_1540,N_1510);
and U1646 (N_1646,N_1501,N_1527);
nand U1647 (N_1647,N_1550,N_1562);
and U1648 (N_1648,N_1549,N_1535);
or U1649 (N_1649,N_1541,N_1538);
nand U1650 (N_1650,N_1600,N_1635);
and U1651 (N_1651,N_1629,N_1632);
nor U1652 (N_1652,N_1617,N_1586);
xnor U1653 (N_1653,N_1601,N_1603);
and U1654 (N_1654,N_1644,N_1577);
and U1655 (N_1655,N_1636,N_1597);
xnor U1656 (N_1656,N_1590,N_1640);
nor U1657 (N_1657,N_1631,N_1613);
nand U1658 (N_1658,N_1641,N_1607);
and U1659 (N_1659,N_1579,N_1618);
nor U1660 (N_1660,N_1634,N_1625);
or U1661 (N_1661,N_1612,N_1642);
xor U1662 (N_1662,N_1621,N_1646);
nor U1663 (N_1663,N_1589,N_1599);
or U1664 (N_1664,N_1649,N_1645);
nand U1665 (N_1665,N_1630,N_1604);
and U1666 (N_1666,N_1575,N_1588);
or U1667 (N_1667,N_1598,N_1585);
or U1668 (N_1668,N_1615,N_1614);
or U1669 (N_1669,N_1591,N_1622);
and U1670 (N_1670,N_1624,N_1578);
nor U1671 (N_1671,N_1609,N_1594);
or U1672 (N_1672,N_1611,N_1633);
or U1673 (N_1673,N_1639,N_1580);
and U1674 (N_1674,N_1623,N_1648);
or U1675 (N_1675,N_1616,N_1647);
nand U1676 (N_1676,N_1606,N_1602);
xnor U1677 (N_1677,N_1605,N_1627);
nand U1678 (N_1678,N_1593,N_1576);
nor U1679 (N_1679,N_1626,N_1587);
and U1680 (N_1680,N_1620,N_1643);
and U1681 (N_1681,N_1584,N_1592);
nor U1682 (N_1682,N_1637,N_1628);
nand U1683 (N_1683,N_1608,N_1596);
and U1684 (N_1684,N_1582,N_1581);
or U1685 (N_1685,N_1619,N_1638);
nand U1686 (N_1686,N_1595,N_1583);
nand U1687 (N_1687,N_1610,N_1587);
xnor U1688 (N_1688,N_1592,N_1599);
nand U1689 (N_1689,N_1640,N_1595);
nor U1690 (N_1690,N_1631,N_1625);
and U1691 (N_1691,N_1602,N_1607);
nand U1692 (N_1692,N_1622,N_1643);
and U1693 (N_1693,N_1634,N_1640);
and U1694 (N_1694,N_1576,N_1641);
nor U1695 (N_1695,N_1582,N_1598);
and U1696 (N_1696,N_1584,N_1606);
nor U1697 (N_1697,N_1581,N_1593);
and U1698 (N_1698,N_1643,N_1641);
or U1699 (N_1699,N_1581,N_1599);
or U1700 (N_1700,N_1611,N_1602);
and U1701 (N_1701,N_1632,N_1596);
nand U1702 (N_1702,N_1624,N_1597);
and U1703 (N_1703,N_1582,N_1583);
or U1704 (N_1704,N_1602,N_1649);
nor U1705 (N_1705,N_1607,N_1587);
or U1706 (N_1706,N_1592,N_1643);
nor U1707 (N_1707,N_1604,N_1603);
nand U1708 (N_1708,N_1624,N_1618);
or U1709 (N_1709,N_1607,N_1648);
nand U1710 (N_1710,N_1593,N_1595);
and U1711 (N_1711,N_1594,N_1629);
or U1712 (N_1712,N_1605,N_1622);
and U1713 (N_1713,N_1627,N_1598);
and U1714 (N_1714,N_1630,N_1647);
and U1715 (N_1715,N_1625,N_1605);
and U1716 (N_1716,N_1642,N_1647);
nand U1717 (N_1717,N_1590,N_1596);
nor U1718 (N_1718,N_1634,N_1627);
nor U1719 (N_1719,N_1581,N_1590);
and U1720 (N_1720,N_1576,N_1606);
nand U1721 (N_1721,N_1618,N_1639);
nor U1722 (N_1722,N_1629,N_1624);
nand U1723 (N_1723,N_1615,N_1606);
and U1724 (N_1724,N_1627,N_1600);
or U1725 (N_1725,N_1686,N_1714);
nor U1726 (N_1726,N_1695,N_1697);
nor U1727 (N_1727,N_1709,N_1654);
nand U1728 (N_1728,N_1724,N_1719);
and U1729 (N_1729,N_1694,N_1658);
and U1730 (N_1730,N_1673,N_1653);
or U1731 (N_1731,N_1705,N_1722);
or U1732 (N_1732,N_1696,N_1721);
or U1733 (N_1733,N_1688,N_1690);
and U1734 (N_1734,N_1704,N_1665);
nor U1735 (N_1735,N_1651,N_1703);
and U1736 (N_1736,N_1713,N_1723);
nor U1737 (N_1737,N_1683,N_1700);
nor U1738 (N_1738,N_1667,N_1664);
or U1739 (N_1739,N_1720,N_1715);
nor U1740 (N_1740,N_1659,N_1672);
or U1741 (N_1741,N_1701,N_1682);
and U1742 (N_1742,N_1678,N_1660);
or U1743 (N_1743,N_1707,N_1662);
or U1744 (N_1744,N_1708,N_1677);
or U1745 (N_1745,N_1687,N_1670);
nand U1746 (N_1746,N_1684,N_1716);
nand U1747 (N_1747,N_1666,N_1702);
nand U1748 (N_1748,N_1698,N_1655);
or U1749 (N_1749,N_1706,N_1661);
and U1750 (N_1750,N_1685,N_1711);
and U1751 (N_1751,N_1675,N_1712);
nand U1752 (N_1752,N_1663,N_1689);
nor U1753 (N_1753,N_1717,N_1650);
and U1754 (N_1754,N_1671,N_1693);
nand U1755 (N_1755,N_1718,N_1692);
nand U1756 (N_1756,N_1669,N_1676);
and U1757 (N_1757,N_1657,N_1710);
nand U1758 (N_1758,N_1691,N_1680);
nand U1759 (N_1759,N_1668,N_1652);
nand U1760 (N_1760,N_1679,N_1681);
nor U1761 (N_1761,N_1656,N_1699);
nor U1762 (N_1762,N_1674,N_1679);
and U1763 (N_1763,N_1686,N_1653);
and U1764 (N_1764,N_1676,N_1693);
xnor U1765 (N_1765,N_1655,N_1672);
and U1766 (N_1766,N_1671,N_1706);
nor U1767 (N_1767,N_1668,N_1679);
nand U1768 (N_1768,N_1660,N_1652);
nor U1769 (N_1769,N_1680,N_1650);
or U1770 (N_1770,N_1719,N_1702);
and U1771 (N_1771,N_1685,N_1705);
and U1772 (N_1772,N_1663,N_1713);
nor U1773 (N_1773,N_1650,N_1665);
nor U1774 (N_1774,N_1654,N_1693);
nand U1775 (N_1775,N_1669,N_1709);
or U1776 (N_1776,N_1671,N_1707);
nand U1777 (N_1777,N_1681,N_1692);
or U1778 (N_1778,N_1656,N_1696);
or U1779 (N_1779,N_1688,N_1718);
nand U1780 (N_1780,N_1720,N_1653);
or U1781 (N_1781,N_1708,N_1695);
or U1782 (N_1782,N_1720,N_1688);
or U1783 (N_1783,N_1673,N_1703);
nand U1784 (N_1784,N_1719,N_1651);
or U1785 (N_1785,N_1673,N_1710);
nand U1786 (N_1786,N_1697,N_1673);
nand U1787 (N_1787,N_1658,N_1650);
and U1788 (N_1788,N_1709,N_1706);
or U1789 (N_1789,N_1666,N_1665);
xor U1790 (N_1790,N_1685,N_1699);
and U1791 (N_1791,N_1672,N_1670);
nand U1792 (N_1792,N_1690,N_1665);
nand U1793 (N_1793,N_1705,N_1665);
or U1794 (N_1794,N_1694,N_1683);
nor U1795 (N_1795,N_1654,N_1676);
or U1796 (N_1796,N_1654,N_1708);
nor U1797 (N_1797,N_1696,N_1670);
and U1798 (N_1798,N_1698,N_1711);
nand U1799 (N_1799,N_1713,N_1686);
and U1800 (N_1800,N_1727,N_1749);
or U1801 (N_1801,N_1735,N_1754);
or U1802 (N_1802,N_1742,N_1733);
or U1803 (N_1803,N_1729,N_1795);
xnor U1804 (N_1804,N_1756,N_1796);
and U1805 (N_1805,N_1753,N_1755);
and U1806 (N_1806,N_1761,N_1747);
or U1807 (N_1807,N_1748,N_1788);
nand U1808 (N_1808,N_1789,N_1781);
and U1809 (N_1809,N_1798,N_1752);
or U1810 (N_1810,N_1776,N_1732);
xnor U1811 (N_1811,N_1777,N_1785);
nor U1812 (N_1812,N_1772,N_1799);
and U1813 (N_1813,N_1780,N_1737);
nor U1814 (N_1814,N_1797,N_1773);
nor U1815 (N_1815,N_1771,N_1758);
and U1816 (N_1816,N_1770,N_1757);
nand U1817 (N_1817,N_1782,N_1736);
nand U1818 (N_1818,N_1763,N_1746);
nand U1819 (N_1819,N_1786,N_1784);
or U1820 (N_1820,N_1741,N_1750);
nor U1821 (N_1821,N_1759,N_1765);
nor U1822 (N_1822,N_1791,N_1787);
nor U1823 (N_1823,N_1775,N_1731);
nand U1824 (N_1824,N_1734,N_1783);
and U1825 (N_1825,N_1762,N_1728);
nand U1826 (N_1826,N_1743,N_1778);
or U1827 (N_1827,N_1792,N_1768);
nand U1828 (N_1828,N_1739,N_1738);
or U1829 (N_1829,N_1774,N_1779);
nor U1830 (N_1830,N_1769,N_1726);
and U1831 (N_1831,N_1744,N_1766);
and U1832 (N_1832,N_1740,N_1764);
nor U1833 (N_1833,N_1745,N_1790);
and U1834 (N_1834,N_1793,N_1760);
nand U1835 (N_1835,N_1725,N_1794);
nor U1836 (N_1836,N_1751,N_1767);
nor U1837 (N_1837,N_1730,N_1761);
nand U1838 (N_1838,N_1734,N_1793);
or U1839 (N_1839,N_1781,N_1791);
and U1840 (N_1840,N_1727,N_1788);
or U1841 (N_1841,N_1774,N_1764);
nor U1842 (N_1842,N_1770,N_1790);
or U1843 (N_1843,N_1770,N_1798);
or U1844 (N_1844,N_1728,N_1795);
nand U1845 (N_1845,N_1733,N_1798);
nor U1846 (N_1846,N_1741,N_1759);
nor U1847 (N_1847,N_1756,N_1758);
nor U1848 (N_1848,N_1766,N_1731);
nor U1849 (N_1849,N_1758,N_1763);
nor U1850 (N_1850,N_1745,N_1799);
xor U1851 (N_1851,N_1757,N_1733);
nand U1852 (N_1852,N_1763,N_1766);
and U1853 (N_1853,N_1763,N_1765);
xor U1854 (N_1854,N_1794,N_1791);
nor U1855 (N_1855,N_1780,N_1783);
or U1856 (N_1856,N_1740,N_1757);
nand U1857 (N_1857,N_1778,N_1738);
nor U1858 (N_1858,N_1789,N_1788);
xor U1859 (N_1859,N_1777,N_1743);
or U1860 (N_1860,N_1749,N_1761);
or U1861 (N_1861,N_1726,N_1743);
and U1862 (N_1862,N_1746,N_1789);
or U1863 (N_1863,N_1779,N_1738);
and U1864 (N_1864,N_1736,N_1794);
or U1865 (N_1865,N_1793,N_1785);
or U1866 (N_1866,N_1762,N_1771);
nor U1867 (N_1867,N_1798,N_1795);
nor U1868 (N_1868,N_1797,N_1769);
nor U1869 (N_1869,N_1789,N_1770);
and U1870 (N_1870,N_1765,N_1757);
nor U1871 (N_1871,N_1783,N_1760);
and U1872 (N_1872,N_1771,N_1752);
and U1873 (N_1873,N_1734,N_1796);
or U1874 (N_1874,N_1729,N_1790);
or U1875 (N_1875,N_1848,N_1806);
nor U1876 (N_1876,N_1841,N_1861);
and U1877 (N_1877,N_1858,N_1833);
nor U1878 (N_1878,N_1809,N_1868);
nand U1879 (N_1879,N_1855,N_1817);
xnor U1880 (N_1880,N_1807,N_1854);
nand U1881 (N_1881,N_1835,N_1872);
nand U1882 (N_1882,N_1822,N_1862);
or U1883 (N_1883,N_1805,N_1818);
or U1884 (N_1884,N_1812,N_1873);
and U1885 (N_1885,N_1857,N_1840);
nand U1886 (N_1886,N_1859,N_1815);
nor U1887 (N_1887,N_1813,N_1850);
and U1888 (N_1888,N_1871,N_1830);
or U1889 (N_1889,N_1816,N_1804);
nor U1890 (N_1890,N_1838,N_1846);
or U1891 (N_1891,N_1856,N_1810);
nor U1892 (N_1892,N_1820,N_1826);
and U1893 (N_1893,N_1803,N_1831);
nand U1894 (N_1894,N_1863,N_1845);
nor U1895 (N_1895,N_1834,N_1853);
or U1896 (N_1896,N_1874,N_1801);
nor U1897 (N_1897,N_1832,N_1842);
or U1898 (N_1898,N_1802,N_1870);
and U1899 (N_1899,N_1800,N_1839);
nand U1900 (N_1900,N_1836,N_1869);
and U1901 (N_1901,N_1865,N_1866);
or U1902 (N_1902,N_1837,N_1823);
nor U1903 (N_1903,N_1814,N_1829);
nor U1904 (N_1904,N_1827,N_1852);
nand U1905 (N_1905,N_1851,N_1808);
nand U1906 (N_1906,N_1819,N_1864);
nand U1907 (N_1907,N_1821,N_1811);
or U1908 (N_1908,N_1825,N_1849);
xnor U1909 (N_1909,N_1860,N_1847);
nor U1910 (N_1910,N_1824,N_1828);
and U1911 (N_1911,N_1843,N_1867);
nor U1912 (N_1912,N_1844,N_1857);
nor U1913 (N_1913,N_1836,N_1870);
and U1914 (N_1914,N_1874,N_1852);
nor U1915 (N_1915,N_1849,N_1837);
nand U1916 (N_1916,N_1826,N_1872);
nand U1917 (N_1917,N_1853,N_1828);
or U1918 (N_1918,N_1871,N_1845);
and U1919 (N_1919,N_1849,N_1803);
or U1920 (N_1920,N_1867,N_1873);
or U1921 (N_1921,N_1837,N_1817);
and U1922 (N_1922,N_1839,N_1829);
and U1923 (N_1923,N_1839,N_1840);
and U1924 (N_1924,N_1830,N_1849);
nor U1925 (N_1925,N_1815,N_1801);
and U1926 (N_1926,N_1814,N_1839);
and U1927 (N_1927,N_1811,N_1858);
or U1928 (N_1928,N_1811,N_1836);
nand U1929 (N_1929,N_1851,N_1806);
nor U1930 (N_1930,N_1812,N_1839);
or U1931 (N_1931,N_1831,N_1858);
nor U1932 (N_1932,N_1824,N_1802);
or U1933 (N_1933,N_1841,N_1820);
nand U1934 (N_1934,N_1856,N_1840);
or U1935 (N_1935,N_1840,N_1806);
or U1936 (N_1936,N_1805,N_1804);
nand U1937 (N_1937,N_1805,N_1837);
and U1938 (N_1938,N_1843,N_1868);
and U1939 (N_1939,N_1802,N_1862);
nand U1940 (N_1940,N_1808,N_1840);
nor U1941 (N_1941,N_1828,N_1873);
or U1942 (N_1942,N_1871,N_1859);
and U1943 (N_1943,N_1811,N_1806);
or U1944 (N_1944,N_1819,N_1854);
and U1945 (N_1945,N_1818,N_1815);
nor U1946 (N_1946,N_1838,N_1844);
or U1947 (N_1947,N_1859,N_1808);
nand U1948 (N_1948,N_1829,N_1871);
and U1949 (N_1949,N_1869,N_1843);
nor U1950 (N_1950,N_1946,N_1922);
nand U1951 (N_1951,N_1880,N_1934);
nor U1952 (N_1952,N_1916,N_1935);
nand U1953 (N_1953,N_1891,N_1903);
nand U1954 (N_1954,N_1905,N_1948);
and U1955 (N_1955,N_1894,N_1907);
or U1956 (N_1956,N_1924,N_1913);
nand U1957 (N_1957,N_1926,N_1941);
or U1958 (N_1958,N_1931,N_1896);
and U1959 (N_1959,N_1887,N_1892);
or U1960 (N_1960,N_1875,N_1925);
nor U1961 (N_1961,N_1885,N_1940);
nor U1962 (N_1962,N_1898,N_1921);
or U1963 (N_1963,N_1930,N_1888);
xor U1964 (N_1964,N_1889,N_1904);
nor U1965 (N_1965,N_1879,N_1895);
nand U1966 (N_1966,N_1876,N_1897);
xor U1967 (N_1967,N_1902,N_1901);
nand U1968 (N_1968,N_1927,N_1890);
and U1969 (N_1969,N_1900,N_1899);
nand U1970 (N_1970,N_1915,N_1929);
nand U1971 (N_1971,N_1877,N_1947);
nand U1972 (N_1972,N_1932,N_1928);
nor U1973 (N_1973,N_1937,N_1943);
nand U1974 (N_1974,N_1942,N_1919);
nand U1975 (N_1975,N_1911,N_1906);
or U1976 (N_1976,N_1936,N_1912);
nand U1977 (N_1977,N_1884,N_1886);
or U1978 (N_1978,N_1918,N_1881);
or U1979 (N_1979,N_1933,N_1945);
and U1980 (N_1980,N_1923,N_1882);
and U1981 (N_1981,N_1920,N_1908);
and U1982 (N_1982,N_1878,N_1917);
nand U1983 (N_1983,N_1949,N_1939);
nor U1984 (N_1984,N_1944,N_1914);
nor U1985 (N_1985,N_1938,N_1893);
or U1986 (N_1986,N_1883,N_1909);
and U1987 (N_1987,N_1910,N_1931);
or U1988 (N_1988,N_1934,N_1946);
nand U1989 (N_1989,N_1940,N_1878);
and U1990 (N_1990,N_1904,N_1897);
and U1991 (N_1991,N_1888,N_1926);
nand U1992 (N_1992,N_1880,N_1913);
nand U1993 (N_1993,N_1876,N_1908);
nand U1994 (N_1994,N_1915,N_1940);
or U1995 (N_1995,N_1882,N_1922);
and U1996 (N_1996,N_1933,N_1907);
and U1997 (N_1997,N_1897,N_1925);
nand U1998 (N_1998,N_1906,N_1879);
and U1999 (N_1999,N_1926,N_1880);
nand U2000 (N_2000,N_1919,N_1898);
and U2001 (N_2001,N_1907,N_1945);
and U2002 (N_2002,N_1886,N_1948);
or U2003 (N_2003,N_1936,N_1942);
and U2004 (N_2004,N_1903,N_1901);
or U2005 (N_2005,N_1915,N_1896);
and U2006 (N_2006,N_1911,N_1909);
xor U2007 (N_2007,N_1903,N_1907);
nor U2008 (N_2008,N_1889,N_1881);
or U2009 (N_2009,N_1923,N_1879);
or U2010 (N_2010,N_1899,N_1934);
nand U2011 (N_2011,N_1908,N_1925);
nand U2012 (N_2012,N_1939,N_1885);
or U2013 (N_2013,N_1891,N_1937);
and U2014 (N_2014,N_1918,N_1893);
nand U2015 (N_2015,N_1943,N_1898);
and U2016 (N_2016,N_1877,N_1921);
or U2017 (N_2017,N_1885,N_1924);
nor U2018 (N_2018,N_1878,N_1938);
nand U2019 (N_2019,N_1917,N_1898);
and U2020 (N_2020,N_1885,N_1918);
and U2021 (N_2021,N_1909,N_1877);
nand U2022 (N_2022,N_1933,N_1886);
or U2023 (N_2023,N_1893,N_1923);
nand U2024 (N_2024,N_1942,N_1928);
nor U2025 (N_2025,N_1982,N_2014);
nand U2026 (N_2026,N_1985,N_1956);
or U2027 (N_2027,N_1984,N_1989);
or U2028 (N_2028,N_2000,N_2002);
nor U2029 (N_2029,N_1979,N_1969);
nand U2030 (N_2030,N_1992,N_1953);
nand U2031 (N_2031,N_1983,N_1958);
nand U2032 (N_2032,N_1981,N_1960);
nor U2033 (N_2033,N_1991,N_2008);
nor U2034 (N_2034,N_2017,N_1988);
nor U2035 (N_2035,N_1957,N_1993);
and U2036 (N_2036,N_1994,N_2019);
or U2037 (N_2037,N_2005,N_2004);
xor U2038 (N_2038,N_2023,N_2012);
or U2039 (N_2039,N_2020,N_1997);
nor U2040 (N_2040,N_1952,N_1954);
or U2041 (N_2041,N_1967,N_1964);
nor U2042 (N_2042,N_1968,N_1973);
and U2043 (N_2043,N_2006,N_1961);
or U2044 (N_2044,N_1972,N_1951);
and U2045 (N_2045,N_2013,N_2024);
or U2046 (N_2046,N_1996,N_2010);
or U2047 (N_2047,N_1976,N_1980);
nand U2048 (N_2048,N_1971,N_1963);
and U2049 (N_2049,N_2016,N_2009);
nand U2050 (N_2050,N_2015,N_1955);
nor U2051 (N_2051,N_1966,N_1959);
or U2052 (N_2052,N_1975,N_1950);
nor U2053 (N_2053,N_2021,N_1977);
and U2054 (N_2054,N_1995,N_2022);
and U2055 (N_2055,N_2018,N_1978);
or U2056 (N_2056,N_1974,N_1987);
nor U2057 (N_2057,N_2011,N_1990);
nor U2058 (N_2058,N_1998,N_1970);
or U2059 (N_2059,N_1962,N_1965);
or U2060 (N_2060,N_2001,N_1986);
and U2061 (N_2061,N_1999,N_2003);
or U2062 (N_2062,N_2007,N_2024);
nor U2063 (N_2063,N_2008,N_1971);
or U2064 (N_2064,N_1992,N_1971);
nor U2065 (N_2065,N_1959,N_1957);
and U2066 (N_2066,N_1996,N_1978);
nand U2067 (N_2067,N_1958,N_1969);
nand U2068 (N_2068,N_2006,N_2001);
and U2069 (N_2069,N_2022,N_2019);
or U2070 (N_2070,N_2019,N_2006);
or U2071 (N_2071,N_2023,N_1961);
nor U2072 (N_2072,N_1957,N_2008);
and U2073 (N_2073,N_1954,N_2021);
or U2074 (N_2074,N_1995,N_2012);
nor U2075 (N_2075,N_1952,N_2001);
or U2076 (N_2076,N_1986,N_1984);
xor U2077 (N_2077,N_1954,N_1988);
nor U2078 (N_2078,N_2004,N_1999);
and U2079 (N_2079,N_1972,N_2002);
nand U2080 (N_2080,N_1979,N_1956);
nor U2081 (N_2081,N_2019,N_1991);
or U2082 (N_2082,N_1980,N_1970);
or U2083 (N_2083,N_2002,N_2024);
nor U2084 (N_2084,N_1970,N_2024);
and U2085 (N_2085,N_1953,N_1993);
nand U2086 (N_2086,N_1960,N_2009);
nor U2087 (N_2087,N_2020,N_2001);
nand U2088 (N_2088,N_2020,N_2010);
nor U2089 (N_2089,N_1972,N_1980);
nor U2090 (N_2090,N_2003,N_1990);
and U2091 (N_2091,N_2000,N_2004);
nand U2092 (N_2092,N_1993,N_2014);
nor U2093 (N_2093,N_2013,N_1980);
or U2094 (N_2094,N_1998,N_1990);
or U2095 (N_2095,N_1967,N_2009);
nand U2096 (N_2096,N_1986,N_1992);
and U2097 (N_2097,N_1981,N_2022);
nand U2098 (N_2098,N_1987,N_2018);
nand U2099 (N_2099,N_1987,N_1964);
or U2100 (N_2100,N_2074,N_2080);
nand U2101 (N_2101,N_2073,N_2094);
nor U2102 (N_2102,N_2026,N_2069);
and U2103 (N_2103,N_2029,N_2082);
nor U2104 (N_2104,N_2060,N_2065);
and U2105 (N_2105,N_2033,N_2031);
nand U2106 (N_2106,N_2053,N_2058);
nor U2107 (N_2107,N_2048,N_2089);
nor U2108 (N_2108,N_2057,N_2038);
or U2109 (N_2109,N_2071,N_2028);
and U2110 (N_2110,N_2095,N_2086);
or U2111 (N_2111,N_2040,N_2059);
nand U2112 (N_2112,N_2054,N_2052);
nand U2113 (N_2113,N_2092,N_2055);
nand U2114 (N_2114,N_2041,N_2072);
and U2115 (N_2115,N_2037,N_2079);
and U2116 (N_2116,N_2063,N_2068);
nand U2117 (N_2117,N_2078,N_2088);
nor U2118 (N_2118,N_2036,N_2087);
or U2119 (N_2119,N_2047,N_2066);
xor U2120 (N_2120,N_2044,N_2098);
or U2121 (N_2121,N_2090,N_2067);
and U2122 (N_2122,N_2025,N_2027);
nand U2123 (N_2123,N_2075,N_2096);
nor U2124 (N_2124,N_2085,N_2061);
and U2125 (N_2125,N_2056,N_2064);
nor U2126 (N_2126,N_2042,N_2081);
nor U2127 (N_2127,N_2030,N_2032);
nor U2128 (N_2128,N_2051,N_2091);
nor U2129 (N_2129,N_2039,N_2070);
nor U2130 (N_2130,N_2043,N_2034);
nand U2131 (N_2131,N_2077,N_2093);
nor U2132 (N_2132,N_2084,N_2045);
nand U2133 (N_2133,N_2097,N_2099);
nor U2134 (N_2134,N_2050,N_2062);
nand U2135 (N_2135,N_2083,N_2035);
or U2136 (N_2136,N_2046,N_2049);
nand U2137 (N_2137,N_2076,N_2030);
nand U2138 (N_2138,N_2028,N_2070);
and U2139 (N_2139,N_2051,N_2085);
nor U2140 (N_2140,N_2032,N_2044);
or U2141 (N_2141,N_2069,N_2061);
nor U2142 (N_2142,N_2090,N_2031);
or U2143 (N_2143,N_2096,N_2054);
or U2144 (N_2144,N_2048,N_2090);
and U2145 (N_2145,N_2053,N_2086);
nand U2146 (N_2146,N_2069,N_2031);
or U2147 (N_2147,N_2035,N_2095);
and U2148 (N_2148,N_2066,N_2095);
nand U2149 (N_2149,N_2091,N_2093);
nor U2150 (N_2150,N_2081,N_2026);
nor U2151 (N_2151,N_2081,N_2034);
nor U2152 (N_2152,N_2062,N_2066);
or U2153 (N_2153,N_2026,N_2034);
nor U2154 (N_2154,N_2099,N_2036);
nand U2155 (N_2155,N_2096,N_2031);
or U2156 (N_2156,N_2064,N_2089);
or U2157 (N_2157,N_2083,N_2064);
nor U2158 (N_2158,N_2080,N_2061);
or U2159 (N_2159,N_2089,N_2076);
nand U2160 (N_2160,N_2053,N_2085);
xnor U2161 (N_2161,N_2030,N_2082);
nand U2162 (N_2162,N_2025,N_2056);
and U2163 (N_2163,N_2067,N_2030);
nand U2164 (N_2164,N_2039,N_2083);
nor U2165 (N_2165,N_2075,N_2031);
and U2166 (N_2166,N_2089,N_2028);
nand U2167 (N_2167,N_2035,N_2034);
nor U2168 (N_2168,N_2056,N_2039);
nor U2169 (N_2169,N_2088,N_2044);
and U2170 (N_2170,N_2095,N_2057);
nand U2171 (N_2171,N_2063,N_2073);
or U2172 (N_2172,N_2068,N_2076);
and U2173 (N_2173,N_2095,N_2098);
nand U2174 (N_2174,N_2050,N_2083);
nor U2175 (N_2175,N_2145,N_2119);
xor U2176 (N_2176,N_2171,N_2129);
nor U2177 (N_2177,N_2139,N_2121);
or U2178 (N_2178,N_2144,N_2109);
or U2179 (N_2179,N_2136,N_2150);
or U2180 (N_2180,N_2137,N_2114);
or U2181 (N_2181,N_2141,N_2142);
and U2182 (N_2182,N_2118,N_2152);
or U2183 (N_2183,N_2103,N_2130);
nor U2184 (N_2184,N_2167,N_2124);
nand U2185 (N_2185,N_2111,N_2158);
and U2186 (N_2186,N_2115,N_2163);
nor U2187 (N_2187,N_2107,N_2156);
or U2188 (N_2188,N_2108,N_2113);
nor U2189 (N_2189,N_2164,N_2153);
and U2190 (N_2190,N_2173,N_2117);
nor U2191 (N_2191,N_2161,N_2165);
nor U2192 (N_2192,N_2143,N_2146);
or U2193 (N_2193,N_2116,N_2169);
or U2194 (N_2194,N_2133,N_2159);
nor U2195 (N_2195,N_2101,N_2148);
or U2196 (N_2196,N_2100,N_2168);
nor U2197 (N_2197,N_2102,N_2127);
nor U2198 (N_2198,N_2128,N_2157);
or U2199 (N_2199,N_2162,N_2126);
or U2200 (N_2200,N_2106,N_2140);
or U2201 (N_2201,N_2132,N_2120);
and U2202 (N_2202,N_2104,N_2122);
nor U2203 (N_2203,N_2170,N_2134);
nand U2204 (N_2204,N_2112,N_2147);
nand U2205 (N_2205,N_2125,N_2160);
and U2206 (N_2206,N_2174,N_2135);
nand U2207 (N_2207,N_2172,N_2149);
xor U2208 (N_2208,N_2131,N_2110);
nand U2209 (N_2209,N_2138,N_2123);
nor U2210 (N_2210,N_2105,N_2155);
and U2211 (N_2211,N_2166,N_2154);
nor U2212 (N_2212,N_2151,N_2106);
nor U2213 (N_2213,N_2158,N_2109);
xnor U2214 (N_2214,N_2165,N_2139);
or U2215 (N_2215,N_2129,N_2161);
or U2216 (N_2216,N_2111,N_2151);
and U2217 (N_2217,N_2106,N_2164);
nor U2218 (N_2218,N_2126,N_2110);
nor U2219 (N_2219,N_2172,N_2102);
nor U2220 (N_2220,N_2156,N_2149);
or U2221 (N_2221,N_2107,N_2154);
nand U2222 (N_2222,N_2152,N_2171);
nand U2223 (N_2223,N_2157,N_2144);
or U2224 (N_2224,N_2166,N_2132);
nor U2225 (N_2225,N_2133,N_2170);
or U2226 (N_2226,N_2124,N_2136);
nand U2227 (N_2227,N_2106,N_2155);
or U2228 (N_2228,N_2125,N_2161);
and U2229 (N_2229,N_2150,N_2145);
or U2230 (N_2230,N_2112,N_2149);
nor U2231 (N_2231,N_2147,N_2146);
or U2232 (N_2232,N_2129,N_2170);
nand U2233 (N_2233,N_2108,N_2123);
xor U2234 (N_2234,N_2115,N_2156);
nor U2235 (N_2235,N_2168,N_2152);
xnor U2236 (N_2236,N_2112,N_2103);
xnor U2237 (N_2237,N_2119,N_2109);
nand U2238 (N_2238,N_2122,N_2101);
nor U2239 (N_2239,N_2100,N_2139);
and U2240 (N_2240,N_2134,N_2152);
nor U2241 (N_2241,N_2162,N_2113);
nand U2242 (N_2242,N_2144,N_2111);
nand U2243 (N_2243,N_2151,N_2121);
nand U2244 (N_2244,N_2110,N_2165);
or U2245 (N_2245,N_2117,N_2129);
nand U2246 (N_2246,N_2172,N_2167);
nand U2247 (N_2247,N_2120,N_2117);
and U2248 (N_2248,N_2167,N_2101);
nor U2249 (N_2249,N_2127,N_2136);
and U2250 (N_2250,N_2249,N_2175);
or U2251 (N_2251,N_2200,N_2183);
nand U2252 (N_2252,N_2247,N_2229);
nand U2253 (N_2253,N_2240,N_2178);
nor U2254 (N_2254,N_2243,N_2196);
or U2255 (N_2255,N_2205,N_2180);
nand U2256 (N_2256,N_2207,N_2232);
or U2257 (N_2257,N_2238,N_2176);
nand U2258 (N_2258,N_2188,N_2204);
nor U2259 (N_2259,N_2186,N_2218);
nand U2260 (N_2260,N_2181,N_2203);
nor U2261 (N_2261,N_2224,N_2236);
nor U2262 (N_2262,N_2223,N_2190);
nor U2263 (N_2263,N_2216,N_2187);
nor U2264 (N_2264,N_2198,N_2195);
or U2265 (N_2265,N_2230,N_2237);
or U2266 (N_2266,N_2209,N_2208);
nand U2267 (N_2267,N_2212,N_2213);
nor U2268 (N_2268,N_2201,N_2210);
nand U2269 (N_2269,N_2242,N_2245);
nand U2270 (N_2270,N_2220,N_2182);
nand U2271 (N_2271,N_2185,N_2239);
and U2272 (N_2272,N_2191,N_2199);
nor U2273 (N_2273,N_2221,N_2177);
and U2274 (N_2274,N_2228,N_2206);
nand U2275 (N_2275,N_2211,N_2226);
nor U2276 (N_2276,N_2179,N_2241);
nand U2277 (N_2277,N_2193,N_2215);
nor U2278 (N_2278,N_2233,N_2244);
and U2279 (N_2279,N_2217,N_2189);
and U2280 (N_2280,N_2235,N_2197);
nor U2281 (N_2281,N_2234,N_2202);
and U2282 (N_2282,N_2231,N_2219);
xor U2283 (N_2283,N_2246,N_2227);
and U2284 (N_2284,N_2225,N_2184);
nor U2285 (N_2285,N_2192,N_2194);
nor U2286 (N_2286,N_2214,N_2222);
nor U2287 (N_2287,N_2248,N_2180);
and U2288 (N_2288,N_2220,N_2200);
and U2289 (N_2289,N_2183,N_2223);
and U2290 (N_2290,N_2227,N_2226);
and U2291 (N_2291,N_2199,N_2235);
and U2292 (N_2292,N_2177,N_2244);
and U2293 (N_2293,N_2180,N_2189);
nand U2294 (N_2294,N_2249,N_2235);
or U2295 (N_2295,N_2234,N_2232);
and U2296 (N_2296,N_2203,N_2225);
and U2297 (N_2297,N_2177,N_2195);
nor U2298 (N_2298,N_2192,N_2208);
or U2299 (N_2299,N_2201,N_2207);
nor U2300 (N_2300,N_2180,N_2224);
or U2301 (N_2301,N_2190,N_2192);
and U2302 (N_2302,N_2199,N_2247);
or U2303 (N_2303,N_2234,N_2219);
and U2304 (N_2304,N_2196,N_2234);
or U2305 (N_2305,N_2204,N_2247);
nand U2306 (N_2306,N_2208,N_2205);
nor U2307 (N_2307,N_2196,N_2185);
xor U2308 (N_2308,N_2248,N_2189);
nand U2309 (N_2309,N_2221,N_2234);
nand U2310 (N_2310,N_2184,N_2223);
nand U2311 (N_2311,N_2210,N_2241);
or U2312 (N_2312,N_2198,N_2189);
nor U2313 (N_2313,N_2178,N_2232);
nor U2314 (N_2314,N_2232,N_2219);
nor U2315 (N_2315,N_2247,N_2215);
nand U2316 (N_2316,N_2239,N_2188);
and U2317 (N_2317,N_2231,N_2200);
nor U2318 (N_2318,N_2209,N_2215);
nand U2319 (N_2319,N_2231,N_2188);
nor U2320 (N_2320,N_2204,N_2234);
nand U2321 (N_2321,N_2184,N_2222);
or U2322 (N_2322,N_2216,N_2227);
and U2323 (N_2323,N_2247,N_2206);
nand U2324 (N_2324,N_2234,N_2207);
nand U2325 (N_2325,N_2279,N_2309);
and U2326 (N_2326,N_2290,N_2299);
nor U2327 (N_2327,N_2256,N_2306);
nand U2328 (N_2328,N_2261,N_2263);
or U2329 (N_2329,N_2311,N_2298);
or U2330 (N_2330,N_2313,N_2252);
nand U2331 (N_2331,N_2315,N_2269);
nor U2332 (N_2332,N_2296,N_2267);
nand U2333 (N_2333,N_2282,N_2319);
and U2334 (N_2334,N_2255,N_2322);
nand U2335 (N_2335,N_2250,N_2317);
nand U2336 (N_2336,N_2253,N_2314);
and U2337 (N_2337,N_2303,N_2257);
nand U2338 (N_2338,N_2285,N_2280);
nand U2339 (N_2339,N_2262,N_2265);
nand U2340 (N_2340,N_2324,N_2302);
or U2341 (N_2341,N_2266,N_2274);
nor U2342 (N_2342,N_2268,N_2271);
and U2343 (N_2343,N_2304,N_2312);
and U2344 (N_2344,N_2308,N_2260);
nor U2345 (N_2345,N_2251,N_2316);
or U2346 (N_2346,N_2281,N_2293);
nand U2347 (N_2347,N_2254,N_2318);
and U2348 (N_2348,N_2323,N_2264);
and U2349 (N_2349,N_2288,N_2292);
nor U2350 (N_2350,N_2321,N_2258);
or U2351 (N_2351,N_2291,N_2320);
nor U2352 (N_2352,N_2286,N_2270);
nand U2353 (N_2353,N_2289,N_2278);
nor U2354 (N_2354,N_2294,N_2276);
or U2355 (N_2355,N_2277,N_2287);
nor U2356 (N_2356,N_2300,N_2301);
nand U2357 (N_2357,N_2275,N_2283);
and U2358 (N_2358,N_2305,N_2284);
or U2359 (N_2359,N_2295,N_2297);
nand U2360 (N_2360,N_2310,N_2272);
nor U2361 (N_2361,N_2259,N_2307);
and U2362 (N_2362,N_2273,N_2251);
and U2363 (N_2363,N_2294,N_2277);
and U2364 (N_2364,N_2316,N_2253);
and U2365 (N_2365,N_2309,N_2256);
or U2366 (N_2366,N_2314,N_2275);
nor U2367 (N_2367,N_2298,N_2312);
and U2368 (N_2368,N_2291,N_2265);
and U2369 (N_2369,N_2296,N_2318);
and U2370 (N_2370,N_2283,N_2280);
and U2371 (N_2371,N_2279,N_2269);
nor U2372 (N_2372,N_2260,N_2277);
nand U2373 (N_2373,N_2281,N_2306);
or U2374 (N_2374,N_2316,N_2299);
nor U2375 (N_2375,N_2322,N_2288);
nor U2376 (N_2376,N_2324,N_2308);
and U2377 (N_2377,N_2291,N_2275);
nand U2378 (N_2378,N_2309,N_2305);
and U2379 (N_2379,N_2275,N_2259);
nor U2380 (N_2380,N_2299,N_2293);
and U2381 (N_2381,N_2270,N_2262);
or U2382 (N_2382,N_2317,N_2273);
and U2383 (N_2383,N_2300,N_2303);
and U2384 (N_2384,N_2292,N_2252);
nor U2385 (N_2385,N_2287,N_2250);
and U2386 (N_2386,N_2293,N_2258);
and U2387 (N_2387,N_2280,N_2270);
nand U2388 (N_2388,N_2322,N_2290);
or U2389 (N_2389,N_2290,N_2263);
nand U2390 (N_2390,N_2303,N_2312);
nor U2391 (N_2391,N_2308,N_2278);
nand U2392 (N_2392,N_2272,N_2289);
and U2393 (N_2393,N_2260,N_2253);
nor U2394 (N_2394,N_2287,N_2291);
or U2395 (N_2395,N_2251,N_2299);
and U2396 (N_2396,N_2275,N_2284);
or U2397 (N_2397,N_2277,N_2309);
nor U2398 (N_2398,N_2280,N_2276);
and U2399 (N_2399,N_2258,N_2270);
and U2400 (N_2400,N_2348,N_2390);
nor U2401 (N_2401,N_2353,N_2327);
nand U2402 (N_2402,N_2398,N_2362);
xor U2403 (N_2403,N_2330,N_2356);
nor U2404 (N_2404,N_2361,N_2337);
nor U2405 (N_2405,N_2378,N_2397);
nor U2406 (N_2406,N_2367,N_2387);
and U2407 (N_2407,N_2355,N_2366);
nor U2408 (N_2408,N_2358,N_2325);
nand U2409 (N_2409,N_2332,N_2385);
or U2410 (N_2410,N_2336,N_2394);
or U2411 (N_2411,N_2351,N_2359);
nand U2412 (N_2412,N_2388,N_2386);
nor U2413 (N_2413,N_2393,N_2339);
nor U2414 (N_2414,N_2368,N_2370);
or U2415 (N_2415,N_2350,N_2363);
nand U2416 (N_2416,N_2349,N_2352);
and U2417 (N_2417,N_2382,N_2375);
or U2418 (N_2418,N_2328,N_2344);
nor U2419 (N_2419,N_2395,N_2392);
nor U2420 (N_2420,N_2383,N_2360);
nand U2421 (N_2421,N_2364,N_2346);
or U2422 (N_2422,N_2389,N_2399);
nand U2423 (N_2423,N_2326,N_2357);
and U2424 (N_2424,N_2329,N_2335);
and U2425 (N_2425,N_2347,N_2333);
or U2426 (N_2426,N_2380,N_2373);
xor U2427 (N_2427,N_2343,N_2374);
and U2428 (N_2428,N_2381,N_2391);
or U2429 (N_2429,N_2345,N_2371);
nor U2430 (N_2430,N_2334,N_2377);
or U2431 (N_2431,N_2369,N_2372);
nand U2432 (N_2432,N_2354,N_2331);
or U2433 (N_2433,N_2338,N_2342);
nor U2434 (N_2434,N_2384,N_2340);
and U2435 (N_2435,N_2376,N_2396);
nand U2436 (N_2436,N_2341,N_2365);
and U2437 (N_2437,N_2379,N_2392);
or U2438 (N_2438,N_2357,N_2377);
nand U2439 (N_2439,N_2398,N_2369);
or U2440 (N_2440,N_2362,N_2349);
xnor U2441 (N_2441,N_2340,N_2389);
or U2442 (N_2442,N_2396,N_2384);
and U2443 (N_2443,N_2325,N_2326);
and U2444 (N_2444,N_2386,N_2384);
or U2445 (N_2445,N_2399,N_2391);
nor U2446 (N_2446,N_2329,N_2345);
nor U2447 (N_2447,N_2336,N_2339);
nand U2448 (N_2448,N_2333,N_2359);
or U2449 (N_2449,N_2353,N_2372);
and U2450 (N_2450,N_2375,N_2369);
or U2451 (N_2451,N_2354,N_2329);
nand U2452 (N_2452,N_2366,N_2388);
or U2453 (N_2453,N_2374,N_2376);
or U2454 (N_2454,N_2384,N_2351);
nand U2455 (N_2455,N_2347,N_2397);
nand U2456 (N_2456,N_2333,N_2395);
or U2457 (N_2457,N_2357,N_2360);
and U2458 (N_2458,N_2373,N_2328);
nand U2459 (N_2459,N_2348,N_2373);
nand U2460 (N_2460,N_2343,N_2387);
nand U2461 (N_2461,N_2377,N_2340);
nor U2462 (N_2462,N_2377,N_2347);
and U2463 (N_2463,N_2350,N_2337);
xor U2464 (N_2464,N_2336,N_2376);
and U2465 (N_2465,N_2362,N_2334);
nor U2466 (N_2466,N_2345,N_2350);
nand U2467 (N_2467,N_2392,N_2371);
nand U2468 (N_2468,N_2329,N_2347);
nor U2469 (N_2469,N_2381,N_2377);
nand U2470 (N_2470,N_2369,N_2384);
and U2471 (N_2471,N_2382,N_2369);
xnor U2472 (N_2472,N_2360,N_2356);
nor U2473 (N_2473,N_2346,N_2382);
nor U2474 (N_2474,N_2367,N_2328);
nand U2475 (N_2475,N_2446,N_2436);
nor U2476 (N_2476,N_2409,N_2406);
nor U2477 (N_2477,N_2422,N_2474);
nand U2478 (N_2478,N_2465,N_2413);
nor U2479 (N_2479,N_2454,N_2411);
or U2480 (N_2480,N_2407,N_2443);
and U2481 (N_2481,N_2415,N_2429);
or U2482 (N_2482,N_2417,N_2467);
and U2483 (N_2483,N_2412,N_2458);
or U2484 (N_2484,N_2452,N_2455);
or U2485 (N_2485,N_2440,N_2469);
or U2486 (N_2486,N_2444,N_2430);
and U2487 (N_2487,N_2449,N_2468);
nand U2488 (N_2488,N_2405,N_2427);
nand U2489 (N_2489,N_2441,N_2418);
or U2490 (N_2490,N_2470,N_2431);
nor U2491 (N_2491,N_2442,N_2421);
and U2492 (N_2492,N_2453,N_2447);
and U2493 (N_2493,N_2424,N_2437);
nor U2494 (N_2494,N_2460,N_2432);
nor U2495 (N_2495,N_2439,N_2400);
nand U2496 (N_2496,N_2403,N_2438);
and U2497 (N_2497,N_2456,N_2434);
nand U2498 (N_2498,N_2445,N_2426);
nor U2499 (N_2499,N_2473,N_2472);
nor U2500 (N_2500,N_2450,N_2423);
and U2501 (N_2501,N_2457,N_2408);
and U2502 (N_2502,N_2425,N_2461);
nor U2503 (N_2503,N_2419,N_2463);
nand U2504 (N_2504,N_2448,N_2433);
or U2505 (N_2505,N_2402,N_2451);
and U2506 (N_2506,N_2410,N_2464);
nand U2507 (N_2507,N_2420,N_2428);
nor U2508 (N_2508,N_2466,N_2416);
nor U2509 (N_2509,N_2435,N_2459);
nor U2510 (N_2510,N_2401,N_2414);
nor U2511 (N_2511,N_2462,N_2404);
or U2512 (N_2512,N_2471,N_2414);
or U2513 (N_2513,N_2457,N_2428);
and U2514 (N_2514,N_2441,N_2429);
and U2515 (N_2515,N_2427,N_2436);
nand U2516 (N_2516,N_2428,N_2443);
or U2517 (N_2517,N_2425,N_2455);
or U2518 (N_2518,N_2459,N_2470);
or U2519 (N_2519,N_2433,N_2434);
nor U2520 (N_2520,N_2417,N_2428);
or U2521 (N_2521,N_2464,N_2407);
nor U2522 (N_2522,N_2447,N_2405);
and U2523 (N_2523,N_2425,N_2463);
or U2524 (N_2524,N_2437,N_2405);
nand U2525 (N_2525,N_2461,N_2465);
or U2526 (N_2526,N_2404,N_2410);
nor U2527 (N_2527,N_2413,N_2471);
and U2528 (N_2528,N_2446,N_2448);
nand U2529 (N_2529,N_2426,N_2406);
or U2530 (N_2530,N_2426,N_2460);
and U2531 (N_2531,N_2430,N_2459);
and U2532 (N_2532,N_2436,N_2430);
or U2533 (N_2533,N_2419,N_2409);
nand U2534 (N_2534,N_2463,N_2472);
and U2535 (N_2535,N_2422,N_2447);
or U2536 (N_2536,N_2433,N_2429);
nor U2537 (N_2537,N_2461,N_2414);
nor U2538 (N_2538,N_2402,N_2409);
and U2539 (N_2539,N_2404,N_2413);
and U2540 (N_2540,N_2464,N_2469);
nand U2541 (N_2541,N_2434,N_2436);
or U2542 (N_2542,N_2445,N_2446);
or U2543 (N_2543,N_2415,N_2450);
nand U2544 (N_2544,N_2433,N_2422);
and U2545 (N_2545,N_2474,N_2413);
nand U2546 (N_2546,N_2452,N_2425);
nor U2547 (N_2547,N_2415,N_2420);
nand U2548 (N_2548,N_2407,N_2426);
or U2549 (N_2549,N_2439,N_2442);
nand U2550 (N_2550,N_2544,N_2497);
nand U2551 (N_2551,N_2501,N_2496);
or U2552 (N_2552,N_2529,N_2483);
and U2553 (N_2553,N_2548,N_2540);
nor U2554 (N_2554,N_2535,N_2539);
nand U2555 (N_2555,N_2503,N_2528);
nand U2556 (N_2556,N_2532,N_2487);
nand U2557 (N_2557,N_2507,N_2520);
xnor U2558 (N_2558,N_2509,N_2506);
nor U2559 (N_2559,N_2489,N_2536);
and U2560 (N_2560,N_2495,N_2543);
or U2561 (N_2561,N_2534,N_2493);
nor U2562 (N_2562,N_2476,N_2511);
or U2563 (N_2563,N_2521,N_2490);
and U2564 (N_2564,N_2475,N_2499);
nor U2565 (N_2565,N_2515,N_2542);
nor U2566 (N_2566,N_2524,N_2492);
and U2567 (N_2567,N_2498,N_2533);
nor U2568 (N_2568,N_2538,N_2549);
and U2569 (N_2569,N_2477,N_2510);
or U2570 (N_2570,N_2547,N_2526);
nand U2571 (N_2571,N_2541,N_2505);
and U2572 (N_2572,N_2518,N_2546);
or U2573 (N_2573,N_2484,N_2531);
nor U2574 (N_2574,N_2545,N_2480);
or U2575 (N_2575,N_2514,N_2479);
or U2576 (N_2576,N_2500,N_2481);
or U2577 (N_2577,N_2502,N_2491);
and U2578 (N_2578,N_2525,N_2512);
and U2579 (N_2579,N_2517,N_2513);
or U2580 (N_2580,N_2488,N_2527);
nor U2581 (N_2581,N_2516,N_2482);
or U2582 (N_2582,N_2530,N_2494);
nor U2583 (N_2583,N_2523,N_2478);
or U2584 (N_2584,N_2508,N_2485);
nand U2585 (N_2585,N_2537,N_2486);
nor U2586 (N_2586,N_2519,N_2522);
nor U2587 (N_2587,N_2504,N_2481);
nand U2588 (N_2588,N_2544,N_2534);
xor U2589 (N_2589,N_2504,N_2516);
nor U2590 (N_2590,N_2482,N_2515);
nand U2591 (N_2591,N_2544,N_2493);
nand U2592 (N_2592,N_2494,N_2511);
or U2593 (N_2593,N_2491,N_2534);
or U2594 (N_2594,N_2547,N_2543);
nor U2595 (N_2595,N_2537,N_2515);
and U2596 (N_2596,N_2541,N_2491);
and U2597 (N_2597,N_2519,N_2536);
nand U2598 (N_2598,N_2542,N_2541);
nor U2599 (N_2599,N_2482,N_2534);
or U2600 (N_2600,N_2541,N_2478);
or U2601 (N_2601,N_2501,N_2542);
or U2602 (N_2602,N_2512,N_2520);
and U2603 (N_2603,N_2544,N_2539);
nor U2604 (N_2604,N_2512,N_2507);
or U2605 (N_2605,N_2488,N_2494);
nand U2606 (N_2606,N_2545,N_2514);
nor U2607 (N_2607,N_2534,N_2521);
or U2608 (N_2608,N_2508,N_2540);
or U2609 (N_2609,N_2523,N_2513);
and U2610 (N_2610,N_2477,N_2532);
nand U2611 (N_2611,N_2487,N_2499);
or U2612 (N_2612,N_2486,N_2507);
nor U2613 (N_2613,N_2485,N_2531);
nor U2614 (N_2614,N_2547,N_2503);
and U2615 (N_2615,N_2483,N_2501);
nor U2616 (N_2616,N_2495,N_2522);
xnor U2617 (N_2617,N_2547,N_2491);
and U2618 (N_2618,N_2514,N_2530);
and U2619 (N_2619,N_2489,N_2515);
or U2620 (N_2620,N_2487,N_2536);
nand U2621 (N_2621,N_2496,N_2498);
or U2622 (N_2622,N_2500,N_2527);
nand U2623 (N_2623,N_2499,N_2489);
nand U2624 (N_2624,N_2496,N_2512);
and U2625 (N_2625,N_2565,N_2587);
or U2626 (N_2626,N_2592,N_2550);
nor U2627 (N_2627,N_2563,N_2607);
or U2628 (N_2628,N_2598,N_2551);
and U2629 (N_2629,N_2572,N_2604);
xnor U2630 (N_2630,N_2561,N_2601);
nand U2631 (N_2631,N_2588,N_2622);
or U2632 (N_2632,N_2564,N_2575);
and U2633 (N_2633,N_2624,N_2577);
or U2634 (N_2634,N_2583,N_2597);
or U2635 (N_2635,N_2556,N_2552);
nor U2636 (N_2636,N_2619,N_2616);
and U2637 (N_2637,N_2580,N_2600);
nand U2638 (N_2638,N_2566,N_2555);
nor U2639 (N_2639,N_2617,N_2620);
nor U2640 (N_2640,N_2614,N_2609);
nand U2641 (N_2641,N_2594,N_2570);
nor U2642 (N_2642,N_2590,N_2559);
xor U2643 (N_2643,N_2578,N_2603);
or U2644 (N_2644,N_2595,N_2606);
nor U2645 (N_2645,N_2613,N_2567);
nand U2646 (N_2646,N_2576,N_2612);
nor U2647 (N_2647,N_2596,N_2615);
nand U2648 (N_2648,N_2608,N_2582);
nor U2649 (N_2649,N_2618,N_2602);
nand U2650 (N_2650,N_2553,N_2610);
or U2651 (N_2651,N_2558,N_2605);
nand U2652 (N_2652,N_2557,N_2571);
nor U2653 (N_2653,N_2585,N_2581);
nand U2654 (N_2654,N_2569,N_2562);
or U2655 (N_2655,N_2621,N_2560);
nor U2656 (N_2656,N_2593,N_2574);
or U2657 (N_2657,N_2554,N_2611);
and U2658 (N_2658,N_2584,N_2579);
nor U2659 (N_2659,N_2573,N_2591);
nand U2660 (N_2660,N_2568,N_2586);
and U2661 (N_2661,N_2623,N_2589);
or U2662 (N_2662,N_2599,N_2578);
and U2663 (N_2663,N_2568,N_2582);
nor U2664 (N_2664,N_2622,N_2562);
and U2665 (N_2665,N_2558,N_2613);
nor U2666 (N_2666,N_2614,N_2556);
nand U2667 (N_2667,N_2616,N_2589);
nor U2668 (N_2668,N_2609,N_2605);
nor U2669 (N_2669,N_2592,N_2576);
nor U2670 (N_2670,N_2613,N_2560);
and U2671 (N_2671,N_2604,N_2597);
and U2672 (N_2672,N_2556,N_2618);
and U2673 (N_2673,N_2569,N_2585);
nor U2674 (N_2674,N_2584,N_2556);
nand U2675 (N_2675,N_2555,N_2584);
or U2676 (N_2676,N_2567,N_2578);
xor U2677 (N_2677,N_2581,N_2599);
xnor U2678 (N_2678,N_2620,N_2574);
or U2679 (N_2679,N_2575,N_2558);
or U2680 (N_2680,N_2576,N_2574);
or U2681 (N_2681,N_2571,N_2618);
or U2682 (N_2682,N_2621,N_2567);
and U2683 (N_2683,N_2602,N_2566);
and U2684 (N_2684,N_2621,N_2580);
nand U2685 (N_2685,N_2622,N_2595);
nor U2686 (N_2686,N_2567,N_2620);
or U2687 (N_2687,N_2614,N_2603);
nor U2688 (N_2688,N_2569,N_2556);
nand U2689 (N_2689,N_2597,N_2607);
or U2690 (N_2690,N_2559,N_2614);
or U2691 (N_2691,N_2591,N_2620);
and U2692 (N_2692,N_2590,N_2581);
nand U2693 (N_2693,N_2577,N_2588);
or U2694 (N_2694,N_2596,N_2587);
nor U2695 (N_2695,N_2594,N_2592);
nand U2696 (N_2696,N_2613,N_2608);
and U2697 (N_2697,N_2589,N_2601);
or U2698 (N_2698,N_2557,N_2586);
nand U2699 (N_2699,N_2564,N_2567);
and U2700 (N_2700,N_2675,N_2690);
nand U2701 (N_2701,N_2641,N_2665);
or U2702 (N_2702,N_2660,N_2696);
nor U2703 (N_2703,N_2653,N_2637);
and U2704 (N_2704,N_2671,N_2654);
nand U2705 (N_2705,N_2638,N_2646);
and U2706 (N_2706,N_2625,N_2670);
or U2707 (N_2707,N_2686,N_2648);
or U2708 (N_2708,N_2632,N_2673);
and U2709 (N_2709,N_2658,N_2693);
or U2710 (N_2710,N_2699,N_2628);
nor U2711 (N_2711,N_2668,N_2691);
nor U2712 (N_2712,N_2651,N_2636);
xor U2713 (N_2713,N_2682,N_2639);
nand U2714 (N_2714,N_2657,N_2672);
nand U2715 (N_2715,N_2695,N_2640);
xnor U2716 (N_2716,N_2645,N_2683);
or U2717 (N_2717,N_2688,N_2685);
and U2718 (N_2718,N_2642,N_2661);
or U2719 (N_2719,N_2629,N_2644);
nor U2720 (N_2720,N_2669,N_2647);
and U2721 (N_2721,N_2694,N_2634);
nor U2722 (N_2722,N_2687,N_2662);
or U2723 (N_2723,N_2659,N_2666);
or U2724 (N_2724,N_2635,N_2676);
or U2725 (N_2725,N_2649,N_2633);
or U2726 (N_2726,N_2692,N_2689);
and U2727 (N_2727,N_2698,N_2679);
and U2728 (N_2728,N_2627,N_2663);
or U2729 (N_2729,N_2643,N_2650);
nor U2730 (N_2730,N_2678,N_2656);
nand U2731 (N_2731,N_2681,N_2667);
and U2732 (N_2732,N_2626,N_2680);
nor U2733 (N_2733,N_2630,N_2631);
nand U2734 (N_2734,N_2664,N_2655);
nor U2735 (N_2735,N_2674,N_2677);
and U2736 (N_2736,N_2652,N_2697);
and U2737 (N_2737,N_2684,N_2685);
or U2738 (N_2738,N_2626,N_2674);
nor U2739 (N_2739,N_2676,N_2695);
nand U2740 (N_2740,N_2652,N_2675);
and U2741 (N_2741,N_2697,N_2636);
nand U2742 (N_2742,N_2661,N_2668);
or U2743 (N_2743,N_2635,N_2685);
nand U2744 (N_2744,N_2643,N_2675);
and U2745 (N_2745,N_2684,N_2626);
and U2746 (N_2746,N_2680,N_2676);
and U2747 (N_2747,N_2663,N_2660);
xor U2748 (N_2748,N_2664,N_2650);
and U2749 (N_2749,N_2674,N_2690);
and U2750 (N_2750,N_2666,N_2658);
nand U2751 (N_2751,N_2681,N_2680);
nor U2752 (N_2752,N_2633,N_2689);
nor U2753 (N_2753,N_2657,N_2699);
xor U2754 (N_2754,N_2697,N_2639);
or U2755 (N_2755,N_2661,N_2681);
nor U2756 (N_2756,N_2645,N_2662);
or U2757 (N_2757,N_2644,N_2641);
and U2758 (N_2758,N_2667,N_2690);
and U2759 (N_2759,N_2647,N_2687);
or U2760 (N_2760,N_2656,N_2663);
or U2761 (N_2761,N_2690,N_2687);
nand U2762 (N_2762,N_2629,N_2640);
nor U2763 (N_2763,N_2641,N_2680);
or U2764 (N_2764,N_2669,N_2666);
and U2765 (N_2765,N_2663,N_2648);
nor U2766 (N_2766,N_2693,N_2630);
and U2767 (N_2767,N_2670,N_2628);
or U2768 (N_2768,N_2645,N_2679);
and U2769 (N_2769,N_2627,N_2680);
or U2770 (N_2770,N_2698,N_2688);
and U2771 (N_2771,N_2679,N_2672);
or U2772 (N_2772,N_2646,N_2627);
and U2773 (N_2773,N_2660,N_2650);
and U2774 (N_2774,N_2662,N_2643);
or U2775 (N_2775,N_2756,N_2773);
or U2776 (N_2776,N_2709,N_2706);
and U2777 (N_2777,N_2762,N_2720);
nor U2778 (N_2778,N_2704,N_2749);
or U2779 (N_2779,N_2743,N_2771);
nand U2780 (N_2780,N_2738,N_2764);
and U2781 (N_2781,N_2730,N_2745);
nor U2782 (N_2782,N_2750,N_2726);
and U2783 (N_2783,N_2707,N_2754);
or U2784 (N_2784,N_2711,N_2729);
or U2785 (N_2785,N_2718,N_2716);
or U2786 (N_2786,N_2765,N_2733);
nand U2787 (N_2787,N_2742,N_2741);
nand U2788 (N_2788,N_2731,N_2753);
and U2789 (N_2789,N_2770,N_2752);
and U2790 (N_2790,N_2772,N_2736);
and U2791 (N_2791,N_2705,N_2768);
nand U2792 (N_2792,N_2763,N_2751);
nand U2793 (N_2793,N_2766,N_2725);
and U2794 (N_2794,N_2735,N_2703);
and U2795 (N_2795,N_2760,N_2722);
and U2796 (N_2796,N_2719,N_2723);
nand U2797 (N_2797,N_2755,N_2732);
or U2798 (N_2798,N_2717,N_2737);
nand U2799 (N_2799,N_2757,N_2728);
nor U2800 (N_2800,N_2701,N_2739);
or U2801 (N_2801,N_2774,N_2747);
xnor U2802 (N_2802,N_2734,N_2761);
or U2803 (N_2803,N_2744,N_2712);
or U2804 (N_2804,N_2724,N_2708);
nor U2805 (N_2805,N_2740,N_2748);
or U2806 (N_2806,N_2710,N_2769);
xor U2807 (N_2807,N_2700,N_2714);
nor U2808 (N_2808,N_2727,N_2702);
nor U2809 (N_2809,N_2746,N_2713);
nand U2810 (N_2810,N_2758,N_2767);
xnor U2811 (N_2811,N_2715,N_2721);
and U2812 (N_2812,N_2759,N_2751);
and U2813 (N_2813,N_2756,N_2734);
or U2814 (N_2814,N_2724,N_2739);
and U2815 (N_2815,N_2738,N_2747);
nor U2816 (N_2816,N_2727,N_2713);
nor U2817 (N_2817,N_2727,N_2724);
nand U2818 (N_2818,N_2737,N_2709);
nor U2819 (N_2819,N_2716,N_2714);
or U2820 (N_2820,N_2746,N_2718);
nand U2821 (N_2821,N_2757,N_2727);
or U2822 (N_2822,N_2765,N_2706);
nor U2823 (N_2823,N_2764,N_2735);
nand U2824 (N_2824,N_2725,N_2735);
and U2825 (N_2825,N_2708,N_2725);
nand U2826 (N_2826,N_2727,N_2740);
nor U2827 (N_2827,N_2729,N_2706);
nand U2828 (N_2828,N_2756,N_2736);
nor U2829 (N_2829,N_2715,N_2753);
and U2830 (N_2830,N_2761,N_2722);
and U2831 (N_2831,N_2709,N_2721);
nand U2832 (N_2832,N_2767,N_2761);
xnor U2833 (N_2833,N_2753,N_2720);
nor U2834 (N_2834,N_2718,N_2769);
and U2835 (N_2835,N_2705,N_2700);
or U2836 (N_2836,N_2764,N_2763);
nand U2837 (N_2837,N_2737,N_2731);
or U2838 (N_2838,N_2739,N_2760);
or U2839 (N_2839,N_2714,N_2713);
nand U2840 (N_2840,N_2744,N_2774);
and U2841 (N_2841,N_2721,N_2724);
and U2842 (N_2842,N_2718,N_2756);
nand U2843 (N_2843,N_2737,N_2708);
nand U2844 (N_2844,N_2731,N_2752);
and U2845 (N_2845,N_2707,N_2766);
or U2846 (N_2846,N_2753,N_2707);
or U2847 (N_2847,N_2701,N_2717);
nor U2848 (N_2848,N_2708,N_2750);
nand U2849 (N_2849,N_2754,N_2741);
and U2850 (N_2850,N_2805,N_2807);
or U2851 (N_2851,N_2819,N_2784);
nor U2852 (N_2852,N_2777,N_2804);
nand U2853 (N_2853,N_2781,N_2811);
or U2854 (N_2854,N_2793,N_2812);
and U2855 (N_2855,N_2826,N_2814);
or U2856 (N_2856,N_2836,N_2797);
nand U2857 (N_2857,N_2779,N_2790);
or U2858 (N_2858,N_2810,N_2822);
and U2859 (N_2859,N_2827,N_2833);
nor U2860 (N_2860,N_2834,N_2823);
nor U2861 (N_2861,N_2789,N_2782);
nor U2862 (N_2862,N_2813,N_2840);
nand U2863 (N_2863,N_2824,N_2828);
and U2864 (N_2864,N_2841,N_2849);
and U2865 (N_2865,N_2847,N_2788);
nor U2866 (N_2866,N_2825,N_2816);
and U2867 (N_2867,N_2815,N_2839);
or U2868 (N_2868,N_2829,N_2848);
and U2869 (N_2869,N_2785,N_2801);
nand U2870 (N_2870,N_2803,N_2796);
nor U2871 (N_2871,N_2809,N_2843);
and U2872 (N_2872,N_2791,N_2846);
nor U2873 (N_2873,N_2831,N_2786);
nor U2874 (N_2874,N_2775,N_2799);
or U2875 (N_2875,N_2798,N_2844);
and U2876 (N_2876,N_2778,N_2783);
nor U2877 (N_2877,N_2838,N_2795);
or U2878 (N_2878,N_2818,N_2787);
nor U2879 (N_2879,N_2842,N_2794);
or U2880 (N_2880,N_2776,N_2817);
and U2881 (N_2881,N_2835,N_2821);
or U2882 (N_2882,N_2806,N_2830);
or U2883 (N_2883,N_2780,N_2802);
nand U2884 (N_2884,N_2837,N_2808);
nor U2885 (N_2885,N_2832,N_2792);
nor U2886 (N_2886,N_2845,N_2820);
nor U2887 (N_2887,N_2800,N_2811);
nand U2888 (N_2888,N_2823,N_2779);
nor U2889 (N_2889,N_2796,N_2847);
or U2890 (N_2890,N_2794,N_2819);
and U2891 (N_2891,N_2801,N_2787);
or U2892 (N_2892,N_2782,N_2833);
and U2893 (N_2893,N_2794,N_2805);
and U2894 (N_2894,N_2832,N_2787);
or U2895 (N_2895,N_2831,N_2823);
nor U2896 (N_2896,N_2842,N_2822);
nand U2897 (N_2897,N_2814,N_2819);
nor U2898 (N_2898,N_2844,N_2802);
nand U2899 (N_2899,N_2846,N_2833);
and U2900 (N_2900,N_2810,N_2779);
nand U2901 (N_2901,N_2815,N_2779);
and U2902 (N_2902,N_2844,N_2836);
or U2903 (N_2903,N_2805,N_2806);
and U2904 (N_2904,N_2805,N_2776);
nor U2905 (N_2905,N_2831,N_2842);
nor U2906 (N_2906,N_2788,N_2846);
or U2907 (N_2907,N_2832,N_2794);
and U2908 (N_2908,N_2813,N_2834);
or U2909 (N_2909,N_2834,N_2802);
xor U2910 (N_2910,N_2838,N_2817);
and U2911 (N_2911,N_2841,N_2846);
and U2912 (N_2912,N_2834,N_2788);
and U2913 (N_2913,N_2811,N_2821);
nand U2914 (N_2914,N_2797,N_2787);
and U2915 (N_2915,N_2792,N_2826);
or U2916 (N_2916,N_2809,N_2810);
nand U2917 (N_2917,N_2812,N_2808);
nand U2918 (N_2918,N_2817,N_2796);
and U2919 (N_2919,N_2780,N_2782);
nand U2920 (N_2920,N_2787,N_2799);
nor U2921 (N_2921,N_2825,N_2845);
or U2922 (N_2922,N_2795,N_2801);
and U2923 (N_2923,N_2828,N_2848);
nand U2924 (N_2924,N_2821,N_2817);
nand U2925 (N_2925,N_2879,N_2870);
or U2926 (N_2926,N_2863,N_2877);
nor U2927 (N_2927,N_2866,N_2922);
and U2928 (N_2928,N_2909,N_2873);
or U2929 (N_2929,N_2902,N_2882);
and U2930 (N_2930,N_2860,N_2906);
nand U2931 (N_2931,N_2869,N_2894);
and U2932 (N_2932,N_2886,N_2903);
nor U2933 (N_2933,N_2867,N_2878);
or U2934 (N_2934,N_2900,N_2858);
and U2935 (N_2935,N_2921,N_2872);
xnor U2936 (N_2936,N_2865,N_2899);
xnor U2937 (N_2937,N_2892,N_2871);
nand U2938 (N_2938,N_2907,N_2912);
nor U2939 (N_2939,N_2853,N_2881);
nor U2940 (N_2940,N_2852,N_2893);
and U2941 (N_2941,N_2918,N_2875);
nor U2942 (N_2942,N_2889,N_2908);
or U2943 (N_2943,N_2883,N_2859);
nand U2944 (N_2944,N_2854,N_2916);
or U2945 (N_2945,N_2901,N_2861);
nor U2946 (N_2946,N_2857,N_2862);
and U2947 (N_2947,N_2888,N_2856);
and U2948 (N_2948,N_2880,N_2876);
and U2949 (N_2949,N_2919,N_2855);
nor U2950 (N_2950,N_2850,N_2885);
nor U2951 (N_2951,N_2868,N_2898);
nand U2952 (N_2952,N_2890,N_2887);
and U2953 (N_2953,N_2911,N_2905);
or U2954 (N_2954,N_2896,N_2915);
nor U2955 (N_2955,N_2920,N_2924);
nand U2956 (N_2956,N_2910,N_2897);
nand U2957 (N_2957,N_2904,N_2895);
nand U2958 (N_2958,N_2874,N_2923);
and U2959 (N_2959,N_2917,N_2864);
or U2960 (N_2960,N_2914,N_2851);
or U2961 (N_2961,N_2891,N_2884);
and U2962 (N_2962,N_2913,N_2895);
and U2963 (N_2963,N_2908,N_2911);
xnor U2964 (N_2964,N_2876,N_2888);
nand U2965 (N_2965,N_2907,N_2866);
nand U2966 (N_2966,N_2869,N_2858);
and U2967 (N_2967,N_2891,N_2893);
or U2968 (N_2968,N_2902,N_2870);
nor U2969 (N_2969,N_2896,N_2875);
or U2970 (N_2970,N_2861,N_2863);
nand U2971 (N_2971,N_2920,N_2852);
nor U2972 (N_2972,N_2902,N_2891);
or U2973 (N_2973,N_2865,N_2888);
or U2974 (N_2974,N_2913,N_2864);
or U2975 (N_2975,N_2890,N_2921);
nand U2976 (N_2976,N_2906,N_2861);
nor U2977 (N_2977,N_2893,N_2920);
nand U2978 (N_2978,N_2880,N_2860);
nor U2979 (N_2979,N_2852,N_2866);
nor U2980 (N_2980,N_2851,N_2886);
and U2981 (N_2981,N_2860,N_2912);
and U2982 (N_2982,N_2900,N_2922);
or U2983 (N_2983,N_2876,N_2855);
or U2984 (N_2984,N_2912,N_2867);
nor U2985 (N_2985,N_2857,N_2905);
nand U2986 (N_2986,N_2866,N_2869);
nand U2987 (N_2987,N_2870,N_2853);
and U2988 (N_2988,N_2876,N_2869);
nor U2989 (N_2989,N_2873,N_2882);
or U2990 (N_2990,N_2917,N_2901);
or U2991 (N_2991,N_2852,N_2873);
or U2992 (N_2992,N_2868,N_2908);
or U2993 (N_2993,N_2901,N_2900);
nor U2994 (N_2994,N_2918,N_2863);
nand U2995 (N_2995,N_2855,N_2852);
nor U2996 (N_2996,N_2852,N_2896);
and U2997 (N_2997,N_2922,N_2851);
nor U2998 (N_2998,N_2859,N_2860);
or U2999 (N_2999,N_2923,N_2881);
nor UO_0 (O_0,N_2958,N_2952);
or UO_1 (O_1,N_2960,N_2964);
nor UO_2 (O_2,N_2957,N_2988);
nand UO_3 (O_3,N_2962,N_2925);
and UO_4 (O_4,N_2966,N_2932);
nand UO_5 (O_5,N_2998,N_2986);
nand UO_6 (O_6,N_2955,N_2977);
or UO_7 (O_7,N_2963,N_2967);
nand UO_8 (O_8,N_2975,N_2979);
nor UO_9 (O_9,N_2965,N_2978);
nor UO_10 (O_10,N_2992,N_2999);
or UO_11 (O_11,N_2972,N_2985);
and UO_12 (O_12,N_2940,N_2989);
nand UO_13 (O_13,N_2997,N_2931);
nand UO_14 (O_14,N_2974,N_2982);
or UO_15 (O_15,N_2950,N_2980);
nand UO_16 (O_16,N_2944,N_2943);
nor UO_17 (O_17,N_2946,N_2926);
nor UO_18 (O_18,N_2983,N_2971);
nor UO_19 (O_19,N_2969,N_2945);
nor UO_20 (O_20,N_2973,N_2991);
and UO_21 (O_21,N_2947,N_2995);
and UO_22 (O_22,N_2927,N_2953);
or UO_23 (O_23,N_2961,N_2956);
nand UO_24 (O_24,N_2937,N_2941);
or UO_25 (O_25,N_2981,N_2993);
and UO_26 (O_26,N_2949,N_2935);
nand UO_27 (O_27,N_2984,N_2959);
nand UO_28 (O_28,N_2948,N_2929);
nand UO_29 (O_29,N_2939,N_2987);
nor UO_30 (O_30,N_2936,N_2994);
or UO_31 (O_31,N_2938,N_2933);
or UO_32 (O_32,N_2942,N_2968);
or UO_33 (O_33,N_2954,N_2951);
nor UO_34 (O_34,N_2976,N_2928);
nand UO_35 (O_35,N_2996,N_2970);
nor UO_36 (O_36,N_2934,N_2990);
and UO_37 (O_37,N_2930,N_2932);
or UO_38 (O_38,N_2940,N_2974);
nand UO_39 (O_39,N_2927,N_2999);
and UO_40 (O_40,N_2941,N_2954);
or UO_41 (O_41,N_2934,N_2941);
or UO_42 (O_42,N_2928,N_2968);
nor UO_43 (O_43,N_2933,N_2960);
and UO_44 (O_44,N_2929,N_2998);
nand UO_45 (O_45,N_2951,N_2940);
nor UO_46 (O_46,N_2997,N_2951);
nor UO_47 (O_47,N_2948,N_2988);
or UO_48 (O_48,N_2991,N_2960);
nand UO_49 (O_49,N_2948,N_2931);
and UO_50 (O_50,N_2956,N_2960);
and UO_51 (O_51,N_2972,N_2975);
nor UO_52 (O_52,N_2984,N_2980);
or UO_53 (O_53,N_2949,N_2941);
xor UO_54 (O_54,N_2930,N_2994);
nor UO_55 (O_55,N_2949,N_2944);
or UO_56 (O_56,N_2992,N_2932);
or UO_57 (O_57,N_2935,N_2940);
nor UO_58 (O_58,N_2955,N_2932);
nand UO_59 (O_59,N_2961,N_2973);
nand UO_60 (O_60,N_2948,N_2982);
and UO_61 (O_61,N_2951,N_2976);
nand UO_62 (O_62,N_2978,N_2952);
or UO_63 (O_63,N_2931,N_2965);
and UO_64 (O_64,N_2938,N_2932);
and UO_65 (O_65,N_2936,N_2983);
nor UO_66 (O_66,N_2995,N_2927);
nor UO_67 (O_67,N_2991,N_2999);
nor UO_68 (O_68,N_2987,N_2956);
and UO_69 (O_69,N_2943,N_2950);
and UO_70 (O_70,N_2941,N_2944);
nand UO_71 (O_71,N_2953,N_2957);
or UO_72 (O_72,N_2950,N_2984);
and UO_73 (O_73,N_2973,N_2954);
and UO_74 (O_74,N_2969,N_2985);
nand UO_75 (O_75,N_2972,N_2940);
nand UO_76 (O_76,N_2980,N_2998);
or UO_77 (O_77,N_2928,N_2926);
xor UO_78 (O_78,N_2946,N_2995);
or UO_79 (O_79,N_2953,N_2949);
and UO_80 (O_80,N_2998,N_2937);
nor UO_81 (O_81,N_2966,N_2995);
nor UO_82 (O_82,N_2926,N_2934);
and UO_83 (O_83,N_2938,N_2976);
nor UO_84 (O_84,N_2940,N_2942);
nand UO_85 (O_85,N_2959,N_2940);
nor UO_86 (O_86,N_2987,N_2978);
and UO_87 (O_87,N_2952,N_2990);
nand UO_88 (O_88,N_2971,N_2935);
or UO_89 (O_89,N_2981,N_2990);
or UO_90 (O_90,N_2969,N_2929);
or UO_91 (O_91,N_2962,N_2953);
and UO_92 (O_92,N_2931,N_2980);
or UO_93 (O_93,N_2948,N_2978);
nand UO_94 (O_94,N_2927,N_2943);
and UO_95 (O_95,N_2948,N_2938);
and UO_96 (O_96,N_2973,N_2979);
nor UO_97 (O_97,N_2952,N_2994);
and UO_98 (O_98,N_2988,N_2944);
nand UO_99 (O_99,N_2985,N_2925);
nand UO_100 (O_100,N_2952,N_2972);
or UO_101 (O_101,N_2969,N_2951);
xor UO_102 (O_102,N_2932,N_2975);
nor UO_103 (O_103,N_2936,N_2938);
and UO_104 (O_104,N_2930,N_2959);
nor UO_105 (O_105,N_2983,N_2987);
nor UO_106 (O_106,N_2928,N_2937);
nand UO_107 (O_107,N_2994,N_2972);
or UO_108 (O_108,N_2975,N_2940);
and UO_109 (O_109,N_2991,N_2965);
or UO_110 (O_110,N_2946,N_2943);
nor UO_111 (O_111,N_2992,N_2930);
nor UO_112 (O_112,N_2983,N_2982);
or UO_113 (O_113,N_2980,N_2972);
nor UO_114 (O_114,N_2958,N_2944);
nand UO_115 (O_115,N_2934,N_2935);
and UO_116 (O_116,N_2996,N_2951);
nor UO_117 (O_117,N_2978,N_2983);
nand UO_118 (O_118,N_2953,N_2998);
nand UO_119 (O_119,N_2980,N_2990);
and UO_120 (O_120,N_2974,N_2956);
and UO_121 (O_121,N_2942,N_2950);
and UO_122 (O_122,N_2931,N_2985);
or UO_123 (O_123,N_2949,N_2963);
and UO_124 (O_124,N_2974,N_2958);
nor UO_125 (O_125,N_2997,N_2943);
and UO_126 (O_126,N_2940,N_2986);
nand UO_127 (O_127,N_2984,N_2947);
nor UO_128 (O_128,N_2952,N_2979);
or UO_129 (O_129,N_2935,N_2957);
or UO_130 (O_130,N_2934,N_2939);
and UO_131 (O_131,N_2976,N_2950);
nand UO_132 (O_132,N_2965,N_2959);
nor UO_133 (O_133,N_2970,N_2977);
nor UO_134 (O_134,N_2988,N_2983);
nor UO_135 (O_135,N_2964,N_2966);
and UO_136 (O_136,N_2965,N_2992);
nand UO_137 (O_137,N_2968,N_2988);
nand UO_138 (O_138,N_2950,N_2949);
or UO_139 (O_139,N_2996,N_2974);
or UO_140 (O_140,N_2950,N_2931);
or UO_141 (O_141,N_2968,N_2962);
nor UO_142 (O_142,N_2934,N_2991);
or UO_143 (O_143,N_2930,N_2984);
or UO_144 (O_144,N_2944,N_2984);
or UO_145 (O_145,N_2936,N_2990);
nor UO_146 (O_146,N_2953,N_2977);
and UO_147 (O_147,N_2961,N_2997);
nor UO_148 (O_148,N_2939,N_2954);
nor UO_149 (O_149,N_2940,N_2995);
nor UO_150 (O_150,N_2938,N_2944);
or UO_151 (O_151,N_2950,N_2933);
nand UO_152 (O_152,N_2947,N_2952);
and UO_153 (O_153,N_2952,N_2943);
nand UO_154 (O_154,N_2934,N_2947);
or UO_155 (O_155,N_2931,N_2975);
nor UO_156 (O_156,N_2963,N_2985);
or UO_157 (O_157,N_2977,N_2959);
nor UO_158 (O_158,N_2945,N_2936);
and UO_159 (O_159,N_2952,N_2946);
xnor UO_160 (O_160,N_2964,N_2994);
nand UO_161 (O_161,N_2970,N_2998);
nor UO_162 (O_162,N_2933,N_2931);
and UO_163 (O_163,N_2939,N_2978);
or UO_164 (O_164,N_2997,N_2974);
nand UO_165 (O_165,N_2985,N_2983);
nand UO_166 (O_166,N_2973,N_2932);
nand UO_167 (O_167,N_2973,N_2970);
and UO_168 (O_168,N_2942,N_2978);
nand UO_169 (O_169,N_2952,N_2951);
and UO_170 (O_170,N_2928,N_2927);
nand UO_171 (O_171,N_2988,N_2978);
or UO_172 (O_172,N_2950,N_2975);
and UO_173 (O_173,N_2954,N_2952);
nand UO_174 (O_174,N_2999,N_2951);
nand UO_175 (O_175,N_2953,N_2983);
nand UO_176 (O_176,N_2966,N_2974);
and UO_177 (O_177,N_2963,N_2992);
nand UO_178 (O_178,N_2997,N_2964);
nor UO_179 (O_179,N_2948,N_2975);
nand UO_180 (O_180,N_2951,N_2932);
and UO_181 (O_181,N_2970,N_2930);
nand UO_182 (O_182,N_2938,N_2993);
nor UO_183 (O_183,N_2997,N_2955);
nand UO_184 (O_184,N_2956,N_2970);
nor UO_185 (O_185,N_2985,N_2993);
and UO_186 (O_186,N_2947,N_2963);
and UO_187 (O_187,N_2961,N_2933);
or UO_188 (O_188,N_2989,N_2995);
and UO_189 (O_189,N_2979,N_2935);
xor UO_190 (O_190,N_2964,N_2952);
or UO_191 (O_191,N_2945,N_2972);
nand UO_192 (O_192,N_2974,N_2973);
nand UO_193 (O_193,N_2952,N_2968);
xor UO_194 (O_194,N_2944,N_2995);
or UO_195 (O_195,N_2927,N_2941);
nand UO_196 (O_196,N_2954,N_2932);
nor UO_197 (O_197,N_2954,N_2938);
nor UO_198 (O_198,N_2979,N_2933);
nor UO_199 (O_199,N_2930,N_2999);
or UO_200 (O_200,N_2944,N_2939);
and UO_201 (O_201,N_2980,N_2944);
nor UO_202 (O_202,N_2992,N_2964);
nor UO_203 (O_203,N_2933,N_2983);
and UO_204 (O_204,N_2983,N_2962);
and UO_205 (O_205,N_2983,N_2948);
nor UO_206 (O_206,N_2960,N_2970);
nand UO_207 (O_207,N_2933,N_2990);
nand UO_208 (O_208,N_2943,N_2938);
nand UO_209 (O_209,N_2926,N_2986);
or UO_210 (O_210,N_2992,N_2967);
nor UO_211 (O_211,N_2972,N_2937);
nor UO_212 (O_212,N_2969,N_2976);
nand UO_213 (O_213,N_2925,N_2927);
and UO_214 (O_214,N_2956,N_2959);
and UO_215 (O_215,N_2979,N_2980);
and UO_216 (O_216,N_2966,N_2968);
and UO_217 (O_217,N_2990,N_2932);
nor UO_218 (O_218,N_2998,N_2938);
and UO_219 (O_219,N_2972,N_2968);
or UO_220 (O_220,N_2983,N_2937);
nand UO_221 (O_221,N_2986,N_2969);
nor UO_222 (O_222,N_2996,N_2944);
and UO_223 (O_223,N_2952,N_2983);
nor UO_224 (O_224,N_2978,N_2998);
or UO_225 (O_225,N_2946,N_2954);
nand UO_226 (O_226,N_2925,N_2947);
or UO_227 (O_227,N_2936,N_2996);
nor UO_228 (O_228,N_2988,N_2936);
and UO_229 (O_229,N_2955,N_2966);
and UO_230 (O_230,N_2996,N_2983);
or UO_231 (O_231,N_2946,N_2962);
or UO_232 (O_232,N_2959,N_2986);
and UO_233 (O_233,N_2953,N_2926);
nand UO_234 (O_234,N_2952,N_2935);
nor UO_235 (O_235,N_2973,N_2935);
nor UO_236 (O_236,N_2986,N_2979);
or UO_237 (O_237,N_2990,N_2998);
nand UO_238 (O_238,N_2979,N_2995);
nand UO_239 (O_239,N_2958,N_2983);
and UO_240 (O_240,N_2971,N_2980);
nand UO_241 (O_241,N_2963,N_2946);
and UO_242 (O_242,N_2954,N_2984);
or UO_243 (O_243,N_2964,N_2978);
and UO_244 (O_244,N_2932,N_2931);
or UO_245 (O_245,N_2968,N_2979);
nand UO_246 (O_246,N_2957,N_2971);
nand UO_247 (O_247,N_2951,N_2977);
nor UO_248 (O_248,N_2928,N_2950);
and UO_249 (O_249,N_2985,N_2948);
xor UO_250 (O_250,N_2992,N_2971);
nand UO_251 (O_251,N_2976,N_2982);
or UO_252 (O_252,N_2933,N_2946);
nor UO_253 (O_253,N_2988,N_2979);
nor UO_254 (O_254,N_2976,N_2931);
nand UO_255 (O_255,N_2933,N_2958);
and UO_256 (O_256,N_2964,N_2926);
nor UO_257 (O_257,N_2927,N_2934);
and UO_258 (O_258,N_2934,N_2963);
or UO_259 (O_259,N_2948,N_2986);
nand UO_260 (O_260,N_2949,N_2933);
nor UO_261 (O_261,N_2967,N_2982);
nand UO_262 (O_262,N_2965,N_2985);
xor UO_263 (O_263,N_2972,N_2982);
or UO_264 (O_264,N_2933,N_2998);
and UO_265 (O_265,N_2955,N_2976);
xor UO_266 (O_266,N_2966,N_2952);
or UO_267 (O_267,N_2958,N_2960);
xnor UO_268 (O_268,N_2936,N_2982);
nand UO_269 (O_269,N_2975,N_2983);
nor UO_270 (O_270,N_2925,N_2975);
or UO_271 (O_271,N_2951,N_2987);
nand UO_272 (O_272,N_2989,N_2935);
and UO_273 (O_273,N_2982,N_2980);
and UO_274 (O_274,N_2965,N_2960);
nand UO_275 (O_275,N_2937,N_2934);
nand UO_276 (O_276,N_2956,N_2932);
and UO_277 (O_277,N_2965,N_2943);
or UO_278 (O_278,N_2979,N_2947);
nor UO_279 (O_279,N_2983,N_2998);
and UO_280 (O_280,N_2999,N_2978);
nor UO_281 (O_281,N_2999,N_2983);
or UO_282 (O_282,N_2954,N_2936);
or UO_283 (O_283,N_2951,N_2942);
and UO_284 (O_284,N_2983,N_2992);
nand UO_285 (O_285,N_2986,N_2932);
nor UO_286 (O_286,N_2975,N_2974);
nor UO_287 (O_287,N_2948,N_2979);
and UO_288 (O_288,N_2949,N_2998);
and UO_289 (O_289,N_2930,N_2966);
nand UO_290 (O_290,N_2956,N_2965);
nand UO_291 (O_291,N_2970,N_2971);
and UO_292 (O_292,N_2934,N_2946);
nor UO_293 (O_293,N_2961,N_2953);
nor UO_294 (O_294,N_2985,N_2966);
or UO_295 (O_295,N_2956,N_2948);
nor UO_296 (O_296,N_2952,N_2961);
or UO_297 (O_297,N_2956,N_2988);
nand UO_298 (O_298,N_2952,N_2930);
xor UO_299 (O_299,N_2962,N_2949);
nor UO_300 (O_300,N_2944,N_2940);
or UO_301 (O_301,N_2958,N_2981);
and UO_302 (O_302,N_2944,N_2993);
nand UO_303 (O_303,N_2984,N_2955);
or UO_304 (O_304,N_2995,N_2999);
xnor UO_305 (O_305,N_2990,N_2963);
or UO_306 (O_306,N_2979,N_2949);
nor UO_307 (O_307,N_2999,N_2947);
nand UO_308 (O_308,N_2925,N_2960);
and UO_309 (O_309,N_2930,N_2956);
nand UO_310 (O_310,N_2925,N_2973);
nand UO_311 (O_311,N_2957,N_2961);
and UO_312 (O_312,N_2962,N_2970);
nand UO_313 (O_313,N_2948,N_2932);
nand UO_314 (O_314,N_2934,N_2955);
and UO_315 (O_315,N_2965,N_2947);
nand UO_316 (O_316,N_2958,N_2993);
and UO_317 (O_317,N_2971,N_2930);
or UO_318 (O_318,N_2963,N_2975);
or UO_319 (O_319,N_2944,N_2983);
or UO_320 (O_320,N_2984,N_2981);
xnor UO_321 (O_321,N_2994,N_2976);
and UO_322 (O_322,N_2986,N_2991);
nor UO_323 (O_323,N_2968,N_2956);
or UO_324 (O_324,N_2999,N_2966);
or UO_325 (O_325,N_2931,N_2955);
nor UO_326 (O_326,N_2944,N_2969);
and UO_327 (O_327,N_2981,N_2955);
or UO_328 (O_328,N_2985,N_2946);
nand UO_329 (O_329,N_2931,N_2944);
nand UO_330 (O_330,N_2980,N_2978);
and UO_331 (O_331,N_2998,N_2960);
nand UO_332 (O_332,N_2951,N_2947);
and UO_333 (O_333,N_2953,N_2960);
and UO_334 (O_334,N_2942,N_2976);
nand UO_335 (O_335,N_2945,N_2990);
and UO_336 (O_336,N_2976,N_2964);
or UO_337 (O_337,N_2982,N_2957);
and UO_338 (O_338,N_2953,N_2950);
nor UO_339 (O_339,N_2938,N_2992);
nand UO_340 (O_340,N_2960,N_2946);
nor UO_341 (O_341,N_2970,N_2961);
and UO_342 (O_342,N_2992,N_2995);
and UO_343 (O_343,N_2933,N_2981);
or UO_344 (O_344,N_2933,N_2951);
nand UO_345 (O_345,N_2957,N_2981);
nor UO_346 (O_346,N_2968,N_2963);
nor UO_347 (O_347,N_2926,N_2960);
nand UO_348 (O_348,N_2963,N_2952);
nand UO_349 (O_349,N_2938,N_2942);
and UO_350 (O_350,N_2970,N_2958);
nor UO_351 (O_351,N_2965,N_2949);
nor UO_352 (O_352,N_2979,N_2965);
nand UO_353 (O_353,N_2979,N_2969);
nor UO_354 (O_354,N_2969,N_2989);
or UO_355 (O_355,N_2971,N_2965);
nand UO_356 (O_356,N_2961,N_2985);
and UO_357 (O_357,N_2939,N_2970);
nor UO_358 (O_358,N_2960,N_2967);
and UO_359 (O_359,N_2971,N_2933);
nor UO_360 (O_360,N_2963,N_2988);
nor UO_361 (O_361,N_2939,N_2985);
nor UO_362 (O_362,N_2981,N_2967);
nor UO_363 (O_363,N_2994,N_2982);
nor UO_364 (O_364,N_2980,N_2995);
nand UO_365 (O_365,N_2951,N_2963);
and UO_366 (O_366,N_2966,N_2960);
or UO_367 (O_367,N_2972,N_2963);
xor UO_368 (O_368,N_2953,N_2939);
or UO_369 (O_369,N_2956,N_2969);
nand UO_370 (O_370,N_2992,N_2937);
or UO_371 (O_371,N_2989,N_2929);
nand UO_372 (O_372,N_2989,N_2998);
nor UO_373 (O_373,N_2938,N_2927);
nor UO_374 (O_374,N_2961,N_2967);
or UO_375 (O_375,N_2992,N_2986);
and UO_376 (O_376,N_2946,N_2945);
nand UO_377 (O_377,N_2934,N_2985);
nor UO_378 (O_378,N_2945,N_2933);
or UO_379 (O_379,N_2991,N_2930);
and UO_380 (O_380,N_2981,N_2999);
nand UO_381 (O_381,N_2951,N_2975);
nand UO_382 (O_382,N_2943,N_2967);
nor UO_383 (O_383,N_2999,N_2980);
or UO_384 (O_384,N_2957,N_2939);
nor UO_385 (O_385,N_2948,N_2951);
nor UO_386 (O_386,N_2945,N_2953);
or UO_387 (O_387,N_2984,N_2968);
nand UO_388 (O_388,N_2971,N_2991);
or UO_389 (O_389,N_2995,N_2983);
or UO_390 (O_390,N_2937,N_2999);
nand UO_391 (O_391,N_2929,N_2938);
nor UO_392 (O_392,N_2931,N_2978);
nor UO_393 (O_393,N_2956,N_2977);
xnor UO_394 (O_394,N_2986,N_2947);
and UO_395 (O_395,N_2990,N_2946);
and UO_396 (O_396,N_2926,N_2944);
and UO_397 (O_397,N_2942,N_2929);
or UO_398 (O_398,N_2982,N_2997);
nand UO_399 (O_399,N_2960,N_2988);
xor UO_400 (O_400,N_2925,N_2990);
nor UO_401 (O_401,N_2928,N_2983);
or UO_402 (O_402,N_2960,N_2982);
or UO_403 (O_403,N_2958,N_2948);
or UO_404 (O_404,N_2942,N_2955);
or UO_405 (O_405,N_2928,N_2998);
and UO_406 (O_406,N_2929,N_2986);
or UO_407 (O_407,N_2938,N_2973);
nor UO_408 (O_408,N_2941,N_2980);
nor UO_409 (O_409,N_2966,N_2984);
and UO_410 (O_410,N_2928,N_2986);
or UO_411 (O_411,N_2949,N_2972);
or UO_412 (O_412,N_2992,N_2954);
nor UO_413 (O_413,N_2944,N_2966);
nand UO_414 (O_414,N_2999,N_2931);
nor UO_415 (O_415,N_2998,N_2943);
or UO_416 (O_416,N_2953,N_2996);
or UO_417 (O_417,N_2962,N_2964);
and UO_418 (O_418,N_2990,N_2964);
or UO_419 (O_419,N_2945,N_2963);
nor UO_420 (O_420,N_2979,N_2962);
nor UO_421 (O_421,N_2987,N_2971);
and UO_422 (O_422,N_2957,N_2950);
nor UO_423 (O_423,N_2948,N_2996);
nor UO_424 (O_424,N_2963,N_2978);
nand UO_425 (O_425,N_2940,N_2929);
nand UO_426 (O_426,N_2944,N_2994);
nor UO_427 (O_427,N_2945,N_2927);
nand UO_428 (O_428,N_2977,N_2939);
and UO_429 (O_429,N_2934,N_2932);
and UO_430 (O_430,N_2946,N_2973);
and UO_431 (O_431,N_2957,N_2944);
or UO_432 (O_432,N_2956,N_2999);
xor UO_433 (O_433,N_2971,N_2979);
nor UO_434 (O_434,N_2974,N_2985);
and UO_435 (O_435,N_2992,N_2998);
nand UO_436 (O_436,N_2976,N_2966);
nand UO_437 (O_437,N_2951,N_2970);
and UO_438 (O_438,N_2925,N_2955);
or UO_439 (O_439,N_2949,N_2959);
nand UO_440 (O_440,N_2943,N_2960);
and UO_441 (O_441,N_2950,N_2995);
nor UO_442 (O_442,N_2987,N_2995);
or UO_443 (O_443,N_2990,N_2967);
or UO_444 (O_444,N_2960,N_2927);
or UO_445 (O_445,N_2926,N_2991);
and UO_446 (O_446,N_2965,N_2944);
nand UO_447 (O_447,N_2972,N_2990);
or UO_448 (O_448,N_2980,N_2976);
nor UO_449 (O_449,N_2977,N_2988);
nand UO_450 (O_450,N_2928,N_2970);
nand UO_451 (O_451,N_2998,N_2963);
nand UO_452 (O_452,N_2939,N_2946);
and UO_453 (O_453,N_2989,N_2974);
nor UO_454 (O_454,N_2985,N_2945);
xor UO_455 (O_455,N_2969,N_2974);
and UO_456 (O_456,N_2994,N_2942);
or UO_457 (O_457,N_2982,N_2966);
xor UO_458 (O_458,N_2993,N_2978);
nor UO_459 (O_459,N_2991,N_2978);
nand UO_460 (O_460,N_2942,N_2995);
and UO_461 (O_461,N_2979,N_2964);
and UO_462 (O_462,N_2978,N_2992);
or UO_463 (O_463,N_2975,N_2978);
or UO_464 (O_464,N_2968,N_2929);
xor UO_465 (O_465,N_2998,N_2956);
and UO_466 (O_466,N_2995,N_2988);
and UO_467 (O_467,N_2937,N_2944);
and UO_468 (O_468,N_2952,N_2981);
or UO_469 (O_469,N_2925,N_2982);
nor UO_470 (O_470,N_2965,N_2998);
nor UO_471 (O_471,N_2941,N_2990);
or UO_472 (O_472,N_2983,N_2946);
nor UO_473 (O_473,N_2978,N_2925);
and UO_474 (O_474,N_2929,N_2958);
and UO_475 (O_475,N_2993,N_2925);
nor UO_476 (O_476,N_2936,N_2979);
or UO_477 (O_477,N_2949,N_2946);
nand UO_478 (O_478,N_2983,N_2938);
nand UO_479 (O_479,N_2982,N_2977);
or UO_480 (O_480,N_2942,N_2980);
and UO_481 (O_481,N_2973,N_2953);
xor UO_482 (O_482,N_2996,N_2931);
and UO_483 (O_483,N_2949,N_2955);
or UO_484 (O_484,N_2926,N_2925);
nor UO_485 (O_485,N_2985,N_2936);
nand UO_486 (O_486,N_2973,N_2943);
nor UO_487 (O_487,N_2986,N_2936);
and UO_488 (O_488,N_2947,N_2980);
nand UO_489 (O_489,N_2942,N_2926);
and UO_490 (O_490,N_2979,N_2929);
or UO_491 (O_491,N_2926,N_2976);
or UO_492 (O_492,N_2949,N_2987);
nor UO_493 (O_493,N_2997,N_2939);
nand UO_494 (O_494,N_2957,N_2955);
and UO_495 (O_495,N_2966,N_2959);
or UO_496 (O_496,N_2938,N_2926);
nor UO_497 (O_497,N_2956,N_2929);
and UO_498 (O_498,N_2977,N_2993);
nor UO_499 (O_499,N_2945,N_2940);
endmodule