module basic_1500_15000_2000_15_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_935,In_176);
and U1 (N_1,In_867,In_668);
or U2 (N_2,In_1117,In_1377);
or U3 (N_3,In_1242,In_308);
and U4 (N_4,In_798,In_158);
nor U5 (N_5,In_173,In_315);
and U6 (N_6,In_1128,In_43);
or U7 (N_7,In_889,In_672);
and U8 (N_8,In_351,In_575);
xor U9 (N_9,In_1475,In_1032);
xnor U10 (N_10,In_13,In_615);
and U11 (N_11,In_1161,In_451);
or U12 (N_12,In_390,In_535);
nand U13 (N_13,In_807,In_1402);
nor U14 (N_14,In_311,In_322);
or U15 (N_15,In_374,In_826);
nor U16 (N_16,In_104,In_1290);
xnor U17 (N_17,In_1422,In_1202);
xor U18 (N_18,In_1177,In_1064);
nor U19 (N_19,In_181,In_458);
nand U20 (N_20,In_248,In_1237);
nand U21 (N_21,In_1364,In_1277);
or U22 (N_22,In_369,In_1391);
or U23 (N_23,In_1266,In_534);
nand U24 (N_24,In_985,In_671);
nand U25 (N_25,In_942,In_790);
nand U26 (N_26,In_992,In_1334);
or U27 (N_27,In_366,In_1424);
and U28 (N_28,In_258,In_1447);
nor U29 (N_29,In_741,In_268);
nor U30 (N_30,In_1168,In_1122);
xor U31 (N_31,In_878,In_1390);
nand U32 (N_32,In_519,In_1256);
nor U33 (N_33,In_674,In_170);
or U34 (N_34,In_513,In_302);
nor U35 (N_35,In_250,In_1329);
and U36 (N_36,In_617,In_404);
nor U37 (N_37,In_386,In_740);
xnor U38 (N_38,In_1164,In_1467);
nor U39 (N_39,In_205,In_953);
nor U40 (N_40,In_445,In_321);
and U41 (N_41,In_1121,In_1474);
and U42 (N_42,In_262,In_33);
xnor U43 (N_43,In_1248,In_1131);
xor U44 (N_44,In_304,In_1196);
or U45 (N_45,In_1144,In_742);
nand U46 (N_46,In_324,In_1332);
and U47 (N_47,In_1333,In_138);
or U48 (N_48,In_466,In_804);
nor U49 (N_49,In_578,In_845);
or U50 (N_50,In_773,In_212);
or U51 (N_51,In_666,In_385);
or U52 (N_52,In_616,In_726);
and U53 (N_53,In_1240,In_633);
nand U54 (N_54,In_518,In_1407);
nand U55 (N_55,In_1146,In_236);
xor U56 (N_56,In_541,In_1452);
nor U57 (N_57,In_1254,In_344);
nand U58 (N_58,In_689,In_673);
nand U59 (N_59,In_407,In_749);
or U60 (N_60,In_787,In_101);
or U61 (N_61,In_995,In_871);
or U62 (N_62,In_36,In_486);
and U63 (N_63,In_1001,In_1033);
nor U64 (N_64,In_405,In_1035);
and U65 (N_65,In_1220,In_201);
nor U66 (N_66,In_166,In_1318);
nand U67 (N_67,In_1116,In_148);
or U68 (N_68,In_903,In_493);
xnor U69 (N_69,In_877,In_572);
or U70 (N_70,In_610,In_1322);
or U71 (N_71,In_1173,In_940);
and U72 (N_72,In_454,In_1295);
and U73 (N_73,In_1478,In_630);
nand U74 (N_74,In_1065,In_1142);
xnor U75 (N_75,In_655,In_664);
and U76 (N_76,In_766,In_1075);
and U77 (N_77,In_1100,In_930);
nor U78 (N_78,In_890,In_881);
nor U79 (N_79,In_844,In_542);
and U80 (N_80,In_1021,In_1313);
or U81 (N_81,In_135,In_154);
or U82 (N_82,In_1077,In_1463);
and U83 (N_83,In_1355,In_478);
nand U84 (N_84,In_1468,In_1388);
nor U85 (N_85,In_342,In_932);
or U86 (N_86,In_1190,In_1079);
nor U87 (N_87,In_1280,In_1425);
and U88 (N_88,In_720,In_159);
or U89 (N_89,In_1345,In_1435);
xnor U90 (N_90,In_1323,In_708);
nand U91 (N_91,In_208,In_1484);
nor U92 (N_92,In_241,In_1274);
nor U93 (N_93,In_1238,In_169);
and U94 (N_94,In_1357,In_294);
nor U95 (N_95,In_437,In_243);
nand U96 (N_96,In_937,In_913);
or U97 (N_97,In_1119,In_783);
nor U98 (N_98,In_533,In_1459);
nor U99 (N_99,In_511,In_204);
nor U100 (N_100,In_363,In_996);
nand U101 (N_101,In_1171,In_450);
nand U102 (N_102,In_748,In_1465);
nor U103 (N_103,In_719,In_1443);
xor U104 (N_104,In_131,In_382);
or U105 (N_105,In_1051,In_866);
or U106 (N_106,In_834,In_207);
nor U107 (N_107,In_143,In_1108);
nand U108 (N_108,In_1175,In_1047);
nor U109 (N_109,In_1304,In_288);
nand U110 (N_110,In_603,In_1339);
or U111 (N_111,In_232,In_239);
and U112 (N_112,In_1412,In_191);
and U113 (N_113,In_147,In_1136);
nor U114 (N_114,In_1058,In_1192);
and U115 (N_115,In_987,In_141);
nor U116 (N_116,In_1247,In_1342);
nand U117 (N_117,In_216,In_669);
and U118 (N_118,In_563,In_904);
or U119 (N_119,In_32,In_1034);
nor U120 (N_120,In_576,In_1103);
nand U121 (N_121,In_957,In_1135);
and U122 (N_122,In_984,In_361);
nor U123 (N_123,In_403,In_1480);
or U124 (N_124,In_416,In_53);
and U125 (N_125,In_1036,In_1227);
nor U126 (N_126,In_730,In_125);
xor U127 (N_127,In_958,In_851);
and U128 (N_128,In_1455,In_1004);
or U129 (N_129,In_1385,In_1260);
or U130 (N_130,In_22,In_156);
nor U131 (N_131,In_811,In_5);
and U132 (N_132,In_1104,In_1207);
nor U133 (N_133,In_92,In_298);
and U134 (N_134,In_571,In_246);
nand U135 (N_135,In_864,In_1160);
or U136 (N_136,In_1460,In_38);
xnor U137 (N_137,In_856,In_10);
or U138 (N_138,In_1113,In_658);
nand U139 (N_139,In_1255,In_75);
and U140 (N_140,In_446,In_1178);
and U141 (N_141,In_601,In_1226);
nor U142 (N_142,In_1386,In_1107);
nor U143 (N_143,In_31,In_1366);
nor U144 (N_144,In_1257,In_414);
nand U145 (N_145,In_725,In_182);
xnor U146 (N_146,In_728,In_1246);
nor U147 (N_147,In_1456,In_1496);
and U148 (N_148,In_1201,In_49);
nand U149 (N_149,In_819,In_897);
and U150 (N_150,In_544,In_251);
nand U151 (N_151,In_636,In_499);
and U152 (N_152,In_642,In_1090);
xnor U153 (N_153,In_312,In_1370);
nand U154 (N_154,In_1265,In_313);
or U155 (N_155,In_1013,In_799);
nand U156 (N_156,In_74,In_402);
and U157 (N_157,In_554,In_1045);
nand U158 (N_158,In_825,In_295);
and U159 (N_159,In_120,In_183);
or U160 (N_160,In_793,In_384);
nand U161 (N_161,In_52,In_801);
and U162 (N_162,In_1138,In_46);
nor U163 (N_163,In_230,In_235);
nand U164 (N_164,In_918,In_178);
or U165 (N_165,In_1092,In_398);
and U166 (N_166,In_1403,In_60);
and U167 (N_167,In_967,In_539);
or U168 (N_168,In_772,In_164);
and U169 (N_169,In_912,In_528);
and U170 (N_170,In_471,In_15);
nand U171 (N_171,In_1182,In_660);
nor U172 (N_172,In_203,In_1423);
nor U173 (N_173,In_1413,In_430);
and U174 (N_174,In_1387,In_1314);
or U175 (N_175,In_911,In_439);
nand U176 (N_176,In_1352,In_775);
nor U177 (N_177,In_589,In_1378);
or U178 (N_178,In_452,In_1353);
or U179 (N_179,In_596,In_401);
and U180 (N_180,In_1427,In_1258);
and U181 (N_181,In_139,In_475);
or U182 (N_182,In_1395,In_1315);
nand U183 (N_183,In_480,In_1231);
or U184 (N_184,In_1197,In_1338);
or U185 (N_185,In_778,In_1252);
and U186 (N_186,In_691,In_956);
xnor U187 (N_187,In_192,In_194);
nor U188 (N_188,In_562,In_1063);
nand U189 (N_189,In_745,In_955);
and U190 (N_190,In_1477,In_245);
and U191 (N_191,In_365,In_222);
nor U192 (N_192,In_1458,In_1291);
nand U193 (N_193,In_490,In_160);
nor U194 (N_194,In_1199,In_1470);
nand U195 (N_195,In_434,In_17);
or U196 (N_196,In_1433,In_928);
nor U197 (N_197,In_214,In_512);
nor U198 (N_198,In_659,In_282);
and U199 (N_199,In_1055,In_989);
nand U200 (N_200,In_371,In_1417);
nand U201 (N_201,In_1054,In_1219);
or U202 (N_202,In_522,In_1328);
or U203 (N_203,In_827,In_98);
nor U204 (N_204,In_808,In_784);
and U205 (N_205,In_517,In_1272);
or U206 (N_206,In_1066,In_21);
or U207 (N_207,In_732,In_558);
xor U208 (N_208,In_1230,In_11);
or U209 (N_209,In_635,In_1420);
or U210 (N_210,In_1008,In_71);
and U211 (N_211,In_61,In_907);
and U212 (N_212,In_153,In_638);
nor U213 (N_213,In_947,In_108);
and U214 (N_214,In_564,In_79);
nor U215 (N_215,In_595,In_714);
nor U216 (N_216,In_893,In_682);
nor U217 (N_217,In_1335,In_149);
and U218 (N_218,In_196,In_584);
nand U219 (N_219,In_946,In_829);
and U220 (N_220,In_1158,In_1261);
nand U221 (N_221,In_1437,In_19);
and U222 (N_222,In_1349,In_1012);
nor U223 (N_223,In_25,In_1046);
nand U224 (N_224,In_543,In_656);
xnor U225 (N_225,In_604,In_694);
or U226 (N_226,In_1371,In_1030);
nand U227 (N_227,In_1101,In_926);
nand U228 (N_228,In_249,In_972);
nor U229 (N_229,In_593,In_1466);
or U230 (N_230,In_359,In_6);
nor U231 (N_231,In_455,In_1384);
nand U232 (N_232,In_1244,In_1074);
or U233 (N_233,In_474,In_838);
nand U234 (N_234,In_858,In_1099);
or U235 (N_235,In_1180,In_1485);
and U236 (N_236,In_1147,In_443);
or U237 (N_237,In_1085,In_355);
nand U238 (N_238,In_209,In_8);
and U239 (N_239,In_77,In_1234);
and U240 (N_240,In_252,In_550);
or U241 (N_241,In_698,In_277);
and U242 (N_242,In_89,In_1123);
or U243 (N_243,In_628,In_137);
nor U244 (N_244,In_715,In_72);
nand U245 (N_245,In_679,In_622);
or U246 (N_246,In_1471,In_530);
or U247 (N_247,In_1473,In_1208);
or U248 (N_248,In_332,In_140);
nand U249 (N_249,In_1203,In_822);
and U250 (N_250,In_527,In_1376);
nor U251 (N_251,In_1091,In_1059);
nand U252 (N_252,In_1186,In_1404);
nor U253 (N_253,In_45,In_435);
or U254 (N_254,In_651,In_662);
nor U255 (N_255,In_65,In_389);
nor U256 (N_256,In_696,In_494);
nand U257 (N_257,In_1169,In_950);
xnor U258 (N_258,In_335,In_739);
nand U259 (N_259,In_1102,In_1129);
or U260 (N_260,In_328,In_1118);
and U261 (N_261,In_503,In_1341);
nand U262 (N_262,In_266,In_665);
nand U263 (N_263,In_1462,In_1279);
nor U264 (N_264,In_861,In_1301);
xor U265 (N_265,In_1394,In_12);
nand U266 (N_266,In_1003,In_297);
xor U267 (N_267,In_1297,In_456);
or U268 (N_268,In_1027,In_614);
xnor U269 (N_269,In_1336,In_599);
nor U270 (N_270,In_1011,In_915);
and U271 (N_271,In_1200,In_105);
and U272 (N_272,In_1292,In_1262);
and U273 (N_273,In_1451,In_1356);
and U274 (N_274,In_1294,In_830);
or U275 (N_275,In_1491,In_1428);
and U276 (N_276,In_1082,In_738);
nor U277 (N_277,In_538,In_1414);
and U278 (N_278,In_35,In_555);
nor U279 (N_279,In_531,In_949);
xnor U280 (N_280,In_260,In_1213);
nand U281 (N_281,In_350,In_1039);
nand U282 (N_282,In_647,In_1159);
nand U283 (N_283,In_704,In_796);
or U284 (N_284,In_1347,In_870);
nor U285 (N_285,In_56,In_96);
nand U286 (N_286,In_358,In_1499);
or U287 (N_287,In_1211,In_901);
or U288 (N_288,In_577,In_293);
and U289 (N_289,In_795,In_805);
nor U290 (N_290,In_1259,In_1450);
or U291 (N_291,In_379,In_1195);
nor U292 (N_292,In_1096,In_899);
nand U293 (N_293,In_195,In_1249);
and U294 (N_294,In_1124,In_1320);
and U295 (N_295,In_945,In_217);
or U296 (N_296,In_353,In_661);
xnor U297 (N_297,In_1080,In_300);
or U298 (N_298,In_174,In_921);
nor U299 (N_299,In_469,In_373);
or U300 (N_300,In_134,In_1139);
xor U301 (N_301,In_270,In_168);
or U302 (N_302,In_994,In_1167);
nand U303 (N_303,In_917,In_1327);
or U304 (N_304,In_352,In_591);
or U305 (N_305,In_1461,In_255);
nand U306 (N_306,In_1087,In_1067);
or U307 (N_307,In_892,In_496);
nor U308 (N_308,In_94,In_582);
nand U309 (N_309,In_1094,In_187);
nor U310 (N_310,In_378,In_1454);
and U311 (N_311,In_525,In_1125);
nor U312 (N_312,In_447,In_1325);
xnor U313 (N_313,In_676,In_343);
nor U314 (N_314,In_185,In_145);
nor U315 (N_315,In_800,In_78);
xnor U316 (N_316,In_1287,In_1204);
nand U317 (N_317,In_197,In_687);
xor U318 (N_318,In_476,In_1050);
nand U319 (N_319,In_1269,In_1106);
nor U320 (N_320,In_1495,In_1312);
or U321 (N_321,In_296,In_898);
and U322 (N_322,In_1410,In_833);
or U323 (N_323,In_498,In_1326);
or U324 (N_324,In_2,In_634);
and U325 (N_325,In_1056,In_916);
and U326 (N_326,In_329,In_975);
nand U327 (N_327,In_712,In_1038);
or U328 (N_328,In_684,In_960);
nand U329 (N_329,In_1097,In_1156);
xor U330 (N_330,In_423,In_175);
and U331 (N_331,In_1439,In_485);
or U332 (N_332,In_372,In_1088);
or U333 (N_333,In_1148,In_63);
and U334 (N_334,In_1093,In_567);
nand U335 (N_335,In_1276,In_210);
or U336 (N_336,In_73,In_62);
nor U337 (N_337,In_623,In_42);
and U338 (N_338,In_310,In_1379);
xnor U339 (N_339,In_1264,In_1105);
nor U340 (N_340,In_460,In_242);
nand U341 (N_341,In_316,In_882);
or U342 (N_342,In_1221,In_1133);
and U343 (N_343,In_1014,In_1445);
nor U344 (N_344,In_184,In_637);
or U345 (N_345,In_1408,In_639);
xnor U346 (N_346,In_349,In_247);
nor U347 (N_347,In_448,In_648);
and U348 (N_348,In_763,In_261);
or U349 (N_349,In_1193,In_132);
nand U350 (N_350,In_317,In_991);
and U351 (N_351,In_504,In_1049);
or U352 (N_352,In_717,In_670);
nand U353 (N_353,In_919,In_1432);
or U354 (N_354,In_115,In_767);
xor U355 (N_355,In_570,In_357);
and U356 (N_356,In_723,In_1078);
nand U357 (N_357,In_981,In_1155);
nor U358 (N_358,In_280,In_1188);
nor U359 (N_359,In_399,In_377);
nand U360 (N_360,In_1253,In_133);
xnor U361 (N_361,In_769,In_100);
and U362 (N_362,In_26,In_453);
or U363 (N_363,In_397,In_237);
and U364 (N_364,In_320,In_863);
or U365 (N_365,In_274,In_1281);
xnor U366 (N_366,In_388,In_1271);
xnor U367 (N_367,In_983,In_393);
nand U368 (N_368,In_1263,In_548);
nand U369 (N_369,In_611,In_961);
xnor U370 (N_370,In_1163,In_449);
nand U371 (N_371,In_161,In_1019);
nand U372 (N_372,In_218,In_1498);
nor U373 (N_373,In_536,In_685);
nor U374 (N_374,In_57,In_1134);
nor U375 (N_375,In_1351,In_198);
nor U376 (N_376,In_223,In_1006);
or U377 (N_377,In_905,In_747);
or U378 (N_378,In_1375,In_1072);
xor U379 (N_379,In_716,In_1037);
and U380 (N_380,In_428,In_1126);
or U381 (N_381,In_607,In_1380);
nand U382 (N_382,In_1298,In_869);
nor U383 (N_383,In_566,In_663);
and U384 (N_384,In_1153,In_4);
nand U385 (N_385,In_1415,In_1229);
nor U386 (N_386,In_922,In_29);
or U387 (N_387,In_121,In_495);
nor U388 (N_388,In_1140,In_228);
xnor U389 (N_389,In_586,In_400);
or U390 (N_390,In_1409,In_188);
or U391 (N_391,In_227,In_23);
nor U392 (N_392,In_421,In_920);
nor U393 (N_393,In_839,In_1358);
nand U394 (N_394,In_180,In_1282);
and U395 (N_395,In_618,In_348);
nand U396 (N_396,In_18,In_1112);
and U397 (N_397,In_1296,In_1053);
xor U398 (N_398,In_1024,In_1215);
nor U399 (N_399,In_1194,In_1440);
xor U400 (N_400,In_76,In_1218);
nand U401 (N_401,In_284,In_1368);
nand U402 (N_402,In_997,In_9);
and U403 (N_403,In_1250,In_307);
and U404 (N_404,In_318,In_692);
nand U405 (N_405,In_954,In_816);
nand U406 (N_406,In_1115,In_1483);
nand U407 (N_407,In_557,In_1348);
nand U408 (N_408,In_757,In_3);
xnor U409 (N_409,In_116,In_1273);
nor U410 (N_410,In_523,In_1225);
nor U411 (N_411,In_467,In_986);
or U412 (N_412,In_883,In_1383);
nand U413 (N_413,In_632,In_552);
or U414 (N_414,In_142,In_1493);
and U415 (N_415,In_506,In_1166);
nand U416 (N_416,In_934,In_752);
nand U417 (N_417,In_884,In_1040);
and U418 (N_418,In_1154,In_966);
nor U419 (N_419,In_1185,In_713);
nor U420 (N_420,In_1464,In_820);
and U421 (N_421,In_483,In_1340);
nor U422 (N_422,In_760,In_432);
or U423 (N_423,In_370,In_1494);
nor U424 (N_424,In_1191,In_1365);
or U425 (N_425,In_843,In_1084);
nand U426 (N_426,In_224,In_0);
and U427 (N_427,In_1187,In_1223);
and U428 (N_428,In_254,In_380);
or U429 (N_429,In_276,In_257);
or U430 (N_430,In_734,In_505);
nand U431 (N_431,In_526,In_433);
or U432 (N_432,In_477,In_409);
or U433 (N_433,In_337,In_1350);
nor U434 (N_434,In_289,In_590);
nor U435 (N_435,In_597,In_462);
and U436 (N_436,In_650,In_900);
nand U437 (N_437,In_818,In_292);
nor U438 (N_438,In_718,In_362);
or U439 (N_439,In_1243,In_649);
nor U440 (N_440,In_625,In_1170);
and U441 (N_441,In_700,In_110);
and U442 (N_442,In_1145,In_724);
or U443 (N_443,In_1081,In_95);
nor U444 (N_444,In_964,In_1111);
or U445 (N_445,In_529,In_427);
nor U446 (N_446,In_14,In_47);
xor U447 (N_447,In_1233,In_1236);
and U448 (N_448,In_514,In_761);
and U449 (N_449,In_44,In_190);
nand U450 (N_450,In_678,In_396);
and U451 (N_451,In_109,In_39);
xor U452 (N_452,In_1083,In_220);
and U453 (N_453,In_1141,In_225);
nand U454 (N_454,In_1354,In_319);
and U455 (N_455,In_341,In_1310);
or U456 (N_456,In_1162,In_547);
or U457 (N_457,In_463,In_1399);
and U458 (N_458,In_206,In_420);
nor U459 (N_459,In_944,In_551);
and U460 (N_460,In_693,In_1306);
or U461 (N_461,In_1017,In_613);
nor U462 (N_462,In_931,In_872);
and U463 (N_463,In_37,In_976);
xnor U464 (N_464,In_97,In_1275);
and U465 (N_465,In_338,In_1206);
nor U466 (N_466,In_1209,In_1241);
xor U467 (N_467,In_1028,In_102);
or U468 (N_468,In_1007,In_891);
nor U469 (N_469,In_736,In_1374);
and U470 (N_470,In_1303,In_765);
or U471 (N_471,In_792,In_273);
nor U472 (N_472,In_1150,In_906);
and U473 (N_473,In_1453,In_20);
or U474 (N_474,In_640,In_1482);
nand U475 (N_475,In_1109,In_59);
nor U476 (N_476,In_1041,In_707);
or U477 (N_477,In_1232,In_123);
nor U478 (N_478,In_779,In_112);
xnor U479 (N_479,In_291,In_457);
and U480 (N_480,In_524,In_325);
nor U481 (N_481,In_786,In_202);
and U482 (N_482,In_813,In_1284);
or U483 (N_483,In_1143,In_709);
and U484 (N_484,In_810,In_814);
or U485 (N_485,In_1481,In_737);
nand U486 (N_486,In_1278,In_417);
nand U487 (N_487,In_213,In_619);
and U488 (N_488,In_1469,In_520);
nor U489 (N_489,In_1308,In_626);
nand U490 (N_490,In_83,In_303);
nor U491 (N_491,In_1288,In_269);
nand U492 (N_492,In_68,In_970);
nor U493 (N_493,In_1398,In_67);
or U494 (N_494,In_1405,In_1172);
nor U495 (N_495,In_809,In_492);
nor U496 (N_496,In_126,In_1337);
and U497 (N_497,In_1070,In_1005);
and U498 (N_498,In_272,In_165);
or U499 (N_499,In_546,In_959);
nand U500 (N_500,In_424,In_860);
xor U501 (N_501,In_873,In_581);
and U502 (N_502,In_330,In_438);
nand U503 (N_503,In_472,In_130);
and U504 (N_504,In_501,In_1361);
and U505 (N_505,In_1367,In_620);
or U506 (N_506,In_560,In_1015);
and U507 (N_507,In_782,In_1132);
xor U508 (N_508,In_1189,In_680);
or U509 (N_509,In_629,In_797);
or U510 (N_510,In_88,In_128);
and U511 (N_511,In_1057,In_697);
xnor U512 (N_512,In_200,In_914);
nand U513 (N_513,In_806,In_1235);
nor U514 (N_514,In_146,In_287);
nand U515 (N_515,In_86,In_842);
nand U516 (N_516,In_1490,In_952);
or U517 (N_517,In_1344,In_106);
xnor U518 (N_518,In_340,In_831);
nor U519 (N_519,In_886,In_426);
or U520 (N_520,In_1359,In_510);
xnor U521 (N_521,In_862,In_240);
nand U522 (N_522,In_1489,In_621);
and U523 (N_523,In_848,In_482);
and U524 (N_524,In_1000,In_774);
nor U525 (N_525,In_179,In_1393);
nor U526 (N_526,In_387,In_58);
nor U527 (N_527,In_1307,In_821);
and U528 (N_528,In_1343,In_653);
nor U529 (N_529,In_1174,In_1149);
or U530 (N_530,In_817,In_602);
nand U531 (N_531,In_1486,In_326);
xor U532 (N_532,In_144,In_189);
nor U533 (N_533,In_122,In_1089);
or U534 (N_534,In_729,In_751);
xnor U535 (N_535,In_124,In_755);
nand U536 (N_536,In_933,In_1060);
and U537 (N_537,In_418,In_1086);
and U538 (N_538,In_977,In_444);
nor U539 (N_539,In_537,In_1448);
nand U540 (N_540,In_929,In_777);
nor U541 (N_541,In_327,In_233);
xnor U542 (N_542,In_971,In_978);
nand U543 (N_543,In_103,In_815);
nand U544 (N_544,In_391,In_231);
and U545 (N_545,In_832,In_733);
or U546 (N_546,In_837,In_367);
xnor U547 (N_547,In_1176,In_1114);
or U548 (N_548,In_885,In_114);
nand U549 (N_549,In_1363,In_285);
or U550 (N_550,In_481,In_186);
nor U551 (N_551,In_908,In_731);
or U552 (N_552,In_1022,In_951);
and U553 (N_553,In_167,In_1095);
nor U554 (N_554,In_1245,In_1009);
nand U555 (N_555,In_759,In_941);
and U556 (N_556,In_1311,In_841);
and U557 (N_557,In_93,In_677);
nand U558 (N_558,In_1042,In_854);
nand U559 (N_559,In_1411,In_1382);
xnor U560 (N_560,In_681,In_119);
nor U561 (N_561,In_857,In_721);
nand U562 (N_562,In_1073,In_612);
or U563 (N_563,In_939,In_540);
and U564 (N_564,In_64,In_1324);
nand U565 (N_565,In_1472,In_990);
xnor U566 (N_566,In_113,In_177);
xor U567 (N_567,In_1362,In_768);
or U568 (N_568,In_1492,In_334);
nand U569 (N_569,In_1419,In_152);
and U570 (N_570,In_598,In_1010);
nand U571 (N_571,In_646,In_1429);
nor U572 (N_572,In_868,In_735);
xnor U573 (N_573,In_70,In_383);
nand U574 (N_574,In_1426,In_275);
or U575 (N_575,In_1205,In_641);
nor U576 (N_576,In_896,In_1268);
and U577 (N_577,In_545,In_1479);
or U578 (N_578,In_1421,In_1069);
nand U579 (N_579,In_502,In_394);
and U580 (N_580,In_419,In_436);
or U581 (N_581,In_835,In_608);
nand U582 (N_582,In_1389,In_1210);
nand U583 (N_583,In_34,In_746);
and U584 (N_584,In_1446,In_556);
or U585 (N_585,In_253,In_500);
xor U586 (N_586,In_155,In_118);
and U587 (N_587,In_1316,In_1224);
or U588 (N_588,In_1397,In_1309);
nand U589 (N_589,In_219,In_171);
and U590 (N_590,In_605,In_157);
and U591 (N_591,In_758,In_24);
nand U592 (N_592,In_336,In_299);
nand U593 (N_593,In_1023,In_1302);
or U594 (N_594,In_887,In_654);
or U595 (N_595,In_345,In_1476);
and U596 (N_596,In_583,In_744);
nand U597 (N_597,In_594,In_413);
nand U598 (N_598,In_1016,In_375);
or U599 (N_599,In_703,In_1181);
or U600 (N_600,In_461,In_853);
or U601 (N_601,In_770,In_1025);
or U602 (N_602,In_1434,In_27);
xor U603 (N_603,In_789,In_695);
nand U604 (N_604,In_585,In_1416);
nand U605 (N_605,In_1373,In_410);
nand U606 (N_606,In_286,In_229);
or U607 (N_607,In_50,In_82);
nor U608 (N_608,In_41,In_846);
nor U609 (N_609,In_1043,In_1137);
xnor U610 (N_610,In_559,In_487);
nand U611 (N_611,In_1183,In_465);
nor U612 (N_612,In_753,In_1031);
nand U613 (N_613,In_722,In_412);
xnor U614 (N_614,In_66,In_99);
nor U615 (N_615,In_962,In_1110);
or U616 (N_616,In_172,In_376);
nand U617 (N_617,In_982,In_1270);
and U618 (N_618,In_163,In_422);
and U619 (N_619,In_283,In_1392);
nor U620 (N_620,In_1438,In_279);
or U621 (N_621,In_993,In_234);
and U622 (N_622,In_55,In_600);
nor U623 (N_623,In_1251,In_812);
or U624 (N_624,In_354,In_411);
xnor U625 (N_625,In_479,In_368);
xor U626 (N_626,In_690,In_1372);
or U627 (N_627,In_894,In_624);
or U628 (N_628,In_515,In_855);
and U629 (N_629,In_823,In_1018);
xnor U630 (N_630,In_587,In_743);
xor U631 (N_631,In_553,In_936);
and U632 (N_632,In_1330,In_1);
or U633 (N_633,In_910,In_794);
nor U634 (N_634,In_150,In_323);
nor U635 (N_635,In_1267,In_701);
and U636 (N_636,In_580,In_998);
xor U637 (N_637,In_1152,In_1406);
nor U638 (N_638,In_431,In_573);
nand U639 (N_639,In_346,In_588);
nor U640 (N_640,In_1048,In_969);
or U641 (N_641,In_1052,In_1212);
nand U642 (N_642,In_1120,In_1239);
and U643 (N_643,In_1198,In_781);
or U644 (N_644,In_470,In_710);
and U645 (N_645,In_1076,In_705);
nor U646 (N_646,In_1044,In_925);
and U647 (N_647,In_309,In_429);
and U648 (N_648,In_574,In_923);
and U649 (N_649,In_771,In_927);
nand U650 (N_650,In_1487,In_151);
nor U651 (N_651,In_1228,In_1300);
nand U652 (N_652,In_281,In_1289);
or U653 (N_653,In_1068,In_688);
or U654 (N_654,In_836,In_727);
and U655 (N_655,In_532,In_521);
and U656 (N_656,In_497,In_1157);
xnor U657 (N_657,In_263,In_28);
or U658 (N_658,In_1321,In_754);
xor U659 (N_659,In_16,In_762);
xnor U660 (N_660,In_974,In_271);
or U661 (N_661,In_702,In_1061);
xnor U662 (N_662,In_948,In_306);
or U663 (N_663,In_999,In_1317);
nor U664 (N_664,In_776,In_764);
nand U665 (N_665,In_699,In_569);
or U666 (N_666,In_468,In_1293);
and U667 (N_667,In_489,In_667);
nand U668 (N_668,In_1400,In_507);
nor U669 (N_669,In_1283,In_516);
nand U670 (N_670,In_364,In_1026);
or U671 (N_671,In_30,In_256);
and U672 (N_672,In_803,In_965);
nor U673 (N_673,In_644,In_988);
and U674 (N_674,In_938,In_1488);
or U675 (N_675,In_69,In_963);
or U676 (N_676,In_865,In_879);
or U677 (N_677,In_968,In_91);
nand U678 (N_678,In_80,In_706);
nor U679 (N_679,In_631,In_127);
nor U680 (N_680,In_943,In_1029);
nor U681 (N_681,In_1431,In_645);
nor U682 (N_682,In_1299,In_117);
or U683 (N_683,In_888,In_1071);
and U684 (N_684,In_392,In_301);
or U685 (N_685,In_267,In_828);
nand U686 (N_686,In_1369,In_609);
nand U687 (N_687,In_484,In_579);
nor U688 (N_688,In_565,In_791);
and U689 (N_689,In_314,In_408);
xnor U690 (N_690,In_1319,In_652);
nor U691 (N_691,In_1331,In_1360);
nand U692 (N_692,In_973,In_244);
or U693 (N_693,In_1381,In_51);
nand U694 (N_694,In_1184,In_1222);
or U695 (N_695,In_561,In_87);
nor U696 (N_696,In_1151,In_592);
nand U697 (N_697,In_215,In_459);
nor U698 (N_698,In_199,In_491);
nand U699 (N_699,In_1002,In_1127);
and U700 (N_700,In_1217,In_1179);
xor U701 (N_701,In_850,In_162);
and U702 (N_702,In_107,In_627);
or U703 (N_703,In_278,In_226);
nand U704 (N_704,In_979,In_683);
and U705 (N_705,In_90,In_440);
and U706 (N_706,In_395,In_1214);
or U707 (N_707,In_1216,In_40);
nand U708 (N_708,In_895,In_902);
xor U709 (N_709,In_136,In_1286);
nor U710 (N_710,In_360,In_1346);
nor U711 (N_711,In_193,In_750);
and U712 (N_712,In_1444,In_415);
or U713 (N_713,In_464,In_211);
or U714 (N_714,In_1401,In_54);
and U715 (N_715,In_1130,In_1020);
nor U716 (N_716,In_1165,In_788);
nor U717 (N_717,In_785,In_924);
nor U718 (N_718,In_780,In_347);
or U719 (N_719,In_802,In_509);
or U720 (N_720,In_339,In_81);
nand U721 (N_721,In_643,In_238);
or U722 (N_722,In_290,In_1062);
and U723 (N_723,In_381,In_441);
nor U724 (N_724,In_264,In_356);
or U725 (N_725,In_1305,In_331);
or U726 (N_726,In_425,In_852);
or U727 (N_727,In_1457,In_980);
or U728 (N_728,In_875,In_657);
nor U729 (N_729,In_824,In_549);
xnor U730 (N_730,In_849,In_1285);
xnor U731 (N_731,In_1418,In_568);
nand U732 (N_732,In_675,In_85);
and U733 (N_733,In_111,In_711);
or U734 (N_734,In_265,In_859);
nand U735 (N_735,In_1442,In_259);
nand U736 (N_736,In_876,In_305);
and U737 (N_737,In_847,In_880);
and U738 (N_738,In_442,In_488);
and U739 (N_739,In_909,In_1497);
nand U740 (N_740,In_84,In_606);
or U741 (N_741,In_1436,In_473);
nand U742 (N_742,In_129,In_1449);
nor U743 (N_743,In_1098,In_1441);
nand U744 (N_744,In_333,In_1430);
xor U745 (N_745,In_686,In_874);
and U746 (N_746,In_1396,In_406);
and U747 (N_747,In_840,In_508);
or U748 (N_748,In_221,In_7);
nand U749 (N_749,In_48,In_756);
nor U750 (N_750,In_1448,In_895);
xor U751 (N_751,In_699,In_653);
nor U752 (N_752,In_1319,In_1291);
and U753 (N_753,In_273,In_76);
nand U754 (N_754,In_705,In_281);
nand U755 (N_755,In_1261,In_1402);
nor U756 (N_756,In_140,In_765);
or U757 (N_757,In_783,In_1101);
or U758 (N_758,In_1480,In_1280);
or U759 (N_759,In_1073,In_111);
nor U760 (N_760,In_995,In_988);
or U761 (N_761,In_1258,In_1409);
and U762 (N_762,In_1082,In_906);
xor U763 (N_763,In_862,In_730);
nand U764 (N_764,In_1153,In_967);
nor U765 (N_765,In_1110,In_1094);
nor U766 (N_766,In_943,In_608);
xnor U767 (N_767,In_1473,In_113);
or U768 (N_768,In_1053,In_1331);
and U769 (N_769,In_710,In_610);
nor U770 (N_770,In_876,In_66);
or U771 (N_771,In_1467,In_1495);
nand U772 (N_772,In_626,In_1078);
nand U773 (N_773,In_1130,In_601);
or U774 (N_774,In_1425,In_310);
and U775 (N_775,In_709,In_1213);
nand U776 (N_776,In_1338,In_1476);
and U777 (N_777,In_261,In_1151);
or U778 (N_778,In_1335,In_613);
or U779 (N_779,In_1278,In_787);
nand U780 (N_780,In_1257,In_1094);
nor U781 (N_781,In_1011,In_36);
nor U782 (N_782,In_802,In_173);
nor U783 (N_783,In_732,In_910);
or U784 (N_784,In_1207,In_207);
nand U785 (N_785,In_1490,In_196);
nand U786 (N_786,In_708,In_183);
and U787 (N_787,In_1214,In_630);
and U788 (N_788,In_376,In_466);
and U789 (N_789,In_1186,In_1400);
and U790 (N_790,In_1344,In_726);
nor U791 (N_791,In_493,In_982);
and U792 (N_792,In_1085,In_927);
and U793 (N_793,In_342,In_365);
or U794 (N_794,In_1123,In_85);
and U795 (N_795,In_663,In_474);
or U796 (N_796,In_172,In_333);
or U797 (N_797,In_124,In_1114);
xor U798 (N_798,In_363,In_759);
or U799 (N_799,In_1420,In_948);
or U800 (N_800,In_1088,In_880);
nand U801 (N_801,In_1281,In_332);
nor U802 (N_802,In_1154,In_1160);
nor U803 (N_803,In_1133,In_384);
and U804 (N_804,In_1306,In_1257);
xnor U805 (N_805,In_792,In_387);
nor U806 (N_806,In_211,In_512);
nand U807 (N_807,In_1326,In_934);
or U808 (N_808,In_368,In_116);
nor U809 (N_809,In_1105,In_909);
nor U810 (N_810,In_1368,In_1357);
nand U811 (N_811,In_249,In_1081);
and U812 (N_812,In_1280,In_30);
nand U813 (N_813,In_304,In_1039);
or U814 (N_814,In_528,In_1343);
nand U815 (N_815,In_49,In_563);
nor U816 (N_816,In_918,In_627);
and U817 (N_817,In_1310,In_1022);
nand U818 (N_818,In_357,In_1493);
nor U819 (N_819,In_1173,In_550);
nor U820 (N_820,In_1461,In_407);
and U821 (N_821,In_1212,In_1072);
and U822 (N_822,In_717,In_294);
or U823 (N_823,In_1047,In_1220);
and U824 (N_824,In_52,In_1389);
nand U825 (N_825,In_545,In_387);
or U826 (N_826,In_1038,In_623);
nand U827 (N_827,In_805,In_1198);
nor U828 (N_828,In_124,In_1015);
nor U829 (N_829,In_594,In_1159);
nand U830 (N_830,In_427,In_1104);
and U831 (N_831,In_672,In_133);
nor U832 (N_832,In_432,In_167);
nand U833 (N_833,In_187,In_672);
nand U834 (N_834,In_216,In_668);
nand U835 (N_835,In_566,In_1194);
nand U836 (N_836,In_1125,In_1144);
nand U837 (N_837,In_1475,In_1004);
nor U838 (N_838,In_1083,In_312);
nand U839 (N_839,In_141,In_465);
and U840 (N_840,In_190,In_1033);
and U841 (N_841,In_822,In_430);
and U842 (N_842,In_457,In_1373);
nand U843 (N_843,In_606,In_885);
and U844 (N_844,In_495,In_1294);
or U845 (N_845,In_675,In_127);
and U846 (N_846,In_945,In_960);
and U847 (N_847,In_1373,In_284);
nand U848 (N_848,In_392,In_212);
and U849 (N_849,In_1356,In_1013);
and U850 (N_850,In_1419,In_121);
nor U851 (N_851,In_371,In_384);
and U852 (N_852,In_1003,In_1376);
nor U853 (N_853,In_572,In_321);
xnor U854 (N_854,In_1123,In_311);
nand U855 (N_855,In_1124,In_1244);
nand U856 (N_856,In_36,In_122);
nor U857 (N_857,In_926,In_695);
and U858 (N_858,In_334,In_324);
nor U859 (N_859,In_415,In_913);
nand U860 (N_860,In_1078,In_36);
nor U861 (N_861,In_469,In_739);
or U862 (N_862,In_776,In_173);
or U863 (N_863,In_1001,In_680);
and U864 (N_864,In_1148,In_489);
and U865 (N_865,In_391,In_542);
nand U866 (N_866,In_621,In_223);
xor U867 (N_867,In_134,In_633);
xnor U868 (N_868,In_470,In_646);
and U869 (N_869,In_982,In_112);
nand U870 (N_870,In_445,In_1170);
or U871 (N_871,In_507,In_912);
or U872 (N_872,In_1030,In_777);
and U873 (N_873,In_150,In_106);
nor U874 (N_874,In_1268,In_786);
nand U875 (N_875,In_466,In_1048);
xnor U876 (N_876,In_1086,In_591);
nor U877 (N_877,In_1257,In_95);
and U878 (N_878,In_228,In_639);
nand U879 (N_879,In_655,In_205);
xor U880 (N_880,In_616,In_1215);
and U881 (N_881,In_815,In_1080);
xnor U882 (N_882,In_32,In_1211);
nor U883 (N_883,In_829,In_459);
and U884 (N_884,In_190,In_1130);
xor U885 (N_885,In_704,In_459);
and U886 (N_886,In_668,In_552);
or U887 (N_887,In_1142,In_871);
nand U888 (N_888,In_830,In_1346);
nor U889 (N_889,In_1253,In_457);
or U890 (N_890,In_1353,In_1297);
nand U891 (N_891,In_234,In_842);
or U892 (N_892,In_800,In_323);
and U893 (N_893,In_400,In_959);
and U894 (N_894,In_1380,In_188);
and U895 (N_895,In_723,In_485);
nor U896 (N_896,In_451,In_747);
or U897 (N_897,In_1055,In_1099);
nor U898 (N_898,In_1095,In_1038);
nor U899 (N_899,In_644,In_92);
nor U900 (N_900,In_750,In_245);
and U901 (N_901,In_427,In_1211);
nor U902 (N_902,In_51,In_80);
nand U903 (N_903,In_1307,In_1407);
and U904 (N_904,In_167,In_332);
and U905 (N_905,In_1220,In_642);
and U906 (N_906,In_911,In_1422);
xnor U907 (N_907,In_1412,In_1086);
nand U908 (N_908,In_695,In_351);
and U909 (N_909,In_893,In_1120);
nand U910 (N_910,In_816,In_1149);
nand U911 (N_911,In_652,In_1154);
nor U912 (N_912,In_126,In_1072);
and U913 (N_913,In_218,In_268);
nor U914 (N_914,In_253,In_860);
and U915 (N_915,In_1165,In_1017);
nor U916 (N_916,In_179,In_1382);
nor U917 (N_917,In_739,In_677);
and U918 (N_918,In_998,In_1216);
xor U919 (N_919,In_928,In_1079);
nor U920 (N_920,In_405,In_906);
nand U921 (N_921,In_374,In_1083);
or U922 (N_922,In_1480,In_942);
nand U923 (N_923,In_8,In_1054);
nor U924 (N_924,In_814,In_1226);
nand U925 (N_925,In_218,In_667);
and U926 (N_926,In_1095,In_873);
nand U927 (N_927,In_127,In_714);
xor U928 (N_928,In_682,In_683);
nor U929 (N_929,In_759,In_927);
nor U930 (N_930,In_477,In_545);
nor U931 (N_931,In_420,In_1262);
nand U932 (N_932,In_1114,In_785);
or U933 (N_933,In_753,In_525);
nor U934 (N_934,In_56,In_363);
and U935 (N_935,In_1056,In_888);
and U936 (N_936,In_424,In_1478);
and U937 (N_937,In_1497,In_14);
or U938 (N_938,In_1001,In_1489);
and U939 (N_939,In_187,In_860);
and U940 (N_940,In_652,In_131);
nor U941 (N_941,In_421,In_843);
nand U942 (N_942,In_558,In_872);
or U943 (N_943,In_1100,In_792);
nor U944 (N_944,In_897,In_279);
nand U945 (N_945,In_1252,In_799);
nor U946 (N_946,In_436,In_443);
nor U947 (N_947,In_600,In_1222);
nor U948 (N_948,In_1001,In_259);
nor U949 (N_949,In_1262,In_810);
xnor U950 (N_950,In_305,In_879);
and U951 (N_951,In_495,In_1459);
xor U952 (N_952,In_1428,In_331);
or U953 (N_953,In_41,In_336);
nor U954 (N_954,In_34,In_1465);
and U955 (N_955,In_1394,In_269);
nor U956 (N_956,In_1378,In_742);
or U957 (N_957,In_978,In_770);
or U958 (N_958,In_1060,In_1132);
xor U959 (N_959,In_8,In_1069);
nand U960 (N_960,In_621,In_656);
or U961 (N_961,In_6,In_1490);
and U962 (N_962,In_1452,In_1239);
or U963 (N_963,In_187,In_1437);
or U964 (N_964,In_1241,In_1465);
nand U965 (N_965,In_1225,In_604);
nor U966 (N_966,In_333,In_1177);
and U967 (N_967,In_1388,In_1225);
nand U968 (N_968,In_1452,In_1208);
nor U969 (N_969,In_1367,In_1275);
nor U970 (N_970,In_1306,In_961);
xor U971 (N_971,In_1488,In_173);
and U972 (N_972,In_396,In_443);
and U973 (N_973,In_1259,In_226);
and U974 (N_974,In_350,In_1199);
or U975 (N_975,In_664,In_1199);
nor U976 (N_976,In_1414,In_378);
or U977 (N_977,In_1162,In_383);
nand U978 (N_978,In_1355,In_836);
or U979 (N_979,In_1465,In_1020);
or U980 (N_980,In_456,In_778);
nand U981 (N_981,In_126,In_403);
nand U982 (N_982,In_363,In_1420);
and U983 (N_983,In_162,In_338);
nor U984 (N_984,In_1084,In_1401);
and U985 (N_985,In_1095,In_20);
xnor U986 (N_986,In_0,In_592);
and U987 (N_987,In_638,In_1499);
or U988 (N_988,In_969,In_677);
nor U989 (N_989,In_710,In_352);
xor U990 (N_990,In_41,In_399);
and U991 (N_991,In_351,In_1233);
or U992 (N_992,In_1030,In_1254);
nand U993 (N_993,In_632,In_355);
nand U994 (N_994,In_1238,In_1201);
nor U995 (N_995,In_639,In_415);
and U996 (N_996,In_777,In_941);
and U997 (N_997,In_369,In_1029);
nand U998 (N_998,In_1058,In_1235);
and U999 (N_999,In_835,In_228);
nand U1000 (N_1000,N_604,N_830);
nand U1001 (N_1001,N_399,N_737);
and U1002 (N_1002,N_435,N_122);
nand U1003 (N_1003,N_194,N_350);
nor U1004 (N_1004,N_3,N_902);
xnor U1005 (N_1005,N_425,N_772);
nand U1006 (N_1006,N_33,N_837);
and U1007 (N_1007,N_372,N_219);
or U1008 (N_1008,N_386,N_643);
xor U1009 (N_1009,N_956,N_584);
nor U1010 (N_1010,N_87,N_396);
nand U1011 (N_1011,N_319,N_984);
nor U1012 (N_1012,N_145,N_909);
nand U1013 (N_1013,N_193,N_630);
nor U1014 (N_1014,N_88,N_920);
xnor U1015 (N_1015,N_439,N_79);
or U1016 (N_1016,N_445,N_916);
and U1017 (N_1017,N_656,N_705);
nor U1018 (N_1018,N_817,N_397);
or U1019 (N_1019,N_696,N_436);
and U1020 (N_1020,N_796,N_313);
or U1021 (N_1021,N_881,N_181);
nor U1022 (N_1022,N_317,N_746);
and U1023 (N_1023,N_798,N_934);
or U1024 (N_1024,N_880,N_458);
xnor U1025 (N_1025,N_168,N_167);
or U1026 (N_1026,N_994,N_118);
or U1027 (N_1027,N_421,N_603);
or U1028 (N_1028,N_286,N_676);
and U1029 (N_1029,N_645,N_316);
nor U1030 (N_1030,N_685,N_17);
xnor U1031 (N_1031,N_130,N_366);
or U1032 (N_1032,N_415,N_159);
and U1033 (N_1033,N_708,N_948);
and U1034 (N_1034,N_182,N_358);
nor U1035 (N_1035,N_361,N_7);
and U1036 (N_1036,N_227,N_497);
and U1037 (N_1037,N_689,N_901);
or U1038 (N_1038,N_8,N_155);
nand U1039 (N_1039,N_434,N_897);
and U1040 (N_1040,N_658,N_740);
and U1041 (N_1041,N_276,N_246);
nand U1042 (N_1042,N_250,N_937);
nand U1043 (N_1043,N_736,N_169);
and U1044 (N_1044,N_352,N_154);
nor U1045 (N_1045,N_252,N_983);
or U1046 (N_1046,N_573,N_999);
xnor U1047 (N_1047,N_476,N_259);
and U1048 (N_1048,N_48,N_75);
nand U1049 (N_1049,N_290,N_453);
nand U1050 (N_1050,N_581,N_23);
nor U1051 (N_1051,N_918,N_303);
nor U1052 (N_1052,N_221,N_549);
or U1053 (N_1053,N_185,N_432);
or U1054 (N_1054,N_474,N_892);
nor U1055 (N_1055,N_917,N_776);
nor U1056 (N_1056,N_546,N_300);
nor U1057 (N_1057,N_4,N_534);
or U1058 (N_1058,N_959,N_92);
and U1059 (N_1059,N_975,N_761);
or U1060 (N_1060,N_200,N_30);
nor U1061 (N_1061,N_839,N_512);
nand U1062 (N_1062,N_642,N_707);
or U1063 (N_1063,N_894,N_601);
nand U1064 (N_1064,N_203,N_560);
nand U1065 (N_1065,N_282,N_280);
nor U1066 (N_1066,N_868,N_283);
nor U1067 (N_1067,N_364,N_569);
or U1068 (N_1068,N_813,N_617);
nor U1069 (N_1069,N_623,N_873);
nor U1070 (N_1070,N_940,N_392);
and U1071 (N_1071,N_787,N_405);
nor U1072 (N_1072,N_258,N_624);
xor U1073 (N_1073,N_416,N_359);
or U1074 (N_1074,N_106,N_292);
nand U1075 (N_1075,N_719,N_35);
and U1076 (N_1076,N_733,N_236);
nand U1077 (N_1077,N_235,N_807);
xnor U1078 (N_1078,N_988,N_144);
or U1079 (N_1079,N_655,N_251);
nor U1080 (N_1080,N_793,N_117);
xor U1081 (N_1081,N_137,N_32);
nand U1082 (N_1082,N_472,N_856);
and U1083 (N_1083,N_694,N_9);
nor U1084 (N_1084,N_382,N_874);
nand U1085 (N_1085,N_487,N_634);
and U1086 (N_1086,N_993,N_278);
nand U1087 (N_1087,N_866,N_955);
or U1088 (N_1088,N_102,N_215);
or U1089 (N_1089,N_263,N_844);
nor U1090 (N_1090,N_343,N_321);
xnor U1091 (N_1091,N_893,N_172);
nor U1092 (N_1092,N_522,N_93);
nor U1093 (N_1093,N_70,N_532);
nand U1094 (N_1094,N_490,N_843);
and U1095 (N_1095,N_489,N_401);
nand U1096 (N_1096,N_407,N_121);
nand U1097 (N_1097,N_377,N_500);
or U1098 (N_1098,N_295,N_675);
or U1099 (N_1099,N_845,N_179);
and U1100 (N_1100,N_331,N_550);
nor U1101 (N_1101,N_391,N_759);
nor U1102 (N_1102,N_922,N_139);
xor U1103 (N_1103,N_848,N_61);
and U1104 (N_1104,N_644,N_944);
nand U1105 (N_1105,N_91,N_113);
or U1106 (N_1106,N_34,N_89);
nor U1107 (N_1107,N_29,N_0);
xor U1108 (N_1108,N_621,N_771);
and U1109 (N_1109,N_38,N_367);
xor U1110 (N_1110,N_820,N_677);
or U1111 (N_1111,N_270,N_688);
nor U1112 (N_1112,N_703,N_561);
and U1113 (N_1113,N_20,N_697);
and U1114 (N_1114,N_978,N_556);
or U1115 (N_1115,N_484,N_201);
and U1116 (N_1116,N_333,N_731);
nand U1117 (N_1117,N_790,N_199);
nor U1118 (N_1118,N_562,N_808);
nor U1119 (N_1119,N_724,N_190);
and U1120 (N_1120,N_143,N_509);
nor U1121 (N_1121,N_60,N_39);
or U1122 (N_1122,N_387,N_729);
or U1123 (N_1123,N_234,N_513);
and U1124 (N_1124,N_131,N_570);
or U1125 (N_1125,N_629,N_368);
or U1126 (N_1126,N_46,N_18);
nand U1127 (N_1127,N_175,N_10);
and U1128 (N_1128,N_51,N_402);
or U1129 (N_1129,N_204,N_803);
nor U1130 (N_1130,N_478,N_197);
nor U1131 (N_1131,N_899,N_142);
or U1132 (N_1132,N_721,N_492);
nor U1133 (N_1133,N_557,N_363);
and U1134 (N_1134,N_53,N_441);
nand U1135 (N_1135,N_173,N_637);
or U1136 (N_1136,N_424,N_298);
and U1137 (N_1137,N_751,N_690);
nand U1138 (N_1138,N_68,N_429);
and U1139 (N_1139,N_611,N_58);
and U1140 (N_1140,N_612,N_997);
or U1141 (N_1141,N_277,N_180);
nor U1142 (N_1142,N_886,N_548);
nand U1143 (N_1143,N_198,N_25);
or U1144 (N_1144,N_320,N_247);
or U1145 (N_1145,N_608,N_470);
or U1146 (N_1146,N_946,N_165);
and U1147 (N_1147,N_895,N_791);
nand U1148 (N_1148,N_882,N_646);
or U1149 (N_1149,N_834,N_832);
nor U1150 (N_1150,N_765,N_720);
nor U1151 (N_1151,N_539,N_430);
xor U1152 (N_1152,N_704,N_285);
or U1153 (N_1153,N_481,N_691);
nor U1154 (N_1154,N_462,N_528);
nor U1155 (N_1155,N_157,N_908);
xor U1156 (N_1156,N_96,N_328);
and U1157 (N_1157,N_717,N_241);
nand U1158 (N_1158,N_739,N_592);
or U1159 (N_1159,N_757,N_14);
nor U1160 (N_1160,N_433,N_580);
nor U1161 (N_1161,N_884,N_632);
or U1162 (N_1162,N_887,N_210);
or U1163 (N_1163,N_390,N_888);
nand U1164 (N_1164,N_465,N_495);
nor U1165 (N_1165,N_599,N_176);
or U1166 (N_1166,N_951,N_510);
nor U1167 (N_1167,N_456,N_915);
nand U1168 (N_1168,N_544,N_311);
nand U1169 (N_1169,N_289,N_622);
nand U1170 (N_1170,N_716,N_47);
nand U1171 (N_1171,N_523,N_558);
nor U1172 (N_1172,N_596,N_961);
and U1173 (N_1173,N_755,N_141);
and U1174 (N_1174,N_954,N_28);
nor U1175 (N_1175,N_507,N_602);
nor U1176 (N_1176,N_450,N_340);
and U1177 (N_1177,N_756,N_413);
and U1178 (N_1178,N_861,N_446);
and U1179 (N_1179,N_384,N_448);
xnor U1180 (N_1180,N_239,N_949);
nand U1181 (N_1181,N_52,N_437);
nor U1182 (N_1182,N_62,N_499);
and U1183 (N_1183,N_552,N_981);
nor U1184 (N_1184,N_906,N_305);
nand U1185 (N_1185,N_670,N_55);
nand U1186 (N_1186,N_606,N_875);
or U1187 (N_1187,N_823,N_971);
nor U1188 (N_1188,N_885,N_191);
xnor U1189 (N_1189,N_326,N_864);
nor U1190 (N_1190,N_511,N_45);
or U1191 (N_1191,N_930,N_164);
nor U1192 (N_1192,N_941,N_957);
or U1193 (N_1193,N_105,N_442);
nor U1194 (N_1194,N_712,N_578);
nand U1195 (N_1195,N_403,N_248);
nor U1196 (N_1196,N_799,N_473);
or U1197 (N_1197,N_543,N_393);
or U1198 (N_1198,N_794,N_825);
and U1199 (N_1199,N_620,N_95);
nand U1200 (N_1200,N_222,N_878);
nand U1201 (N_1201,N_78,N_395);
or U1202 (N_1202,N_394,N_341);
or U1203 (N_1203,N_19,N_447);
or U1204 (N_1204,N_564,N_668);
nand U1205 (N_1205,N_809,N_152);
and U1206 (N_1206,N_347,N_572);
nor U1207 (N_1207,N_346,N_695);
and U1208 (N_1208,N_466,N_710);
nand U1209 (N_1209,N_800,N_26);
or U1210 (N_1210,N_650,N_972);
nor U1211 (N_1211,N_388,N_503);
and U1212 (N_1212,N_992,N_715);
xnor U1213 (N_1213,N_400,N_618);
or U1214 (N_1214,N_269,N_980);
nand U1215 (N_1215,N_370,N_281);
nand U1216 (N_1216,N_590,N_15);
or U1217 (N_1217,N_815,N_110);
or U1218 (N_1218,N_336,N_230);
nand U1219 (N_1219,N_711,N_22);
or U1220 (N_1220,N_745,N_936);
nand U1221 (N_1221,N_664,N_898);
or U1222 (N_1222,N_74,N_312);
or U1223 (N_1223,N_174,N_551);
xnor U1224 (N_1224,N_730,N_126);
xnor U1225 (N_1225,N_767,N_267);
or U1226 (N_1226,N_903,N_841);
xor U1227 (N_1227,N_699,N_412);
nor U1228 (N_1228,N_431,N_187);
nor U1229 (N_1229,N_272,N_826);
or U1230 (N_1230,N_207,N_659);
and U1231 (N_1231,N_138,N_802);
nor U1232 (N_1232,N_594,N_789);
nor U1233 (N_1233,N_968,N_297);
nand U1234 (N_1234,N_108,N_50);
nand U1235 (N_1235,N_376,N_764);
or U1236 (N_1236,N_970,N_140);
nand U1237 (N_1237,N_967,N_527);
or U1238 (N_1238,N_455,N_196);
and U1239 (N_1239,N_821,N_208);
nor U1240 (N_1240,N_567,N_274);
nor U1241 (N_1241,N_480,N_666);
or U1242 (N_1242,N_260,N_132);
or U1243 (N_1243,N_64,N_502);
nand U1244 (N_1244,N_762,N_582);
or U1245 (N_1245,N_869,N_890);
or U1246 (N_1246,N_964,N_133);
or U1247 (N_1247,N_750,N_12);
nor U1248 (N_1248,N_850,N_738);
and U1249 (N_1249,N_342,N_995);
nand U1250 (N_1250,N_872,N_498);
xor U1251 (N_1251,N_104,N_942);
nor U1252 (N_1252,N_846,N_408);
and U1253 (N_1253,N_785,N_797);
nor U1254 (N_1254,N_86,N_100);
xnor U1255 (N_1255,N_538,N_440);
or U1256 (N_1256,N_907,N_784);
nand U1257 (N_1257,N_160,N_709);
nor U1258 (N_1258,N_6,N_354);
nor U1259 (N_1259,N_833,N_211);
nor U1260 (N_1260,N_398,N_414);
and U1261 (N_1261,N_647,N_186);
and U1262 (N_1262,N_103,N_979);
and U1263 (N_1263,N_31,N_587);
nand U1264 (N_1264,N_355,N_362);
or U1265 (N_1265,N_693,N_589);
or U1266 (N_1266,N_614,N_56);
and U1267 (N_1267,N_444,N_44);
nor U1268 (N_1268,N_774,N_610);
and U1269 (N_1269,N_452,N_322);
and U1270 (N_1270,N_945,N_849);
xor U1271 (N_1271,N_982,N_518);
nand U1272 (N_1272,N_905,N_149);
and U1273 (N_1273,N_728,N_989);
nor U1274 (N_1274,N_919,N_508);
nor U1275 (N_1275,N_679,N_555);
nor U1276 (N_1276,N_667,N_741);
nand U1277 (N_1277,N_747,N_744);
nand U1278 (N_1278,N_706,N_684);
or U1279 (N_1279,N_521,N_559);
nor U1280 (N_1280,N_279,N_947);
nor U1281 (N_1281,N_883,N_49);
xnor U1282 (N_1282,N_101,N_483);
nor U1283 (N_1283,N_129,N_485);
and U1284 (N_1284,N_324,N_37);
nor U1285 (N_1285,N_847,N_98);
or U1286 (N_1286,N_330,N_170);
nand U1287 (N_1287,N_375,N_344);
nand U1288 (N_1288,N_545,N_921);
nor U1289 (N_1289,N_763,N_422);
nand U1290 (N_1290,N_212,N_43);
or U1291 (N_1291,N_287,N_85);
and U1292 (N_1292,N_127,N_600);
nor U1293 (N_1293,N_753,N_526);
nand U1294 (N_1294,N_163,N_640);
nand U1295 (N_1295,N_966,N_770);
xor U1296 (N_1296,N_648,N_309);
and U1297 (N_1297,N_879,N_304);
and U1298 (N_1298,N_229,N_926);
or U1299 (N_1299,N_912,N_353);
and U1300 (N_1300,N_109,N_795);
nand U1301 (N_1301,N_698,N_209);
nand U1302 (N_1302,N_974,N_952);
nor U1303 (N_1303,N_871,N_77);
nor U1304 (N_1304,N_726,N_649);
nor U1305 (N_1305,N_925,N_59);
nor U1306 (N_1306,N_334,N_619);
xor U1307 (N_1307,N_24,N_124);
xnor U1308 (N_1308,N_520,N_976);
or U1309 (N_1309,N_257,N_13);
nor U1310 (N_1310,N_380,N_579);
or U1311 (N_1311,N_842,N_780);
nor U1312 (N_1312,N_296,N_438);
and U1313 (N_1313,N_27,N_97);
or U1314 (N_1314,N_80,N_428);
nor U1315 (N_1315,N_517,N_566);
and U1316 (N_1316,N_758,N_116);
or U1317 (N_1317,N_238,N_598);
xor U1318 (N_1318,N_914,N_775);
nand U1319 (N_1319,N_778,N_242);
and U1320 (N_1320,N_254,N_877);
nor U1321 (N_1321,N_913,N_865);
or U1322 (N_1322,N_525,N_410);
or U1323 (N_1323,N_781,N_991);
xnor U1324 (N_1324,N_595,N_669);
nand U1325 (N_1325,N_672,N_732);
and U1326 (N_1326,N_963,N_325);
nand U1327 (N_1327,N_651,N_654);
nor U1328 (N_1328,N_423,N_218);
xnor U1329 (N_1329,N_475,N_853);
or U1330 (N_1330,N_404,N_535);
nor U1331 (N_1331,N_529,N_680);
nor U1332 (N_1332,N_256,N_749);
nand U1333 (N_1333,N_674,N_192);
or U1334 (N_1334,N_625,N_563);
and U1335 (N_1335,N_818,N_504);
or U1336 (N_1336,N_686,N_700);
or U1337 (N_1337,N_301,N_125);
and U1338 (N_1338,N_638,N_41);
nand U1339 (N_1339,N_381,N_588);
nand U1340 (N_1340,N_206,N_851);
or U1341 (N_1341,N_858,N_904);
and U1342 (N_1342,N_16,N_687);
xor U1343 (N_1343,N_107,N_216);
and U1344 (N_1344,N_801,N_501);
and U1345 (N_1345,N_760,N_123);
and U1346 (N_1346,N_468,N_530);
xnor U1347 (N_1347,N_547,N_542);
and U1348 (N_1348,N_662,N_863);
or U1349 (N_1349,N_768,N_929);
xnor U1350 (N_1350,N_805,N_65);
and U1351 (N_1351,N_162,N_639);
or U1352 (N_1352,N_299,N_120);
nand U1353 (N_1353,N_253,N_536);
nand U1354 (N_1354,N_838,N_244);
xnor U1355 (N_1355,N_461,N_819);
xor U1356 (N_1356,N_153,N_486);
and U1357 (N_1357,N_420,N_213);
and U1358 (N_1358,N_577,N_943);
nand U1359 (N_1359,N_933,N_824);
xnor U1360 (N_1360,N_339,N_488);
xnor U1361 (N_1361,N_571,N_42);
or U1362 (N_1362,N_240,N_822);
nor U1363 (N_1363,N_810,N_938);
xnor U1364 (N_1364,N_302,N_973);
nor U1365 (N_1365,N_73,N_814);
nor U1366 (N_1366,N_119,N_816);
nand U1367 (N_1367,N_493,N_718);
and U1368 (N_1368,N_953,N_245);
nand U1369 (N_1369,N_482,N_636);
or U1370 (N_1370,N_653,N_965);
or U1371 (N_1371,N_870,N_337);
and U1372 (N_1372,N_626,N_840);
nand U1373 (N_1373,N_852,N_226);
and U1374 (N_1374,N_896,N_683);
nor U1375 (N_1375,N_635,N_958);
nor U1376 (N_1376,N_752,N_2);
nor U1377 (N_1377,N_171,N_67);
and U1378 (N_1378,N_494,N_115);
nand U1379 (N_1379,N_335,N_867);
or U1380 (N_1380,N_479,N_537);
nor U1381 (N_1381,N_161,N_356);
xor U1382 (N_1382,N_345,N_891);
nor U1383 (N_1383,N_417,N_998);
or U1384 (N_1384,N_722,N_275);
or U1385 (N_1385,N_931,N_315);
nand U1386 (N_1386,N_323,N_111);
xnor U1387 (N_1387,N_205,N_63);
nand U1388 (N_1388,N_189,N_950);
nand U1389 (N_1389,N_40,N_188);
or U1390 (N_1390,N_271,N_568);
nor U1391 (N_1391,N_860,N_792);
or U1392 (N_1392,N_713,N_373);
or U1393 (N_1393,N_702,N_379);
or U1394 (N_1394,N_723,N_924);
or U1395 (N_1395,N_288,N_217);
nand U1396 (N_1396,N_927,N_318);
nand U1397 (N_1397,N_613,N_977);
and U1398 (N_1398,N_663,N_294);
xnor U1399 (N_1399,N_349,N_932);
nor U1400 (N_1400,N_609,N_385);
or U1401 (N_1401,N_268,N_962);
and U1402 (N_1402,N_678,N_616);
nor U1403 (N_1403,N_540,N_471);
nor U1404 (N_1404,N_427,N_1);
nand U1405 (N_1405,N_985,N_565);
nand U1406 (N_1406,N_491,N_83);
nand U1407 (N_1407,N_284,N_506);
nor U1408 (N_1408,N_128,N_960);
nor U1409 (N_1409,N_112,N_151);
or U1410 (N_1410,N_516,N_574);
or U1411 (N_1411,N_836,N_255);
or U1412 (N_1412,N_660,N_533);
nand U1413 (N_1413,N_314,N_969);
or U1414 (N_1414,N_69,N_36);
or U1415 (N_1415,N_293,N_348);
and U1416 (N_1416,N_779,N_811);
or U1417 (N_1417,N_214,N_714);
nand U1418 (N_1418,N_990,N_641);
xor U1419 (N_1419,N_519,N_835);
and U1420 (N_1420,N_82,N_859);
and U1421 (N_1421,N_692,N_332);
nor U1422 (N_1422,N_682,N_773);
nor U1423 (N_1423,N_627,N_734);
nand U1424 (N_1424,N_135,N_607);
nor U1425 (N_1425,N_505,N_464);
nor U1426 (N_1426,N_575,N_114);
and U1427 (N_1427,N_806,N_876);
nand U1428 (N_1428,N_5,N_329);
xnor U1429 (N_1429,N_409,N_671);
nor U1430 (N_1430,N_597,N_804);
and U1431 (N_1431,N_986,N_419);
nor U1432 (N_1432,N_769,N_457);
nor U1433 (N_1433,N_76,N_195);
and U1434 (N_1434,N_360,N_21);
nor U1435 (N_1435,N_743,N_725);
and U1436 (N_1436,N_310,N_665);
nor U1437 (N_1437,N_177,N_54);
nand U1438 (N_1438,N_224,N_593);
nand U1439 (N_1439,N_443,N_291);
nor U1440 (N_1440,N_66,N_265);
nand U1441 (N_1441,N_829,N_146);
and U1442 (N_1442,N_911,N_266);
or U1443 (N_1443,N_84,N_262);
and U1444 (N_1444,N_812,N_661);
and U1445 (N_1445,N_754,N_515);
nand U1446 (N_1446,N_553,N_351);
and U1447 (N_1447,N_166,N_338);
and U1448 (N_1448,N_460,N_243);
nor U1449 (N_1449,N_273,N_615);
nor U1450 (N_1450,N_220,N_233);
nor U1451 (N_1451,N_628,N_786);
and U1452 (N_1452,N_459,N_910);
or U1453 (N_1453,N_585,N_147);
nor U1454 (N_1454,N_463,N_81);
nand U1455 (N_1455,N_406,N_148);
or U1456 (N_1456,N_857,N_369);
xor U1457 (N_1457,N_374,N_928);
and U1458 (N_1458,N_855,N_449);
nor U1459 (N_1459,N_454,N_389);
or U1460 (N_1460,N_923,N_605);
and U1461 (N_1461,N_514,N_554);
or U1462 (N_1462,N_378,N_652);
nand U1463 (N_1463,N_223,N_94);
and U1464 (N_1464,N_633,N_742);
and U1465 (N_1465,N_72,N_996);
or U1466 (N_1466,N_156,N_854);
nor U1467 (N_1467,N_183,N_935);
and U1468 (N_1468,N_184,N_327);
nor U1469 (N_1469,N_426,N_71);
nor U1470 (N_1470,N_777,N_237);
and U1471 (N_1471,N_631,N_782);
xor U1472 (N_1472,N_889,N_496);
nor U1473 (N_1473,N_231,N_225);
or U1474 (N_1474,N_586,N_99);
nor U1475 (N_1475,N_158,N_727);
nor U1476 (N_1476,N_307,N_576);
or U1477 (N_1477,N_228,N_987);
and U1478 (N_1478,N_900,N_591);
nand U1479 (N_1479,N_583,N_150);
nor U1480 (N_1480,N_365,N_57);
and U1481 (N_1481,N_264,N_783);
or U1482 (N_1482,N_90,N_657);
nor U1483 (N_1483,N_788,N_673);
nor U1484 (N_1484,N_467,N_202);
nor U1485 (N_1485,N_828,N_232);
and U1486 (N_1486,N_306,N_531);
and U1487 (N_1487,N_178,N_451);
nand U1488 (N_1488,N_411,N_418);
nand U1489 (N_1489,N_357,N_524);
nand U1490 (N_1490,N_134,N_308);
and U1491 (N_1491,N_701,N_261);
nor U1492 (N_1492,N_681,N_371);
nand U1493 (N_1493,N_469,N_541);
and U1494 (N_1494,N_735,N_831);
nand U1495 (N_1495,N_939,N_748);
nor U1496 (N_1496,N_477,N_136);
or U1497 (N_1497,N_11,N_249);
and U1498 (N_1498,N_766,N_383);
nand U1499 (N_1499,N_827,N_862);
nand U1500 (N_1500,N_226,N_186);
nand U1501 (N_1501,N_963,N_272);
and U1502 (N_1502,N_714,N_597);
xor U1503 (N_1503,N_584,N_302);
nor U1504 (N_1504,N_210,N_763);
nand U1505 (N_1505,N_115,N_445);
nor U1506 (N_1506,N_645,N_723);
and U1507 (N_1507,N_640,N_900);
nand U1508 (N_1508,N_633,N_381);
nor U1509 (N_1509,N_872,N_496);
and U1510 (N_1510,N_203,N_19);
nand U1511 (N_1511,N_927,N_132);
nor U1512 (N_1512,N_659,N_919);
nand U1513 (N_1513,N_284,N_815);
nor U1514 (N_1514,N_294,N_587);
nand U1515 (N_1515,N_478,N_982);
nand U1516 (N_1516,N_914,N_261);
nand U1517 (N_1517,N_340,N_76);
and U1518 (N_1518,N_444,N_593);
nand U1519 (N_1519,N_110,N_995);
and U1520 (N_1520,N_583,N_126);
nor U1521 (N_1521,N_50,N_658);
or U1522 (N_1522,N_888,N_432);
nor U1523 (N_1523,N_691,N_564);
nor U1524 (N_1524,N_317,N_160);
and U1525 (N_1525,N_839,N_190);
and U1526 (N_1526,N_382,N_988);
nor U1527 (N_1527,N_442,N_291);
nand U1528 (N_1528,N_286,N_609);
xor U1529 (N_1529,N_673,N_865);
nand U1530 (N_1530,N_450,N_994);
and U1531 (N_1531,N_203,N_226);
nor U1532 (N_1532,N_478,N_248);
nand U1533 (N_1533,N_794,N_258);
nor U1534 (N_1534,N_947,N_211);
nor U1535 (N_1535,N_62,N_771);
and U1536 (N_1536,N_141,N_702);
nor U1537 (N_1537,N_98,N_197);
nand U1538 (N_1538,N_804,N_838);
nand U1539 (N_1539,N_183,N_247);
and U1540 (N_1540,N_926,N_312);
nor U1541 (N_1541,N_549,N_445);
xnor U1542 (N_1542,N_771,N_156);
nor U1543 (N_1543,N_777,N_599);
or U1544 (N_1544,N_14,N_52);
or U1545 (N_1545,N_532,N_33);
or U1546 (N_1546,N_310,N_463);
and U1547 (N_1547,N_254,N_154);
or U1548 (N_1548,N_271,N_316);
or U1549 (N_1549,N_578,N_564);
nor U1550 (N_1550,N_458,N_160);
or U1551 (N_1551,N_650,N_37);
nand U1552 (N_1552,N_553,N_239);
xnor U1553 (N_1553,N_330,N_451);
nand U1554 (N_1554,N_167,N_302);
or U1555 (N_1555,N_839,N_472);
nor U1556 (N_1556,N_304,N_647);
or U1557 (N_1557,N_6,N_981);
nand U1558 (N_1558,N_578,N_869);
nand U1559 (N_1559,N_362,N_584);
nor U1560 (N_1560,N_594,N_113);
nor U1561 (N_1561,N_567,N_974);
xnor U1562 (N_1562,N_978,N_743);
nor U1563 (N_1563,N_125,N_849);
nor U1564 (N_1564,N_834,N_839);
or U1565 (N_1565,N_998,N_187);
and U1566 (N_1566,N_457,N_52);
or U1567 (N_1567,N_768,N_144);
nor U1568 (N_1568,N_167,N_541);
and U1569 (N_1569,N_349,N_936);
or U1570 (N_1570,N_940,N_629);
nand U1571 (N_1571,N_581,N_976);
and U1572 (N_1572,N_431,N_390);
and U1573 (N_1573,N_339,N_491);
nand U1574 (N_1574,N_715,N_49);
or U1575 (N_1575,N_103,N_357);
nor U1576 (N_1576,N_671,N_465);
or U1577 (N_1577,N_89,N_733);
nand U1578 (N_1578,N_245,N_384);
or U1579 (N_1579,N_397,N_346);
and U1580 (N_1580,N_252,N_328);
or U1581 (N_1581,N_906,N_627);
and U1582 (N_1582,N_560,N_691);
nand U1583 (N_1583,N_924,N_157);
and U1584 (N_1584,N_340,N_0);
or U1585 (N_1585,N_160,N_176);
nor U1586 (N_1586,N_936,N_486);
or U1587 (N_1587,N_467,N_634);
and U1588 (N_1588,N_770,N_357);
nand U1589 (N_1589,N_663,N_336);
nand U1590 (N_1590,N_690,N_194);
or U1591 (N_1591,N_86,N_10);
or U1592 (N_1592,N_39,N_422);
nor U1593 (N_1593,N_183,N_918);
and U1594 (N_1594,N_367,N_175);
and U1595 (N_1595,N_932,N_619);
and U1596 (N_1596,N_486,N_878);
nor U1597 (N_1597,N_804,N_532);
or U1598 (N_1598,N_645,N_225);
nor U1599 (N_1599,N_503,N_416);
and U1600 (N_1600,N_847,N_668);
and U1601 (N_1601,N_462,N_938);
or U1602 (N_1602,N_926,N_84);
nor U1603 (N_1603,N_307,N_148);
nand U1604 (N_1604,N_733,N_258);
nor U1605 (N_1605,N_177,N_649);
or U1606 (N_1606,N_736,N_293);
and U1607 (N_1607,N_693,N_32);
nor U1608 (N_1608,N_685,N_807);
nand U1609 (N_1609,N_708,N_924);
xor U1610 (N_1610,N_183,N_869);
and U1611 (N_1611,N_97,N_748);
nand U1612 (N_1612,N_477,N_155);
nand U1613 (N_1613,N_458,N_598);
xor U1614 (N_1614,N_976,N_287);
or U1615 (N_1615,N_434,N_618);
nor U1616 (N_1616,N_497,N_995);
and U1617 (N_1617,N_592,N_528);
nor U1618 (N_1618,N_383,N_976);
and U1619 (N_1619,N_735,N_969);
or U1620 (N_1620,N_46,N_709);
and U1621 (N_1621,N_397,N_197);
nand U1622 (N_1622,N_526,N_325);
nor U1623 (N_1623,N_425,N_120);
nor U1624 (N_1624,N_235,N_851);
and U1625 (N_1625,N_309,N_68);
or U1626 (N_1626,N_394,N_526);
or U1627 (N_1627,N_129,N_513);
and U1628 (N_1628,N_888,N_114);
or U1629 (N_1629,N_147,N_592);
and U1630 (N_1630,N_778,N_894);
nand U1631 (N_1631,N_327,N_599);
and U1632 (N_1632,N_820,N_597);
and U1633 (N_1633,N_860,N_830);
and U1634 (N_1634,N_512,N_318);
nor U1635 (N_1635,N_657,N_673);
nor U1636 (N_1636,N_735,N_51);
nor U1637 (N_1637,N_836,N_778);
or U1638 (N_1638,N_757,N_119);
nor U1639 (N_1639,N_868,N_622);
or U1640 (N_1640,N_788,N_656);
and U1641 (N_1641,N_142,N_674);
nor U1642 (N_1642,N_299,N_336);
or U1643 (N_1643,N_865,N_578);
nand U1644 (N_1644,N_475,N_720);
or U1645 (N_1645,N_947,N_751);
or U1646 (N_1646,N_645,N_321);
xor U1647 (N_1647,N_916,N_830);
nand U1648 (N_1648,N_596,N_936);
xnor U1649 (N_1649,N_519,N_147);
nor U1650 (N_1650,N_652,N_113);
and U1651 (N_1651,N_89,N_229);
or U1652 (N_1652,N_658,N_952);
nor U1653 (N_1653,N_220,N_428);
and U1654 (N_1654,N_985,N_505);
nand U1655 (N_1655,N_516,N_570);
nand U1656 (N_1656,N_924,N_604);
xnor U1657 (N_1657,N_894,N_335);
and U1658 (N_1658,N_174,N_539);
or U1659 (N_1659,N_439,N_126);
nand U1660 (N_1660,N_435,N_116);
and U1661 (N_1661,N_413,N_90);
or U1662 (N_1662,N_665,N_244);
xnor U1663 (N_1663,N_51,N_192);
nand U1664 (N_1664,N_652,N_871);
nor U1665 (N_1665,N_810,N_851);
or U1666 (N_1666,N_761,N_89);
and U1667 (N_1667,N_303,N_515);
nand U1668 (N_1668,N_7,N_339);
or U1669 (N_1669,N_588,N_127);
xnor U1670 (N_1670,N_508,N_714);
or U1671 (N_1671,N_965,N_996);
nand U1672 (N_1672,N_129,N_478);
or U1673 (N_1673,N_26,N_535);
nand U1674 (N_1674,N_382,N_464);
or U1675 (N_1675,N_914,N_457);
nor U1676 (N_1676,N_121,N_375);
and U1677 (N_1677,N_78,N_948);
nor U1678 (N_1678,N_752,N_481);
nand U1679 (N_1679,N_679,N_394);
or U1680 (N_1680,N_21,N_898);
xor U1681 (N_1681,N_824,N_280);
and U1682 (N_1682,N_796,N_333);
xnor U1683 (N_1683,N_468,N_867);
or U1684 (N_1684,N_34,N_261);
and U1685 (N_1685,N_621,N_233);
or U1686 (N_1686,N_621,N_828);
or U1687 (N_1687,N_784,N_36);
or U1688 (N_1688,N_701,N_840);
xor U1689 (N_1689,N_85,N_551);
nand U1690 (N_1690,N_630,N_58);
and U1691 (N_1691,N_488,N_318);
nand U1692 (N_1692,N_827,N_436);
nand U1693 (N_1693,N_684,N_711);
and U1694 (N_1694,N_487,N_528);
xor U1695 (N_1695,N_644,N_351);
nor U1696 (N_1696,N_100,N_77);
or U1697 (N_1697,N_499,N_667);
nor U1698 (N_1698,N_531,N_825);
nor U1699 (N_1699,N_479,N_122);
and U1700 (N_1700,N_975,N_600);
or U1701 (N_1701,N_692,N_456);
and U1702 (N_1702,N_933,N_499);
and U1703 (N_1703,N_639,N_656);
and U1704 (N_1704,N_130,N_873);
and U1705 (N_1705,N_51,N_932);
nor U1706 (N_1706,N_600,N_589);
or U1707 (N_1707,N_24,N_137);
or U1708 (N_1708,N_613,N_907);
and U1709 (N_1709,N_279,N_396);
or U1710 (N_1710,N_41,N_565);
nor U1711 (N_1711,N_906,N_296);
nand U1712 (N_1712,N_963,N_105);
or U1713 (N_1713,N_606,N_705);
nand U1714 (N_1714,N_827,N_893);
nor U1715 (N_1715,N_627,N_7);
and U1716 (N_1716,N_266,N_508);
xor U1717 (N_1717,N_2,N_149);
or U1718 (N_1718,N_726,N_33);
nor U1719 (N_1719,N_100,N_292);
nor U1720 (N_1720,N_670,N_699);
nor U1721 (N_1721,N_454,N_102);
nor U1722 (N_1722,N_453,N_331);
nor U1723 (N_1723,N_983,N_147);
or U1724 (N_1724,N_296,N_966);
and U1725 (N_1725,N_230,N_755);
nor U1726 (N_1726,N_725,N_726);
nand U1727 (N_1727,N_929,N_844);
nor U1728 (N_1728,N_446,N_284);
nand U1729 (N_1729,N_321,N_78);
or U1730 (N_1730,N_19,N_386);
and U1731 (N_1731,N_283,N_630);
and U1732 (N_1732,N_609,N_6);
nand U1733 (N_1733,N_578,N_341);
and U1734 (N_1734,N_198,N_528);
or U1735 (N_1735,N_747,N_48);
or U1736 (N_1736,N_685,N_238);
nand U1737 (N_1737,N_998,N_327);
or U1738 (N_1738,N_403,N_38);
and U1739 (N_1739,N_60,N_246);
nand U1740 (N_1740,N_859,N_87);
nor U1741 (N_1741,N_596,N_763);
nand U1742 (N_1742,N_695,N_60);
nand U1743 (N_1743,N_703,N_37);
or U1744 (N_1744,N_972,N_800);
nand U1745 (N_1745,N_413,N_867);
nand U1746 (N_1746,N_824,N_481);
nand U1747 (N_1747,N_905,N_240);
nand U1748 (N_1748,N_317,N_383);
and U1749 (N_1749,N_691,N_303);
or U1750 (N_1750,N_953,N_707);
nand U1751 (N_1751,N_897,N_327);
and U1752 (N_1752,N_289,N_768);
nand U1753 (N_1753,N_733,N_382);
nor U1754 (N_1754,N_422,N_183);
nor U1755 (N_1755,N_195,N_379);
and U1756 (N_1756,N_590,N_503);
xnor U1757 (N_1757,N_125,N_650);
and U1758 (N_1758,N_784,N_841);
or U1759 (N_1759,N_850,N_820);
and U1760 (N_1760,N_931,N_163);
nor U1761 (N_1761,N_864,N_447);
nand U1762 (N_1762,N_302,N_119);
or U1763 (N_1763,N_11,N_690);
xnor U1764 (N_1764,N_547,N_688);
nor U1765 (N_1765,N_969,N_931);
nand U1766 (N_1766,N_494,N_328);
or U1767 (N_1767,N_126,N_632);
and U1768 (N_1768,N_901,N_277);
nor U1769 (N_1769,N_64,N_595);
and U1770 (N_1770,N_320,N_862);
nor U1771 (N_1771,N_317,N_423);
xnor U1772 (N_1772,N_149,N_107);
or U1773 (N_1773,N_571,N_737);
or U1774 (N_1774,N_532,N_681);
or U1775 (N_1775,N_645,N_249);
nand U1776 (N_1776,N_900,N_108);
and U1777 (N_1777,N_937,N_394);
and U1778 (N_1778,N_336,N_809);
nand U1779 (N_1779,N_770,N_874);
and U1780 (N_1780,N_544,N_272);
nor U1781 (N_1781,N_437,N_770);
or U1782 (N_1782,N_806,N_862);
or U1783 (N_1783,N_275,N_80);
and U1784 (N_1784,N_144,N_984);
or U1785 (N_1785,N_441,N_927);
and U1786 (N_1786,N_677,N_62);
and U1787 (N_1787,N_701,N_466);
and U1788 (N_1788,N_962,N_282);
nor U1789 (N_1789,N_268,N_267);
nand U1790 (N_1790,N_157,N_611);
and U1791 (N_1791,N_1,N_628);
or U1792 (N_1792,N_387,N_918);
nor U1793 (N_1793,N_856,N_705);
and U1794 (N_1794,N_478,N_225);
nor U1795 (N_1795,N_430,N_582);
xor U1796 (N_1796,N_75,N_643);
and U1797 (N_1797,N_132,N_705);
or U1798 (N_1798,N_16,N_166);
nor U1799 (N_1799,N_263,N_313);
nand U1800 (N_1800,N_532,N_510);
nand U1801 (N_1801,N_165,N_236);
nand U1802 (N_1802,N_898,N_10);
xor U1803 (N_1803,N_37,N_367);
and U1804 (N_1804,N_697,N_400);
nand U1805 (N_1805,N_285,N_921);
or U1806 (N_1806,N_718,N_190);
nor U1807 (N_1807,N_120,N_716);
or U1808 (N_1808,N_865,N_501);
nand U1809 (N_1809,N_720,N_402);
and U1810 (N_1810,N_190,N_859);
and U1811 (N_1811,N_569,N_47);
nor U1812 (N_1812,N_153,N_370);
or U1813 (N_1813,N_778,N_83);
xor U1814 (N_1814,N_630,N_772);
nor U1815 (N_1815,N_603,N_905);
and U1816 (N_1816,N_449,N_480);
nor U1817 (N_1817,N_883,N_138);
or U1818 (N_1818,N_878,N_594);
nand U1819 (N_1819,N_58,N_300);
or U1820 (N_1820,N_881,N_845);
and U1821 (N_1821,N_361,N_654);
and U1822 (N_1822,N_985,N_369);
or U1823 (N_1823,N_158,N_498);
and U1824 (N_1824,N_701,N_599);
or U1825 (N_1825,N_20,N_253);
nor U1826 (N_1826,N_535,N_794);
and U1827 (N_1827,N_540,N_563);
or U1828 (N_1828,N_118,N_572);
nand U1829 (N_1829,N_623,N_222);
nor U1830 (N_1830,N_530,N_443);
and U1831 (N_1831,N_78,N_618);
nor U1832 (N_1832,N_781,N_876);
and U1833 (N_1833,N_452,N_485);
or U1834 (N_1834,N_636,N_192);
and U1835 (N_1835,N_528,N_172);
or U1836 (N_1836,N_587,N_506);
xnor U1837 (N_1837,N_987,N_325);
nand U1838 (N_1838,N_218,N_606);
and U1839 (N_1839,N_851,N_554);
nand U1840 (N_1840,N_535,N_610);
nor U1841 (N_1841,N_54,N_972);
nand U1842 (N_1842,N_454,N_861);
or U1843 (N_1843,N_663,N_919);
nor U1844 (N_1844,N_566,N_551);
and U1845 (N_1845,N_909,N_411);
and U1846 (N_1846,N_544,N_674);
nor U1847 (N_1847,N_865,N_927);
nand U1848 (N_1848,N_130,N_62);
nor U1849 (N_1849,N_79,N_590);
and U1850 (N_1850,N_410,N_88);
nor U1851 (N_1851,N_768,N_76);
xor U1852 (N_1852,N_394,N_407);
nand U1853 (N_1853,N_790,N_811);
and U1854 (N_1854,N_931,N_471);
and U1855 (N_1855,N_280,N_412);
or U1856 (N_1856,N_308,N_317);
nor U1857 (N_1857,N_691,N_835);
or U1858 (N_1858,N_22,N_252);
or U1859 (N_1859,N_833,N_473);
nor U1860 (N_1860,N_735,N_276);
nand U1861 (N_1861,N_960,N_882);
nand U1862 (N_1862,N_691,N_810);
or U1863 (N_1863,N_152,N_199);
or U1864 (N_1864,N_424,N_276);
nand U1865 (N_1865,N_575,N_617);
or U1866 (N_1866,N_918,N_173);
nand U1867 (N_1867,N_937,N_731);
nand U1868 (N_1868,N_470,N_524);
nand U1869 (N_1869,N_50,N_286);
and U1870 (N_1870,N_836,N_828);
and U1871 (N_1871,N_280,N_257);
nor U1872 (N_1872,N_847,N_397);
nand U1873 (N_1873,N_102,N_295);
nand U1874 (N_1874,N_293,N_221);
nand U1875 (N_1875,N_103,N_855);
and U1876 (N_1876,N_952,N_290);
nor U1877 (N_1877,N_550,N_926);
nor U1878 (N_1878,N_547,N_824);
nor U1879 (N_1879,N_328,N_189);
nand U1880 (N_1880,N_41,N_883);
nor U1881 (N_1881,N_273,N_807);
and U1882 (N_1882,N_627,N_492);
or U1883 (N_1883,N_323,N_449);
or U1884 (N_1884,N_91,N_707);
or U1885 (N_1885,N_41,N_486);
or U1886 (N_1886,N_593,N_352);
nor U1887 (N_1887,N_706,N_766);
xnor U1888 (N_1888,N_34,N_579);
or U1889 (N_1889,N_761,N_755);
nor U1890 (N_1890,N_397,N_60);
nor U1891 (N_1891,N_510,N_243);
nor U1892 (N_1892,N_988,N_881);
nor U1893 (N_1893,N_174,N_275);
nor U1894 (N_1894,N_70,N_881);
and U1895 (N_1895,N_254,N_319);
or U1896 (N_1896,N_465,N_905);
or U1897 (N_1897,N_952,N_665);
and U1898 (N_1898,N_934,N_547);
and U1899 (N_1899,N_364,N_867);
and U1900 (N_1900,N_339,N_320);
nor U1901 (N_1901,N_581,N_335);
nand U1902 (N_1902,N_542,N_496);
nand U1903 (N_1903,N_423,N_646);
nor U1904 (N_1904,N_770,N_79);
or U1905 (N_1905,N_474,N_273);
nor U1906 (N_1906,N_357,N_620);
and U1907 (N_1907,N_562,N_135);
xnor U1908 (N_1908,N_588,N_546);
xor U1909 (N_1909,N_577,N_281);
nor U1910 (N_1910,N_477,N_475);
or U1911 (N_1911,N_145,N_295);
nand U1912 (N_1912,N_947,N_734);
or U1913 (N_1913,N_801,N_252);
or U1914 (N_1914,N_610,N_256);
nand U1915 (N_1915,N_636,N_169);
and U1916 (N_1916,N_147,N_245);
or U1917 (N_1917,N_272,N_297);
and U1918 (N_1918,N_498,N_155);
or U1919 (N_1919,N_135,N_246);
xnor U1920 (N_1920,N_45,N_778);
nor U1921 (N_1921,N_443,N_518);
or U1922 (N_1922,N_747,N_455);
and U1923 (N_1923,N_543,N_485);
nand U1924 (N_1924,N_430,N_800);
nor U1925 (N_1925,N_811,N_652);
or U1926 (N_1926,N_946,N_485);
and U1927 (N_1927,N_911,N_54);
and U1928 (N_1928,N_577,N_696);
or U1929 (N_1929,N_671,N_8);
nor U1930 (N_1930,N_242,N_808);
xnor U1931 (N_1931,N_503,N_676);
and U1932 (N_1932,N_541,N_670);
and U1933 (N_1933,N_543,N_835);
nor U1934 (N_1934,N_303,N_67);
and U1935 (N_1935,N_498,N_873);
and U1936 (N_1936,N_369,N_544);
nor U1937 (N_1937,N_652,N_464);
and U1938 (N_1938,N_704,N_34);
nand U1939 (N_1939,N_724,N_236);
nor U1940 (N_1940,N_435,N_166);
and U1941 (N_1941,N_998,N_167);
nor U1942 (N_1942,N_94,N_849);
nand U1943 (N_1943,N_486,N_140);
nor U1944 (N_1944,N_616,N_574);
nor U1945 (N_1945,N_322,N_881);
and U1946 (N_1946,N_918,N_518);
nor U1947 (N_1947,N_302,N_601);
nand U1948 (N_1948,N_590,N_871);
xor U1949 (N_1949,N_647,N_923);
nand U1950 (N_1950,N_463,N_991);
and U1951 (N_1951,N_819,N_334);
and U1952 (N_1952,N_880,N_57);
and U1953 (N_1953,N_12,N_65);
or U1954 (N_1954,N_743,N_762);
nor U1955 (N_1955,N_642,N_190);
nand U1956 (N_1956,N_215,N_239);
or U1957 (N_1957,N_237,N_683);
and U1958 (N_1958,N_775,N_673);
nor U1959 (N_1959,N_851,N_734);
and U1960 (N_1960,N_100,N_96);
and U1961 (N_1961,N_938,N_638);
nand U1962 (N_1962,N_422,N_518);
nor U1963 (N_1963,N_73,N_938);
nand U1964 (N_1964,N_583,N_236);
nand U1965 (N_1965,N_242,N_328);
and U1966 (N_1966,N_350,N_822);
or U1967 (N_1967,N_96,N_930);
or U1968 (N_1968,N_244,N_126);
or U1969 (N_1969,N_227,N_456);
nand U1970 (N_1970,N_676,N_218);
and U1971 (N_1971,N_853,N_354);
nor U1972 (N_1972,N_160,N_346);
nor U1973 (N_1973,N_853,N_296);
nand U1974 (N_1974,N_57,N_556);
or U1975 (N_1975,N_849,N_794);
nand U1976 (N_1976,N_678,N_863);
xnor U1977 (N_1977,N_436,N_274);
or U1978 (N_1978,N_409,N_429);
or U1979 (N_1979,N_759,N_957);
nand U1980 (N_1980,N_78,N_370);
xnor U1981 (N_1981,N_62,N_271);
or U1982 (N_1982,N_530,N_556);
or U1983 (N_1983,N_139,N_547);
and U1984 (N_1984,N_511,N_180);
or U1985 (N_1985,N_735,N_446);
nand U1986 (N_1986,N_357,N_592);
xnor U1987 (N_1987,N_89,N_199);
nand U1988 (N_1988,N_231,N_639);
and U1989 (N_1989,N_198,N_956);
nor U1990 (N_1990,N_660,N_753);
and U1991 (N_1991,N_98,N_89);
nor U1992 (N_1992,N_251,N_321);
nand U1993 (N_1993,N_791,N_258);
nand U1994 (N_1994,N_474,N_25);
nand U1995 (N_1995,N_152,N_253);
and U1996 (N_1996,N_516,N_244);
xor U1997 (N_1997,N_877,N_242);
nor U1998 (N_1998,N_885,N_336);
and U1999 (N_1999,N_822,N_410);
and U2000 (N_2000,N_1962,N_1731);
xnor U2001 (N_2001,N_1887,N_1653);
and U2002 (N_2002,N_1659,N_1335);
and U2003 (N_2003,N_1904,N_1798);
nand U2004 (N_2004,N_1632,N_1138);
and U2005 (N_2005,N_1586,N_1840);
and U2006 (N_2006,N_1427,N_1555);
and U2007 (N_2007,N_1537,N_1194);
nor U2008 (N_2008,N_1108,N_1684);
nand U2009 (N_2009,N_1815,N_1738);
and U2010 (N_2010,N_1508,N_1912);
nand U2011 (N_2011,N_1472,N_1379);
and U2012 (N_2012,N_1679,N_1979);
or U2013 (N_2013,N_1836,N_1564);
nor U2014 (N_2014,N_1263,N_1676);
nand U2015 (N_2015,N_1809,N_1035);
nor U2016 (N_2016,N_1707,N_1987);
nor U2017 (N_2017,N_1961,N_1055);
and U2018 (N_2018,N_1341,N_1473);
or U2019 (N_2019,N_1140,N_1506);
xor U2020 (N_2020,N_1838,N_1526);
and U2021 (N_2021,N_1163,N_1323);
nor U2022 (N_2022,N_1441,N_1629);
or U2023 (N_2023,N_1375,N_1688);
or U2024 (N_2024,N_1767,N_1092);
nor U2025 (N_2025,N_1068,N_1534);
nor U2026 (N_2026,N_1876,N_1805);
nor U2027 (N_2027,N_1978,N_1937);
or U2028 (N_2028,N_1089,N_1737);
nand U2029 (N_2029,N_1248,N_1336);
xnor U2030 (N_2030,N_1439,N_1061);
or U2031 (N_2031,N_1647,N_1057);
or U2032 (N_2032,N_1743,N_1875);
nand U2033 (N_2033,N_1954,N_1400);
nand U2034 (N_2034,N_1371,N_1255);
or U2035 (N_2035,N_1114,N_1939);
and U2036 (N_2036,N_1696,N_1643);
nand U2037 (N_2037,N_1626,N_1167);
or U2038 (N_2038,N_1952,N_1530);
xor U2039 (N_2039,N_1617,N_1386);
or U2040 (N_2040,N_1514,N_1548);
and U2041 (N_2041,N_1000,N_1218);
nor U2042 (N_2042,N_1656,N_1118);
nor U2043 (N_2043,N_1816,N_1121);
or U2044 (N_2044,N_1338,N_1886);
and U2045 (N_2045,N_1628,N_1977);
nor U2046 (N_2046,N_1754,N_1773);
and U2047 (N_2047,N_1370,N_1151);
or U2048 (N_2048,N_1863,N_1732);
or U2049 (N_2049,N_1851,N_1869);
nand U2050 (N_2050,N_1148,N_1559);
nand U2051 (N_2051,N_1858,N_1931);
nor U2052 (N_2052,N_1631,N_1162);
nor U2053 (N_2053,N_1137,N_1608);
nor U2054 (N_2054,N_1367,N_1822);
nand U2055 (N_2055,N_1919,N_1704);
nor U2056 (N_2056,N_1466,N_1281);
and U2057 (N_2057,N_1694,N_1106);
nor U2058 (N_2058,N_1357,N_1397);
or U2059 (N_2059,N_1495,N_1844);
xnor U2060 (N_2060,N_1882,N_1591);
and U2061 (N_2061,N_1158,N_1657);
nor U2062 (N_2062,N_1053,N_1031);
and U2063 (N_2063,N_1193,N_1999);
nand U2064 (N_2064,N_1642,N_1139);
or U2065 (N_2065,N_1319,N_1006);
xnor U2066 (N_2066,N_1761,N_1959);
and U2067 (N_2067,N_1475,N_1180);
nor U2068 (N_2068,N_1669,N_1906);
nand U2069 (N_2069,N_1685,N_1860);
and U2070 (N_2070,N_1077,N_1871);
xor U2071 (N_2071,N_1995,N_1101);
and U2072 (N_2072,N_1376,N_1533);
or U2073 (N_2073,N_1556,N_1010);
and U2074 (N_2074,N_1607,N_1346);
xnor U2075 (N_2075,N_1081,N_1490);
nor U2076 (N_2076,N_1765,N_1426);
nor U2077 (N_2077,N_1269,N_1394);
and U2078 (N_2078,N_1799,N_1115);
xor U2079 (N_2079,N_1476,N_1445);
or U2080 (N_2080,N_1678,N_1976);
and U2081 (N_2081,N_1098,N_1576);
or U2082 (N_2082,N_1827,N_1278);
or U2083 (N_2083,N_1048,N_1191);
nand U2084 (N_2084,N_1440,N_1717);
or U2085 (N_2085,N_1615,N_1360);
or U2086 (N_2086,N_1549,N_1909);
and U2087 (N_2087,N_1347,N_1627);
or U2088 (N_2088,N_1129,N_1892);
or U2089 (N_2089,N_1926,N_1254);
and U2090 (N_2090,N_1601,N_1308);
or U2091 (N_2091,N_1786,N_1412);
nand U2092 (N_2092,N_1214,N_1491);
nor U2093 (N_2093,N_1710,N_1333);
and U2094 (N_2094,N_1522,N_1618);
or U2095 (N_2095,N_1787,N_1573);
xor U2096 (N_2096,N_1368,N_1947);
or U2097 (N_2097,N_1009,N_1093);
nor U2098 (N_2098,N_1784,N_1410);
nor U2099 (N_2099,N_1974,N_1890);
or U2100 (N_2100,N_1049,N_1437);
or U2101 (N_2101,N_1293,N_1750);
or U2102 (N_2102,N_1971,N_1467);
and U2103 (N_2103,N_1966,N_1861);
and U2104 (N_2104,N_1528,N_1870);
nor U2105 (N_2105,N_1791,N_1880);
and U2106 (N_2106,N_1905,N_1488);
or U2107 (N_2107,N_1111,N_1683);
and U2108 (N_2108,N_1503,N_1550);
nor U2109 (N_2109,N_1337,N_1675);
nor U2110 (N_2110,N_1328,N_1087);
nand U2111 (N_2111,N_1431,N_1759);
nor U2112 (N_2112,N_1334,N_1982);
nand U2113 (N_2113,N_1687,N_1568);
nor U2114 (N_2114,N_1170,N_1945);
and U2115 (N_2115,N_1258,N_1243);
nand U2116 (N_2116,N_1249,N_1105);
and U2117 (N_2117,N_1998,N_1079);
nor U2118 (N_2118,N_1990,N_1135);
and U2119 (N_2119,N_1125,N_1877);
xor U2120 (N_2120,N_1157,N_1830);
nor U2121 (N_2121,N_1173,N_1078);
or U2122 (N_2122,N_1563,N_1814);
and U2123 (N_2123,N_1824,N_1419);
nand U2124 (N_2124,N_1235,N_1463);
nor U2125 (N_2125,N_1358,N_1697);
nor U2126 (N_2126,N_1505,N_1110);
or U2127 (N_2127,N_1407,N_1800);
and U2128 (N_2128,N_1690,N_1853);
nor U2129 (N_2129,N_1658,N_1525);
nor U2130 (N_2130,N_1315,N_1342);
or U2131 (N_2131,N_1794,N_1282);
and U2132 (N_2132,N_1655,N_1229);
nor U2133 (N_2133,N_1022,N_1044);
and U2134 (N_2134,N_1780,N_1703);
nand U2135 (N_2135,N_1545,N_1480);
and U2136 (N_2136,N_1382,N_1291);
or U2137 (N_2137,N_1438,N_1202);
or U2138 (N_2138,N_1963,N_1789);
xnor U2139 (N_2139,N_1872,N_1065);
or U2140 (N_2140,N_1884,N_1186);
or U2141 (N_2141,N_1973,N_1856);
and U2142 (N_2142,N_1728,N_1517);
or U2143 (N_2143,N_1693,N_1562);
nor U2144 (N_2144,N_1641,N_1741);
nand U2145 (N_2145,N_1623,N_1908);
nand U2146 (N_2146,N_1625,N_1147);
and U2147 (N_2147,N_1262,N_1819);
or U2148 (N_2148,N_1064,N_1590);
nor U2149 (N_2149,N_1459,N_1435);
nor U2150 (N_2150,N_1211,N_1016);
xor U2151 (N_2151,N_1721,N_1175);
and U2152 (N_2152,N_1216,N_1801);
and U2153 (N_2153,N_1510,N_1025);
xor U2154 (N_2154,N_1897,N_1793);
nor U2155 (N_2155,N_1661,N_1471);
and U2156 (N_2156,N_1402,N_1462);
nand U2157 (N_2157,N_1399,N_1667);
xor U2158 (N_2158,N_1456,N_1825);
and U2159 (N_2159,N_1726,N_1958);
and U2160 (N_2160,N_1640,N_1302);
nand U2161 (N_2161,N_1091,N_1239);
nand U2162 (N_2162,N_1415,N_1232);
or U2163 (N_2163,N_1578,N_1066);
and U2164 (N_2164,N_1390,N_1889);
and U2165 (N_2165,N_1881,N_1305);
nand U2166 (N_2166,N_1646,N_1117);
nor U2167 (N_2167,N_1088,N_1541);
and U2168 (N_2168,N_1544,N_1972);
and U2169 (N_2169,N_1828,N_1478);
and U2170 (N_2170,N_1532,N_1320);
nand U2171 (N_2171,N_1458,N_1953);
nor U2172 (N_2172,N_1206,N_1256);
nand U2173 (N_2173,N_1387,N_1233);
and U2174 (N_2174,N_1190,N_1352);
nor U2175 (N_2175,N_1936,N_1014);
xor U2176 (N_2176,N_1602,N_1662);
and U2177 (N_2177,N_1265,N_1705);
or U2178 (N_2178,N_1502,N_1450);
xor U2179 (N_2179,N_1489,N_1365);
nor U2180 (N_2180,N_1848,N_1831);
xnor U2181 (N_2181,N_1418,N_1635);
xnor U2182 (N_2182,N_1321,N_1547);
and U2183 (N_2183,N_1200,N_1046);
nand U2184 (N_2184,N_1969,N_1546);
and U2185 (N_2185,N_1454,N_1422);
and U2186 (N_2186,N_1424,N_1245);
nor U2187 (N_2187,N_1294,N_1901);
nand U2188 (N_2188,N_1330,N_1383);
xnor U2189 (N_2189,N_1501,N_1145);
nand U2190 (N_2190,N_1583,N_1090);
nand U2191 (N_2191,N_1482,N_1005);
nand U2192 (N_2192,N_1907,N_1063);
nor U2193 (N_2193,N_1826,N_1264);
xnor U2194 (N_2194,N_1497,N_1327);
xor U2195 (N_2195,N_1648,N_1485);
and U2196 (N_2196,N_1416,N_1771);
nor U2197 (N_2197,N_1981,N_1113);
or U2198 (N_2198,N_1509,N_1398);
or U2199 (N_2199,N_1748,N_1516);
or U2200 (N_2200,N_1785,N_1343);
and U2201 (N_2201,N_1774,N_1587);
nor U2202 (N_2202,N_1991,N_1701);
and U2203 (N_2203,N_1823,N_1080);
or U2204 (N_2204,N_1050,N_1592);
nor U2205 (N_2205,N_1266,N_1421);
and U2206 (N_2206,N_1849,N_1989);
nand U2207 (N_2207,N_1353,N_1363);
nor U2208 (N_2208,N_1192,N_1839);
nor U2209 (N_2209,N_1920,N_1900);
xnor U2210 (N_2210,N_1762,N_1613);
or U2211 (N_2211,N_1189,N_1130);
or U2212 (N_2212,N_1569,N_1903);
xnor U2213 (N_2213,N_1709,N_1700);
or U2214 (N_2214,N_1724,N_1252);
or U2215 (N_2215,N_1637,N_1520);
nand U2216 (N_2216,N_1619,N_1605);
or U2217 (N_2217,N_1116,N_1680);
nand U2218 (N_2218,N_1539,N_1795);
or U2219 (N_2219,N_1287,N_1841);
xor U2220 (N_2220,N_1301,N_1986);
or U2221 (N_2221,N_1408,N_1835);
nor U2222 (N_2222,N_1855,N_1925);
nand U2223 (N_2223,N_1146,N_1722);
nor U2224 (N_2224,N_1388,N_1150);
or U2225 (N_2225,N_1272,N_1362);
nand U2226 (N_2226,N_1531,N_1187);
nand U2227 (N_2227,N_1689,N_1873);
or U2228 (N_2228,N_1460,N_1013);
xor U2229 (N_2229,N_1734,N_1240);
nand U2230 (N_2230,N_1444,N_1120);
or U2231 (N_2231,N_1561,N_1716);
nor U2232 (N_2232,N_1712,N_1425);
and U2233 (N_2233,N_1535,N_1492);
and U2234 (N_2234,N_1723,N_1284);
nand U2235 (N_2235,N_1434,N_1949);
nand U2236 (N_2236,N_1332,N_1760);
nor U2237 (N_2237,N_1178,N_1843);
nand U2238 (N_2238,N_1040,N_1893);
nor U2239 (N_2239,N_1001,N_1599);
nor U2240 (N_2240,N_1913,N_1654);
and U2241 (N_2241,N_1630,N_1603);
or U2242 (N_2242,N_1929,N_1259);
nand U2243 (N_2243,N_1739,N_1725);
and U2244 (N_2244,N_1127,N_1477);
and U2245 (N_2245,N_1847,N_1677);
and U2246 (N_2246,N_1339,N_1985);
and U2247 (N_2247,N_1695,N_1666);
or U2248 (N_2248,N_1777,N_1983);
or U2249 (N_2249,N_1238,N_1567);
or U2250 (N_2250,N_1744,N_1234);
and U2251 (N_2251,N_1208,N_1711);
nor U2252 (N_2252,N_1638,N_1829);
or U2253 (N_2253,N_1496,N_1296);
and U2254 (N_2254,N_1279,N_1228);
or U2255 (N_2255,N_1404,N_1935);
nor U2256 (N_2256,N_1071,N_1790);
nand U2257 (N_2257,N_1042,N_1597);
nor U2258 (N_2258,N_1527,N_1915);
and U2259 (N_2259,N_1649,N_1409);
and U2260 (N_2260,N_1834,N_1176);
nand U2261 (N_2261,N_1275,N_1536);
nor U2262 (N_2262,N_1033,N_1928);
nand U2263 (N_2263,N_1751,N_1980);
nor U2264 (N_2264,N_1779,N_1134);
nor U2265 (N_2265,N_1310,N_1029);
and U2266 (N_2266,N_1883,N_1165);
xnor U2267 (N_2267,N_1644,N_1498);
or U2268 (N_2268,N_1833,N_1085);
xnor U2269 (N_2269,N_1560,N_1024);
and U2270 (N_2270,N_1359,N_1166);
xor U2271 (N_2271,N_1523,N_1914);
and U2272 (N_2272,N_1372,N_1624);
xor U2273 (N_2273,N_1464,N_1714);
and U2274 (N_2274,N_1069,N_1924);
and U2275 (N_2275,N_1699,N_1204);
nor U2276 (N_2276,N_1512,N_1420);
nor U2277 (N_2277,N_1210,N_1778);
and U2278 (N_2278,N_1572,N_1126);
and U2279 (N_2279,N_1933,N_1182);
nand U2280 (N_2280,N_1312,N_1131);
and U2281 (N_2281,N_1414,N_1538);
xor U2282 (N_2282,N_1322,N_1885);
and U2283 (N_2283,N_1988,N_1850);
nand U2284 (N_2284,N_1236,N_1852);
or U2285 (N_2285,N_1832,N_1329);
or U2286 (N_2286,N_1225,N_1610);
nand U2287 (N_2287,N_1045,N_1673);
and U2288 (N_2288,N_1486,N_1067);
xnor U2289 (N_2289,N_1529,N_1558);
or U2290 (N_2290,N_1300,N_1455);
nor U2291 (N_2291,N_1195,N_1465);
nor U2292 (N_2292,N_1447,N_1217);
nor U2293 (N_2293,N_1212,N_1096);
nor U2294 (N_2294,N_1348,N_1574);
nand U2295 (N_2295,N_1996,N_1027);
nor U2296 (N_2296,N_1866,N_1878);
nand U2297 (N_2297,N_1378,N_1566);
nor U2298 (N_2298,N_1749,N_1369);
xnor U2299 (N_2299,N_1059,N_1395);
nor U2300 (N_2300,N_1314,N_1956);
and U2301 (N_2301,N_1896,N_1161);
and U2302 (N_2302,N_1468,N_1316);
nor U2303 (N_2303,N_1804,N_1041);
or U2304 (N_2304,N_1168,N_1948);
xnor U2305 (N_2305,N_1060,N_1344);
nor U2306 (N_2306,N_1571,N_1902);
xnor U2307 (N_2307,N_1706,N_1413);
and U2308 (N_2308,N_1797,N_1788);
nor U2309 (N_2309,N_1614,N_1772);
nand U2310 (N_2310,N_1396,N_1012);
or U2311 (N_2311,N_1740,N_1224);
and U2312 (N_2312,N_1524,N_1201);
or U2313 (N_2313,N_1251,N_1997);
and U2314 (N_2314,N_1733,N_1433);
nand U2315 (N_2315,N_1663,N_1768);
and U2316 (N_2316,N_1008,N_1405);
nor U2317 (N_2317,N_1636,N_1250);
and U2318 (N_2318,N_1753,N_1515);
and U2319 (N_2319,N_1253,N_1283);
and U2320 (N_2320,N_1325,N_1718);
nand U2321 (N_2321,N_1155,N_1854);
and U2322 (N_2322,N_1598,N_1318);
and U2323 (N_2323,N_1209,N_1288);
or U2324 (N_2324,N_1719,N_1864);
or U2325 (N_2325,N_1109,N_1355);
nand U2326 (N_2326,N_1746,N_1557);
nand U2327 (N_2327,N_1796,N_1494);
nor U2328 (N_2328,N_1975,N_1241);
nand U2329 (N_2329,N_1374,N_1955);
nor U2330 (N_2330,N_1019,N_1859);
and U2331 (N_2331,N_1922,N_1286);
nand U2332 (N_2332,N_1713,N_1203);
xor U2333 (N_2333,N_1616,N_1609);
or U2334 (N_2334,N_1671,N_1682);
or U2335 (N_2335,N_1306,N_1917);
or U2336 (N_2336,N_1304,N_1645);
or U2337 (N_2337,N_1112,N_1226);
or U2338 (N_2338,N_1513,N_1152);
and U2339 (N_2339,N_1595,N_1075);
or U2340 (N_2340,N_1317,N_1992);
or U2341 (N_2341,N_1708,N_1715);
and U2342 (N_2342,N_1373,N_1073);
nand U2343 (N_2343,N_1199,N_1289);
nand U2344 (N_2344,N_1620,N_1303);
xnor U2345 (N_2345,N_1401,N_1132);
or U2346 (N_2346,N_1107,N_1076);
and U2347 (N_2347,N_1285,N_1565);
nand U2348 (N_2348,N_1361,N_1086);
or U2349 (N_2349,N_1895,N_1354);
nand U2350 (N_2350,N_1393,N_1257);
nand U2351 (N_2351,N_1820,N_1036);
or U2352 (N_2352,N_1807,N_1142);
nand U2353 (N_2353,N_1596,N_1461);
and U2354 (N_2354,N_1207,N_1391);
nand U2355 (N_2355,N_1552,N_1588);
nand U2356 (N_2356,N_1349,N_1702);
nand U2357 (N_2357,N_1582,N_1429);
and U2358 (N_2358,N_1551,N_1639);
and U2359 (N_2359,N_1965,N_1670);
nand U2360 (N_2360,N_1752,N_1198);
nor U2361 (N_2361,N_1943,N_1633);
nand U2362 (N_2362,N_1600,N_1769);
or U2363 (N_2363,N_1326,N_1665);
or U2364 (N_2364,N_1899,N_1857);
or U2365 (N_2365,N_1842,N_1280);
and U2366 (N_2366,N_1651,N_1222);
or U2367 (N_2367,N_1729,N_1011);
or U2368 (N_2368,N_1692,N_1944);
or U2369 (N_2369,N_1197,N_1023);
xor U2370 (N_2370,N_1570,N_1417);
or U2371 (N_2371,N_1385,N_1865);
or U2372 (N_2372,N_1575,N_1811);
nor U2373 (N_2373,N_1149,N_1124);
nor U2374 (N_2374,N_1058,N_1803);
and U2375 (N_2375,N_1470,N_1141);
nand U2376 (N_2376,N_1062,N_1122);
or U2377 (N_2377,N_1083,N_1755);
nand U2378 (N_2378,N_1172,N_1164);
or U2379 (N_2379,N_1862,N_1691);
nand U2380 (N_2380,N_1177,N_1313);
nand U2381 (N_2381,N_1698,N_1946);
and U2382 (N_2382,N_1812,N_1356);
and U2383 (N_2383,N_1584,N_1757);
nor U2384 (N_2384,N_1763,N_1039);
nor U2385 (N_2385,N_1964,N_1018);
xnor U2386 (N_2386,N_1507,N_1267);
nand U2387 (N_2387,N_1276,N_1518);
nor U2388 (N_2388,N_1521,N_1776);
nor U2389 (N_2389,N_1021,N_1268);
nor U2390 (N_2390,N_1867,N_1580);
nor U2391 (N_2391,N_1668,N_1511);
nor U2392 (N_2392,N_1674,N_1221);
nand U2393 (N_2393,N_1612,N_1123);
nand U2394 (N_2394,N_1951,N_1967);
nand U2395 (N_2395,N_1143,N_1481);
nor U2396 (N_2396,N_1542,N_1446);
nor U2397 (N_2397,N_1219,N_1934);
or U2398 (N_2398,N_1984,N_1270);
and U2399 (N_2399,N_1295,N_1099);
nor U2400 (N_2400,N_1103,N_1783);
and U2401 (N_2401,N_1084,N_1821);
xnor U2402 (N_2402,N_1894,N_1868);
nor U2403 (N_2403,N_1100,N_1766);
xnor U2404 (N_2404,N_1493,N_1891);
nand U2405 (N_2405,N_1730,N_1888);
or U2406 (N_2406,N_1043,N_1727);
and U2407 (N_2407,N_1652,N_1457);
nor U2408 (N_2408,N_1810,N_1030);
nand U2409 (N_2409,N_1171,N_1159);
nor U2410 (N_2410,N_1581,N_1664);
and U2411 (N_2411,N_1519,N_1994);
and U2412 (N_2412,N_1802,N_1156);
or U2413 (N_2413,N_1846,N_1593);
or U2414 (N_2414,N_1938,N_1781);
nand U2415 (N_2415,N_1183,N_1144);
nor U2416 (N_2416,N_1443,N_1927);
and U2417 (N_2417,N_1817,N_1735);
nor U2418 (N_2418,N_1188,N_1921);
nor U2419 (N_2419,N_1960,N_1451);
xor U2420 (N_2420,N_1324,N_1034);
nor U2421 (N_2421,N_1585,N_1345);
xor U2422 (N_2422,N_1104,N_1095);
nand U2423 (N_2423,N_1003,N_1020);
nor U2424 (N_2424,N_1277,N_1589);
xnor U2425 (N_2425,N_1350,N_1453);
nand U2426 (N_2426,N_1553,N_1056);
nand U2427 (N_2427,N_1950,N_1611);
or U2428 (N_2428,N_1923,N_1879);
and U2429 (N_2429,N_1579,N_1381);
nand U2430 (N_2430,N_1227,N_1745);
nand U2431 (N_2431,N_1968,N_1377);
or U2432 (N_2432,N_1051,N_1017);
nand U2433 (N_2433,N_1244,N_1004);
nand U2434 (N_2434,N_1340,N_1594);
nor U2435 (N_2435,N_1423,N_1160);
nor U2436 (N_2436,N_1634,N_1436);
or U2437 (N_2437,N_1543,N_1185);
or U2438 (N_2438,N_1054,N_1411);
and U2439 (N_2439,N_1430,N_1932);
nand U2440 (N_2440,N_1384,N_1174);
and U2441 (N_2441,N_1184,N_1213);
or U2442 (N_2442,N_1499,N_1271);
nor U2443 (N_2443,N_1366,N_1940);
and U2444 (N_2444,N_1299,N_1782);
and U2445 (N_2445,N_1230,N_1038);
nor U2446 (N_2446,N_1577,N_1364);
and U2447 (N_2447,N_1942,N_1500);
nand U2448 (N_2448,N_1392,N_1970);
nor U2449 (N_2449,N_1874,N_1898);
and U2450 (N_2450,N_1941,N_1205);
and U2451 (N_2451,N_1448,N_1102);
or U2452 (N_2452,N_1309,N_1806);
or U2453 (N_2453,N_1179,N_1169);
nand U2454 (N_2454,N_1479,N_1911);
nand U2455 (N_2455,N_1916,N_1604);
xor U2456 (N_2456,N_1736,N_1672);
or U2457 (N_2457,N_1153,N_1813);
nand U2458 (N_2458,N_1047,N_1311);
or U2459 (N_2459,N_1845,N_1052);
nor U2460 (N_2460,N_1442,N_1483);
nand U2461 (N_2461,N_1403,N_1260);
nand U2462 (N_2462,N_1072,N_1351);
nand U2463 (N_2463,N_1775,N_1136);
nor U2464 (N_2464,N_1792,N_1196);
nand U2465 (N_2465,N_1261,N_1380);
and U2466 (N_2466,N_1428,N_1007);
and U2467 (N_2467,N_1070,N_1215);
or U2468 (N_2468,N_1469,N_1742);
xnor U2469 (N_2469,N_1770,N_1837);
xor U2470 (N_2470,N_1406,N_1720);
and U2471 (N_2471,N_1181,N_1242);
nand U2472 (N_2472,N_1930,N_1133);
or U2473 (N_2473,N_1290,N_1119);
or U2474 (N_2474,N_1307,N_1273);
nand U2475 (N_2475,N_1237,N_1231);
nor U2476 (N_2476,N_1432,N_1247);
nor U2477 (N_2477,N_1622,N_1487);
and U2478 (N_2478,N_1660,N_1910);
nor U2479 (N_2479,N_1298,N_1606);
or U2480 (N_2480,N_1747,N_1621);
or U2481 (N_2481,N_1540,N_1015);
nand U2482 (N_2482,N_1918,N_1128);
or U2483 (N_2483,N_1554,N_1756);
and U2484 (N_2484,N_1074,N_1082);
nor U2485 (N_2485,N_1331,N_1094);
nand U2486 (N_2486,N_1686,N_1389);
nand U2487 (N_2487,N_1274,N_1028);
or U2488 (N_2488,N_1026,N_1818);
xnor U2489 (N_2489,N_1246,N_1650);
nor U2490 (N_2490,N_1292,N_1032);
nor U2491 (N_2491,N_1764,N_1452);
nand U2492 (N_2492,N_1097,N_1297);
nor U2493 (N_2493,N_1504,N_1220);
xnor U2494 (N_2494,N_1484,N_1154);
and U2495 (N_2495,N_1758,N_1993);
or U2496 (N_2496,N_1474,N_1037);
nor U2497 (N_2497,N_1808,N_1957);
nand U2498 (N_2498,N_1223,N_1002);
and U2499 (N_2499,N_1449,N_1681);
nor U2500 (N_2500,N_1566,N_1632);
or U2501 (N_2501,N_1426,N_1913);
and U2502 (N_2502,N_1062,N_1590);
nand U2503 (N_2503,N_1396,N_1673);
and U2504 (N_2504,N_1596,N_1437);
and U2505 (N_2505,N_1612,N_1552);
and U2506 (N_2506,N_1250,N_1280);
nand U2507 (N_2507,N_1585,N_1252);
nand U2508 (N_2508,N_1718,N_1590);
xnor U2509 (N_2509,N_1061,N_1938);
and U2510 (N_2510,N_1218,N_1260);
nor U2511 (N_2511,N_1950,N_1400);
and U2512 (N_2512,N_1588,N_1631);
nand U2513 (N_2513,N_1084,N_1950);
nand U2514 (N_2514,N_1432,N_1556);
nand U2515 (N_2515,N_1576,N_1974);
nand U2516 (N_2516,N_1835,N_1154);
nand U2517 (N_2517,N_1088,N_1476);
xnor U2518 (N_2518,N_1300,N_1980);
and U2519 (N_2519,N_1129,N_1012);
and U2520 (N_2520,N_1784,N_1022);
or U2521 (N_2521,N_1924,N_1277);
or U2522 (N_2522,N_1213,N_1144);
nor U2523 (N_2523,N_1701,N_1146);
nand U2524 (N_2524,N_1781,N_1969);
and U2525 (N_2525,N_1482,N_1657);
nand U2526 (N_2526,N_1301,N_1878);
xnor U2527 (N_2527,N_1024,N_1931);
nor U2528 (N_2528,N_1708,N_1076);
nand U2529 (N_2529,N_1704,N_1458);
nor U2530 (N_2530,N_1125,N_1370);
and U2531 (N_2531,N_1464,N_1100);
nand U2532 (N_2532,N_1505,N_1807);
nand U2533 (N_2533,N_1086,N_1221);
or U2534 (N_2534,N_1591,N_1901);
nor U2535 (N_2535,N_1722,N_1340);
nor U2536 (N_2536,N_1336,N_1005);
and U2537 (N_2537,N_1321,N_1428);
nand U2538 (N_2538,N_1355,N_1161);
nor U2539 (N_2539,N_1275,N_1087);
or U2540 (N_2540,N_1586,N_1987);
or U2541 (N_2541,N_1044,N_1005);
nor U2542 (N_2542,N_1545,N_1152);
xor U2543 (N_2543,N_1175,N_1521);
and U2544 (N_2544,N_1605,N_1823);
or U2545 (N_2545,N_1683,N_1344);
xnor U2546 (N_2546,N_1403,N_1549);
and U2547 (N_2547,N_1136,N_1164);
and U2548 (N_2548,N_1491,N_1628);
or U2549 (N_2549,N_1356,N_1848);
nand U2550 (N_2550,N_1075,N_1701);
nor U2551 (N_2551,N_1854,N_1646);
nand U2552 (N_2552,N_1979,N_1664);
nand U2553 (N_2553,N_1887,N_1495);
and U2554 (N_2554,N_1732,N_1825);
nor U2555 (N_2555,N_1226,N_1720);
xor U2556 (N_2556,N_1454,N_1955);
nand U2557 (N_2557,N_1519,N_1513);
nor U2558 (N_2558,N_1252,N_1299);
and U2559 (N_2559,N_1556,N_1894);
xnor U2560 (N_2560,N_1817,N_1696);
or U2561 (N_2561,N_1812,N_1315);
nand U2562 (N_2562,N_1421,N_1106);
nand U2563 (N_2563,N_1408,N_1523);
nor U2564 (N_2564,N_1705,N_1922);
nor U2565 (N_2565,N_1304,N_1985);
and U2566 (N_2566,N_1117,N_1662);
and U2567 (N_2567,N_1935,N_1991);
and U2568 (N_2568,N_1517,N_1190);
nor U2569 (N_2569,N_1480,N_1075);
and U2570 (N_2570,N_1897,N_1847);
or U2571 (N_2571,N_1541,N_1985);
nand U2572 (N_2572,N_1904,N_1634);
nand U2573 (N_2573,N_1080,N_1544);
and U2574 (N_2574,N_1294,N_1894);
or U2575 (N_2575,N_1312,N_1688);
or U2576 (N_2576,N_1018,N_1500);
nor U2577 (N_2577,N_1080,N_1176);
or U2578 (N_2578,N_1013,N_1170);
xnor U2579 (N_2579,N_1743,N_1764);
and U2580 (N_2580,N_1114,N_1669);
or U2581 (N_2581,N_1712,N_1816);
or U2582 (N_2582,N_1941,N_1956);
nand U2583 (N_2583,N_1043,N_1407);
nor U2584 (N_2584,N_1180,N_1680);
nor U2585 (N_2585,N_1156,N_1876);
or U2586 (N_2586,N_1790,N_1679);
nand U2587 (N_2587,N_1996,N_1505);
nor U2588 (N_2588,N_1382,N_1595);
nor U2589 (N_2589,N_1258,N_1556);
nand U2590 (N_2590,N_1946,N_1811);
xor U2591 (N_2591,N_1424,N_1009);
or U2592 (N_2592,N_1178,N_1425);
nor U2593 (N_2593,N_1901,N_1238);
and U2594 (N_2594,N_1993,N_1721);
or U2595 (N_2595,N_1507,N_1239);
nor U2596 (N_2596,N_1977,N_1270);
nor U2597 (N_2597,N_1139,N_1797);
or U2598 (N_2598,N_1171,N_1415);
nor U2599 (N_2599,N_1209,N_1213);
nor U2600 (N_2600,N_1276,N_1600);
xnor U2601 (N_2601,N_1120,N_1144);
or U2602 (N_2602,N_1504,N_1487);
and U2603 (N_2603,N_1899,N_1717);
nand U2604 (N_2604,N_1547,N_1002);
nor U2605 (N_2605,N_1341,N_1664);
xor U2606 (N_2606,N_1589,N_1054);
nand U2607 (N_2607,N_1597,N_1575);
nand U2608 (N_2608,N_1913,N_1243);
xor U2609 (N_2609,N_1659,N_1412);
or U2610 (N_2610,N_1550,N_1163);
nand U2611 (N_2611,N_1611,N_1642);
or U2612 (N_2612,N_1571,N_1757);
nand U2613 (N_2613,N_1737,N_1577);
nor U2614 (N_2614,N_1317,N_1402);
nor U2615 (N_2615,N_1909,N_1581);
nand U2616 (N_2616,N_1612,N_1570);
xnor U2617 (N_2617,N_1491,N_1076);
nand U2618 (N_2618,N_1522,N_1141);
and U2619 (N_2619,N_1975,N_1553);
and U2620 (N_2620,N_1090,N_1556);
nor U2621 (N_2621,N_1577,N_1157);
nand U2622 (N_2622,N_1871,N_1055);
and U2623 (N_2623,N_1772,N_1304);
or U2624 (N_2624,N_1325,N_1124);
or U2625 (N_2625,N_1054,N_1092);
nor U2626 (N_2626,N_1916,N_1280);
and U2627 (N_2627,N_1671,N_1496);
xnor U2628 (N_2628,N_1755,N_1979);
or U2629 (N_2629,N_1606,N_1723);
or U2630 (N_2630,N_1953,N_1167);
and U2631 (N_2631,N_1876,N_1989);
and U2632 (N_2632,N_1788,N_1204);
and U2633 (N_2633,N_1104,N_1321);
or U2634 (N_2634,N_1082,N_1922);
nor U2635 (N_2635,N_1879,N_1339);
nor U2636 (N_2636,N_1646,N_1071);
xnor U2637 (N_2637,N_1152,N_1644);
xnor U2638 (N_2638,N_1239,N_1159);
nand U2639 (N_2639,N_1444,N_1600);
or U2640 (N_2640,N_1021,N_1095);
nand U2641 (N_2641,N_1942,N_1293);
and U2642 (N_2642,N_1640,N_1217);
xnor U2643 (N_2643,N_1440,N_1806);
or U2644 (N_2644,N_1477,N_1405);
nand U2645 (N_2645,N_1517,N_1100);
and U2646 (N_2646,N_1917,N_1112);
nand U2647 (N_2647,N_1645,N_1029);
nor U2648 (N_2648,N_1687,N_1048);
nand U2649 (N_2649,N_1305,N_1287);
nor U2650 (N_2650,N_1431,N_1853);
nand U2651 (N_2651,N_1185,N_1124);
nand U2652 (N_2652,N_1001,N_1671);
and U2653 (N_2653,N_1295,N_1020);
or U2654 (N_2654,N_1827,N_1047);
or U2655 (N_2655,N_1161,N_1685);
nor U2656 (N_2656,N_1555,N_1263);
or U2657 (N_2657,N_1377,N_1927);
or U2658 (N_2658,N_1767,N_1027);
or U2659 (N_2659,N_1701,N_1516);
or U2660 (N_2660,N_1926,N_1755);
and U2661 (N_2661,N_1341,N_1053);
nor U2662 (N_2662,N_1915,N_1304);
nor U2663 (N_2663,N_1943,N_1334);
nand U2664 (N_2664,N_1681,N_1486);
nand U2665 (N_2665,N_1971,N_1634);
or U2666 (N_2666,N_1315,N_1231);
xor U2667 (N_2667,N_1397,N_1059);
and U2668 (N_2668,N_1520,N_1841);
xnor U2669 (N_2669,N_1803,N_1795);
nor U2670 (N_2670,N_1746,N_1947);
and U2671 (N_2671,N_1819,N_1110);
and U2672 (N_2672,N_1905,N_1860);
or U2673 (N_2673,N_1044,N_1941);
or U2674 (N_2674,N_1991,N_1642);
nor U2675 (N_2675,N_1061,N_1303);
and U2676 (N_2676,N_1878,N_1461);
or U2677 (N_2677,N_1578,N_1805);
or U2678 (N_2678,N_1762,N_1399);
or U2679 (N_2679,N_1634,N_1901);
or U2680 (N_2680,N_1735,N_1542);
and U2681 (N_2681,N_1737,N_1556);
and U2682 (N_2682,N_1424,N_1023);
and U2683 (N_2683,N_1520,N_1792);
or U2684 (N_2684,N_1593,N_1869);
nor U2685 (N_2685,N_1556,N_1414);
xnor U2686 (N_2686,N_1216,N_1091);
nand U2687 (N_2687,N_1355,N_1882);
nand U2688 (N_2688,N_1934,N_1500);
xor U2689 (N_2689,N_1378,N_1805);
and U2690 (N_2690,N_1718,N_1238);
or U2691 (N_2691,N_1886,N_1352);
or U2692 (N_2692,N_1309,N_1877);
nand U2693 (N_2693,N_1572,N_1780);
nand U2694 (N_2694,N_1264,N_1413);
or U2695 (N_2695,N_1347,N_1324);
and U2696 (N_2696,N_1657,N_1650);
or U2697 (N_2697,N_1803,N_1512);
and U2698 (N_2698,N_1216,N_1404);
nand U2699 (N_2699,N_1801,N_1194);
nor U2700 (N_2700,N_1009,N_1017);
xor U2701 (N_2701,N_1572,N_1477);
nand U2702 (N_2702,N_1309,N_1009);
nand U2703 (N_2703,N_1218,N_1550);
and U2704 (N_2704,N_1370,N_1169);
nor U2705 (N_2705,N_1573,N_1921);
or U2706 (N_2706,N_1244,N_1232);
or U2707 (N_2707,N_1434,N_1430);
and U2708 (N_2708,N_1007,N_1878);
nand U2709 (N_2709,N_1250,N_1216);
or U2710 (N_2710,N_1195,N_1880);
nor U2711 (N_2711,N_1462,N_1308);
or U2712 (N_2712,N_1159,N_1752);
nand U2713 (N_2713,N_1255,N_1167);
nor U2714 (N_2714,N_1284,N_1955);
xnor U2715 (N_2715,N_1183,N_1584);
xor U2716 (N_2716,N_1721,N_1964);
nor U2717 (N_2717,N_1669,N_1947);
xor U2718 (N_2718,N_1982,N_1333);
and U2719 (N_2719,N_1057,N_1282);
and U2720 (N_2720,N_1882,N_1736);
nand U2721 (N_2721,N_1953,N_1113);
nor U2722 (N_2722,N_1659,N_1068);
xor U2723 (N_2723,N_1504,N_1583);
and U2724 (N_2724,N_1342,N_1956);
or U2725 (N_2725,N_1452,N_1658);
and U2726 (N_2726,N_1955,N_1978);
or U2727 (N_2727,N_1201,N_1279);
nand U2728 (N_2728,N_1694,N_1165);
or U2729 (N_2729,N_1610,N_1937);
xnor U2730 (N_2730,N_1254,N_1260);
nor U2731 (N_2731,N_1327,N_1426);
or U2732 (N_2732,N_1998,N_1733);
and U2733 (N_2733,N_1781,N_1120);
or U2734 (N_2734,N_1469,N_1887);
nand U2735 (N_2735,N_1072,N_1558);
or U2736 (N_2736,N_1320,N_1890);
and U2737 (N_2737,N_1167,N_1829);
or U2738 (N_2738,N_1282,N_1850);
nand U2739 (N_2739,N_1486,N_1286);
and U2740 (N_2740,N_1206,N_1138);
nand U2741 (N_2741,N_1830,N_1467);
nand U2742 (N_2742,N_1479,N_1870);
nor U2743 (N_2743,N_1885,N_1196);
nor U2744 (N_2744,N_1350,N_1123);
nand U2745 (N_2745,N_1635,N_1085);
nand U2746 (N_2746,N_1088,N_1578);
or U2747 (N_2747,N_1024,N_1719);
nand U2748 (N_2748,N_1483,N_1958);
nand U2749 (N_2749,N_1542,N_1063);
or U2750 (N_2750,N_1186,N_1698);
or U2751 (N_2751,N_1276,N_1644);
nor U2752 (N_2752,N_1545,N_1846);
nand U2753 (N_2753,N_1275,N_1249);
nand U2754 (N_2754,N_1382,N_1734);
and U2755 (N_2755,N_1686,N_1405);
or U2756 (N_2756,N_1857,N_1036);
nor U2757 (N_2757,N_1667,N_1046);
nand U2758 (N_2758,N_1400,N_1136);
and U2759 (N_2759,N_1414,N_1167);
and U2760 (N_2760,N_1854,N_1049);
nand U2761 (N_2761,N_1133,N_1856);
nand U2762 (N_2762,N_1087,N_1134);
nand U2763 (N_2763,N_1037,N_1451);
nor U2764 (N_2764,N_1951,N_1971);
xnor U2765 (N_2765,N_1460,N_1714);
nor U2766 (N_2766,N_1261,N_1736);
nand U2767 (N_2767,N_1286,N_1133);
xor U2768 (N_2768,N_1405,N_1806);
nor U2769 (N_2769,N_1611,N_1721);
nand U2770 (N_2770,N_1747,N_1668);
or U2771 (N_2771,N_1319,N_1637);
nor U2772 (N_2772,N_1518,N_1901);
or U2773 (N_2773,N_1429,N_1342);
nor U2774 (N_2774,N_1950,N_1643);
nor U2775 (N_2775,N_1208,N_1147);
nor U2776 (N_2776,N_1377,N_1638);
and U2777 (N_2777,N_1327,N_1038);
or U2778 (N_2778,N_1706,N_1660);
nor U2779 (N_2779,N_1421,N_1944);
and U2780 (N_2780,N_1994,N_1837);
xor U2781 (N_2781,N_1952,N_1326);
nand U2782 (N_2782,N_1380,N_1019);
and U2783 (N_2783,N_1953,N_1352);
or U2784 (N_2784,N_1870,N_1330);
or U2785 (N_2785,N_1698,N_1603);
nand U2786 (N_2786,N_1504,N_1946);
nor U2787 (N_2787,N_1750,N_1418);
nand U2788 (N_2788,N_1181,N_1078);
nand U2789 (N_2789,N_1962,N_1457);
or U2790 (N_2790,N_1868,N_1472);
xnor U2791 (N_2791,N_1956,N_1267);
nand U2792 (N_2792,N_1592,N_1698);
and U2793 (N_2793,N_1392,N_1695);
or U2794 (N_2794,N_1928,N_1071);
nand U2795 (N_2795,N_1141,N_1927);
nor U2796 (N_2796,N_1791,N_1782);
xnor U2797 (N_2797,N_1952,N_1426);
or U2798 (N_2798,N_1035,N_1946);
and U2799 (N_2799,N_1776,N_1772);
and U2800 (N_2800,N_1421,N_1366);
nand U2801 (N_2801,N_1082,N_1662);
nor U2802 (N_2802,N_1481,N_1973);
nor U2803 (N_2803,N_1794,N_1736);
nand U2804 (N_2804,N_1644,N_1317);
nor U2805 (N_2805,N_1800,N_1978);
nand U2806 (N_2806,N_1052,N_1431);
and U2807 (N_2807,N_1171,N_1958);
and U2808 (N_2808,N_1661,N_1455);
nand U2809 (N_2809,N_1071,N_1123);
or U2810 (N_2810,N_1775,N_1265);
xnor U2811 (N_2811,N_1426,N_1820);
nor U2812 (N_2812,N_1893,N_1453);
nor U2813 (N_2813,N_1639,N_1798);
nand U2814 (N_2814,N_1388,N_1410);
or U2815 (N_2815,N_1026,N_1116);
or U2816 (N_2816,N_1509,N_1715);
or U2817 (N_2817,N_1749,N_1127);
and U2818 (N_2818,N_1421,N_1343);
nor U2819 (N_2819,N_1568,N_1846);
nand U2820 (N_2820,N_1429,N_1386);
and U2821 (N_2821,N_1194,N_1043);
nor U2822 (N_2822,N_1977,N_1785);
nand U2823 (N_2823,N_1609,N_1718);
nor U2824 (N_2824,N_1708,N_1167);
nor U2825 (N_2825,N_1779,N_1923);
or U2826 (N_2826,N_1742,N_1797);
and U2827 (N_2827,N_1196,N_1736);
nand U2828 (N_2828,N_1986,N_1977);
and U2829 (N_2829,N_1927,N_1919);
or U2830 (N_2830,N_1378,N_1714);
nor U2831 (N_2831,N_1192,N_1033);
nor U2832 (N_2832,N_1069,N_1020);
nor U2833 (N_2833,N_1406,N_1917);
or U2834 (N_2834,N_1964,N_1615);
or U2835 (N_2835,N_1572,N_1506);
and U2836 (N_2836,N_1405,N_1591);
xor U2837 (N_2837,N_1402,N_1805);
nand U2838 (N_2838,N_1119,N_1635);
nand U2839 (N_2839,N_1623,N_1155);
nor U2840 (N_2840,N_1928,N_1609);
nand U2841 (N_2841,N_1011,N_1717);
or U2842 (N_2842,N_1738,N_1564);
nand U2843 (N_2843,N_1215,N_1524);
nor U2844 (N_2844,N_1128,N_1332);
or U2845 (N_2845,N_1993,N_1043);
and U2846 (N_2846,N_1312,N_1656);
and U2847 (N_2847,N_1186,N_1431);
nand U2848 (N_2848,N_1165,N_1986);
nor U2849 (N_2849,N_1362,N_1732);
and U2850 (N_2850,N_1077,N_1354);
xor U2851 (N_2851,N_1858,N_1415);
and U2852 (N_2852,N_1250,N_1495);
nor U2853 (N_2853,N_1748,N_1545);
or U2854 (N_2854,N_1448,N_1376);
nand U2855 (N_2855,N_1448,N_1031);
and U2856 (N_2856,N_1938,N_1673);
and U2857 (N_2857,N_1992,N_1412);
or U2858 (N_2858,N_1005,N_1353);
xor U2859 (N_2859,N_1785,N_1565);
nor U2860 (N_2860,N_1758,N_1640);
or U2861 (N_2861,N_1266,N_1630);
nand U2862 (N_2862,N_1693,N_1151);
or U2863 (N_2863,N_1112,N_1792);
and U2864 (N_2864,N_1182,N_1812);
and U2865 (N_2865,N_1562,N_1709);
nor U2866 (N_2866,N_1145,N_1553);
nand U2867 (N_2867,N_1428,N_1461);
nor U2868 (N_2868,N_1718,N_1715);
nand U2869 (N_2869,N_1770,N_1502);
and U2870 (N_2870,N_1755,N_1427);
nor U2871 (N_2871,N_1486,N_1096);
nand U2872 (N_2872,N_1239,N_1285);
xor U2873 (N_2873,N_1679,N_1783);
nand U2874 (N_2874,N_1734,N_1685);
nor U2875 (N_2875,N_1389,N_1507);
xnor U2876 (N_2876,N_1793,N_1130);
and U2877 (N_2877,N_1244,N_1566);
nor U2878 (N_2878,N_1723,N_1540);
nor U2879 (N_2879,N_1586,N_1422);
or U2880 (N_2880,N_1608,N_1583);
nor U2881 (N_2881,N_1546,N_1859);
and U2882 (N_2882,N_1079,N_1124);
and U2883 (N_2883,N_1727,N_1774);
xor U2884 (N_2884,N_1892,N_1294);
nand U2885 (N_2885,N_1067,N_1677);
xor U2886 (N_2886,N_1196,N_1120);
nor U2887 (N_2887,N_1802,N_1051);
and U2888 (N_2888,N_1985,N_1169);
nor U2889 (N_2889,N_1606,N_1259);
nor U2890 (N_2890,N_1923,N_1991);
xor U2891 (N_2891,N_1297,N_1149);
nand U2892 (N_2892,N_1915,N_1065);
or U2893 (N_2893,N_1529,N_1225);
xor U2894 (N_2894,N_1232,N_1250);
and U2895 (N_2895,N_1549,N_1180);
nand U2896 (N_2896,N_1762,N_1834);
or U2897 (N_2897,N_1495,N_1290);
and U2898 (N_2898,N_1664,N_1050);
and U2899 (N_2899,N_1381,N_1557);
or U2900 (N_2900,N_1403,N_1331);
nor U2901 (N_2901,N_1028,N_1397);
nor U2902 (N_2902,N_1956,N_1527);
or U2903 (N_2903,N_1442,N_1729);
xnor U2904 (N_2904,N_1928,N_1077);
or U2905 (N_2905,N_1825,N_1890);
nand U2906 (N_2906,N_1924,N_1973);
nor U2907 (N_2907,N_1439,N_1320);
nand U2908 (N_2908,N_1685,N_1549);
nor U2909 (N_2909,N_1029,N_1422);
or U2910 (N_2910,N_1129,N_1493);
nor U2911 (N_2911,N_1803,N_1157);
and U2912 (N_2912,N_1810,N_1181);
nor U2913 (N_2913,N_1912,N_1265);
nor U2914 (N_2914,N_1793,N_1119);
or U2915 (N_2915,N_1573,N_1758);
nor U2916 (N_2916,N_1923,N_1378);
nor U2917 (N_2917,N_1148,N_1633);
or U2918 (N_2918,N_1688,N_1231);
nor U2919 (N_2919,N_1629,N_1787);
or U2920 (N_2920,N_1721,N_1824);
xnor U2921 (N_2921,N_1418,N_1217);
or U2922 (N_2922,N_1270,N_1508);
and U2923 (N_2923,N_1177,N_1122);
or U2924 (N_2924,N_1755,N_1993);
xor U2925 (N_2925,N_1328,N_1842);
or U2926 (N_2926,N_1826,N_1852);
nand U2927 (N_2927,N_1292,N_1065);
xor U2928 (N_2928,N_1280,N_1439);
nor U2929 (N_2929,N_1177,N_1591);
and U2930 (N_2930,N_1272,N_1090);
nor U2931 (N_2931,N_1942,N_1759);
xnor U2932 (N_2932,N_1904,N_1937);
nor U2933 (N_2933,N_1829,N_1450);
nand U2934 (N_2934,N_1711,N_1986);
nor U2935 (N_2935,N_1256,N_1339);
or U2936 (N_2936,N_1312,N_1702);
nand U2937 (N_2937,N_1699,N_1826);
nor U2938 (N_2938,N_1549,N_1599);
or U2939 (N_2939,N_1952,N_1366);
and U2940 (N_2940,N_1974,N_1772);
and U2941 (N_2941,N_1074,N_1880);
and U2942 (N_2942,N_1160,N_1494);
nor U2943 (N_2943,N_1382,N_1706);
nor U2944 (N_2944,N_1583,N_1953);
nand U2945 (N_2945,N_1474,N_1541);
nand U2946 (N_2946,N_1920,N_1131);
nand U2947 (N_2947,N_1256,N_1808);
and U2948 (N_2948,N_1785,N_1667);
nand U2949 (N_2949,N_1474,N_1944);
nand U2950 (N_2950,N_1214,N_1280);
and U2951 (N_2951,N_1537,N_1799);
and U2952 (N_2952,N_1215,N_1648);
and U2953 (N_2953,N_1088,N_1648);
and U2954 (N_2954,N_1768,N_1388);
or U2955 (N_2955,N_1106,N_1286);
nor U2956 (N_2956,N_1626,N_1505);
nor U2957 (N_2957,N_1413,N_1785);
nor U2958 (N_2958,N_1828,N_1526);
and U2959 (N_2959,N_1410,N_1545);
nor U2960 (N_2960,N_1747,N_1699);
xnor U2961 (N_2961,N_1806,N_1654);
or U2962 (N_2962,N_1873,N_1665);
nand U2963 (N_2963,N_1969,N_1778);
nor U2964 (N_2964,N_1818,N_1904);
and U2965 (N_2965,N_1251,N_1633);
nand U2966 (N_2966,N_1968,N_1199);
or U2967 (N_2967,N_1640,N_1274);
nor U2968 (N_2968,N_1349,N_1046);
nor U2969 (N_2969,N_1712,N_1494);
or U2970 (N_2970,N_1639,N_1656);
and U2971 (N_2971,N_1497,N_1210);
nor U2972 (N_2972,N_1943,N_1052);
or U2973 (N_2973,N_1231,N_1233);
xor U2974 (N_2974,N_1476,N_1170);
and U2975 (N_2975,N_1006,N_1052);
or U2976 (N_2976,N_1290,N_1034);
or U2977 (N_2977,N_1965,N_1980);
nor U2978 (N_2978,N_1568,N_1031);
or U2979 (N_2979,N_1452,N_1013);
nor U2980 (N_2980,N_1609,N_1812);
and U2981 (N_2981,N_1569,N_1763);
or U2982 (N_2982,N_1818,N_1848);
and U2983 (N_2983,N_1465,N_1426);
nand U2984 (N_2984,N_1917,N_1669);
nor U2985 (N_2985,N_1700,N_1113);
nand U2986 (N_2986,N_1113,N_1562);
xnor U2987 (N_2987,N_1602,N_1941);
and U2988 (N_2988,N_1816,N_1245);
and U2989 (N_2989,N_1517,N_1660);
nand U2990 (N_2990,N_1946,N_1431);
or U2991 (N_2991,N_1917,N_1769);
nand U2992 (N_2992,N_1632,N_1248);
nor U2993 (N_2993,N_1352,N_1337);
nor U2994 (N_2994,N_1432,N_1614);
or U2995 (N_2995,N_1240,N_1180);
nor U2996 (N_2996,N_1430,N_1423);
nand U2997 (N_2997,N_1844,N_1210);
and U2998 (N_2998,N_1092,N_1957);
nor U2999 (N_2999,N_1659,N_1270);
and U3000 (N_3000,N_2137,N_2093);
nand U3001 (N_3001,N_2324,N_2491);
or U3002 (N_3002,N_2277,N_2727);
nor U3003 (N_3003,N_2524,N_2446);
or U3004 (N_3004,N_2669,N_2150);
xor U3005 (N_3005,N_2144,N_2356);
xor U3006 (N_3006,N_2950,N_2306);
xnor U3007 (N_3007,N_2741,N_2906);
and U3008 (N_3008,N_2748,N_2660);
or U3009 (N_3009,N_2156,N_2280);
nor U3010 (N_3010,N_2212,N_2803);
and U3011 (N_3011,N_2094,N_2370);
nand U3012 (N_3012,N_2722,N_2486);
and U3013 (N_3013,N_2469,N_2892);
nand U3014 (N_3014,N_2301,N_2537);
nand U3015 (N_3015,N_2864,N_2412);
nor U3016 (N_3016,N_2082,N_2522);
nand U3017 (N_3017,N_2159,N_2059);
and U3018 (N_3018,N_2237,N_2939);
nor U3019 (N_3019,N_2207,N_2139);
nor U3020 (N_3020,N_2954,N_2378);
nor U3021 (N_3021,N_2201,N_2514);
or U3022 (N_3022,N_2585,N_2229);
nand U3023 (N_3023,N_2163,N_2015);
nand U3024 (N_3024,N_2965,N_2712);
nand U3025 (N_3025,N_2467,N_2307);
and U3026 (N_3026,N_2521,N_2393);
and U3027 (N_3027,N_2036,N_2647);
and U3028 (N_3028,N_2010,N_2335);
or U3029 (N_3029,N_2990,N_2291);
xor U3030 (N_3030,N_2988,N_2331);
nand U3031 (N_3031,N_2102,N_2615);
xor U3032 (N_3032,N_2287,N_2679);
or U3033 (N_3033,N_2725,N_2018);
xnor U3034 (N_3034,N_2786,N_2969);
and U3035 (N_3035,N_2643,N_2011);
or U3036 (N_3036,N_2194,N_2758);
and U3037 (N_3037,N_2596,N_2557);
nor U3038 (N_3038,N_2401,N_2891);
nor U3039 (N_3039,N_2184,N_2410);
xor U3040 (N_3040,N_2633,N_2685);
nand U3041 (N_3041,N_2162,N_2536);
nor U3042 (N_3042,N_2048,N_2802);
or U3043 (N_3043,N_2027,N_2723);
and U3044 (N_3044,N_2610,N_2987);
nor U3045 (N_3045,N_2661,N_2859);
or U3046 (N_3046,N_2628,N_2520);
and U3047 (N_3047,N_2947,N_2456);
and U3048 (N_3048,N_2533,N_2756);
nand U3049 (N_3049,N_2636,N_2471);
or U3050 (N_3050,N_2149,N_2500);
nand U3051 (N_3051,N_2224,N_2871);
nand U3052 (N_3052,N_2659,N_2665);
and U3053 (N_3053,N_2769,N_2840);
nand U3054 (N_3054,N_2733,N_2957);
or U3055 (N_3055,N_2921,N_2885);
or U3056 (N_3056,N_2562,N_2364);
xnor U3057 (N_3057,N_2927,N_2234);
and U3058 (N_3058,N_2826,N_2454);
and U3059 (N_3059,N_2991,N_2470);
xor U3060 (N_3060,N_2645,N_2038);
nand U3061 (N_3061,N_2004,N_2377);
or U3062 (N_3062,N_2369,N_2457);
nand U3063 (N_3063,N_2421,N_2692);
nand U3064 (N_3064,N_2680,N_2602);
nor U3065 (N_3065,N_2126,N_2781);
or U3066 (N_3066,N_2613,N_2641);
nor U3067 (N_3067,N_2134,N_2542);
and U3068 (N_3068,N_2616,N_2075);
and U3069 (N_3069,N_2091,N_2180);
xnor U3070 (N_3070,N_2772,N_2822);
nor U3071 (N_3071,N_2030,N_2831);
nand U3072 (N_3072,N_2812,N_2190);
nand U3073 (N_3073,N_2933,N_2193);
or U3074 (N_3074,N_2972,N_2977);
or U3075 (N_3075,N_2409,N_2848);
and U3076 (N_3076,N_2600,N_2763);
xor U3077 (N_3077,N_2925,N_2583);
or U3078 (N_3078,N_2886,N_2153);
or U3079 (N_3079,N_2687,N_2926);
or U3080 (N_3080,N_2718,N_2223);
xnor U3081 (N_3081,N_2172,N_2061);
and U3082 (N_3082,N_2586,N_2876);
and U3083 (N_3083,N_2941,N_2415);
nand U3084 (N_3084,N_2841,N_2313);
or U3085 (N_3085,N_2762,N_2515);
or U3086 (N_3086,N_2942,N_2380);
nand U3087 (N_3087,N_2423,N_2414);
or U3088 (N_3088,N_2448,N_2254);
and U3089 (N_3089,N_2986,N_2123);
or U3090 (N_3090,N_2654,N_2773);
or U3091 (N_3091,N_2080,N_2870);
nor U3092 (N_3092,N_2098,N_2345);
nand U3093 (N_3093,N_2006,N_2084);
nand U3094 (N_3094,N_2746,N_2671);
and U3095 (N_3095,N_2328,N_2239);
nand U3096 (N_3096,N_2106,N_2706);
or U3097 (N_3097,N_2477,N_2397);
nand U3098 (N_3098,N_2145,N_2069);
nand U3099 (N_3099,N_2753,N_2517);
xnor U3100 (N_3100,N_2131,N_2961);
nor U3101 (N_3101,N_2319,N_2089);
or U3102 (N_3102,N_2649,N_2262);
or U3103 (N_3103,N_2973,N_2785);
nor U3104 (N_3104,N_2386,N_2064);
nand U3105 (N_3105,N_2512,N_2304);
nor U3106 (N_3106,N_2407,N_2581);
and U3107 (N_3107,N_2196,N_2099);
and U3108 (N_3108,N_2593,N_2315);
and U3109 (N_3109,N_2952,N_2399);
or U3110 (N_3110,N_2735,N_2547);
or U3111 (N_3111,N_2868,N_2005);
and U3112 (N_3112,N_2427,N_2998);
nor U3113 (N_3113,N_2571,N_2035);
nor U3114 (N_3114,N_2717,N_2187);
or U3115 (N_3115,N_2323,N_2857);
nor U3116 (N_3116,N_2340,N_2129);
nand U3117 (N_3117,N_2248,N_2627);
nor U3118 (N_3118,N_2700,N_2917);
nor U3119 (N_3119,N_2031,N_2809);
nor U3120 (N_3120,N_2525,N_2049);
or U3121 (N_3121,N_2856,N_2824);
xor U3122 (N_3122,N_2657,N_2865);
nor U3123 (N_3123,N_2016,N_2890);
xor U3124 (N_3124,N_2750,N_2757);
nor U3125 (N_3125,N_2632,N_2160);
nor U3126 (N_3126,N_2853,N_2435);
nand U3127 (N_3127,N_2249,N_2862);
or U3128 (N_3128,N_2481,N_2815);
nand U3129 (N_3129,N_2033,N_2359);
or U3130 (N_3130,N_2041,N_2157);
nand U3131 (N_3131,N_2771,N_2151);
or U3132 (N_3132,N_2598,N_2014);
nand U3133 (N_3133,N_2795,N_2579);
or U3134 (N_3134,N_2424,N_2352);
nand U3135 (N_3135,N_2716,N_2449);
xor U3136 (N_3136,N_2147,N_2710);
and U3137 (N_3137,N_2419,N_2425);
xor U3138 (N_3138,N_2278,N_2541);
xor U3139 (N_3139,N_2836,N_2071);
or U3140 (N_3140,N_2979,N_2827);
xor U3141 (N_3141,N_2243,N_2932);
xnor U3142 (N_3142,N_2357,N_2624);
nor U3143 (N_3143,N_2440,N_2487);
and U3144 (N_3144,N_2852,N_2349);
or U3145 (N_3145,N_2749,N_2165);
nor U3146 (N_3146,N_2776,N_2026);
nor U3147 (N_3147,N_2231,N_2755);
nor U3148 (N_3148,N_2232,N_2971);
nor U3149 (N_3149,N_2945,N_2325);
nor U3150 (N_3150,N_2404,N_2678);
or U3151 (N_3151,N_2247,N_2078);
and U3152 (N_3152,N_2213,N_2204);
xor U3153 (N_3153,N_2850,N_2108);
or U3154 (N_3154,N_2317,N_2400);
xor U3155 (N_3155,N_2726,N_2907);
and U3156 (N_3156,N_2743,N_2416);
and U3157 (N_3157,N_2731,N_2576);
nor U3158 (N_3158,N_2299,N_2902);
and U3159 (N_3159,N_2001,N_2117);
nand U3160 (N_3160,N_2745,N_2518);
nor U3161 (N_3161,N_2334,N_2839);
nand U3162 (N_3162,N_2188,N_2588);
nor U3163 (N_3163,N_2119,N_2691);
xor U3164 (N_3164,N_2601,N_2813);
nor U3165 (N_3165,N_2504,N_2042);
and U3166 (N_3166,N_2553,N_2493);
nor U3167 (N_3167,N_2385,N_2963);
nor U3168 (N_3168,N_2447,N_2931);
or U3169 (N_3169,N_2663,N_2432);
or U3170 (N_3170,N_2483,N_2637);
nand U3171 (N_3171,N_2511,N_2845);
nand U3172 (N_3172,N_2490,N_2582);
and U3173 (N_3173,N_2697,N_2915);
and U3174 (N_3174,N_2185,N_2916);
and U3175 (N_3175,N_2210,N_2312);
and U3176 (N_3176,N_2076,N_2279);
or U3177 (N_3177,N_2173,N_2496);
or U3178 (N_3178,N_2439,N_2854);
or U3179 (N_3179,N_2888,N_2573);
and U3180 (N_3180,N_2810,N_2882);
or U3181 (N_3181,N_2164,N_2684);
and U3182 (N_3182,N_2120,N_2696);
nor U3183 (N_3183,N_2214,N_2079);
and U3184 (N_3184,N_2189,N_2318);
nand U3185 (N_3185,N_2855,N_2460);
and U3186 (N_3186,N_2097,N_2568);
and U3187 (N_3187,N_2689,N_2127);
and U3188 (N_3188,N_2782,N_2801);
nand U3189 (N_3189,N_2115,N_2251);
or U3190 (N_3190,N_2132,N_2630);
xnor U3191 (N_3191,N_2371,N_2740);
or U3192 (N_3192,N_2430,N_2937);
nor U3193 (N_3193,N_2494,N_2192);
or U3194 (N_3194,N_2653,N_2374);
and U3195 (N_3195,N_2730,N_2779);
xor U3196 (N_3196,N_2436,N_2903);
and U3197 (N_3197,N_2395,N_2209);
nand U3198 (N_3198,N_2881,N_2866);
or U3199 (N_3199,N_2221,N_2737);
or U3200 (N_3200,N_2250,N_2474);
xor U3201 (N_3201,N_2113,N_2170);
nor U3202 (N_3202,N_2365,N_2981);
and U3203 (N_3203,N_2580,N_2047);
nor U3204 (N_3204,N_2434,N_2914);
or U3205 (N_3205,N_2354,N_2342);
and U3206 (N_3206,N_2675,N_2202);
or U3207 (N_3207,N_2233,N_2353);
nor U3208 (N_3208,N_2200,N_2732);
and U3209 (N_3209,N_2565,N_2452);
or U3210 (N_3210,N_2936,N_2244);
and U3211 (N_3211,N_2215,N_2245);
nor U3212 (N_3212,N_2887,N_2455);
or U3213 (N_3213,N_2022,N_2056);
nor U3214 (N_3214,N_2955,N_2003);
and U3215 (N_3215,N_2044,N_2253);
nand U3216 (N_3216,N_2333,N_2308);
or U3217 (N_3217,N_2849,N_2721);
or U3218 (N_3218,N_2843,N_2595);
nand U3219 (N_3219,N_2897,N_2282);
xnor U3220 (N_3220,N_2577,N_2607);
xnor U3221 (N_3221,N_2550,N_2505);
or U3222 (N_3222,N_2516,N_2219);
or U3223 (N_3223,N_2818,N_2808);
nor U3224 (N_3224,N_2274,N_2688);
and U3225 (N_3225,N_2842,N_2297);
and U3226 (N_3226,N_2968,N_2922);
and U3227 (N_3227,N_2655,N_2107);
xnor U3228 (N_3228,N_2008,N_2996);
or U3229 (N_3229,N_2437,N_2951);
nor U3230 (N_3230,N_2392,N_2530);
nor U3231 (N_3231,N_2833,N_2337);
nand U3232 (N_3232,N_2208,N_2799);
and U3233 (N_3233,N_2478,N_2154);
nand U3234 (N_3234,N_2584,N_2125);
nor U3235 (N_3235,N_2388,N_2873);
and U3236 (N_3236,N_2513,N_2711);
xnor U3237 (N_3237,N_2362,N_2896);
or U3238 (N_3238,N_2465,N_2567);
nor U3239 (N_3239,N_2350,N_2012);
xnor U3240 (N_3240,N_2908,N_2860);
and U3241 (N_3241,N_2648,N_2570);
nor U3242 (N_3242,N_2442,N_2422);
and U3243 (N_3243,N_2806,N_2555);
nor U3244 (N_3244,N_2072,N_2495);
xor U3245 (N_3245,N_2472,N_2501);
and U3246 (N_3246,N_2976,N_2889);
nand U3247 (N_3247,N_2715,N_2719);
xor U3248 (N_3248,N_2441,N_2905);
and U3249 (N_3249,N_2777,N_2389);
nand U3250 (N_3250,N_2646,N_2956);
or U3251 (N_3251,N_2528,N_2703);
nor U3252 (N_3252,N_2970,N_2285);
nand U3253 (N_3253,N_2043,N_2152);
and U3254 (N_3254,N_2029,N_2713);
and U3255 (N_3255,N_2911,N_2418);
and U3256 (N_3256,N_2928,N_2060);
nand U3257 (N_3257,N_2677,N_2834);
and U3258 (N_3258,N_2024,N_2546);
nor U3259 (N_3259,N_2784,N_2070);
nor U3260 (N_3260,N_2109,N_2742);
and U3261 (N_3261,N_2791,N_2556);
and U3262 (N_3262,N_2166,N_2623);
or U3263 (N_3263,N_2054,N_2321);
and U3264 (N_3264,N_2794,N_2235);
xnor U3265 (N_3265,N_2569,N_2461);
or U3266 (N_3266,N_2087,N_2605);
or U3267 (N_3267,N_2480,N_2114);
and U3268 (N_3268,N_2899,N_2893);
or U3269 (N_3269,N_2199,N_2747);
xor U3270 (N_3270,N_2376,N_2609);
and U3271 (N_3271,N_2445,N_2037);
and U3272 (N_3272,N_2384,N_2240);
nor U3273 (N_3273,N_2062,N_2751);
and U3274 (N_3274,N_2264,N_2290);
or U3275 (N_3275,N_2411,N_2217);
xnor U3276 (N_3276,N_2475,N_2046);
nor U3277 (N_3277,N_2343,N_2174);
or U3278 (N_3278,N_2551,N_2608);
nand U3279 (N_3279,N_2989,N_2666);
xor U3280 (N_3280,N_2629,N_2330);
nor U3281 (N_3281,N_2529,N_2203);
nor U3282 (N_3282,N_2704,N_2499);
or U3283 (N_3283,N_2462,N_2527);
nor U3284 (N_3284,N_2261,N_2363);
nand U3285 (N_3285,N_2817,N_2158);
or U3286 (N_3286,N_2545,N_2708);
and U3287 (N_3287,N_2774,N_2761);
and U3288 (N_3288,N_2695,N_2877);
or U3289 (N_3289,N_2265,N_2997);
and U3290 (N_3290,N_2316,N_2765);
nand U3291 (N_3291,N_2367,N_2993);
and U3292 (N_3292,N_2405,N_2975);
nor U3293 (N_3293,N_2720,N_2398);
xor U3294 (N_3294,N_2104,N_2130);
xor U3295 (N_3295,N_2861,N_2355);
and U3296 (N_3296,N_2760,N_2724);
and U3297 (N_3297,N_2110,N_2532);
xor U3298 (N_3298,N_2566,N_2728);
nor U3299 (N_3299,N_2816,N_2428);
nand U3300 (N_3300,N_2281,N_2590);
nor U3301 (N_3301,N_2182,N_2292);
nor U3302 (N_3302,N_2672,N_2895);
nor U3303 (N_3303,N_2293,N_2348);
nor U3304 (N_3304,N_2694,N_2403);
nor U3305 (N_3305,N_2420,N_2040);
or U3306 (N_3306,N_2216,N_2175);
or U3307 (N_3307,N_2701,N_2631);
nand U3308 (N_3308,N_2266,N_2081);
nand U3309 (N_3309,N_2510,N_2574);
xnor U3310 (N_3310,N_2314,N_2429);
and U3311 (N_3311,N_2994,N_2039);
nand U3312 (N_3312,N_2966,N_2179);
nand U3313 (N_3313,N_2488,N_2055);
nand U3314 (N_3314,N_2358,N_2073);
and U3315 (N_3315,N_2155,N_2057);
and U3316 (N_3316,N_2744,N_2652);
and U3317 (N_3317,N_2883,N_2270);
xor U3318 (N_3318,N_2962,N_2832);
or U3319 (N_3319,N_2273,N_2327);
and U3320 (N_3320,N_2322,N_2148);
nand U3321 (N_3321,N_2978,N_2045);
or U3322 (N_3322,N_2549,N_2181);
or U3323 (N_3323,N_2620,N_2768);
nand U3324 (N_3324,N_2621,N_2116);
nand U3325 (N_3325,N_2787,N_2206);
nor U3326 (N_3326,N_2662,N_2225);
and U3327 (N_3327,N_2009,N_2980);
or U3328 (N_3328,N_2508,N_2468);
nand U3329 (N_3329,N_2382,N_2938);
or U3330 (N_3330,N_2958,N_2919);
xnor U3331 (N_3331,N_2111,N_2366);
and U3332 (N_3332,N_2238,N_2778);
nor U3333 (N_3333,N_2698,N_2667);
or U3334 (N_3334,N_2589,N_2453);
or U3335 (N_3335,N_2092,N_2286);
and U3336 (N_3336,N_2523,N_2417);
or U3337 (N_3337,N_2020,N_2368);
and U3338 (N_3338,N_2544,N_2729);
nor U3339 (N_3339,N_2869,N_2912);
nand U3340 (N_3340,N_2433,N_2985);
and U3341 (N_3341,N_2819,N_2142);
or U3342 (N_3342,N_2141,N_2361);
nand U3343 (N_3343,N_2476,N_2105);
xnor U3344 (N_3344,N_2823,N_2909);
nor U3345 (N_3345,N_2390,N_2485);
nor U3346 (N_3346,N_2880,N_2051);
xor U3347 (N_3347,N_2699,N_2458);
nand U3348 (N_3348,N_2775,N_2095);
nor U3349 (N_3349,N_2614,N_2948);
or U3350 (N_3350,N_2302,N_2268);
or U3351 (N_3351,N_2228,N_2683);
or U3352 (N_3352,N_2300,N_2028);
and U3353 (N_3353,N_2619,N_2186);
and U3354 (N_3354,N_2227,N_2121);
or U3355 (N_3355,N_2575,N_2940);
nand U3356 (N_3356,N_2935,N_2066);
or U3357 (N_3357,N_2792,N_2426);
and U3358 (N_3358,N_2642,N_2197);
nor U3359 (N_3359,N_2288,N_2143);
and U3360 (N_3360,N_2373,N_2846);
and U3361 (N_3361,N_2133,N_2591);
nor U3362 (N_3362,N_2686,N_2707);
nor U3363 (N_3363,N_2884,N_2705);
nor U3364 (N_3364,N_2320,N_2714);
or U3365 (N_3365,N_2934,N_2820);
or U3366 (N_3366,N_2258,N_2920);
nand U3367 (N_3367,N_2329,N_2263);
or U3368 (N_3368,N_2236,N_2289);
nand U3369 (N_3369,N_2738,N_2644);
and U3370 (N_3370,N_2339,N_2053);
or U3371 (N_3371,N_2351,N_2558);
and U3372 (N_3372,N_2086,N_2526);
or U3373 (N_3373,N_2171,N_2807);
and U3374 (N_3374,N_2538,N_2503);
and U3375 (N_3375,N_2379,N_2220);
xnor U3376 (N_3376,N_2112,N_2752);
or U3377 (N_3377,N_2269,N_2176);
or U3378 (N_3378,N_2222,N_2296);
nand U3379 (N_3379,N_2205,N_2984);
or U3380 (N_3380,N_2394,N_2021);
nor U3381 (N_3381,N_2754,N_2198);
or U3382 (N_3382,N_2275,N_2668);
nand U3383 (N_3383,N_2944,N_2497);
nor U3384 (N_3384,N_2611,N_2664);
nand U3385 (N_3385,N_2800,N_2177);
nor U3386 (N_3386,N_2599,N_2587);
nand U3387 (N_3387,N_2543,N_2879);
xnor U3388 (N_3388,N_2077,N_2019);
or U3389 (N_3389,N_2519,N_2492);
or U3390 (N_3390,N_2796,N_2535);
nand U3391 (N_3391,N_2498,N_2995);
nor U3392 (N_3392,N_2068,N_2169);
nand U3393 (N_3393,N_2612,N_2548);
nor U3394 (N_3394,N_2797,N_2858);
nand U3395 (N_3395,N_2676,N_2790);
and U3396 (N_3396,N_2252,N_2242);
xor U3397 (N_3397,N_2058,N_2597);
or U3398 (N_3398,N_2381,N_2878);
xnor U3399 (N_3399,N_2618,N_2682);
nor U3400 (N_3400,N_2502,N_2604);
nand U3401 (N_3401,N_2168,N_2413);
nand U3402 (N_3402,N_2067,N_2391);
and U3403 (N_3403,N_2964,N_2088);
or U3404 (N_3404,N_2847,N_2982);
nand U3405 (N_3405,N_2625,N_2167);
xnor U3406 (N_3406,N_2375,N_2910);
nor U3407 (N_3407,N_2539,N_2780);
or U3408 (N_3408,N_2178,N_2838);
or U3409 (N_3409,N_2992,N_2444);
nand U3410 (N_3410,N_2276,N_2594);
and U3411 (N_3411,N_2128,N_2626);
nor U3412 (N_3412,N_2872,N_2479);
or U3413 (N_3413,N_2930,N_2634);
or U3414 (N_3414,N_2821,N_2974);
or U3415 (N_3415,N_2656,N_2267);
nor U3416 (N_3416,N_2336,N_2867);
or U3417 (N_3417,N_2635,N_2272);
or U3418 (N_3418,N_2875,N_2256);
nand U3419 (N_3419,N_2913,N_2310);
nor U3420 (N_3420,N_2191,N_2999);
nand U3421 (N_3421,N_2759,N_2805);
nand U3422 (N_3422,N_2923,N_2298);
or U3423 (N_3423,N_2767,N_2309);
or U3424 (N_3424,N_2459,N_2804);
and U3425 (N_3425,N_2770,N_2140);
and U3426 (N_3426,N_2690,N_2900);
or U3427 (N_3427,N_2681,N_2793);
or U3428 (N_3428,N_2002,N_2564);
nor U3429 (N_3429,N_2118,N_2898);
nor U3430 (N_3430,N_2617,N_2034);
or U3431 (N_3431,N_2482,N_2943);
nor U3432 (N_3432,N_2894,N_2346);
xnor U3433 (N_3433,N_2814,N_2226);
xor U3434 (N_3434,N_2788,N_2146);
or U3435 (N_3435,N_2450,N_2063);
xnor U3436 (N_3436,N_2183,N_2326);
and U3437 (N_3437,N_2709,N_2837);
and U3438 (N_3438,N_2658,N_2096);
nand U3439 (N_3439,N_2561,N_2013);
or U3440 (N_3440,N_2443,N_2959);
and U3441 (N_3441,N_2484,N_2844);
xor U3442 (N_3442,N_2534,N_2830);
nand U3443 (N_3443,N_2074,N_2829);
nand U3444 (N_3444,N_2195,N_2025);
and U3445 (N_3445,N_2507,N_2101);
and U3446 (N_3446,N_2764,N_2789);
or U3447 (N_3447,N_2603,N_2967);
nor U3448 (N_3448,N_2578,N_2766);
and U3449 (N_3449,N_2100,N_2811);
xnor U3450 (N_3450,N_2135,N_2559);
nor U3451 (N_3451,N_2929,N_2983);
or U3452 (N_3452,N_2103,N_2260);
or U3453 (N_3453,N_2924,N_2408);
and U3454 (N_3454,N_2953,N_2332);
or U3455 (N_3455,N_2835,N_2639);
nand U3456 (N_3456,N_2473,N_2383);
or U3457 (N_3457,N_2257,N_2798);
nand U3458 (N_3458,N_2007,N_2466);
nor U3459 (N_3459,N_2638,N_2065);
and U3460 (N_3460,N_2736,N_2949);
nand U3461 (N_3461,N_2739,N_2651);
and U3462 (N_3462,N_2000,N_2946);
nand U3463 (N_3463,N_2734,N_2825);
or U3464 (N_3464,N_2406,N_2693);
xor U3465 (N_3465,N_2305,N_2640);
and U3466 (N_3466,N_2552,N_2303);
nand U3467 (N_3467,N_2918,N_2402);
or U3468 (N_3468,N_2563,N_2673);
and U3469 (N_3469,N_2230,N_2211);
and U3470 (N_3470,N_2396,N_2560);
nand U3471 (N_3471,N_2506,N_2341);
or U3472 (N_3472,N_2124,N_2572);
nand U3473 (N_3473,N_2023,N_2431);
nor U3474 (N_3474,N_2360,N_2592);
nor U3475 (N_3475,N_2674,N_2531);
or U3476 (N_3476,N_2464,N_2032);
and U3477 (N_3477,N_2622,N_2161);
nor U3478 (N_3478,N_2828,N_2255);
and U3479 (N_3479,N_2509,N_2085);
nand U3480 (N_3480,N_2489,N_2295);
nor U3481 (N_3481,N_2451,N_2017);
nand U3482 (N_3482,N_2387,N_2294);
or U3483 (N_3483,N_2271,N_2259);
or U3484 (N_3484,N_2650,N_2901);
or U3485 (N_3485,N_2246,N_2372);
nand U3486 (N_3486,N_2052,N_2136);
or U3487 (N_3487,N_2138,N_2344);
or U3488 (N_3488,N_2311,N_2083);
and U3489 (N_3489,N_2122,N_2904);
or U3490 (N_3490,N_2347,N_2090);
nand U3491 (N_3491,N_2702,N_2241);
or U3492 (N_3492,N_2540,N_2050);
or U3493 (N_3493,N_2874,N_2606);
xnor U3494 (N_3494,N_2670,N_2218);
nor U3495 (N_3495,N_2438,N_2783);
nor U3496 (N_3496,N_2851,N_2284);
nand U3497 (N_3497,N_2283,N_2863);
nor U3498 (N_3498,N_2463,N_2338);
or U3499 (N_3499,N_2554,N_2960);
or U3500 (N_3500,N_2776,N_2581);
nand U3501 (N_3501,N_2596,N_2612);
xnor U3502 (N_3502,N_2326,N_2517);
nor U3503 (N_3503,N_2063,N_2214);
xnor U3504 (N_3504,N_2779,N_2786);
or U3505 (N_3505,N_2961,N_2598);
and U3506 (N_3506,N_2991,N_2205);
and U3507 (N_3507,N_2183,N_2874);
and U3508 (N_3508,N_2653,N_2040);
nor U3509 (N_3509,N_2919,N_2647);
nand U3510 (N_3510,N_2910,N_2605);
or U3511 (N_3511,N_2187,N_2002);
xor U3512 (N_3512,N_2270,N_2317);
nor U3513 (N_3513,N_2964,N_2604);
and U3514 (N_3514,N_2499,N_2228);
or U3515 (N_3515,N_2275,N_2904);
nor U3516 (N_3516,N_2143,N_2944);
and U3517 (N_3517,N_2413,N_2641);
or U3518 (N_3518,N_2236,N_2479);
nor U3519 (N_3519,N_2206,N_2528);
nand U3520 (N_3520,N_2495,N_2733);
or U3521 (N_3521,N_2768,N_2152);
xor U3522 (N_3522,N_2320,N_2865);
or U3523 (N_3523,N_2221,N_2573);
nand U3524 (N_3524,N_2899,N_2573);
and U3525 (N_3525,N_2803,N_2706);
and U3526 (N_3526,N_2232,N_2797);
nor U3527 (N_3527,N_2036,N_2886);
xor U3528 (N_3528,N_2129,N_2695);
and U3529 (N_3529,N_2858,N_2630);
nand U3530 (N_3530,N_2291,N_2436);
nand U3531 (N_3531,N_2729,N_2522);
nand U3532 (N_3532,N_2948,N_2157);
nand U3533 (N_3533,N_2543,N_2387);
and U3534 (N_3534,N_2023,N_2110);
nor U3535 (N_3535,N_2837,N_2398);
nor U3536 (N_3536,N_2129,N_2354);
and U3537 (N_3537,N_2364,N_2438);
or U3538 (N_3538,N_2528,N_2125);
nor U3539 (N_3539,N_2657,N_2936);
nor U3540 (N_3540,N_2182,N_2554);
nand U3541 (N_3541,N_2018,N_2785);
nor U3542 (N_3542,N_2040,N_2730);
nor U3543 (N_3543,N_2617,N_2326);
and U3544 (N_3544,N_2017,N_2720);
or U3545 (N_3545,N_2408,N_2360);
xnor U3546 (N_3546,N_2438,N_2827);
and U3547 (N_3547,N_2285,N_2476);
nand U3548 (N_3548,N_2848,N_2323);
or U3549 (N_3549,N_2267,N_2071);
nor U3550 (N_3550,N_2643,N_2705);
or U3551 (N_3551,N_2125,N_2424);
nor U3552 (N_3552,N_2095,N_2620);
or U3553 (N_3553,N_2940,N_2932);
nand U3554 (N_3554,N_2312,N_2518);
nand U3555 (N_3555,N_2925,N_2956);
nand U3556 (N_3556,N_2541,N_2114);
or U3557 (N_3557,N_2490,N_2273);
nand U3558 (N_3558,N_2756,N_2243);
and U3559 (N_3559,N_2237,N_2716);
nor U3560 (N_3560,N_2993,N_2291);
nand U3561 (N_3561,N_2137,N_2091);
nor U3562 (N_3562,N_2990,N_2147);
or U3563 (N_3563,N_2833,N_2960);
nor U3564 (N_3564,N_2026,N_2596);
nor U3565 (N_3565,N_2491,N_2558);
or U3566 (N_3566,N_2837,N_2979);
nor U3567 (N_3567,N_2193,N_2534);
xnor U3568 (N_3568,N_2840,N_2316);
xnor U3569 (N_3569,N_2795,N_2393);
nor U3570 (N_3570,N_2740,N_2261);
nor U3571 (N_3571,N_2481,N_2966);
nand U3572 (N_3572,N_2162,N_2926);
nand U3573 (N_3573,N_2329,N_2631);
nand U3574 (N_3574,N_2045,N_2604);
or U3575 (N_3575,N_2351,N_2836);
and U3576 (N_3576,N_2916,N_2229);
nand U3577 (N_3577,N_2435,N_2930);
xnor U3578 (N_3578,N_2661,N_2418);
nand U3579 (N_3579,N_2312,N_2542);
or U3580 (N_3580,N_2071,N_2494);
and U3581 (N_3581,N_2000,N_2957);
nand U3582 (N_3582,N_2275,N_2156);
nand U3583 (N_3583,N_2096,N_2128);
nand U3584 (N_3584,N_2622,N_2092);
or U3585 (N_3585,N_2077,N_2051);
nor U3586 (N_3586,N_2837,N_2944);
nor U3587 (N_3587,N_2502,N_2377);
or U3588 (N_3588,N_2516,N_2218);
or U3589 (N_3589,N_2598,N_2829);
and U3590 (N_3590,N_2523,N_2286);
nor U3591 (N_3591,N_2440,N_2653);
or U3592 (N_3592,N_2085,N_2272);
and U3593 (N_3593,N_2428,N_2576);
or U3594 (N_3594,N_2093,N_2878);
or U3595 (N_3595,N_2693,N_2808);
and U3596 (N_3596,N_2485,N_2620);
xnor U3597 (N_3597,N_2794,N_2096);
nor U3598 (N_3598,N_2512,N_2379);
nand U3599 (N_3599,N_2745,N_2102);
nand U3600 (N_3600,N_2456,N_2855);
or U3601 (N_3601,N_2860,N_2986);
or U3602 (N_3602,N_2463,N_2265);
nand U3603 (N_3603,N_2888,N_2222);
nand U3604 (N_3604,N_2411,N_2761);
nor U3605 (N_3605,N_2006,N_2033);
nand U3606 (N_3606,N_2875,N_2476);
or U3607 (N_3607,N_2408,N_2338);
and U3608 (N_3608,N_2305,N_2327);
nor U3609 (N_3609,N_2184,N_2256);
nand U3610 (N_3610,N_2199,N_2443);
nor U3611 (N_3611,N_2771,N_2533);
xor U3612 (N_3612,N_2767,N_2406);
nand U3613 (N_3613,N_2811,N_2415);
nor U3614 (N_3614,N_2434,N_2246);
xor U3615 (N_3615,N_2013,N_2744);
or U3616 (N_3616,N_2122,N_2352);
nand U3617 (N_3617,N_2503,N_2534);
or U3618 (N_3618,N_2157,N_2047);
or U3619 (N_3619,N_2559,N_2306);
or U3620 (N_3620,N_2278,N_2513);
nor U3621 (N_3621,N_2003,N_2378);
xor U3622 (N_3622,N_2209,N_2580);
nand U3623 (N_3623,N_2479,N_2488);
nor U3624 (N_3624,N_2353,N_2996);
or U3625 (N_3625,N_2584,N_2224);
nand U3626 (N_3626,N_2563,N_2976);
and U3627 (N_3627,N_2524,N_2090);
or U3628 (N_3628,N_2366,N_2032);
and U3629 (N_3629,N_2245,N_2980);
nor U3630 (N_3630,N_2057,N_2537);
and U3631 (N_3631,N_2181,N_2090);
and U3632 (N_3632,N_2356,N_2645);
or U3633 (N_3633,N_2534,N_2935);
nor U3634 (N_3634,N_2660,N_2882);
nand U3635 (N_3635,N_2189,N_2630);
and U3636 (N_3636,N_2093,N_2405);
and U3637 (N_3637,N_2435,N_2171);
and U3638 (N_3638,N_2572,N_2654);
nor U3639 (N_3639,N_2195,N_2671);
nor U3640 (N_3640,N_2884,N_2416);
xnor U3641 (N_3641,N_2757,N_2114);
and U3642 (N_3642,N_2629,N_2129);
nand U3643 (N_3643,N_2867,N_2335);
nor U3644 (N_3644,N_2678,N_2324);
nor U3645 (N_3645,N_2869,N_2528);
nand U3646 (N_3646,N_2866,N_2343);
nand U3647 (N_3647,N_2098,N_2879);
nand U3648 (N_3648,N_2951,N_2242);
or U3649 (N_3649,N_2312,N_2228);
nand U3650 (N_3650,N_2950,N_2942);
and U3651 (N_3651,N_2148,N_2229);
and U3652 (N_3652,N_2812,N_2492);
or U3653 (N_3653,N_2517,N_2461);
nand U3654 (N_3654,N_2686,N_2430);
and U3655 (N_3655,N_2838,N_2101);
nand U3656 (N_3656,N_2938,N_2083);
and U3657 (N_3657,N_2639,N_2203);
nor U3658 (N_3658,N_2426,N_2014);
and U3659 (N_3659,N_2429,N_2558);
nor U3660 (N_3660,N_2538,N_2062);
nor U3661 (N_3661,N_2657,N_2808);
and U3662 (N_3662,N_2788,N_2977);
and U3663 (N_3663,N_2658,N_2478);
and U3664 (N_3664,N_2222,N_2119);
xnor U3665 (N_3665,N_2123,N_2295);
xnor U3666 (N_3666,N_2798,N_2442);
or U3667 (N_3667,N_2013,N_2206);
or U3668 (N_3668,N_2726,N_2822);
or U3669 (N_3669,N_2693,N_2583);
and U3670 (N_3670,N_2879,N_2041);
nor U3671 (N_3671,N_2666,N_2098);
nor U3672 (N_3672,N_2772,N_2454);
nand U3673 (N_3673,N_2769,N_2143);
nand U3674 (N_3674,N_2238,N_2783);
nor U3675 (N_3675,N_2543,N_2348);
nand U3676 (N_3676,N_2466,N_2464);
nand U3677 (N_3677,N_2827,N_2588);
and U3678 (N_3678,N_2196,N_2077);
nor U3679 (N_3679,N_2638,N_2665);
nor U3680 (N_3680,N_2020,N_2114);
xor U3681 (N_3681,N_2569,N_2965);
and U3682 (N_3682,N_2052,N_2043);
or U3683 (N_3683,N_2513,N_2862);
nor U3684 (N_3684,N_2967,N_2477);
nand U3685 (N_3685,N_2558,N_2983);
nand U3686 (N_3686,N_2527,N_2360);
or U3687 (N_3687,N_2671,N_2531);
nor U3688 (N_3688,N_2750,N_2251);
xor U3689 (N_3689,N_2496,N_2936);
and U3690 (N_3690,N_2000,N_2157);
nand U3691 (N_3691,N_2637,N_2776);
xor U3692 (N_3692,N_2894,N_2146);
or U3693 (N_3693,N_2041,N_2099);
and U3694 (N_3694,N_2188,N_2493);
nand U3695 (N_3695,N_2707,N_2773);
nor U3696 (N_3696,N_2747,N_2115);
nand U3697 (N_3697,N_2847,N_2382);
nor U3698 (N_3698,N_2200,N_2343);
nor U3699 (N_3699,N_2803,N_2289);
nand U3700 (N_3700,N_2492,N_2296);
nor U3701 (N_3701,N_2300,N_2263);
nor U3702 (N_3702,N_2756,N_2126);
and U3703 (N_3703,N_2618,N_2335);
or U3704 (N_3704,N_2815,N_2762);
and U3705 (N_3705,N_2479,N_2077);
nor U3706 (N_3706,N_2492,N_2715);
and U3707 (N_3707,N_2318,N_2274);
nand U3708 (N_3708,N_2120,N_2683);
nor U3709 (N_3709,N_2388,N_2346);
xnor U3710 (N_3710,N_2499,N_2180);
or U3711 (N_3711,N_2538,N_2246);
nor U3712 (N_3712,N_2060,N_2212);
nor U3713 (N_3713,N_2018,N_2569);
and U3714 (N_3714,N_2087,N_2366);
nor U3715 (N_3715,N_2253,N_2295);
nand U3716 (N_3716,N_2552,N_2114);
or U3717 (N_3717,N_2492,N_2379);
xor U3718 (N_3718,N_2508,N_2697);
xnor U3719 (N_3719,N_2430,N_2744);
and U3720 (N_3720,N_2033,N_2510);
and U3721 (N_3721,N_2962,N_2107);
xnor U3722 (N_3722,N_2492,N_2989);
nor U3723 (N_3723,N_2923,N_2690);
nand U3724 (N_3724,N_2524,N_2768);
nand U3725 (N_3725,N_2909,N_2878);
and U3726 (N_3726,N_2673,N_2748);
and U3727 (N_3727,N_2798,N_2477);
and U3728 (N_3728,N_2197,N_2604);
nand U3729 (N_3729,N_2552,N_2365);
or U3730 (N_3730,N_2225,N_2529);
or U3731 (N_3731,N_2940,N_2356);
nor U3732 (N_3732,N_2112,N_2554);
nand U3733 (N_3733,N_2779,N_2793);
xor U3734 (N_3734,N_2576,N_2772);
xnor U3735 (N_3735,N_2621,N_2703);
nor U3736 (N_3736,N_2167,N_2386);
nand U3737 (N_3737,N_2017,N_2581);
and U3738 (N_3738,N_2459,N_2719);
and U3739 (N_3739,N_2582,N_2304);
xnor U3740 (N_3740,N_2364,N_2088);
nand U3741 (N_3741,N_2358,N_2158);
and U3742 (N_3742,N_2712,N_2419);
xnor U3743 (N_3743,N_2779,N_2002);
or U3744 (N_3744,N_2209,N_2315);
or U3745 (N_3745,N_2060,N_2967);
nor U3746 (N_3746,N_2411,N_2421);
and U3747 (N_3747,N_2537,N_2315);
or U3748 (N_3748,N_2085,N_2923);
nand U3749 (N_3749,N_2561,N_2706);
xor U3750 (N_3750,N_2400,N_2326);
or U3751 (N_3751,N_2965,N_2120);
nand U3752 (N_3752,N_2710,N_2369);
xnor U3753 (N_3753,N_2102,N_2646);
and U3754 (N_3754,N_2247,N_2982);
and U3755 (N_3755,N_2885,N_2304);
and U3756 (N_3756,N_2659,N_2126);
nand U3757 (N_3757,N_2333,N_2964);
or U3758 (N_3758,N_2387,N_2596);
and U3759 (N_3759,N_2086,N_2193);
and U3760 (N_3760,N_2794,N_2319);
or U3761 (N_3761,N_2971,N_2427);
nor U3762 (N_3762,N_2626,N_2865);
xor U3763 (N_3763,N_2224,N_2637);
nand U3764 (N_3764,N_2290,N_2233);
nor U3765 (N_3765,N_2196,N_2805);
nor U3766 (N_3766,N_2185,N_2536);
or U3767 (N_3767,N_2994,N_2091);
nand U3768 (N_3768,N_2733,N_2714);
nand U3769 (N_3769,N_2533,N_2820);
and U3770 (N_3770,N_2479,N_2870);
xnor U3771 (N_3771,N_2210,N_2696);
nor U3772 (N_3772,N_2846,N_2489);
nor U3773 (N_3773,N_2809,N_2849);
xnor U3774 (N_3774,N_2615,N_2642);
nand U3775 (N_3775,N_2747,N_2136);
or U3776 (N_3776,N_2727,N_2142);
nor U3777 (N_3777,N_2264,N_2352);
or U3778 (N_3778,N_2293,N_2776);
and U3779 (N_3779,N_2099,N_2573);
and U3780 (N_3780,N_2266,N_2672);
nor U3781 (N_3781,N_2498,N_2724);
nor U3782 (N_3782,N_2944,N_2221);
nand U3783 (N_3783,N_2955,N_2855);
xor U3784 (N_3784,N_2051,N_2418);
and U3785 (N_3785,N_2119,N_2137);
and U3786 (N_3786,N_2100,N_2000);
nor U3787 (N_3787,N_2944,N_2923);
nand U3788 (N_3788,N_2599,N_2882);
or U3789 (N_3789,N_2722,N_2178);
nor U3790 (N_3790,N_2971,N_2612);
or U3791 (N_3791,N_2950,N_2766);
or U3792 (N_3792,N_2245,N_2254);
nor U3793 (N_3793,N_2232,N_2888);
nor U3794 (N_3794,N_2365,N_2727);
and U3795 (N_3795,N_2831,N_2822);
and U3796 (N_3796,N_2344,N_2122);
or U3797 (N_3797,N_2274,N_2545);
and U3798 (N_3798,N_2691,N_2296);
nor U3799 (N_3799,N_2679,N_2499);
nor U3800 (N_3800,N_2282,N_2757);
or U3801 (N_3801,N_2395,N_2587);
xor U3802 (N_3802,N_2086,N_2575);
nor U3803 (N_3803,N_2373,N_2843);
or U3804 (N_3804,N_2599,N_2217);
or U3805 (N_3805,N_2476,N_2094);
and U3806 (N_3806,N_2838,N_2443);
nor U3807 (N_3807,N_2506,N_2520);
xnor U3808 (N_3808,N_2815,N_2016);
nor U3809 (N_3809,N_2615,N_2921);
nor U3810 (N_3810,N_2064,N_2090);
or U3811 (N_3811,N_2980,N_2772);
nand U3812 (N_3812,N_2516,N_2498);
nand U3813 (N_3813,N_2374,N_2137);
nand U3814 (N_3814,N_2940,N_2059);
nand U3815 (N_3815,N_2173,N_2120);
or U3816 (N_3816,N_2748,N_2944);
xnor U3817 (N_3817,N_2245,N_2048);
xor U3818 (N_3818,N_2891,N_2500);
or U3819 (N_3819,N_2530,N_2279);
xnor U3820 (N_3820,N_2761,N_2858);
and U3821 (N_3821,N_2893,N_2576);
and U3822 (N_3822,N_2202,N_2661);
xor U3823 (N_3823,N_2772,N_2059);
or U3824 (N_3824,N_2247,N_2330);
nor U3825 (N_3825,N_2735,N_2497);
nor U3826 (N_3826,N_2912,N_2652);
and U3827 (N_3827,N_2074,N_2683);
nand U3828 (N_3828,N_2374,N_2288);
and U3829 (N_3829,N_2148,N_2061);
and U3830 (N_3830,N_2138,N_2763);
nor U3831 (N_3831,N_2281,N_2060);
nor U3832 (N_3832,N_2277,N_2788);
nand U3833 (N_3833,N_2986,N_2238);
xnor U3834 (N_3834,N_2942,N_2250);
xor U3835 (N_3835,N_2434,N_2589);
nor U3836 (N_3836,N_2238,N_2386);
or U3837 (N_3837,N_2641,N_2146);
and U3838 (N_3838,N_2125,N_2987);
or U3839 (N_3839,N_2987,N_2381);
or U3840 (N_3840,N_2962,N_2994);
nand U3841 (N_3841,N_2693,N_2266);
nand U3842 (N_3842,N_2926,N_2930);
nor U3843 (N_3843,N_2060,N_2500);
or U3844 (N_3844,N_2179,N_2304);
nand U3845 (N_3845,N_2230,N_2875);
or U3846 (N_3846,N_2758,N_2954);
and U3847 (N_3847,N_2151,N_2301);
nor U3848 (N_3848,N_2407,N_2814);
nor U3849 (N_3849,N_2329,N_2673);
and U3850 (N_3850,N_2070,N_2825);
nand U3851 (N_3851,N_2221,N_2617);
or U3852 (N_3852,N_2421,N_2076);
nand U3853 (N_3853,N_2219,N_2276);
and U3854 (N_3854,N_2008,N_2782);
or U3855 (N_3855,N_2404,N_2939);
nor U3856 (N_3856,N_2408,N_2376);
nor U3857 (N_3857,N_2951,N_2469);
nand U3858 (N_3858,N_2760,N_2617);
and U3859 (N_3859,N_2348,N_2418);
xor U3860 (N_3860,N_2082,N_2574);
nand U3861 (N_3861,N_2666,N_2200);
or U3862 (N_3862,N_2867,N_2826);
or U3863 (N_3863,N_2535,N_2556);
nand U3864 (N_3864,N_2824,N_2210);
or U3865 (N_3865,N_2749,N_2287);
nand U3866 (N_3866,N_2548,N_2660);
nor U3867 (N_3867,N_2290,N_2662);
xor U3868 (N_3868,N_2363,N_2839);
nand U3869 (N_3869,N_2270,N_2204);
or U3870 (N_3870,N_2638,N_2871);
nor U3871 (N_3871,N_2184,N_2650);
nand U3872 (N_3872,N_2575,N_2529);
nor U3873 (N_3873,N_2361,N_2924);
nor U3874 (N_3874,N_2933,N_2432);
nand U3875 (N_3875,N_2448,N_2641);
or U3876 (N_3876,N_2525,N_2543);
nand U3877 (N_3877,N_2938,N_2429);
or U3878 (N_3878,N_2901,N_2021);
nor U3879 (N_3879,N_2364,N_2246);
nor U3880 (N_3880,N_2277,N_2818);
nor U3881 (N_3881,N_2734,N_2472);
xnor U3882 (N_3882,N_2556,N_2823);
or U3883 (N_3883,N_2216,N_2599);
nor U3884 (N_3884,N_2537,N_2143);
and U3885 (N_3885,N_2627,N_2625);
nand U3886 (N_3886,N_2195,N_2372);
and U3887 (N_3887,N_2547,N_2734);
or U3888 (N_3888,N_2716,N_2639);
xnor U3889 (N_3889,N_2545,N_2655);
and U3890 (N_3890,N_2127,N_2012);
or U3891 (N_3891,N_2671,N_2003);
and U3892 (N_3892,N_2002,N_2647);
nand U3893 (N_3893,N_2633,N_2056);
nand U3894 (N_3894,N_2018,N_2907);
and U3895 (N_3895,N_2825,N_2952);
or U3896 (N_3896,N_2866,N_2941);
xnor U3897 (N_3897,N_2377,N_2403);
nor U3898 (N_3898,N_2654,N_2401);
nand U3899 (N_3899,N_2645,N_2702);
or U3900 (N_3900,N_2001,N_2287);
nor U3901 (N_3901,N_2698,N_2680);
nand U3902 (N_3902,N_2068,N_2676);
or U3903 (N_3903,N_2225,N_2950);
or U3904 (N_3904,N_2243,N_2334);
nor U3905 (N_3905,N_2943,N_2199);
nand U3906 (N_3906,N_2335,N_2912);
and U3907 (N_3907,N_2738,N_2837);
nor U3908 (N_3908,N_2207,N_2918);
and U3909 (N_3909,N_2529,N_2377);
nor U3910 (N_3910,N_2684,N_2592);
or U3911 (N_3911,N_2839,N_2543);
or U3912 (N_3912,N_2456,N_2490);
or U3913 (N_3913,N_2457,N_2994);
and U3914 (N_3914,N_2672,N_2362);
nand U3915 (N_3915,N_2478,N_2970);
xor U3916 (N_3916,N_2549,N_2988);
nand U3917 (N_3917,N_2503,N_2826);
nand U3918 (N_3918,N_2663,N_2270);
nor U3919 (N_3919,N_2692,N_2651);
nor U3920 (N_3920,N_2580,N_2422);
nand U3921 (N_3921,N_2163,N_2980);
xnor U3922 (N_3922,N_2090,N_2926);
or U3923 (N_3923,N_2672,N_2052);
nor U3924 (N_3924,N_2069,N_2304);
or U3925 (N_3925,N_2906,N_2068);
xor U3926 (N_3926,N_2374,N_2822);
or U3927 (N_3927,N_2417,N_2477);
and U3928 (N_3928,N_2614,N_2161);
nand U3929 (N_3929,N_2787,N_2507);
nor U3930 (N_3930,N_2387,N_2070);
and U3931 (N_3931,N_2678,N_2812);
and U3932 (N_3932,N_2490,N_2043);
or U3933 (N_3933,N_2503,N_2913);
and U3934 (N_3934,N_2032,N_2147);
nor U3935 (N_3935,N_2648,N_2934);
nor U3936 (N_3936,N_2157,N_2232);
or U3937 (N_3937,N_2946,N_2999);
xnor U3938 (N_3938,N_2460,N_2291);
nor U3939 (N_3939,N_2061,N_2062);
or U3940 (N_3940,N_2206,N_2282);
and U3941 (N_3941,N_2560,N_2399);
nor U3942 (N_3942,N_2133,N_2845);
nor U3943 (N_3943,N_2822,N_2817);
nand U3944 (N_3944,N_2441,N_2655);
and U3945 (N_3945,N_2389,N_2634);
nand U3946 (N_3946,N_2323,N_2901);
nand U3947 (N_3947,N_2258,N_2752);
nor U3948 (N_3948,N_2474,N_2258);
nand U3949 (N_3949,N_2436,N_2360);
and U3950 (N_3950,N_2798,N_2260);
nand U3951 (N_3951,N_2573,N_2746);
or U3952 (N_3952,N_2784,N_2367);
nor U3953 (N_3953,N_2760,N_2926);
nor U3954 (N_3954,N_2496,N_2473);
nand U3955 (N_3955,N_2541,N_2951);
nand U3956 (N_3956,N_2862,N_2003);
xnor U3957 (N_3957,N_2312,N_2583);
xnor U3958 (N_3958,N_2520,N_2494);
or U3959 (N_3959,N_2646,N_2112);
or U3960 (N_3960,N_2822,N_2531);
nor U3961 (N_3961,N_2531,N_2512);
nand U3962 (N_3962,N_2614,N_2650);
and U3963 (N_3963,N_2295,N_2833);
or U3964 (N_3964,N_2495,N_2679);
xnor U3965 (N_3965,N_2520,N_2933);
nand U3966 (N_3966,N_2022,N_2874);
or U3967 (N_3967,N_2472,N_2838);
or U3968 (N_3968,N_2122,N_2584);
nor U3969 (N_3969,N_2542,N_2751);
nor U3970 (N_3970,N_2339,N_2747);
xor U3971 (N_3971,N_2330,N_2131);
xor U3972 (N_3972,N_2813,N_2579);
or U3973 (N_3973,N_2095,N_2600);
or U3974 (N_3974,N_2530,N_2865);
xor U3975 (N_3975,N_2412,N_2954);
nor U3976 (N_3976,N_2185,N_2939);
or U3977 (N_3977,N_2261,N_2512);
or U3978 (N_3978,N_2618,N_2697);
and U3979 (N_3979,N_2697,N_2962);
nand U3980 (N_3980,N_2932,N_2682);
or U3981 (N_3981,N_2091,N_2902);
nand U3982 (N_3982,N_2070,N_2179);
and U3983 (N_3983,N_2217,N_2886);
nand U3984 (N_3984,N_2338,N_2803);
nand U3985 (N_3985,N_2921,N_2937);
or U3986 (N_3986,N_2311,N_2112);
nor U3987 (N_3987,N_2755,N_2858);
nand U3988 (N_3988,N_2083,N_2186);
nor U3989 (N_3989,N_2693,N_2632);
and U3990 (N_3990,N_2166,N_2981);
or U3991 (N_3991,N_2572,N_2412);
nand U3992 (N_3992,N_2129,N_2776);
nand U3993 (N_3993,N_2819,N_2330);
and U3994 (N_3994,N_2439,N_2324);
or U3995 (N_3995,N_2460,N_2902);
nand U3996 (N_3996,N_2309,N_2488);
nand U3997 (N_3997,N_2489,N_2443);
and U3998 (N_3998,N_2908,N_2777);
nor U3999 (N_3999,N_2456,N_2749);
nor U4000 (N_4000,N_3442,N_3473);
nand U4001 (N_4001,N_3106,N_3949);
and U4002 (N_4002,N_3320,N_3109);
nand U4003 (N_4003,N_3686,N_3034);
and U4004 (N_4004,N_3703,N_3646);
and U4005 (N_4005,N_3950,N_3581);
xnor U4006 (N_4006,N_3188,N_3823);
xnor U4007 (N_4007,N_3710,N_3381);
nand U4008 (N_4008,N_3286,N_3216);
nor U4009 (N_4009,N_3443,N_3709);
nor U4010 (N_4010,N_3358,N_3923);
nand U4011 (N_4011,N_3400,N_3053);
nand U4012 (N_4012,N_3002,N_3575);
and U4013 (N_4013,N_3343,N_3087);
or U4014 (N_4014,N_3127,N_3198);
or U4015 (N_4015,N_3839,N_3677);
or U4016 (N_4016,N_3678,N_3071);
nor U4017 (N_4017,N_3281,N_3701);
nor U4018 (N_4018,N_3972,N_3757);
or U4019 (N_4019,N_3321,N_3656);
nand U4020 (N_4020,N_3328,N_3136);
nor U4021 (N_4021,N_3290,N_3333);
nand U4022 (N_4022,N_3612,N_3593);
xnor U4023 (N_4023,N_3821,N_3461);
xnor U4024 (N_4024,N_3687,N_3205);
and U4025 (N_4025,N_3438,N_3012);
nand U4026 (N_4026,N_3406,N_3111);
nand U4027 (N_4027,N_3984,N_3768);
nand U4028 (N_4028,N_3148,N_3896);
and U4029 (N_4029,N_3526,N_3561);
and U4030 (N_4030,N_3669,N_3805);
nand U4031 (N_4031,N_3201,N_3969);
nor U4032 (N_4032,N_3022,N_3624);
or U4033 (N_4033,N_3738,N_3857);
and U4034 (N_4034,N_3781,N_3184);
xnor U4035 (N_4035,N_3001,N_3737);
nand U4036 (N_4036,N_3691,N_3030);
or U4037 (N_4037,N_3342,N_3484);
or U4038 (N_4038,N_3700,N_3415);
nand U4039 (N_4039,N_3660,N_3636);
or U4040 (N_4040,N_3579,N_3200);
and U4041 (N_4041,N_3645,N_3414);
nand U4042 (N_4042,N_3763,N_3297);
nor U4043 (N_4043,N_3684,N_3621);
or U4044 (N_4044,N_3331,N_3867);
xnor U4045 (N_4045,N_3880,N_3661);
and U4046 (N_4046,N_3471,N_3982);
xnor U4047 (N_4047,N_3528,N_3132);
nand U4048 (N_4048,N_3427,N_3514);
nor U4049 (N_4049,N_3971,N_3488);
and U4050 (N_4050,N_3441,N_3147);
or U4051 (N_4051,N_3954,N_3233);
nand U4052 (N_4052,N_3634,N_3827);
nand U4053 (N_4053,N_3329,N_3498);
or U4054 (N_4054,N_3830,N_3919);
or U4055 (N_4055,N_3892,N_3614);
and U4056 (N_4056,N_3081,N_3855);
or U4057 (N_4057,N_3067,N_3435);
nor U4058 (N_4058,N_3878,N_3596);
and U4059 (N_4059,N_3074,N_3274);
or U4060 (N_4060,N_3393,N_3941);
nand U4061 (N_4061,N_3631,N_3327);
and U4062 (N_4062,N_3080,N_3772);
nor U4063 (N_4063,N_3815,N_3480);
nand U4064 (N_4064,N_3503,N_3576);
or U4065 (N_4065,N_3792,N_3760);
nand U4066 (N_4066,N_3913,N_3103);
xor U4067 (N_4067,N_3440,N_3856);
nand U4068 (N_4068,N_3428,N_3330);
nand U4069 (N_4069,N_3886,N_3871);
nand U4070 (N_4070,N_3016,N_3762);
and U4071 (N_4071,N_3072,N_3653);
or U4072 (N_4072,N_3448,N_3311);
and U4073 (N_4073,N_3552,N_3719);
xnor U4074 (N_4074,N_3953,N_3056);
nor U4075 (N_4075,N_3199,N_3625);
nand U4076 (N_4076,N_3387,N_3345);
nor U4077 (N_4077,N_3996,N_3234);
or U4078 (N_4078,N_3603,N_3287);
xnor U4079 (N_4079,N_3325,N_3549);
and U4080 (N_4080,N_3690,N_3938);
nor U4081 (N_4081,N_3567,N_3492);
nor U4082 (N_4082,N_3064,N_3644);
nand U4083 (N_4083,N_3726,N_3041);
nor U4084 (N_4084,N_3899,N_3613);
or U4085 (N_4085,N_3648,N_3024);
nand U4086 (N_4086,N_3209,N_3778);
nand U4087 (N_4087,N_3776,N_3332);
xor U4088 (N_4088,N_3957,N_3883);
nand U4089 (N_4089,N_3229,N_3992);
or U4090 (N_4090,N_3548,N_3456);
nor U4091 (N_4091,N_3800,N_3693);
and U4092 (N_4092,N_3202,N_3521);
nand U4093 (N_4093,N_3974,N_3812);
nand U4094 (N_4094,N_3591,N_3252);
or U4095 (N_4095,N_3091,N_3215);
and U4096 (N_4096,N_3973,N_3824);
nand U4097 (N_4097,N_3918,N_3172);
or U4098 (N_4098,N_3247,N_3110);
nand U4099 (N_4099,N_3152,N_3657);
or U4100 (N_4100,N_3866,N_3518);
nor U4101 (N_4101,N_3217,N_3970);
or U4102 (N_4102,N_3711,N_3566);
nor U4103 (N_4103,N_3031,N_3910);
xnor U4104 (N_4104,N_3154,N_3500);
nor U4105 (N_4105,N_3997,N_3529);
or U4106 (N_4106,N_3742,N_3003);
nor U4107 (N_4107,N_3294,N_3512);
nand U4108 (N_4108,N_3336,N_3846);
nand U4109 (N_4109,N_3135,N_3707);
or U4110 (N_4110,N_3039,N_3679);
and U4111 (N_4111,N_3494,N_3164);
or U4112 (N_4112,N_3683,N_3338);
nand U4113 (N_4113,N_3043,N_3813);
nor U4114 (N_4114,N_3520,N_3817);
nor U4115 (N_4115,N_3370,N_3635);
nor U4116 (N_4116,N_3902,N_3452);
nor U4117 (N_4117,N_3623,N_3755);
and U4118 (N_4118,N_3680,N_3782);
nand U4119 (N_4119,N_3582,N_3479);
or U4120 (N_4120,N_3218,N_3079);
xnor U4121 (N_4121,N_3809,N_3238);
and U4122 (N_4122,N_3371,N_3227);
or U4123 (N_4123,N_3667,N_3725);
xnor U4124 (N_4124,N_3605,N_3951);
nand U4125 (N_4125,N_3573,N_3875);
nand U4126 (N_4126,N_3570,N_3303);
and U4127 (N_4127,N_3754,N_3354);
nand U4128 (N_4128,N_3751,N_3788);
and U4129 (N_4129,N_3253,N_3716);
or U4130 (N_4130,N_3681,N_3543);
nor U4131 (N_4131,N_3270,N_3697);
xor U4132 (N_4132,N_3365,N_3946);
or U4133 (N_4133,N_3028,N_3746);
and U4134 (N_4134,N_3908,N_3068);
nand U4135 (N_4135,N_3884,N_3374);
nand U4136 (N_4136,N_3586,N_3534);
and U4137 (N_4137,N_3865,N_3640);
nor U4138 (N_4138,N_3096,N_3465);
or U4139 (N_4139,N_3999,N_3531);
or U4140 (N_4140,N_3010,N_3998);
nor U4141 (N_4141,N_3149,N_3504);
or U4142 (N_4142,N_3276,N_3120);
or U4143 (N_4143,N_3437,N_3904);
nand U4144 (N_4144,N_3541,N_3363);
and U4145 (N_4145,N_3568,N_3078);
nor U4146 (N_4146,N_3392,N_3059);
nor U4147 (N_4147,N_3008,N_3611);
nor U4148 (N_4148,N_3806,N_3965);
nand U4149 (N_4149,N_3811,N_3366);
and U4150 (N_4150,N_3167,N_3930);
nor U4151 (N_4151,N_3237,N_3991);
or U4152 (N_4152,N_3487,N_3670);
nor U4153 (N_4153,N_3840,N_3787);
and U4154 (N_4154,N_3535,N_3774);
nand U4155 (N_4155,N_3826,N_3181);
nand U4156 (N_4156,N_3718,N_3594);
or U4157 (N_4157,N_3000,N_3391);
nand U4158 (N_4158,N_3352,N_3242);
xnor U4159 (N_4159,N_3993,N_3523);
and U4160 (N_4160,N_3731,N_3100);
nand U4161 (N_4161,N_3418,N_3493);
nand U4162 (N_4162,N_3672,N_3983);
nand U4163 (N_4163,N_3639,N_3407);
or U4164 (N_4164,N_3663,N_3183);
and U4165 (N_4165,N_3419,N_3720);
nor U4166 (N_4166,N_3089,N_3159);
or U4167 (N_4167,N_3887,N_3278);
and U4168 (N_4168,N_3517,N_3906);
nor U4169 (N_4169,N_3143,N_3530);
and U4170 (N_4170,N_3942,N_3712);
and U4171 (N_4171,N_3061,N_3060);
or U4172 (N_4172,N_3769,N_3869);
nand U4173 (N_4173,N_3313,N_3650);
nor U4174 (N_4174,N_3544,N_3565);
nand U4175 (N_4175,N_3472,N_3094);
and U4176 (N_4176,N_3900,N_3372);
nor U4177 (N_4177,N_3542,N_3128);
xor U4178 (N_4178,N_3162,N_3430);
or U4179 (N_4179,N_3626,N_3622);
nand U4180 (N_4180,N_3481,N_3533);
or U4181 (N_4181,N_3397,N_3194);
nor U4182 (N_4182,N_3467,N_3125);
and U4183 (N_4183,N_3936,N_3717);
xnor U4184 (N_4184,N_3099,N_3584);
xnor U4185 (N_4185,N_3761,N_3850);
or U4186 (N_4186,N_3791,N_3583);
nor U4187 (N_4187,N_3416,N_3015);
xnor U4188 (N_4188,N_3083,N_3799);
or U4189 (N_4189,N_3018,N_3102);
and U4190 (N_4190,N_3863,N_3457);
or U4191 (N_4191,N_3251,N_3532);
and U4192 (N_4192,N_3505,N_3967);
nand U4193 (N_4193,N_3318,N_3478);
xor U4194 (N_4194,N_3411,N_3302);
nor U4195 (N_4195,N_3752,N_3741);
nor U4196 (N_4196,N_3050,N_3468);
nand U4197 (N_4197,N_3685,N_3191);
or U4198 (N_4198,N_3312,N_3864);
nor U4199 (N_4199,N_3203,N_3554);
nand U4200 (N_4200,N_3577,N_3597);
or U4201 (N_4201,N_3046,N_3309);
nor U4202 (N_4202,N_3429,N_3353);
nor U4203 (N_4203,N_3268,N_3119);
nor U4204 (N_4204,N_3168,N_3985);
or U4205 (N_4205,N_3295,N_3696);
or U4206 (N_4206,N_3893,N_3364);
and U4207 (N_4207,N_3379,N_3901);
nand U4208 (N_4208,N_3334,N_3383);
nand U4209 (N_4209,N_3315,N_3296);
or U4210 (N_4210,N_3727,N_3054);
or U4211 (N_4211,N_3322,N_3140);
nor U4212 (N_4212,N_3642,N_3265);
or U4213 (N_4213,N_3260,N_3641);
xor U4214 (N_4214,N_3658,N_3748);
nor U4215 (N_4215,N_3272,N_3066);
nand U4216 (N_4216,N_3454,N_3004);
or U4217 (N_4217,N_3537,N_3256);
xnor U4218 (N_4218,N_3835,N_3927);
or U4219 (N_4219,N_3178,N_3126);
nor U4220 (N_4220,N_3065,N_3513);
nand U4221 (N_4221,N_3786,N_3705);
or U4222 (N_4222,N_3466,N_3314);
or U4223 (N_4223,N_3917,N_3652);
and U4224 (N_4224,N_3615,N_3986);
and U4225 (N_4225,N_3134,N_3453);
or U4226 (N_4226,N_3356,N_3052);
or U4227 (N_4227,N_3196,N_3121);
or U4228 (N_4228,N_3212,N_3283);
nor U4229 (N_4229,N_3525,N_3695);
nand U4230 (N_4230,N_3747,N_3714);
and U4231 (N_4231,N_3350,N_3834);
or U4232 (N_4232,N_3422,N_3486);
nand U4233 (N_4233,N_3417,N_3469);
nand U4234 (N_4234,N_3796,N_3174);
or U4235 (N_4235,N_3035,N_3173);
nor U4236 (N_4236,N_3694,N_3818);
and U4237 (N_4237,N_3849,N_3745);
and U4238 (N_4238,N_3779,N_3920);
and U4239 (N_4239,N_3668,N_3014);
nor U4240 (N_4240,N_3235,N_3398);
or U4241 (N_4241,N_3213,N_3688);
or U4242 (N_4242,N_3876,N_3455);
and U4243 (N_4243,N_3914,N_3775);
nand U4244 (N_4244,N_3929,N_3421);
and U4245 (N_4245,N_3958,N_3193);
or U4246 (N_4246,N_3708,N_3773);
and U4247 (N_4247,N_3562,N_3659);
and U4248 (N_4248,N_3979,N_3836);
nor U4249 (N_4249,N_3859,N_3845);
nand U4250 (N_4250,N_3137,N_3228);
xor U4251 (N_4251,N_3907,N_3423);
nand U4252 (N_4252,N_3916,N_3793);
and U4253 (N_4253,N_3610,N_3524);
nor U4254 (N_4254,N_3843,N_3401);
and U4255 (N_4255,N_3291,N_3104);
and U4256 (N_4256,N_3357,N_3638);
nand U4257 (N_4257,N_3377,N_3507);
or U4258 (N_4258,N_3055,N_3107);
or U4259 (N_4259,N_3807,N_3150);
and U4260 (N_4260,N_3264,N_3163);
xnor U4261 (N_4261,N_3317,N_3601);
or U4262 (N_4262,N_3339,N_3477);
nand U4263 (N_4263,N_3962,N_3151);
or U4264 (N_4264,N_3828,N_3462);
nand U4265 (N_4265,N_3831,N_3898);
and U4266 (N_4266,N_3186,N_3036);
or U4267 (N_4267,N_3651,N_3804);
and U4268 (N_4268,N_3360,N_3964);
and U4269 (N_4269,N_3037,N_3665);
and U4270 (N_4270,N_3058,N_3816);
nor U4271 (N_4271,N_3114,N_3032);
or U4272 (N_4272,N_3223,N_3980);
or U4273 (N_4273,N_3699,N_3380);
and U4274 (N_4274,N_3819,N_3759);
or U4275 (N_4275,N_3225,N_3023);
nand U4276 (N_4276,N_3721,N_3069);
nand U4277 (N_4277,N_3197,N_3399);
or U4278 (N_4278,N_3077,N_3825);
or U4279 (N_4279,N_3637,N_3944);
nor U4280 (N_4280,N_3632,N_3798);
or U4281 (N_4281,N_3758,N_3647);
and U4282 (N_4282,N_3633,N_3446);
or U4283 (N_4283,N_3092,N_3141);
and U4284 (N_4284,N_3617,N_3536);
or U4285 (N_4285,N_3177,N_3861);
or U4286 (N_4286,N_3766,N_3981);
xnor U4287 (N_4287,N_3559,N_3649);
or U4288 (N_4288,N_3966,N_3491);
or U4289 (N_4289,N_3580,N_3405);
nor U4290 (N_4290,N_3232,N_3284);
xor U4291 (N_4291,N_3158,N_3664);
nand U4292 (N_4292,N_3483,N_3226);
or U4293 (N_4293,N_3239,N_3220);
nor U4294 (N_4294,N_3101,N_3978);
and U4295 (N_4295,N_3402,N_3968);
and U4296 (N_4296,N_3947,N_3560);
and U4297 (N_4297,N_3599,N_3038);
or U4298 (N_4298,N_3231,N_3394);
or U4299 (N_4299,N_3113,N_3335);
nand U4300 (N_4300,N_3780,N_3385);
nand U4301 (N_4301,N_3729,N_3123);
nand U4302 (N_4302,N_3540,N_3404);
xor U4303 (N_4303,N_3431,N_3341);
and U4304 (N_4304,N_3689,N_3783);
or U4305 (N_4305,N_3282,N_3439);
nor U4306 (N_4306,N_3890,N_3048);
and U4307 (N_4307,N_3616,N_3271);
nor U4308 (N_4308,N_3359,N_3527);
nor U4309 (N_4309,N_3182,N_3189);
xor U4310 (N_4310,N_3673,N_3367);
nand U4311 (N_4311,N_3165,N_3928);
nand U4312 (N_4312,N_3157,N_3546);
and U4313 (N_4313,N_3948,N_3005);
xor U4314 (N_4314,N_3801,N_3706);
or U4315 (N_4315,N_3262,N_3589);
and U4316 (N_4316,N_3029,N_3230);
or U4317 (N_4317,N_3926,N_3608);
and U4318 (N_4318,N_3937,N_3924);
xor U4319 (N_4319,N_3240,N_3732);
nand U4320 (N_4320,N_3676,N_3743);
or U4321 (N_4321,N_3571,N_3076);
nand U4322 (N_4322,N_3585,N_3692);
nor U4323 (N_4323,N_3085,N_3733);
or U4324 (N_4324,N_3185,N_3447);
xor U4325 (N_4325,N_3837,N_3388);
xnor U4326 (N_4326,N_3368,N_3145);
or U4327 (N_4327,N_3413,N_3822);
and U4328 (N_4328,N_3459,N_3702);
and U4329 (N_4329,N_3389,N_3355);
or U4330 (N_4330,N_3445,N_3460);
and U4331 (N_4331,N_3424,N_3715);
and U4332 (N_4332,N_3275,N_3277);
and U4333 (N_4333,N_3156,N_3187);
or U4334 (N_4334,N_3346,N_3933);
nor U4335 (N_4335,N_3557,N_3166);
and U4336 (N_4336,N_3753,N_3873);
nor U4337 (N_4337,N_3261,N_3221);
and U4338 (N_4338,N_3903,N_3449);
nor U4339 (N_4339,N_3810,N_3988);
nor U4340 (N_4340,N_3310,N_3458);
nand U4341 (N_4341,N_3475,N_3169);
or U4342 (N_4342,N_3619,N_3308);
nor U4343 (N_4343,N_3922,N_3122);
and U4344 (N_4344,N_3326,N_3960);
or U4345 (N_4345,N_3627,N_3082);
nor U4346 (N_4346,N_3502,N_3464);
or U4347 (N_4347,N_3362,N_3877);
nor U4348 (N_4348,N_3739,N_3598);
nor U4349 (N_4349,N_3889,N_3509);
xnor U4350 (N_4350,N_3300,N_3063);
or U4351 (N_4351,N_3872,N_3722);
nand U4352 (N_4352,N_3146,N_3171);
nor U4353 (N_4353,N_3244,N_3307);
or U4354 (N_4354,N_3337,N_3093);
or U4355 (N_4355,N_3316,N_3734);
and U4356 (N_4356,N_3007,N_3208);
nand U4357 (N_4357,N_3129,N_3057);
and U4358 (N_4358,N_3555,N_3841);
nor U4359 (N_4359,N_3820,N_3210);
or U4360 (N_4360,N_3211,N_3153);
or U4361 (N_4361,N_3574,N_3190);
nor U4362 (N_4362,N_3959,N_3558);
nand U4363 (N_4363,N_3797,N_3319);
or U4364 (N_4364,N_3522,N_3386);
nor U4365 (N_4365,N_3306,N_3009);
or U4366 (N_4366,N_3412,N_3222);
nor U4367 (N_4367,N_3086,N_3736);
nor U4368 (N_4368,N_3987,N_3844);
xor U4369 (N_4369,N_3931,N_3019);
nor U4370 (N_4370,N_3934,N_3409);
nor U4371 (N_4371,N_3956,N_3860);
nand U4372 (N_4372,N_3266,N_3133);
or U4373 (N_4373,N_3047,N_3305);
xor U4374 (N_4374,N_3515,N_3155);
nand U4375 (N_4375,N_3425,N_3420);
and U4376 (N_4376,N_3049,N_3070);
xnor U4377 (N_4377,N_3909,N_3600);
nor U4378 (N_4378,N_3740,N_3588);
nor U4379 (N_4379,N_3803,N_3450);
and U4380 (N_4380,N_3257,N_3042);
nor U4381 (N_4381,N_3105,N_3620);
and U4382 (N_4382,N_3744,N_3506);
nand U4383 (N_4383,N_3881,N_3879);
xnor U4384 (N_4384,N_3476,N_3246);
or U4385 (N_4385,N_3433,N_3384);
or U4386 (N_4386,N_3882,N_3847);
and U4387 (N_4387,N_3219,N_3905);
nor U4388 (N_4388,N_3829,N_3292);
xnor U4389 (N_4389,N_3750,N_3375);
and U4390 (N_4390,N_3939,N_3723);
xnor U4391 (N_4391,N_3051,N_3961);
nor U4392 (N_4392,N_3361,N_3943);
nand U4393 (N_4393,N_3547,N_3771);
nand U4394 (N_4394,N_3842,N_3578);
or U4395 (N_4395,N_3426,N_3116);
nand U4396 (N_4396,N_3245,N_3263);
nor U4397 (N_4397,N_3989,N_3858);
and U4398 (N_4398,N_3088,N_3808);
xor U4399 (N_4399,N_3432,N_3299);
or U4400 (N_4400,N_3728,N_3108);
xnor U4401 (N_4401,N_3144,N_3195);
or U4402 (N_4402,N_3990,N_3347);
and U4403 (N_4403,N_3020,N_3204);
nor U4404 (N_4404,N_3767,N_3662);
nor U4405 (N_4405,N_3618,N_3485);
nor U4406 (N_4406,N_3269,N_3090);
nor U4407 (N_4407,N_3258,N_3874);
nor U4408 (N_4408,N_3259,N_3434);
nor U4409 (N_4409,N_3955,N_3564);
nand U4410 (N_4410,N_3130,N_3378);
nor U4411 (N_4411,N_3241,N_3025);
and U4412 (N_4412,N_3925,N_3013);
nor U4413 (N_4413,N_3764,N_3444);
nor U4414 (N_4414,N_3403,N_3395);
nand U4415 (N_4415,N_3324,N_3497);
nand U4416 (N_4416,N_3451,N_3749);
and U4417 (N_4417,N_3551,N_3765);
nand U4418 (N_4418,N_3248,N_3044);
or U4419 (N_4419,N_3894,N_3675);
or U4420 (N_4420,N_3344,N_3040);
and U4421 (N_4421,N_3280,N_3142);
and U4422 (N_4422,N_3897,N_3139);
or U4423 (N_4423,N_3921,N_3501);
nor U4424 (N_4424,N_3853,N_3249);
or U4425 (N_4425,N_3556,N_3496);
nor U4426 (N_4426,N_3490,N_3095);
nor U4427 (N_4427,N_3595,N_3963);
and U4428 (N_4428,N_3790,N_3602);
or U4429 (N_4429,N_3704,N_3868);
and U4430 (N_4430,N_3550,N_3891);
nor U4431 (N_4431,N_3833,N_3643);
nor U4432 (N_4432,N_3519,N_3408);
and U4433 (N_4433,N_3236,N_3118);
xnor U4434 (N_4434,N_3629,N_3323);
nand U4435 (N_4435,N_3569,N_3192);
nand U4436 (N_4436,N_3273,N_3607);
xor U4437 (N_4437,N_3682,N_3124);
nor U4438 (N_4438,N_3976,N_3250);
nor U4439 (N_4439,N_3098,N_3474);
and U4440 (N_4440,N_3062,N_3499);
or U4441 (N_4441,N_3606,N_3084);
and U4442 (N_4442,N_3006,N_3911);
nand U4443 (N_4443,N_3730,N_3770);
or U4444 (N_4444,N_3138,N_3995);
nand U4445 (N_4445,N_3224,N_3671);
or U4446 (N_4446,N_3870,N_3654);
nand U4447 (N_4447,N_3254,N_3539);
or U4448 (N_4448,N_3207,N_3170);
or U4449 (N_4449,N_3482,N_3026);
or U4450 (N_4450,N_3802,N_3795);
nor U4451 (N_4451,N_3590,N_3895);
nor U4452 (N_4452,N_3508,N_3592);
xor U4453 (N_4453,N_3410,N_3011);
or U4454 (N_4454,N_3021,N_3495);
and U4455 (N_4455,N_3553,N_3382);
nor U4456 (N_4456,N_3340,N_3033);
nand U4457 (N_4457,N_3180,N_3538);
nor U4458 (N_4458,N_3852,N_3131);
and U4459 (N_4459,N_3609,N_3285);
nand U4460 (N_4460,N_3587,N_3848);
xnor U4461 (N_4461,N_3470,N_3628);
nand U4462 (N_4462,N_3854,N_3369);
nand U4463 (N_4463,N_3655,N_3572);
and U4464 (N_4464,N_3563,N_3075);
nor U4465 (N_4465,N_3545,N_3713);
nor U4466 (N_4466,N_3376,N_3851);
nand U4467 (N_4467,N_3604,N_3289);
or U4468 (N_4468,N_3862,N_3293);
nand U4469 (N_4469,N_3243,N_3789);
and U4470 (N_4470,N_3489,N_3832);
nor U4471 (N_4471,N_3463,N_3735);
and U4472 (N_4472,N_3112,N_3017);
and U4473 (N_4473,N_3814,N_3912);
nor U4474 (N_4474,N_3301,N_3888);
xor U4475 (N_4475,N_3279,N_3160);
and U4476 (N_4476,N_3975,N_3698);
nand U4477 (N_4477,N_3255,N_3630);
nand U4478 (N_4478,N_3784,N_3977);
nand U4479 (N_4479,N_3994,N_3073);
and U4480 (N_4480,N_3945,N_3175);
and U4481 (N_4481,N_3756,N_3785);
and U4482 (N_4482,N_3348,N_3045);
and U4483 (N_4483,N_3511,N_3373);
nand U4484 (N_4484,N_3267,N_3724);
and U4485 (N_4485,N_3097,N_3298);
nand U4486 (N_4486,N_3666,N_3390);
nor U4487 (N_4487,N_3288,N_3777);
or U4488 (N_4488,N_3351,N_3915);
nor U4489 (N_4489,N_3516,N_3510);
and U4490 (N_4490,N_3206,N_3117);
and U4491 (N_4491,N_3179,N_3940);
nor U4492 (N_4492,N_3794,N_3935);
nor U4493 (N_4493,N_3115,N_3027);
xnor U4494 (N_4494,N_3349,N_3674);
nand U4495 (N_4495,N_3436,N_3838);
and U4496 (N_4496,N_3304,N_3952);
nand U4497 (N_4497,N_3214,N_3932);
nand U4498 (N_4498,N_3396,N_3176);
xnor U4499 (N_4499,N_3161,N_3885);
and U4500 (N_4500,N_3581,N_3016);
nor U4501 (N_4501,N_3654,N_3802);
and U4502 (N_4502,N_3026,N_3331);
nand U4503 (N_4503,N_3808,N_3589);
or U4504 (N_4504,N_3638,N_3067);
and U4505 (N_4505,N_3368,N_3323);
xor U4506 (N_4506,N_3912,N_3544);
nor U4507 (N_4507,N_3340,N_3106);
nand U4508 (N_4508,N_3772,N_3269);
or U4509 (N_4509,N_3987,N_3483);
or U4510 (N_4510,N_3227,N_3969);
or U4511 (N_4511,N_3848,N_3800);
nand U4512 (N_4512,N_3118,N_3696);
nor U4513 (N_4513,N_3836,N_3433);
or U4514 (N_4514,N_3848,N_3973);
or U4515 (N_4515,N_3007,N_3472);
or U4516 (N_4516,N_3663,N_3810);
nand U4517 (N_4517,N_3355,N_3422);
nor U4518 (N_4518,N_3376,N_3291);
nand U4519 (N_4519,N_3659,N_3041);
and U4520 (N_4520,N_3082,N_3263);
or U4521 (N_4521,N_3922,N_3165);
and U4522 (N_4522,N_3727,N_3186);
nand U4523 (N_4523,N_3230,N_3383);
nor U4524 (N_4524,N_3422,N_3541);
or U4525 (N_4525,N_3576,N_3940);
nor U4526 (N_4526,N_3224,N_3514);
nand U4527 (N_4527,N_3884,N_3301);
or U4528 (N_4528,N_3545,N_3477);
nand U4529 (N_4529,N_3843,N_3110);
or U4530 (N_4530,N_3299,N_3671);
nor U4531 (N_4531,N_3794,N_3687);
and U4532 (N_4532,N_3564,N_3641);
and U4533 (N_4533,N_3435,N_3869);
xor U4534 (N_4534,N_3488,N_3198);
xor U4535 (N_4535,N_3771,N_3355);
nor U4536 (N_4536,N_3218,N_3918);
or U4537 (N_4537,N_3084,N_3529);
nand U4538 (N_4538,N_3097,N_3534);
nand U4539 (N_4539,N_3308,N_3016);
and U4540 (N_4540,N_3301,N_3438);
nor U4541 (N_4541,N_3982,N_3997);
xor U4542 (N_4542,N_3805,N_3087);
or U4543 (N_4543,N_3479,N_3436);
nor U4544 (N_4544,N_3870,N_3198);
and U4545 (N_4545,N_3134,N_3143);
nand U4546 (N_4546,N_3322,N_3462);
nor U4547 (N_4547,N_3532,N_3444);
nor U4548 (N_4548,N_3753,N_3886);
nor U4549 (N_4549,N_3634,N_3884);
xnor U4550 (N_4550,N_3098,N_3752);
or U4551 (N_4551,N_3946,N_3716);
or U4552 (N_4552,N_3771,N_3588);
nor U4553 (N_4553,N_3860,N_3466);
and U4554 (N_4554,N_3297,N_3974);
or U4555 (N_4555,N_3124,N_3388);
nor U4556 (N_4556,N_3754,N_3960);
or U4557 (N_4557,N_3389,N_3139);
nor U4558 (N_4558,N_3325,N_3028);
and U4559 (N_4559,N_3815,N_3435);
nand U4560 (N_4560,N_3901,N_3730);
and U4561 (N_4561,N_3204,N_3235);
and U4562 (N_4562,N_3506,N_3007);
nand U4563 (N_4563,N_3377,N_3213);
nand U4564 (N_4564,N_3778,N_3217);
nor U4565 (N_4565,N_3401,N_3406);
or U4566 (N_4566,N_3417,N_3969);
nand U4567 (N_4567,N_3891,N_3304);
nor U4568 (N_4568,N_3936,N_3908);
and U4569 (N_4569,N_3145,N_3482);
or U4570 (N_4570,N_3804,N_3799);
or U4571 (N_4571,N_3426,N_3985);
nor U4572 (N_4572,N_3300,N_3882);
nor U4573 (N_4573,N_3787,N_3270);
xnor U4574 (N_4574,N_3208,N_3633);
nor U4575 (N_4575,N_3574,N_3579);
nor U4576 (N_4576,N_3540,N_3326);
nand U4577 (N_4577,N_3796,N_3411);
and U4578 (N_4578,N_3821,N_3663);
or U4579 (N_4579,N_3097,N_3498);
nor U4580 (N_4580,N_3049,N_3144);
and U4581 (N_4581,N_3993,N_3417);
or U4582 (N_4582,N_3820,N_3391);
and U4583 (N_4583,N_3198,N_3412);
or U4584 (N_4584,N_3269,N_3532);
or U4585 (N_4585,N_3879,N_3404);
and U4586 (N_4586,N_3329,N_3440);
nand U4587 (N_4587,N_3388,N_3806);
xnor U4588 (N_4588,N_3011,N_3342);
or U4589 (N_4589,N_3326,N_3339);
and U4590 (N_4590,N_3114,N_3962);
or U4591 (N_4591,N_3380,N_3169);
and U4592 (N_4592,N_3699,N_3475);
nor U4593 (N_4593,N_3859,N_3656);
and U4594 (N_4594,N_3578,N_3483);
nand U4595 (N_4595,N_3483,N_3054);
or U4596 (N_4596,N_3144,N_3478);
nor U4597 (N_4597,N_3672,N_3464);
or U4598 (N_4598,N_3567,N_3667);
or U4599 (N_4599,N_3163,N_3047);
nor U4600 (N_4600,N_3898,N_3031);
and U4601 (N_4601,N_3112,N_3778);
and U4602 (N_4602,N_3772,N_3712);
or U4603 (N_4603,N_3304,N_3910);
or U4604 (N_4604,N_3758,N_3322);
or U4605 (N_4605,N_3197,N_3931);
nor U4606 (N_4606,N_3021,N_3611);
xnor U4607 (N_4607,N_3150,N_3249);
xor U4608 (N_4608,N_3625,N_3091);
nand U4609 (N_4609,N_3762,N_3217);
or U4610 (N_4610,N_3515,N_3318);
xor U4611 (N_4611,N_3175,N_3088);
nor U4612 (N_4612,N_3034,N_3856);
nor U4613 (N_4613,N_3481,N_3130);
or U4614 (N_4614,N_3485,N_3144);
and U4615 (N_4615,N_3643,N_3517);
or U4616 (N_4616,N_3959,N_3532);
nor U4617 (N_4617,N_3205,N_3552);
and U4618 (N_4618,N_3729,N_3849);
nor U4619 (N_4619,N_3606,N_3483);
and U4620 (N_4620,N_3260,N_3512);
or U4621 (N_4621,N_3157,N_3629);
and U4622 (N_4622,N_3456,N_3696);
nand U4623 (N_4623,N_3402,N_3206);
xnor U4624 (N_4624,N_3271,N_3877);
nor U4625 (N_4625,N_3579,N_3449);
nand U4626 (N_4626,N_3585,N_3491);
nor U4627 (N_4627,N_3883,N_3136);
nor U4628 (N_4628,N_3524,N_3485);
nand U4629 (N_4629,N_3302,N_3752);
xor U4630 (N_4630,N_3901,N_3759);
or U4631 (N_4631,N_3825,N_3967);
and U4632 (N_4632,N_3020,N_3628);
or U4633 (N_4633,N_3235,N_3707);
or U4634 (N_4634,N_3004,N_3030);
or U4635 (N_4635,N_3613,N_3309);
and U4636 (N_4636,N_3808,N_3959);
and U4637 (N_4637,N_3624,N_3944);
or U4638 (N_4638,N_3415,N_3373);
nand U4639 (N_4639,N_3426,N_3787);
and U4640 (N_4640,N_3031,N_3609);
xnor U4641 (N_4641,N_3942,N_3255);
nand U4642 (N_4642,N_3528,N_3499);
and U4643 (N_4643,N_3957,N_3333);
nand U4644 (N_4644,N_3637,N_3660);
or U4645 (N_4645,N_3139,N_3021);
nor U4646 (N_4646,N_3355,N_3621);
nor U4647 (N_4647,N_3035,N_3156);
xor U4648 (N_4648,N_3470,N_3137);
and U4649 (N_4649,N_3419,N_3345);
or U4650 (N_4650,N_3038,N_3864);
nand U4651 (N_4651,N_3250,N_3142);
and U4652 (N_4652,N_3084,N_3602);
and U4653 (N_4653,N_3807,N_3788);
and U4654 (N_4654,N_3219,N_3358);
and U4655 (N_4655,N_3667,N_3206);
nand U4656 (N_4656,N_3961,N_3360);
or U4657 (N_4657,N_3782,N_3615);
nand U4658 (N_4658,N_3891,N_3702);
nand U4659 (N_4659,N_3403,N_3556);
and U4660 (N_4660,N_3522,N_3709);
nand U4661 (N_4661,N_3092,N_3963);
nor U4662 (N_4662,N_3154,N_3507);
nand U4663 (N_4663,N_3380,N_3882);
or U4664 (N_4664,N_3651,N_3294);
xnor U4665 (N_4665,N_3539,N_3829);
and U4666 (N_4666,N_3362,N_3587);
and U4667 (N_4667,N_3763,N_3318);
and U4668 (N_4668,N_3718,N_3144);
or U4669 (N_4669,N_3272,N_3835);
nor U4670 (N_4670,N_3508,N_3351);
and U4671 (N_4671,N_3459,N_3408);
xnor U4672 (N_4672,N_3623,N_3213);
xor U4673 (N_4673,N_3978,N_3006);
nand U4674 (N_4674,N_3313,N_3182);
or U4675 (N_4675,N_3372,N_3801);
nand U4676 (N_4676,N_3220,N_3636);
or U4677 (N_4677,N_3807,N_3366);
or U4678 (N_4678,N_3250,N_3940);
and U4679 (N_4679,N_3852,N_3305);
nor U4680 (N_4680,N_3326,N_3191);
nand U4681 (N_4681,N_3468,N_3371);
or U4682 (N_4682,N_3473,N_3431);
or U4683 (N_4683,N_3413,N_3192);
xor U4684 (N_4684,N_3126,N_3006);
nor U4685 (N_4685,N_3602,N_3604);
nand U4686 (N_4686,N_3469,N_3875);
or U4687 (N_4687,N_3271,N_3749);
nand U4688 (N_4688,N_3210,N_3589);
nor U4689 (N_4689,N_3265,N_3675);
and U4690 (N_4690,N_3007,N_3014);
nor U4691 (N_4691,N_3676,N_3513);
nor U4692 (N_4692,N_3535,N_3006);
nor U4693 (N_4693,N_3044,N_3502);
nand U4694 (N_4694,N_3287,N_3766);
nor U4695 (N_4695,N_3034,N_3446);
nand U4696 (N_4696,N_3244,N_3109);
nor U4697 (N_4697,N_3745,N_3620);
or U4698 (N_4698,N_3703,N_3800);
nor U4699 (N_4699,N_3924,N_3288);
or U4700 (N_4700,N_3390,N_3718);
nand U4701 (N_4701,N_3751,N_3249);
and U4702 (N_4702,N_3329,N_3073);
nor U4703 (N_4703,N_3645,N_3158);
nor U4704 (N_4704,N_3210,N_3074);
or U4705 (N_4705,N_3357,N_3489);
and U4706 (N_4706,N_3661,N_3059);
nor U4707 (N_4707,N_3805,N_3549);
nand U4708 (N_4708,N_3965,N_3876);
or U4709 (N_4709,N_3974,N_3231);
nand U4710 (N_4710,N_3817,N_3731);
and U4711 (N_4711,N_3045,N_3767);
xnor U4712 (N_4712,N_3883,N_3714);
nand U4713 (N_4713,N_3298,N_3700);
nor U4714 (N_4714,N_3581,N_3085);
nand U4715 (N_4715,N_3113,N_3767);
and U4716 (N_4716,N_3828,N_3198);
nor U4717 (N_4717,N_3063,N_3299);
nand U4718 (N_4718,N_3724,N_3289);
nor U4719 (N_4719,N_3613,N_3542);
nand U4720 (N_4720,N_3771,N_3360);
or U4721 (N_4721,N_3196,N_3146);
nor U4722 (N_4722,N_3914,N_3966);
nor U4723 (N_4723,N_3592,N_3002);
or U4724 (N_4724,N_3719,N_3446);
and U4725 (N_4725,N_3635,N_3852);
nand U4726 (N_4726,N_3078,N_3535);
or U4727 (N_4727,N_3874,N_3469);
nor U4728 (N_4728,N_3773,N_3632);
nor U4729 (N_4729,N_3640,N_3641);
or U4730 (N_4730,N_3099,N_3755);
and U4731 (N_4731,N_3819,N_3339);
and U4732 (N_4732,N_3867,N_3248);
and U4733 (N_4733,N_3807,N_3655);
nand U4734 (N_4734,N_3897,N_3946);
nand U4735 (N_4735,N_3454,N_3647);
nor U4736 (N_4736,N_3702,N_3904);
or U4737 (N_4737,N_3264,N_3066);
or U4738 (N_4738,N_3170,N_3819);
and U4739 (N_4739,N_3955,N_3932);
and U4740 (N_4740,N_3210,N_3870);
and U4741 (N_4741,N_3347,N_3454);
nand U4742 (N_4742,N_3420,N_3170);
nor U4743 (N_4743,N_3639,N_3976);
nand U4744 (N_4744,N_3795,N_3603);
nand U4745 (N_4745,N_3406,N_3108);
nand U4746 (N_4746,N_3491,N_3809);
and U4747 (N_4747,N_3784,N_3460);
nor U4748 (N_4748,N_3995,N_3744);
nand U4749 (N_4749,N_3166,N_3453);
nand U4750 (N_4750,N_3856,N_3646);
and U4751 (N_4751,N_3842,N_3232);
and U4752 (N_4752,N_3217,N_3959);
xor U4753 (N_4753,N_3802,N_3844);
or U4754 (N_4754,N_3396,N_3017);
or U4755 (N_4755,N_3602,N_3752);
nor U4756 (N_4756,N_3128,N_3585);
and U4757 (N_4757,N_3198,N_3294);
and U4758 (N_4758,N_3954,N_3669);
nand U4759 (N_4759,N_3080,N_3799);
or U4760 (N_4760,N_3162,N_3398);
xor U4761 (N_4761,N_3855,N_3823);
nor U4762 (N_4762,N_3142,N_3685);
nand U4763 (N_4763,N_3552,N_3301);
and U4764 (N_4764,N_3032,N_3217);
and U4765 (N_4765,N_3212,N_3672);
and U4766 (N_4766,N_3195,N_3226);
and U4767 (N_4767,N_3143,N_3066);
xor U4768 (N_4768,N_3221,N_3496);
and U4769 (N_4769,N_3683,N_3951);
and U4770 (N_4770,N_3398,N_3404);
or U4771 (N_4771,N_3951,N_3070);
nand U4772 (N_4772,N_3743,N_3772);
nand U4773 (N_4773,N_3097,N_3591);
or U4774 (N_4774,N_3647,N_3414);
nor U4775 (N_4775,N_3001,N_3367);
nand U4776 (N_4776,N_3137,N_3362);
or U4777 (N_4777,N_3108,N_3908);
nor U4778 (N_4778,N_3484,N_3449);
and U4779 (N_4779,N_3543,N_3944);
nand U4780 (N_4780,N_3270,N_3525);
nand U4781 (N_4781,N_3137,N_3216);
and U4782 (N_4782,N_3447,N_3514);
nor U4783 (N_4783,N_3788,N_3047);
and U4784 (N_4784,N_3416,N_3126);
and U4785 (N_4785,N_3959,N_3193);
xor U4786 (N_4786,N_3372,N_3695);
nor U4787 (N_4787,N_3819,N_3858);
nor U4788 (N_4788,N_3361,N_3352);
or U4789 (N_4789,N_3126,N_3504);
nor U4790 (N_4790,N_3263,N_3160);
and U4791 (N_4791,N_3855,N_3083);
nor U4792 (N_4792,N_3764,N_3592);
or U4793 (N_4793,N_3611,N_3052);
or U4794 (N_4794,N_3891,N_3364);
or U4795 (N_4795,N_3164,N_3992);
or U4796 (N_4796,N_3388,N_3767);
or U4797 (N_4797,N_3959,N_3972);
and U4798 (N_4798,N_3914,N_3456);
nand U4799 (N_4799,N_3597,N_3612);
nor U4800 (N_4800,N_3950,N_3298);
or U4801 (N_4801,N_3118,N_3653);
and U4802 (N_4802,N_3794,N_3341);
and U4803 (N_4803,N_3096,N_3692);
nand U4804 (N_4804,N_3256,N_3668);
nor U4805 (N_4805,N_3594,N_3789);
nand U4806 (N_4806,N_3194,N_3571);
or U4807 (N_4807,N_3290,N_3304);
xnor U4808 (N_4808,N_3264,N_3549);
and U4809 (N_4809,N_3184,N_3914);
nor U4810 (N_4810,N_3208,N_3120);
nand U4811 (N_4811,N_3082,N_3511);
nor U4812 (N_4812,N_3782,N_3123);
nor U4813 (N_4813,N_3885,N_3827);
nand U4814 (N_4814,N_3175,N_3091);
or U4815 (N_4815,N_3681,N_3800);
or U4816 (N_4816,N_3369,N_3220);
nor U4817 (N_4817,N_3955,N_3354);
or U4818 (N_4818,N_3844,N_3382);
nor U4819 (N_4819,N_3126,N_3305);
or U4820 (N_4820,N_3951,N_3569);
and U4821 (N_4821,N_3124,N_3724);
and U4822 (N_4822,N_3464,N_3859);
and U4823 (N_4823,N_3057,N_3530);
nand U4824 (N_4824,N_3332,N_3833);
or U4825 (N_4825,N_3042,N_3983);
nand U4826 (N_4826,N_3432,N_3730);
and U4827 (N_4827,N_3399,N_3186);
or U4828 (N_4828,N_3761,N_3747);
nor U4829 (N_4829,N_3258,N_3206);
or U4830 (N_4830,N_3592,N_3084);
nand U4831 (N_4831,N_3533,N_3541);
or U4832 (N_4832,N_3205,N_3370);
nand U4833 (N_4833,N_3421,N_3477);
and U4834 (N_4834,N_3263,N_3641);
nor U4835 (N_4835,N_3456,N_3851);
and U4836 (N_4836,N_3916,N_3119);
nand U4837 (N_4837,N_3821,N_3278);
nand U4838 (N_4838,N_3915,N_3754);
and U4839 (N_4839,N_3722,N_3142);
and U4840 (N_4840,N_3775,N_3353);
or U4841 (N_4841,N_3012,N_3282);
or U4842 (N_4842,N_3708,N_3010);
or U4843 (N_4843,N_3554,N_3891);
and U4844 (N_4844,N_3082,N_3594);
or U4845 (N_4845,N_3252,N_3568);
nor U4846 (N_4846,N_3934,N_3400);
or U4847 (N_4847,N_3472,N_3413);
or U4848 (N_4848,N_3766,N_3564);
and U4849 (N_4849,N_3917,N_3035);
nand U4850 (N_4850,N_3494,N_3514);
and U4851 (N_4851,N_3369,N_3632);
or U4852 (N_4852,N_3598,N_3701);
nand U4853 (N_4853,N_3163,N_3509);
xnor U4854 (N_4854,N_3226,N_3601);
nand U4855 (N_4855,N_3885,N_3547);
nand U4856 (N_4856,N_3416,N_3967);
or U4857 (N_4857,N_3818,N_3497);
nand U4858 (N_4858,N_3984,N_3033);
nand U4859 (N_4859,N_3981,N_3246);
nor U4860 (N_4860,N_3068,N_3779);
nand U4861 (N_4861,N_3496,N_3503);
and U4862 (N_4862,N_3216,N_3192);
and U4863 (N_4863,N_3227,N_3223);
nand U4864 (N_4864,N_3212,N_3542);
and U4865 (N_4865,N_3951,N_3284);
nor U4866 (N_4866,N_3459,N_3379);
nand U4867 (N_4867,N_3850,N_3095);
and U4868 (N_4868,N_3999,N_3339);
nor U4869 (N_4869,N_3564,N_3305);
nand U4870 (N_4870,N_3350,N_3337);
nor U4871 (N_4871,N_3765,N_3857);
and U4872 (N_4872,N_3281,N_3333);
nor U4873 (N_4873,N_3918,N_3056);
nor U4874 (N_4874,N_3376,N_3554);
nor U4875 (N_4875,N_3522,N_3814);
nor U4876 (N_4876,N_3239,N_3537);
xor U4877 (N_4877,N_3374,N_3806);
xnor U4878 (N_4878,N_3447,N_3686);
nand U4879 (N_4879,N_3898,N_3145);
xnor U4880 (N_4880,N_3839,N_3964);
nand U4881 (N_4881,N_3300,N_3781);
and U4882 (N_4882,N_3482,N_3204);
or U4883 (N_4883,N_3696,N_3288);
or U4884 (N_4884,N_3209,N_3827);
nor U4885 (N_4885,N_3719,N_3627);
nor U4886 (N_4886,N_3133,N_3183);
nand U4887 (N_4887,N_3065,N_3958);
nor U4888 (N_4888,N_3488,N_3549);
nor U4889 (N_4889,N_3006,N_3685);
nor U4890 (N_4890,N_3389,N_3048);
nand U4891 (N_4891,N_3046,N_3485);
and U4892 (N_4892,N_3009,N_3286);
and U4893 (N_4893,N_3091,N_3047);
and U4894 (N_4894,N_3457,N_3304);
nor U4895 (N_4895,N_3498,N_3571);
xnor U4896 (N_4896,N_3703,N_3273);
nor U4897 (N_4897,N_3731,N_3121);
nor U4898 (N_4898,N_3433,N_3953);
or U4899 (N_4899,N_3957,N_3472);
or U4900 (N_4900,N_3320,N_3133);
nor U4901 (N_4901,N_3161,N_3367);
nand U4902 (N_4902,N_3588,N_3573);
nand U4903 (N_4903,N_3613,N_3044);
nor U4904 (N_4904,N_3692,N_3812);
nor U4905 (N_4905,N_3037,N_3560);
and U4906 (N_4906,N_3847,N_3464);
and U4907 (N_4907,N_3232,N_3558);
nand U4908 (N_4908,N_3437,N_3743);
or U4909 (N_4909,N_3357,N_3165);
and U4910 (N_4910,N_3716,N_3398);
nand U4911 (N_4911,N_3886,N_3123);
nor U4912 (N_4912,N_3953,N_3735);
or U4913 (N_4913,N_3216,N_3630);
or U4914 (N_4914,N_3584,N_3690);
nor U4915 (N_4915,N_3363,N_3538);
nor U4916 (N_4916,N_3982,N_3801);
or U4917 (N_4917,N_3140,N_3651);
and U4918 (N_4918,N_3559,N_3234);
and U4919 (N_4919,N_3514,N_3363);
nand U4920 (N_4920,N_3521,N_3412);
nor U4921 (N_4921,N_3811,N_3768);
xor U4922 (N_4922,N_3564,N_3289);
and U4923 (N_4923,N_3995,N_3757);
nor U4924 (N_4924,N_3341,N_3387);
or U4925 (N_4925,N_3448,N_3332);
nand U4926 (N_4926,N_3598,N_3383);
and U4927 (N_4927,N_3819,N_3936);
xor U4928 (N_4928,N_3936,N_3692);
and U4929 (N_4929,N_3230,N_3033);
nand U4930 (N_4930,N_3877,N_3758);
nand U4931 (N_4931,N_3854,N_3239);
and U4932 (N_4932,N_3061,N_3748);
nor U4933 (N_4933,N_3474,N_3361);
nand U4934 (N_4934,N_3341,N_3570);
or U4935 (N_4935,N_3036,N_3241);
nand U4936 (N_4936,N_3088,N_3062);
and U4937 (N_4937,N_3286,N_3765);
xor U4938 (N_4938,N_3849,N_3439);
nor U4939 (N_4939,N_3082,N_3167);
nand U4940 (N_4940,N_3464,N_3775);
and U4941 (N_4941,N_3678,N_3319);
nor U4942 (N_4942,N_3252,N_3328);
nor U4943 (N_4943,N_3471,N_3871);
xnor U4944 (N_4944,N_3716,N_3545);
or U4945 (N_4945,N_3389,N_3163);
nand U4946 (N_4946,N_3432,N_3740);
or U4947 (N_4947,N_3111,N_3163);
nand U4948 (N_4948,N_3511,N_3140);
nor U4949 (N_4949,N_3562,N_3867);
nor U4950 (N_4950,N_3390,N_3171);
or U4951 (N_4951,N_3908,N_3788);
nand U4952 (N_4952,N_3775,N_3345);
nand U4953 (N_4953,N_3364,N_3140);
and U4954 (N_4954,N_3507,N_3879);
or U4955 (N_4955,N_3475,N_3007);
nand U4956 (N_4956,N_3372,N_3189);
or U4957 (N_4957,N_3793,N_3871);
and U4958 (N_4958,N_3627,N_3359);
or U4959 (N_4959,N_3117,N_3108);
nand U4960 (N_4960,N_3083,N_3216);
and U4961 (N_4961,N_3813,N_3858);
nand U4962 (N_4962,N_3716,N_3726);
nand U4963 (N_4963,N_3210,N_3715);
or U4964 (N_4964,N_3464,N_3927);
nor U4965 (N_4965,N_3711,N_3796);
nor U4966 (N_4966,N_3908,N_3916);
nand U4967 (N_4967,N_3631,N_3299);
nand U4968 (N_4968,N_3948,N_3353);
xnor U4969 (N_4969,N_3806,N_3477);
nand U4970 (N_4970,N_3872,N_3857);
and U4971 (N_4971,N_3503,N_3485);
xor U4972 (N_4972,N_3523,N_3117);
and U4973 (N_4973,N_3938,N_3634);
or U4974 (N_4974,N_3210,N_3214);
or U4975 (N_4975,N_3892,N_3172);
or U4976 (N_4976,N_3796,N_3512);
nand U4977 (N_4977,N_3626,N_3474);
and U4978 (N_4978,N_3108,N_3985);
nand U4979 (N_4979,N_3726,N_3353);
or U4980 (N_4980,N_3606,N_3898);
or U4981 (N_4981,N_3064,N_3213);
nor U4982 (N_4982,N_3541,N_3845);
or U4983 (N_4983,N_3392,N_3033);
xnor U4984 (N_4984,N_3778,N_3714);
xor U4985 (N_4985,N_3845,N_3940);
or U4986 (N_4986,N_3041,N_3515);
and U4987 (N_4987,N_3416,N_3838);
or U4988 (N_4988,N_3294,N_3047);
nor U4989 (N_4989,N_3667,N_3448);
xor U4990 (N_4990,N_3659,N_3914);
nor U4991 (N_4991,N_3696,N_3840);
xnor U4992 (N_4992,N_3541,N_3481);
or U4993 (N_4993,N_3955,N_3709);
nand U4994 (N_4994,N_3494,N_3429);
nand U4995 (N_4995,N_3111,N_3311);
xnor U4996 (N_4996,N_3197,N_3633);
and U4997 (N_4997,N_3278,N_3179);
and U4998 (N_4998,N_3413,N_3090);
and U4999 (N_4999,N_3320,N_3356);
and U5000 (N_5000,N_4824,N_4275);
or U5001 (N_5001,N_4289,N_4148);
and U5002 (N_5002,N_4080,N_4225);
nand U5003 (N_5003,N_4995,N_4720);
nand U5004 (N_5004,N_4870,N_4169);
or U5005 (N_5005,N_4364,N_4372);
nor U5006 (N_5006,N_4749,N_4837);
nor U5007 (N_5007,N_4287,N_4729);
or U5008 (N_5008,N_4133,N_4307);
or U5009 (N_5009,N_4095,N_4861);
nand U5010 (N_5010,N_4213,N_4038);
and U5011 (N_5011,N_4697,N_4295);
and U5012 (N_5012,N_4081,N_4112);
xnor U5013 (N_5013,N_4486,N_4210);
and U5014 (N_5014,N_4231,N_4981);
and U5015 (N_5015,N_4355,N_4468);
or U5016 (N_5016,N_4279,N_4609);
nor U5017 (N_5017,N_4477,N_4363);
nand U5018 (N_5018,N_4379,N_4014);
and U5019 (N_5019,N_4554,N_4828);
nor U5020 (N_5020,N_4124,N_4844);
and U5021 (N_5021,N_4214,N_4751);
or U5022 (N_5022,N_4625,N_4181);
and U5023 (N_5023,N_4251,N_4574);
or U5024 (N_5024,N_4585,N_4805);
nand U5025 (N_5025,N_4977,N_4656);
and U5026 (N_5026,N_4202,N_4387);
xnor U5027 (N_5027,N_4943,N_4592);
nand U5028 (N_5028,N_4176,N_4551);
and U5029 (N_5029,N_4061,N_4817);
and U5030 (N_5030,N_4919,N_4332);
nor U5031 (N_5031,N_4780,N_4561);
nor U5032 (N_5032,N_4060,N_4209);
nand U5033 (N_5033,N_4791,N_4368);
nand U5034 (N_5034,N_4145,N_4555);
nand U5035 (N_5035,N_4036,N_4660);
or U5036 (N_5036,N_4352,N_4503);
and U5037 (N_5037,N_4796,N_4889);
and U5038 (N_5038,N_4255,N_4151);
nor U5039 (N_5039,N_4665,N_4727);
or U5040 (N_5040,N_4589,N_4342);
and U5041 (N_5041,N_4886,N_4435);
xnor U5042 (N_5042,N_4422,N_4630);
and U5043 (N_5043,N_4821,N_4733);
nor U5044 (N_5044,N_4264,N_4516);
or U5045 (N_5045,N_4705,N_4682);
nand U5046 (N_5046,N_4337,N_4678);
nor U5047 (N_5047,N_4427,N_4319);
xnor U5048 (N_5048,N_4167,N_4333);
and U5049 (N_5049,N_4783,N_4543);
or U5050 (N_5050,N_4960,N_4990);
nor U5051 (N_5051,N_4668,N_4715);
and U5052 (N_5052,N_4437,N_4107);
or U5053 (N_5053,N_4792,N_4182);
or U5054 (N_5054,N_4254,N_4766);
nor U5055 (N_5055,N_4966,N_4548);
or U5056 (N_5056,N_4021,N_4082);
nand U5057 (N_5057,N_4987,N_4451);
nand U5058 (N_5058,N_4536,N_4887);
xnor U5059 (N_5059,N_4381,N_4562);
nor U5060 (N_5060,N_4452,N_4146);
xor U5061 (N_5061,N_4747,N_4843);
xor U5062 (N_5062,N_4237,N_4568);
and U5063 (N_5063,N_4076,N_4166);
and U5064 (N_5064,N_4240,N_4773);
and U5065 (N_5065,N_4223,N_4161);
and U5066 (N_5066,N_4593,N_4522);
nor U5067 (N_5067,N_4501,N_4894);
nand U5068 (N_5068,N_4128,N_4612);
and U5069 (N_5069,N_4714,N_4748);
and U5070 (N_5070,N_4155,N_4219);
xor U5071 (N_5071,N_4587,N_4298);
nand U5072 (N_5072,N_4938,N_4511);
nor U5073 (N_5073,N_4781,N_4975);
nor U5074 (N_5074,N_4246,N_4073);
nand U5075 (N_5075,N_4144,N_4353);
xnor U5076 (N_5076,N_4417,N_4470);
nand U5077 (N_5077,N_4633,N_4542);
and U5078 (N_5078,N_4757,N_4496);
nor U5079 (N_5079,N_4461,N_4280);
and U5080 (N_5080,N_4928,N_4389);
nand U5081 (N_5081,N_4644,N_4183);
nor U5082 (N_5082,N_4921,N_4158);
xor U5083 (N_5083,N_4754,N_4740);
nor U5084 (N_5084,N_4838,N_4117);
nand U5085 (N_5085,N_4385,N_4827);
and U5086 (N_5086,N_4340,N_4680);
and U5087 (N_5087,N_4873,N_4839);
xor U5088 (N_5088,N_4926,N_4534);
xnor U5089 (N_5089,N_4573,N_4799);
nand U5090 (N_5090,N_4062,N_4495);
nand U5091 (N_5091,N_4359,N_4742);
nor U5092 (N_5092,N_4878,N_4027);
or U5093 (N_5093,N_4498,N_4002);
or U5094 (N_5094,N_4313,N_4911);
nand U5095 (N_5095,N_4200,N_4947);
and U5096 (N_5096,N_4136,N_4575);
nor U5097 (N_5097,N_4818,N_4604);
or U5098 (N_5098,N_4591,N_4642);
and U5099 (N_5099,N_4283,N_4635);
nor U5100 (N_5100,N_4616,N_4962);
nor U5101 (N_5101,N_4973,N_4518);
and U5102 (N_5102,N_4051,N_4063);
and U5103 (N_5103,N_4583,N_4043);
nor U5104 (N_5104,N_4737,N_4628);
xnor U5105 (N_5105,N_4147,N_4520);
and U5106 (N_5106,N_4571,N_4164);
and U5107 (N_5107,N_4508,N_4707);
and U5108 (N_5108,N_4758,N_4312);
nand U5109 (N_5109,N_4658,N_4946);
xor U5110 (N_5110,N_4929,N_4473);
nor U5111 (N_5111,N_4120,N_4111);
or U5112 (N_5112,N_4141,N_4872);
nor U5113 (N_5113,N_4034,N_4526);
or U5114 (N_5114,N_4205,N_4436);
or U5115 (N_5115,N_4106,N_4521);
nor U5116 (N_5116,N_4922,N_4681);
xnor U5117 (N_5117,N_4581,N_4489);
nand U5118 (N_5118,N_4343,N_4657);
and U5119 (N_5119,N_4101,N_4950);
and U5120 (N_5120,N_4341,N_4937);
nor U5121 (N_5121,N_4252,N_4457);
nand U5122 (N_5122,N_4345,N_4566);
and U5123 (N_5123,N_4853,N_4648);
nor U5124 (N_5124,N_4560,N_4150);
and U5125 (N_5125,N_4413,N_4908);
nand U5126 (N_5126,N_4299,N_4953);
xnor U5127 (N_5127,N_4001,N_4804);
and U5128 (N_5128,N_4645,N_4165);
and U5129 (N_5129,N_4218,N_4374);
or U5130 (N_5130,N_4813,N_4600);
or U5131 (N_5131,N_4685,N_4897);
and U5132 (N_5132,N_4309,N_4539);
nand U5133 (N_5133,N_4550,N_4188);
or U5134 (N_5134,N_4103,N_4208);
nand U5135 (N_5135,N_4003,N_4432);
nand U5136 (N_5136,N_4982,N_4916);
or U5137 (N_5137,N_4471,N_4540);
and U5138 (N_5138,N_4765,N_4871);
and U5139 (N_5139,N_4546,N_4663);
xor U5140 (N_5140,N_4857,N_4722);
nor U5141 (N_5141,N_4405,N_4260);
and U5142 (N_5142,N_4994,N_4371);
and U5143 (N_5143,N_4394,N_4541);
or U5144 (N_5144,N_4608,N_4607);
and U5145 (N_5145,N_4162,N_4986);
xor U5146 (N_5146,N_4819,N_4790);
nand U5147 (N_5147,N_4127,N_4849);
and U5148 (N_5148,N_4274,N_4721);
and U5149 (N_5149,N_4338,N_4528);
and U5150 (N_5150,N_4655,N_4867);
and U5151 (N_5151,N_4463,N_4402);
nand U5152 (N_5152,N_4549,N_4406);
and U5153 (N_5153,N_4807,N_4860);
nand U5154 (N_5154,N_4713,N_4241);
and U5155 (N_5155,N_4840,N_4132);
nor U5156 (N_5156,N_4653,N_4303);
or U5157 (N_5157,N_4997,N_4322);
or U5158 (N_5158,N_4472,N_4684);
and U5159 (N_5159,N_4841,N_4965);
nor U5160 (N_5160,N_4388,N_4315);
and U5161 (N_5161,N_4694,N_4375);
nand U5162 (N_5162,N_4494,N_4203);
nor U5163 (N_5163,N_4830,N_4085);
or U5164 (N_5164,N_4320,N_4438);
or U5165 (N_5165,N_4690,N_4369);
and U5166 (N_5166,N_4601,N_4925);
nand U5167 (N_5167,N_4090,N_4140);
nor U5168 (N_5168,N_4880,N_4940);
xnor U5169 (N_5169,N_4572,N_4440);
nand U5170 (N_5170,N_4262,N_4373);
nor U5171 (N_5171,N_4351,N_4448);
or U5172 (N_5172,N_4157,N_4410);
nor U5173 (N_5173,N_4492,N_4236);
nor U5174 (N_5174,N_4180,N_4088);
nor U5175 (N_5175,N_4286,N_4632);
or U5176 (N_5176,N_4877,N_4918);
or U5177 (N_5177,N_4178,N_4545);
nor U5178 (N_5178,N_4677,N_4057);
and U5179 (N_5179,N_4297,N_4445);
nand U5180 (N_5180,N_4171,N_4862);
or U5181 (N_5181,N_4497,N_4055);
and U5182 (N_5182,N_4578,N_4978);
nor U5183 (N_5183,N_4667,N_4614);
nand U5184 (N_5184,N_4285,N_4414);
or U5185 (N_5185,N_4365,N_4956);
or U5186 (N_5186,N_4970,N_4491);
nor U5187 (N_5187,N_4153,N_4250);
or U5188 (N_5188,N_4199,N_4779);
nand U5189 (N_5189,N_4687,N_4323);
xnor U5190 (N_5190,N_4408,N_4959);
nor U5191 (N_5191,N_4831,N_4113);
nor U5192 (N_5192,N_4895,N_4278);
or U5193 (N_5193,N_4618,N_4039);
nand U5194 (N_5194,N_4137,N_4070);
or U5195 (N_5195,N_4156,N_4458);
nor U5196 (N_5196,N_4159,N_4899);
nand U5197 (N_5197,N_4258,N_4464);
or U5198 (N_5198,N_4370,N_4504);
nor U5199 (N_5199,N_4048,N_4814);
or U5200 (N_5200,N_4400,N_4234);
and U5201 (N_5201,N_4961,N_4666);
nand U5202 (N_5202,N_4290,N_4755);
nand U5203 (N_5203,N_4294,N_4398);
or U5204 (N_5204,N_4671,N_4793);
and U5205 (N_5205,N_4746,N_4778);
nand U5206 (N_5206,N_4367,N_4594);
nand U5207 (N_5207,N_4130,N_4530);
or U5208 (N_5208,N_4196,N_4197);
and U5209 (N_5209,N_4305,N_4270);
xor U5210 (N_5210,N_4598,N_4265);
nand U5211 (N_5211,N_4788,N_4537);
nand U5212 (N_5212,N_4175,N_4361);
nor U5213 (N_5213,N_4505,N_4523);
nand U5214 (N_5214,N_4613,N_4932);
and U5215 (N_5215,N_4507,N_4386);
nor U5216 (N_5216,N_4634,N_4098);
and U5217 (N_5217,N_4775,N_4403);
nand U5218 (N_5218,N_4431,N_4524);
nor U5219 (N_5219,N_4776,N_4579);
or U5220 (N_5220,N_4430,N_4096);
nor U5221 (N_5221,N_4281,N_4753);
or U5222 (N_5222,N_4863,N_4704);
nor U5223 (N_5223,N_4756,N_4284);
and U5224 (N_5224,N_4193,N_4888);
nor U5225 (N_5225,N_4170,N_4446);
nor U5226 (N_5226,N_4514,N_4955);
nor U5227 (N_5227,N_4485,N_4292);
nand U5228 (N_5228,N_4915,N_4835);
and U5229 (N_5229,N_4099,N_4984);
nor U5230 (N_5230,N_4123,N_4669);
nand U5231 (N_5231,N_4611,N_4230);
and U5232 (N_5232,N_4570,N_4763);
nand U5233 (N_5233,N_4736,N_4703);
xnor U5234 (N_5234,N_4890,N_4211);
nand U5235 (N_5235,N_4967,N_4802);
nor U5236 (N_5236,N_4282,N_4565);
nor U5237 (N_5237,N_4009,N_4964);
and U5238 (N_5238,N_4875,N_4362);
xor U5239 (N_5239,N_4621,N_4806);
nor U5240 (N_5240,N_4903,N_4996);
nor U5241 (N_5241,N_4083,N_4808);
and U5242 (N_5242,N_4324,N_4544);
or U5243 (N_5243,N_4771,N_4177);
or U5244 (N_5244,N_4531,N_4856);
and U5245 (N_5245,N_4954,N_4893);
and U5246 (N_5246,N_4515,N_4606);
or U5247 (N_5247,N_4902,N_4479);
and U5248 (N_5248,N_4517,N_4212);
or U5249 (N_5249,N_4195,N_4772);
and U5250 (N_5250,N_4936,N_4941);
xor U5251 (N_5251,N_4138,N_4227);
nand U5252 (N_5252,N_4629,N_4590);
or U5253 (N_5253,N_4826,N_4045);
nor U5254 (N_5254,N_4344,N_4983);
and U5255 (N_5255,N_4253,N_4650);
nand U5256 (N_5256,N_4825,N_4909);
nor U5257 (N_5257,N_4006,N_4030);
or U5258 (N_5258,N_4078,N_4952);
xor U5259 (N_5259,N_4532,N_4268);
xor U5260 (N_5260,N_4718,N_4864);
nand U5261 (N_5261,N_4559,N_4493);
nand U5262 (N_5262,N_4993,N_4444);
nand U5263 (N_5263,N_4393,N_4288);
or U5264 (N_5264,N_4079,N_4201);
and U5265 (N_5265,N_4122,N_4011);
nor U5266 (N_5266,N_4698,N_4453);
or U5267 (N_5267,N_4226,N_4866);
nand U5268 (N_5268,N_4969,N_4163);
or U5269 (N_5269,N_4882,N_4968);
nand U5270 (N_5270,N_4067,N_4896);
nor U5271 (N_5271,N_4052,N_4249);
and U5272 (N_5272,N_4483,N_4071);
and U5273 (N_5273,N_4420,N_4846);
or U5274 (N_5274,N_4092,N_4269);
or U5275 (N_5275,N_4623,N_4743);
xor U5276 (N_5276,N_4366,N_4979);
and U5277 (N_5277,N_4416,N_4725);
nand U5278 (N_5278,N_4302,N_4421);
nand U5279 (N_5279,N_4519,N_4383);
and U5280 (N_5280,N_4951,N_4985);
and U5281 (N_5281,N_4640,N_4190);
or U5282 (N_5282,N_4024,N_4512);
xor U5283 (N_5283,N_4696,N_4626);
nand U5284 (N_5284,N_4649,N_4869);
and U5285 (N_5285,N_4118,N_4646);
xor U5286 (N_5286,N_4506,N_4321);
nand U5287 (N_5287,N_4091,N_4232);
xnor U5288 (N_5288,N_4812,N_4723);
or U5289 (N_5289,N_4104,N_4317);
nor U5290 (N_5290,N_4832,N_4441);
or U5291 (N_5291,N_4142,N_4971);
nor U5292 (N_5292,N_4917,N_4019);
nor U5293 (N_5293,N_4273,N_4418);
nand U5294 (N_5294,N_4741,N_4116);
nor U5295 (N_5295,N_4066,N_4750);
or U5296 (N_5296,N_4467,N_4032);
nand U5297 (N_5297,N_4901,N_4026);
or U5298 (N_5298,N_4046,N_4425);
xor U5299 (N_5299,N_4709,N_4168);
and U5300 (N_5300,N_4174,N_4016);
or U5301 (N_5301,N_4728,N_4850);
nand U5302 (N_5302,N_4336,N_4377);
or U5303 (N_5303,N_4056,N_4930);
nor U5304 (N_5304,N_4217,N_4731);
nor U5305 (N_5305,N_4538,N_4884);
nand U5306 (N_5306,N_4782,N_4459);
nor U5307 (N_5307,N_4025,N_4760);
nor U5308 (N_5308,N_4706,N_4712);
nand U5309 (N_5309,N_4291,N_4711);
nand U5310 (N_5310,N_4910,N_4851);
nand U5311 (N_5311,N_4325,N_4239);
xnor U5312 (N_5312,N_4624,N_4100);
or U5313 (N_5313,N_4272,N_4301);
and U5314 (N_5314,N_4786,N_4173);
or U5315 (N_5315,N_4378,N_4129);
nor U5316 (N_5316,N_4327,N_4848);
nand U5317 (N_5317,N_4350,N_4868);
and U5318 (N_5318,N_4474,N_4184);
or U5319 (N_5319,N_4194,N_4206);
nand U5320 (N_5320,N_4068,N_4801);
nor U5321 (N_5321,N_4636,N_4944);
nand U5322 (N_5322,N_4277,N_4789);
nor U5323 (N_5323,N_4639,N_4502);
xor U5324 (N_5324,N_4022,N_4881);
nand U5325 (N_5325,N_4018,N_4404);
nand U5326 (N_5326,N_4764,N_4439);
and U5327 (N_5327,N_4409,N_4296);
nand U5328 (N_5328,N_4029,N_4105);
nor U5329 (N_5329,N_4809,N_4466);
xor U5330 (N_5330,N_4300,N_4460);
or U5331 (N_5331,N_4401,N_4557);
nor U5332 (N_5332,N_4800,N_4109);
or U5333 (N_5333,N_4735,N_4077);
and U5334 (N_5334,N_4582,N_4724);
and U5335 (N_5335,N_4637,N_4415);
or U5336 (N_5336,N_4615,N_4007);
and U5337 (N_5337,N_4811,N_4834);
or U5338 (N_5338,N_4360,N_4072);
nand U5339 (N_5339,N_4035,N_4662);
and U5340 (N_5340,N_4610,N_4119);
or U5341 (N_5341,N_4186,N_4829);
nor U5342 (N_5342,N_4934,N_4115);
and U5343 (N_5343,N_4822,N_4509);
or U5344 (N_5344,N_4963,N_4094);
and U5345 (N_5345,N_4876,N_4883);
and U5346 (N_5346,N_4042,N_4752);
or U5347 (N_5347,N_4998,N_4126);
and U5348 (N_5348,N_4004,N_4823);
nand U5349 (N_5349,N_4093,N_4972);
nand U5350 (N_5350,N_4008,N_4510);
nand U5351 (N_5351,N_4267,N_4798);
and U5352 (N_5352,N_4652,N_4065);
nand U5353 (N_5353,N_4054,N_4500);
nor U5354 (N_5354,N_4716,N_4097);
or U5355 (N_5355,N_4031,N_4898);
or U5356 (N_5356,N_4139,N_4396);
or U5357 (N_5357,N_4795,N_4597);
and U5358 (N_5358,N_4980,N_4620);
or U5359 (N_5359,N_4143,N_4204);
nand U5360 (N_5360,N_4271,N_4328);
and U5361 (N_5361,N_4276,N_4859);
nor U5362 (N_5362,N_4040,N_4392);
or U5363 (N_5363,N_4058,N_4376);
nor U5364 (N_5364,N_4726,N_4412);
nand U5365 (N_5365,N_4121,N_4064);
nand U5366 (N_5366,N_4912,N_4084);
nand U5367 (N_5367,N_4647,N_4222);
nand U5368 (N_5368,N_4331,N_4033);
or U5369 (N_5369,N_4767,N_4957);
xor U5370 (N_5370,N_4248,N_4261);
nor U5371 (N_5371,N_4670,N_4777);
or U5372 (N_5372,N_4874,N_4855);
nand U5373 (N_5373,N_4339,N_4739);
and U5374 (N_5374,N_4044,N_4487);
or U5375 (N_5375,N_4391,N_4852);
or U5376 (N_5376,N_4905,N_4384);
nor U5377 (N_5377,N_4529,N_4738);
xor U5378 (N_5378,N_4689,N_4428);
or U5379 (N_5379,N_4481,N_4717);
nand U5380 (N_5380,N_4462,N_4224);
nand U5381 (N_5381,N_4395,N_4397);
nand U5382 (N_5382,N_4643,N_4257);
nand U5383 (N_5383,N_4047,N_4220);
and U5384 (N_5384,N_4945,N_4434);
or U5385 (N_5385,N_4759,N_4617);
nor U5386 (N_5386,N_4672,N_4664);
nor U5387 (N_5387,N_4564,N_4456);
or U5388 (N_5388,N_4089,N_4329);
nand U5389 (N_5389,N_4708,N_4683);
and U5390 (N_5390,N_4433,N_4619);
xor U5391 (N_5391,N_4216,N_4651);
nand U5392 (N_5392,N_4892,N_4484);
or U5393 (N_5393,N_4577,N_4730);
or U5394 (N_5394,N_4499,N_4160);
and U5395 (N_5395,N_4992,N_4885);
or U5396 (N_5396,N_4847,N_4074);
nor U5397 (N_5397,N_4335,N_4005);
nor U5398 (N_5398,N_4679,N_4854);
nand U5399 (N_5399,N_4797,N_4768);
and U5400 (N_5400,N_4049,N_4037);
and U5401 (N_5401,N_4306,N_4900);
or U5402 (N_5402,N_4675,N_4803);
and U5403 (N_5403,N_4075,N_4314);
and U5404 (N_5404,N_4215,N_4358);
nand U5405 (N_5405,N_4189,N_4920);
xnor U5406 (N_5406,N_4449,N_4935);
or U5407 (N_5407,N_4429,N_4794);
nor U5408 (N_5408,N_4482,N_4238);
nand U5409 (N_5409,N_4622,N_4556);
nand U5410 (N_5410,N_4599,N_4924);
and U5411 (N_5411,N_4816,N_4244);
and U5412 (N_5412,N_4447,N_4948);
nand U5413 (N_5413,N_4576,N_4357);
nor U5414 (N_5414,N_4185,N_4187);
nor U5415 (N_5415,N_4469,N_4235);
or U5416 (N_5416,N_4638,N_4923);
and U5417 (N_5417,N_4603,N_4784);
xnor U5418 (N_5418,N_4050,N_4013);
nand U5419 (N_5419,N_4426,N_4308);
xor U5420 (N_5420,N_4891,N_4787);
nor U5421 (N_5421,N_4247,N_4454);
and U5422 (N_5422,N_4602,N_4914);
nor U5423 (N_5423,N_4266,N_4933);
or U5424 (N_5424,N_4191,N_4131);
and U5425 (N_5425,N_4533,N_4527);
nand U5426 (N_5426,N_4567,N_4478);
nand U5427 (N_5427,N_4154,N_4242);
and U5428 (N_5428,N_4949,N_4192);
nor U5429 (N_5429,N_4991,N_4135);
nor U5430 (N_5430,N_4547,N_4349);
and U5431 (N_5431,N_4710,N_4488);
and U5432 (N_5432,N_4149,N_4179);
or U5433 (N_5433,N_4020,N_4348);
xor U5434 (N_5434,N_4927,N_4015);
nor U5435 (N_5435,N_4836,N_4525);
or U5436 (N_5436,N_4762,N_4087);
xor U5437 (N_5437,N_4419,N_4931);
or U5438 (N_5438,N_4659,N_4326);
or U5439 (N_5439,N_4976,N_4688);
and U5440 (N_5440,N_4693,N_4442);
nor U5441 (N_5441,N_4745,N_4734);
or U5442 (N_5442,N_4017,N_4553);
and U5443 (N_5443,N_4198,N_4334);
nand U5444 (N_5444,N_4086,N_4152);
nand U5445 (N_5445,N_4761,N_4588);
and U5446 (N_5446,N_4913,N_4311);
xnor U5447 (N_5447,N_4380,N_4785);
and U5448 (N_5448,N_4356,N_4631);
and U5449 (N_5449,N_4347,N_4586);
and U5450 (N_5450,N_4465,N_4535);
and U5451 (N_5451,N_4661,N_4233);
and U5452 (N_5452,N_4480,N_4207);
nor U5453 (N_5453,N_4407,N_4134);
and U5454 (N_5454,N_4641,N_4263);
and U5455 (N_5455,N_4382,N_4125);
or U5456 (N_5456,N_4700,N_4108);
nand U5457 (N_5457,N_4810,N_4774);
and U5458 (N_5458,N_4833,N_4455);
xnor U5459 (N_5459,N_4490,N_4842);
nor U5460 (N_5460,N_4221,N_4069);
or U5461 (N_5461,N_4000,N_4411);
nor U5462 (N_5462,N_4310,N_4702);
and U5463 (N_5463,N_4939,N_4744);
nor U5464 (N_5464,N_4845,N_4595);
nor U5465 (N_5465,N_4475,N_4988);
nor U5466 (N_5466,N_4041,N_4513);
nand U5467 (N_5467,N_4563,N_4243);
or U5468 (N_5468,N_4330,N_4691);
nor U5469 (N_5469,N_4974,N_4906);
xnor U5470 (N_5470,N_4569,N_4695);
or U5471 (N_5471,N_4865,N_4102);
xnor U5472 (N_5472,N_4450,N_4770);
xor U5473 (N_5473,N_4686,N_4701);
and U5474 (N_5474,N_4390,N_4674);
nand U5475 (N_5475,N_4318,N_4989);
or U5476 (N_5476,N_4584,N_4858);
nand U5477 (N_5477,N_4399,N_4354);
and U5478 (N_5478,N_4423,N_4879);
xor U5479 (N_5479,N_4605,N_4654);
nor U5480 (N_5480,N_4627,N_4012);
or U5481 (N_5481,N_4259,N_4053);
and U5482 (N_5482,N_4304,N_4476);
xnor U5483 (N_5483,N_4346,N_4059);
nand U5484 (N_5484,N_4719,N_4228);
and U5485 (N_5485,N_4676,N_4958);
and U5486 (N_5486,N_4942,N_4229);
or U5487 (N_5487,N_4256,N_4110);
and U5488 (N_5488,N_4820,N_4023);
nor U5489 (N_5489,N_4172,N_4245);
and U5490 (N_5490,N_4552,N_4443);
and U5491 (N_5491,N_4316,N_4028);
or U5492 (N_5492,N_4999,N_4424);
or U5493 (N_5493,N_4114,N_4692);
or U5494 (N_5494,N_4580,N_4293);
xor U5495 (N_5495,N_4904,N_4596);
xnor U5496 (N_5496,N_4673,N_4699);
xnor U5497 (N_5497,N_4907,N_4010);
and U5498 (N_5498,N_4558,N_4769);
xor U5499 (N_5499,N_4815,N_4732);
and U5500 (N_5500,N_4153,N_4734);
or U5501 (N_5501,N_4598,N_4044);
and U5502 (N_5502,N_4919,N_4355);
nor U5503 (N_5503,N_4556,N_4834);
xnor U5504 (N_5504,N_4417,N_4450);
nor U5505 (N_5505,N_4151,N_4011);
and U5506 (N_5506,N_4069,N_4144);
nand U5507 (N_5507,N_4801,N_4390);
nand U5508 (N_5508,N_4308,N_4228);
and U5509 (N_5509,N_4052,N_4692);
and U5510 (N_5510,N_4336,N_4926);
nor U5511 (N_5511,N_4327,N_4679);
nand U5512 (N_5512,N_4341,N_4164);
nor U5513 (N_5513,N_4892,N_4913);
and U5514 (N_5514,N_4947,N_4045);
and U5515 (N_5515,N_4988,N_4730);
xor U5516 (N_5516,N_4655,N_4188);
or U5517 (N_5517,N_4371,N_4901);
nand U5518 (N_5518,N_4434,N_4279);
nor U5519 (N_5519,N_4262,N_4341);
nor U5520 (N_5520,N_4467,N_4864);
and U5521 (N_5521,N_4248,N_4555);
or U5522 (N_5522,N_4320,N_4441);
or U5523 (N_5523,N_4080,N_4837);
nand U5524 (N_5524,N_4321,N_4606);
nand U5525 (N_5525,N_4719,N_4518);
nand U5526 (N_5526,N_4353,N_4444);
and U5527 (N_5527,N_4480,N_4814);
or U5528 (N_5528,N_4290,N_4090);
and U5529 (N_5529,N_4430,N_4225);
nand U5530 (N_5530,N_4126,N_4921);
or U5531 (N_5531,N_4779,N_4411);
and U5532 (N_5532,N_4521,N_4764);
nand U5533 (N_5533,N_4633,N_4657);
and U5534 (N_5534,N_4031,N_4498);
nand U5535 (N_5535,N_4216,N_4988);
nand U5536 (N_5536,N_4751,N_4853);
nor U5537 (N_5537,N_4958,N_4077);
xnor U5538 (N_5538,N_4576,N_4676);
and U5539 (N_5539,N_4247,N_4693);
and U5540 (N_5540,N_4650,N_4213);
or U5541 (N_5541,N_4825,N_4600);
nand U5542 (N_5542,N_4003,N_4645);
xnor U5543 (N_5543,N_4952,N_4189);
and U5544 (N_5544,N_4242,N_4492);
nor U5545 (N_5545,N_4167,N_4799);
or U5546 (N_5546,N_4733,N_4772);
and U5547 (N_5547,N_4489,N_4013);
and U5548 (N_5548,N_4181,N_4131);
and U5549 (N_5549,N_4124,N_4157);
and U5550 (N_5550,N_4117,N_4076);
nand U5551 (N_5551,N_4514,N_4932);
nand U5552 (N_5552,N_4078,N_4548);
xnor U5553 (N_5553,N_4865,N_4367);
or U5554 (N_5554,N_4707,N_4466);
or U5555 (N_5555,N_4420,N_4443);
and U5556 (N_5556,N_4892,N_4044);
or U5557 (N_5557,N_4650,N_4032);
and U5558 (N_5558,N_4720,N_4104);
and U5559 (N_5559,N_4987,N_4664);
nor U5560 (N_5560,N_4429,N_4371);
nand U5561 (N_5561,N_4345,N_4987);
xor U5562 (N_5562,N_4597,N_4057);
xor U5563 (N_5563,N_4274,N_4483);
nand U5564 (N_5564,N_4568,N_4343);
nand U5565 (N_5565,N_4989,N_4716);
and U5566 (N_5566,N_4949,N_4269);
nand U5567 (N_5567,N_4194,N_4510);
nor U5568 (N_5568,N_4542,N_4389);
nand U5569 (N_5569,N_4262,N_4745);
or U5570 (N_5570,N_4133,N_4046);
or U5571 (N_5571,N_4890,N_4016);
nor U5572 (N_5572,N_4910,N_4970);
xnor U5573 (N_5573,N_4462,N_4939);
or U5574 (N_5574,N_4854,N_4685);
and U5575 (N_5575,N_4876,N_4965);
or U5576 (N_5576,N_4781,N_4013);
and U5577 (N_5577,N_4952,N_4235);
nand U5578 (N_5578,N_4480,N_4602);
or U5579 (N_5579,N_4687,N_4915);
nand U5580 (N_5580,N_4206,N_4125);
and U5581 (N_5581,N_4782,N_4928);
and U5582 (N_5582,N_4340,N_4215);
nor U5583 (N_5583,N_4868,N_4316);
and U5584 (N_5584,N_4233,N_4645);
nor U5585 (N_5585,N_4261,N_4166);
or U5586 (N_5586,N_4292,N_4386);
nor U5587 (N_5587,N_4124,N_4211);
nor U5588 (N_5588,N_4454,N_4530);
and U5589 (N_5589,N_4696,N_4524);
and U5590 (N_5590,N_4502,N_4834);
nand U5591 (N_5591,N_4454,N_4727);
nor U5592 (N_5592,N_4466,N_4214);
and U5593 (N_5593,N_4847,N_4216);
and U5594 (N_5594,N_4851,N_4999);
and U5595 (N_5595,N_4564,N_4105);
xnor U5596 (N_5596,N_4371,N_4117);
nor U5597 (N_5597,N_4998,N_4718);
nand U5598 (N_5598,N_4652,N_4223);
and U5599 (N_5599,N_4700,N_4262);
xnor U5600 (N_5600,N_4370,N_4218);
or U5601 (N_5601,N_4313,N_4315);
nor U5602 (N_5602,N_4941,N_4142);
and U5603 (N_5603,N_4746,N_4536);
nor U5604 (N_5604,N_4916,N_4246);
or U5605 (N_5605,N_4485,N_4416);
nor U5606 (N_5606,N_4124,N_4904);
nand U5607 (N_5607,N_4555,N_4670);
nor U5608 (N_5608,N_4473,N_4518);
and U5609 (N_5609,N_4194,N_4455);
nand U5610 (N_5610,N_4432,N_4885);
nand U5611 (N_5611,N_4825,N_4726);
nor U5612 (N_5612,N_4269,N_4551);
and U5613 (N_5613,N_4363,N_4580);
or U5614 (N_5614,N_4301,N_4494);
nand U5615 (N_5615,N_4864,N_4398);
nor U5616 (N_5616,N_4593,N_4306);
and U5617 (N_5617,N_4191,N_4821);
nor U5618 (N_5618,N_4304,N_4788);
nor U5619 (N_5619,N_4681,N_4701);
nor U5620 (N_5620,N_4502,N_4686);
or U5621 (N_5621,N_4587,N_4096);
or U5622 (N_5622,N_4430,N_4375);
nor U5623 (N_5623,N_4081,N_4299);
nand U5624 (N_5624,N_4792,N_4989);
and U5625 (N_5625,N_4411,N_4437);
and U5626 (N_5626,N_4218,N_4608);
or U5627 (N_5627,N_4584,N_4863);
nand U5628 (N_5628,N_4268,N_4888);
nand U5629 (N_5629,N_4817,N_4377);
xnor U5630 (N_5630,N_4511,N_4094);
or U5631 (N_5631,N_4109,N_4607);
and U5632 (N_5632,N_4068,N_4484);
or U5633 (N_5633,N_4272,N_4403);
xor U5634 (N_5634,N_4327,N_4872);
or U5635 (N_5635,N_4030,N_4045);
or U5636 (N_5636,N_4848,N_4260);
and U5637 (N_5637,N_4973,N_4270);
nor U5638 (N_5638,N_4466,N_4653);
or U5639 (N_5639,N_4559,N_4947);
nand U5640 (N_5640,N_4261,N_4701);
or U5641 (N_5641,N_4578,N_4169);
nor U5642 (N_5642,N_4161,N_4606);
nand U5643 (N_5643,N_4484,N_4153);
nor U5644 (N_5644,N_4061,N_4660);
nand U5645 (N_5645,N_4319,N_4324);
nand U5646 (N_5646,N_4332,N_4501);
or U5647 (N_5647,N_4771,N_4816);
nand U5648 (N_5648,N_4752,N_4543);
nand U5649 (N_5649,N_4011,N_4428);
nand U5650 (N_5650,N_4046,N_4250);
and U5651 (N_5651,N_4682,N_4226);
or U5652 (N_5652,N_4068,N_4332);
and U5653 (N_5653,N_4669,N_4618);
xor U5654 (N_5654,N_4941,N_4938);
nor U5655 (N_5655,N_4238,N_4211);
or U5656 (N_5656,N_4103,N_4052);
nand U5657 (N_5657,N_4196,N_4171);
nand U5658 (N_5658,N_4281,N_4713);
xor U5659 (N_5659,N_4489,N_4086);
and U5660 (N_5660,N_4485,N_4244);
nand U5661 (N_5661,N_4264,N_4286);
xor U5662 (N_5662,N_4822,N_4883);
nor U5663 (N_5663,N_4359,N_4798);
nor U5664 (N_5664,N_4723,N_4393);
nand U5665 (N_5665,N_4432,N_4251);
and U5666 (N_5666,N_4795,N_4872);
and U5667 (N_5667,N_4406,N_4650);
or U5668 (N_5668,N_4705,N_4622);
nand U5669 (N_5669,N_4641,N_4941);
nand U5670 (N_5670,N_4772,N_4451);
xnor U5671 (N_5671,N_4634,N_4337);
nand U5672 (N_5672,N_4008,N_4944);
and U5673 (N_5673,N_4983,N_4918);
and U5674 (N_5674,N_4397,N_4527);
or U5675 (N_5675,N_4748,N_4414);
and U5676 (N_5676,N_4380,N_4186);
nand U5677 (N_5677,N_4800,N_4225);
nand U5678 (N_5678,N_4953,N_4866);
and U5679 (N_5679,N_4704,N_4614);
and U5680 (N_5680,N_4525,N_4117);
nand U5681 (N_5681,N_4569,N_4841);
xor U5682 (N_5682,N_4774,N_4601);
xnor U5683 (N_5683,N_4611,N_4970);
nand U5684 (N_5684,N_4820,N_4626);
nand U5685 (N_5685,N_4154,N_4189);
and U5686 (N_5686,N_4787,N_4893);
or U5687 (N_5687,N_4390,N_4065);
and U5688 (N_5688,N_4797,N_4478);
nand U5689 (N_5689,N_4660,N_4818);
nand U5690 (N_5690,N_4866,N_4410);
nor U5691 (N_5691,N_4436,N_4281);
or U5692 (N_5692,N_4861,N_4859);
or U5693 (N_5693,N_4763,N_4305);
nor U5694 (N_5694,N_4017,N_4293);
or U5695 (N_5695,N_4586,N_4890);
or U5696 (N_5696,N_4908,N_4313);
nand U5697 (N_5697,N_4139,N_4138);
nand U5698 (N_5698,N_4626,N_4708);
nor U5699 (N_5699,N_4304,N_4925);
and U5700 (N_5700,N_4928,N_4078);
xnor U5701 (N_5701,N_4273,N_4000);
or U5702 (N_5702,N_4185,N_4752);
nor U5703 (N_5703,N_4598,N_4905);
or U5704 (N_5704,N_4635,N_4803);
xnor U5705 (N_5705,N_4529,N_4994);
and U5706 (N_5706,N_4581,N_4151);
nand U5707 (N_5707,N_4002,N_4646);
nor U5708 (N_5708,N_4630,N_4498);
and U5709 (N_5709,N_4966,N_4424);
xnor U5710 (N_5710,N_4176,N_4607);
nor U5711 (N_5711,N_4973,N_4045);
or U5712 (N_5712,N_4518,N_4036);
or U5713 (N_5713,N_4259,N_4566);
and U5714 (N_5714,N_4542,N_4378);
nor U5715 (N_5715,N_4002,N_4839);
nor U5716 (N_5716,N_4536,N_4567);
nor U5717 (N_5717,N_4518,N_4437);
nor U5718 (N_5718,N_4981,N_4110);
nand U5719 (N_5719,N_4016,N_4193);
and U5720 (N_5720,N_4258,N_4281);
nand U5721 (N_5721,N_4808,N_4515);
or U5722 (N_5722,N_4983,N_4376);
or U5723 (N_5723,N_4240,N_4340);
nand U5724 (N_5724,N_4654,N_4486);
nor U5725 (N_5725,N_4303,N_4927);
and U5726 (N_5726,N_4426,N_4915);
nor U5727 (N_5727,N_4444,N_4905);
or U5728 (N_5728,N_4558,N_4776);
nor U5729 (N_5729,N_4346,N_4573);
xor U5730 (N_5730,N_4637,N_4767);
xor U5731 (N_5731,N_4468,N_4753);
or U5732 (N_5732,N_4404,N_4142);
nand U5733 (N_5733,N_4321,N_4137);
nand U5734 (N_5734,N_4700,N_4207);
nand U5735 (N_5735,N_4316,N_4563);
nand U5736 (N_5736,N_4019,N_4921);
xor U5737 (N_5737,N_4825,N_4766);
nand U5738 (N_5738,N_4280,N_4348);
or U5739 (N_5739,N_4673,N_4143);
and U5740 (N_5740,N_4097,N_4516);
and U5741 (N_5741,N_4738,N_4586);
nor U5742 (N_5742,N_4462,N_4920);
and U5743 (N_5743,N_4256,N_4112);
nand U5744 (N_5744,N_4321,N_4374);
or U5745 (N_5745,N_4818,N_4980);
nor U5746 (N_5746,N_4976,N_4768);
and U5747 (N_5747,N_4636,N_4919);
or U5748 (N_5748,N_4424,N_4303);
nand U5749 (N_5749,N_4306,N_4029);
xor U5750 (N_5750,N_4547,N_4515);
nor U5751 (N_5751,N_4026,N_4977);
nand U5752 (N_5752,N_4984,N_4489);
xor U5753 (N_5753,N_4208,N_4899);
and U5754 (N_5754,N_4139,N_4441);
nand U5755 (N_5755,N_4384,N_4162);
or U5756 (N_5756,N_4850,N_4533);
or U5757 (N_5757,N_4654,N_4311);
nor U5758 (N_5758,N_4327,N_4746);
and U5759 (N_5759,N_4249,N_4708);
nor U5760 (N_5760,N_4373,N_4539);
and U5761 (N_5761,N_4726,N_4451);
nand U5762 (N_5762,N_4407,N_4085);
nand U5763 (N_5763,N_4848,N_4285);
and U5764 (N_5764,N_4856,N_4013);
nor U5765 (N_5765,N_4856,N_4213);
nor U5766 (N_5766,N_4038,N_4345);
or U5767 (N_5767,N_4048,N_4063);
nand U5768 (N_5768,N_4422,N_4436);
nor U5769 (N_5769,N_4670,N_4066);
or U5770 (N_5770,N_4417,N_4228);
or U5771 (N_5771,N_4644,N_4135);
and U5772 (N_5772,N_4236,N_4850);
and U5773 (N_5773,N_4303,N_4536);
nand U5774 (N_5774,N_4696,N_4148);
xnor U5775 (N_5775,N_4503,N_4877);
nor U5776 (N_5776,N_4946,N_4197);
nand U5777 (N_5777,N_4912,N_4567);
and U5778 (N_5778,N_4484,N_4601);
or U5779 (N_5779,N_4572,N_4401);
xnor U5780 (N_5780,N_4215,N_4671);
nand U5781 (N_5781,N_4903,N_4573);
or U5782 (N_5782,N_4089,N_4371);
or U5783 (N_5783,N_4413,N_4797);
nand U5784 (N_5784,N_4595,N_4483);
nand U5785 (N_5785,N_4825,N_4454);
or U5786 (N_5786,N_4410,N_4562);
nand U5787 (N_5787,N_4469,N_4641);
and U5788 (N_5788,N_4948,N_4745);
and U5789 (N_5789,N_4745,N_4910);
or U5790 (N_5790,N_4295,N_4419);
nor U5791 (N_5791,N_4828,N_4343);
or U5792 (N_5792,N_4469,N_4596);
nor U5793 (N_5793,N_4642,N_4317);
nor U5794 (N_5794,N_4677,N_4731);
nand U5795 (N_5795,N_4077,N_4751);
nand U5796 (N_5796,N_4444,N_4884);
or U5797 (N_5797,N_4855,N_4314);
xor U5798 (N_5798,N_4677,N_4699);
nor U5799 (N_5799,N_4567,N_4910);
nor U5800 (N_5800,N_4026,N_4560);
nand U5801 (N_5801,N_4663,N_4013);
xnor U5802 (N_5802,N_4657,N_4814);
xnor U5803 (N_5803,N_4608,N_4042);
or U5804 (N_5804,N_4563,N_4728);
or U5805 (N_5805,N_4481,N_4785);
nor U5806 (N_5806,N_4511,N_4957);
nand U5807 (N_5807,N_4548,N_4815);
and U5808 (N_5808,N_4226,N_4382);
nor U5809 (N_5809,N_4901,N_4699);
or U5810 (N_5810,N_4404,N_4807);
or U5811 (N_5811,N_4061,N_4433);
or U5812 (N_5812,N_4699,N_4943);
nor U5813 (N_5813,N_4870,N_4276);
nand U5814 (N_5814,N_4698,N_4711);
and U5815 (N_5815,N_4343,N_4235);
nor U5816 (N_5816,N_4330,N_4723);
nor U5817 (N_5817,N_4388,N_4911);
nor U5818 (N_5818,N_4217,N_4757);
nor U5819 (N_5819,N_4410,N_4849);
nand U5820 (N_5820,N_4637,N_4001);
nor U5821 (N_5821,N_4196,N_4105);
or U5822 (N_5822,N_4790,N_4257);
nor U5823 (N_5823,N_4502,N_4271);
or U5824 (N_5824,N_4053,N_4697);
nand U5825 (N_5825,N_4694,N_4624);
nand U5826 (N_5826,N_4167,N_4260);
nand U5827 (N_5827,N_4359,N_4490);
and U5828 (N_5828,N_4770,N_4230);
xnor U5829 (N_5829,N_4175,N_4384);
nand U5830 (N_5830,N_4966,N_4095);
nand U5831 (N_5831,N_4232,N_4791);
nor U5832 (N_5832,N_4100,N_4745);
or U5833 (N_5833,N_4595,N_4930);
nand U5834 (N_5834,N_4310,N_4434);
and U5835 (N_5835,N_4965,N_4175);
xor U5836 (N_5836,N_4461,N_4595);
nor U5837 (N_5837,N_4442,N_4262);
or U5838 (N_5838,N_4684,N_4923);
nand U5839 (N_5839,N_4170,N_4532);
or U5840 (N_5840,N_4305,N_4268);
or U5841 (N_5841,N_4675,N_4126);
nor U5842 (N_5842,N_4782,N_4044);
or U5843 (N_5843,N_4118,N_4250);
or U5844 (N_5844,N_4219,N_4707);
or U5845 (N_5845,N_4200,N_4986);
and U5846 (N_5846,N_4752,N_4115);
nand U5847 (N_5847,N_4029,N_4864);
nand U5848 (N_5848,N_4595,N_4835);
nand U5849 (N_5849,N_4676,N_4090);
or U5850 (N_5850,N_4362,N_4419);
nor U5851 (N_5851,N_4679,N_4696);
or U5852 (N_5852,N_4645,N_4479);
and U5853 (N_5853,N_4970,N_4172);
nand U5854 (N_5854,N_4787,N_4618);
nor U5855 (N_5855,N_4011,N_4740);
or U5856 (N_5856,N_4724,N_4487);
and U5857 (N_5857,N_4877,N_4030);
or U5858 (N_5858,N_4156,N_4494);
nand U5859 (N_5859,N_4572,N_4474);
nand U5860 (N_5860,N_4664,N_4233);
or U5861 (N_5861,N_4459,N_4426);
or U5862 (N_5862,N_4962,N_4827);
nor U5863 (N_5863,N_4057,N_4649);
xor U5864 (N_5864,N_4826,N_4262);
and U5865 (N_5865,N_4107,N_4064);
nor U5866 (N_5866,N_4914,N_4339);
or U5867 (N_5867,N_4241,N_4773);
xor U5868 (N_5868,N_4962,N_4289);
nand U5869 (N_5869,N_4016,N_4670);
nor U5870 (N_5870,N_4169,N_4999);
nor U5871 (N_5871,N_4630,N_4516);
xor U5872 (N_5872,N_4473,N_4958);
and U5873 (N_5873,N_4834,N_4194);
and U5874 (N_5874,N_4361,N_4737);
and U5875 (N_5875,N_4619,N_4462);
nand U5876 (N_5876,N_4004,N_4998);
xnor U5877 (N_5877,N_4692,N_4471);
nand U5878 (N_5878,N_4738,N_4102);
or U5879 (N_5879,N_4818,N_4734);
nand U5880 (N_5880,N_4662,N_4793);
nor U5881 (N_5881,N_4925,N_4744);
nor U5882 (N_5882,N_4672,N_4614);
and U5883 (N_5883,N_4683,N_4218);
nor U5884 (N_5884,N_4824,N_4108);
nor U5885 (N_5885,N_4322,N_4844);
nand U5886 (N_5886,N_4166,N_4960);
xor U5887 (N_5887,N_4419,N_4397);
and U5888 (N_5888,N_4304,N_4746);
nand U5889 (N_5889,N_4748,N_4615);
nor U5890 (N_5890,N_4555,N_4235);
and U5891 (N_5891,N_4513,N_4299);
xor U5892 (N_5892,N_4747,N_4388);
and U5893 (N_5893,N_4851,N_4799);
xor U5894 (N_5894,N_4762,N_4782);
nand U5895 (N_5895,N_4991,N_4165);
nor U5896 (N_5896,N_4799,N_4419);
and U5897 (N_5897,N_4332,N_4450);
nand U5898 (N_5898,N_4447,N_4794);
nand U5899 (N_5899,N_4419,N_4867);
nor U5900 (N_5900,N_4098,N_4304);
and U5901 (N_5901,N_4112,N_4752);
xnor U5902 (N_5902,N_4423,N_4726);
nor U5903 (N_5903,N_4435,N_4176);
nor U5904 (N_5904,N_4544,N_4439);
xnor U5905 (N_5905,N_4044,N_4909);
and U5906 (N_5906,N_4292,N_4776);
nand U5907 (N_5907,N_4091,N_4384);
nand U5908 (N_5908,N_4282,N_4853);
or U5909 (N_5909,N_4485,N_4006);
or U5910 (N_5910,N_4540,N_4599);
nor U5911 (N_5911,N_4348,N_4568);
nand U5912 (N_5912,N_4767,N_4800);
or U5913 (N_5913,N_4480,N_4106);
nor U5914 (N_5914,N_4845,N_4795);
or U5915 (N_5915,N_4797,N_4829);
and U5916 (N_5916,N_4034,N_4792);
or U5917 (N_5917,N_4078,N_4008);
nand U5918 (N_5918,N_4903,N_4134);
nor U5919 (N_5919,N_4204,N_4731);
nor U5920 (N_5920,N_4055,N_4122);
nor U5921 (N_5921,N_4713,N_4396);
nor U5922 (N_5922,N_4297,N_4600);
xnor U5923 (N_5923,N_4093,N_4123);
or U5924 (N_5924,N_4144,N_4687);
nand U5925 (N_5925,N_4187,N_4767);
or U5926 (N_5926,N_4666,N_4634);
and U5927 (N_5927,N_4507,N_4317);
xnor U5928 (N_5928,N_4259,N_4945);
and U5929 (N_5929,N_4786,N_4590);
and U5930 (N_5930,N_4930,N_4537);
xnor U5931 (N_5931,N_4758,N_4242);
nand U5932 (N_5932,N_4667,N_4841);
nor U5933 (N_5933,N_4124,N_4554);
nor U5934 (N_5934,N_4773,N_4823);
nor U5935 (N_5935,N_4896,N_4389);
or U5936 (N_5936,N_4922,N_4224);
nand U5937 (N_5937,N_4821,N_4227);
or U5938 (N_5938,N_4978,N_4544);
or U5939 (N_5939,N_4893,N_4915);
xnor U5940 (N_5940,N_4614,N_4246);
nand U5941 (N_5941,N_4907,N_4444);
and U5942 (N_5942,N_4933,N_4641);
or U5943 (N_5943,N_4477,N_4729);
nor U5944 (N_5944,N_4268,N_4738);
nor U5945 (N_5945,N_4759,N_4264);
or U5946 (N_5946,N_4820,N_4954);
xor U5947 (N_5947,N_4042,N_4162);
or U5948 (N_5948,N_4476,N_4012);
and U5949 (N_5949,N_4680,N_4297);
nand U5950 (N_5950,N_4153,N_4796);
nand U5951 (N_5951,N_4305,N_4349);
and U5952 (N_5952,N_4012,N_4862);
or U5953 (N_5953,N_4988,N_4962);
nor U5954 (N_5954,N_4606,N_4243);
nand U5955 (N_5955,N_4610,N_4601);
or U5956 (N_5956,N_4822,N_4184);
nor U5957 (N_5957,N_4994,N_4336);
or U5958 (N_5958,N_4536,N_4149);
nand U5959 (N_5959,N_4465,N_4044);
or U5960 (N_5960,N_4228,N_4478);
or U5961 (N_5961,N_4363,N_4092);
xor U5962 (N_5962,N_4681,N_4580);
nor U5963 (N_5963,N_4962,N_4295);
nor U5964 (N_5964,N_4365,N_4790);
nor U5965 (N_5965,N_4948,N_4797);
or U5966 (N_5966,N_4189,N_4486);
nor U5967 (N_5967,N_4395,N_4496);
or U5968 (N_5968,N_4368,N_4317);
or U5969 (N_5969,N_4491,N_4359);
or U5970 (N_5970,N_4581,N_4414);
xor U5971 (N_5971,N_4993,N_4631);
or U5972 (N_5972,N_4490,N_4996);
or U5973 (N_5973,N_4068,N_4284);
and U5974 (N_5974,N_4356,N_4589);
nand U5975 (N_5975,N_4134,N_4436);
and U5976 (N_5976,N_4140,N_4299);
or U5977 (N_5977,N_4263,N_4717);
xnor U5978 (N_5978,N_4520,N_4346);
or U5979 (N_5979,N_4383,N_4409);
and U5980 (N_5980,N_4155,N_4800);
nor U5981 (N_5981,N_4294,N_4529);
and U5982 (N_5982,N_4648,N_4150);
or U5983 (N_5983,N_4141,N_4310);
nor U5984 (N_5984,N_4182,N_4810);
and U5985 (N_5985,N_4688,N_4828);
nor U5986 (N_5986,N_4096,N_4717);
or U5987 (N_5987,N_4286,N_4130);
xor U5988 (N_5988,N_4768,N_4912);
or U5989 (N_5989,N_4430,N_4871);
nand U5990 (N_5990,N_4975,N_4441);
or U5991 (N_5991,N_4948,N_4803);
nand U5992 (N_5992,N_4593,N_4311);
and U5993 (N_5993,N_4040,N_4068);
nand U5994 (N_5994,N_4138,N_4836);
nor U5995 (N_5995,N_4121,N_4915);
and U5996 (N_5996,N_4621,N_4423);
nand U5997 (N_5997,N_4488,N_4682);
nor U5998 (N_5998,N_4787,N_4272);
xor U5999 (N_5999,N_4351,N_4647);
nor U6000 (N_6000,N_5716,N_5012);
nor U6001 (N_6001,N_5817,N_5478);
nand U6002 (N_6002,N_5027,N_5700);
or U6003 (N_6003,N_5321,N_5009);
or U6004 (N_6004,N_5853,N_5756);
and U6005 (N_6005,N_5025,N_5753);
xor U6006 (N_6006,N_5726,N_5952);
nand U6007 (N_6007,N_5649,N_5326);
nand U6008 (N_6008,N_5650,N_5579);
nand U6009 (N_6009,N_5619,N_5112);
nand U6010 (N_6010,N_5209,N_5384);
or U6011 (N_6011,N_5354,N_5253);
nand U6012 (N_6012,N_5260,N_5658);
and U6013 (N_6013,N_5486,N_5656);
nor U6014 (N_6014,N_5095,N_5448);
xor U6015 (N_6015,N_5154,N_5856);
xor U6016 (N_6016,N_5087,N_5008);
nand U6017 (N_6017,N_5996,N_5862);
nor U6018 (N_6018,N_5134,N_5876);
or U6019 (N_6019,N_5231,N_5606);
and U6020 (N_6020,N_5484,N_5139);
nor U6021 (N_6021,N_5600,N_5452);
and U6022 (N_6022,N_5526,N_5041);
nor U6023 (N_6023,N_5084,N_5802);
nor U6024 (N_6024,N_5307,N_5320);
nand U6025 (N_6025,N_5908,N_5182);
xor U6026 (N_6026,N_5325,N_5786);
or U6027 (N_6027,N_5050,N_5754);
and U6028 (N_6028,N_5052,N_5133);
xor U6029 (N_6029,N_5235,N_5468);
nand U6030 (N_6030,N_5106,N_5504);
or U6031 (N_6031,N_5705,N_5437);
and U6032 (N_6032,N_5516,N_5064);
and U6033 (N_6033,N_5434,N_5854);
nand U6034 (N_6034,N_5415,N_5159);
and U6035 (N_6035,N_5342,N_5114);
xnor U6036 (N_6036,N_5568,N_5599);
or U6037 (N_6037,N_5919,N_5279);
and U6038 (N_6038,N_5233,N_5038);
nand U6039 (N_6039,N_5271,N_5804);
and U6040 (N_6040,N_5790,N_5687);
nand U6041 (N_6041,N_5450,N_5514);
nor U6042 (N_6042,N_5751,N_5183);
or U6043 (N_6043,N_5546,N_5783);
nor U6044 (N_6044,N_5000,N_5418);
nand U6045 (N_6045,N_5735,N_5944);
or U6046 (N_6046,N_5767,N_5607);
nor U6047 (N_6047,N_5480,N_5595);
xor U6048 (N_6048,N_5282,N_5147);
or U6049 (N_6049,N_5832,N_5822);
and U6050 (N_6050,N_5552,N_5356);
or U6051 (N_6051,N_5380,N_5160);
xor U6052 (N_6052,N_5058,N_5103);
or U6053 (N_6053,N_5693,N_5431);
or U6054 (N_6054,N_5313,N_5481);
nand U6055 (N_6055,N_5071,N_5789);
nand U6056 (N_6056,N_5033,N_5234);
or U6057 (N_6057,N_5877,N_5244);
and U6058 (N_6058,N_5310,N_5634);
and U6059 (N_6059,N_5685,N_5347);
or U6060 (N_6060,N_5328,N_5392);
and U6061 (N_6061,N_5189,N_5503);
and U6062 (N_6062,N_5333,N_5895);
or U6063 (N_6063,N_5858,N_5156);
or U6064 (N_6064,N_5390,N_5865);
and U6065 (N_6065,N_5602,N_5971);
or U6066 (N_6066,N_5383,N_5273);
or U6067 (N_6067,N_5535,N_5191);
nor U6068 (N_6068,N_5636,N_5592);
nor U6069 (N_6069,N_5699,N_5438);
or U6070 (N_6070,N_5808,N_5293);
or U6071 (N_6071,N_5461,N_5757);
xor U6072 (N_6072,N_5898,N_5662);
nor U6073 (N_6073,N_5522,N_5965);
nor U6074 (N_6074,N_5677,N_5212);
xor U6075 (N_6075,N_5550,N_5957);
or U6076 (N_6076,N_5633,N_5878);
xor U6077 (N_6077,N_5284,N_5985);
xor U6078 (N_6078,N_5304,N_5747);
nand U6079 (N_6079,N_5646,N_5175);
or U6080 (N_6080,N_5974,N_5824);
nor U6081 (N_6081,N_5381,N_5357);
and U6082 (N_6082,N_5143,N_5363);
and U6083 (N_6083,N_5630,N_5533);
xor U6084 (N_6084,N_5412,N_5635);
nor U6085 (N_6085,N_5053,N_5564);
and U6086 (N_6086,N_5648,N_5200);
nand U6087 (N_6087,N_5713,N_5737);
nand U6088 (N_6088,N_5521,N_5286);
nand U6089 (N_6089,N_5849,N_5764);
nor U6090 (N_6090,N_5266,N_5778);
or U6091 (N_6091,N_5332,N_5907);
and U6092 (N_6092,N_5744,N_5509);
nand U6093 (N_6093,N_5097,N_5239);
nand U6094 (N_6094,N_5445,N_5988);
and U6095 (N_6095,N_5351,N_5407);
or U6096 (N_6096,N_5477,N_5995);
or U6097 (N_6097,N_5855,N_5193);
xnor U6098 (N_6098,N_5358,N_5976);
nand U6099 (N_6099,N_5397,N_5834);
and U6100 (N_6100,N_5610,N_5991);
or U6101 (N_6101,N_5639,N_5784);
nor U6102 (N_6102,N_5369,N_5314);
and U6103 (N_6103,N_5119,N_5350);
nor U6104 (N_6104,N_5844,N_5723);
or U6105 (N_6105,N_5872,N_5349);
nand U6106 (N_6106,N_5593,N_5340);
or U6107 (N_6107,N_5946,N_5900);
xor U6108 (N_6108,N_5776,N_5794);
nor U6109 (N_6109,N_5890,N_5303);
nor U6110 (N_6110,N_5501,N_5285);
nor U6111 (N_6111,N_5155,N_5882);
xor U6112 (N_6112,N_5170,N_5616);
xor U6113 (N_6113,N_5839,N_5588);
or U6114 (N_6114,N_5426,N_5935);
or U6115 (N_6115,N_5981,N_5603);
or U6116 (N_6116,N_5423,N_5389);
nand U6117 (N_6117,N_5671,N_5224);
nand U6118 (N_6118,N_5538,N_5933);
xor U6119 (N_6119,N_5246,N_5765);
xor U6120 (N_6120,N_5548,N_5799);
nor U6121 (N_6121,N_5229,N_5888);
nor U6122 (N_6122,N_5572,N_5830);
nor U6123 (N_6123,N_5105,N_5066);
nor U6124 (N_6124,N_5181,N_5018);
or U6125 (N_6125,N_5360,N_5645);
xor U6126 (N_6126,N_5172,N_5518);
nand U6127 (N_6127,N_5682,N_5385);
nor U6128 (N_6128,N_5396,N_5036);
nand U6129 (N_6129,N_5243,N_5267);
or U6130 (N_6130,N_5524,N_5563);
xor U6131 (N_6131,N_5970,N_5044);
nor U6132 (N_6132,N_5746,N_5632);
or U6133 (N_6133,N_5270,N_5777);
and U6134 (N_6134,N_5562,N_5473);
nor U6135 (N_6135,N_5704,N_5037);
or U6136 (N_6136,N_5086,N_5906);
and U6137 (N_6137,N_5128,N_5190);
nand U6138 (N_6138,N_5422,N_5263);
and U6139 (N_6139,N_5821,N_5111);
nand U6140 (N_6140,N_5115,N_5498);
and U6141 (N_6141,N_5057,N_5732);
nor U6142 (N_6142,N_5098,N_5100);
and U6143 (N_6143,N_5462,N_5812);
nand U6144 (N_6144,N_5680,N_5968);
nand U6145 (N_6145,N_5655,N_5034);
and U6146 (N_6146,N_5718,N_5728);
nor U6147 (N_6147,N_5641,N_5251);
and U6148 (N_6148,N_5557,N_5698);
nand U6149 (N_6149,N_5998,N_5219);
or U6150 (N_6150,N_5841,N_5206);
xnor U6151 (N_6151,N_5241,N_5770);
or U6152 (N_6152,N_5060,N_5355);
or U6153 (N_6153,N_5640,N_5923);
xnor U6154 (N_6154,N_5049,N_5963);
nor U6155 (N_6155,N_5814,N_5594);
nor U6156 (N_6156,N_5424,N_5311);
or U6157 (N_6157,N_5712,N_5472);
nor U6158 (N_6158,N_5990,N_5398);
nand U6159 (N_6159,N_5217,N_5379);
or U6160 (N_6160,N_5800,N_5078);
xnor U6161 (N_6161,N_5252,N_5335);
xnor U6162 (N_6162,N_5090,N_5967);
and U6163 (N_6163,N_5318,N_5032);
nor U6164 (N_6164,N_5444,N_5202);
xnor U6165 (N_6165,N_5569,N_5300);
and U6166 (N_6166,N_5555,N_5135);
nor U6167 (N_6167,N_5195,N_5110);
or U6168 (N_6168,N_5317,N_5724);
and U6169 (N_6169,N_5609,N_5443);
xor U6170 (N_6170,N_5059,N_5870);
or U6171 (N_6171,N_5491,N_5945);
and U6172 (N_6172,N_5519,N_5931);
and U6173 (N_6173,N_5177,N_5949);
or U6174 (N_6174,N_5344,N_5955);
and U6175 (N_6175,N_5611,N_5586);
nand U6176 (N_6176,N_5067,N_5912);
or U6177 (N_6177,N_5506,N_5428);
and U6178 (N_6178,N_5301,N_5394);
xor U6179 (N_6179,N_5315,N_5720);
nor U6180 (N_6180,N_5857,N_5406);
nand U6181 (N_6181,N_5710,N_5901);
and U6182 (N_6182,N_5214,N_5675);
nor U6183 (N_6183,N_5487,N_5141);
nor U6184 (N_6184,N_5080,N_5769);
xor U6185 (N_6185,N_5657,N_5883);
and U6186 (N_6186,N_5331,N_5624);
or U6187 (N_6187,N_5176,N_5667);
or U6188 (N_6188,N_5023,N_5204);
nand U6189 (N_6189,N_5823,N_5388);
nand U6190 (N_6190,N_5738,N_5918);
and U6191 (N_6191,N_5021,N_5010);
xnor U6192 (N_6192,N_5911,N_5758);
nor U6193 (N_6193,N_5596,N_5816);
or U6194 (N_6194,N_5489,N_5617);
or U6195 (N_6195,N_5730,N_5168);
and U6196 (N_6196,N_5440,N_5245);
xor U6197 (N_6197,N_5979,N_5375);
xnor U6198 (N_6198,N_5525,N_5850);
and U6199 (N_6199,N_5926,N_5250);
or U6200 (N_6200,N_5948,N_5575);
nor U6201 (N_6201,N_5152,N_5837);
or U6202 (N_6202,N_5161,N_5560);
and U6203 (N_6203,N_5507,N_5618);
and U6204 (N_6204,N_5026,N_5124);
nand U6205 (N_6205,N_5077,N_5275);
nand U6206 (N_6206,N_5294,N_5248);
xor U6207 (N_6207,N_5165,N_5958);
or U6208 (N_6208,N_5120,N_5404);
nand U6209 (N_6209,N_5306,N_5674);
or U6210 (N_6210,N_5162,N_5714);
or U6211 (N_6211,N_5887,N_5631);
or U6212 (N_6212,N_5583,N_5269);
nor U6213 (N_6213,N_5045,N_5016);
and U6214 (N_6214,N_5289,N_5393);
nand U6215 (N_6215,N_5984,N_5915);
or U6216 (N_6216,N_5070,N_5441);
and U6217 (N_6217,N_5413,N_5400);
nand U6218 (N_6218,N_5451,N_5846);
and U6219 (N_6219,N_5411,N_5795);
and U6220 (N_6220,N_5584,N_5527);
or U6221 (N_6221,N_5539,N_5131);
nand U6222 (N_6222,N_5512,N_5924);
nor U6223 (N_6223,N_5199,N_5736);
nor U6224 (N_6224,N_5014,N_5327);
and U6225 (N_6225,N_5893,N_5471);
and U6226 (N_6226,N_5827,N_5806);
nand U6227 (N_6227,N_5669,N_5055);
and U6228 (N_6228,N_5042,N_5683);
nor U6229 (N_6229,N_5140,N_5492);
nor U6230 (N_6230,N_5697,N_5668);
nor U6231 (N_6231,N_5993,N_5566);
and U6232 (N_6232,N_5559,N_5866);
nor U6233 (N_6233,N_5410,N_5421);
and U6234 (N_6234,N_5227,N_5992);
nor U6235 (N_6235,N_5541,N_5715);
nand U6236 (N_6236,N_5366,N_5094);
and U6237 (N_6237,N_5845,N_5659);
or U6238 (N_6238,N_5178,N_5513);
xnor U6239 (N_6239,N_5807,N_5322);
and U6240 (N_6240,N_5851,N_5169);
nor U6241 (N_6241,N_5222,N_5308);
and U6242 (N_6242,N_5734,N_5601);
and U6243 (N_6243,N_5761,N_5242);
nand U6244 (N_6244,N_5030,N_5435);
and U6245 (N_6245,N_5232,N_5654);
or U6246 (N_6246,N_5719,N_5902);
nand U6247 (N_6247,N_5505,N_5585);
nand U6248 (N_6248,N_5947,N_5986);
or U6249 (N_6249,N_5977,N_5517);
nand U6250 (N_6250,N_5561,N_5781);
and U6251 (N_6251,N_5291,N_5035);
and U6252 (N_6252,N_5590,N_5904);
nor U6253 (N_6253,N_5419,N_5678);
nor U6254 (N_6254,N_5909,N_5171);
and U6255 (N_6255,N_5528,N_5651);
or U6256 (N_6256,N_5905,N_5571);
or U6257 (N_6257,N_5281,N_5801);
and U6258 (N_6258,N_5810,N_5129);
or U6259 (N_6259,N_5088,N_5208);
and U6260 (N_6260,N_5386,N_5287);
nor U6261 (N_6261,N_5999,N_5914);
nand U6262 (N_6262,N_5024,N_5576);
or U6263 (N_6263,N_5628,N_5319);
xor U6264 (N_6264,N_5068,N_5056);
nor U6265 (N_6265,N_5614,N_5228);
or U6266 (N_6266,N_5436,N_5701);
nand U6267 (N_6267,N_5006,N_5367);
nand U6268 (N_6268,N_5638,N_5540);
and U6269 (N_6269,N_5475,N_5399);
or U6270 (N_6270,N_5476,N_5828);
xor U6271 (N_6271,N_5929,N_5079);
nand U6272 (N_6272,N_5961,N_5039);
and U6273 (N_6273,N_5694,N_5916);
and U6274 (N_6274,N_5259,N_5690);
or U6275 (N_6275,N_5975,N_5871);
nand U6276 (N_6276,N_5387,N_5686);
or U6277 (N_6277,N_5953,N_5759);
nand U6278 (N_6278,N_5809,N_5791);
and U6279 (N_6279,N_5537,N_5565);
nor U6280 (N_6280,N_5515,N_5278);
nor U6281 (N_6281,N_5479,N_5288);
nor U6282 (N_6282,N_5994,N_5741);
nand U6283 (N_6283,N_5455,N_5198);
xor U6284 (N_6284,N_5420,N_5626);
or U6285 (N_6285,N_5125,N_5706);
nand U6286 (N_6286,N_5729,N_5962);
and U6287 (N_6287,N_5409,N_5458);
nand U6288 (N_6288,N_5230,N_5213);
or U6289 (N_6289,N_5203,N_5063);
nor U6290 (N_6290,N_5752,N_5921);
xnor U6291 (N_6291,N_5109,N_5254);
and U6292 (N_6292,N_5868,N_5427);
nor U6293 (N_6293,N_5612,N_5258);
nor U6294 (N_6294,N_5755,N_5302);
or U6295 (N_6295,N_5329,N_5969);
or U6296 (N_6296,N_5299,N_5932);
or U6297 (N_6297,N_5196,N_5825);
or U6298 (N_6298,N_5913,N_5666);
nor U6299 (N_6299,N_5001,N_5894);
nand U6300 (N_6300,N_5847,N_5889);
xnor U6301 (N_6301,N_5465,N_5076);
nand U6302 (N_6302,N_5605,N_5237);
and U6303 (N_6303,N_5545,N_5733);
xnor U6304 (N_6304,N_5074,N_5376);
and U6305 (N_6305,N_5186,N_5464);
or U6306 (N_6306,N_5779,N_5722);
and U6307 (N_6307,N_5739,N_5928);
nand U6308 (N_6308,N_5951,N_5069);
xnor U6309 (N_6309,N_5938,N_5051);
nor U6310 (N_6310,N_5046,N_5936);
nor U6311 (N_6311,N_5780,N_5925);
and U6312 (N_6312,N_5939,N_5943);
nor U6313 (N_6313,N_5022,N_5922);
and U6314 (N_6314,N_5762,N_5885);
nor U6315 (N_6315,N_5463,N_5166);
nand U6316 (N_6316,N_5276,N_5028);
xnor U6317 (N_6317,N_5280,N_5763);
nor U6318 (N_6318,N_5003,N_5663);
nand U6319 (N_6319,N_5980,N_5277);
nand U6320 (N_6320,N_5771,N_5688);
and U6321 (N_6321,N_5500,N_5373);
or U6322 (N_6322,N_5430,N_5395);
or U6323 (N_6323,N_5150,N_5073);
nand U6324 (N_6324,N_5772,N_5102);
nand U6325 (N_6325,N_5861,N_5615);
nor U6326 (N_6326,N_5247,N_5896);
nor U6327 (N_6327,N_5192,N_5691);
and U6328 (N_6328,N_5092,N_5339);
and U6329 (N_6329,N_5264,N_5265);
nor U6330 (N_6330,N_5742,N_5622);
and U6331 (N_6331,N_5785,N_5581);
and U6332 (N_6332,N_5826,N_5470);
nand U6333 (N_6333,N_5989,N_5972);
nor U6334 (N_6334,N_5323,N_5891);
nor U6335 (N_6335,N_5848,N_5341);
or U6336 (N_6336,N_5973,N_5283);
nand U6337 (N_6337,N_5937,N_5643);
and U6338 (N_6338,N_5884,N_5863);
nor U6339 (N_6339,N_5226,N_5818);
nand U6340 (N_6340,N_5838,N_5910);
or U6341 (N_6341,N_5117,N_5927);
nand U6342 (N_6342,N_5138,N_5708);
xnor U6343 (N_6343,N_5123,N_5833);
and U6344 (N_6344,N_5803,N_5004);
and U6345 (N_6345,N_5960,N_5978);
xnor U6346 (N_6346,N_5627,N_5620);
nand U6347 (N_6347,N_5173,N_5920);
nand U6348 (N_6348,N_5589,N_5859);
or U6349 (N_6349,N_5672,N_5775);
and U6350 (N_6350,N_5474,N_5298);
nor U6351 (N_6351,N_5570,N_5043);
nand U6352 (N_6352,N_5013,N_5748);
nor U6353 (N_6353,N_5787,N_5743);
and U6354 (N_6354,N_5337,N_5544);
nor U6355 (N_6355,N_5613,N_5793);
or U6356 (N_6356,N_5797,N_5136);
or U6357 (N_6357,N_5485,N_5145);
or U6358 (N_6358,N_5835,N_5361);
or U6359 (N_6359,N_5652,N_5151);
nand U6360 (N_6360,N_5144,N_5184);
and U6361 (N_6361,N_5899,N_5020);
and U6362 (N_6362,N_5268,N_5345);
and U6363 (N_6363,N_5494,N_5447);
nor U6364 (N_6364,N_5130,N_5188);
nor U6365 (N_6365,N_5598,N_5083);
xor U6366 (N_6366,N_5163,N_5142);
or U6367 (N_6367,N_5940,N_5295);
or U6368 (N_6368,N_5488,N_5879);
or U6369 (N_6369,N_5180,N_5597);
xnor U6370 (N_6370,N_5343,N_5676);
or U6371 (N_6371,N_5238,N_5749);
or U6372 (N_6372,N_5642,N_5842);
nor U6373 (N_6373,N_5187,N_5623);
nor U6374 (N_6374,N_5364,N_5954);
nor U6375 (N_6375,N_5334,N_5153);
or U6376 (N_6376,N_5829,N_5015);
and U6377 (N_6377,N_5442,N_5950);
and U6378 (N_6378,N_5695,N_5336);
and U6379 (N_6379,N_5460,N_5439);
nor U6380 (N_6380,N_5365,N_5727);
and U6381 (N_6381,N_5530,N_5608);
and U6382 (N_6382,N_5402,N_5121);
xor U6383 (N_6383,N_5567,N_5493);
and U6384 (N_6384,N_5132,N_5256);
or U6385 (N_6385,N_5054,N_5917);
or U6386 (N_6386,N_5553,N_5941);
or U6387 (N_6387,N_5956,N_5881);
nand U6388 (N_6388,N_5127,N_5257);
or U6389 (N_6389,N_5843,N_5348);
nor U6390 (N_6390,N_5903,N_5201);
nand U6391 (N_6391,N_5223,N_5220);
nand U6392 (N_6392,N_5766,N_5118);
or U6393 (N_6393,N_5573,N_5740);
xor U6394 (N_6394,N_5457,N_5296);
nand U6395 (N_6395,N_5216,N_5696);
and U6396 (N_6396,N_5495,N_5017);
and U6397 (N_6397,N_5297,N_5482);
and U6398 (N_6398,N_5401,N_5330);
nand U6399 (N_6399,N_5983,N_5711);
and U6400 (N_6400,N_5637,N_5048);
nand U6401 (N_6401,N_5629,N_5582);
nand U6402 (N_6402,N_5005,N_5108);
nor U6403 (N_6403,N_5886,N_5425);
xnor U6404 (N_6404,N_5496,N_5075);
or U6405 (N_6405,N_5215,N_5673);
xnor U6406 (N_6406,N_5549,N_5371);
and U6407 (N_6407,N_5047,N_5867);
or U6408 (N_6408,N_5930,N_5864);
or U6409 (N_6409,N_5391,N_5508);
or U6410 (N_6410,N_5982,N_5377);
nor U6411 (N_6411,N_5352,N_5255);
xor U6412 (N_6412,N_5236,N_5221);
nor U6413 (N_6413,N_5831,N_5469);
xor U6414 (N_6414,N_5547,N_5065);
nand U6415 (N_6415,N_5207,N_5966);
nor U6416 (N_6416,N_5959,N_5782);
nand U6417 (N_6417,N_5429,N_5353);
xnor U6418 (N_6418,N_5085,N_5194);
nand U6419 (N_6419,N_5745,N_5773);
or U6420 (N_6420,N_5502,N_5653);
nor U6421 (N_6421,N_5490,N_5456);
nor U6422 (N_6422,N_5040,N_5211);
nor U6423 (N_6423,N_5122,N_5378);
or U6424 (N_6424,N_5811,N_5532);
xor U6425 (N_6425,N_5011,N_5146);
or U6426 (N_6426,N_5558,N_5661);
and U6427 (N_6427,N_5689,N_5174);
and U6428 (N_6428,N_5338,N_5551);
and U6429 (N_6429,N_5554,N_5874);
and U6430 (N_6430,N_5520,N_5370);
nand U6431 (N_6431,N_5261,N_5368);
and U6432 (N_6432,N_5019,N_5179);
xor U6433 (N_6433,N_5840,N_5249);
or U6434 (N_6434,N_5099,N_5082);
nand U6435 (N_6435,N_5096,N_5591);
or U6436 (N_6436,N_5309,N_5542);
or U6437 (N_6437,N_5164,N_5942);
nand U6438 (N_6438,N_5240,N_5104);
and U6439 (N_6439,N_5499,N_5072);
or U6440 (N_6440,N_5454,N_5089);
and U6441 (N_6441,N_5197,N_5987);
and U6442 (N_6442,N_5149,N_5324);
xnor U6443 (N_6443,N_5305,N_5113);
nand U6444 (N_6444,N_5934,N_5997);
or U6445 (N_6445,N_5852,N_5792);
nand U6446 (N_6446,N_5819,N_5604);
nor U6447 (N_6447,N_5875,N_5644);
nand U6448 (N_6448,N_5813,N_5274);
or U6449 (N_6449,N_5531,N_5093);
and U6450 (N_6450,N_5483,N_5815);
nand U6451 (N_6451,N_5709,N_5873);
and U6452 (N_6452,N_5466,N_5625);
or U6453 (N_6453,N_5061,N_5262);
xnor U6454 (N_6454,N_5316,N_5869);
and U6455 (N_6455,N_5860,N_5580);
or U6456 (N_6456,N_5167,N_5536);
nand U6457 (N_6457,N_5225,N_5587);
nor U6458 (N_6458,N_5346,N_5692);
nand U6459 (N_6459,N_5453,N_5880);
nor U6460 (N_6460,N_5665,N_5467);
or U6461 (N_6461,N_5205,N_5272);
or U6462 (N_6462,N_5137,N_5107);
nand U6463 (N_6463,N_5403,N_5359);
xor U6464 (N_6464,N_5081,N_5372);
or U6465 (N_6465,N_5731,N_5798);
nand U6466 (N_6466,N_5157,N_5892);
or U6467 (N_6467,N_5684,N_5101);
and U6468 (N_6468,N_5116,N_5964);
xnor U6469 (N_6469,N_5534,N_5446);
xor U6470 (N_6470,N_5408,N_5760);
nand U6471 (N_6471,N_5185,N_5031);
and U6472 (N_6472,N_5523,N_5497);
and U6473 (N_6473,N_5647,N_5029);
xor U6474 (N_6474,N_5836,N_5414);
and U6475 (N_6475,N_5707,N_5416);
and U6476 (N_6476,N_5290,N_5002);
and U6477 (N_6477,N_5511,N_5774);
or U6478 (N_6478,N_5459,N_5432);
xnor U6479 (N_6479,N_5091,N_5703);
or U6480 (N_6480,N_5574,N_5788);
and U6481 (N_6481,N_5578,N_5405);
xnor U6482 (N_6482,N_5210,N_5556);
xnor U6483 (N_6483,N_5577,N_5805);
or U6484 (N_6484,N_5449,N_5750);
nand U6485 (N_6485,N_5681,N_5126);
and U6486 (N_6486,N_5660,N_5721);
and U6487 (N_6487,N_5529,N_5148);
or U6488 (N_6488,N_5670,N_5768);
nand U6489 (N_6489,N_5374,N_5382);
and U6490 (N_6490,N_5543,N_5062);
nand U6491 (N_6491,N_5510,N_5007);
nor U6492 (N_6492,N_5312,N_5621);
nor U6493 (N_6493,N_5717,N_5158);
and U6494 (N_6494,N_5417,N_5702);
and U6495 (N_6495,N_5218,N_5679);
xor U6496 (N_6496,N_5725,N_5433);
and U6497 (N_6497,N_5897,N_5292);
nor U6498 (N_6498,N_5664,N_5796);
nor U6499 (N_6499,N_5362,N_5820);
or U6500 (N_6500,N_5084,N_5819);
nand U6501 (N_6501,N_5128,N_5236);
nand U6502 (N_6502,N_5569,N_5031);
nand U6503 (N_6503,N_5926,N_5079);
or U6504 (N_6504,N_5378,N_5553);
nand U6505 (N_6505,N_5579,N_5049);
and U6506 (N_6506,N_5347,N_5222);
or U6507 (N_6507,N_5073,N_5502);
nor U6508 (N_6508,N_5374,N_5856);
nand U6509 (N_6509,N_5967,N_5497);
or U6510 (N_6510,N_5554,N_5343);
nand U6511 (N_6511,N_5552,N_5481);
nor U6512 (N_6512,N_5727,N_5379);
nand U6513 (N_6513,N_5314,N_5206);
nor U6514 (N_6514,N_5291,N_5487);
and U6515 (N_6515,N_5943,N_5261);
xor U6516 (N_6516,N_5088,N_5036);
or U6517 (N_6517,N_5974,N_5073);
or U6518 (N_6518,N_5881,N_5488);
nand U6519 (N_6519,N_5401,N_5312);
and U6520 (N_6520,N_5011,N_5703);
or U6521 (N_6521,N_5600,N_5426);
or U6522 (N_6522,N_5012,N_5863);
or U6523 (N_6523,N_5683,N_5881);
and U6524 (N_6524,N_5565,N_5245);
nor U6525 (N_6525,N_5203,N_5570);
xor U6526 (N_6526,N_5081,N_5487);
xnor U6527 (N_6527,N_5795,N_5839);
nand U6528 (N_6528,N_5777,N_5246);
xor U6529 (N_6529,N_5368,N_5958);
nand U6530 (N_6530,N_5731,N_5218);
xor U6531 (N_6531,N_5365,N_5558);
nor U6532 (N_6532,N_5838,N_5269);
or U6533 (N_6533,N_5632,N_5785);
or U6534 (N_6534,N_5547,N_5028);
and U6535 (N_6535,N_5289,N_5555);
nand U6536 (N_6536,N_5784,N_5093);
and U6537 (N_6537,N_5573,N_5752);
nand U6538 (N_6538,N_5407,N_5743);
nor U6539 (N_6539,N_5510,N_5415);
xor U6540 (N_6540,N_5552,N_5006);
nor U6541 (N_6541,N_5060,N_5618);
or U6542 (N_6542,N_5547,N_5802);
and U6543 (N_6543,N_5061,N_5354);
or U6544 (N_6544,N_5170,N_5925);
or U6545 (N_6545,N_5972,N_5642);
nand U6546 (N_6546,N_5874,N_5285);
and U6547 (N_6547,N_5700,N_5395);
nand U6548 (N_6548,N_5764,N_5422);
nor U6549 (N_6549,N_5366,N_5274);
nor U6550 (N_6550,N_5740,N_5998);
and U6551 (N_6551,N_5804,N_5923);
nand U6552 (N_6552,N_5896,N_5593);
or U6553 (N_6553,N_5903,N_5092);
and U6554 (N_6554,N_5545,N_5649);
nand U6555 (N_6555,N_5937,N_5783);
or U6556 (N_6556,N_5572,N_5431);
nand U6557 (N_6557,N_5685,N_5684);
or U6558 (N_6558,N_5230,N_5601);
nor U6559 (N_6559,N_5707,N_5596);
and U6560 (N_6560,N_5901,N_5044);
nand U6561 (N_6561,N_5457,N_5611);
nand U6562 (N_6562,N_5733,N_5796);
and U6563 (N_6563,N_5637,N_5572);
or U6564 (N_6564,N_5741,N_5282);
and U6565 (N_6565,N_5615,N_5937);
or U6566 (N_6566,N_5571,N_5836);
and U6567 (N_6567,N_5829,N_5766);
and U6568 (N_6568,N_5490,N_5085);
nand U6569 (N_6569,N_5333,N_5357);
nor U6570 (N_6570,N_5110,N_5113);
xnor U6571 (N_6571,N_5734,N_5633);
xnor U6572 (N_6572,N_5748,N_5049);
xor U6573 (N_6573,N_5663,N_5647);
or U6574 (N_6574,N_5536,N_5557);
or U6575 (N_6575,N_5814,N_5295);
nor U6576 (N_6576,N_5043,N_5921);
nor U6577 (N_6577,N_5534,N_5679);
xnor U6578 (N_6578,N_5700,N_5575);
nand U6579 (N_6579,N_5789,N_5216);
and U6580 (N_6580,N_5865,N_5239);
xnor U6581 (N_6581,N_5694,N_5489);
or U6582 (N_6582,N_5558,N_5829);
xor U6583 (N_6583,N_5310,N_5976);
nand U6584 (N_6584,N_5572,N_5402);
and U6585 (N_6585,N_5482,N_5073);
and U6586 (N_6586,N_5231,N_5059);
nand U6587 (N_6587,N_5904,N_5554);
nand U6588 (N_6588,N_5801,N_5484);
nand U6589 (N_6589,N_5220,N_5142);
xor U6590 (N_6590,N_5222,N_5905);
xnor U6591 (N_6591,N_5593,N_5814);
and U6592 (N_6592,N_5865,N_5574);
or U6593 (N_6593,N_5566,N_5811);
or U6594 (N_6594,N_5747,N_5298);
nand U6595 (N_6595,N_5381,N_5639);
nand U6596 (N_6596,N_5907,N_5799);
or U6597 (N_6597,N_5637,N_5925);
nand U6598 (N_6598,N_5143,N_5896);
nand U6599 (N_6599,N_5759,N_5724);
or U6600 (N_6600,N_5476,N_5561);
and U6601 (N_6601,N_5202,N_5185);
or U6602 (N_6602,N_5364,N_5182);
or U6603 (N_6603,N_5296,N_5721);
and U6604 (N_6604,N_5429,N_5884);
and U6605 (N_6605,N_5764,N_5211);
xor U6606 (N_6606,N_5397,N_5881);
nor U6607 (N_6607,N_5696,N_5683);
nand U6608 (N_6608,N_5917,N_5845);
or U6609 (N_6609,N_5194,N_5186);
and U6610 (N_6610,N_5717,N_5709);
or U6611 (N_6611,N_5887,N_5241);
xor U6612 (N_6612,N_5949,N_5849);
nor U6613 (N_6613,N_5203,N_5273);
nand U6614 (N_6614,N_5466,N_5612);
or U6615 (N_6615,N_5429,N_5890);
nor U6616 (N_6616,N_5505,N_5996);
xnor U6617 (N_6617,N_5447,N_5138);
nand U6618 (N_6618,N_5463,N_5066);
nand U6619 (N_6619,N_5020,N_5206);
nand U6620 (N_6620,N_5331,N_5357);
and U6621 (N_6621,N_5088,N_5325);
xor U6622 (N_6622,N_5617,N_5149);
nor U6623 (N_6623,N_5724,N_5847);
or U6624 (N_6624,N_5617,N_5793);
and U6625 (N_6625,N_5450,N_5586);
or U6626 (N_6626,N_5689,N_5564);
xor U6627 (N_6627,N_5035,N_5552);
or U6628 (N_6628,N_5893,N_5245);
nor U6629 (N_6629,N_5886,N_5771);
and U6630 (N_6630,N_5856,N_5782);
nor U6631 (N_6631,N_5179,N_5938);
nand U6632 (N_6632,N_5578,N_5391);
and U6633 (N_6633,N_5459,N_5670);
or U6634 (N_6634,N_5001,N_5767);
nand U6635 (N_6635,N_5633,N_5970);
nor U6636 (N_6636,N_5114,N_5241);
nor U6637 (N_6637,N_5635,N_5196);
nand U6638 (N_6638,N_5158,N_5969);
or U6639 (N_6639,N_5456,N_5243);
nor U6640 (N_6640,N_5954,N_5806);
and U6641 (N_6641,N_5829,N_5017);
nor U6642 (N_6642,N_5594,N_5445);
and U6643 (N_6643,N_5906,N_5176);
nor U6644 (N_6644,N_5388,N_5528);
nor U6645 (N_6645,N_5984,N_5951);
nor U6646 (N_6646,N_5670,N_5209);
or U6647 (N_6647,N_5913,N_5097);
or U6648 (N_6648,N_5906,N_5343);
nand U6649 (N_6649,N_5608,N_5406);
or U6650 (N_6650,N_5020,N_5494);
and U6651 (N_6651,N_5937,N_5676);
nand U6652 (N_6652,N_5891,N_5303);
xor U6653 (N_6653,N_5319,N_5750);
and U6654 (N_6654,N_5542,N_5777);
or U6655 (N_6655,N_5440,N_5773);
nor U6656 (N_6656,N_5499,N_5047);
nor U6657 (N_6657,N_5616,N_5714);
xor U6658 (N_6658,N_5057,N_5079);
or U6659 (N_6659,N_5388,N_5161);
and U6660 (N_6660,N_5907,N_5702);
nor U6661 (N_6661,N_5749,N_5377);
and U6662 (N_6662,N_5105,N_5294);
nor U6663 (N_6663,N_5942,N_5448);
xnor U6664 (N_6664,N_5977,N_5255);
nor U6665 (N_6665,N_5126,N_5142);
xor U6666 (N_6666,N_5039,N_5006);
and U6667 (N_6667,N_5297,N_5847);
nand U6668 (N_6668,N_5675,N_5375);
nand U6669 (N_6669,N_5477,N_5545);
nand U6670 (N_6670,N_5004,N_5743);
or U6671 (N_6671,N_5467,N_5071);
nor U6672 (N_6672,N_5762,N_5422);
and U6673 (N_6673,N_5529,N_5441);
nor U6674 (N_6674,N_5486,N_5321);
xnor U6675 (N_6675,N_5163,N_5729);
or U6676 (N_6676,N_5508,N_5039);
nor U6677 (N_6677,N_5403,N_5842);
or U6678 (N_6678,N_5792,N_5253);
and U6679 (N_6679,N_5895,N_5399);
and U6680 (N_6680,N_5639,N_5314);
nor U6681 (N_6681,N_5353,N_5594);
nor U6682 (N_6682,N_5289,N_5063);
or U6683 (N_6683,N_5179,N_5750);
nand U6684 (N_6684,N_5550,N_5236);
and U6685 (N_6685,N_5750,N_5951);
or U6686 (N_6686,N_5313,N_5999);
nor U6687 (N_6687,N_5308,N_5050);
or U6688 (N_6688,N_5841,N_5843);
nor U6689 (N_6689,N_5335,N_5020);
or U6690 (N_6690,N_5159,N_5378);
or U6691 (N_6691,N_5092,N_5332);
xor U6692 (N_6692,N_5520,N_5323);
and U6693 (N_6693,N_5458,N_5015);
nand U6694 (N_6694,N_5605,N_5356);
nor U6695 (N_6695,N_5885,N_5367);
or U6696 (N_6696,N_5593,N_5847);
nor U6697 (N_6697,N_5157,N_5541);
nand U6698 (N_6698,N_5662,N_5397);
nor U6699 (N_6699,N_5853,N_5493);
and U6700 (N_6700,N_5534,N_5637);
and U6701 (N_6701,N_5501,N_5210);
nor U6702 (N_6702,N_5598,N_5978);
nand U6703 (N_6703,N_5427,N_5844);
and U6704 (N_6704,N_5100,N_5702);
or U6705 (N_6705,N_5932,N_5432);
nor U6706 (N_6706,N_5007,N_5088);
nor U6707 (N_6707,N_5225,N_5881);
nor U6708 (N_6708,N_5775,N_5044);
nor U6709 (N_6709,N_5901,N_5519);
or U6710 (N_6710,N_5287,N_5078);
nand U6711 (N_6711,N_5154,N_5766);
xor U6712 (N_6712,N_5771,N_5225);
and U6713 (N_6713,N_5758,N_5250);
nor U6714 (N_6714,N_5451,N_5526);
and U6715 (N_6715,N_5222,N_5541);
nand U6716 (N_6716,N_5297,N_5628);
nand U6717 (N_6717,N_5754,N_5182);
xor U6718 (N_6718,N_5533,N_5551);
xnor U6719 (N_6719,N_5261,N_5706);
nand U6720 (N_6720,N_5024,N_5416);
or U6721 (N_6721,N_5070,N_5615);
nand U6722 (N_6722,N_5310,N_5733);
nor U6723 (N_6723,N_5051,N_5116);
and U6724 (N_6724,N_5868,N_5826);
nor U6725 (N_6725,N_5397,N_5167);
and U6726 (N_6726,N_5811,N_5754);
and U6727 (N_6727,N_5757,N_5627);
or U6728 (N_6728,N_5102,N_5677);
or U6729 (N_6729,N_5773,N_5652);
and U6730 (N_6730,N_5686,N_5264);
nor U6731 (N_6731,N_5792,N_5780);
and U6732 (N_6732,N_5416,N_5367);
nor U6733 (N_6733,N_5699,N_5175);
nand U6734 (N_6734,N_5782,N_5611);
xor U6735 (N_6735,N_5482,N_5235);
xnor U6736 (N_6736,N_5077,N_5645);
nor U6737 (N_6737,N_5502,N_5974);
and U6738 (N_6738,N_5187,N_5627);
nor U6739 (N_6739,N_5365,N_5662);
xnor U6740 (N_6740,N_5029,N_5967);
and U6741 (N_6741,N_5068,N_5175);
or U6742 (N_6742,N_5128,N_5517);
nand U6743 (N_6743,N_5606,N_5011);
nor U6744 (N_6744,N_5753,N_5388);
xnor U6745 (N_6745,N_5798,N_5678);
and U6746 (N_6746,N_5938,N_5451);
or U6747 (N_6747,N_5601,N_5432);
and U6748 (N_6748,N_5065,N_5500);
nand U6749 (N_6749,N_5489,N_5054);
xnor U6750 (N_6750,N_5732,N_5044);
and U6751 (N_6751,N_5198,N_5849);
nand U6752 (N_6752,N_5974,N_5343);
or U6753 (N_6753,N_5004,N_5079);
and U6754 (N_6754,N_5118,N_5139);
and U6755 (N_6755,N_5366,N_5192);
and U6756 (N_6756,N_5588,N_5339);
xnor U6757 (N_6757,N_5066,N_5576);
or U6758 (N_6758,N_5816,N_5521);
nand U6759 (N_6759,N_5568,N_5861);
nand U6760 (N_6760,N_5952,N_5326);
xor U6761 (N_6761,N_5569,N_5367);
or U6762 (N_6762,N_5397,N_5616);
nand U6763 (N_6763,N_5233,N_5392);
or U6764 (N_6764,N_5359,N_5782);
nor U6765 (N_6765,N_5373,N_5944);
and U6766 (N_6766,N_5014,N_5511);
and U6767 (N_6767,N_5585,N_5826);
nor U6768 (N_6768,N_5407,N_5679);
or U6769 (N_6769,N_5901,N_5828);
and U6770 (N_6770,N_5077,N_5367);
nor U6771 (N_6771,N_5037,N_5871);
nor U6772 (N_6772,N_5422,N_5691);
nor U6773 (N_6773,N_5065,N_5989);
and U6774 (N_6774,N_5536,N_5681);
or U6775 (N_6775,N_5115,N_5076);
and U6776 (N_6776,N_5102,N_5669);
nand U6777 (N_6777,N_5702,N_5705);
xnor U6778 (N_6778,N_5093,N_5567);
or U6779 (N_6779,N_5273,N_5760);
or U6780 (N_6780,N_5369,N_5356);
and U6781 (N_6781,N_5601,N_5275);
nand U6782 (N_6782,N_5923,N_5210);
and U6783 (N_6783,N_5334,N_5425);
nand U6784 (N_6784,N_5989,N_5165);
and U6785 (N_6785,N_5915,N_5667);
nor U6786 (N_6786,N_5332,N_5392);
nor U6787 (N_6787,N_5886,N_5929);
nor U6788 (N_6788,N_5744,N_5108);
and U6789 (N_6789,N_5728,N_5752);
nand U6790 (N_6790,N_5925,N_5536);
or U6791 (N_6791,N_5656,N_5640);
or U6792 (N_6792,N_5309,N_5147);
nor U6793 (N_6793,N_5382,N_5112);
or U6794 (N_6794,N_5807,N_5148);
and U6795 (N_6795,N_5054,N_5837);
nand U6796 (N_6796,N_5920,N_5620);
nand U6797 (N_6797,N_5204,N_5134);
and U6798 (N_6798,N_5213,N_5699);
and U6799 (N_6799,N_5475,N_5927);
nand U6800 (N_6800,N_5816,N_5279);
or U6801 (N_6801,N_5929,N_5489);
or U6802 (N_6802,N_5011,N_5063);
nor U6803 (N_6803,N_5566,N_5211);
and U6804 (N_6804,N_5897,N_5189);
xor U6805 (N_6805,N_5037,N_5448);
nor U6806 (N_6806,N_5679,N_5828);
nand U6807 (N_6807,N_5301,N_5926);
nand U6808 (N_6808,N_5203,N_5865);
or U6809 (N_6809,N_5891,N_5981);
and U6810 (N_6810,N_5711,N_5930);
xnor U6811 (N_6811,N_5896,N_5964);
xor U6812 (N_6812,N_5477,N_5786);
or U6813 (N_6813,N_5301,N_5310);
or U6814 (N_6814,N_5725,N_5506);
and U6815 (N_6815,N_5155,N_5500);
xor U6816 (N_6816,N_5633,N_5522);
and U6817 (N_6817,N_5831,N_5921);
and U6818 (N_6818,N_5666,N_5268);
nand U6819 (N_6819,N_5016,N_5952);
nor U6820 (N_6820,N_5226,N_5481);
or U6821 (N_6821,N_5940,N_5174);
nor U6822 (N_6822,N_5546,N_5949);
nand U6823 (N_6823,N_5648,N_5350);
nor U6824 (N_6824,N_5383,N_5104);
or U6825 (N_6825,N_5141,N_5409);
xnor U6826 (N_6826,N_5577,N_5201);
nand U6827 (N_6827,N_5623,N_5436);
or U6828 (N_6828,N_5106,N_5703);
nand U6829 (N_6829,N_5593,N_5036);
nor U6830 (N_6830,N_5498,N_5081);
and U6831 (N_6831,N_5660,N_5430);
or U6832 (N_6832,N_5344,N_5623);
and U6833 (N_6833,N_5590,N_5221);
or U6834 (N_6834,N_5901,N_5047);
and U6835 (N_6835,N_5468,N_5908);
nor U6836 (N_6836,N_5901,N_5986);
and U6837 (N_6837,N_5069,N_5809);
or U6838 (N_6838,N_5128,N_5148);
nor U6839 (N_6839,N_5220,N_5383);
or U6840 (N_6840,N_5314,N_5144);
or U6841 (N_6841,N_5614,N_5607);
nor U6842 (N_6842,N_5605,N_5010);
and U6843 (N_6843,N_5264,N_5711);
nand U6844 (N_6844,N_5222,N_5511);
nand U6845 (N_6845,N_5104,N_5065);
or U6846 (N_6846,N_5096,N_5482);
nor U6847 (N_6847,N_5201,N_5685);
nand U6848 (N_6848,N_5777,N_5656);
or U6849 (N_6849,N_5189,N_5454);
nor U6850 (N_6850,N_5131,N_5468);
nor U6851 (N_6851,N_5548,N_5275);
nor U6852 (N_6852,N_5101,N_5599);
nand U6853 (N_6853,N_5070,N_5542);
xor U6854 (N_6854,N_5894,N_5641);
and U6855 (N_6855,N_5409,N_5646);
nor U6856 (N_6856,N_5738,N_5234);
or U6857 (N_6857,N_5597,N_5638);
and U6858 (N_6858,N_5153,N_5879);
nand U6859 (N_6859,N_5428,N_5908);
or U6860 (N_6860,N_5959,N_5896);
nor U6861 (N_6861,N_5938,N_5034);
or U6862 (N_6862,N_5755,N_5270);
nand U6863 (N_6863,N_5259,N_5064);
xnor U6864 (N_6864,N_5605,N_5923);
nor U6865 (N_6865,N_5043,N_5804);
or U6866 (N_6866,N_5715,N_5059);
nor U6867 (N_6867,N_5216,N_5947);
xnor U6868 (N_6868,N_5302,N_5542);
or U6869 (N_6869,N_5708,N_5488);
and U6870 (N_6870,N_5729,N_5570);
and U6871 (N_6871,N_5546,N_5262);
or U6872 (N_6872,N_5623,N_5749);
or U6873 (N_6873,N_5976,N_5616);
nand U6874 (N_6874,N_5346,N_5409);
and U6875 (N_6875,N_5442,N_5802);
and U6876 (N_6876,N_5533,N_5045);
nand U6877 (N_6877,N_5589,N_5383);
and U6878 (N_6878,N_5172,N_5714);
nor U6879 (N_6879,N_5206,N_5776);
nor U6880 (N_6880,N_5866,N_5191);
nor U6881 (N_6881,N_5313,N_5415);
nor U6882 (N_6882,N_5367,N_5446);
nor U6883 (N_6883,N_5808,N_5058);
or U6884 (N_6884,N_5409,N_5746);
and U6885 (N_6885,N_5929,N_5374);
nand U6886 (N_6886,N_5088,N_5274);
or U6887 (N_6887,N_5130,N_5634);
nand U6888 (N_6888,N_5565,N_5598);
nor U6889 (N_6889,N_5924,N_5727);
nor U6890 (N_6890,N_5498,N_5566);
nand U6891 (N_6891,N_5049,N_5282);
and U6892 (N_6892,N_5243,N_5857);
nand U6893 (N_6893,N_5293,N_5136);
and U6894 (N_6894,N_5725,N_5622);
and U6895 (N_6895,N_5300,N_5591);
nand U6896 (N_6896,N_5903,N_5051);
or U6897 (N_6897,N_5123,N_5395);
nand U6898 (N_6898,N_5328,N_5949);
nor U6899 (N_6899,N_5269,N_5197);
and U6900 (N_6900,N_5083,N_5906);
nor U6901 (N_6901,N_5344,N_5293);
nor U6902 (N_6902,N_5688,N_5839);
nor U6903 (N_6903,N_5795,N_5969);
or U6904 (N_6904,N_5699,N_5839);
or U6905 (N_6905,N_5878,N_5117);
xnor U6906 (N_6906,N_5837,N_5014);
and U6907 (N_6907,N_5050,N_5554);
nand U6908 (N_6908,N_5831,N_5216);
nor U6909 (N_6909,N_5022,N_5481);
nand U6910 (N_6910,N_5067,N_5788);
and U6911 (N_6911,N_5232,N_5399);
and U6912 (N_6912,N_5546,N_5221);
or U6913 (N_6913,N_5462,N_5426);
xor U6914 (N_6914,N_5661,N_5452);
nand U6915 (N_6915,N_5034,N_5328);
and U6916 (N_6916,N_5049,N_5704);
nand U6917 (N_6917,N_5074,N_5121);
xor U6918 (N_6918,N_5586,N_5917);
or U6919 (N_6919,N_5824,N_5761);
nor U6920 (N_6920,N_5036,N_5161);
or U6921 (N_6921,N_5824,N_5318);
nor U6922 (N_6922,N_5391,N_5417);
nand U6923 (N_6923,N_5385,N_5878);
nor U6924 (N_6924,N_5027,N_5180);
or U6925 (N_6925,N_5893,N_5404);
nor U6926 (N_6926,N_5582,N_5673);
and U6927 (N_6927,N_5444,N_5722);
nor U6928 (N_6928,N_5638,N_5164);
nand U6929 (N_6929,N_5143,N_5023);
or U6930 (N_6930,N_5433,N_5879);
nand U6931 (N_6931,N_5324,N_5335);
and U6932 (N_6932,N_5762,N_5377);
and U6933 (N_6933,N_5211,N_5170);
and U6934 (N_6934,N_5286,N_5712);
or U6935 (N_6935,N_5436,N_5999);
nand U6936 (N_6936,N_5777,N_5074);
nand U6937 (N_6937,N_5018,N_5169);
xor U6938 (N_6938,N_5017,N_5602);
nor U6939 (N_6939,N_5384,N_5327);
xor U6940 (N_6940,N_5753,N_5533);
or U6941 (N_6941,N_5448,N_5262);
xnor U6942 (N_6942,N_5786,N_5797);
xnor U6943 (N_6943,N_5147,N_5396);
nand U6944 (N_6944,N_5670,N_5040);
nor U6945 (N_6945,N_5060,N_5904);
xor U6946 (N_6946,N_5076,N_5155);
xor U6947 (N_6947,N_5291,N_5784);
nor U6948 (N_6948,N_5567,N_5742);
and U6949 (N_6949,N_5613,N_5233);
nand U6950 (N_6950,N_5295,N_5929);
or U6951 (N_6951,N_5821,N_5244);
nor U6952 (N_6952,N_5718,N_5200);
nor U6953 (N_6953,N_5636,N_5206);
nor U6954 (N_6954,N_5995,N_5481);
nor U6955 (N_6955,N_5797,N_5737);
and U6956 (N_6956,N_5477,N_5788);
nor U6957 (N_6957,N_5849,N_5148);
and U6958 (N_6958,N_5641,N_5394);
and U6959 (N_6959,N_5293,N_5735);
nand U6960 (N_6960,N_5689,N_5646);
nand U6961 (N_6961,N_5905,N_5243);
or U6962 (N_6962,N_5398,N_5319);
and U6963 (N_6963,N_5564,N_5864);
nand U6964 (N_6964,N_5200,N_5696);
or U6965 (N_6965,N_5304,N_5894);
and U6966 (N_6966,N_5774,N_5349);
xnor U6967 (N_6967,N_5529,N_5952);
nor U6968 (N_6968,N_5071,N_5949);
and U6969 (N_6969,N_5727,N_5376);
nor U6970 (N_6970,N_5286,N_5105);
nor U6971 (N_6971,N_5051,N_5090);
xor U6972 (N_6972,N_5355,N_5167);
nand U6973 (N_6973,N_5594,N_5583);
or U6974 (N_6974,N_5963,N_5289);
nor U6975 (N_6975,N_5792,N_5378);
nor U6976 (N_6976,N_5961,N_5549);
nor U6977 (N_6977,N_5066,N_5598);
nand U6978 (N_6978,N_5295,N_5985);
nor U6979 (N_6979,N_5867,N_5559);
and U6980 (N_6980,N_5833,N_5121);
and U6981 (N_6981,N_5841,N_5142);
or U6982 (N_6982,N_5630,N_5193);
and U6983 (N_6983,N_5156,N_5863);
and U6984 (N_6984,N_5079,N_5569);
nand U6985 (N_6985,N_5414,N_5971);
nor U6986 (N_6986,N_5270,N_5404);
nor U6987 (N_6987,N_5863,N_5649);
nor U6988 (N_6988,N_5358,N_5002);
and U6989 (N_6989,N_5460,N_5609);
or U6990 (N_6990,N_5973,N_5159);
or U6991 (N_6991,N_5191,N_5122);
and U6992 (N_6992,N_5182,N_5464);
nor U6993 (N_6993,N_5714,N_5274);
and U6994 (N_6994,N_5363,N_5415);
and U6995 (N_6995,N_5292,N_5610);
nor U6996 (N_6996,N_5967,N_5872);
xor U6997 (N_6997,N_5596,N_5457);
nor U6998 (N_6998,N_5315,N_5782);
nor U6999 (N_6999,N_5481,N_5315);
nand U7000 (N_7000,N_6698,N_6215);
and U7001 (N_7001,N_6543,N_6103);
nand U7002 (N_7002,N_6686,N_6405);
nor U7003 (N_7003,N_6579,N_6236);
nand U7004 (N_7004,N_6251,N_6800);
or U7005 (N_7005,N_6984,N_6211);
nand U7006 (N_7006,N_6998,N_6752);
nor U7007 (N_7007,N_6704,N_6390);
nand U7008 (N_7008,N_6824,N_6745);
nor U7009 (N_7009,N_6900,N_6261);
nor U7010 (N_7010,N_6365,N_6339);
and U7011 (N_7011,N_6217,N_6844);
or U7012 (N_7012,N_6239,N_6645);
and U7013 (N_7013,N_6833,N_6568);
xor U7014 (N_7014,N_6722,N_6626);
and U7015 (N_7015,N_6969,N_6266);
nand U7016 (N_7016,N_6385,N_6581);
and U7017 (N_7017,N_6601,N_6078);
nor U7018 (N_7018,N_6506,N_6249);
nand U7019 (N_7019,N_6308,N_6946);
xnor U7020 (N_7020,N_6286,N_6797);
xnor U7021 (N_7021,N_6038,N_6693);
xor U7022 (N_7022,N_6167,N_6348);
nor U7023 (N_7023,N_6003,N_6812);
nand U7024 (N_7024,N_6298,N_6886);
nand U7025 (N_7025,N_6632,N_6110);
and U7026 (N_7026,N_6245,N_6045);
nand U7027 (N_7027,N_6063,N_6054);
nor U7028 (N_7028,N_6403,N_6374);
nand U7029 (N_7029,N_6491,N_6004);
and U7030 (N_7030,N_6237,N_6960);
or U7031 (N_7031,N_6591,N_6860);
nor U7032 (N_7032,N_6639,N_6838);
nor U7033 (N_7033,N_6707,N_6633);
and U7034 (N_7034,N_6762,N_6387);
or U7035 (N_7035,N_6612,N_6642);
xor U7036 (N_7036,N_6470,N_6914);
nor U7037 (N_7037,N_6803,N_6573);
nor U7038 (N_7038,N_6848,N_6233);
nor U7039 (N_7039,N_6616,N_6561);
nor U7040 (N_7040,N_6257,N_6418);
or U7041 (N_7041,N_6501,N_6330);
nand U7042 (N_7042,N_6505,N_6148);
nand U7043 (N_7043,N_6867,N_6728);
nand U7044 (N_7044,N_6450,N_6185);
nor U7045 (N_7045,N_6893,N_6120);
xor U7046 (N_7046,N_6849,N_6615);
and U7047 (N_7047,N_6021,N_6278);
nand U7048 (N_7048,N_6794,N_6388);
or U7049 (N_7049,N_6084,N_6309);
nand U7050 (N_7050,N_6820,N_6143);
xor U7051 (N_7051,N_6892,N_6454);
nor U7052 (N_7052,N_6764,N_6293);
or U7053 (N_7053,N_6911,N_6191);
or U7054 (N_7054,N_6464,N_6182);
nand U7055 (N_7055,N_6953,N_6985);
or U7056 (N_7056,N_6748,N_6956);
or U7057 (N_7057,N_6509,N_6497);
nand U7058 (N_7058,N_6075,N_6052);
xnor U7059 (N_7059,N_6354,N_6066);
nor U7060 (N_7060,N_6146,N_6362);
xor U7061 (N_7061,N_6444,N_6877);
nor U7062 (N_7062,N_6888,N_6381);
xnor U7063 (N_7063,N_6687,N_6252);
nor U7064 (N_7064,N_6258,N_6917);
nand U7065 (N_7065,N_6739,N_6829);
and U7066 (N_7066,N_6993,N_6370);
nand U7067 (N_7067,N_6098,N_6119);
nor U7068 (N_7068,N_6578,N_6656);
nand U7069 (N_7069,N_6696,N_6475);
and U7070 (N_7070,N_6720,N_6706);
nand U7071 (N_7071,N_6708,N_6316);
nor U7072 (N_7072,N_6826,N_6876);
nor U7073 (N_7073,N_6015,N_6373);
or U7074 (N_7074,N_6600,N_6778);
and U7075 (N_7075,N_6662,N_6836);
or U7076 (N_7076,N_6093,N_6407);
and U7077 (N_7077,N_6436,N_6256);
nand U7078 (N_7078,N_6223,N_6253);
nand U7079 (N_7079,N_6187,N_6401);
and U7080 (N_7080,N_6856,N_6898);
nor U7081 (N_7081,N_6306,N_6839);
nor U7082 (N_7082,N_6209,N_6212);
nand U7083 (N_7083,N_6482,N_6392);
nor U7084 (N_7084,N_6446,N_6071);
nand U7085 (N_7085,N_6205,N_6344);
nand U7086 (N_7086,N_6942,N_6040);
or U7087 (N_7087,N_6636,N_6835);
or U7088 (N_7088,N_6731,N_6281);
and U7089 (N_7089,N_6398,N_6810);
or U7090 (N_7090,N_6654,N_6109);
and U7091 (N_7091,N_6978,N_6628);
nand U7092 (N_7092,N_6010,N_6831);
nand U7093 (N_7093,N_6840,N_6743);
or U7094 (N_7094,N_6496,N_6709);
and U7095 (N_7095,N_6235,N_6389);
or U7096 (N_7096,N_6524,N_6866);
nand U7097 (N_7097,N_6299,N_6129);
or U7098 (N_7098,N_6250,N_6819);
nand U7099 (N_7099,N_6366,N_6472);
and U7100 (N_7100,N_6283,N_6000);
or U7101 (N_7101,N_6772,N_6945);
and U7102 (N_7102,N_6319,N_6691);
nor U7103 (N_7103,N_6567,N_6882);
nor U7104 (N_7104,N_6260,N_6897);
xnor U7105 (N_7105,N_6666,N_6254);
nor U7106 (N_7106,N_6396,N_6044);
and U7107 (N_7107,N_6345,N_6268);
nand U7108 (N_7108,N_6150,N_6011);
or U7109 (N_7109,N_6913,N_6437);
and U7110 (N_7110,N_6463,N_6132);
nor U7111 (N_7111,N_6314,N_6466);
nand U7112 (N_7112,N_6342,N_6753);
nor U7113 (N_7113,N_6697,N_6548);
xor U7114 (N_7114,N_6959,N_6043);
or U7115 (N_7115,N_6777,N_6486);
nor U7116 (N_7116,N_6551,N_6380);
and U7117 (N_7117,N_6881,N_6830);
nand U7118 (N_7118,N_6779,N_6858);
nor U7119 (N_7119,N_6822,N_6188);
nor U7120 (N_7120,N_6972,N_6030);
or U7121 (N_7121,N_6163,N_6789);
or U7122 (N_7122,N_6766,N_6340);
and U7123 (N_7123,N_6775,N_6383);
nor U7124 (N_7124,N_6622,N_6134);
nand U7125 (N_7125,N_6242,N_6783);
nand U7126 (N_7126,N_6039,N_6028);
nand U7127 (N_7127,N_6008,N_6462);
or U7128 (N_7128,N_6750,N_6871);
and U7129 (N_7129,N_6417,N_6857);
nor U7130 (N_7130,N_6983,N_6801);
nor U7131 (N_7131,N_6790,N_6080);
or U7132 (N_7132,N_6767,N_6776);
and U7133 (N_7133,N_6199,N_6246);
nor U7134 (N_7134,N_6138,N_6979);
nand U7135 (N_7135,N_6473,N_6145);
xnor U7136 (N_7136,N_6657,N_6841);
nor U7137 (N_7137,N_6035,N_6869);
nor U7138 (N_7138,N_6599,N_6522);
or U7139 (N_7139,N_6087,N_6925);
and U7140 (N_7140,N_6863,N_6057);
and U7141 (N_7141,N_6310,N_6369);
nor U7142 (N_7142,N_6910,N_6349);
nor U7143 (N_7143,N_6602,N_6048);
nor U7144 (N_7144,N_6156,N_6516);
nor U7145 (N_7145,N_6255,N_6029);
xor U7146 (N_7146,N_6042,N_6224);
and U7147 (N_7147,N_6170,N_6695);
and U7148 (N_7148,N_6670,N_6449);
nor U7149 (N_7149,N_6901,N_6807);
and U7150 (N_7150,N_6603,N_6174);
or U7151 (N_7151,N_6429,N_6701);
or U7152 (N_7152,N_6685,N_6872);
and U7153 (N_7153,N_6041,N_6500);
and U7154 (N_7154,N_6991,N_6555);
nor U7155 (N_7155,N_6711,N_6977);
and U7156 (N_7156,N_6171,N_6336);
or U7157 (N_7157,N_6435,N_6202);
nor U7158 (N_7158,N_6438,N_6853);
nor U7159 (N_7159,N_6520,N_6510);
nand U7160 (N_7160,N_6915,N_6890);
and U7161 (N_7161,N_6355,N_6937);
nand U7162 (N_7162,N_6391,N_6741);
xor U7163 (N_7163,N_6154,N_6232);
nand U7164 (N_7164,N_6318,N_6056);
or U7165 (N_7165,N_6049,N_6606);
or U7166 (N_7166,N_6575,N_6372);
nor U7167 (N_7167,N_6175,N_6586);
nor U7168 (N_7168,N_6907,N_6448);
nor U7169 (N_7169,N_6584,N_6082);
and U7170 (N_7170,N_6733,N_6465);
nor U7171 (N_7171,N_6992,N_6494);
nor U7172 (N_7172,N_6289,N_6222);
xnor U7173 (N_7173,N_6854,N_6196);
nor U7174 (N_7174,N_6664,N_6271);
and U7175 (N_7175,N_6288,N_6924);
or U7176 (N_7176,N_6136,N_6069);
xor U7177 (N_7177,N_6141,N_6195);
xor U7178 (N_7178,N_6988,N_6780);
or U7179 (N_7179,N_6804,N_6311);
nor U7180 (N_7180,N_6007,N_6483);
nand U7181 (N_7181,N_6851,N_6144);
nor U7182 (N_7182,N_6047,N_6507);
nor U7183 (N_7183,N_6891,N_6495);
nor U7184 (N_7184,N_6105,N_6763);
and U7185 (N_7185,N_6430,N_6447);
xnor U7186 (N_7186,N_6903,N_6719);
or U7187 (N_7187,N_6880,N_6861);
or U7188 (N_7188,N_6453,N_6798);
nor U7189 (N_7189,N_6213,N_6059);
nand U7190 (N_7190,N_6926,N_6458);
nand U7191 (N_7191,N_6884,N_6557);
and U7192 (N_7192,N_6050,N_6131);
or U7193 (N_7193,N_6104,N_6062);
or U7194 (N_7194,N_6574,N_6658);
or U7195 (N_7195,N_6668,N_6186);
nor U7196 (N_7196,N_6569,N_6335);
nand U7197 (N_7197,N_6220,N_6096);
nor U7198 (N_7198,N_6139,N_6259);
and U7199 (N_7199,N_6729,N_6244);
nand U7200 (N_7200,N_6346,N_6845);
nor U7201 (N_7201,N_6016,N_6815);
or U7202 (N_7202,N_6808,N_6802);
and U7203 (N_7203,N_6712,N_6963);
nand U7204 (N_7204,N_6558,N_6406);
nor U7205 (N_7205,N_6634,N_6547);
xnor U7206 (N_7206,N_6416,N_6751);
and U7207 (N_7207,N_6981,N_6617);
nand U7208 (N_7208,N_6582,N_6895);
and U7209 (N_7209,N_6530,N_6031);
xor U7210 (N_7210,N_6147,N_6967);
or U7211 (N_7211,N_6452,N_6460);
or U7212 (N_7212,N_6002,N_6535);
nor U7213 (N_7213,N_6116,N_6420);
xor U7214 (N_7214,N_6275,N_6122);
nand U7215 (N_7215,N_6787,N_6760);
and U7216 (N_7216,N_6843,N_6534);
or U7217 (N_7217,N_6512,N_6742);
nand U7218 (N_7218,N_6994,N_6596);
and U7219 (N_7219,N_6208,N_6537);
nor U7220 (N_7220,N_6688,N_6672);
and U7221 (N_7221,N_6832,N_6594);
nand U7222 (N_7222,N_6367,N_6061);
and U7223 (N_7223,N_6409,N_6734);
or U7224 (N_7224,N_6746,N_6546);
or U7225 (N_7225,N_6083,N_6936);
and U7226 (N_7226,N_6651,N_6717);
xor U7227 (N_7227,N_6284,N_6912);
nand U7228 (N_7228,N_6627,N_6210);
nand U7229 (N_7229,N_6181,N_6100);
and U7230 (N_7230,N_6929,N_6592);
or U7231 (N_7231,N_6587,N_6177);
nand U7232 (N_7232,N_6456,N_6487);
or U7233 (N_7233,N_6037,N_6590);
nor U7234 (N_7234,N_6060,N_6230);
xor U7235 (N_7235,N_6559,N_6878);
nor U7236 (N_7236,N_6142,N_6492);
and U7237 (N_7237,N_6908,N_6939);
nor U7238 (N_7238,N_6736,N_6655);
or U7239 (N_7239,N_6221,N_6611);
nor U7240 (N_7240,N_6428,N_6862);
nor U7241 (N_7241,N_6153,N_6508);
or U7242 (N_7242,N_6353,N_6513);
nand U7243 (N_7243,N_6542,N_6677);
nor U7244 (N_7244,N_6192,N_6846);
nor U7245 (N_7245,N_6184,N_6480);
nor U7246 (N_7246,N_6997,N_6646);
nand U7247 (N_7247,N_6713,N_6650);
xor U7248 (N_7248,N_6784,N_6905);
nand U7249 (N_7249,N_6757,N_6619);
nor U7250 (N_7250,N_6197,N_6478);
or U7251 (N_7251,N_6887,N_6644);
xnor U7252 (N_7252,N_6160,N_6613);
nand U7253 (N_7253,N_6287,N_6539);
and U7254 (N_7254,N_6541,N_6768);
or U7255 (N_7255,N_6352,N_6243);
and U7256 (N_7256,N_6540,N_6005);
and U7257 (N_7257,N_6471,N_6999);
and U7258 (N_7258,N_6957,N_6921);
and U7259 (N_7259,N_6785,N_6827);
and U7260 (N_7260,N_6502,N_6950);
xor U7261 (N_7261,N_6609,N_6771);
and U7262 (N_7262,N_6598,N_6324);
and U7263 (N_7263,N_6386,N_6665);
nor U7264 (N_7264,N_6941,N_6358);
nor U7265 (N_7265,N_6976,N_6681);
and U7266 (N_7266,N_6621,N_6427);
nand U7267 (N_7267,N_6629,N_6770);
nand U7268 (N_7268,N_6519,N_6928);
nand U7269 (N_7269,N_6393,N_6111);
nand U7270 (N_7270,N_6818,N_6809);
nor U7271 (N_7271,N_6269,N_6415);
nand U7272 (N_7272,N_6097,N_6904);
and U7273 (N_7273,N_6842,N_6610);
nand U7274 (N_7274,N_6285,N_6282);
or U7275 (N_7275,N_6326,N_6490);
and U7276 (N_7276,N_6828,N_6019);
xor U7277 (N_7277,N_6576,N_6813);
and U7278 (N_7278,N_6067,N_6341);
nand U7279 (N_7279,N_6761,N_6457);
xnor U7280 (N_7280,N_6200,N_6909);
xor U7281 (N_7281,N_6248,N_6273);
nand U7282 (N_7282,N_6414,N_6749);
and U7283 (N_7283,N_6423,N_6489);
xor U7284 (N_7284,N_6012,N_6680);
or U7285 (N_7285,N_6678,N_6943);
nand U7286 (N_7286,N_6441,N_6765);
and U7287 (N_7287,N_6889,N_6025);
nor U7288 (N_7288,N_6321,N_6952);
or U7289 (N_7289,N_6206,N_6618);
and U7290 (N_7290,N_6408,N_6837);
nand U7291 (N_7291,N_6238,N_6161);
and U7292 (N_7292,N_6477,N_6975);
nor U7293 (N_7293,N_6550,N_6026);
nand U7294 (N_7294,N_6605,N_6874);
or U7295 (N_7295,N_6363,N_6511);
and U7296 (N_7296,N_6570,N_6305);
xnor U7297 (N_7297,N_6679,N_6536);
or U7298 (N_7298,N_6690,N_6865);
nand U7299 (N_7299,N_6431,N_6689);
and U7300 (N_7300,N_6528,N_6811);
or U7301 (N_7301,N_6461,N_6549);
nand U7302 (N_7302,N_6919,N_6614);
nor U7303 (N_7303,N_6443,N_6424);
xor U7304 (N_7304,N_6973,N_6518);
nor U7305 (N_7305,N_6323,N_6128);
xor U7306 (N_7306,N_6079,N_6394);
and U7307 (N_7307,N_6661,N_6034);
or U7308 (N_7308,N_6379,N_6737);
nor U7309 (N_7309,N_6364,N_6726);
nand U7310 (N_7310,N_6955,N_6724);
nand U7311 (N_7311,N_6411,N_6747);
or U7312 (N_7312,N_6607,N_6404);
or U7313 (N_7313,N_6328,N_6126);
or U7314 (N_7314,N_6343,N_6117);
or U7315 (N_7315,N_6902,N_6873);
xor U7316 (N_7316,N_6203,N_6674);
or U7317 (N_7317,N_6413,N_6479);
and U7318 (N_7318,N_6759,N_6152);
and U7319 (N_7319,N_6572,N_6938);
nand U7320 (N_7320,N_6375,N_6327);
nor U7321 (N_7321,N_6920,N_6225);
and U7322 (N_7322,N_6755,N_6357);
xnor U7323 (N_7323,N_6868,N_6013);
nor U7324 (N_7324,N_6402,N_6521);
nor U7325 (N_7325,N_6799,N_6962);
and U7326 (N_7326,N_6421,N_6730);
nand U7327 (N_7327,N_6108,N_6927);
and U7328 (N_7328,N_6556,N_6320);
and U7329 (N_7329,N_6190,N_6964);
nand U7330 (N_7330,N_6683,N_6334);
or U7331 (N_7331,N_6371,N_6422);
nor U7332 (N_7332,N_6638,N_6085);
or U7333 (N_7333,N_6870,N_6292);
and U7334 (N_7334,N_6932,N_6137);
xor U7335 (N_7335,N_6425,N_6183);
nor U7336 (N_7336,N_6162,N_6313);
or U7337 (N_7337,N_6459,N_6935);
and U7338 (N_7338,N_6155,N_6947);
and U7339 (N_7339,N_6089,N_6064);
nand U7340 (N_7340,N_6961,N_6648);
nor U7341 (N_7341,N_6032,N_6692);
nand U7342 (N_7342,N_6980,N_6127);
nand U7343 (N_7343,N_6700,N_6971);
xor U7344 (N_7344,N_6280,N_6296);
nand U7345 (N_7345,N_6671,N_6159);
or U7346 (N_7346,N_6538,N_6172);
and U7347 (N_7347,N_6635,N_6023);
xor U7348 (N_7348,N_6276,N_6279);
and U7349 (N_7349,N_6589,N_6474);
or U7350 (N_7350,N_6219,N_6652);
and U7351 (N_7351,N_6916,N_6118);
xnor U7352 (N_7352,N_6774,N_6451);
and U7353 (N_7353,N_6982,N_6263);
xnor U7354 (N_7354,N_6165,N_6329);
nor U7355 (N_7355,N_6918,N_6970);
nand U7356 (N_7356,N_6485,N_6356);
nand U7357 (N_7357,N_6958,N_6124);
and U7358 (N_7358,N_6906,N_6554);
nor U7359 (N_7359,N_6732,N_6095);
and U7360 (N_7360,N_6699,N_6229);
xor U7361 (N_7361,N_6498,N_6267);
and U7362 (N_7362,N_6989,N_6740);
and U7363 (N_7363,N_6930,N_6940);
nor U7364 (N_7364,N_6262,N_6673);
or U7365 (N_7365,N_6168,N_6608);
nand U7366 (N_7366,N_6410,N_6986);
nor U7367 (N_7367,N_6481,N_6382);
or U7368 (N_7368,N_6455,N_6725);
nand U7369 (N_7369,N_6265,N_6158);
nor U7370 (N_7370,N_6966,N_6552);
nor U7371 (N_7371,N_6659,N_6623);
nor U7372 (N_7372,N_6504,N_6001);
and U7373 (N_7373,N_6377,N_6176);
nand U7374 (N_7374,N_6566,N_6426);
or U7375 (N_7375,N_6684,N_6376);
nor U7376 (N_7376,N_6499,N_6164);
nor U7377 (N_7377,N_6036,N_6805);
or U7378 (N_7378,N_6133,N_6715);
and U7379 (N_7379,N_6527,N_6051);
nand U7380 (N_7380,N_6068,N_6018);
nor U7381 (N_7381,N_6081,N_6476);
nand U7382 (N_7382,N_6675,N_6545);
nor U7383 (N_7383,N_6304,N_6332);
or U7384 (N_7384,N_6247,N_6796);
nor U7385 (N_7385,N_6562,N_6922);
nor U7386 (N_7386,N_6523,N_6710);
nor U7387 (N_7387,N_6821,N_6337);
nor U7388 (N_7388,N_6620,N_6317);
nand U7389 (N_7389,N_6140,N_6643);
nand U7390 (N_7390,N_6351,N_6834);
and U7391 (N_7391,N_6359,N_6149);
and U7392 (N_7392,N_6580,N_6577);
xor U7393 (N_7393,N_6113,N_6923);
nor U7394 (N_7394,N_6291,N_6218);
xor U7395 (N_7395,N_6467,N_6397);
and U7396 (N_7396,N_6315,N_6272);
xor U7397 (N_7397,N_6151,N_6951);
nand U7398 (N_7398,N_6974,N_6526);
and U7399 (N_7399,N_6274,N_6663);
nand U7400 (N_7400,N_6954,N_6855);
nand U7401 (N_7401,N_6434,N_6123);
or U7402 (N_7402,N_6076,N_6440);
nand U7403 (N_7403,N_6702,N_6864);
and U7404 (N_7404,N_6020,N_6361);
xor U7405 (N_7405,N_6055,N_6825);
nand U7406 (N_7406,N_6157,N_6009);
nand U7407 (N_7407,N_6086,N_6077);
xnor U7408 (N_7408,N_6640,N_6852);
or U7409 (N_7409,N_6121,N_6791);
nor U7410 (N_7410,N_6676,N_6788);
or U7411 (N_7411,N_6234,N_6583);
nand U7412 (N_7412,N_6107,N_6301);
nand U7413 (N_7413,N_6703,N_6585);
and U7414 (N_7414,N_6027,N_6207);
xor U7415 (N_7415,N_6944,N_6968);
nor U7416 (N_7416,N_6816,N_6216);
and U7417 (N_7417,N_6948,N_6934);
nor U7418 (N_7418,N_6488,N_6295);
or U7419 (N_7419,N_6115,N_6338);
and U7420 (N_7420,N_6419,N_6017);
and U7421 (N_7421,N_6647,N_6694);
xor U7422 (N_7422,N_6649,N_6933);
and U7423 (N_7423,N_6294,N_6046);
nor U7424 (N_7424,N_6931,N_6065);
and U7425 (N_7425,N_6588,N_6102);
and U7426 (N_7426,N_6006,N_6368);
and U7427 (N_7427,N_6718,N_6723);
xnor U7428 (N_7428,N_6300,N_6899);
nand U7429 (N_7429,N_6094,N_6439);
nand U7430 (N_7430,N_6312,N_6302);
nand U7431 (N_7431,N_6503,N_6194);
and U7432 (N_7432,N_6073,N_6885);
nand U7433 (N_7433,N_6987,N_6226);
nor U7434 (N_7434,N_6099,N_6179);
nand U7435 (N_7435,N_6178,N_6637);
and U7436 (N_7436,N_6625,N_6201);
nor U7437 (N_7437,N_6641,N_6773);
and U7438 (N_7438,N_6756,N_6277);
nand U7439 (N_7439,N_6735,N_6597);
or U7440 (N_7440,N_6024,N_6493);
xor U7441 (N_7441,N_6850,N_6669);
nor U7442 (N_7442,N_6544,N_6173);
or U7443 (N_7443,N_6525,N_6814);
or U7444 (N_7444,N_6270,N_6563);
or U7445 (N_7445,N_6445,N_6331);
or U7446 (N_7446,N_6074,N_6995);
xnor U7447 (N_7447,N_6727,N_6879);
nor U7448 (N_7448,N_6896,N_6180);
or U7449 (N_7449,N_6307,N_6297);
nor U7450 (N_7450,N_6198,N_6604);
and U7451 (N_7451,N_6264,N_6241);
or U7452 (N_7452,N_6092,N_6795);
or U7453 (N_7453,N_6228,N_6949);
and U7454 (N_7454,N_6412,N_6721);
and U7455 (N_7455,N_6469,N_6769);
nor U7456 (N_7456,N_6758,N_6378);
nor U7457 (N_7457,N_6514,N_6135);
nand U7458 (N_7458,N_6014,N_6705);
nand U7459 (N_7459,N_6593,N_6360);
or U7460 (N_7460,N_6738,N_6806);
nand U7461 (N_7461,N_6792,N_6214);
and U7462 (N_7462,N_6101,N_6847);
and U7463 (N_7463,N_6682,N_6240);
and U7464 (N_7464,N_6130,N_6894);
xor U7465 (N_7465,N_6817,N_6624);
and U7466 (N_7466,N_6532,N_6660);
or U7467 (N_7467,N_6204,N_6531);
nand U7468 (N_7468,N_6823,N_6189);
or U7469 (N_7469,N_6303,N_6786);
nand U7470 (N_7470,N_6072,N_6529);
nand U7471 (N_7471,N_6565,N_6560);
or U7472 (N_7472,N_6169,N_6564);
nor U7473 (N_7473,N_6106,N_6347);
nor U7474 (N_7474,N_6395,N_6781);
and U7475 (N_7475,N_6965,N_6166);
nand U7476 (N_7476,N_6112,N_6990);
or U7477 (N_7477,N_6442,N_6553);
xnor U7478 (N_7478,N_6290,N_6754);
nand U7479 (N_7479,N_6595,N_6744);
nand U7480 (N_7480,N_6058,N_6515);
nor U7481 (N_7481,N_6333,N_6400);
nor U7482 (N_7482,N_6468,N_6875);
xnor U7483 (N_7483,N_6517,N_6325);
nand U7484 (N_7484,N_6033,N_6667);
nor U7485 (N_7485,N_6091,N_6090);
and U7486 (N_7486,N_6231,N_6782);
nand U7487 (N_7487,N_6432,N_6533);
or U7488 (N_7488,N_6322,N_6399);
xor U7489 (N_7489,N_6053,N_6114);
nand U7490 (N_7490,N_6653,N_6793);
nand U7491 (N_7491,N_6883,N_6125);
or U7492 (N_7492,N_6384,N_6859);
or U7493 (N_7493,N_6350,N_6227);
and U7494 (N_7494,N_6716,N_6484);
and U7495 (N_7495,N_6088,N_6571);
nand U7496 (N_7496,N_6070,N_6433);
nand U7497 (N_7497,N_6714,N_6631);
nor U7498 (N_7498,N_6022,N_6630);
or U7499 (N_7499,N_6193,N_6996);
or U7500 (N_7500,N_6256,N_6399);
nor U7501 (N_7501,N_6664,N_6028);
nand U7502 (N_7502,N_6285,N_6712);
nand U7503 (N_7503,N_6681,N_6780);
xnor U7504 (N_7504,N_6257,N_6849);
and U7505 (N_7505,N_6376,N_6803);
nor U7506 (N_7506,N_6783,N_6776);
nand U7507 (N_7507,N_6678,N_6898);
and U7508 (N_7508,N_6597,N_6702);
nor U7509 (N_7509,N_6047,N_6362);
xnor U7510 (N_7510,N_6115,N_6856);
or U7511 (N_7511,N_6537,N_6302);
and U7512 (N_7512,N_6480,N_6452);
xnor U7513 (N_7513,N_6813,N_6681);
or U7514 (N_7514,N_6561,N_6808);
and U7515 (N_7515,N_6334,N_6850);
or U7516 (N_7516,N_6651,N_6661);
nand U7517 (N_7517,N_6753,N_6487);
or U7518 (N_7518,N_6262,N_6747);
nor U7519 (N_7519,N_6084,N_6092);
xor U7520 (N_7520,N_6907,N_6210);
and U7521 (N_7521,N_6439,N_6772);
nand U7522 (N_7522,N_6814,N_6118);
or U7523 (N_7523,N_6575,N_6343);
nand U7524 (N_7524,N_6326,N_6568);
nand U7525 (N_7525,N_6199,N_6133);
and U7526 (N_7526,N_6286,N_6205);
nand U7527 (N_7527,N_6640,N_6771);
nor U7528 (N_7528,N_6103,N_6771);
nand U7529 (N_7529,N_6367,N_6170);
and U7530 (N_7530,N_6179,N_6645);
nand U7531 (N_7531,N_6672,N_6945);
xnor U7532 (N_7532,N_6528,N_6110);
and U7533 (N_7533,N_6177,N_6690);
nor U7534 (N_7534,N_6578,N_6119);
and U7535 (N_7535,N_6873,N_6249);
xor U7536 (N_7536,N_6146,N_6703);
and U7537 (N_7537,N_6474,N_6765);
xor U7538 (N_7538,N_6168,N_6046);
or U7539 (N_7539,N_6817,N_6329);
or U7540 (N_7540,N_6834,N_6405);
and U7541 (N_7541,N_6296,N_6062);
and U7542 (N_7542,N_6981,N_6524);
nor U7543 (N_7543,N_6785,N_6823);
and U7544 (N_7544,N_6476,N_6600);
or U7545 (N_7545,N_6821,N_6128);
nor U7546 (N_7546,N_6187,N_6774);
nor U7547 (N_7547,N_6589,N_6535);
or U7548 (N_7548,N_6611,N_6619);
and U7549 (N_7549,N_6176,N_6427);
xnor U7550 (N_7550,N_6395,N_6328);
nor U7551 (N_7551,N_6995,N_6276);
nor U7552 (N_7552,N_6724,N_6337);
nor U7553 (N_7553,N_6956,N_6019);
nand U7554 (N_7554,N_6318,N_6023);
or U7555 (N_7555,N_6584,N_6359);
nor U7556 (N_7556,N_6528,N_6169);
or U7557 (N_7557,N_6722,N_6529);
or U7558 (N_7558,N_6061,N_6377);
nor U7559 (N_7559,N_6443,N_6665);
or U7560 (N_7560,N_6777,N_6476);
or U7561 (N_7561,N_6106,N_6851);
nor U7562 (N_7562,N_6591,N_6634);
or U7563 (N_7563,N_6393,N_6338);
nand U7564 (N_7564,N_6368,N_6287);
and U7565 (N_7565,N_6102,N_6552);
nor U7566 (N_7566,N_6894,N_6971);
and U7567 (N_7567,N_6035,N_6440);
and U7568 (N_7568,N_6433,N_6841);
and U7569 (N_7569,N_6351,N_6149);
nor U7570 (N_7570,N_6610,N_6757);
nor U7571 (N_7571,N_6595,N_6010);
or U7572 (N_7572,N_6690,N_6038);
and U7573 (N_7573,N_6327,N_6647);
nor U7574 (N_7574,N_6944,N_6425);
xnor U7575 (N_7575,N_6838,N_6853);
or U7576 (N_7576,N_6157,N_6115);
or U7577 (N_7577,N_6944,N_6004);
nor U7578 (N_7578,N_6679,N_6094);
nand U7579 (N_7579,N_6901,N_6750);
or U7580 (N_7580,N_6355,N_6423);
and U7581 (N_7581,N_6317,N_6785);
and U7582 (N_7582,N_6158,N_6461);
or U7583 (N_7583,N_6197,N_6556);
nand U7584 (N_7584,N_6167,N_6985);
and U7585 (N_7585,N_6322,N_6695);
or U7586 (N_7586,N_6747,N_6751);
nand U7587 (N_7587,N_6784,N_6982);
nor U7588 (N_7588,N_6886,N_6623);
nand U7589 (N_7589,N_6995,N_6668);
and U7590 (N_7590,N_6508,N_6261);
or U7591 (N_7591,N_6478,N_6808);
and U7592 (N_7592,N_6062,N_6555);
or U7593 (N_7593,N_6036,N_6615);
nand U7594 (N_7594,N_6239,N_6490);
xnor U7595 (N_7595,N_6159,N_6027);
nand U7596 (N_7596,N_6440,N_6466);
nand U7597 (N_7597,N_6969,N_6606);
or U7598 (N_7598,N_6110,N_6500);
nor U7599 (N_7599,N_6084,N_6434);
nor U7600 (N_7600,N_6964,N_6105);
nand U7601 (N_7601,N_6088,N_6794);
nor U7602 (N_7602,N_6189,N_6229);
nor U7603 (N_7603,N_6680,N_6002);
xor U7604 (N_7604,N_6463,N_6596);
nor U7605 (N_7605,N_6953,N_6833);
and U7606 (N_7606,N_6862,N_6189);
or U7607 (N_7607,N_6558,N_6585);
and U7608 (N_7608,N_6287,N_6561);
and U7609 (N_7609,N_6874,N_6908);
or U7610 (N_7610,N_6587,N_6959);
nand U7611 (N_7611,N_6687,N_6392);
nor U7612 (N_7612,N_6609,N_6434);
and U7613 (N_7613,N_6083,N_6721);
or U7614 (N_7614,N_6216,N_6587);
nor U7615 (N_7615,N_6389,N_6847);
or U7616 (N_7616,N_6462,N_6799);
nand U7617 (N_7617,N_6784,N_6693);
and U7618 (N_7618,N_6078,N_6068);
nand U7619 (N_7619,N_6242,N_6344);
or U7620 (N_7620,N_6694,N_6655);
and U7621 (N_7621,N_6908,N_6895);
nand U7622 (N_7622,N_6119,N_6156);
nor U7623 (N_7623,N_6938,N_6369);
and U7624 (N_7624,N_6884,N_6824);
or U7625 (N_7625,N_6360,N_6160);
and U7626 (N_7626,N_6520,N_6831);
and U7627 (N_7627,N_6054,N_6828);
nand U7628 (N_7628,N_6882,N_6415);
nor U7629 (N_7629,N_6456,N_6087);
nand U7630 (N_7630,N_6102,N_6386);
nand U7631 (N_7631,N_6827,N_6824);
and U7632 (N_7632,N_6955,N_6205);
or U7633 (N_7633,N_6474,N_6226);
nand U7634 (N_7634,N_6075,N_6379);
and U7635 (N_7635,N_6375,N_6289);
and U7636 (N_7636,N_6256,N_6038);
nand U7637 (N_7637,N_6356,N_6134);
xnor U7638 (N_7638,N_6012,N_6948);
nor U7639 (N_7639,N_6564,N_6921);
nor U7640 (N_7640,N_6616,N_6671);
and U7641 (N_7641,N_6479,N_6330);
nand U7642 (N_7642,N_6607,N_6755);
or U7643 (N_7643,N_6395,N_6840);
nor U7644 (N_7644,N_6285,N_6644);
and U7645 (N_7645,N_6215,N_6020);
or U7646 (N_7646,N_6481,N_6290);
or U7647 (N_7647,N_6872,N_6405);
nor U7648 (N_7648,N_6002,N_6571);
or U7649 (N_7649,N_6234,N_6834);
nand U7650 (N_7650,N_6398,N_6659);
nor U7651 (N_7651,N_6572,N_6083);
and U7652 (N_7652,N_6629,N_6068);
and U7653 (N_7653,N_6149,N_6943);
and U7654 (N_7654,N_6857,N_6185);
xnor U7655 (N_7655,N_6417,N_6631);
nor U7656 (N_7656,N_6498,N_6871);
nor U7657 (N_7657,N_6640,N_6589);
nand U7658 (N_7658,N_6280,N_6852);
xor U7659 (N_7659,N_6290,N_6892);
or U7660 (N_7660,N_6258,N_6339);
nand U7661 (N_7661,N_6367,N_6155);
xnor U7662 (N_7662,N_6951,N_6597);
and U7663 (N_7663,N_6986,N_6697);
and U7664 (N_7664,N_6866,N_6955);
nor U7665 (N_7665,N_6601,N_6289);
nor U7666 (N_7666,N_6670,N_6781);
nand U7667 (N_7667,N_6794,N_6247);
or U7668 (N_7668,N_6715,N_6155);
or U7669 (N_7669,N_6487,N_6777);
and U7670 (N_7670,N_6643,N_6367);
nand U7671 (N_7671,N_6744,N_6298);
nand U7672 (N_7672,N_6456,N_6994);
or U7673 (N_7673,N_6740,N_6657);
xnor U7674 (N_7674,N_6523,N_6365);
and U7675 (N_7675,N_6454,N_6462);
or U7676 (N_7676,N_6327,N_6398);
nor U7677 (N_7677,N_6355,N_6400);
or U7678 (N_7678,N_6372,N_6631);
nor U7679 (N_7679,N_6440,N_6351);
nand U7680 (N_7680,N_6604,N_6592);
or U7681 (N_7681,N_6200,N_6591);
nand U7682 (N_7682,N_6711,N_6202);
xnor U7683 (N_7683,N_6842,N_6307);
or U7684 (N_7684,N_6195,N_6198);
and U7685 (N_7685,N_6706,N_6745);
and U7686 (N_7686,N_6904,N_6412);
nand U7687 (N_7687,N_6445,N_6320);
and U7688 (N_7688,N_6511,N_6303);
xor U7689 (N_7689,N_6123,N_6253);
nand U7690 (N_7690,N_6557,N_6449);
nand U7691 (N_7691,N_6867,N_6830);
nand U7692 (N_7692,N_6082,N_6789);
or U7693 (N_7693,N_6183,N_6692);
nand U7694 (N_7694,N_6582,N_6029);
and U7695 (N_7695,N_6729,N_6310);
xor U7696 (N_7696,N_6762,N_6260);
nand U7697 (N_7697,N_6154,N_6688);
or U7698 (N_7698,N_6566,N_6181);
or U7699 (N_7699,N_6038,N_6120);
nand U7700 (N_7700,N_6809,N_6609);
nand U7701 (N_7701,N_6568,N_6358);
or U7702 (N_7702,N_6531,N_6089);
nand U7703 (N_7703,N_6229,N_6557);
or U7704 (N_7704,N_6573,N_6295);
and U7705 (N_7705,N_6783,N_6619);
nand U7706 (N_7706,N_6548,N_6657);
nand U7707 (N_7707,N_6218,N_6154);
and U7708 (N_7708,N_6507,N_6613);
nor U7709 (N_7709,N_6136,N_6070);
xor U7710 (N_7710,N_6046,N_6948);
and U7711 (N_7711,N_6070,N_6853);
or U7712 (N_7712,N_6563,N_6387);
nor U7713 (N_7713,N_6261,N_6965);
nand U7714 (N_7714,N_6673,N_6547);
nor U7715 (N_7715,N_6261,N_6599);
or U7716 (N_7716,N_6820,N_6726);
nand U7717 (N_7717,N_6784,N_6282);
and U7718 (N_7718,N_6943,N_6425);
and U7719 (N_7719,N_6584,N_6372);
nand U7720 (N_7720,N_6625,N_6018);
and U7721 (N_7721,N_6904,N_6557);
or U7722 (N_7722,N_6430,N_6120);
and U7723 (N_7723,N_6090,N_6044);
nand U7724 (N_7724,N_6309,N_6478);
nor U7725 (N_7725,N_6610,N_6948);
or U7726 (N_7726,N_6130,N_6461);
and U7727 (N_7727,N_6916,N_6077);
nand U7728 (N_7728,N_6376,N_6501);
and U7729 (N_7729,N_6260,N_6292);
xor U7730 (N_7730,N_6911,N_6278);
nor U7731 (N_7731,N_6197,N_6104);
or U7732 (N_7732,N_6487,N_6588);
xor U7733 (N_7733,N_6274,N_6418);
nand U7734 (N_7734,N_6842,N_6304);
and U7735 (N_7735,N_6337,N_6986);
xor U7736 (N_7736,N_6258,N_6778);
or U7737 (N_7737,N_6062,N_6999);
and U7738 (N_7738,N_6145,N_6899);
or U7739 (N_7739,N_6779,N_6693);
or U7740 (N_7740,N_6052,N_6267);
or U7741 (N_7741,N_6762,N_6614);
nor U7742 (N_7742,N_6417,N_6299);
nand U7743 (N_7743,N_6994,N_6532);
nor U7744 (N_7744,N_6013,N_6066);
and U7745 (N_7745,N_6665,N_6782);
or U7746 (N_7746,N_6381,N_6689);
nor U7747 (N_7747,N_6297,N_6373);
or U7748 (N_7748,N_6615,N_6014);
nor U7749 (N_7749,N_6182,N_6282);
nor U7750 (N_7750,N_6463,N_6710);
xnor U7751 (N_7751,N_6083,N_6840);
and U7752 (N_7752,N_6181,N_6288);
and U7753 (N_7753,N_6988,N_6121);
or U7754 (N_7754,N_6655,N_6909);
and U7755 (N_7755,N_6469,N_6795);
nor U7756 (N_7756,N_6170,N_6239);
and U7757 (N_7757,N_6617,N_6854);
and U7758 (N_7758,N_6553,N_6890);
nand U7759 (N_7759,N_6809,N_6995);
and U7760 (N_7760,N_6790,N_6825);
and U7761 (N_7761,N_6195,N_6296);
or U7762 (N_7762,N_6793,N_6926);
nand U7763 (N_7763,N_6645,N_6378);
and U7764 (N_7764,N_6363,N_6685);
nor U7765 (N_7765,N_6536,N_6117);
and U7766 (N_7766,N_6179,N_6030);
nand U7767 (N_7767,N_6580,N_6530);
or U7768 (N_7768,N_6088,N_6617);
nor U7769 (N_7769,N_6957,N_6415);
nand U7770 (N_7770,N_6031,N_6441);
and U7771 (N_7771,N_6174,N_6645);
and U7772 (N_7772,N_6220,N_6070);
nor U7773 (N_7773,N_6303,N_6277);
nand U7774 (N_7774,N_6464,N_6976);
nand U7775 (N_7775,N_6364,N_6847);
nand U7776 (N_7776,N_6858,N_6835);
xnor U7777 (N_7777,N_6828,N_6907);
xnor U7778 (N_7778,N_6127,N_6968);
and U7779 (N_7779,N_6968,N_6623);
nor U7780 (N_7780,N_6105,N_6775);
xnor U7781 (N_7781,N_6393,N_6048);
and U7782 (N_7782,N_6307,N_6924);
nand U7783 (N_7783,N_6919,N_6215);
and U7784 (N_7784,N_6160,N_6078);
nand U7785 (N_7785,N_6798,N_6487);
nand U7786 (N_7786,N_6466,N_6479);
and U7787 (N_7787,N_6806,N_6169);
nand U7788 (N_7788,N_6416,N_6196);
or U7789 (N_7789,N_6193,N_6005);
nor U7790 (N_7790,N_6684,N_6453);
nand U7791 (N_7791,N_6458,N_6625);
and U7792 (N_7792,N_6732,N_6217);
and U7793 (N_7793,N_6296,N_6736);
nand U7794 (N_7794,N_6305,N_6597);
xnor U7795 (N_7795,N_6674,N_6356);
nand U7796 (N_7796,N_6046,N_6348);
or U7797 (N_7797,N_6291,N_6568);
nor U7798 (N_7798,N_6875,N_6279);
and U7799 (N_7799,N_6870,N_6555);
xor U7800 (N_7800,N_6391,N_6819);
nor U7801 (N_7801,N_6981,N_6501);
nand U7802 (N_7802,N_6063,N_6282);
and U7803 (N_7803,N_6747,N_6119);
or U7804 (N_7804,N_6152,N_6827);
or U7805 (N_7805,N_6495,N_6998);
and U7806 (N_7806,N_6480,N_6200);
nor U7807 (N_7807,N_6101,N_6889);
nand U7808 (N_7808,N_6787,N_6395);
or U7809 (N_7809,N_6625,N_6173);
or U7810 (N_7810,N_6794,N_6750);
or U7811 (N_7811,N_6323,N_6650);
or U7812 (N_7812,N_6148,N_6135);
and U7813 (N_7813,N_6963,N_6175);
nor U7814 (N_7814,N_6789,N_6663);
and U7815 (N_7815,N_6831,N_6298);
and U7816 (N_7816,N_6247,N_6810);
nand U7817 (N_7817,N_6408,N_6329);
nand U7818 (N_7818,N_6720,N_6665);
nand U7819 (N_7819,N_6673,N_6911);
nand U7820 (N_7820,N_6476,N_6623);
nor U7821 (N_7821,N_6462,N_6450);
nand U7822 (N_7822,N_6177,N_6920);
nor U7823 (N_7823,N_6623,N_6410);
xnor U7824 (N_7824,N_6864,N_6372);
or U7825 (N_7825,N_6667,N_6550);
nor U7826 (N_7826,N_6409,N_6266);
nor U7827 (N_7827,N_6159,N_6693);
nand U7828 (N_7828,N_6577,N_6030);
nand U7829 (N_7829,N_6009,N_6693);
or U7830 (N_7830,N_6746,N_6724);
nor U7831 (N_7831,N_6445,N_6636);
nor U7832 (N_7832,N_6815,N_6637);
nor U7833 (N_7833,N_6826,N_6187);
nor U7834 (N_7834,N_6757,N_6704);
and U7835 (N_7835,N_6847,N_6186);
or U7836 (N_7836,N_6793,N_6019);
and U7837 (N_7837,N_6974,N_6516);
nor U7838 (N_7838,N_6458,N_6215);
nand U7839 (N_7839,N_6444,N_6200);
xor U7840 (N_7840,N_6634,N_6182);
nand U7841 (N_7841,N_6440,N_6040);
and U7842 (N_7842,N_6262,N_6081);
nand U7843 (N_7843,N_6890,N_6038);
or U7844 (N_7844,N_6162,N_6484);
xnor U7845 (N_7845,N_6669,N_6136);
nor U7846 (N_7846,N_6370,N_6599);
xnor U7847 (N_7847,N_6507,N_6484);
xnor U7848 (N_7848,N_6842,N_6150);
or U7849 (N_7849,N_6766,N_6924);
and U7850 (N_7850,N_6064,N_6078);
nand U7851 (N_7851,N_6485,N_6401);
xor U7852 (N_7852,N_6293,N_6285);
nor U7853 (N_7853,N_6713,N_6017);
nand U7854 (N_7854,N_6818,N_6270);
nand U7855 (N_7855,N_6387,N_6594);
and U7856 (N_7856,N_6598,N_6107);
and U7857 (N_7857,N_6501,N_6695);
and U7858 (N_7858,N_6258,N_6725);
xnor U7859 (N_7859,N_6001,N_6960);
and U7860 (N_7860,N_6895,N_6021);
xor U7861 (N_7861,N_6205,N_6492);
nand U7862 (N_7862,N_6948,N_6038);
and U7863 (N_7863,N_6225,N_6551);
nor U7864 (N_7864,N_6232,N_6479);
nand U7865 (N_7865,N_6005,N_6806);
nand U7866 (N_7866,N_6406,N_6560);
nand U7867 (N_7867,N_6262,N_6863);
nand U7868 (N_7868,N_6735,N_6914);
xnor U7869 (N_7869,N_6082,N_6525);
or U7870 (N_7870,N_6413,N_6694);
nand U7871 (N_7871,N_6002,N_6986);
nand U7872 (N_7872,N_6015,N_6900);
xnor U7873 (N_7873,N_6634,N_6821);
or U7874 (N_7874,N_6531,N_6850);
nor U7875 (N_7875,N_6477,N_6356);
or U7876 (N_7876,N_6462,N_6523);
and U7877 (N_7877,N_6955,N_6632);
xor U7878 (N_7878,N_6810,N_6231);
or U7879 (N_7879,N_6927,N_6000);
nand U7880 (N_7880,N_6065,N_6611);
nand U7881 (N_7881,N_6401,N_6313);
nor U7882 (N_7882,N_6850,N_6575);
nor U7883 (N_7883,N_6342,N_6639);
and U7884 (N_7884,N_6943,N_6539);
nor U7885 (N_7885,N_6798,N_6781);
and U7886 (N_7886,N_6843,N_6428);
xnor U7887 (N_7887,N_6050,N_6553);
or U7888 (N_7888,N_6263,N_6693);
nand U7889 (N_7889,N_6379,N_6632);
and U7890 (N_7890,N_6879,N_6934);
and U7891 (N_7891,N_6733,N_6422);
nand U7892 (N_7892,N_6938,N_6436);
xor U7893 (N_7893,N_6014,N_6903);
and U7894 (N_7894,N_6475,N_6490);
or U7895 (N_7895,N_6621,N_6180);
and U7896 (N_7896,N_6368,N_6073);
or U7897 (N_7897,N_6332,N_6749);
xnor U7898 (N_7898,N_6383,N_6656);
nand U7899 (N_7899,N_6455,N_6786);
nand U7900 (N_7900,N_6686,N_6566);
or U7901 (N_7901,N_6793,N_6072);
nand U7902 (N_7902,N_6586,N_6320);
nand U7903 (N_7903,N_6890,N_6962);
xor U7904 (N_7904,N_6355,N_6832);
xnor U7905 (N_7905,N_6476,N_6988);
nor U7906 (N_7906,N_6557,N_6624);
xor U7907 (N_7907,N_6163,N_6340);
nand U7908 (N_7908,N_6340,N_6339);
or U7909 (N_7909,N_6688,N_6860);
nor U7910 (N_7910,N_6658,N_6832);
nor U7911 (N_7911,N_6997,N_6832);
and U7912 (N_7912,N_6145,N_6186);
or U7913 (N_7913,N_6877,N_6764);
xor U7914 (N_7914,N_6062,N_6485);
nand U7915 (N_7915,N_6716,N_6092);
or U7916 (N_7916,N_6554,N_6141);
xnor U7917 (N_7917,N_6051,N_6582);
nand U7918 (N_7918,N_6338,N_6400);
or U7919 (N_7919,N_6495,N_6847);
and U7920 (N_7920,N_6240,N_6631);
and U7921 (N_7921,N_6036,N_6721);
nand U7922 (N_7922,N_6479,N_6325);
or U7923 (N_7923,N_6693,N_6754);
and U7924 (N_7924,N_6691,N_6656);
nor U7925 (N_7925,N_6687,N_6353);
and U7926 (N_7926,N_6668,N_6264);
or U7927 (N_7927,N_6184,N_6108);
nor U7928 (N_7928,N_6278,N_6735);
and U7929 (N_7929,N_6499,N_6696);
nand U7930 (N_7930,N_6939,N_6623);
or U7931 (N_7931,N_6204,N_6666);
and U7932 (N_7932,N_6919,N_6556);
and U7933 (N_7933,N_6754,N_6096);
or U7934 (N_7934,N_6617,N_6728);
and U7935 (N_7935,N_6038,N_6490);
nor U7936 (N_7936,N_6222,N_6331);
xor U7937 (N_7937,N_6880,N_6672);
nor U7938 (N_7938,N_6690,N_6672);
and U7939 (N_7939,N_6852,N_6979);
nor U7940 (N_7940,N_6456,N_6689);
nand U7941 (N_7941,N_6692,N_6603);
or U7942 (N_7942,N_6000,N_6421);
nor U7943 (N_7943,N_6017,N_6334);
nand U7944 (N_7944,N_6472,N_6775);
nand U7945 (N_7945,N_6285,N_6698);
or U7946 (N_7946,N_6082,N_6278);
nand U7947 (N_7947,N_6597,N_6206);
nand U7948 (N_7948,N_6412,N_6451);
and U7949 (N_7949,N_6166,N_6318);
and U7950 (N_7950,N_6473,N_6545);
xor U7951 (N_7951,N_6605,N_6658);
and U7952 (N_7952,N_6672,N_6553);
xnor U7953 (N_7953,N_6208,N_6109);
nand U7954 (N_7954,N_6508,N_6878);
nor U7955 (N_7955,N_6503,N_6474);
xnor U7956 (N_7956,N_6299,N_6118);
xor U7957 (N_7957,N_6933,N_6524);
and U7958 (N_7958,N_6834,N_6174);
and U7959 (N_7959,N_6138,N_6092);
xor U7960 (N_7960,N_6466,N_6665);
nor U7961 (N_7961,N_6517,N_6622);
nand U7962 (N_7962,N_6700,N_6446);
and U7963 (N_7963,N_6363,N_6422);
xor U7964 (N_7964,N_6115,N_6387);
nor U7965 (N_7965,N_6831,N_6454);
nand U7966 (N_7966,N_6124,N_6615);
nor U7967 (N_7967,N_6345,N_6754);
nor U7968 (N_7968,N_6016,N_6155);
nand U7969 (N_7969,N_6784,N_6971);
or U7970 (N_7970,N_6569,N_6820);
nor U7971 (N_7971,N_6904,N_6763);
nor U7972 (N_7972,N_6702,N_6199);
and U7973 (N_7973,N_6629,N_6110);
nor U7974 (N_7974,N_6439,N_6680);
xnor U7975 (N_7975,N_6904,N_6643);
nor U7976 (N_7976,N_6164,N_6619);
nor U7977 (N_7977,N_6772,N_6624);
and U7978 (N_7978,N_6284,N_6890);
xnor U7979 (N_7979,N_6023,N_6266);
xor U7980 (N_7980,N_6427,N_6023);
nand U7981 (N_7981,N_6757,N_6606);
and U7982 (N_7982,N_6270,N_6951);
nand U7983 (N_7983,N_6889,N_6119);
nor U7984 (N_7984,N_6191,N_6959);
and U7985 (N_7985,N_6771,N_6869);
nand U7986 (N_7986,N_6310,N_6108);
nand U7987 (N_7987,N_6088,N_6772);
and U7988 (N_7988,N_6497,N_6483);
or U7989 (N_7989,N_6554,N_6403);
nor U7990 (N_7990,N_6625,N_6647);
and U7991 (N_7991,N_6672,N_6812);
and U7992 (N_7992,N_6355,N_6201);
nand U7993 (N_7993,N_6318,N_6528);
nand U7994 (N_7994,N_6566,N_6270);
nand U7995 (N_7995,N_6507,N_6573);
xnor U7996 (N_7996,N_6221,N_6528);
nor U7997 (N_7997,N_6414,N_6368);
nor U7998 (N_7998,N_6799,N_6673);
nand U7999 (N_7999,N_6780,N_6589);
or U8000 (N_8000,N_7213,N_7767);
or U8001 (N_8001,N_7676,N_7906);
or U8002 (N_8002,N_7430,N_7204);
and U8003 (N_8003,N_7777,N_7363);
xnor U8004 (N_8004,N_7976,N_7815);
and U8005 (N_8005,N_7952,N_7257);
nor U8006 (N_8006,N_7969,N_7281);
or U8007 (N_8007,N_7594,N_7998);
xnor U8008 (N_8008,N_7378,N_7251);
and U8009 (N_8009,N_7657,N_7694);
nor U8010 (N_8010,N_7505,N_7894);
xor U8011 (N_8011,N_7396,N_7724);
and U8012 (N_8012,N_7375,N_7580);
nor U8013 (N_8013,N_7726,N_7042);
or U8014 (N_8014,N_7974,N_7552);
or U8015 (N_8015,N_7265,N_7899);
nand U8016 (N_8016,N_7658,N_7308);
nor U8017 (N_8017,N_7855,N_7092);
nand U8018 (N_8018,N_7354,N_7255);
or U8019 (N_8019,N_7020,N_7350);
nand U8020 (N_8020,N_7644,N_7884);
or U8021 (N_8021,N_7837,N_7423);
and U8022 (N_8022,N_7557,N_7065);
and U8023 (N_8023,N_7599,N_7037);
nor U8024 (N_8024,N_7043,N_7618);
or U8025 (N_8025,N_7493,N_7157);
nor U8026 (N_8026,N_7611,N_7848);
and U8027 (N_8027,N_7847,N_7639);
or U8028 (N_8028,N_7756,N_7929);
and U8029 (N_8029,N_7287,N_7347);
nand U8030 (N_8030,N_7061,N_7192);
or U8031 (N_8031,N_7302,N_7652);
nor U8032 (N_8032,N_7366,N_7584);
or U8033 (N_8033,N_7443,N_7259);
or U8034 (N_8034,N_7547,N_7314);
and U8035 (N_8035,N_7900,N_7253);
xnor U8036 (N_8036,N_7151,N_7235);
and U8037 (N_8037,N_7395,N_7181);
nor U8038 (N_8038,N_7244,N_7967);
nor U8039 (N_8039,N_7706,N_7663);
nor U8040 (N_8040,N_7785,N_7982);
or U8041 (N_8041,N_7217,N_7172);
and U8042 (N_8042,N_7937,N_7691);
or U8043 (N_8043,N_7093,N_7765);
xor U8044 (N_8044,N_7530,N_7579);
nand U8045 (N_8045,N_7955,N_7523);
and U8046 (N_8046,N_7797,N_7809);
or U8047 (N_8047,N_7304,N_7510);
nand U8048 (N_8048,N_7773,N_7185);
nand U8049 (N_8049,N_7176,N_7054);
and U8050 (N_8050,N_7410,N_7620);
nand U8051 (N_8051,N_7112,N_7002);
and U8052 (N_8052,N_7492,N_7124);
and U8053 (N_8053,N_7254,N_7017);
nand U8054 (N_8054,N_7509,N_7223);
or U8055 (N_8055,N_7716,N_7108);
nor U8056 (N_8056,N_7193,N_7865);
or U8057 (N_8057,N_7048,N_7438);
nand U8058 (N_8058,N_7041,N_7384);
or U8059 (N_8059,N_7299,N_7078);
nand U8060 (N_8060,N_7806,N_7852);
nor U8061 (N_8061,N_7480,N_7717);
nand U8062 (N_8062,N_7524,N_7592);
or U8063 (N_8063,N_7913,N_7886);
or U8064 (N_8064,N_7590,N_7989);
or U8065 (N_8065,N_7935,N_7850);
nand U8066 (N_8066,N_7619,N_7686);
and U8067 (N_8067,N_7024,N_7623);
nand U8068 (N_8068,N_7285,N_7490);
nor U8069 (N_8069,N_7883,N_7573);
and U8070 (N_8070,N_7332,N_7392);
xnor U8071 (N_8071,N_7648,N_7402);
nor U8072 (N_8072,N_7985,N_7868);
or U8073 (N_8073,N_7803,N_7635);
nand U8074 (N_8074,N_7858,N_7113);
xnor U8075 (N_8075,N_7519,N_7687);
nor U8076 (N_8076,N_7000,N_7117);
xnor U8077 (N_8077,N_7545,N_7533);
nor U8078 (N_8078,N_7636,N_7907);
and U8079 (N_8079,N_7928,N_7925);
nor U8080 (N_8080,N_7548,N_7664);
nand U8081 (N_8081,N_7436,N_7058);
or U8082 (N_8082,N_7578,N_7760);
or U8083 (N_8083,N_7381,N_7497);
nor U8084 (N_8084,N_7066,N_7056);
and U8085 (N_8085,N_7129,N_7435);
and U8086 (N_8086,N_7359,N_7529);
and U8087 (N_8087,N_7645,N_7753);
or U8088 (N_8088,N_7307,N_7301);
nor U8089 (N_8089,N_7946,N_7555);
nor U8090 (N_8090,N_7322,N_7534);
and U8091 (N_8091,N_7703,N_7214);
nand U8092 (N_8092,N_7241,N_7426);
nor U8093 (N_8093,N_7881,N_7541);
xor U8094 (N_8094,N_7387,N_7627);
nor U8095 (N_8095,N_7477,N_7422);
xor U8096 (N_8096,N_7641,N_7382);
xor U8097 (N_8097,N_7938,N_7038);
xnor U8098 (N_8098,N_7771,N_7064);
nand U8099 (N_8099,N_7310,N_7236);
nand U8100 (N_8100,N_7574,N_7692);
and U8101 (N_8101,N_7197,N_7072);
nor U8102 (N_8102,N_7804,N_7001);
and U8103 (N_8103,N_7588,N_7252);
xor U8104 (N_8104,N_7950,N_7247);
xnor U8105 (N_8105,N_7857,N_7734);
nand U8106 (N_8106,N_7059,N_7032);
and U8107 (N_8107,N_7186,N_7010);
nand U8108 (N_8108,N_7246,N_7601);
and U8109 (N_8109,N_7418,N_7680);
nand U8110 (N_8110,N_7282,N_7099);
and U8111 (N_8111,N_7256,N_7147);
or U8112 (N_8112,N_7461,N_7604);
nor U8113 (N_8113,N_7261,N_7788);
nor U8114 (N_8114,N_7828,N_7669);
nand U8115 (N_8115,N_7207,N_7709);
nand U8116 (N_8116,N_7927,N_7429);
and U8117 (N_8117,N_7637,N_7999);
nor U8118 (N_8118,N_7923,N_7475);
nor U8119 (N_8119,N_7810,N_7587);
and U8120 (N_8120,N_7311,N_7144);
nor U8121 (N_8121,N_7075,N_7374);
nor U8122 (N_8122,N_7120,N_7388);
and U8123 (N_8123,N_7714,N_7672);
nand U8124 (N_8124,N_7393,N_7919);
or U8125 (N_8125,N_7980,N_7459);
nor U8126 (N_8126,N_7630,N_7634);
nor U8127 (N_8127,N_7211,N_7462);
and U8128 (N_8128,N_7216,N_7478);
nand U8129 (N_8129,N_7448,N_7715);
nor U8130 (N_8130,N_7428,N_7812);
nand U8131 (N_8131,N_7445,N_7051);
xnor U8132 (N_8132,N_7508,N_7165);
xnor U8133 (N_8133,N_7011,N_7902);
or U8134 (N_8134,N_7646,N_7289);
or U8135 (N_8135,N_7476,N_7668);
and U8136 (N_8136,N_7559,N_7158);
nand U8137 (N_8137,N_7409,N_7647);
or U8138 (N_8138,N_7349,N_7153);
nor U8139 (N_8139,N_7598,N_7926);
nor U8140 (N_8140,N_7231,N_7954);
xor U8141 (N_8141,N_7738,N_7102);
nand U8142 (N_8142,N_7199,N_7903);
or U8143 (N_8143,N_7135,N_7162);
nor U8144 (N_8144,N_7786,N_7411);
xnor U8145 (N_8145,N_7468,N_7007);
or U8146 (N_8146,N_7737,N_7205);
nor U8147 (N_8147,N_7016,N_7425);
xor U8148 (N_8148,N_7667,N_7170);
nand U8149 (N_8149,N_7684,N_7596);
nor U8150 (N_8150,N_7296,N_7187);
and U8151 (N_8151,N_7867,N_7401);
nor U8152 (N_8152,N_7990,N_7670);
or U8153 (N_8153,N_7626,N_7142);
and U8154 (N_8154,N_7368,N_7437);
nor U8155 (N_8155,N_7965,N_7742);
nor U8156 (N_8156,N_7780,N_7964);
and U8157 (N_8157,N_7528,N_7538);
nor U8158 (N_8158,N_7696,N_7268);
and U8159 (N_8159,N_7267,N_7063);
nor U8160 (N_8160,N_7233,N_7270);
nand U8161 (N_8161,N_7609,N_7139);
nor U8162 (N_8162,N_7708,N_7227);
xnor U8163 (N_8163,N_7355,N_7602);
and U8164 (N_8164,N_7249,N_7732);
nor U8165 (N_8165,N_7278,N_7431);
or U8166 (N_8166,N_7793,N_7330);
and U8167 (N_8167,N_7128,N_7957);
nor U8168 (N_8168,N_7918,N_7665);
nor U8169 (N_8169,N_7491,N_7939);
and U8170 (N_8170,N_7380,N_7503);
nand U8171 (N_8171,N_7705,N_7420);
and U8172 (N_8172,N_7184,N_7895);
nand U8173 (N_8173,N_7313,N_7791);
and U8174 (N_8174,N_7277,N_7309);
xnor U8175 (N_8175,N_7878,N_7546);
nand U8176 (N_8176,N_7603,N_7838);
nor U8177 (N_8177,N_7383,N_7678);
nand U8178 (N_8178,N_7076,N_7130);
nor U8179 (N_8179,N_7829,N_7198);
and U8180 (N_8180,N_7103,N_7394);
or U8181 (N_8181,N_7452,N_7605);
nand U8182 (N_8182,N_7718,N_7994);
xnor U8183 (N_8183,N_7606,N_7098);
nor U8184 (N_8184,N_7360,N_7479);
and U8185 (N_8185,N_7224,N_7434);
and U8186 (N_8186,N_7303,N_7004);
or U8187 (N_8187,N_7370,N_7173);
and U8188 (N_8188,N_7553,N_7518);
or U8189 (N_8189,N_7498,N_7229);
nor U8190 (N_8190,N_7874,N_7014);
nand U8191 (N_8191,N_7975,N_7472);
nor U8192 (N_8192,N_7700,N_7835);
or U8193 (N_8193,N_7564,N_7915);
xnor U8194 (N_8194,N_7450,N_7013);
nor U8195 (N_8195,N_7306,N_7962);
xor U8196 (N_8196,N_7221,N_7416);
or U8197 (N_8197,N_7209,N_7496);
nand U8198 (N_8198,N_7447,N_7789);
or U8199 (N_8199,N_7225,N_7543);
xnor U8200 (N_8200,N_7695,N_7140);
xnor U8201 (N_8201,N_7909,N_7084);
or U8202 (N_8202,N_7683,N_7454);
or U8203 (N_8203,N_7615,N_7196);
or U8204 (N_8204,N_7854,N_7822);
and U8205 (N_8205,N_7266,N_7551);
and U8206 (N_8206,N_7271,N_7910);
xnor U8207 (N_8207,N_7203,N_7086);
and U8208 (N_8208,N_7693,N_7662);
nand U8209 (N_8209,N_7487,N_7179);
xnor U8210 (N_8210,N_7081,N_7782);
nand U8211 (N_8211,N_7045,N_7134);
nand U8212 (N_8212,N_7333,N_7770);
or U8213 (N_8213,N_7862,N_7525);
or U8214 (N_8214,N_7284,N_7844);
nand U8215 (N_8215,N_7677,N_7190);
nor U8216 (N_8216,N_7743,N_7331);
or U8217 (N_8217,N_7466,N_7337);
nor U8218 (N_8218,N_7115,N_7515);
nor U8219 (N_8219,N_7589,N_7792);
nor U8220 (N_8220,N_7039,N_7653);
and U8221 (N_8221,N_7276,N_7567);
nand U8222 (N_8222,N_7164,N_7730);
nor U8223 (N_8223,N_7751,N_7890);
and U8224 (N_8224,N_7062,N_7960);
or U8225 (N_8225,N_7210,N_7202);
xnor U8226 (N_8226,N_7326,N_7335);
or U8227 (N_8227,N_7568,N_7397);
or U8228 (N_8228,N_7018,N_7876);
and U8229 (N_8229,N_7825,N_7094);
nand U8230 (N_8230,N_7150,N_7549);
nor U8231 (N_8231,N_7631,N_7712);
or U8232 (N_8232,N_7071,N_7433);
nand U8233 (N_8233,N_7177,N_7872);
or U8234 (N_8234,N_7986,N_7080);
and U8235 (N_8235,N_7860,N_7775);
nor U8236 (N_8236,N_7853,N_7188);
nand U8237 (N_8237,N_7898,N_7735);
nand U8238 (N_8238,N_7167,N_7485);
or U8239 (N_8239,N_7174,N_7940);
nor U8240 (N_8240,N_7660,N_7339);
nor U8241 (N_8241,N_7463,N_7704);
or U8242 (N_8242,N_7869,N_7215);
nor U8243 (N_8243,N_7100,N_7951);
nor U8244 (N_8244,N_7352,N_7357);
nand U8245 (N_8245,N_7467,N_7095);
xor U8246 (N_8246,N_7364,N_7377);
nand U8247 (N_8247,N_7319,N_7323);
xor U8248 (N_8248,N_7572,N_7522);
and U8249 (N_8249,N_7550,N_7591);
and U8250 (N_8250,N_7930,N_7741);
nand U8251 (N_8251,N_7707,N_7995);
nor U8252 (N_8252,N_7554,N_7273);
nand U8253 (N_8253,N_7556,N_7840);
nand U8254 (N_8254,N_7212,N_7312);
and U8255 (N_8255,N_7324,N_7517);
or U8256 (N_8256,N_7819,N_7661);
and U8257 (N_8257,N_7798,N_7507);
nor U8258 (N_8258,N_7628,N_7759);
nand U8259 (N_8259,N_7947,N_7656);
xnor U8260 (N_8260,N_7453,N_7739);
nor U8261 (N_8261,N_7168,N_7346);
or U8262 (N_8262,N_7943,N_7784);
or U8263 (N_8263,N_7090,N_7750);
or U8264 (N_8264,N_7219,N_7633);
nand U8265 (N_8265,N_7026,N_7079);
xor U8266 (N_8266,N_7945,N_7908);
or U8267 (N_8267,N_7222,N_7801);
or U8268 (N_8268,N_7713,N_7889);
and U8269 (N_8269,N_7571,N_7089);
and U8270 (N_8270,N_7022,N_7096);
nor U8271 (N_8271,N_7725,N_7027);
xnor U8272 (N_8272,N_7916,N_7827);
and U8273 (N_8273,N_7892,N_7414);
xnor U8274 (N_8274,N_7893,N_7563);
nand U8275 (N_8275,N_7195,N_7575);
and U8276 (N_8276,N_7012,N_7710);
nor U8277 (N_8277,N_7651,N_7036);
xnor U8278 (N_8278,N_7851,N_7116);
and U8279 (N_8279,N_7484,N_7031);
nor U8280 (N_8280,N_7841,N_7914);
nand U8281 (N_8281,N_7028,N_7228);
and U8282 (N_8282,N_7649,N_7444);
or U8283 (N_8283,N_7582,N_7040);
or U8284 (N_8284,N_7060,N_7156);
or U8285 (N_8285,N_7379,N_7009);
and U8286 (N_8286,N_7754,N_7871);
and U8287 (N_8287,N_7432,N_7755);
xor U8288 (N_8288,N_7640,N_7617);
or U8289 (N_8289,N_7681,N_7023);
or U8290 (N_8290,N_7632,N_7757);
or U8291 (N_8291,N_7736,N_7486);
nand U8292 (N_8292,N_7136,N_7149);
nand U8293 (N_8293,N_7966,N_7465);
and U8294 (N_8294,N_7279,N_7146);
or U8295 (N_8295,N_7520,N_7991);
or U8296 (N_8296,N_7794,N_7417);
and U8297 (N_8297,N_7440,N_7327);
nor U8298 (N_8298,N_7406,N_7817);
or U8299 (N_8299,N_7183,N_7237);
xnor U8300 (N_8300,N_7931,N_7118);
or U8301 (N_8301,N_7544,N_7805);
and U8302 (N_8302,N_7180,N_7131);
or U8303 (N_8303,N_7861,N_7234);
nand U8304 (N_8304,N_7141,N_7050);
or U8305 (N_8305,N_7154,N_7842);
and U8306 (N_8306,N_7344,N_7539);
nor U8307 (N_8307,N_7272,N_7200);
and U8308 (N_8308,N_7220,N_7351);
nor U8309 (N_8309,N_7949,N_7356);
and U8310 (N_8310,N_7015,N_7566);
nand U8311 (N_8311,N_7082,N_7160);
or U8312 (N_8312,N_7125,N_7911);
nand U8313 (N_8313,N_7897,N_7362);
nand U8314 (N_8314,N_7796,N_7029);
nor U8315 (N_8315,N_7451,N_7389);
and U8316 (N_8316,N_7823,N_7845);
nand U8317 (N_8317,N_7159,N_7722);
nor U8318 (N_8318,N_7248,N_7148);
or U8319 (N_8319,N_7442,N_7540);
or U8320 (N_8320,N_7856,N_7821);
or U8321 (N_8321,N_7948,N_7882);
nand U8322 (N_8322,N_7600,N_7673);
nand U8323 (N_8323,N_7329,N_7521);
and U8324 (N_8324,N_7761,N_7781);
or U8325 (N_8325,N_7240,N_7297);
nor U8326 (N_8326,N_7537,N_7025);
and U8327 (N_8327,N_7610,N_7972);
or U8328 (N_8328,N_7504,N_7934);
and U8329 (N_8329,N_7057,N_7390);
nor U8330 (N_8330,N_7182,N_7629);
xnor U8331 (N_8331,N_7321,N_7888);
or U8332 (N_8332,N_7483,N_7752);
xnor U8333 (N_8333,N_7859,N_7398);
or U8334 (N_8334,N_7833,N_7325);
xor U8335 (N_8335,N_7532,N_7373);
and U8336 (N_8336,N_7201,N_7818);
or U8337 (N_8337,N_7073,N_7811);
and U8338 (N_8338,N_7728,N_7824);
and U8339 (N_8339,N_7361,N_7400);
xor U8340 (N_8340,N_7997,N_7005);
or U8341 (N_8341,N_7993,N_7415);
xnor U8342 (N_8342,N_7904,N_7593);
or U8343 (N_8343,N_7105,N_7449);
nand U8344 (N_8344,N_7772,N_7191);
or U8345 (N_8345,N_7258,N_7682);
nand U8346 (N_8346,N_7034,N_7795);
nand U8347 (N_8347,N_7880,N_7419);
and U8348 (N_8348,N_7455,N_7345);
or U8349 (N_8349,N_7961,N_7624);
nand U8350 (N_8350,N_7123,N_7787);
and U8351 (N_8351,N_7679,N_7298);
nand U8352 (N_8352,N_7053,N_7376);
and U8353 (N_8353,N_7959,N_7614);
nand U8354 (N_8354,N_7671,N_7456);
nand U8355 (N_8355,N_7175,N_7953);
xnor U8356 (N_8356,N_7132,N_7161);
nor U8357 (N_8357,N_7920,N_7341);
and U8358 (N_8358,N_7896,N_7643);
and U8359 (N_8359,N_7399,N_7807);
nand U8360 (N_8360,N_7612,N_7260);
nand U8361 (N_8361,N_7119,N_7625);
and U8362 (N_8362,N_7570,N_7763);
or U8363 (N_8363,N_7674,N_7166);
and U8364 (N_8364,N_7501,N_7597);
nor U8365 (N_8365,N_7405,N_7250);
nor U8366 (N_8366,N_7879,N_7049);
nand U8367 (N_8367,N_7666,N_7870);
nor U8368 (N_8368,N_7992,N_7699);
or U8369 (N_8369,N_7638,N_7077);
nor U8370 (N_8370,N_7971,N_7471);
or U8371 (N_8371,N_7981,N_7689);
and U8372 (N_8372,N_7866,N_7813);
or U8373 (N_8373,N_7274,N_7746);
and U8374 (N_8374,N_7328,N_7145);
and U8375 (N_8375,N_7372,N_7558);
xnor U8376 (N_8376,N_7107,N_7748);
nor U8377 (N_8377,N_7996,N_7963);
nand U8378 (N_8378,N_7283,N_7178);
and U8379 (N_8379,N_7055,N_7917);
nor U8380 (N_8380,N_7239,N_7412);
and U8381 (N_8381,N_7316,N_7122);
or U8382 (N_8382,N_7243,N_7973);
nand U8383 (N_8383,N_7542,N_7275);
or U8384 (N_8384,N_7369,N_7106);
or U8385 (N_8385,N_7527,N_7336);
nor U8386 (N_8386,N_7968,N_7046);
and U8387 (N_8387,N_7458,N_7232);
and U8388 (N_8388,N_7690,N_7218);
nor U8389 (N_8389,N_7836,N_7800);
and U8390 (N_8390,N_7280,N_7408);
and U8391 (N_8391,N_7887,N_7155);
nor U8392 (N_8392,N_7021,N_7747);
nand U8393 (N_8393,N_7052,N_7121);
or U8394 (N_8394,N_7044,N_7758);
nand U8395 (N_8395,N_7473,N_7740);
and U8396 (N_8396,N_7901,N_7585);
xor U8397 (N_8397,N_7245,N_7942);
nor U8398 (N_8398,N_7292,N_7729);
and U8399 (N_8399,N_7169,N_7814);
and U8400 (N_8400,N_7839,N_7526);
nand U8401 (N_8401,N_7922,N_7936);
or U8402 (N_8402,N_7097,N_7494);
nand U8403 (N_8403,N_7305,N_7269);
nor U8404 (N_8404,N_7650,N_7834);
nand U8405 (N_8405,N_7688,N_7502);
or U8406 (N_8406,N_7262,N_7830);
nor U8407 (N_8407,N_7424,N_7749);
or U8408 (N_8408,N_7933,N_7385);
nor U8409 (N_8409,N_7970,N_7745);
nor U8410 (N_8410,N_7189,N_7413);
nand U8411 (N_8411,N_7286,N_7295);
and U8412 (N_8412,N_7242,N_7315);
nand U8413 (N_8413,N_7560,N_7941);
nand U8414 (N_8414,N_7642,N_7733);
nor U8415 (N_8415,N_7912,N_7358);
and U8416 (N_8416,N_7873,N_7863);
nand U8417 (N_8417,N_7565,N_7404);
nand U8418 (N_8418,N_7654,N_7264);
nor U8419 (N_8419,N_7230,N_7109);
nor U8420 (N_8420,N_7849,N_7616);
nor U8421 (N_8421,N_7226,N_7586);
and U8422 (N_8422,N_7831,N_7343);
and U8423 (N_8423,N_7386,N_7790);
nand U8424 (N_8424,N_7104,N_7003);
nand U8425 (N_8425,N_7047,N_7291);
or U8426 (N_8426,N_7769,N_7832);
nor U8427 (N_8427,N_7489,N_7067);
or U8428 (N_8428,N_7138,N_7338);
nor U8429 (N_8429,N_7768,N_7562);
and U8430 (N_8430,N_7514,N_7511);
and U8431 (N_8431,N_7403,N_7595);
nand U8432 (N_8432,N_7019,N_7799);
or U8433 (N_8433,N_7727,N_7816);
nand U8434 (N_8434,N_7983,N_7208);
nand U8435 (N_8435,N_7607,N_7290);
and U8436 (N_8436,N_7008,N_7720);
xor U8437 (N_8437,N_7126,N_7101);
xnor U8438 (N_8438,N_7988,N_7334);
nor U8439 (N_8439,N_7342,N_7320);
nor U8440 (N_8440,N_7068,N_7697);
or U8441 (N_8441,N_7365,N_7137);
nor U8442 (N_8442,N_7621,N_7846);
nor U8443 (N_8443,N_7685,N_7074);
and U8444 (N_8444,N_7583,N_7576);
nand U8445 (N_8445,N_7163,N_7977);
nor U8446 (N_8446,N_7110,N_7348);
nand U8447 (N_8447,N_7085,N_7495);
nand U8448 (N_8448,N_7764,N_7877);
nand U8449 (N_8449,N_7317,N_7469);
nand U8450 (N_8450,N_7608,N_7723);
or U8451 (N_8451,N_7006,N_7783);
and U8452 (N_8452,N_7655,N_7512);
nor U8453 (N_8453,N_7294,N_7774);
nor U8454 (N_8454,N_7675,N_7875);
nor U8455 (N_8455,N_7924,N_7087);
and U8456 (N_8456,N_7561,N_7516);
nor U8457 (N_8457,N_7905,N_7802);
nand U8458 (N_8458,N_7318,N_7391);
xor U8459 (N_8459,N_7531,N_7488);
nand U8460 (N_8460,N_7263,N_7978);
nand U8461 (N_8461,N_7932,N_7439);
xor U8462 (N_8462,N_7921,N_7194);
xnor U8463 (N_8463,N_7958,N_7464);
xnor U8464 (N_8464,N_7152,N_7088);
and U8465 (N_8465,N_7171,N_7701);
and U8466 (N_8466,N_7127,N_7698);
and U8467 (N_8467,N_7744,N_7460);
nand U8468 (N_8468,N_7030,N_7033);
nor U8469 (N_8469,N_7731,N_7826);
and U8470 (N_8470,N_7427,N_7659);
or U8471 (N_8471,N_7470,N_7288);
nor U8472 (N_8472,N_7778,N_7808);
or U8473 (N_8473,N_7293,N_7864);
or U8474 (N_8474,N_7481,N_7820);
and U8475 (N_8475,N_7956,N_7613);
and U8476 (N_8476,N_7577,N_7371);
or U8477 (N_8477,N_7111,N_7206);
and U8478 (N_8478,N_7407,N_7441);
nor U8479 (N_8479,N_7482,N_7083);
nand U8480 (N_8480,N_7353,N_7987);
and U8481 (N_8481,N_7984,N_7300);
and U8482 (N_8482,N_7979,N_7513);
nor U8483 (N_8483,N_7885,N_7776);
xnor U8484 (N_8484,N_7367,N_7114);
nand U8485 (N_8485,N_7944,N_7702);
or U8486 (N_8486,N_7719,N_7506);
nand U8487 (N_8487,N_7891,N_7779);
or U8488 (N_8488,N_7133,N_7143);
and U8489 (N_8489,N_7474,N_7569);
nand U8490 (N_8490,N_7581,N_7843);
nor U8491 (N_8491,N_7070,N_7091);
xor U8492 (N_8492,N_7535,N_7622);
nand U8493 (N_8493,N_7238,N_7762);
nor U8494 (N_8494,N_7457,N_7340);
or U8495 (N_8495,N_7766,N_7536);
and U8496 (N_8496,N_7500,N_7069);
nand U8497 (N_8497,N_7446,N_7421);
and U8498 (N_8498,N_7035,N_7711);
nor U8499 (N_8499,N_7499,N_7721);
or U8500 (N_8500,N_7323,N_7113);
or U8501 (N_8501,N_7332,N_7383);
nor U8502 (N_8502,N_7030,N_7706);
or U8503 (N_8503,N_7691,N_7936);
nand U8504 (N_8504,N_7727,N_7376);
xnor U8505 (N_8505,N_7580,N_7160);
nand U8506 (N_8506,N_7926,N_7769);
or U8507 (N_8507,N_7575,N_7646);
nor U8508 (N_8508,N_7075,N_7223);
nor U8509 (N_8509,N_7510,N_7753);
nor U8510 (N_8510,N_7098,N_7431);
nand U8511 (N_8511,N_7374,N_7437);
nand U8512 (N_8512,N_7584,N_7065);
nor U8513 (N_8513,N_7938,N_7286);
or U8514 (N_8514,N_7376,N_7849);
and U8515 (N_8515,N_7902,N_7161);
nand U8516 (N_8516,N_7404,N_7507);
and U8517 (N_8517,N_7615,N_7679);
xnor U8518 (N_8518,N_7429,N_7096);
and U8519 (N_8519,N_7750,N_7323);
xor U8520 (N_8520,N_7085,N_7814);
xor U8521 (N_8521,N_7013,N_7205);
or U8522 (N_8522,N_7986,N_7051);
xnor U8523 (N_8523,N_7096,N_7510);
xor U8524 (N_8524,N_7983,N_7667);
and U8525 (N_8525,N_7255,N_7149);
and U8526 (N_8526,N_7390,N_7586);
nand U8527 (N_8527,N_7007,N_7581);
nor U8528 (N_8528,N_7577,N_7879);
nand U8529 (N_8529,N_7212,N_7705);
nor U8530 (N_8530,N_7786,N_7222);
nand U8531 (N_8531,N_7154,N_7826);
nand U8532 (N_8532,N_7692,N_7965);
nor U8533 (N_8533,N_7254,N_7760);
nor U8534 (N_8534,N_7169,N_7978);
nor U8535 (N_8535,N_7541,N_7096);
or U8536 (N_8536,N_7555,N_7746);
and U8537 (N_8537,N_7342,N_7995);
or U8538 (N_8538,N_7321,N_7624);
nand U8539 (N_8539,N_7816,N_7414);
nor U8540 (N_8540,N_7497,N_7478);
nor U8541 (N_8541,N_7058,N_7554);
nand U8542 (N_8542,N_7698,N_7123);
nor U8543 (N_8543,N_7921,N_7941);
or U8544 (N_8544,N_7531,N_7061);
and U8545 (N_8545,N_7235,N_7799);
nor U8546 (N_8546,N_7419,N_7631);
nor U8547 (N_8547,N_7608,N_7694);
xnor U8548 (N_8548,N_7084,N_7108);
nor U8549 (N_8549,N_7311,N_7472);
nor U8550 (N_8550,N_7724,N_7578);
nor U8551 (N_8551,N_7244,N_7395);
nor U8552 (N_8552,N_7100,N_7794);
or U8553 (N_8553,N_7064,N_7265);
or U8554 (N_8554,N_7435,N_7982);
and U8555 (N_8555,N_7804,N_7101);
and U8556 (N_8556,N_7186,N_7018);
or U8557 (N_8557,N_7193,N_7755);
or U8558 (N_8558,N_7253,N_7496);
and U8559 (N_8559,N_7360,N_7297);
nand U8560 (N_8560,N_7936,N_7969);
nor U8561 (N_8561,N_7840,N_7396);
and U8562 (N_8562,N_7888,N_7861);
nor U8563 (N_8563,N_7086,N_7332);
nor U8564 (N_8564,N_7107,N_7638);
or U8565 (N_8565,N_7563,N_7989);
xor U8566 (N_8566,N_7868,N_7584);
nand U8567 (N_8567,N_7652,N_7738);
nand U8568 (N_8568,N_7953,N_7103);
xnor U8569 (N_8569,N_7937,N_7577);
or U8570 (N_8570,N_7503,N_7197);
and U8571 (N_8571,N_7003,N_7772);
nor U8572 (N_8572,N_7015,N_7092);
or U8573 (N_8573,N_7679,N_7162);
and U8574 (N_8574,N_7328,N_7541);
or U8575 (N_8575,N_7019,N_7459);
or U8576 (N_8576,N_7998,N_7211);
nor U8577 (N_8577,N_7859,N_7828);
or U8578 (N_8578,N_7200,N_7415);
xor U8579 (N_8579,N_7402,N_7765);
nand U8580 (N_8580,N_7509,N_7898);
nand U8581 (N_8581,N_7575,N_7923);
nor U8582 (N_8582,N_7441,N_7120);
or U8583 (N_8583,N_7034,N_7986);
xor U8584 (N_8584,N_7539,N_7470);
xor U8585 (N_8585,N_7815,N_7993);
nand U8586 (N_8586,N_7024,N_7208);
or U8587 (N_8587,N_7542,N_7756);
nand U8588 (N_8588,N_7768,N_7795);
xor U8589 (N_8589,N_7193,N_7649);
or U8590 (N_8590,N_7737,N_7679);
nand U8591 (N_8591,N_7861,N_7588);
nand U8592 (N_8592,N_7370,N_7907);
or U8593 (N_8593,N_7963,N_7797);
nor U8594 (N_8594,N_7054,N_7241);
or U8595 (N_8595,N_7340,N_7962);
nor U8596 (N_8596,N_7468,N_7738);
and U8597 (N_8597,N_7545,N_7017);
or U8598 (N_8598,N_7347,N_7479);
and U8599 (N_8599,N_7116,N_7346);
nand U8600 (N_8600,N_7549,N_7051);
or U8601 (N_8601,N_7884,N_7301);
or U8602 (N_8602,N_7914,N_7232);
or U8603 (N_8603,N_7923,N_7632);
nand U8604 (N_8604,N_7803,N_7062);
nand U8605 (N_8605,N_7519,N_7066);
and U8606 (N_8606,N_7290,N_7044);
xor U8607 (N_8607,N_7640,N_7512);
or U8608 (N_8608,N_7274,N_7116);
nor U8609 (N_8609,N_7906,N_7420);
nand U8610 (N_8610,N_7919,N_7244);
and U8611 (N_8611,N_7833,N_7582);
xnor U8612 (N_8612,N_7527,N_7220);
and U8613 (N_8613,N_7016,N_7284);
xor U8614 (N_8614,N_7516,N_7974);
or U8615 (N_8615,N_7224,N_7555);
xor U8616 (N_8616,N_7181,N_7546);
nand U8617 (N_8617,N_7919,N_7617);
nor U8618 (N_8618,N_7737,N_7639);
xnor U8619 (N_8619,N_7322,N_7007);
and U8620 (N_8620,N_7095,N_7219);
or U8621 (N_8621,N_7999,N_7410);
nor U8622 (N_8622,N_7618,N_7985);
and U8623 (N_8623,N_7242,N_7423);
or U8624 (N_8624,N_7114,N_7577);
and U8625 (N_8625,N_7983,N_7702);
xor U8626 (N_8626,N_7821,N_7530);
or U8627 (N_8627,N_7322,N_7186);
nand U8628 (N_8628,N_7830,N_7544);
nor U8629 (N_8629,N_7307,N_7774);
nor U8630 (N_8630,N_7454,N_7685);
nand U8631 (N_8631,N_7079,N_7987);
nor U8632 (N_8632,N_7148,N_7581);
or U8633 (N_8633,N_7461,N_7174);
and U8634 (N_8634,N_7748,N_7249);
nand U8635 (N_8635,N_7262,N_7765);
nand U8636 (N_8636,N_7946,N_7464);
nor U8637 (N_8637,N_7503,N_7580);
xor U8638 (N_8638,N_7959,N_7294);
and U8639 (N_8639,N_7291,N_7552);
nand U8640 (N_8640,N_7767,N_7869);
xor U8641 (N_8641,N_7810,N_7979);
xor U8642 (N_8642,N_7938,N_7010);
xnor U8643 (N_8643,N_7113,N_7647);
nor U8644 (N_8644,N_7005,N_7693);
nor U8645 (N_8645,N_7691,N_7205);
or U8646 (N_8646,N_7712,N_7681);
or U8647 (N_8647,N_7235,N_7600);
or U8648 (N_8648,N_7793,N_7385);
or U8649 (N_8649,N_7651,N_7868);
or U8650 (N_8650,N_7206,N_7475);
nand U8651 (N_8651,N_7783,N_7819);
or U8652 (N_8652,N_7541,N_7584);
nand U8653 (N_8653,N_7141,N_7137);
and U8654 (N_8654,N_7096,N_7750);
nor U8655 (N_8655,N_7798,N_7481);
and U8656 (N_8656,N_7113,N_7588);
or U8657 (N_8657,N_7063,N_7036);
and U8658 (N_8658,N_7233,N_7421);
nand U8659 (N_8659,N_7980,N_7041);
xor U8660 (N_8660,N_7577,N_7329);
and U8661 (N_8661,N_7081,N_7179);
or U8662 (N_8662,N_7323,N_7429);
nand U8663 (N_8663,N_7670,N_7372);
nor U8664 (N_8664,N_7430,N_7042);
nor U8665 (N_8665,N_7579,N_7274);
or U8666 (N_8666,N_7785,N_7985);
nand U8667 (N_8667,N_7920,N_7031);
nor U8668 (N_8668,N_7355,N_7731);
or U8669 (N_8669,N_7253,N_7894);
and U8670 (N_8670,N_7994,N_7089);
nor U8671 (N_8671,N_7292,N_7720);
nor U8672 (N_8672,N_7862,N_7049);
or U8673 (N_8673,N_7073,N_7488);
nand U8674 (N_8674,N_7760,N_7192);
nor U8675 (N_8675,N_7645,N_7997);
and U8676 (N_8676,N_7347,N_7087);
or U8677 (N_8677,N_7380,N_7434);
nor U8678 (N_8678,N_7656,N_7516);
nor U8679 (N_8679,N_7120,N_7949);
nand U8680 (N_8680,N_7527,N_7840);
or U8681 (N_8681,N_7356,N_7786);
xnor U8682 (N_8682,N_7606,N_7056);
and U8683 (N_8683,N_7399,N_7264);
nor U8684 (N_8684,N_7117,N_7584);
xor U8685 (N_8685,N_7001,N_7066);
nand U8686 (N_8686,N_7245,N_7596);
and U8687 (N_8687,N_7030,N_7974);
nor U8688 (N_8688,N_7463,N_7115);
and U8689 (N_8689,N_7199,N_7020);
and U8690 (N_8690,N_7960,N_7203);
or U8691 (N_8691,N_7863,N_7129);
nor U8692 (N_8692,N_7088,N_7255);
or U8693 (N_8693,N_7539,N_7535);
nand U8694 (N_8694,N_7243,N_7142);
and U8695 (N_8695,N_7760,N_7935);
and U8696 (N_8696,N_7718,N_7961);
nand U8697 (N_8697,N_7618,N_7726);
or U8698 (N_8698,N_7860,N_7310);
xnor U8699 (N_8699,N_7641,N_7402);
or U8700 (N_8700,N_7016,N_7203);
nand U8701 (N_8701,N_7374,N_7002);
and U8702 (N_8702,N_7431,N_7399);
or U8703 (N_8703,N_7715,N_7781);
nand U8704 (N_8704,N_7021,N_7906);
nor U8705 (N_8705,N_7930,N_7049);
xor U8706 (N_8706,N_7951,N_7075);
nand U8707 (N_8707,N_7083,N_7959);
nand U8708 (N_8708,N_7002,N_7274);
nor U8709 (N_8709,N_7048,N_7003);
or U8710 (N_8710,N_7111,N_7268);
or U8711 (N_8711,N_7017,N_7855);
xnor U8712 (N_8712,N_7822,N_7203);
nand U8713 (N_8713,N_7495,N_7527);
nand U8714 (N_8714,N_7229,N_7362);
xor U8715 (N_8715,N_7155,N_7097);
xor U8716 (N_8716,N_7918,N_7169);
nor U8717 (N_8717,N_7099,N_7106);
or U8718 (N_8718,N_7574,N_7043);
nor U8719 (N_8719,N_7392,N_7683);
and U8720 (N_8720,N_7434,N_7110);
nand U8721 (N_8721,N_7779,N_7581);
nand U8722 (N_8722,N_7646,N_7184);
nand U8723 (N_8723,N_7976,N_7531);
or U8724 (N_8724,N_7720,N_7131);
nor U8725 (N_8725,N_7612,N_7710);
nor U8726 (N_8726,N_7761,N_7139);
nor U8727 (N_8727,N_7853,N_7474);
nand U8728 (N_8728,N_7072,N_7413);
nand U8729 (N_8729,N_7613,N_7849);
and U8730 (N_8730,N_7098,N_7214);
or U8731 (N_8731,N_7814,N_7064);
nand U8732 (N_8732,N_7277,N_7164);
nor U8733 (N_8733,N_7177,N_7748);
nand U8734 (N_8734,N_7911,N_7742);
nor U8735 (N_8735,N_7039,N_7640);
nand U8736 (N_8736,N_7666,N_7174);
nor U8737 (N_8737,N_7160,N_7516);
and U8738 (N_8738,N_7472,N_7192);
or U8739 (N_8739,N_7742,N_7253);
or U8740 (N_8740,N_7990,N_7112);
or U8741 (N_8741,N_7695,N_7242);
nor U8742 (N_8742,N_7612,N_7771);
or U8743 (N_8743,N_7964,N_7595);
and U8744 (N_8744,N_7258,N_7607);
and U8745 (N_8745,N_7545,N_7607);
nand U8746 (N_8746,N_7503,N_7886);
nor U8747 (N_8747,N_7645,N_7968);
nand U8748 (N_8748,N_7602,N_7392);
and U8749 (N_8749,N_7127,N_7692);
xnor U8750 (N_8750,N_7420,N_7855);
and U8751 (N_8751,N_7441,N_7810);
nand U8752 (N_8752,N_7979,N_7463);
nand U8753 (N_8753,N_7178,N_7475);
nand U8754 (N_8754,N_7577,N_7802);
nor U8755 (N_8755,N_7963,N_7981);
nand U8756 (N_8756,N_7045,N_7179);
nor U8757 (N_8757,N_7694,N_7356);
and U8758 (N_8758,N_7418,N_7168);
nor U8759 (N_8759,N_7202,N_7997);
nor U8760 (N_8760,N_7289,N_7927);
nand U8761 (N_8761,N_7647,N_7404);
nor U8762 (N_8762,N_7358,N_7312);
xnor U8763 (N_8763,N_7663,N_7126);
nand U8764 (N_8764,N_7899,N_7147);
and U8765 (N_8765,N_7686,N_7244);
nor U8766 (N_8766,N_7805,N_7070);
and U8767 (N_8767,N_7492,N_7459);
nand U8768 (N_8768,N_7504,N_7913);
nor U8769 (N_8769,N_7812,N_7295);
and U8770 (N_8770,N_7459,N_7069);
and U8771 (N_8771,N_7103,N_7368);
or U8772 (N_8772,N_7743,N_7113);
nor U8773 (N_8773,N_7343,N_7604);
or U8774 (N_8774,N_7441,N_7174);
xor U8775 (N_8775,N_7069,N_7305);
nand U8776 (N_8776,N_7880,N_7965);
nand U8777 (N_8777,N_7724,N_7351);
nand U8778 (N_8778,N_7837,N_7094);
xnor U8779 (N_8779,N_7361,N_7599);
nand U8780 (N_8780,N_7724,N_7883);
nand U8781 (N_8781,N_7102,N_7814);
or U8782 (N_8782,N_7567,N_7235);
and U8783 (N_8783,N_7972,N_7552);
and U8784 (N_8784,N_7129,N_7857);
nand U8785 (N_8785,N_7498,N_7846);
nand U8786 (N_8786,N_7162,N_7674);
or U8787 (N_8787,N_7871,N_7590);
nor U8788 (N_8788,N_7348,N_7042);
nand U8789 (N_8789,N_7642,N_7328);
or U8790 (N_8790,N_7624,N_7141);
nor U8791 (N_8791,N_7069,N_7577);
nand U8792 (N_8792,N_7669,N_7508);
nand U8793 (N_8793,N_7303,N_7057);
nand U8794 (N_8794,N_7294,N_7983);
nor U8795 (N_8795,N_7322,N_7247);
or U8796 (N_8796,N_7140,N_7008);
nand U8797 (N_8797,N_7204,N_7403);
nor U8798 (N_8798,N_7010,N_7495);
nand U8799 (N_8799,N_7348,N_7729);
nand U8800 (N_8800,N_7348,N_7618);
nand U8801 (N_8801,N_7947,N_7590);
nor U8802 (N_8802,N_7777,N_7859);
xor U8803 (N_8803,N_7186,N_7642);
nor U8804 (N_8804,N_7638,N_7509);
and U8805 (N_8805,N_7634,N_7275);
or U8806 (N_8806,N_7580,N_7628);
nand U8807 (N_8807,N_7998,N_7906);
and U8808 (N_8808,N_7325,N_7850);
nand U8809 (N_8809,N_7573,N_7168);
or U8810 (N_8810,N_7569,N_7102);
nand U8811 (N_8811,N_7419,N_7810);
nand U8812 (N_8812,N_7186,N_7429);
or U8813 (N_8813,N_7706,N_7891);
xor U8814 (N_8814,N_7516,N_7921);
xnor U8815 (N_8815,N_7672,N_7653);
and U8816 (N_8816,N_7972,N_7225);
nor U8817 (N_8817,N_7114,N_7573);
nand U8818 (N_8818,N_7580,N_7049);
nor U8819 (N_8819,N_7674,N_7789);
and U8820 (N_8820,N_7518,N_7915);
nand U8821 (N_8821,N_7607,N_7516);
or U8822 (N_8822,N_7471,N_7717);
or U8823 (N_8823,N_7316,N_7908);
or U8824 (N_8824,N_7219,N_7296);
nand U8825 (N_8825,N_7668,N_7113);
and U8826 (N_8826,N_7305,N_7766);
nand U8827 (N_8827,N_7381,N_7336);
and U8828 (N_8828,N_7224,N_7249);
nor U8829 (N_8829,N_7093,N_7050);
or U8830 (N_8830,N_7538,N_7824);
nand U8831 (N_8831,N_7558,N_7201);
or U8832 (N_8832,N_7985,N_7039);
nor U8833 (N_8833,N_7426,N_7500);
and U8834 (N_8834,N_7638,N_7120);
nand U8835 (N_8835,N_7808,N_7398);
and U8836 (N_8836,N_7176,N_7076);
nand U8837 (N_8837,N_7915,N_7855);
nor U8838 (N_8838,N_7461,N_7353);
or U8839 (N_8839,N_7342,N_7122);
nor U8840 (N_8840,N_7518,N_7051);
or U8841 (N_8841,N_7735,N_7673);
or U8842 (N_8842,N_7778,N_7563);
nor U8843 (N_8843,N_7897,N_7444);
xor U8844 (N_8844,N_7286,N_7703);
xor U8845 (N_8845,N_7543,N_7936);
or U8846 (N_8846,N_7217,N_7068);
or U8847 (N_8847,N_7556,N_7424);
or U8848 (N_8848,N_7491,N_7864);
and U8849 (N_8849,N_7129,N_7799);
or U8850 (N_8850,N_7797,N_7366);
nor U8851 (N_8851,N_7660,N_7758);
xor U8852 (N_8852,N_7972,N_7036);
and U8853 (N_8853,N_7078,N_7954);
nor U8854 (N_8854,N_7255,N_7483);
nand U8855 (N_8855,N_7892,N_7666);
nand U8856 (N_8856,N_7698,N_7581);
and U8857 (N_8857,N_7166,N_7357);
xor U8858 (N_8858,N_7980,N_7782);
nor U8859 (N_8859,N_7866,N_7956);
nor U8860 (N_8860,N_7736,N_7599);
xor U8861 (N_8861,N_7668,N_7205);
and U8862 (N_8862,N_7168,N_7817);
and U8863 (N_8863,N_7494,N_7917);
and U8864 (N_8864,N_7609,N_7752);
nor U8865 (N_8865,N_7610,N_7450);
xnor U8866 (N_8866,N_7041,N_7398);
and U8867 (N_8867,N_7925,N_7172);
and U8868 (N_8868,N_7816,N_7854);
nor U8869 (N_8869,N_7480,N_7074);
or U8870 (N_8870,N_7948,N_7921);
nand U8871 (N_8871,N_7228,N_7607);
nor U8872 (N_8872,N_7386,N_7909);
or U8873 (N_8873,N_7041,N_7943);
nand U8874 (N_8874,N_7706,N_7817);
nand U8875 (N_8875,N_7062,N_7392);
or U8876 (N_8876,N_7438,N_7681);
xor U8877 (N_8877,N_7836,N_7385);
and U8878 (N_8878,N_7763,N_7810);
xnor U8879 (N_8879,N_7894,N_7412);
nor U8880 (N_8880,N_7896,N_7600);
nand U8881 (N_8881,N_7316,N_7005);
xor U8882 (N_8882,N_7867,N_7794);
xnor U8883 (N_8883,N_7842,N_7127);
and U8884 (N_8884,N_7446,N_7787);
or U8885 (N_8885,N_7953,N_7182);
and U8886 (N_8886,N_7823,N_7348);
nor U8887 (N_8887,N_7807,N_7808);
and U8888 (N_8888,N_7021,N_7963);
or U8889 (N_8889,N_7640,N_7069);
and U8890 (N_8890,N_7678,N_7632);
xor U8891 (N_8891,N_7356,N_7838);
and U8892 (N_8892,N_7728,N_7142);
and U8893 (N_8893,N_7125,N_7516);
nand U8894 (N_8894,N_7056,N_7317);
xnor U8895 (N_8895,N_7718,N_7515);
or U8896 (N_8896,N_7828,N_7267);
nand U8897 (N_8897,N_7249,N_7062);
and U8898 (N_8898,N_7125,N_7646);
nand U8899 (N_8899,N_7562,N_7999);
nand U8900 (N_8900,N_7412,N_7172);
nand U8901 (N_8901,N_7428,N_7885);
and U8902 (N_8902,N_7469,N_7700);
nand U8903 (N_8903,N_7522,N_7431);
or U8904 (N_8904,N_7757,N_7370);
nand U8905 (N_8905,N_7405,N_7842);
xnor U8906 (N_8906,N_7318,N_7822);
xnor U8907 (N_8907,N_7150,N_7807);
nand U8908 (N_8908,N_7396,N_7969);
and U8909 (N_8909,N_7883,N_7317);
nor U8910 (N_8910,N_7745,N_7390);
nand U8911 (N_8911,N_7712,N_7857);
nor U8912 (N_8912,N_7349,N_7738);
and U8913 (N_8913,N_7318,N_7087);
xnor U8914 (N_8914,N_7331,N_7298);
nor U8915 (N_8915,N_7488,N_7392);
xnor U8916 (N_8916,N_7586,N_7088);
and U8917 (N_8917,N_7041,N_7310);
nand U8918 (N_8918,N_7021,N_7214);
or U8919 (N_8919,N_7501,N_7108);
nor U8920 (N_8920,N_7699,N_7584);
and U8921 (N_8921,N_7881,N_7342);
nand U8922 (N_8922,N_7531,N_7461);
and U8923 (N_8923,N_7191,N_7986);
xor U8924 (N_8924,N_7105,N_7740);
nand U8925 (N_8925,N_7626,N_7421);
and U8926 (N_8926,N_7738,N_7920);
or U8927 (N_8927,N_7461,N_7346);
nand U8928 (N_8928,N_7970,N_7535);
and U8929 (N_8929,N_7511,N_7466);
nor U8930 (N_8930,N_7115,N_7439);
or U8931 (N_8931,N_7277,N_7149);
or U8932 (N_8932,N_7830,N_7158);
nor U8933 (N_8933,N_7676,N_7215);
or U8934 (N_8934,N_7497,N_7490);
nand U8935 (N_8935,N_7348,N_7739);
nand U8936 (N_8936,N_7298,N_7254);
or U8937 (N_8937,N_7730,N_7142);
and U8938 (N_8938,N_7754,N_7104);
xor U8939 (N_8939,N_7006,N_7214);
or U8940 (N_8940,N_7680,N_7262);
nand U8941 (N_8941,N_7690,N_7302);
nand U8942 (N_8942,N_7319,N_7807);
or U8943 (N_8943,N_7398,N_7356);
and U8944 (N_8944,N_7500,N_7044);
nand U8945 (N_8945,N_7369,N_7347);
or U8946 (N_8946,N_7667,N_7964);
nor U8947 (N_8947,N_7420,N_7637);
or U8948 (N_8948,N_7139,N_7104);
nor U8949 (N_8949,N_7148,N_7692);
or U8950 (N_8950,N_7999,N_7235);
nor U8951 (N_8951,N_7561,N_7263);
or U8952 (N_8952,N_7156,N_7264);
and U8953 (N_8953,N_7839,N_7093);
or U8954 (N_8954,N_7105,N_7868);
nor U8955 (N_8955,N_7066,N_7814);
and U8956 (N_8956,N_7478,N_7004);
and U8957 (N_8957,N_7880,N_7755);
nand U8958 (N_8958,N_7026,N_7190);
nor U8959 (N_8959,N_7375,N_7534);
nor U8960 (N_8960,N_7170,N_7848);
or U8961 (N_8961,N_7915,N_7851);
nor U8962 (N_8962,N_7818,N_7121);
nand U8963 (N_8963,N_7731,N_7042);
and U8964 (N_8964,N_7576,N_7817);
nor U8965 (N_8965,N_7135,N_7133);
xnor U8966 (N_8966,N_7594,N_7826);
xnor U8967 (N_8967,N_7209,N_7056);
nor U8968 (N_8968,N_7274,N_7688);
or U8969 (N_8969,N_7353,N_7855);
nor U8970 (N_8970,N_7408,N_7377);
nand U8971 (N_8971,N_7565,N_7569);
and U8972 (N_8972,N_7684,N_7383);
xor U8973 (N_8973,N_7816,N_7393);
or U8974 (N_8974,N_7337,N_7548);
nor U8975 (N_8975,N_7800,N_7214);
and U8976 (N_8976,N_7098,N_7482);
and U8977 (N_8977,N_7260,N_7438);
and U8978 (N_8978,N_7195,N_7564);
or U8979 (N_8979,N_7470,N_7978);
xnor U8980 (N_8980,N_7579,N_7762);
or U8981 (N_8981,N_7615,N_7833);
or U8982 (N_8982,N_7227,N_7866);
nor U8983 (N_8983,N_7194,N_7624);
nor U8984 (N_8984,N_7915,N_7346);
or U8985 (N_8985,N_7711,N_7343);
or U8986 (N_8986,N_7615,N_7309);
nand U8987 (N_8987,N_7008,N_7036);
and U8988 (N_8988,N_7013,N_7582);
xor U8989 (N_8989,N_7215,N_7312);
or U8990 (N_8990,N_7114,N_7448);
or U8991 (N_8991,N_7425,N_7841);
nand U8992 (N_8992,N_7709,N_7206);
nand U8993 (N_8993,N_7928,N_7667);
and U8994 (N_8994,N_7743,N_7602);
and U8995 (N_8995,N_7293,N_7791);
nand U8996 (N_8996,N_7936,N_7712);
and U8997 (N_8997,N_7545,N_7427);
nor U8998 (N_8998,N_7453,N_7648);
nor U8999 (N_8999,N_7516,N_7350);
nand U9000 (N_9000,N_8010,N_8671);
nand U9001 (N_9001,N_8889,N_8607);
nor U9002 (N_9002,N_8481,N_8108);
or U9003 (N_9003,N_8610,N_8325);
xnor U9004 (N_9004,N_8077,N_8960);
and U9005 (N_9005,N_8296,N_8052);
and U9006 (N_9006,N_8716,N_8431);
and U9007 (N_9007,N_8830,N_8099);
nor U9008 (N_9008,N_8012,N_8947);
and U9009 (N_9009,N_8323,N_8213);
nor U9010 (N_9010,N_8111,N_8879);
and U9011 (N_9011,N_8191,N_8138);
and U9012 (N_9012,N_8819,N_8901);
and U9013 (N_9013,N_8432,N_8676);
and U9014 (N_9014,N_8264,N_8083);
or U9015 (N_9015,N_8789,N_8686);
and U9016 (N_9016,N_8179,N_8496);
and U9017 (N_9017,N_8275,N_8386);
nand U9018 (N_9018,N_8519,N_8524);
and U9019 (N_9019,N_8211,N_8096);
nand U9020 (N_9020,N_8482,N_8982);
nand U9021 (N_9021,N_8801,N_8362);
or U9022 (N_9022,N_8422,N_8187);
nand U9023 (N_9023,N_8469,N_8377);
xor U9024 (N_9024,N_8603,N_8932);
xor U9025 (N_9025,N_8375,N_8544);
nand U9026 (N_9026,N_8502,N_8844);
nor U9027 (N_9027,N_8445,N_8641);
nor U9028 (N_9028,N_8270,N_8841);
or U9029 (N_9029,N_8669,N_8295);
nand U9030 (N_9030,N_8221,N_8451);
and U9031 (N_9031,N_8708,N_8692);
nor U9032 (N_9032,N_8536,N_8132);
or U9033 (N_9033,N_8137,N_8840);
or U9034 (N_9034,N_8910,N_8929);
and U9035 (N_9035,N_8827,N_8113);
nand U9036 (N_9036,N_8399,N_8691);
nor U9037 (N_9037,N_8870,N_8144);
and U9038 (N_9038,N_8632,N_8517);
nand U9039 (N_9039,N_8775,N_8157);
nor U9040 (N_9040,N_8437,N_8250);
or U9041 (N_9041,N_8762,N_8049);
or U9042 (N_9042,N_8571,N_8036);
and U9043 (N_9043,N_8050,N_8882);
nand U9044 (N_9044,N_8467,N_8818);
and U9045 (N_9045,N_8635,N_8204);
and U9046 (N_9046,N_8913,N_8555);
xor U9047 (N_9047,N_8575,N_8673);
or U9048 (N_9048,N_8232,N_8890);
nand U9049 (N_9049,N_8941,N_8547);
nand U9050 (N_9050,N_8243,N_8118);
or U9051 (N_9051,N_8831,N_8230);
nor U9052 (N_9052,N_8951,N_8989);
nand U9053 (N_9053,N_8699,N_8900);
nand U9054 (N_9054,N_8899,N_8715);
nand U9055 (N_9055,N_8606,N_8219);
and U9056 (N_9056,N_8659,N_8744);
or U9057 (N_9057,N_8043,N_8513);
xnor U9058 (N_9058,N_8350,N_8162);
and U9059 (N_9059,N_8442,N_8920);
nor U9060 (N_9060,N_8541,N_8944);
nand U9061 (N_9061,N_8631,N_8680);
or U9062 (N_9062,N_8364,N_8074);
nand U9063 (N_9063,N_8620,N_8226);
xnor U9064 (N_9064,N_8491,N_8551);
and U9065 (N_9065,N_8282,N_8312);
nand U9066 (N_9066,N_8493,N_8064);
and U9067 (N_9067,N_8189,N_8988);
xor U9068 (N_9068,N_8199,N_8034);
nand U9069 (N_9069,N_8112,N_8134);
and U9070 (N_9070,N_8133,N_8677);
xor U9071 (N_9071,N_8568,N_8795);
and U9072 (N_9072,N_8057,N_8749);
and U9073 (N_9073,N_8105,N_8478);
or U9074 (N_9074,N_8558,N_8760);
nor U9075 (N_9075,N_8060,N_8942);
nand U9076 (N_9076,N_8499,N_8367);
and U9077 (N_9077,N_8428,N_8014);
nor U9078 (N_9078,N_8661,N_8436);
and U9079 (N_9079,N_8704,N_8776);
or U9080 (N_9080,N_8463,N_8668);
or U9081 (N_9081,N_8266,N_8412);
nor U9082 (N_9082,N_8100,N_8928);
nor U9083 (N_9083,N_8015,N_8905);
and U9084 (N_9084,N_8486,N_8679);
and U9085 (N_9085,N_8806,N_8538);
or U9086 (N_9086,N_8921,N_8156);
nor U9087 (N_9087,N_8590,N_8797);
nor U9088 (N_9088,N_8949,N_8021);
and U9089 (N_9089,N_8670,N_8962);
nand U9090 (N_9090,N_8549,N_8912);
nor U9091 (N_9091,N_8414,N_8824);
nand U9092 (N_9092,N_8505,N_8585);
nand U9093 (N_9093,N_8039,N_8868);
or U9094 (N_9094,N_8176,N_8572);
or U9095 (N_9095,N_8365,N_8835);
nand U9096 (N_9096,N_8854,N_8820);
or U9097 (N_9097,N_8031,N_8847);
xnor U9098 (N_9098,N_8542,N_8501);
or U9099 (N_9099,N_8244,N_8896);
and U9100 (N_9100,N_8135,N_8618);
or U9101 (N_9101,N_8209,N_8790);
and U9102 (N_9102,N_8201,N_8294);
xor U9103 (N_9103,N_8041,N_8741);
or U9104 (N_9104,N_8088,N_8403);
nand U9105 (N_9105,N_8914,N_8602);
nand U9106 (N_9106,N_8061,N_8999);
or U9107 (N_9107,N_8177,N_8883);
nand U9108 (N_9108,N_8884,N_8344);
nand U9109 (N_9109,N_8856,N_8102);
nor U9110 (N_9110,N_8101,N_8146);
and U9111 (N_9111,N_8598,N_8685);
and U9112 (N_9112,N_8843,N_8907);
or U9113 (N_9113,N_8583,N_8340);
or U9114 (N_9114,N_8167,N_8268);
nand U9115 (N_9115,N_8004,N_8131);
nor U9116 (N_9116,N_8527,N_8310);
and U9117 (N_9117,N_8263,N_8522);
or U9118 (N_9118,N_8233,N_8466);
or U9119 (N_9119,N_8056,N_8755);
and U9120 (N_9120,N_8611,N_8409);
and U9121 (N_9121,N_8357,N_8448);
and U9122 (N_9122,N_8277,N_8693);
nand U9123 (N_9123,N_8290,N_8013);
and U9124 (N_9124,N_8750,N_8609);
and U9125 (N_9125,N_8302,N_8867);
or U9126 (N_9126,N_8717,N_8588);
nor U9127 (N_9127,N_8161,N_8805);
and U9128 (N_9128,N_8388,N_8695);
and U9129 (N_9129,N_8361,N_8175);
and U9130 (N_9130,N_8044,N_8553);
or U9131 (N_9131,N_8022,N_8887);
nand U9132 (N_9132,N_8577,N_8576);
and U9133 (N_9133,N_8771,N_8550);
and U9134 (N_9134,N_8793,N_8308);
nor U9135 (N_9135,N_8279,N_8997);
or U9136 (N_9136,N_8153,N_8791);
and U9137 (N_9137,N_8053,N_8251);
or U9138 (N_9138,N_8981,N_8188);
nor U9139 (N_9139,N_8915,N_8166);
nor U9140 (N_9140,N_8616,N_8121);
nor U9141 (N_9141,N_8589,N_8937);
or U9142 (N_9142,N_8648,N_8378);
xor U9143 (N_9143,N_8712,N_8332);
or U9144 (N_9144,N_8086,N_8666);
xnor U9145 (N_9145,N_8515,N_8816);
nand U9146 (N_9146,N_8371,N_8390);
xor U9147 (N_9147,N_8238,N_8778);
or U9148 (N_9148,N_8169,N_8917);
nor U9149 (N_9149,N_8823,N_8028);
nor U9150 (N_9150,N_8253,N_8278);
nor U9151 (N_9151,N_8009,N_8126);
nor U9152 (N_9152,N_8461,N_8506);
nand U9153 (N_9153,N_8207,N_8338);
nor U9154 (N_9154,N_8069,N_8785);
and U9155 (N_9155,N_8281,N_8839);
or U9156 (N_9156,N_8368,N_8995);
nand U9157 (N_9157,N_8956,N_8392);
xor U9158 (N_9158,N_8435,N_8065);
and U9159 (N_9159,N_8430,N_8600);
nor U9160 (N_9160,N_8417,N_8683);
xor U9161 (N_9161,N_8614,N_8552);
nand U9162 (N_9162,N_8411,N_8051);
or U9163 (N_9163,N_8406,N_8173);
or U9164 (N_9164,N_8186,N_8834);
nand U9165 (N_9165,N_8045,N_8407);
and U9166 (N_9166,N_8998,N_8694);
nor U9167 (N_9167,N_8143,N_8637);
or U9168 (N_9168,N_8617,N_8892);
nor U9169 (N_9169,N_8927,N_8678);
or U9170 (N_9170,N_8537,N_8684);
or U9171 (N_9171,N_8489,N_8347);
or U9172 (N_9172,N_8986,N_8713);
nand U9173 (N_9173,N_8287,N_8836);
nor U9174 (N_9174,N_8525,N_8581);
nor U9175 (N_9175,N_8540,N_8814);
nand U9176 (N_9176,N_8545,N_8740);
or U9177 (N_9177,N_8218,N_8151);
nor U9178 (N_9178,N_8688,N_8971);
xnor U9179 (N_9179,N_8701,N_8654);
and U9180 (N_9180,N_8756,N_8376);
and U9181 (N_9181,N_8068,N_8649);
or U9182 (N_9182,N_8359,N_8363);
nor U9183 (N_9183,N_8297,N_8024);
nor U9184 (N_9184,N_8252,N_8935);
and U9185 (N_9185,N_8301,N_8825);
nand U9186 (N_9186,N_8745,N_8521);
or U9187 (N_9187,N_8107,N_8786);
and U9188 (N_9188,N_8062,N_8084);
or U9189 (N_9189,N_8863,N_8950);
and U9190 (N_9190,N_8869,N_8122);
xnor U9191 (N_9191,N_8384,N_8289);
nor U9192 (N_9192,N_8815,N_8042);
and U9193 (N_9193,N_8373,N_8063);
or U9194 (N_9194,N_8897,N_8002);
nand U9195 (N_9195,N_8656,N_8346);
nor U9196 (N_9196,N_8738,N_8228);
and U9197 (N_9197,N_8531,N_8405);
and U9198 (N_9198,N_8242,N_8873);
xor U9199 (N_9199,N_8647,N_8240);
and U9200 (N_9200,N_8416,N_8858);
xnor U9201 (N_9201,N_8706,N_8546);
or U9202 (N_9202,N_8994,N_8705);
nand U9203 (N_9203,N_8509,N_8163);
and U9204 (N_9204,N_8198,N_8339);
nand U9205 (N_9205,N_8450,N_8140);
nor U9206 (N_9206,N_8639,N_8098);
and U9207 (N_9207,N_8970,N_8472);
nor U9208 (N_9208,N_8774,N_8474);
nand U9209 (N_9209,N_8303,N_8514);
nor U9210 (N_9210,N_8352,N_8492);
or U9211 (N_9211,N_8440,N_8732);
nand U9212 (N_9212,N_8961,N_8237);
nand U9213 (N_9213,N_8728,N_8424);
or U9214 (N_9214,N_8979,N_8320);
xor U9215 (N_9215,N_8154,N_8192);
and U9216 (N_9216,N_8908,N_8016);
nand U9217 (N_9217,N_8798,N_8828);
and U9218 (N_9218,N_8934,N_8566);
nor U9219 (N_9219,N_8120,N_8066);
or U9220 (N_9220,N_8996,N_8646);
nor U9221 (N_9221,N_8473,N_8922);
or U9222 (N_9222,N_8626,N_8599);
and U9223 (N_9223,N_8909,N_8202);
and U9224 (N_9224,N_8484,N_8130);
nand U9225 (N_9225,N_8342,N_8300);
nand U9226 (N_9226,N_8220,N_8718);
nand U9227 (N_9227,N_8249,N_8773);
nor U9228 (N_9228,N_8963,N_8259);
nor U9229 (N_9229,N_8597,N_8413);
nor U9230 (N_9230,N_8579,N_8565);
and U9231 (N_9231,N_8807,N_8800);
and U9232 (N_9232,N_8593,N_8382);
and U9233 (N_9233,N_8817,N_8345);
or U9234 (N_9234,N_8214,N_8256);
nor U9235 (N_9235,N_8168,N_8073);
and U9236 (N_9236,N_8881,N_8980);
or U9237 (N_9237,N_8293,N_8488);
xor U9238 (N_9238,N_8324,N_8257);
xor U9239 (N_9239,N_8385,N_8446);
or U9240 (N_9240,N_8005,N_8076);
nor U9241 (N_9241,N_8660,N_8203);
or U9242 (N_9242,N_8563,N_8742);
nand U9243 (N_9243,N_8709,N_8562);
and U9244 (N_9244,N_8337,N_8753);
nor U9245 (N_9245,N_8075,N_8178);
or U9246 (N_9246,N_8781,N_8370);
nand U9247 (N_9247,N_8149,N_8878);
or U9248 (N_9248,N_8276,N_8967);
and U9249 (N_9249,N_8707,N_8723);
or U9250 (N_9250,N_8595,N_8148);
nand U9251 (N_9251,N_8852,N_8846);
nand U9252 (N_9252,N_8080,N_8453);
or U9253 (N_9253,N_8480,N_8455);
or U9254 (N_9254,N_8059,N_8658);
nand U9255 (N_9255,N_8622,N_8040);
and U9256 (N_9256,N_8369,N_8582);
and U9257 (N_9257,N_8283,N_8530);
or U9258 (N_9258,N_8485,N_8425);
and U9259 (N_9259,N_8462,N_8439);
and U9260 (N_9260,N_8821,N_8444);
or U9261 (N_9261,N_8808,N_8532);
xor U9262 (N_9262,N_8398,N_8212);
or U9263 (N_9263,N_8174,N_8329);
xnor U9264 (N_9264,N_8700,N_8615);
or U9265 (N_9265,N_8939,N_8751);
nor U9266 (N_9266,N_8930,N_8667);
nor U9267 (N_9267,N_8159,N_8262);
nor U9268 (N_9268,N_8826,N_8833);
and U9269 (N_9269,N_8001,N_8458);
and U9270 (N_9270,N_8861,N_8341);
and U9271 (N_9271,N_8427,N_8477);
xor U9272 (N_9272,N_8587,N_8292);
nor U9273 (N_9273,N_8507,N_8539);
nand U9274 (N_9274,N_8965,N_8418);
nor U9275 (N_9275,N_8011,N_8943);
nand U9276 (N_9276,N_8327,N_8594);
nand U9277 (N_9277,N_8619,N_8229);
and U9278 (N_9278,N_8623,N_8239);
nor U9279 (N_9279,N_8383,N_8419);
nand U9280 (N_9280,N_8802,N_8360);
nand U9281 (N_9281,N_8969,N_8196);
nor U9282 (N_9282,N_8983,N_8812);
xnor U9283 (N_9283,N_8380,N_8119);
nor U9284 (N_9284,N_8125,N_8772);
and U9285 (N_9285,N_8180,N_8567);
nand U9286 (N_9286,N_8330,N_8271);
or U9287 (N_9287,N_8093,N_8464);
and U9288 (N_9288,N_8946,N_8309);
and U9289 (N_9289,N_8494,N_8316);
or U9290 (N_9290,N_8813,N_8027);
nor U9291 (N_9291,N_8657,N_8497);
or U9292 (N_9292,N_8636,N_8629);
nor U9293 (N_9293,N_8460,N_8698);
and U9294 (N_9294,N_8182,N_8903);
and U9295 (N_9295,N_8246,N_8940);
nand U9296 (N_9296,N_8895,N_8644);
or U9297 (N_9297,N_8006,N_8394);
and U9298 (N_9298,N_8033,N_8334);
xnor U9299 (N_9299,N_8569,N_8029);
nor U9300 (N_9300,N_8945,N_8048);
and U9301 (N_9301,N_8205,N_8315);
nor U9302 (N_9302,N_8089,N_8170);
nor U9303 (N_9303,N_8248,N_8675);
or U9304 (N_9304,N_8952,N_8366);
nand U9305 (N_9305,N_8613,N_8853);
nand U9306 (N_9306,N_8008,N_8110);
xor U9307 (N_9307,N_8880,N_8722);
nor U9308 (N_9308,N_8231,N_8779);
nand U9309 (N_9309,N_8559,N_8328);
nand U9310 (N_9310,N_8643,N_8020);
nand U9311 (N_9311,N_8687,N_8272);
or U9312 (N_9312,N_8142,N_8987);
or U9313 (N_9313,N_8591,N_8862);
nand U9314 (N_9314,N_8782,N_8254);
and U9315 (N_9315,N_8580,N_8193);
xor U9316 (N_9316,N_8739,N_8794);
or U9317 (N_9317,N_8586,N_8314);
and U9318 (N_9318,N_8288,N_8109);
or U9319 (N_9319,N_8465,N_8087);
and U9320 (N_9320,N_8627,N_8351);
nor U9321 (N_9321,N_8702,N_8401);
xor U9322 (N_9322,N_8958,N_8150);
nor U9323 (N_9323,N_8933,N_8495);
nor U9324 (N_9324,N_8047,N_8396);
or U9325 (N_9325,N_8387,N_8926);
or U9326 (N_9326,N_8007,N_8758);
nor U9327 (N_9327,N_8936,N_8025);
or U9328 (N_9328,N_8748,N_8645);
nand U9329 (N_9329,N_8037,N_8190);
nand U9330 (N_9330,N_8759,N_8129);
xnor U9331 (N_9331,N_8886,N_8145);
nor U9332 (N_9332,N_8117,N_8092);
nand U9333 (N_9333,N_8333,N_8877);
xnor U9334 (N_9334,N_8682,N_8054);
or U9335 (N_9335,N_8754,N_8625);
and U9336 (N_9336,N_8978,N_8311);
nand U9337 (N_9337,N_8123,N_8402);
nor U9338 (N_9338,N_8181,N_8690);
nor U9339 (N_9339,N_8662,N_8959);
nand U9340 (N_9340,N_8924,N_8822);
or U9341 (N_9341,N_8026,N_8584);
nor U9342 (N_9342,N_8923,N_8955);
nor U9343 (N_9343,N_8269,N_8761);
nor U9344 (N_9344,N_8734,N_8479);
nor U9345 (N_9345,N_8082,N_8948);
nor U9346 (N_9346,N_8245,N_8318);
and U9347 (N_9347,N_8729,N_8765);
and U9348 (N_9348,N_8714,N_8938);
or U9349 (N_9349,N_8184,N_8395);
nand U9350 (N_9350,N_8183,N_8236);
or U9351 (N_9351,N_8993,N_8067);
or U9352 (N_9352,N_8106,N_8241);
nand U9353 (N_9353,N_8898,N_8261);
xnor U9354 (N_9354,N_8857,N_8404);
nor U9355 (N_9355,N_8234,N_8449);
or U9356 (N_9356,N_8274,N_8511);
and U9357 (N_9357,N_8185,N_8094);
and U9358 (N_9358,N_8003,N_8888);
nand U9359 (N_9359,N_8265,N_8114);
nor U9360 (N_9360,N_8503,N_8991);
nor U9361 (N_9361,N_8103,N_8291);
nor U9362 (N_9362,N_8650,N_8916);
nor U9363 (N_9363,N_8267,N_8116);
or U9364 (N_9364,N_8307,N_8608);
xor U9365 (N_9365,N_8689,N_8072);
and U9366 (N_9366,N_8508,N_8780);
nand U9367 (N_9367,N_8319,N_8784);
and U9368 (N_9368,N_8984,N_8459);
nand U9369 (N_9369,N_8306,N_8443);
or U9370 (N_9370,N_8736,N_8155);
nor U9371 (N_9371,N_8866,N_8533);
nand U9372 (N_9372,N_8516,N_8968);
nor U9373 (N_9373,N_8849,N_8476);
xor U9374 (N_9374,N_8438,N_8081);
xor U9375 (N_9375,N_8735,N_8726);
and U9376 (N_9376,N_8147,N_8719);
nand U9377 (N_9377,N_8850,N_8095);
nand U9378 (N_9378,N_8642,N_8408);
or U9379 (N_9379,N_8127,N_8766);
nand U9380 (N_9380,N_8681,N_8456);
nor U9381 (N_9381,N_8471,N_8421);
nor U9382 (N_9382,N_8195,N_8372);
nor U9383 (N_9383,N_8071,N_8804);
nor U9384 (N_9384,N_8845,N_8038);
nor U9385 (N_9385,N_8746,N_8796);
nor U9386 (N_9386,N_8526,N_8215);
nor U9387 (N_9387,N_8604,N_8304);
and U9388 (N_9388,N_8097,N_8397);
and U9389 (N_9389,N_8326,N_8902);
and U9390 (N_9390,N_8470,N_8543);
nor U9391 (N_9391,N_8447,N_8172);
nor U9392 (N_9392,N_8454,N_8090);
nand U9393 (N_9393,N_8079,N_8764);
nand U9394 (N_9394,N_8855,N_8574);
and U9395 (N_9395,N_8721,N_8224);
and U9396 (N_9396,N_8355,N_8731);
or U9397 (N_9397,N_8596,N_8058);
and U9398 (N_9398,N_8164,N_8356);
nand U9399 (N_9399,N_8621,N_8730);
xor U9400 (N_9400,N_8299,N_8322);
nand U9401 (N_9401,N_8379,N_8055);
nand U9402 (N_9402,N_8030,N_8354);
or U9403 (N_9403,N_8792,N_8518);
or U9404 (N_9404,N_8872,N_8415);
nor U9405 (N_9405,N_8353,N_8601);
or U9406 (N_9406,N_8017,N_8752);
and U9407 (N_9407,N_8141,N_8763);
nor U9408 (N_9408,N_8768,N_8628);
or U9409 (N_9409,N_8651,N_8115);
nand U9410 (N_9410,N_8535,N_8992);
or U9411 (N_9411,N_8504,N_8925);
nor U9412 (N_9412,N_8973,N_8223);
and U9413 (N_9413,N_8227,N_8358);
nor U9414 (N_9414,N_8953,N_8556);
or U9415 (N_9415,N_8788,N_8838);
nand U9416 (N_9416,N_8078,N_8018);
or U9417 (N_9417,N_8171,N_8743);
nor U9418 (N_9418,N_8554,N_8747);
xnor U9419 (N_9419,N_8674,N_8136);
nor U9420 (N_9420,N_8457,N_8349);
and U9421 (N_9421,N_8104,N_8975);
and U9422 (N_9422,N_8313,N_8640);
xnor U9423 (N_9423,N_8957,N_8410);
xor U9424 (N_9424,N_8570,N_8864);
nor U9425 (N_9425,N_8810,N_8860);
and U9426 (N_9426,N_8548,N_8255);
and U9427 (N_9427,N_8468,N_8510);
or U9428 (N_9428,N_8208,N_8720);
nor U9429 (N_9429,N_8974,N_8483);
and U9430 (N_9430,N_8335,N_8634);
nor U9431 (N_9431,N_8298,N_8966);
or U9432 (N_9432,N_8128,N_8000);
or U9433 (N_9433,N_8770,N_8200);
nand U9434 (N_9434,N_8194,N_8964);
and U9435 (N_9435,N_8954,N_8217);
nand U9436 (N_9436,N_8235,N_8703);
nor U9437 (N_9437,N_8529,N_8523);
nor U9438 (N_9438,N_8374,N_8725);
or U9439 (N_9439,N_8837,N_8919);
nand U9440 (N_9440,N_8787,N_8124);
and U9441 (N_9441,N_8139,N_8475);
nor U9442 (N_9442,N_8612,N_8985);
xor U9443 (N_9443,N_8336,N_8737);
or U9444 (N_9444,N_8871,N_8560);
xor U9445 (N_9445,N_8769,N_8767);
and U9446 (N_9446,N_8803,N_8697);
nand U9447 (N_9447,N_8441,N_8592);
and U9448 (N_9448,N_8976,N_8799);
or U9449 (N_9449,N_8225,N_8426);
nor U9450 (N_9450,N_8733,N_8783);
or U9451 (N_9451,N_8757,N_8032);
or U9452 (N_9452,N_8520,N_8423);
nor U9453 (N_9453,N_8885,N_8876);
nand U9454 (N_9454,N_8904,N_8894);
nand U9455 (N_9455,N_8906,N_8638);
nand U9456 (N_9456,N_8724,N_8665);
and U9457 (N_9457,N_8165,N_8777);
or U9458 (N_9458,N_8972,N_8400);
nor U9459 (N_9459,N_8711,N_8809);
nor U9460 (N_9460,N_8664,N_8655);
and U9461 (N_9461,N_8534,N_8498);
or U9462 (N_9462,N_8990,N_8696);
nor U9463 (N_9463,N_8023,N_8393);
and U9464 (N_9464,N_8893,N_8222);
nor U9465 (N_9465,N_8273,N_8605);
xor U9466 (N_9466,N_8260,N_8490);
nor U9467 (N_9467,N_8197,N_8091);
and U9468 (N_9468,N_8381,N_8848);
nand U9469 (N_9469,N_8500,N_8210);
and U9470 (N_9470,N_8653,N_8557);
and U9471 (N_9471,N_8389,N_8811);
or U9472 (N_9472,N_8832,N_8578);
and U9473 (N_9473,N_8842,N_8727);
nor U9474 (N_9474,N_8152,N_8891);
and U9475 (N_9475,N_8286,N_8085);
xnor U9476 (N_9476,N_8829,N_8630);
nor U9477 (N_9477,N_8859,N_8317);
and U9478 (N_9478,N_8035,N_8216);
or U9479 (N_9479,N_8343,N_8046);
and U9480 (N_9480,N_8348,N_8977);
nor U9481 (N_9481,N_8874,N_8452);
nor U9482 (N_9482,N_8865,N_8573);
nor U9483 (N_9483,N_8875,N_8512);
nor U9484 (N_9484,N_8331,N_8663);
xnor U9485 (N_9485,N_8911,N_8710);
nand U9486 (N_9486,N_8420,N_8433);
nand U9487 (N_9487,N_8624,N_8019);
and U9488 (N_9488,N_8247,N_8160);
nand U9489 (N_9489,N_8528,N_8321);
or U9490 (N_9490,N_8429,N_8931);
and U9491 (N_9491,N_8284,N_8851);
or U9492 (N_9492,N_8305,N_8158);
or U9493 (N_9493,N_8285,N_8206);
nand U9494 (N_9494,N_8918,N_8564);
or U9495 (N_9495,N_8487,N_8070);
nor U9496 (N_9496,N_8391,N_8280);
nand U9497 (N_9497,N_8434,N_8652);
nand U9498 (N_9498,N_8561,N_8672);
nor U9499 (N_9499,N_8633,N_8258);
or U9500 (N_9500,N_8570,N_8223);
and U9501 (N_9501,N_8864,N_8464);
and U9502 (N_9502,N_8817,N_8851);
nand U9503 (N_9503,N_8600,N_8606);
nand U9504 (N_9504,N_8405,N_8420);
and U9505 (N_9505,N_8087,N_8147);
and U9506 (N_9506,N_8559,N_8254);
or U9507 (N_9507,N_8234,N_8684);
nor U9508 (N_9508,N_8876,N_8859);
or U9509 (N_9509,N_8575,N_8582);
or U9510 (N_9510,N_8167,N_8896);
and U9511 (N_9511,N_8492,N_8016);
and U9512 (N_9512,N_8504,N_8106);
nand U9513 (N_9513,N_8059,N_8363);
nor U9514 (N_9514,N_8872,N_8349);
and U9515 (N_9515,N_8669,N_8621);
xor U9516 (N_9516,N_8706,N_8191);
nor U9517 (N_9517,N_8923,N_8047);
xor U9518 (N_9518,N_8311,N_8451);
xor U9519 (N_9519,N_8032,N_8732);
nand U9520 (N_9520,N_8378,N_8198);
xnor U9521 (N_9521,N_8517,N_8624);
or U9522 (N_9522,N_8375,N_8237);
nor U9523 (N_9523,N_8130,N_8619);
and U9524 (N_9524,N_8116,N_8269);
nor U9525 (N_9525,N_8061,N_8995);
or U9526 (N_9526,N_8619,N_8623);
xor U9527 (N_9527,N_8590,N_8883);
nor U9528 (N_9528,N_8921,N_8205);
nand U9529 (N_9529,N_8405,N_8956);
nand U9530 (N_9530,N_8319,N_8137);
or U9531 (N_9531,N_8969,N_8008);
and U9532 (N_9532,N_8866,N_8282);
xor U9533 (N_9533,N_8539,N_8187);
nand U9534 (N_9534,N_8923,N_8795);
or U9535 (N_9535,N_8798,N_8808);
or U9536 (N_9536,N_8518,N_8458);
nand U9537 (N_9537,N_8565,N_8209);
nor U9538 (N_9538,N_8144,N_8267);
and U9539 (N_9539,N_8096,N_8623);
or U9540 (N_9540,N_8004,N_8608);
nand U9541 (N_9541,N_8368,N_8897);
or U9542 (N_9542,N_8817,N_8730);
and U9543 (N_9543,N_8027,N_8122);
xor U9544 (N_9544,N_8489,N_8373);
xor U9545 (N_9545,N_8186,N_8584);
nand U9546 (N_9546,N_8383,N_8502);
nand U9547 (N_9547,N_8933,N_8462);
xor U9548 (N_9548,N_8006,N_8014);
nor U9549 (N_9549,N_8290,N_8462);
and U9550 (N_9550,N_8004,N_8136);
and U9551 (N_9551,N_8326,N_8999);
nand U9552 (N_9552,N_8972,N_8141);
nand U9553 (N_9553,N_8825,N_8086);
and U9554 (N_9554,N_8192,N_8122);
or U9555 (N_9555,N_8060,N_8793);
or U9556 (N_9556,N_8284,N_8944);
xor U9557 (N_9557,N_8188,N_8830);
and U9558 (N_9558,N_8913,N_8078);
or U9559 (N_9559,N_8969,N_8725);
or U9560 (N_9560,N_8017,N_8580);
and U9561 (N_9561,N_8295,N_8697);
xor U9562 (N_9562,N_8887,N_8003);
and U9563 (N_9563,N_8092,N_8555);
nor U9564 (N_9564,N_8702,N_8241);
and U9565 (N_9565,N_8058,N_8564);
and U9566 (N_9566,N_8957,N_8012);
and U9567 (N_9567,N_8209,N_8011);
nand U9568 (N_9568,N_8382,N_8376);
and U9569 (N_9569,N_8559,N_8182);
or U9570 (N_9570,N_8196,N_8505);
nand U9571 (N_9571,N_8694,N_8627);
nand U9572 (N_9572,N_8782,N_8921);
nor U9573 (N_9573,N_8762,N_8048);
or U9574 (N_9574,N_8111,N_8181);
or U9575 (N_9575,N_8516,N_8996);
and U9576 (N_9576,N_8549,N_8674);
and U9577 (N_9577,N_8667,N_8949);
nand U9578 (N_9578,N_8116,N_8516);
nor U9579 (N_9579,N_8040,N_8984);
nand U9580 (N_9580,N_8894,N_8061);
nor U9581 (N_9581,N_8635,N_8747);
or U9582 (N_9582,N_8440,N_8731);
nand U9583 (N_9583,N_8161,N_8588);
nor U9584 (N_9584,N_8983,N_8533);
or U9585 (N_9585,N_8792,N_8836);
or U9586 (N_9586,N_8434,N_8859);
or U9587 (N_9587,N_8526,N_8135);
nor U9588 (N_9588,N_8537,N_8348);
and U9589 (N_9589,N_8269,N_8108);
and U9590 (N_9590,N_8975,N_8311);
nor U9591 (N_9591,N_8271,N_8521);
or U9592 (N_9592,N_8793,N_8673);
and U9593 (N_9593,N_8717,N_8538);
nand U9594 (N_9594,N_8513,N_8324);
or U9595 (N_9595,N_8388,N_8694);
nand U9596 (N_9596,N_8870,N_8329);
nor U9597 (N_9597,N_8824,N_8095);
or U9598 (N_9598,N_8864,N_8283);
or U9599 (N_9599,N_8423,N_8956);
nor U9600 (N_9600,N_8092,N_8249);
xnor U9601 (N_9601,N_8707,N_8228);
nand U9602 (N_9602,N_8225,N_8570);
and U9603 (N_9603,N_8271,N_8853);
nor U9604 (N_9604,N_8923,N_8685);
or U9605 (N_9605,N_8366,N_8587);
xor U9606 (N_9606,N_8962,N_8693);
nor U9607 (N_9607,N_8128,N_8349);
nor U9608 (N_9608,N_8877,N_8960);
or U9609 (N_9609,N_8452,N_8033);
or U9610 (N_9610,N_8970,N_8454);
or U9611 (N_9611,N_8944,N_8482);
or U9612 (N_9612,N_8089,N_8395);
nand U9613 (N_9613,N_8236,N_8062);
nand U9614 (N_9614,N_8460,N_8381);
or U9615 (N_9615,N_8186,N_8181);
nor U9616 (N_9616,N_8162,N_8243);
nand U9617 (N_9617,N_8406,N_8258);
nor U9618 (N_9618,N_8159,N_8596);
nor U9619 (N_9619,N_8699,N_8337);
and U9620 (N_9620,N_8415,N_8144);
nand U9621 (N_9621,N_8832,N_8928);
and U9622 (N_9622,N_8524,N_8279);
nand U9623 (N_9623,N_8274,N_8829);
xor U9624 (N_9624,N_8245,N_8041);
and U9625 (N_9625,N_8168,N_8814);
or U9626 (N_9626,N_8068,N_8875);
and U9627 (N_9627,N_8739,N_8259);
nor U9628 (N_9628,N_8934,N_8619);
or U9629 (N_9629,N_8045,N_8053);
xor U9630 (N_9630,N_8038,N_8252);
and U9631 (N_9631,N_8255,N_8023);
and U9632 (N_9632,N_8567,N_8044);
and U9633 (N_9633,N_8673,N_8735);
or U9634 (N_9634,N_8481,N_8900);
nor U9635 (N_9635,N_8467,N_8782);
and U9636 (N_9636,N_8623,N_8193);
nor U9637 (N_9637,N_8127,N_8800);
nand U9638 (N_9638,N_8549,N_8193);
and U9639 (N_9639,N_8649,N_8027);
or U9640 (N_9640,N_8039,N_8327);
nor U9641 (N_9641,N_8955,N_8734);
and U9642 (N_9642,N_8519,N_8188);
and U9643 (N_9643,N_8650,N_8819);
nor U9644 (N_9644,N_8737,N_8759);
nand U9645 (N_9645,N_8596,N_8627);
and U9646 (N_9646,N_8044,N_8660);
and U9647 (N_9647,N_8989,N_8460);
or U9648 (N_9648,N_8660,N_8550);
nand U9649 (N_9649,N_8663,N_8984);
or U9650 (N_9650,N_8257,N_8461);
nand U9651 (N_9651,N_8850,N_8595);
nor U9652 (N_9652,N_8642,N_8952);
xor U9653 (N_9653,N_8154,N_8002);
nand U9654 (N_9654,N_8100,N_8650);
nand U9655 (N_9655,N_8288,N_8201);
and U9656 (N_9656,N_8234,N_8932);
nor U9657 (N_9657,N_8197,N_8702);
or U9658 (N_9658,N_8479,N_8439);
or U9659 (N_9659,N_8462,N_8841);
nor U9660 (N_9660,N_8978,N_8058);
or U9661 (N_9661,N_8612,N_8867);
and U9662 (N_9662,N_8113,N_8467);
or U9663 (N_9663,N_8563,N_8113);
nor U9664 (N_9664,N_8013,N_8212);
and U9665 (N_9665,N_8609,N_8709);
and U9666 (N_9666,N_8777,N_8476);
nor U9667 (N_9667,N_8563,N_8071);
and U9668 (N_9668,N_8777,N_8891);
nor U9669 (N_9669,N_8282,N_8028);
and U9670 (N_9670,N_8821,N_8581);
nand U9671 (N_9671,N_8036,N_8670);
nor U9672 (N_9672,N_8179,N_8001);
and U9673 (N_9673,N_8115,N_8670);
and U9674 (N_9674,N_8265,N_8762);
and U9675 (N_9675,N_8615,N_8054);
and U9676 (N_9676,N_8297,N_8472);
nand U9677 (N_9677,N_8551,N_8241);
nor U9678 (N_9678,N_8287,N_8853);
nor U9679 (N_9679,N_8167,N_8045);
and U9680 (N_9680,N_8587,N_8749);
xor U9681 (N_9681,N_8568,N_8236);
nand U9682 (N_9682,N_8171,N_8057);
nand U9683 (N_9683,N_8714,N_8051);
nor U9684 (N_9684,N_8715,N_8788);
nor U9685 (N_9685,N_8361,N_8470);
and U9686 (N_9686,N_8771,N_8311);
and U9687 (N_9687,N_8688,N_8325);
nor U9688 (N_9688,N_8530,N_8815);
or U9689 (N_9689,N_8470,N_8828);
xor U9690 (N_9690,N_8848,N_8153);
or U9691 (N_9691,N_8686,N_8141);
nand U9692 (N_9692,N_8907,N_8821);
nand U9693 (N_9693,N_8858,N_8259);
and U9694 (N_9694,N_8036,N_8357);
or U9695 (N_9695,N_8884,N_8645);
and U9696 (N_9696,N_8543,N_8685);
or U9697 (N_9697,N_8425,N_8666);
or U9698 (N_9698,N_8972,N_8091);
nand U9699 (N_9699,N_8170,N_8045);
xnor U9700 (N_9700,N_8958,N_8870);
and U9701 (N_9701,N_8391,N_8844);
or U9702 (N_9702,N_8243,N_8841);
or U9703 (N_9703,N_8821,N_8842);
nor U9704 (N_9704,N_8757,N_8459);
nand U9705 (N_9705,N_8513,N_8738);
nand U9706 (N_9706,N_8610,N_8542);
and U9707 (N_9707,N_8840,N_8578);
nand U9708 (N_9708,N_8599,N_8281);
or U9709 (N_9709,N_8736,N_8789);
and U9710 (N_9710,N_8508,N_8447);
nand U9711 (N_9711,N_8323,N_8269);
nand U9712 (N_9712,N_8051,N_8889);
or U9713 (N_9713,N_8045,N_8591);
or U9714 (N_9714,N_8237,N_8065);
nand U9715 (N_9715,N_8240,N_8705);
xor U9716 (N_9716,N_8718,N_8259);
or U9717 (N_9717,N_8939,N_8635);
and U9718 (N_9718,N_8167,N_8297);
nand U9719 (N_9719,N_8143,N_8428);
nor U9720 (N_9720,N_8348,N_8137);
or U9721 (N_9721,N_8865,N_8375);
nand U9722 (N_9722,N_8870,N_8878);
nor U9723 (N_9723,N_8141,N_8504);
nand U9724 (N_9724,N_8829,N_8559);
nor U9725 (N_9725,N_8125,N_8721);
or U9726 (N_9726,N_8428,N_8080);
nor U9727 (N_9727,N_8677,N_8436);
nor U9728 (N_9728,N_8350,N_8693);
nand U9729 (N_9729,N_8624,N_8963);
and U9730 (N_9730,N_8260,N_8122);
nand U9731 (N_9731,N_8393,N_8966);
nor U9732 (N_9732,N_8065,N_8918);
xnor U9733 (N_9733,N_8056,N_8553);
nand U9734 (N_9734,N_8863,N_8724);
nand U9735 (N_9735,N_8230,N_8093);
nor U9736 (N_9736,N_8865,N_8938);
or U9737 (N_9737,N_8452,N_8214);
nor U9738 (N_9738,N_8208,N_8467);
or U9739 (N_9739,N_8966,N_8170);
or U9740 (N_9740,N_8439,N_8003);
or U9741 (N_9741,N_8787,N_8984);
nor U9742 (N_9742,N_8236,N_8995);
or U9743 (N_9743,N_8169,N_8086);
nand U9744 (N_9744,N_8530,N_8235);
nor U9745 (N_9745,N_8978,N_8387);
xor U9746 (N_9746,N_8476,N_8322);
and U9747 (N_9747,N_8468,N_8545);
xnor U9748 (N_9748,N_8718,N_8880);
and U9749 (N_9749,N_8753,N_8030);
or U9750 (N_9750,N_8790,N_8727);
or U9751 (N_9751,N_8158,N_8521);
nor U9752 (N_9752,N_8164,N_8286);
or U9753 (N_9753,N_8865,N_8110);
nand U9754 (N_9754,N_8798,N_8593);
nor U9755 (N_9755,N_8175,N_8463);
nand U9756 (N_9756,N_8231,N_8642);
or U9757 (N_9757,N_8359,N_8751);
and U9758 (N_9758,N_8305,N_8719);
or U9759 (N_9759,N_8594,N_8875);
xnor U9760 (N_9760,N_8560,N_8562);
nand U9761 (N_9761,N_8186,N_8691);
xor U9762 (N_9762,N_8591,N_8662);
or U9763 (N_9763,N_8076,N_8069);
nand U9764 (N_9764,N_8529,N_8565);
and U9765 (N_9765,N_8493,N_8710);
or U9766 (N_9766,N_8200,N_8224);
and U9767 (N_9767,N_8222,N_8869);
nor U9768 (N_9768,N_8449,N_8684);
nor U9769 (N_9769,N_8988,N_8337);
nor U9770 (N_9770,N_8412,N_8490);
and U9771 (N_9771,N_8874,N_8538);
nor U9772 (N_9772,N_8547,N_8219);
or U9773 (N_9773,N_8082,N_8122);
or U9774 (N_9774,N_8322,N_8611);
nand U9775 (N_9775,N_8722,N_8400);
and U9776 (N_9776,N_8052,N_8411);
and U9777 (N_9777,N_8868,N_8989);
nor U9778 (N_9778,N_8070,N_8241);
xnor U9779 (N_9779,N_8474,N_8076);
or U9780 (N_9780,N_8705,N_8640);
or U9781 (N_9781,N_8097,N_8793);
nor U9782 (N_9782,N_8005,N_8132);
and U9783 (N_9783,N_8107,N_8360);
nand U9784 (N_9784,N_8415,N_8155);
nand U9785 (N_9785,N_8599,N_8812);
nand U9786 (N_9786,N_8461,N_8900);
nor U9787 (N_9787,N_8877,N_8228);
or U9788 (N_9788,N_8900,N_8987);
or U9789 (N_9789,N_8794,N_8017);
and U9790 (N_9790,N_8184,N_8828);
nor U9791 (N_9791,N_8285,N_8939);
or U9792 (N_9792,N_8012,N_8964);
and U9793 (N_9793,N_8023,N_8984);
and U9794 (N_9794,N_8266,N_8998);
and U9795 (N_9795,N_8217,N_8046);
or U9796 (N_9796,N_8576,N_8233);
nor U9797 (N_9797,N_8606,N_8016);
and U9798 (N_9798,N_8515,N_8885);
nand U9799 (N_9799,N_8731,N_8299);
xnor U9800 (N_9800,N_8937,N_8998);
nor U9801 (N_9801,N_8273,N_8715);
or U9802 (N_9802,N_8122,N_8009);
nand U9803 (N_9803,N_8684,N_8952);
nor U9804 (N_9804,N_8969,N_8358);
and U9805 (N_9805,N_8778,N_8097);
nand U9806 (N_9806,N_8624,N_8159);
nor U9807 (N_9807,N_8713,N_8468);
or U9808 (N_9808,N_8969,N_8747);
or U9809 (N_9809,N_8189,N_8638);
and U9810 (N_9810,N_8766,N_8529);
nand U9811 (N_9811,N_8211,N_8992);
nor U9812 (N_9812,N_8770,N_8766);
nor U9813 (N_9813,N_8689,N_8834);
nand U9814 (N_9814,N_8183,N_8150);
nor U9815 (N_9815,N_8692,N_8875);
xnor U9816 (N_9816,N_8147,N_8496);
or U9817 (N_9817,N_8445,N_8419);
nor U9818 (N_9818,N_8776,N_8284);
nor U9819 (N_9819,N_8084,N_8069);
or U9820 (N_9820,N_8332,N_8502);
nor U9821 (N_9821,N_8643,N_8962);
nor U9822 (N_9822,N_8379,N_8426);
nor U9823 (N_9823,N_8407,N_8743);
xnor U9824 (N_9824,N_8698,N_8246);
nand U9825 (N_9825,N_8675,N_8059);
xor U9826 (N_9826,N_8511,N_8283);
nor U9827 (N_9827,N_8339,N_8938);
and U9828 (N_9828,N_8993,N_8769);
nor U9829 (N_9829,N_8057,N_8841);
or U9830 (N_9830,N_8379,N_8983);
nor U9831 (N_9831,N_8565,N_8074);
nor U9832 (N_9832,N_8413,N_8661);
nor U9833 (N_9833,N_8663,N_8196);
xor U9834 (N_9834,N_8100,N_8475);
nor U9835 (N_9835,N_8687,N_8458);
nand U9836 (N_9836,N_8598,N_8792);
nand U9837 (N_9837,N_8136,N_8189);
nor U9838 (N_9838,N_8940,N_8822);
and U9839 (N_9839,N_8092,N_8969);
or U9840 (N_9840,N_8707,N_8686);
nand U9841 (N_9841,N_8721,N_8674);
nand U9842 (N_9842,N_8493,N_8676);
nor U9843 (N_9843,N_8841,N_8292);
and U9844 (N_9844,N_8429,N_8961);
nand U9845 (N_9845,N_8156,N_8535);
nor U9846 (N_9846,N_8904,N_8544);
xor U9847 (N_9847,N_8152,N_8313);
nor U9848 (N_9848,N_8901,N_8026);
nor U9849 (N_9849,N_8868,N_8016);
nor U9850 (N_9850,N_8869,N_8739);
or U9851 (N_9851,N_8062,N_8136);
and U9852 (N_9852,N_8650,N_8351);
nor U9853 (N_9853,N_8572,N_8643);
nor U9854 (N_9854,N_8288,N_8677);
nor U9855 (N_9855,N_8635,N_8812);
and U9856 (N_9856,N_8689,N_8377);
or U9857 (N_9857,N_8275,N_8955);
or U9858 (N_9858,N_8887,N_8101);
and U9859 (N_9859,N_8232,N_8039);
nand U9860 (N_9860,N_8271,N_8466);
or U9861 (N_9861,N_8383,N_8432);
nor U9862 (N_9862,N_8283,N_8884);
or U9863 (N_9863,N_8453,N_8672);
and U9864 (N_9864,N_8260,N_8798);
nor U9865 (N_9865,N_8604,N_8763);
xor U9866 (N_9866,N_8643,N_8065);
and U9867 (N_9867,N_8521,N_8141);
nor U9868 (N_9868,N_8759,N_8279);
nor U9869 (N_9869,N_8348,N_8061);
nor U9870 (N_9870,N_8601,N_8703);
or U9871 (N_9871,N_8021,N_8887);
nand U9872 (N_9872,N_8569,N_8724);
or U9873 (N_9873,N_8361,N_8296);
and U9874 (N_9874,N_8799,N_8656);
nand U9875 (N_9875,N_8562,N_8540);
nand U9876 (N_9876,N_8077,N_8866);
nand U9877 (N_9877,N_8221,N_8857);
or U9878 (N_9878,N_8366,N_8128);
and U9879 (N_9879,N_8710,N_8158);
nor U9880 (N_9880,N_8147,N_8084);
xnor U9881 (N_9881,N_8000,N_8907);
nor U9882 (N_9882,N_8616,N_8307);
xor U9883 (N_9883,N_8631,N_8758);
xnor U9884 (N_9884,N_8922,N_8175);
nand U9885 (N_9885,N_8339,N_8812);
and U9886 (N_9886,N_8034,N_8723);
nand U9887 (N_9887,N_8601,N_8024);
nor U9888 (N_9888,N_8951,N_8952);
nor U9889 (N_9889,N_8202,N_8640);
and U9890 (N_9890,N_8472,N_8750);
and U9891 (N_9891,N_8985,N_8212);
or U9892 (N_9892,N_8206,N_8366);
xor U9893 (N_9893,N_8765,N_8962);
nand U9894 (N_9894,N_8846,N_8556);
nor U9895 (N_9895,N_8958,N_8574);
or U9896 (N_9896,N_8549,N_8228);
or U9897 (N_9897,N_8805,N_8740);
nor U9898 (N_9898,N_8077,N_8937);
and U9899 (N_9899,N_8842,N_8488);
or U9900 (N_9900,N_8554,N_8660);
nor U9901 (N_9901,N_8452,N_8084);
and U9902 (N_9902,N_8551,N_8707);
xor U9903 (N_9903,N_8534,N_8778);
nand U9904 (N_9904,N_8966,N_8164);
nor U9905 (N_9905,N_8858,N_8025);
nand U9906 (N_9906,N_8098,N_8907);
or U9907 (N_9907,N_8296,N_8379);
nor U9908 (N_9908,N_8487,N_8694);
and U9909 (N_9909,N_8649,N_8371);
xor U9910 (N_9910,N_8687,N_8081);
nand U9911 (N_9911,N_8776,N_8794);
and U9912 (N_9912,N_8496,N_8601);
nand U9913 (N_9913,N_8656,N_8598);
nand U9914 (N_9914,N_8561,N_8689);
and U9915 (N_9915,N_8675,N_8685);
nand U9916 (N_9916,N_8500,N_8445);
and U9917 (N_9917,N_8482,N_8074);
nand U9918 (N_9918,N_8844,N_8783);
or U9919 (N_9919,N_8038,N_8832);
nand U9920 (N_9920,N_8353,N_8006);
nor U9921 (N_9921,N_8874,N_8978);
nand U9922 (N_9922,N_8433,N_8466);
xnor U9923 (N_9923,N_8223,N_8089);
or U9924 (N_9924,N_8795,N_8548);
or U9925 (N_9925,N_8303,N_8532);
nand U9926 (N_9926,N_8310,N_8862);
or U9927 (N_9927,N_8088,N_8637);
or U9928 (N_9928,N_8660,N_8095);
nand U9929 (N_9929,N_8538,N_8330);
xnor U9930 (N_9930,N_8382,N_8836);
and U9931 (N_9931,N_8301,N_8645);
nor U9932 (N_9932,N_8293,N_8872);
or U9933 (N_9933,N_8812,N_8720);
nor U9934 (N_9934,N_8964,N_8531);
nand U9935 (N_9935,N_8216,N_8262);
or U9936 (N_9936,N_8911,N_8147);
nor U9937 (N_9937,N_8121,N_8159);
and U9938 (N_9938,N_8727,N_8583);
nand U9939 (N_9939,N_8844,N_8492);
or U9940 (N_9940,N_8388,N_8687);
nor U9941 (N_9941,N_8627,N_8256);
nand U9942 (N_9942,N_8703,N_8440);
nor U9943 (N_9943,N_8346,N_8941);
nand U9944 (N_9944,N_8732,N_8737);
or U9945 (N_9945,N_8087,N_8130);
nor U9946 (N_9946,N_8012,N_8332);
or U9947 (N_9947,N_8416,N_8703);
xor U9948 (N_9948,N_8244,N_8825);
and U9949 (N_9949,N_8033,N_8213);
nand U9950 (N_9950,N_8633,N_8457);
nor U9951 (N_9951,N_8319,N_8529);
nand U9952 (N_9952,N_8793,N_8547);
nor U9953 (N_9953,N_8302,N_8888);
or U9954 (N_9954,N_8591,N_8201);
nand U9955 (N_9955,N_8642,N_8558);
nand U9956 (N_9956,N_8261,N_8877);
and U9957 (N_9957,N_8053,N_8487);
nor U9958 (N_9958,N_8652,N_8188);
or U9959 (N_9959,N_8301,N_8930);
or U9960 (N_9960,N_8161,N_8190);
or U9961 (N_9961,N_8854,N_8951);
nor U9962 (N_9962,N_8730,N_8447);
or U9963 (N_9963,N_8856,N_8545);
or U9964 (N_9964,N_8982,N_8869);
or U9965 (N_9965,N_8255,N_8261);
nor U9966 (N_9966,N_8017,N_8717);
nand U9967 (N_9967,N_8294,N_8235);
or U9968 (N_9968,N_8645,N_8551);
nand U9969 (N_9969,N_8075,N_8576);
and U9970 (N_9970,N_8890,N_8544);
or U9971 (N_9971,N_8326,N_8419);
nor U9972 (N_9972,N_8984,N_8708);
nor U9973 (N_9973,N_8891,N_8815);
and U9974 (N_9974,N_8072,N_8806);
or U9975 (N_9975,N_8119,N_8136);
or U9976 (N_9976,N_8980,N_8863);
nand U9977 (N_9977,N_8540,N_8326);
nor U9978 (N_9978,N_8635,N_8110);
xnor U9979 (N_9979,N_8286,N_8042);
or U9980 (N_9980,N_8136,N_8222);
nor U9981 (N_9981,N_8138,N_8392);
nor U9982 (N_9982,N_8567,N_8038);
and U9983 (N_9983,N_8993,N_8974);
nor U9984 (N_9984,N_8719,N_8844);
and U9985 (N_9985,N_8025,N_8620);
nand U9986 (N_9986,N_8500,N_8352);
and U9987 (N_9987,N_8793,N_8830);
or U9988 (N_9988,N_8941,N_8185);
nand U9989 (N_9989,N_8488,N_8410);
and U9990 (N_9990,N_8420,N_8025);
nand U9991 (N_9991,N_8231,N_8475);
nand U9992 (N_9992,N_8765,N_8778);
xnor U9993 (N_9993,N_8215,N_8498);
nor U9994 (N_9994,N_8612,N_8077);
nand U9995 (N_9995,N_8333,N_8370);
and U9996 (N_9996,N_8506,N_8541);
nand U9997 (N_9997,N_8773,N_8540);
nor U9998 (N_9998,N_8194,N_8417);
nand U9999 (N_9999,N_8852,N_8241);
nand U10000 (N_10000,N_9637,N_9631);
and U10001 (N_10001,N_9462,N_9788);
or U10002 (N_10002,N_9095,N_9804);
and U10003 (N_10003,N_9246,N_9103);
and U10004 (N_10004,N_9740,N_9266);
and U10005 (N_10005,N_9743,N_9510);
xor U10006 (N_10006,N_9512,N_9161);
nand U10007 (N_10007,N_9793,N_9338);
or U10008 (N_10008,N_9550,N_9972);
nor U10009 (N_10009,N_9597,N_9548);
nor U10010 (N_10010,N_9998,N_9670);
and U10011 (N_10011,N_9953,N_9215);
and U10012 (N_10012,N_9817,N_9206);
nand U10013 (N_10013,N_9237,N_9946);
or U10014 (N_10014,N_9049,N_9652);
and U10015 (N_10015,N_9030,N_9446);
nand U10016 (N_10016,N_9473,N_9481);
nand U10017 (N_10017,N_9287,N_9411);
nor U10018 (N_10018,N_9355,N_9459);
nor U10019 (N_10019,N_9828,N_9630);
or U10020 (N_10020,N_9056,N_9307);
nand U10021 (N_10021,N_9867,N_9838);
and U10022 (N_10022,N_9109,N_9780);
nand U10023 (N_10023,N_9233,N_9656);
xnor U10024 (N_10024,N_9094,N_9377);
nand U10025 (N_10025,N_9019,N_9876);
nor U10026 (N_10026,N_9697,N_9937);
nand U10027 (N_10027,N_9032,N_9556);
or U10028 (N_10028,N_9523,N_9826);
and U10029 (N_10029,N_9698,N_9469);
nor U10030 (N_10030,N_9378,N_9269);
xor U10031 (N_10031,N_9513,N_9488);
and U10032 (N_10032,N_9101,N_9615);
nor U10033 (N_10033,N_9391,N_9767);
and U10034 (N_10034,N_9211,N_9640);
nor U10035 (N_10035,N_9626,N_9433);
nor U10036 (N_10036,N_9877,N_9686);
nor U10037 (N_10037,N_9969,N_9560);
or U10038 (N_10038,N_9245,N_9899);
nor U10039 (N_10039,N_9999,N_9555);
and U10040 (N_10040,N_9799,N_9334);
and U10041 (N_10041,N_9116,N_9144);
nor U10042 (N_10042,N_9022,N_9710);
nor U10043 (N_10043,N_9566,N_9408);
and U10044 (N_10044,N_9420,N_9417);
xor U10045 (N_10045,N_9127,N_9790);
nand U10046 (N_10046,N_9609,N_9750);
and U10047 (N_10047,N_9791,N_9259);
nor U10048 (N_10048,N_9718,N_9938);
nand U10049 (N_10049,N_9492,N_9039);
or U10050 (N_10050,N_9502,N_9222);
nand U10051 (N_10051,N_9661,N_9415);
nor U10052 (N_10052,N_9011,N_9342);
or U10053 (N_10053,N_9447,N_9827);
and U10054 (N_10054,N_9467,N_9141);
or U10055 (N_10055,N_9293,N_9143);
or U10056 (N_10056,N_9148,N_9238);
nand U10057 (N_10057,N_9240,N_9763);
nor U10058 (N_10058,N_9778,N_9118);
nand U10059 (N_10059,N_9450,N_9235);
and U10060 (N_10060,N_9859,N_9326);
nor U10061 (N_10061,N_9115,N_9785);
nand U10062 (N_10062,N_9691,N_9603);
nand U10063 (N_10063,N_9028,N_9419);
nand U10064 (N_10064,N_9675,N_9762);
nor U10065 (N_10065,N_9313,N_9782);
or U10066 (N_10066,N_9059,N_9552);
xnor U10067 (N_10067,N_9400,N_9715);
and U10068 (N_10068,N_9303,N_9988);
nand U10069 (N_10069,N_9783,N_9044);
xor U10070 (N_10070,N_9409,N_9163);
or U10071 (N_10071,N_9494,N_9731);
or U10072 (N_10072,N_9832,N_9021);
xnor U10073 (N_10073,N_9327,N_9680);
and U10074 (N_10074,N_9607,N_9744);
nand U10075 (N_10075,N_9191,N_9739);
or U10076 (N_10076,N_9578,N_9038);
or U10077 (N_10077,N_9296,N_9764);
nand U10078 (N_10078,N_9860,N_9166);
and U10079 (N_10079,N_9167,N_9498);
or U10080 (N_10080,N_9214,N_9186);
or U10081 (N_10081,N_9930,N_9009);
or U10082 (N_10082,N_9439,N_9920);
xnor U10083 (N_10083,N_9511,N_9933);
nand U10084 (N_10084,N_9333,N_9110);
nor U10085 (N_10085,N_9643,N_9694);
and U10086 (N_10086,N_9653,N_9903);
or U10087 (N_10087,N_9170,N_9064);
and U10088 (N_10088,N_9944,N_9181);
or U10089 (N_10089,N_9616,N_9781);
nand U10090 (N_10090,N_9406,N_9673);
and U10091 (N_10091,N_9884,N_9539);
nand U10092 (N_10092,N_9658,N_9968);
or U10093 (N_10093,N_9868,N_9445);
or U10094 (N_10094,N_9267,N_9208);
and U10095 (N_10095,N_9573,N_9225);
nand U10096 (N_10096,N_9907,N_9761);
xnor U10097 (N_10097,N_9505,N_9641);
and U10098 (N_10098,N_9796,N_9047);
nor U10099 (N_10099,N_9217,N_9325);
xnor U10100 (N_10100,N_9773,N_9986);
and U10101 (N_10101,N_9098,N_9608);
nor U10102 (N_10102,N_9332,N_9553);
nand U10103 (N_10103,N_9295,N_9359);
and U10104 (N_10104,N_9236,N_9478);
and U10105 (N_10105,N_9220,N_9557);
xor U10106 (N_10106,N_9519,N_9251);
nor U10107 (N_10107,N_9271,N_9104);
or U10108 (N_10108,N_9210,N_9702);
nor U10109 (N_10109,N_9897,N_9729);
and U10110 (N_10110,N_9132,N_9456);
nand U10111 (N_10111,N_9562,N_9894);
or U10112 (N_10112,N_9401,N_9984);
xnor U10113 (N_10113,N_9034,N_9335);
and U10114 (N_10114,N_9466,N_9169);
nor U10115 (N_10115,N_9171,N_9316);
or U10116 (N_10116,N_9881,N_9939);
or U10117 (N_10117,N_9843,N_9769);
nand U10118 (N_10118,N_9414,N_9657);
or U10119 (N_10119,N_9193,N_9042);
or U10120 (N_10120,N_9199,N_9912);
or U10121 (N_10121,N_9353,N_9974);
or U10122 (N_10122,N_9276,N_9863);
or U10123 (N_10123,N_9845,N_9412);
nor U10124 (N_10124,N_9090,N_9809);
nand U10125 (N_10125,N_9079,N_9304);
and U10126 (N_10126,N_9617,N_9003);
or U10127 (N_10127,N_9035,N_9581);
nor U10128 (N_10128,N_9213,N_9575);
nand U10129 (N_10129,N_9454,N_9219);
nand U10130 (N_10130,N_9960,N_9921);
xor U10131 (N_10131,N_9943,N_9389);
or U10132 (N_10132,N_9951,N_9465);
nor U10133 (N_10133,N_9484,N_9150);
and U10134 (N_10134,N_9458,N_9570);
nand U10135 (N_10135,N_9126,N_9544);
or U10136 (N_10136,N_9100,N_9814);
xnor U10137 (N_10137,N_9971,N_9275);
nor U10138 (N_10138,N_9692,N_9125);
nor U10139 (N_10139,N_9192,N_9178);
nand U10140 (N_10140,N_9844,N_9797);
and U10141 (N_10141,N_9298,N_9373);
or U10142 (N_10142,N_9393,N_9959);
nand U10143 (N_10143,N_9917,N_9547);
nor U10144 (N_10144,N_9374,N_9654);
or U10145 (N_10145,N_9349,N_9441);
xor U10146 (N_10146,N_9248,N_9551);
or U10147 (N_10147,N_9704,N_9591);
nand U10148 (N_10148,N_9936,N_9108);
nand U10149 (N_10149,N_9530,N_9900);
and U10150 (N_10150,N_9117,N_9932);
nand U10151 (N_10151,N_9501,N_9156);
and U10152 (N_10152,N_9157,N_9518);
or U10153 (N_10153,N_9754,N_9701);
nand U10154 (N_10154,N_9668,N_9836);
and U10155 (N_10155,N_9007,N_9075);
or U10156 (N_10156,N_9541,N_9243);
nand U10157 (N_10157,N_9872,N_9046);
nand U10158 (N_10158,N_9160,N_9187);
and U10159 (N_10159,N_9745,N_9810);
and U10160 (N_10160,N_9614,N_9565);
nor U10161 (N_10161,N_9913,N_9395);
nor U10162 (N_10162,N_9084,N_9037);
and U10163 (N_10163,N_9291,N_9436);
nand U10164 (N_10164,N_9721,N_9134);
or U10165 (N_10165,N_9283,N_9524);
nand U10166 (N_10166,N_9487,N_9013);
nor U10167 (N_10167,N_9351,N_9593);
nor U10168 (N_10168,N_9529,N_9983);
nand U10169 (N_10169,N_9674,N_9130);
nand U10170 (N_10170,N_9730,N_9273);
nor U10171 (N_10171,N_9665,N_9197);
or U10172 (N_10172,N_9711,N_9598);
and U10173 (N_10173,N_9734,N_9979);
xnor U10174 (N_10174,N_9604,N_9712);
and U10175 (N_10175,N_9212,N_9752);
nor U10176 (N_10176,N_9677,N_9423);
or U10177 (N_10177,N_9599,N_9693);
nor U10178 (N_10178,N_9493,N_9074);
or U10179 (N_10179,N_9396,N_9319);
nand U10180 (N_10180,N_9048,N_9542);
and U10181 (N_10181,N_9375,N_9128);
or U10182 (N_10182,N_9977,N_9496);
nor U10183 (N_10183,N_9757,N_9962);
and U10184 (N_10184,N_9873,N_9713);
and U10185 (N_10185,N_9402,N_9645);
or U10186 (N_10186,N_9367,N_9747);
nand U10187 (N_10187,N_9735,N_9777);
and U10188 (N_10188,N_9952,N_9310);
and U10189 (N_10189,N_9154,N_9925);
nor U10190 (N_10190,N_9870,N_9644);
and U10191 (N_10191,N_9318,N_9923);
and U10192 (N_10192,N_9379,N_9112);
xnor U10193 (N_10193,N_9250,N_9798);
nor U10194 (N_10194,N_9151,N_9323);
nand U10195 (N_10195,N_9321,N_9350);
nor U10196 (N_10196,N_9386,N_9159);
nor U10197 (N_10197,N_9795,N_9308);
nand U10198 (N_10198,N_9516,N_9070);
and U10199 (N_10199,N_9435,N_9639);
nand U10200 (N_10200,N_9619,N_9891);
or U10201 (N_10201,N_9055,N_9633);
or U10202 (N_10202,N_9612,N_9954);
nor U10203 (N_10203,N_9371,N_9239);
and U10204 (N_10204,N_9689,N_9786);
xnor U10205 (N_10205,N_9973,N_9390);
and U10206 (N_10206,N_9231,N_9669);
xnor U10207 (N_10207,N_9392,N_9878);
nand U10208 (N_10208,N_9486,N_9229);
nand U10209 (N_10209,N_9980,N_9746);
xnor U10210 (N_10210,N_9006,N_9733);
and U10211 (N_10211,N_9587,N_9164);
and U10212 (N_10212,N_9073,N_9341);
or U10213 (N_10213,N_9340,N_9787);
nand U10214 (N_10214,N_9683,N_9568);
or U10215 (N_10215,N_9531,N_9540);
nor U10216 (N_10216,N_9422,N_9289);
xor U10217 (N_10217,N_9475,N_9312);
nor U10218 (N_10218,N_9268,N_9534);
nor U10219 (N_10219,N_9260,N_9725);
xnor U10220 (N_10220,N_9583,N_9227);
nand U10221 (N_10221,N_9483,N_9088);
nor U10222 (N_10222,N_9472,N_9053);
xnor U10223 (N_10223,N_9136,N_9914);
nor U10224 (N_10224,N_9172,N_9966);
or U10225 (N_10225,N_9324,N_9057);
nand U10226 (N_10226,N_9142,N_9398);
or U10227 (N_10227,N_9620,N_9982);
or U10228 (N_10228,N_9184,N_9311);
nor U10229 (N_10229,N_9285,N_9480);
nor U10230 (N_10230,N_9723,N_9354);
xor U10231 (N_10231,N_9532,N_9470);
and U10232 (N_10232,N_9571,N_9122);
nand U10233 (N_10233,N_9660,N_9708);
nor U10234 (N_10234,N_9522,N_9203);
nor U10235 (N_10235,N_9457,N_9854);
xor U10236 (N_10236,N_9448,N_9662);
and U10237 (N_10237,N_9366,N_9594);
and U10238 (N_10238,N_9589,N_9440);
nand U10239 (N_10239,N_9145,N_9282);
xor U10240 (N_10240,N_9842,N_9947);
nor U10241 (N_10241,N_9299,N_9045);
nand U10242 (N_10242,N_9363,N_9058);
and U10243 (N_10243,N_9800,N_9040);
and U10244 (N_10244,N_9737,N_9429);
nor U10245 (N_10245,N_9671,N_9759);
nor U10246 (N_10246,N_9024,N_9270);
or U10247 (N_10247,N_9699,N_9432);
and U10248 (N_10248,N_9789,N_9538);
nor U10249 (N_10249,N_9705,N_9768);
nand U10250 (N_10250,N_9405,N_9137);
nor U10251 (N_10251,N_9678,N_9188);
xnor U10252 (N_10252,N_9202,N_9455);
and U10253 (N_10253,N_9749,N_9895);
xnor U10254 (N_10254,N_9012,N_9066);
xnor U10255 (N_10255,N_9076,N_9092);
nor U10256 (N_10256,N_9317,N_9833);
or U10257 (N_10257,N_9086,N_9452);
nor U10258 (N_10258,N_9033,N_9360);
and U10259 (N_10259,N_9286,N_9302);
xnor U10260 (N_10260,N_9714,N_9765);
nand U10261 (N_10261,N_9893,N_9940);
nor U10262 (N_10262,N_9177,N_9794);
nand U10263 (N_10263,N_9062,N_9183);
nand U10264 (N_10264,N_9272,N_9111);
or U10265 (N_10265,N_9080,N_9911);
xnor U10266 (N_10266,N_9265,N_9625);
and U10267 (N_10267,N_9606,N_9537);
or U10268 (N_10268,N_9461,N_9784);
nand U10269 (N_10269,N_9449,N_9495);
or U10270 (N_10270,N_9682,N_9016);
and U10271 (N_10271,N_9105,N_9474);
nor U10272 (N_10272,N_9152,N_9834);
or U10273 (N_10273,N_9315,N_9218);
and U10274 (N_10274,N_9162,N_9010);
or U10275 (N_10275,N_9929,N_9482);
nor U10276 (N_10276,N_9856,N_9802);
nand U10277 (N_10277,N_9898,N_9464);
nand U10278 (N_10278,N_9124,N_9370);
and U10279 (N_10279,N_9774,N_9029);
or U10280 (N_10280,N_9403,N_9862);
nand U10281 (N_10281,N_9020,N_9135);
nor U10282 (N_10282,N_9300,N_9822);
and U10283 (N_10283,N_9427,N_9666);
and U10284 (N_10284,N_9685,N_9054);
or U10285 (N_10285,N_9352,N_9471);
and U10286 (N_10286,N_9981,N_9394);
nor U10287 (N_10287,N_9189,N_9085);
and U10288 (N_10288,N_9185,N_9228);
nor U10289 (N_10289,N_9558,N_9650);
xnor U10290 (N_10290,N_9087,N_9613);
and U10291 (N_10291,N_9902,N_9015);
nor U10292 (N_10292,N_9543,N_9348);
nor U10293 (N_10293,N_9175,N_9506);
and U10294 (N_10294,N_9935,N_9663);
or U10295 (N_10295,N_9824,N_9805);
nor U10296 (N_10296,N_9060,N_9890);
nor U10297 (N_10297,N_9910,N_9577);
nand U10298 (N_10298,N_9430,N_9949);
nor U10299 (N_10299,N_9437,N_9888);
and U10300 (N_10300,N_9065,N_9083);
or U10301 (N_10301,N_9106,N_9851);
nor U10302 (N_10302,N_9072,N_9629);
nand U10303 (N_10303,N_9091,N_9372);
nor U10304 (N_10304,N_9853,N_9816);
and U10305 (N_10305,N_9008,N_9165);
nor U10306 (N_10306,N_9242,N_9365);
xor U10307 (N_10307,N_9941,N_9113);
and U10308 (N_10308,N_9089,N_9590);
and U10309 (N_10309,N_9956,N_9861);
and U10310 (N_10310,N_9232,N_9887);
or U10311 (N_10311,N_9582,N_9803);
nor U10312 (N_10312,N_9527,N_9336);
or U10313 (N_10313,N_9438,N_9847);
and U10314 (N_10314,N_9528,N_9444);
nand U10315 (N_10315,N_9052,N_9892);
and U10316 (N_10316,N_9918,N_9525);
nand U10317 (N_10317,N_9463,N_9741);
nor U10318 (N_10318,N_9955,N_9549);
or U10319 (N_10319,N_9667,N_9831);
and U10320 (N_10320,N_9601,N_9244);
and U10321 (N_10321,N_9041,N_9726);
nand U10322 (N_10322,N_9533,N_9153);
or U10323 (N_10323,N_9385,N_9451);
nand U10324 (N_10324,N_9627,N_9345);
xnor U10325 (N_10325,N_9753,N_9277);
or U10326 (N_10326,N_9168,N_9642);
nand U10327 (N_10327,N_9875,N_9155);
or U10328 (N_10328,N_9292,N_9179);
or U10329 (N_10329,N_9031,N_9257);
and U10330 (N_10330,N_9418,N_9600);
or U10331 (N_10331,N_9479,N_9119);
nand U10332 (N_10332,N_9027,N_9958);
and U10333 (N_10333,N_9499,N_9772);
or U10334 (N_10334,N_9564,N_9840);
and U10335 (N_10335,N_9306,N_9063);
nor U10336 (N_10336,N_9879,N_9905);
nand U10337 (N_10337,N_9942,N_9659);
and U10338 (N_10338,N_9380,N_9945);
nor U10339 (N_10339,N_9869,N_9965);
or U10340 (N_10340,N_9230,N_9508);
and U10341 (N_10341,N_9755,N_9381);
nor U10342 (N_10342,N_9792,N_9611);
nor U10343 (N_10343,N_9280,N_9618);
xor U10344 (N_10344,N_9655,N_9736);
nor U10345 (N_10345,N_9256,N_9138);
or U10346 (N_10346,N_9382,N_9688);
or U10347 (N_10347,N_9706,N_9812);
nor U10348 (N_10348,N_9255,N_9477);
nand U10349 (N_10349,N_9707,N_9975);
xor U10350 (N_10350,N_9443,N_9885);
or U10351 (N_10351,N_9919,N_9536);
nand U10352 (N_10352,N_9262,N_9837);
and U10353 (N_10353,N_9017,N_9004);
and U10354 (N_10354,N_9247,N_9358);
nor U10355 (N_10355,N_9069,N_9624);
xnor U10356 (N_10356,N_9849,N_9036);
or U10357 (N_10357,N_9281,N_9476);
and U10358 (N_10358,N_9716,N_9278);
nand U10359 (N_10359,N_9928,N_9807);
nor U10360 (N_10360,N_9368,N_9226);
xor U10361 (N_10361,N_9301,N_9829);
nor U10362 (N_10362,N_9093,N_9346);
and U10363 (N_10363,N_9976,N_9821);
and U10364 (N_10364,N_9364,N_9068);
xor U10365 (N_10365,N_9290,N_9811);
nor U10366 (N_10366,N_9279,N_9099);
and U10367 (N_10367,N_9241,N_9407);
and U10368 (N_10368,N_9649,N_9567);
nor U10369 (N_10369,N_9563,N_9889);
or U10370 (N_10370,N_9114,N_9216);
nor U10371 (N_10371,N_9067,N_9320);
nor U10372 (N_10372,N_9078,N_9018);
and U10373 (N_10373,N_9173,N_9096);
and U10374 (N_10374,N_9948,N_9825);
or U10375 (N_10375,N_9638,N_9703);
and U10376 (N_10376,N_9223,N_9294);
or U10377 (N_10377,N_9727,N_9554);
nand U10378 (N_10378,N_9331,N_9133);
xor U10379 (N_10379,N_9194,N_9904);
nor U10380 (N_10380,N_9131,N_9107);
xor U10381 (N_10381,N_9361,N_9857);
nor U10382 (N_10382,N_9249,N_9748);
xnor U10383 (N_10383,N_9695,N_9329);
or U10384 (N_10384,N_9684,N_9404);
nand U10385 (N_10385,N_9717,N_9991);
xnor U10386 (N_10386,N_9841,N_9874);
and U10387 (N_10387,N_9916,N_9254);
nand U10388 (N_10388,N_9005,N_9209);
and U10389 (N_10389,N_9738,N_9742);
and U10390 (N_10390,N_9830,N_9535);
or U10391 (N_10391,N_9081,N_9410);
nor U10392 (N_10392,N_9201,N_9337);
nand U10393 (N_10393,N_9198,N_9681);
and U10394 (N_10394,N_9071,N_9442);
or U10395 (N_10395,N_9635,N_9526);
or U10396 (N_10396,N_9413,N_9623);
or U10397 (N_10397,N_9728,N_9284);
or U10398 (N_10398,N_9204,N_9632);
nand U10399 (N_10399,N_9751,N_9061);
or U10400 (N_10400,N_9839,N_9963);
xnor U10401 (N_10401,N_9343,N_9621);
or U10402 (N_10402,N_9023,N_9961);
nor U10403 (N_10403,N_9924,N_9077);
nand U10404 (N_10404,N_9221,N_9174);
nor U10405 (N_10405,N_9775,N_9504);
and U10406 (N_10406,N_9521,N_9871);
nor U10407 (N_10407,N_9700,N_9182);
and U10408 (N_10408,N_9901,N_9813);
nor U10409 (N_10409,N_9001,N_9149);
xnor U10410 (N_10410,N_9672,N_9636);
nor U10411 (N_10411,N_9180,N_9514);
nor U10412 (N_10412,N_9634,N_9545);
nor U10413 (N_10413,N_9460,N_9820);
nand U10414 (N_10414,N_9000,N_9421);
nand U10415 (N_10415,N_9610,N_9909);
nand U10416 (N_10416,N_9176,N_9855);
and U10417 (N_10417,N_9097,N_9996);
and U10418 (N_10418,N_9576,N_9934);
nor U10419 (N_10419,N_9520,N_9043);
and U10420 (N_10420,N_9139,N_9428);
and U10421 (N_10421,N_9200,N_9517);
nor U10422 (N_10422,N_9766,N_9994);
or U10423 (N_10423,N_9500,N_9258);
or U10424 (N_10424,N_9102,N_9651);
xnor U10425 (N_10425,N_9322,N_9261);
nand U10426 (N_10426,N_9388,N_9196);
xor U10427 (N_10427,N_9823,N_9586);
and U10428 (N_10428,N_9416,N_9140);
nand U10429 (N_10429,N_9383,N_9546);
nor U10430 (N_10430,N_9964,N_9896);
xor U10431 (N_10431,N_9927,N_9801);
nand U10432 (N_10432,N_9347,N_9050);
and U10433 (N_10433,N_9605,N_9992);
nor U10434 (N_10434,N_9595,N_9709);
nand U10435 (N_10435,N_9574,N_9288);
and U10436 (N_10436,N_9957,N_9648);
nor U10437 (N_10437,N_9082,N_9453);
or U10438 (N_10438,N_9397,N_9305);
nor U10439 (N_10439,N_9509,N_9931);
or U10440 (N_10440,N_9357,N_9489);
nor U10441 (N_10441,N_9886,N_9263);
or U10442 (N_10442,N_9362,N_9720);
nand U10443 (N_10443,N_9858,N_9344);
nor U10444 (N_10444,N_9970,N_9399);
xnor U10445 (N_10445,N_9234,N_9569);
and U10446 (N_10446,N_9880,N_9026);
nor U10447 (N_10447,N_9760,N_9770);
nor U10448 (N_10448,N_9835,N_9580);
or U10449 (N_10449,N_9997,N_9883);
or U10450 (N_10450,N_9297,N_9376);
and U10451 (N_10451,N_9915,N_9309);
nor U10452 (N_10452,N_9121,N_9724);
and U10453 (N_10453,N_9579,N_9926);
nand U10454 (N_10454,N_9756,N_9771);
or U10455 (N_10455,N_9646,N_9561);
nor U10456 (N_10456,N_9129,N_9676);
or U10457 (N_10457,N_9864,N_9722);
or U10458 (N_10458,N_9985,N_9719);
xor U10459 (N_10459,N_9596,N_9882);
nor U10460 (N_10460,N_9602,N_9491);
nand U10461 (N_10461,N_9848,N_9387);
and U10462 (N_10462,N_9051,N_9818);
or U10463 (N_10463,N_9806,N_9485);
and U10464 (N_10464,N_9025,N_9384);
or U10465 (N_10465,N_9314,N_9758);
nand U10466 (N_10466,N_9865,N_9190);
or U10467 (N_10467,N_9993,N_9922);
nand U10468 (N_10468,N_9622,N_9815);
or U10469 (N_10469,N_9588,N_9490);
or U10470 (N_10470,N_9990,N_9950);
nor U10471 (N_10471,N_9585,N_9274);
or U10472 (N_10472,N_9426,N_9507);
and U10473 (N_10473,N_9158,N_9207);
xor U10474 (N_10474,N_9906,N_9014);
and U10475 (N_10475,N_9967,N_9852);
nand U10476 (N_10476,N_9664,N_9779);
and U10477 (N_10477,N_9978,N_9369);
or U10478 (N_10478,N_9592,N_9987);
or U10479 (N_10479,N_9808,N_9468);
or U10480 (N_10480,N_9120,N_9002);
and U10481 (N_10481,N_9687,N_9572);
nand U10482 (N_10482,N_9431,N_9776);
nand U10483 (N_10483,N_9224,N_9584);
nand U10484 (N_10484,N_9123,N_9497);
or U10485 (N_10485,N_9647,N_9205);
nor U10486 (N_10486,N_9908,N_9146);
nor U10487 (N_10487,N_9995,N_9253);
nor U10488 (N_10488,N_9850,N_9819);
nand U10489 (N_10489,N_9503,N_9328);
or U10490 (N_10490,N_9195,N_9866);
nor U10491 (N_10491,N_9628,N_9434);
or U10492 (N_10492,N_9690,N_9732);
and U10493 (N_10493,N_9330,N_9515);
nor U10494 (N_10494,N_9989,N_9696);
or U10495 (N_10495,N_9846,N_9424);
nor U10496 (N_10496,N_9264,N_9339);
or U10497 (N_10497,N_9252,N_9425);
xnor U10498 (N_10498,N_9559,N_9679);
and U10499 (N_10499,N_9356,N_9147);
or U10500 (N_10500,N_9310,N_9188);
nor U10501 (N_10501,N_9211,N_9076);
nor U10502 (N_10502,N_9836,N_9411);
nor U10503 (N_10503,N_9167,N_9229);
nor U10504 (N_10504,N_9459,N_9811);
and U10505 (N_10505,N_9891,N_9968);
or U10506 (N_10506,N_9615,N_9014);
or U10507 (N_10507,N_9363,N_9706);
xnor U10508 (N_10508,N_9223,N_9322);
nand U10509 (N_10509,N_9398,N_9405);
and U10510 (N_10510,N_9012,N_9227);
and U10511 (N_10511,N_9919,N_9352);
xnor U10512 (N_10512,N_9117,N_9197);
or U10513 (N_10513,N_9801,N_9321);
nand U10514 (N_10514,N_9424,N_9097);
nand U10515 (N_10515,N_9903,N_9745);
and U10516 (N_10516,N_9920,N_9199);
nand U10517 (N_10517,N_9749,N_9161);
or U10518 (N_10518,N_9472,N_9132);
and U10519 (N_10519,N_9707,N_9886);
or U10520 (N_10520,N_9456,N_9024);
and U10521 (N_10521,N_9968,N_9924);
nor U10522 (N_10522,N_9555,N_9996);
and U10523 (N_10523,N_9714,N_9375);
nor U10524 (N_10524,N_9494,N_9044);
nor U10525 (N_10525,N_9639,N_9354);
and U10526 (N_10526,N_9137,N_9191);
nand U10527 (N_10527,N_9998,N_9576);
or U10528 (N_10528,N_9748,N_9931);
and U10529 (N_10529,N_9201,N_9907);
and U10530 (N_10530,N_9955,N_9489);
xnor U10531 (N_10531,N_9195,N_9068);
nor U10532 (N_10532,N_9873,N_9101);
or U10533 (N_10533,N_9827,N_9561);
nand U10534 (N_10534,N_9361,N_9602);
or U10535 (N_10535,N_9842,N_9629);
nor U10536 (N_10536,N_9016,N_9012);
nor U10537 (N_10537,N_9433,N_9986);
xor U10538 (N_10538,N_9426,N_9029);
nand U10539 (N_10539,N_9626,N_9440);
nor U10540 (N_10540,N_9509,N_9787);
and U10541 (N_10541,N_9155,N_9698);
or U10542 (N_10542,N_9235,N_9811);
xor U10543 (N_10543,N_9201,N_9133);
nor U10544 (N_10544,N_9944,N_9718);
nand U10545 (N_10545,N_9401,N_9136);
or U10546 (N_10546,N_9094,N_9078);
nor U10547 (N_10547,N_9970,N_9435);
and U10548 (N_10548,N_9040,N_9638);
xor U10549 (N_10549,N_9601,N_9421);
nand U10550 (N_10550,N_9349,N_9961);
and U10551 (N_10551,N_9538,N_9173);
nand U10552 (N_10552,N_9695,N_9983);
and U10553 (N_10553,N_9925,N_9591);
or U10554 (N_10554,N_9861,N_9705);
nand U10555 (N_10555,N_9248,N_9615);
nand U10556 (N_10556,N_9681,N_9090);
and U10557 (N_10557,N_9018,N_9231);
nor U10558 (N_10558,N_9370,N_9831);
nand U10559 (N_10559,N_9816,N_9286);
nand U10560 (N_10560,N_9446,N_9058);
or U10561 (N_10561,N_9515,N_9626);
nor U10562 (N_10562,N_9007,N_9086);
or U10563 (N_10563,N_9007,N_9735);
nor U10564 (N_10564,N_9165,N_9245);
xor U10565 (N_10565,N_9898,N_9475);
and U10566 (N_10566,N_9504,N_9118);
or U10567 (N_10567,N_9363,N_9777);
nand U10568 (N_10568,N_9683,N_9671);
nand U10569 (N_10569,N_9385,N_9212);
and U10570 (N_10570,N_9836,N_9817);
nor U10571 (N_10571,N_9398,N_9726);
xor U10572 (N_10572,N_9503,N_9109);
and U10573 (N_10573,N_9711,N_9118);
nor U10574 (N_10574,N_9055,N_9330);
xnor U10575 (N_10575,N_9462,N_9488);
nand U10576 (N_10576,N_9852,N_9020);
xor U10577 (N_10577,N_9915,N_9287);
or U10578 (N_10578,N_9421,N_9286);
and U10579 (N_10579,N_9182,N_9495);
nand U10580 (N_10580,N_9839,N_9391);
nor U10581 (N_10581,N_9653,N_9385);
nor U10582 (N_10582,N_9862,N_9782);
or U10583 (N_10583,N_9703,N_9579);
or U10584 (N_10584,N_9257,N_9006);
nor U10585 (N_10585,N_9753,N_9703);
xnor U10586 (N_10586,N_9993,N_9771);
and U10587 (N_10587,N_9997,N_9387);
and U10588 (N_10588,N_9161,N_9352);
xnor U10589 (N_10589,N_9970,N_9394);
xnor U10590 (N_10590,N_9112,N_9623);
or U10591 (N_10591,N_9268,N_9381);
and U10592 (N_10592,N_9012,N_9361);
xnor U10593 (N_10593,N_9287,N_9439);
nor U10594 (N_10594,N_9715,N_9553);
xor U10595 (N_10595,N_9386,N_9187);
nand U10596 (N_10596,N_9411,N_9459);
and U10597 (N_10597,N_9203,N_9979);
nor U10598 (N_10598,N_9981,N_9581);
nor U10599 (N_10599,N_9241,N_9849);
and U10600 (N_10600,N_9628,N_9732);
nor U10601 (N_10601,N_9609,N_9745);
nor U10602 (N_10602,N_9761,N_9970);
nor U10603 (N_10603,N_9975,N_9521);
nand U10604 (N_10604,N_9376,N_9474);
and U10605 (N_10605,N_9261,N_9675);
nor U10606 (N_10606,N_9539,N_9303);
nand U10607 (N_10607,N_9956,N_9836);
nand U10608 (N_10608,N_9505,N_9541);
or U10609 (N_10609,N_9978,N_9667);
nand U10610 (N_10610,N_9862,N_9519);
xor U10611 (N_10611,N_9397,N_9577);
xor U10612 (N_10612,N_9964,N_9125);
nand U10613 (N_10613,N_9928,N_9788);
nand U10614 (N_10614,N_9707,N_9173);
xor U10615 (N_10615,N_9058,N_9624);
and U10616 (N_10616,N_9797,N_9075);
and U10617 (N_10617,N_9439,N_9482);
or U10618 (N_10618,N_9040,N_9653);
nor U10619 (N_10619,N_9219,N_9544);
and U10620 (N_10620,N_9318,N_9916);
nor U10621 (N_10621,N_9920,N_9135);
and U10622 (N_10622,N_9894,N_9210);
nor U10623 (N_10623,N_9631,N_9304);
xnor U10624 (N_10624,N_9928,N_9256);
nor U10625 (N_10625,N_9988,N_9552);
or U10626 (N_10626,N_9383,N_9496);
nand U10627 (N_10627,N_9522,N_9598);
nand U10628 (N_10628,N_9338,N_9885);
nor U10629 (N_10629,N_9396,N_9696);
nand U10630 (N_10630,N_9997,N_9901);
nand U10631 (N_10631,N_9407,N_9826);
nand U10632 (N_10632,N_9024,N_9023);
or U10633 (N_10633,N_9469,N_9551);
xnor U10634 (N_10634,N_9798,N_9117);
and U10635 (N_10635,N_9133,N_9167);
nand U10636 (N_10636,N_9194,N_9628);
nor U10637 (N_10637,N_9122,N_9568);
nand U10638 (N_10638,N_9958,N_9450);
and U10639 (N_10639,N_9340,N_9360);
nor U10640 (N_10640,N_9473,N_9340);
nand U10641 (N_10641,N_9142,N_9290);
nor U10642 (N_10642,N_9783,N_9033);
or U10643 (N_10643,N_9723,N_9789);
and U10644 (N_10644,N_9656,N_9690);
and U10645 (N_10645,N_9516,N_9563);
nand U10646 (N_10646,N_9839,N_9456);
nor U10647 (N_10647,N_9607,N_9753);
and U10648 (N_10648,N_9110,N_9876);
nor U10649 (N_10649,N_9077,N_9519);
nor U10650 (N_10650,N_9563,N_9122);
or U10651 (N_10651,N_9005,N_9474);
and U10652 (N_10652,N_9921,N_9312);
or U10653 (N_10653,N_9722,N_9034);
nand U10654 (N_10654,N_9380,N_9864);
and U10655 (N_10655,N_9175,N_9052);
and U10656 (N_10656,N_9776,N_9063);
nand U10657 (N_10657,N_9655,N_9871);
nor U10658 (N_10658,N_9315,N_9553);
nor U10659 (N_10659,N_9660,N_9826);
or U10660 (N_10660,N_9517,N_9041);
nor U10661 (N_10661,N_9654,N_9458);
nand U10662 (N_10662,N_9792,N_9359);
and U10663 (N_10663,N_9951,N_9823);
nand U10664 (N_10664,N_9721,N_9093);
nand U10665 (N_10665,N_9608,N_9132);
or U10666 (N_10666,N_9874,N_9455);
and U10667 (N_10667,N_9581,N_9254);
or U10668 (N_10668,N_9102,N_9762);
nor U10669 (N_10669,N_9226,N_9466);
or U10670 (N_10670,N_9886,N_9968);
nor U10671 (N_10671,N_9703,N_9310);
nor U10672 (N_10672,N_9590,N_9633);
nor U10673 (N_10673,N_9747,N_9647);
or U10674 (N_10674,N_9227,N_9939);
or U10675 (N_10675,N_9064,N_9317);
and U10676 (N_10676,N_9665,N_9582);
nand U10677 (N_10677,N_9166,N_9322);
or U10678 (N_10678,N_9331,N_9164);
nand U10679 (N_10679,N_9019,N_9214);
nand U10680 (N_10680,N_9808,N_9343);
nand U10681 (N_10681,N_9306,N_9932);
or U10682 (N_10682,N_9852,N_9891);
nor U10683 (N_10683,N_9255,N_9783);
or U10684 (N_10684,N_9771,N_9403);
xnor U10685 (N_10685,N_9216,N_9294);
or U10686 (N_10686,N_9637,N_9409);
and U10687 (N_10687,N_9308,N_9387);
and U10688 (N_10688,N_9584,N_9435);
nand U10689 (N_10689,N_9918,N_9998);
and U10690 (N_10690,N_9296,N_9271);
nand U10691 (N_10691,N_9145,N_9004);
or U10692 (N_10692,N_9577,N_9153);
or U10693 (N_10693,N_9225,N_9470);
nand U10694 (N_10694,N_9742,N_9941);
nand U10695 (N_10695,N_9562,N_9986);
nor U10696 (N_10696,N_9015,N_9385);
and U10697 (N_10697,N_9811,N_9645);
and U10698 (N_10698,N_9198,N_9824);
nor U10699 (N_10699,N_9548,N_9466);
nor U10700 (N_10700,N_9184,N_9934);
nor U10701 (N_10701,N_9159,N_9090);
nor U10702 (N_10702,N_9598,N_9660);
nand U10703 (N_10703,N_9196,N_9888);
nor U10704 (N_10704,N_9250,N_9397);
and U10705 (N_10705,N_9160,N_9247);
nand U10706 (N_10706,N_9992,N_9545);
and U10707 (N_10707,N_9845,N_9695);
nand U10708 (N_10708,N_9773,N_9367);
nor U10709 (N_10709,N_9074,N_9004);
nor U10710 (N_10710,N_9216,N_9187);
and U10711 (N_10711,N_9259,N_9214);
nand U10712 (N_10712,N_9174,N_9973);
nor U10713 (N_10713,N_9362,N_9456);
or U10714 (N_10714,N_9107,N_9308);
nor U10715 (N_10715,N_9740,N_9728);
nand U10716 (N_10716,N_9258,N_9900);
nor U10717 (N_10717,N_9572,N_9816);
or U10718 (N_10718,N_9141,N_9320);
nand U10719 (N_10719,N_9305,N_9615);
or U10720 (N_10720,N_9348,N_9023);
and U10721 (N_10721,N_9661,N_9536);
nor U10722 (N_10722,N_9662,N_9257);
or U10723 (N_10723,N_9369,N_9296);
or U10724 (N_10724,N_9994,N_9938);
or U10725 (N_10725,N_9819,N_9051);
and U10726 (N_10726,N_9022,N_9838);
and U10727 (N_10727,N_9044,N_9050);
nand U10728 (N_10728,N_9969,N_9788);
nor U10729 (N_10729,N_9413,N_9078);
and U10730 (N_10730,N_9174,N_9663);
xnor U10731 (N_10731,N_9382,N_9822);
nor U10732 (N_10732,N_9379,N_9697);
or U10733 (N_10733,N_9480,N_9556);
nor U10734 (N_10734,N_9353,N_9178);
or U10735 (N_10735,N_9081,N_9764);
and U10736 (N_10736,N_9773,N_9713);
nand U10737 (N_10737,N_9537,N_9950);
nor U10738 (N_10738,N_9594,N_9874);
xnor U10739 (N_10739,N_9839,N_9820);
or U10740 (N_10740,N_9168,N_9788);
and U10741 (N_10741,N_9270,N_9020);
nor U10742 (N_10742,N_9698,N_9090);
or U10743 (N_10743,N_9219,N_9568);
nor U10744 (N_10744,N_9222,N_9965);
and U10745 (N_10745,N_9401,N_9931);
nand U10746 (N_10746,N_9320,N_9485);
xnor U10747 (N_10747,N_9242,N_9199);
xor U10748 (N_10748,N_9730,N_9247);
nand U10749 (N_10749,N_9460,N_9322);
nand U10750 (N_10750,N_9847,N_9136);
nand U10751 (N_10751,N_9446,N_9410);
and U10752 (N_10752,N_9465,N_9029);
or U10753 (N_10753,N_9038,N_9612);
nand U10754 (N_10754,N_9827,N_9792);
and U10755 (N_10755,N_9185,N_9232);
nand U10756 (N_10756,N_9827,N_9972);
and U10757 (N_10757,N_9945,N_9669);
or U10758 (N_10758,N_9159,N_9844);
nor U10759 (N_10759,N_9236,N_9645);
and U10760 (N_10760,N_9253,N_9406);
and U10761 (N_10761,N_9824,N_9407);
nand U10762 (N_10762,N_9562,N_9201);
nand U10763 (N_10763,N_9243,N_9347);
and U10764 (N_10764,N_9221,N_9150);
or U10765 (N_10765,N_9453,N_9174);
nor U10766 (N_10766,N_9041,N_9845);
nand U10767 (N_10767,N_9260,N_9198);
nand U10768 (N_10768,N_9590,N_9302);
xnor U10769 (N_10769,N_9205,N_9514);
or U10770 (N_10770,N_9528,N_9076);
nor U10771 (N_10771,N_9626,N_9600);
and U10772 (N_10772,N_9257,N_9647);
nand U10773 (N_10773,N_9272,N_9491);
or U10774 (N_10774,N_9045,N_9487);
and U10775 (N_10775,N_9280,N_9818);
xnor U10776 (N_10776,N_9785,N_9712);
nand U10777 (N_10777,N_9177,N_9750);
nor U10778 (N_10778,N_9493,N_9472);
or U10779 (N_10779,N_9984,N_9274);
nor U10780 (N_10780,N_9186,N_9923);
xor U10781 (N_10781,N_9818,N_9829);
or U10782 (N_10782,N_9375,N_9518);
nor U10783 (N_10783,N_9494,N_9030);
xor U10784 (N_10784,N_9495,N_9530);
or U10785 (N_10785,N_9556,N_9450);
nor U10786 (N_10786,N_9450,N_9357);
nand U10787 (N_10787,N_9773,N_9458);
or U10788 (N_10788,N_9556,N_9998);
and U10789 (N_10789,N_9843,N_9288);
xor U10790 (N_10790,N_9149,N_9458);
nor U10791 (N_10791,N_9491,N_9189);
and U10792 (N_10792,N_9061,N_9797);
nor U10793 (N_10793,N_9403,N_9173);
nand U10794 (N_10794,N_9767,N_9463);
or U10795 (N_10795,N_9489,N_9021);
nor U10796 (N_10796,N_9803,N_9445);
nand U10797 (N_10797,N_9172,N_9561);
and U10798 (N_10798,N_9123,N_9546);
nor U10799 (N_10799,N_9026,N_9421);
and U10800 (N_10800,N_9860,N_9151);
and U10801 (N_10801,N_9858,N_9918);
nand U10802 (N_10802,N_9337,N_9663);
and U10803 (N_10803,N_9835,N_9476);
or U10804 (N_10804,N_9543,N_9626);
and U10805 (N_10805,N_9561,N_9505);
xor U10806 (N_10806,N_9369,N_9706);
nor U10807 (N_10807,N_9614,N_9345);
nand U10808 (N_10808,N_9318,N_9913);
nor U10809 (N_10809,N_9683,N_9624);
or U10810 (N_10810,N_9807,N_9234);
nor U10811 (N_10811,N_9212,N_9900);
nor U10812 (N_10812,N_9542,N_9509);
nand U10813 (N_10813,N_9386,N_9368);
nand U10814 (N_10814,N_9539,N_9452);
xor U10815 (N_10815,N_9758,N_9716);
nor U10816 (N_10816,N_9868,N_9577);
or U10817 (N_10817,N_9624,N_9040);
nor U10818 (N_10818,N_9065,N_9511);
nor U10819 (N_10819,N_9137,N_9270);
nand U10820 (N_10820,N_9060,N_9732);
or U10821 (N_10821,N_9807,N_9108);
nor U10822 (N_10822,N_9665,N_9378);
nand U10823 (N_10823,N_9010,N_9392);
or U10824 (N_10824,N_9449,N_9058);
nor U10825 (N_10825,N_9321,N_9223);
or U10826 (N_10826,N_9923,N_9664);
and U10827 (N_10827,N_9846,N_9845);
and U10828 (N_10828,N_9434,N_9503);
nand U10829 (N_10829,N_9487,N_9292);
nand U10830 (N_10830,N_9847,N_9992);
or U10831 (N_10831,N_9585,N_9281);
nor U10832 (N_10832,N_9519,N_9633);
xor U10833 (N_10833,N_9579,N_9702);
and U10834 (N_10834,N_9655,N_9223);
nand U10835 (N_10835,N_9826,N_9715);
nor U10836 (N_10836,N_9008,N_9152);
nand U10837 (N_10837,N_9201,N_9667);
and U10838 (N_10838,N_9570,N_9020);
or U10839 (N_10839,N_9967,N_9562);
nor U10840 (N_10840,N_9286,N_9071);
and U10841 (N_10841,N_9670,N_9347);
or U10842 (N_10842,N_9991,N_9060);
or U10843 (N_10843,N_9777,N_9035);
xor U10844 (N_10844,N_9800,N_9075);
or U10845 (N_10845,N_9552,N_9775);
and U10846 (N_10846,N_9997,N_9675);
and U10847 (N_10847,N_9891,N_9143);
xnor U10848 (N_10848,N_9660,N_9222);
xnor U10849 (N_10849,N_9554,N_9573);
and U10850 (N_10850,N_9118,N_9221);
and U10851 (N_10851,N_9957,N_9046);
xor U10852 (N_10852,N_9666,N_9388);
or U10853 (N_10853,N_9150,N_9999);
or U10854 (N_10854,N_9718,N_9070);
nand U10855 (N_10855,N_9063,N_9877);
nor U10856 (N_10856,N_9108,N_9131);
or U10857 (N_10857,N_9777,N_9454);
nand U10858 (N_10858,N_9563,N_9912);
nor U10859 (N_10859,N_9001,N_9124);
nand U10860 (N_10860,N_9279,N_9063);
and U10861 (N_10861,N_9064,N_9124);
xor U10862 (N_10862,N_9612,N_9566);
xor U10863 (N_10863,N_9530,N_9448);
and U10864 (N_10864,N_9107,N_9820);
nor U10865 (N_10865,N_9572,N_9856);
xor U10866 (N_10866,N_9101,N_9046);
and U10867 (N_10867,N_9662,N_9721);
nor U10868 (N_10868,N_9171,N_9259);
nand U10869 (N_10869,N_9125,N_9585);
or U10870 (N_10870,N_9072,N_9100);
and U10871 (N_10871,N_9500,N_9299);
xnor U10872 (N_10872,N_9556,N_9821);
or U10873 (N_10873,N_9709,N_9312);
nor U10874 (N_10874,N_9706,N_9320);
nor U10875 (N_10875,N_9786,N_9620);
and U10876 (N_10876,N_9354,N_9442);
and U10877 (N_10877,N_9586,N_9420);
and U10878 (N_10878,N_9648,N_9971);
xnor U10879 (N_10879,N_9160,N_9488);
or U10880 (N_10880,N_9805,N_9077);
nand U10881 (N_10881,N_9560,N_9686);
or U10882 (N_10882,N_9663,N_9451);
nand U10883 (N_10883,N_9751,N_9515);
nand U10884 (N_10884,N_9319,N_9784);
nor U10885 (N_10885,N_9079,N_9798);
nand U10886 (N_10886,N_9626,N_9246);
or U10887 (N_10887,N_9647,N_9849);
and U10888 (N_10888,N_9245,N_9714);
nor U10889 (N_10889,N_9425,N_9304);
or U10890 (N_10890,N_9413,N_9503);
nor U10891 (N_10891,N_9701,N_9020);
or U10892 (N_10892,N_9803,N_9748);
or U10893 (N_10893,N_9488,N_9143);
and U10894 (N_10894,N_9734,N_9634);
xnor U10895 (N_10895,N_9604,N_9945);
nor U10896 (N_10896,N_9572,N_9756);
nor U10897 (N_10897,N_9114,N_9253);
nor U10898 (N_10898,N_9387,N_9980);
and U10899 (N_10899,N_9940,N_9672);
nand U10900 (N_10900,N_9215,N_9761);
or U10901 (N_10901,N_9737,N_9757);
nor U10902 (N_10902,N_9794,N_9394);
or U10903 (N_10903,N_9695,N_9612);
and U10904 (N_10904,N_9785,N_9657);
nor U10905 (N_10905,N_9247,N_9086);
nand U10906 (N_10906,N_9773,N_9959);
and U10907 (N_10907,N_9377,N_9561);
or U10908 (N_10908,N_9335,N_9194);
nor U10909 (N_10909,N_9164,N_9514);
nand U10910 (N_10910,N_9349,N_9330);
nor U10911 (N_10911,N_9788,N_9841);
or U10912 (N_10912,N_9927,N_9073);
nand U10913 (N_10913,N_9885,N_9606);
and U10914 (N_10914,N_9596,N_9273);
nand U10915 (N_10915,N_9340,N_9633);
nor U10916 (N_10916,N_9978,N_9545);
nand U10917 (N_10917,N_9521,N_9409);
nor U10918 (N_10918,N_9416,N_9916);
xnor U10919 (N_10919,N_9562,N_9951);
nand U10920 (N_10920,N_9720,N_9603);
and U10921 (N_10921,N_9777,N_9599);
nand U10922 (N_10922,N_9523,N_9401);
or U10923 (N_10923,N_9818,N_9150);
or U10924 (N_10924,N_9852,N_9445);
nand U10925 (N_10925,N_9973,N_9365);
and U10926 (N_10926,N_9261,N_9719);
nor U10927 (N_10927,N_9526,N_9805);
and U10928 (N_10928,N_9973,N_9175);
nand U10929 (N_10929,N_9841,N_9991);
nand U10930 (N_10930,N_9340,N_9796);
and U10931 (N_10931,N_9149,N_9131);
and U10932 (N_10932,N_9632,N_9194);
nor U10933 (N_10933,N_9807,N_9547);
or U10934 (N_10934,N_9900,N_9729);
xor U10935 (N_10935,N_9174,N_9805);
xor U10936 (N_10936,N_9561,N_9674);
nand U10937 (N_10937,N_9385,N_9002);
or U10938 (N_10938,N_9001,N_9732);
nor U10939 (N_10939,N_9112,N_9026);
nand U10940 (N_10940,N_9739,N_9024);
or U10941 (N_10941,N_9512,N_9432);
or U10942 (N_10942,N_9889,N_9430);
or U10943 (N_10943,N_9128,N_9919);
and U10944 (N_10944,N_9208,N_9289);
nand U10945 (N_10945,N_9077,N_9129);
xnor U10946 (N_10946,N_9879,N_9221);
nor U10947 (N_10947,N_9818,N_9941);
or U10948 (N_10948,N_9400,N_9964);
or U10949 (N_10949,N_9894,N_9124);
and U10950 (N_10950,N_9842,N_9482);
nor U10951 (N_10951,N_9458,N_9575);
and U10952 (N_10952,N_9229,N_9572);
nand U10953 (N_10953,N_9035,N_9393);
or U10954 (N_10954,N_9604,N_9253);
and U10955 (N_10955,N_9411,N_9804);
and U10956 (N_10956,N_9916,N_9444);
and U10957 (N_10957,N_9768,N_9683);
or U10958 (N_10958,N_9241,N_9993);
nor U10959 (N_10959,N_9115,N_9866);
nor U10960 (N_10960,N_9087,N_9376);
xor U10961 (N_10961,N_9367,N_9094);
or U10962 (N_10962,N_9969,N_9035);
and U10963 (N_10963,N_9856,N_9066);
or U10964 (N_10964,N_9781,N_9042);
nor U10965 (N_10965,N_9396,N_9014);
or U10966 (N_10966,N_9770,N_9384);
nor U10967 (N_10967,N_9316,N_9065);
nand U10968 (N_10968,N_9006,N_9073);
nor U10969 (N_10969,N_9830,N_9324);
and U10970 (N_10970,N_9384,N_9879);
and U10971 (N_10971,N_9688,N_9984);
and U10972 (N_10972,N_9405,N_9773);
nand U10973 (N_10973,N_9402,N_9416);
and U10974 (N_10974,N_9631,N_9301);
or U10975 (N_10975,N_9702,N_9465);
and U10976 (N_10976,N_9297,N_9739);
and U10977 (N_10977,N_9771,N_9849);
or U10978 (N_10978,N_9062,N_9452);
xor U10979 (N_10979,N_9284,N_9113);
or U10980 (N_10980,N_9192,N_9873);
or U10981 (N_10981,N_9144,N_9533);
and U10982 (N_10982,N_9610,N_9530);
xnor U10983 (N_10983,N_9990,N_9984);
or U10984 (N_10984,N_9520,N_9092);
and U10985 (N_10985,N_9887,N_9154);
and U10986 (N_10986,N_9281,N_9511);
nand U10987 (N_10987,N_9711,N_9248);
nor U10988 (N_10988,N_9216,N_9115);
nand U10989 (N_10989,N_9412,N_9907);
nor U10990 (N_10990,N_9346,N_9030);
or U10991 (N_10991,N_9989,N_9475);
nand U10992 (N_10992,N_9331,N_9747);
or U10993 (N_10993,N_9132,N_9553);
nor U10994 (N_10994,N_9097,N_9441);
and U10995 (N_10995,N_9012,N_9884);
nor U10996 (N_10996,N_9409,N_9690);
nand U10997 (N_10997,N_9132,N_9905);
nand U10998 (N_10998,N_9754,N_9993);
nand U10999 (N_10999,N_9837,N_9046);
nand U11000 (N_11000,N_10474,N_10125);
and U11001 (N_11001,N_10534,N_10448);
or U11002 (N_11002,N_10453,N_10146);
or U11003 (N_11003,N_10233,N_10095);
or U11004 (N_11004,N_10944,N_10622);
or U11005 (N_11005,N_10470,N_10952);
and U11006 (N_11006,N_10954,N_10787);
and U11007 (N_11007,N_10253,N_10298);
nand U11008 (N_11008,N_10627,N_10162);
or U11009 (N_11009,N_10390,N_10873);
or U11010 (N_11010,N_10172,N_10316);
and U11011 (N_11011,N_10027,N_10338);
or U11012 (N_11012,N_10708,N_10893);
xor U11013 (N_11013,N_10420,N_10018);
nand U11014 (N_11014,N_10114,N_10511);
nor U11015 (N_11015,N_10090,N_10078);
nor U11016 (N_11016,N_10762,N_10686);
xor U11017 (N_11017,N_10823,N_10718);
or U11018 (N_11018,N_10207,N_10303);
nor U11019 (N_11019,N_10309,N_10360);
and U11020 (N_11020,N_10574,N_10838);
xnor U11021 (N_11021,N_10350,N_10830);
and U11022 (N_11022,N_10806,N_10123);
nor U11023 (N_11023,N_10184,N_10737);
and U11024 (N_11024,N_10249,N_10417);
or U11025 (N_11025,N_10937,N_10908);
nand U11026 (N_11026,N_10901,N_10043);
and U11027 (N_11027,N_10799,N_10518);
nand U11028 (N_11028,N_10913,N_10914);
and U11029 (N_11029,N_10811,N_10835);
nor U11030 (N_11030,N_10365,N_10634);
nor U11031 (N_11031,N_10802,N_10803);
and U11032 (N_11032,N_10773,N_10493);
or U11033 (N_11033,N_10280,N_10814);
nand U11034 (N_11034,N_10101,N_10150);
xor U11035 (N_11035,N_10371,N_10515);
nor U11036 (N_11036,N_10600,N_10267);
or U11037 (N_11037,N_10575,N_10542);
nand U11038 (N_11038,N_10969,N_10058);
and U11039 (N_11039,N_10130,N_10675);
xor U11040 (N_11040,N_10537,N_10100);
nand U11041 (N_11041,N_10254,N_10116);
nor U11042 (N_11042,N_10421,N_10591);
or U11043 (N_11043,N_10775,N_10483);
nor U11044 (N_11044,N_10195,N_10003);
nor U11045 (N_11045,N_10331,N_10782);
nor U11046 (N_11046,N_10990,N_10953);
and U11047 (N_11047,N_10526,N_10250);
or U11048 (N_11048,N_10946,N_10978);
and U11049 (N_11049,N_10970,N_10340);
and U11050 (N_11050,N_10963,N_10728);
and U11051 (N_11051,N_10696,N_10785);
nand U11052 (N_11052,N_10452,N_10241);
xor U11053 (N_11053,N_10900,N_10874);
nand U11054 (N_11054,N_10403,N_10377);
xor U11055 (N_11055,N_10805,N_10834);
nand U11056 (N_11056,N_10159,N_10044);
nand U11057 (N_11057,N_10294,N_10468);
xor U11058 (N_11058,N_10170,N_10618);
xor U11059 (N_11059,N_10567,N_10083);
nand U11060 (N_11060,N_10692,N_10664);
or U11061 (N_11061,N_10405,N_10629);
nor U11062 (N_11062,N_10311,N_10810);
nand U11063 (N_11063,N_10177,N_10579);
nand U11064 (N_11064,N_10726,N_10875);
or U11065 (N_11065,N_10394,N_10282);
and U11066 (N_11066,N_10107,N_10216);
and U11067 (N_11067,N_10804,N_10509);
nand U11068 (N_11068,N_10244,N_10186);
xor U11069 (N_11069,N_10842,N_10995);
nor U11070 (N_11070,N_10919,N_10770);
or U11071 (N_11071,N_10673,N_10632);
or U11072 (N_11072,N_10722,N_10736);
nor U11073 (N_11073,N_10516,N_10813);
or U11074 (N_11074,N_10147,N_10368);
or U11075 (N_11075,N_10760,N_10662);
nand U11076 (N_11076,N_10149,N_10559);
or U11077 (N_11077,N_10084,N_10108);
nor U11078 (N_11078,N_10157,N_10698);
and U11079 (N_11079,N_10507,N_10642);
nor U11080 (N_11080,N_10684,N_10426);
and U11081 (N_11081,N_10866,N_10134);
nor U11082 (N_11082,N_10174,N_10307);
nor U11083 (N_11083,N_10293,N_10755);
nand U11084 (N_11084,N_10208,N_10945);
nand U11085 (N_11085,N_10401,N_10073);
or U11086 (N_11086,N_10991,N_10329);
or U11087 (N_11087,N_10353,N_10603);
and U11088 (N_11088,N_10702,N_10308);
nor U11089 (N_11089,N_10711,N_10502);
nand U11090 (N_11090,N_10148,N_10409);
and U11091 (N_11091,N_10735,N_10580);
or U11092 (N_11092,N_10975,N_10938);
xnor U11093 (N_11093,N_10732,N_10626);
and U11094 (N_11094,N_10021,N_10712);
xnor U11095 (N_11095,N_10318,N_10747);
nand U11096 (N_11096,N_10270,N_10440);
and U11097 (N_11097,N_10503,N_10817);
or U11098 (N_11098,N_10521,N_10678);
nand U11099 (N_11099,N_10129,N_10410);
xor U11100 (N_11100,N_10927,N_10964);
and U11101 (N_11101,N_10120,N_10774);
or U11102 (N_11102,N_10202,N_10020);
or U11103 (N_11103,N_10248,N_10751);
and U11104 (N_11104,N_10392,N_10665);
and U11105 (N_11105,N_10533,N_10654);
or U11106 (N_11106,N_10441,N_10994);
or U11107 (N_11107,N_10843,N_10277);
xnor U11108 (N_11108,N_10458,N_10539);
and U11109 (N_11109,N_10047,N_10887);
nand U11110 (N_11110,N_10156,N_10776);
or U11111 (N_11111,N_10789,N_10436);
nand U11112 (N_11112,N_10480,N_10546);
or U11113 (N_11113,N_10781,N_10034);
nand U11114 (N_11114,N_10570,N_10608);
and U11115 (N_11115,N_10029,N_10278);
nor U11116 (N_11116,N_10976,N_10204);
nand U11117 (N_11117,N_10829,N_10336);
nand U11118 (N_11118,N_10222,N_10869);
and U11119 (N_11119,N_10973,N_10089);
nand U11120 (N_11120,N_10880,N_10158);
or U11121 (N_11121,N_10258,N_10636);
and U11122 (N_11122,N_10142,N_10897);
nor U11123 (N_11123,N_10131,N_10934);
and U11124 (N_11124,N_10955,N_10765);
or U11125 (N_11125,N_10399,N_10815);
nand U11126 (N_11126,N_10757,N_10788);
and U11127 (N_11127,N_10532,N_10323);
or U11128 (N_11128,N_10314,N_10260);
nor U11129 (N_11129,N_10556,N_10681);
and U11130 (N_11130,N_10651,N_10167);
nor U11131 (N_11131,N_10427,N_10614);
and U11132 (N_11132,N_10807,N_10265);
nor U11133 (N_11133,N_10469,N_10597);
or U11134 (N_11134,N_10552,N_10564);
and U11135 (N_11135,N_10040,N_10193);
and U11136 (N_11136,N_10137,N_10959);
or U11137 (N_11137,N_10463,N_10205);
and U11138 (N_11138,N_10855,N_10358);
and U11139 (N_11139,N_10498,N_10062);
or U11140 (N_11140,N_10431,N_10848);
nor U11141 (N_11141,N_10752,N_10647);
nor U11142 (N_11142,N_10444,N_10355);
and U11143 (N_11143,N_10612,N_10850);
nor U11144 (N_11144,N_10327,N_10962);
nor U11145 (N_11145,N_10911,N_10272);
and U11146 (N_11146,N_10933,N_10950);
nor U11147 (N_11147,N_10871,N_10190);
nand U11148 (N_11148,N_10001,N_10569);
nor U11149 (N_11149,N_10139,N_10416);
and U11150 (N_11150,N_10854,N_10987);
nor U11151 (N_11151,N_10831,N_10916);
nand U11152 (N_11152,N_10461,N_10052);
or U11153 (N_11153,N_10103,N_10734);
or U11154 (N_11154,N_10283,N_10827);
nor U11155 (N_11155,N_10422,N_10361);
or U11156 (N_11156,N_10085,N_10198);
nor U11157 (N_11157,N_10902,N_10197);
or U11158 (N_11158,N_10921,N_10345);
nand U11159 (N_11159,N_10445,N_10816);
and U11160 (N_11160,N_10941,N_10408);
nor U11161 (N_11161,N_10160,N_10562);
or U11162 (N_11162,N_10727,N_10883);
and U11163 (N_11163,N_10906,N_10086);
or U11164 (N_11164,N_10217,N_10928);
xnor U11165 (N_11165,N_10002,N_10032);
nand U11166 (N_11166,N_10800,N_10189);
or U11167 (N_11167,N_10840,N_10457);
nor U11168 (N_11168,N_10153,N_10046);
and U11169 (N_11169,N_10106,N_10140);
nor U11170 (N_11170,N_10402,N_10793);
and U11171 (N_11171,N_10476,N_10545);
nor U11172 (N_11172,N_10364,N_10663);
or U11173 (N_11173,N_10943,N_10847);
and U11174 (N_11174,N_10211,N_10650);
nand U11175 (N_11175,N_10375,N_10301);
nor U11176 (N_11176,N_10033,N_10263);
or U11177 (N_11177,N_10404,N_10386);
xnor U11178 (N_11178,N_10742,N_10879);
xnor U11179 (N_11179,N_10864,N_10219);
nand U11180 (N_11180,N_10535,N_10929);
or U11181 (N_11181,N_10281,N_10400);
nand U11182 (N_11182,N_10004,N_10669);
nand U11183 (N_11183,N_10312,N_10454);
nand U11184 (N_11184,N_10997,N_10287);
xor U11185 (N_11185,N_10598,N_10342);
nand U11186 (N_11186,N_10910,N_10753);
nand U11187 (N_11187,N_10924,N_10014);
nor U11188 (N_11188,N_10853,N_10746);
nand U11189 (N_11189,N_10667,N_10699);
and U11190 (N_11190,N_10035,N_10676);
and U11191 (N_11191,N_10315,N_10583);
nand U11192 (N_11192,N_10517,N_10382);
and U11193 (N_11193,N_10284,N_10655);
or U11194 (N_11194,N_10749,N_10661);
or U11195 (N_11195,N_10641,N_10707);
nand U11196 (N_11196,N_10931,N_10473);
and U11197 (N_11197,N_10939,N_10333);
and U11198 (N_11198,N_10660,N_10719);
or U11199 (N_11199,N_10859,N_10031);
nor U11200 (N_11200,N_10522,N_10892);
or U11201 (N_11201,N_10993,N_10234);
nor U11202 (N_11202,N_10111,N_10885);
nor U11203 (N_11203,N_10487,N_10981);
or U11204 (N_11204,N_10909,N_10347);
nor U11205 (N_11205,N_10601,N_10500);
or U11206 (N_11206,N_10604,N_10703);
and U11207 (N_11207,N_10767,N_10586);
or U11208 (N_11208,N_10239,N_10743);
xor U11209 (N_11209,N_10630,N_10538);
nor U11210 (N_11210,N_10363,N_10151);
nor U11211 (N_11211,N_10467,N_10479);
or U11212 (N_11212,N_10966,N_10819);
or U11213 (N_11213,N_10602,N_10109);
nand U11214 (N_11214,N_10482,N_10940);
xnor U11215 (N_11215,N_10888,N_10616);
xnor U11216 (N_11216,N_10112,N_10985);
and U11217 (N_11217,N_10224,N_10433);
nand U11218 (N_11218,N_10132,N_10412);
or U11219 (N_11219,N_10242,N_10037);
nor U11220 (N_11220,N_10229,N_10143);
nor U11221 (N_11221,N_10074,N_10594);
xor U11222 (N_11222,N_10247,N_10704);
or U11223 (N_11223,N_10974,N_10808);
or U11224 (N_11224,N_10080,N_10841);
nand U11225 (N_11225,N_10890,N_10872);
nand U11226 (N_11226,N_10983,N_10024);
or U11227 (N_11227,N_10395,N_10235);
and U11228 (N_11228,N_10064,N_10961);
nand U11229 (N_11229,N_10012,N_10756);
and U11230 (N_11230,N_10212,N_10209);
or U11231 (N_11231,N_10741,N_10508);
nand U11232 (N_11232,N_10297,N_10724);
nor U11233 (N_11233,N_10530,N_10429);
or U11234 (N_11234,N_10339,N_10464);
or U11235 (N_11235,N_10268,N_10956);
nand U11236 (N_11236,N_10185,N_10439);
nand U11237 (N_11237,N_10288,N_10481);
nor U11238 (N_11238,N_10649,N_10419);
or U11239 (N_11239,N_10206,N_10820);
xnor U11240 (N_11240,N_10764,N_10477);
nor U11241 (N_11241,N_10356,N_10446);
nand U11242 (N_11242,N_10173,N_10379);
and U11243 (N_11243,N_10889,N_10652);
or U11244 (N_11244,N_10540,N_10346);
and U11245 (N_11245,N_10279,N_10777);
nand U11246 (N_11246,N_10447,N_10054);
nand U11247 (N_11247,N_10243,N_10745);
nand U11248 (N_11248,N_10894,N_10682);
nor U11249 (N_11249,N_10648,N_10677);
or U11250 (N_11250,N_10826,N_10589);
xnor U11251 (N_11251,N_10486,N_10475);
nor U11252 (N_11252,N_10462,N_10450);
nor U11253 (N_11253,N_10877,N_10920);
xnor U11254 (N_11254,N_10196,N_10918);
or U11255 (N_11255,N_10484,N_10768);
xor U11256 (N_11256,N_10466,N_10178);
nand U11257 (N_11257,N_10126,N_10796);
or U11258 (N_11258,N_10615,N_10388);
nor U11259 (N_11259,N_10972,N_10194);
nand U11260 (N_11260,N_10896,N_10011);
xnor U11261 (N_11261,N_10723,N_10668);
nor U11262 (N_11262,N_10895,N_10369);
or U11263 (N_11263,N_10320,N_10659);
and U11264 (N_11264,N_10273,N_10366);
or U11265 (N_11265,N_10304,N_10882);
nand U11266 (N_11266,N_10124,N_10519);
or U11267 (N_11267,N_10513,N_10551);
nand U11268 (N_11268,N_10053,N_10863);
and U11269 (N_11269,N_10341,N_10082);
nor U11270 (N_11270,N_10261,N_10958);
nor U11271 (N_11271,N_10354,N_10631);
nor U11272 (N_11272,N_10117,N_10182);
xnor U11273 (N_11273,N_10442,N_10451);
xor U11274 (N_11274,N_10010,N_10227);
and U11275 (N_11275,N_10541,N_10725);
nor U11276 (N_11276,N_10305,N_10693);
nand U11277 (N_11277,N_10061,N_10754);
nand U11278 (N_11278,N_10771,N_10790);
and U11279 (N_11279,N_10657,N_10565);
or U11280 (N_11280,N_10857,N_10700);
and U11281 (N_11281,N_10965,N_10821);
nand U11282 (N_11282,N_10245,N_10013);
nor U11283 (N_11283,N_10015,N_10334);
xnor U11284 (N_11284,N_10759,N_10128);
nor U11285 (N_11285,N_10671,N_10495);
or U11286 (N_11286,N_10512,N_10070);
and U11287 (N_11287,N_10494,N_10465);
or U11288 (N_11288,N_10325,N_10772);
nand U11289 (N_11289,N_10582,N_10936);
nand U11290 (N_11290,N_10285,N_10915);
nor U11291 (N_11291,N_10060,N_10057);
nand U11292 (N_11292,N_10504,N_10544);
xor U11293 (N_11293,N_10059,N_10091);
nor U11294 (N_11294,N_10118,N_10335);
or U11295 (N_11295,N_10948,N_10592);
and U11296 (N_11296,N_10766,N_10731);
nor U11297 (N_11297,N_10729,N_10349);
nor U11298 (N_11298,N_10846,N_10694);
nor U11299 (N_11299,N_10397,N_10324);
nand U11300 (N_11300,N_10683,N_10098);
or U11301 (N_11301,N_10296,N_10845);
or U11302 (N_11302,N_10175,N_10769);
and U11303 (N_11303,N_10501,N_10210);
nor U11304 (N_11304,N_10870,N_10554);
nand U11305 (N_11305,N_10520,N_10374);
nand U11306 (N_11306,N_10343,N_10437);
nor U11307 (N_11307,N_10606,N_10624);
nand U11308 (N_11308,N_10230,N_10471);
nand U11309 (N_11309,N_10192,N_10670);
or U11310 (N_11310,N_10917,N_10351);
and U11311 (N_11311,N_10218,N_10069);
or U11312 (N_11312,N_10274,N_10555);
nor U11313 (N_11313,N_10007,N_10240);
and U11314 (N_11314,N_10104,N_10935);
nor U11315 (N_11315,N_10373,N_10259);
or U11316 (N_11316,N_10418,N_10133);
nand U11317 (N_11317,N_10051,N_10638);
nor U11318 (N_11318,N_10572,N_10068);
nor U11319 (N_11319,N_10075,N_10337);
nor U11320 (N_11320,N_10529,N_10856);
or U11321 (N_11321,N_10348,N_10949);
or U11322 (N_11322,N_10844,N_10063);
nor U11323 (N_11323,N_10036,N_10531);
nor U11324 (N_11324,N_10784,N_10135);
or U11325 (N_11325,N_10472,N_10982);
and U11326 (N_11326,N_10947,N_10645);
xor U11327 (N_11327,N_10049,N_10378);
nand U11328 (N_11328,N_10867,N_10023);
and U11329 (N_11329,N_10275,N_10792);
xnor U11330 (N_11330,N_10705,N_10653);
nor U11331 (N_11331,N_10127,N_10865);
nand U11332 (N_11332,N_10191,N_10758);
nand U11333 (N_11333,N_10903,N_10658);
nor U11334 (N_11334,N_10593,N_10607);
nand U11335 (N_11335,N_10590,N_10822);
or U11336 (N_11336,N_10038,N_10706);
or U11337 (N_11337,N_10621,N_10860);
nand U11338 (N_11338,N_10092,N_10605);
nor U11339 (N_11339,N_10884,N_10999);
nand U11340 (N_11340,N_10171,N_10491);
and U11341 (N_11341,N_10271,N_10306);
nand U11342 (N_11342,N_10791,N_10858);
nand U11343 (N_11343,N_10907,N_10188);
xor U11344 (N_11344,N_10048,N_10951);
and U11345 (N_11345,N_10079,N_10330);
nand U11346 (N_11346,N_10674,N_10839);
nor U11347 (N_11347,N_10640,N_10362);
xnor U11348 (N_11348,N_10372,N_10102);
and U11349 (N_11349,N_10276,N_10055);
nand U11350 (N_11350,N_10425,N_10812);
xnor U11351 (N_11351,N_10214,N_10381);
nor U11352 (N_11352,N_10628,N_10113);
nor U11353 (N_11353,N_10709,N_10459);
or U11354 (N_11354,N_10563,N_10322);
xnor U11355 (N_11355,N_10837,N_10609);
nand U11356 (N_11356,N_10566,N_10971);
nor U11357 (N_11357,N_10203,N_10490);
nor U11358 (N_11358,N_10666,N_10795);
and U11359 (N_11359,N_10223,N_10169);
or U11360 (N_11360,N_10317,N_10411);
nand U11361 (N_11361,N_10625,N_10376);
nor U11362 (N_11362,N_10187,N_10988);
nor U11363 (N_11363,N_10794,N_10221);
or U11364 (N_11364,N_10558,N_10656);
nor U11365 (N_11365,N_10215,N_10691);
nand U11366 (N_11366,N_10585,N_10455);
nor U11367 (N_11367,N_10290,N_10492);
nor U11368 (N_11368,N_10423,N_10923);
and U11369 (N_11369,N_10016,N_10161);
or U11370 (N_11370,N_10721,N_10398);
xor U11371 (N_11371,N_10041,N_10144);
or U11372 (N_11372,N_10536,N_10071);
and U11373 (N_11373,N_10733,N_10688);
nor U11374 (N_11374,N_10415,N_10039);
and U11375 (N_11375,N_10154,N_10028);
xor U11376 (N_11376,N_10499,N_10783);
nand U11377 (N_11377,N_10695,N_10300);
xor U11378 (N_11378,N_10299,N_10960);
nand U11379 (N_11379,N_10543,N_10136);
nor U11380 (N_11380,N_10199,N_10163);
nor U11381 (N_11381,N_10026,N_10828);
nand U11382 (N_11382,N_10228,N_10849);
nor U11383 (N_11383,N_10017,N_10852);
and U11384 (N_11384,N_10319,N_10967);
or U11385 (N_11385,N_10672,N_10942);
nor U11386 (N_11386,N_10438,N_10635);
nand U11387 (N_11387,N_10687,N_10099);
nor U11388 (N_11388,N_10344,N_10778);
nand U11389 (N_11389,N_10525,N_10779);
and U11390 (N_11390,N_10328,N_10549);
or U11391 (N_11391,N_10380,N_10025);
or U11392 (N_11392,N_10710,N_10977);
and U11393 (N_11393,N_10256,N_10155);
nor U11394 (N_11394,N_10321,N_10286);
nor U11395 (N_11395,N_10005,N_10088);
and U11396 (N_11396,N_10213,N_10644);
or U11397 (N_11397,N_10527,N_10701);
and U11398 (N_11398,N_10430,N_10717);
and U11399 (N_11399,N_10180,N_10886);
and U11400 (N_11400,N_10930,N_10022);
nor U11401 (N_11401,N_10291,N_10008);
xor U11402 (N_11402,N_10310,N_10548);
and U11403 (N_11403,N_10833,N_10257);
and U11404 (N_11404,N_10201,N_10251);
xor U11405 (N_11405,N_10183,N_10689);
nor U11406 (N_11406,N_10269,N_10434);
or U11407 (N_11407,N_10238,N_10748);
and U11408 (N_11408,N_10138,N_10876);
or U11409 (N_11409,N_10680,N_10152);
nor U11410 (N_11410,N_10176,N_10096);
nor U11411 (N_11411,N_10391,N_10697);
xor U11412 (N_11412,N_10714,N_10489);
or U11413 (N_11413,N_10456,N_10617);
nand U11414 (N_11414,N_10359,N_10744);
nand U11415 (N_11415,N_10087,N_10357);
nor U11416 (N_11416,N_10119,N_10164);
or U11417 (N_11417,N_10313,N_10998);
nand U11418 (N_11418,N_10045,N_10679);
or U11419 (N_11419,N_10578,N_10352);
or U11420 (N_11420,N_10851,N_10019);
or U11421 (N_11421,N_10497,N_10389);
nand U11422 (N_11422,N_10832,N_10485);
or U11423 (N_11423,N_10443,N_10514);
xnor U11424 (N_11424,N_10878,N_10006);
and U11425 (N_11425,N_10868,N_10740);
and U11426 (N_11426,N_10761,N_10818);
nor U11427 (N_11427,N_10925,N_10825);
and U11428 (N_11428,N_10926,N_10065);
and U11429 (N_11429,N_10384,N_10449);
and U11430 (N_11430,N_10488,N_10553);
or U11431 (N_11431,N_10577,N_10560);
and U11432 (N_11432,N_10122,N_10809);
and U11433 (N_11433,N_10246,N_10181);
and U11434 (N_11434,N_10989,N_10797);
xnor U11435 (N_11435,N_10110,N_10596);
nor U11436 (N_11436,N_10407,N_10370);
nand U11437 (N_11437,N_10385,N_10432);
and U11438 (N_11438,N_10413,N_10332);
or U11439 (N_11439,N_10367,N_10168);
and U11440 (N_11440,N_10715,N_10225);
and U11441 (N_11441,N_10292,N_10121);
and U11442 (N_11442,N_10496,N_10326);
or U11443 (N_11443,N_10620,N_10510);
and U11444 (N_11444,N_10236,N_10979);
or U11445 (N_11445,N_10266,N_10097);
and U11446 (N_11446,N_10387,N_10861);
nand U11447 (N_11447,N_10093,N_10619);
or U11448 (N_11448,N_10528,N_10523);
xor U11449 (N_11449,N_10478,N_10165);
or U11450 (N_11450,N_10623,N_10393);
or U11451 (N_11451,N_10094,N_10588);
nand U11452 (N_11452,N_10611,N_10220);
and U11453 (N_11453,N_10289,N_10406);
or U11454 (N_11454,N_10738,N_10424);
nor U11455 (N_11455,N_10862,N_10584);
nor U11456 (N_11456,N_10685,N_10639);
and U11457 (N_11457,N_10557,N_10262);
nor U11458 (N_11458,N_10836,N_10996);
nand U11459 (N_11459,N_10050,N_10505);
or U11460 (N_11460,N_10166,N_10081);
and U11461 (N_11461,N_10587,N_10524);
and U11462 (N_11462,N_10763,N_10798);
or U11463 (N_11463,N_10066,N_10396);
or U11464 (N_11464,N_10547,N_10042);
nand U11465 (N_11465,N_10179,N_10435);
and U11466 (N_11466,N_10613,N_10231);
nor U11467 (N_11467,N_10237,N_10891);
or U11468 (N_11468,N_10992,N_10571);
nor U11469 (N_11469,N_10968,N_10739);
nor U11470 (N_11470,N_10690,N_10986);
nand U11471 (N_11471,N_10904,N_10801);
xor U11472 (N_11472,N_10599,N_10984);
xnor U11473 (N_11473,N_10030,N_10076);
nor U11474 (N_11474,N_10141,N_10750);
nand U11475 (N_11475,N_10720,N_10595);
xor U11476 (N_11476,N_10226,N_10264);
and U11477 (N_11477,N_10610,N_10200);
or U11478 (N_11478,N_10561,N_10633);
or U11479 (N_11479,N_10905,N_10105);
nor U11480 (N_11480,N_10716,N_10898);
nand U11481 (N_11481,N_10145,N_10302);
xor U11482 (N_11482,N_10786,N_10922);
nor U11483 (N_11483,N_10899,N_10255);
nor U11484 (N_11484,N_10730,N_10881);
and U11485 (N_11485,N_10072,N_10056);
and U11486 (N_11486,N_10824,N_10646);
nand U11487 (N_11487,N_10428,N_10713);
nand U11488 (N_11488,N_10077,N_10115);
nor U11489 (N_11489,N_10550,N_10232);
nor U11490 (N_11490,N_10383,N_10980);
nor U11491 (N_11491,N_10637,N_10957);
nand U11492 (N_11492,N_10000,N_10460);
and U11493 (N_11493,N_10414,N_10009);
or U11494 (N_11494,N_10912,N_10581);
nor U11495 (N_11495,N_10576,N_10573);
nor U11496 (N_11496,N_10780,N_10568);
nor U11497 (N_11497,N_10506,N_10295);
nand U11498 (N_11498,N_10067,N_10932);
nor U11499 (N_11499,N_10252,N_10643);
or U11500 (N_11500,N_10301,N_10577);
nor U11501 (N_11501,N_10444,N_10706);
and U11502 (N_11502,N_10440,N_10724);
or U11503 (N_11503,N_10366,N_10058);
nor U11504 (N_11504,N_10948,N_10937);
and U11505 (N_11505,N_10580,N_10957);
nor U11506 (N_11506,N_10931,N_10681);
and U11507 (N_11507,N_10381,N_10003);
xor U11508 (N_11508,N_10807,N_10465);
or U11509 (N_11509,N_10531,N_10147);
and U11510 (N_11510,N_10344,N_10733);
or U11511 (N_11511,N_10240,N_10055);
nor U11512 (N_11512,N_10858,N_10102);
and U11513 (N_11513,N_10726,N_10133);
nand U11514 (N_11514,N_10145,N_10917);
nor U11515 (N_11515,N_10700,N_10498);
or U11516 (N_11516,N_10312,N_10940);
nand U11517 (N_11517,N_10618,N_10527);
xnor U11518 (N_11518,N_10208,N_10811);
nor U11519 (N_11519,N_10615,N_10844);
nand U11520 (N_11520,N_10479,N_10295);
nor U11521 (N_11521,N_10239,N_10236);
or U11522 (N_11522,N_10518,N_10216);
or U11523 (N_11523,N_10957,N_10272);
or U11524 (N_11524,N_10271,N_10384);
xor U11525 (N_11525,N_10859,N_10515);
nand U11526 (N_11526,N_10439,N_10833);
and U11527 (N_11527,N_10227,N_10422);
or U11528 (N_11528,N_10064,N_10095);
nand U11529 (N_11529,N_10084,N_10802);
and U11530 (N_11530,N_10063,N_10770);
xor U11531 (N_11531,N_10004,N_10050);
nand U11532 (N_11532,N_10123,N_10020);
and U11533 (N_11533,N_10818,N_10202);
or U11534 (N_11534,N_10894,N_10721);
nand U11535 (N_11535,N_10154,N_10808);
xor U11536 (N_11536,N_10765,N_10767);
and U11537 (N_11537,N_10271,N_10489);
nand U11538 (N_11538,N_10835,N_10983);
nor U11539 (N_11539,N_10688,N_10029);
nand U11540 (N_11540,N_10995,N_10563);
nand U11541 (N_11541,N_10193,N_10340);
or U11542 (N_11542,N_10256,N_10492);
xnor U11543 (N_11543,N_10746,N_10935);
and U11544 (N_11544,N_10407,N_10280);
nand U11545 (N_11545,N_10289,N_10304);
or U11546 (N_11546,N_10394,N_10757);
nand U11547 (N_11547,N_10853,N_10096);
or U11548 (N_11548,N_10922,N_10167);
xor U11549 (N_11549,N_10854,N_10363);
and U11550 (N_11550,N_10388,N_10202);
xor U11551 (N_11551,N_10484,N_10728);
nand U11552 (N_11552,N_10953,N_10282);
or U11553 (N_11553,N_10780,N_10831);
or U11554 (N_11554,N_10286,N_10723);
or U11555 (N_11555,N_10477,N_10962);
nand U11556 (N_11556,N_10708,N_10084);
nand U11557 (N_11557,N_10238,N_10153);
xnor U11558 (N_11558,N_10350,N_10871);
and U11559 (N_11559,N_10321,N_10322);
and U11560 (N_11560,N_10229,N_10880);
nor U11561 (N_11561,N_10087,N_10061);
nor U11562 (N_11562,N_10721,N_10364);
nor U11563 (N_11563,N_10863,N_10371);
xor U11564 (N_11564,N_10304,N_10978);
nand U11565 (N_11565,N_10260,N_10717);
nand U11566 (N_11566,N_10555,N_10093);
and U11567 (N_11567,N_10347,N_10780);
or U11568 (N_11568,N_10311,N_10533);
and U11569 (N_11569,N_10232,N_10158);
nand U11570 (N_11570,N_10611,N_10049);
nand U11571 (N_11571,N_10924,N_10152);
nand U11572 (N_11572,N_10958,N_10576);
nand U11573 (N_11573,N_10461,N_10275);
nand U11574 (N_11574,N_10059,N_10894);
xor U11575 (N_11575,N_10638,N_10834);
nor U11576 (N_11576,N_10392,N_10422);
or U11577 (N_11577,N_10306,N_10281);
and U11578 (N_11578,N_10553,N_10130);
or U11579 (N_11579,N_10655,N_10623);
and U11580 (N_11580,N_10668,N_10542);
nor U11581 (N_11581,N_10004,N_10480);
and U11582 (N_11582,N_10244,N_10867);
or U11583 (N_11583,N_10762,N_10330);
and U11584 (N_11584,N_10356,N_10596);
nor U11585 (N_11585,N_10156,N_10495);
nor U11586 (N_11586,N_10426,N_10139);
nor U11587 (N_11587,N_10547,N_10104);
nand U11588 (N_11588,N_10377,N_10862);
or U11589 (N_11589,N_10486,N_10617);
nor U11590 (N_11590,N_10978,N_10386);
nand U11591 (N_11591,N_10996,N_10988);
nand U11592 (N_11592,N_10092,N_10935);
nand U11593 (N_11593,N_10709,N_10235);
and U11594 (N_11594,N_10989,N_10718);
or U11595 (N_11595,N_10358,N_10716);
nor U11596 (N_11596,N_10009,N_10987);
or U11597 (N_11597,N_10767,N_10740);
and U11598 (N_11598,N_10438,N_10607);
or U11599 (N_11599,N_10966,N_10455);
nand U11600 (N_11600,N_10453,N_10551);
or U11601 (N_11601,N_10823,N_10431);
xnor U11602 (N_11602,N_10206,N_10273);
or U11603 (N_11603,N_10434,N_10375);
or U11604 (N_11604,N_10775,N_10558);
nand U11605 (N_11605,N_10311,N_10832);
nand U11606 (N_11606,N_10559,N_10998);
xor U11607 (N_11607,N_10954,N_10237);
and U11608 (N_11608,N_10585,N_10314);
xor U11609 (N_11609,N_10951,N_10983);
and U11610 (N_11610,N_10156,N_10352);
and U11611 (N_11611,N_10031,N_10196);
xnor U11612 (N_11612,N_10663,N_10568);
nand U11613 (N_11613,N_10120,N_10043);
nor U11614 (N_11614,N_10629,N_10417);
nand U11615 (N_11615,N_10094,N_10365);
and U11616 (N_11616,N_10065,N_10048);
nor U11617 (N_11617,N_10929,N_10832);
nand U11618 (N_11618,N_10925,N_10665);
and U11619 (N_11619,N_10701,N_10697);
nand U11620 (N_11620,N_10687,N_10363);
and U11621 (N_11621,N_10984,N_10987);
xor U11622 (N_11622,N_10807,N_10926);
and U11623 (N_11623,N_10189,N_10338);
or U11624 (N_11624,N_10132,N_10608);
or U11625 (N_11625,N_10075,N_10178);
and U11626 (N_11626,N_10548,N_10886);
xnor U11627 (N_11627,N_10749,N_10243);
nand U11628 (N_11628,N_10046,N_10752);
nand U11629 (N_11629,N_10827,N_10844);
nand U11630 (N_11630,N_10154,N_10799);
and U11631 (N_11631,N_10589,N_10281);
xnor U11632 (N_11632,N_10469,N_10131);
nand U11633 (N_11633,N_10820,N_10830);
nor U11634 (N_11634,N_10724,N_10184);
nor U11635 (N_11635,N_10298,N_10972);
and U11636 (N_11636,N_10872,N_10302);
nand U11637 (N_11637,N_10390,N_10879);
and U11638 (N_11638,N_10715,N_10639);
or U11639 (N_11639,N_10526,N_10350);
or U11640 (N_11640,N_10964,N_10907);
nand U11641 (N_11641,N_10315,N_10550);
or U11642 (N_11642,N_10123,N_10765);
or U11643 (N_11643,N_10784,N_10988);
nor U11644 (N_11644,N_10656,N_10118);
nand U11645 (N_11645,N_10276,N_10416);
and U11646 (N_11646,N_10630,N_10367);
or U11647 (N_11647,N_10254,N_10500);
or U11648 (N_11648,N_10668,N_10956);
or U11649 (N_11649,N_10782,N_10068);
and U11650 (N_11650,N_10785,N_10005);
nor U11651 (N_11651,N_10466,N_10372);
xor U11652 (N_11652,N_10711,N_10862);
nand U11653 (N_11653,N_10045,N_10450);
and U11654 (N_11654,N_10174,N_10688);
xor U11655 (N_11655,N_10914,N_10543);
and U11656 (N_11656,N_10731,N_10680);
and U11657 (N_11657,N_10076,N_10654);
nand U11658 (N_11658,N_10468,N_10647);
nor U11659 (N_11659,N_10311,N_10839);
nand U11660 (N_11660,N_10085,N_10306);
and U11661 (N_11661,N_10954,N_10321);
nand U11662 (N_11662,N_10285,N_10606);
nand U11663 (N_11663,N_10709,N_10404);
and U11664 (N_11664,N_10722,N_10973);
or U11665 (N_11665,N_10490,N_10984);
or U11666 (N_11666,N_10662,N_10892);
nand U11667 (N_11667,N_10243,N_10228);
nor U11668 (N_11668,N_10295,N_10645);
or U11669 (N_11669,N_10961,N_10437);
nor U11670 (N_11670,N_10048,N_10303);
or U11671 (N_11671,N_10764,N_10982);
nor U11672 (N_11672,N_10997,N_10503);
nand U11673 (N_11673,N_10946,N_10819);
nand U11674 (N_11674,N_10485,N_10614);
nor U11675 (N_11675,N_10213,N_10027);
nor U11676 (N_11676,N_10424,N_10034);
nor U11677 (N_11677,N_10945,N_10551);
and U11678 (N_11678,N_10254,N_10852);
and U11679 (N_11679,N_10071,N_10977);
and U11680 (N_11680,N_10480,N_10453);
nand U11681 (N_11681,N_10844,N_10498);
and U11682 (N_11682,N_10957,N_10331);
or U11683 (N_11683,N_10064,N_10723);
or U11684 (N_11684,N_10607,N_10576);
or U11685 (N_11685,N_10351,N_10057);
and U11686 (N_11686,N_10122,N_10916);
and U11687 (N_11687,N_10476,N_10867);
or U11688 (N_11688,N_10301,N_10027);
nor U11689 (N_11689,N_10945,N_10381);
and U11690 (N_11690,N_10520,N_10383);
or U11691 (N_11691,N_10793,N_10753);
nand U11692 (N_11692,N_10432,N_10378);
or U11693 (N_11693,N_10081,N_10033);
nand U11694 (N_11694,N_10902,N_10435);
xor U11695 (N_11695,N_10953,N_10736);
or U11696 (N_11696,N_10570,N_10089);
nand U11697 (N_11697,N_10664,N_10415);
nor U11698 (N_11698,N_10883,N_10852);
nor U11699 (N_11699,N_10071,N_10228);
nand U11700 (N_11700,N_10932,N_10401);
and U11701 (N_11701,N_10605,N_10342);
nand U11702 (N_11702,N_10146,N_10895);
nand U11703 (N_11703,N_10364,N_10564);
and U11704 (N_11704,N_10347,N_10129);
or U11705 (N_11705,N_10943,N_10658);
and U11706 (N_11706,N_10880,N_10146);
or U11707 (N_11707,N_10004,N_10350);
and U11708 (N_11708,N_10846,N_10438);
xnor U11709 (N_11709,N_10783,N_10379);
or U11710 (N_11710,N_10307,N_10204);
or U11711 (N_11711,N_10453,N_10745);
nor U11712 (N_11712,N_10495,N_10374);
nor U11713 (N_11713,N_10920,N_10539);
xnor U11714 (N_11714,N_10649,N_10545);
and U11715 (N_11715,N_10361,N_10883);
and U11716 (N_11716,N_10034,N_10791);
or U11717 (N_11717,N_10039,N_10249);
and U11718 (N_11718,N_10492,N_10128);
and U11719 (N_11719,N_10089,N_10572);
and U11720 (N_11720,N_10486,N_10750);
xnor U11721 (N_11721,N_10055,N_10507);
xnor U11722 (N_11722,N_10927,N_10055);
nand U11723 (N_11723,N_10613,N_10000);
nand U11724 (N_11724,N_10657,N_10995);
nand U11725 (N_11725,N_10605,N_10860);
or U11726 (N_11726,N_10137,N_10346);
nand U11727 (N_11727,N_10080,N_10821);
xor U11728 (N_11728,N_10472,N_10069);
nand U11729 (N_11729,N_10678,N_10401);
nor U11730 (N_11730,N_10483,N_10974);
or U11731 (N_11731,N_10326,N_10381);
or U11732 (N_11732,N_10823,N_10807);
or U11733 (N_11733,N_10933,N_10939);
nand U11734 (N_11734,N_10998,N_10036);
nor U11735 (N_11735,N_10956,N_10613);
nand U11736 (N_11736,N_10062,N_10569);
nand U11737 (N_11737,N_10281,N_10425);
nor U11738 (N_11738,N_10529,N_10580);
and U11739 (N_11739,N_10258,N_10206);
nand U11740 (N_11740,N_10181,N_10171);
and U11741 (N_11741,N_10514,N_10077);
and U11742 (N_11742,N_10999,N_10397);
nand U11743 (N_11743,N_10564,N_10828);
nor U11744 (N_11744,N_10359,N_10105);
or U11745 (N_11745,N_10530,N_10686);
nand U11746 (N_11746,N_10891,N_10164);
or U11747 (N_11747,N_10787,N_10719);
nand U11748 (N_11748,N_10814,N_10828);
or U11749 (N_11749,N_10969,N_10223);
and U11750 (N_11750,N_10571,N_10783);
or U11751 (N_11751,N_10436,N_10672);
nand U11752 (N_11752,N_10137,N_10444);
nor U11753 (N_11753,N_10639,N_10304);
nand U11754 (N_11754,N_10366,N_10577);
and U11755 (N_11755,N_10945,N_10514);
or U11756 (N_11756,N_10335,N_10314);
nand U11757 (N_11757,N_10764,N_10466);
nand U11758 (N_11758,N_10322,N_10341);
nor U11759 (N_11759,N_10208,N_10558);
or U11760 (N_11760,N_10073,N_10270);
or U11761 (N_11761,N_10382,N_10174);
xor U11762 (N_11762,N_10579,N_10559);
xor U11763 (N_11763,N_10744,N_10522);
xnor U11764 (N_11764,N_10459,N_10272);
or U11765 (N_11765,N_10340,N_10471);
or U11766 (N_11766,N_10980,N_10786);
or U11767 (N_11767,N_10003,N_10267);
nor U11768 (N_11768,N_10476,N_10281);
nand U11769 (N_11769,N_10595,N_10994);
or U11770 (N_11770,N_10334,N_10501);
and U11771 (N_11771,N_10228,N_10998);
xor U11772 (N_11772,N_10091,N_10678);
or U11773 (N_11773,N_10410,N_10988);
nor U11774 (N_11774,N_10693,N_10555);
or U11775 (N_11775,N_10518,N_10909);
nand U11776 (N_11776,N_10319,N_10343);
nor U11777 (N_11777,N_10946,N_10431);
xor U11778 (N_11778,N_10851,N_10556);
and U11779 (N_11779,N_10900,N_10884);
nor U11780 (N_11780,N_10601,N_10070);
or U11781 (N_11781,N_10896,N_10608);
and U11782 (N_11782,N_10839,N_10537);
nand U11783 (N_11783,N_10835,N_10695);
or U11784 (N_11784,N_10371,N_10454);
xnor U11785 (N_11785,N_10010,N_10941);
nor U11786 (N_11786,N_10169,N_10550);
nor U11787 (N_11787,N_10031,N_10995);
nor U11788 (N_11788,N_10797,N_10430);
nand U11789 (N_11789,N_10300,N_10628);
nand U11790 (N_11790,N_10407,N_10648);
nor U11791 (N_11791,N_10086,N_10265);
or U11792 (N_11792,N_10168,N_10038);
or U11793 (N_11793,N_10454,N_10259);
and U11794 (N_11794,N_10160,N_10486);
or U11795 (N_11795,N_10827,N_10600);
nand U11796 (N_11796,N_10497,N_10843);
and U11797 (N_11797,N_10700,N_10772);
nor U11798 (N_11798,N_10713,N_10727);
nand U11799 (N_11799,N_10145,N_10194);
nand U11800 (N_11800,N_10385,N_10183);
and U11801 (N_11801,N_10272,N_10345);
and U11802 (N_11802,N_10091,N_10198);
or U11803 (N_11803,N_10743,N_10428);
and U11804 (N_11804,N_10817,N_10602);
nand U11805 (N_11805,N_10265,N_10340);
or U11806 (N_11806,N_10091,N_10223);
and U11807 (N_11807,N_10283,N_10976);
xnor U11808 (N_11808,N_10549,N_10346);
nor U11809 (N_11809,N_10574,N_10903);
nand U11810 (N_11810,N_10841,N_10852);
xnor U11811 (N_11811,N_10834,N_10807);
and U11812 (N_11812,N_10302,N_10227);
nand U11813 (N_11813,N_10850,N_10497);
nand U11814 (N_11814,N_10375,N_10838);
and U11815 (N_11815,N_10860,N_10689);
and U11816 (N_11816,N_10097,N_10370);
and U11817 (N_11817,N_10104,N_10047);
xnor U11818 (N_11818,N_10852,N_10052);
or U11819 (N_11819,N_10674,N_10321);
nand U11820 (N_11820,N_10557,N_10189);
and U11821 (N_11821,N_10664,N_10269);
nor U11822 (N_11822,N_10772,N_10623);
nand U11823 (N_11823,N_10985,N_10195);
and U11824 (N_11824,N_10383,N_10197);
nand U11825 (N_11825,N_10382,N_10953);
or U11826 (N_11826,N_10521,N_10740);
nor U11827 (N_11827,N_10798,N_10969);
or U11828 (N_11828,N_10173,N_10343);
nand U11829 (N_11829,N_10899,N_10468);
and U11830 (N_11830,N_10072,N_10722);
or U11831 (N_11831,N_10455,N_10866);
nand U11832 (N_11832,N_10859,N_10649);
or U11833 (N_11833,N_10872,N_10194);
nand U11834 (N_11834,N_10999,N_10039);
nor U11835 (N_11835,N_10057,N_10328);
or U11836 (N_11836,N_10083,N_10112);
nor U11837 (N_11837,N_10247,N_10464);
or U11838 (N_11838,N_10424,N_10980);
and U11839 (N_11839,N_10453,N_10121);
and U11840 (N_11840,N_10868,N_10761);
nor U11841 (N_11841,N_10560,N_10564);
or U11842 (N_11842,N_10399,N_10014);
nand U11843 (N_11843,N_10941,N_10460);
xnor U11844 (N_11844,N_10336,N_10070);
nor U11845 (N_11845,N_10970,N_10894);
nand U11846 (N_11846,N_10852,N_10886);
and U11847 (N_11847,N_10133,N_10012);
or U11848 (N_11848,N_10296,N_10333);
and U11849 (N_11849,N_10604,N_10713);
nand U11850 (N_11850,N_10219,N_10372);
nor U11851 (N_11851,N_10552,N_10668);
and U11852 (N_11852,N_10490,N_10890);
or U11853 (N_11853,N_10029,N_10785);
and U11854 (N_11854,N_10625,N_10397);
or U11855 (N_11855,N_10542,N_10752);
nand U11856 (N_11856,N_10842,N_10778);
and U11857 (N_11857,N_10674,N_10040);
or U11858 (N_11858,N_10751,N_10318);
or U11859 (N_11859,N_10174,N_10383);
and U11860 (N_11860,N_10899,N_10675);
and U11861 (N_11861,N_10752,N_10155);
nor U11862 (N_11862,N_10732,N_10341);
or U11863 (N_11863,N_10980,N_10173);
or U11864 (N_11864,N_10732,N_10156);
xor U11865 (N_11865,N_10856,N_10787);
or U11866 (N_11866,N_10103,N_10901);
nor U11867 (N_11867,N_10889,N_10869);
nand U11868 (N_11868,N_10429,N_10754);
and U11869 (N_11869,N_10836,N_10375);
xor U11870 (N_11870,N_10750,N_10919);
nor U11871 (N_11871,N_10450,N_10197);
nand U11872 (N_11872,N_10102,N_10063);
xnor U11873 (N_11873,N_10170,N_10042);
xor U11874 (N_11874,N_10256,N_10497);
nor U11875 (N_11875,N_10068,N_10421);
and U11876 (N_11876,N_10881,N_10293);
or U11877 (N_11877,N_10037,N_10343);
or U11878 (N_11878,N_10646,N_10431);
xnor U11879 (N_11879,N_10064,N_10366);
nor U11880 (N_11880,N_10053,N_10942);
or U11881 (N_11881,N_10655,N_10565);
xor U11882 (N_11882,N_10521,N_10714);
or U11883 (N_11883,N_10046,N_10109);
nand U11884 (N_11884,N_10237,N_10393);
nor U11885 (N_11885,N_10367,N_10050);
xor U11886 (N_11886,N_10405,N_10156);
nand U11887 (N_11887,N_10740,N_10268);
or U11888 (N_11888,N_10177,N_10049);
nor U11889 (N_11889,N_10255,N_10876);
or U11890 (N_11890,N_10252,N_10605);
nand U11891 (N_11891,N_10534,N_10779);
nand U11892 (N_11892,N_10400,N_10820);
or U11893 (N_11893,N_10031,N_10923);
nand U11894 (N_11894,N_10872,N_10214);
xnor U11895 (N_11895,N_10621,N_10357);
and U11896 (N_11896,N_10155,N_10889);
and U11897 (N_11897,N_10547,N_10996);
nand U11898 (N_11898,N_10558,N_10259);
and U11899 (N_11899,N_10852,N_10008);
nand U11900 (N_11900,N_10311,N_10740);
and U11901 (N_11901,N_10348,N_10547);
nand U11902 (N_11902,N_10437,N_10661);
nand U11903 (N_11903,N_10632,N_10625);
nand U11904 (N_11904,N_10121,N_10025);
or U11905 (N_11905,N_10093,N_10961);
and U11906 (N_11906,N_10664,N_10793);
nor U11907 (N_11907,N_10257,N_10217);
nand U11908 (N_11908,N_10706,N_10837);
nand U11909 (N_11909,N_10932,N_10114);
and U11910 (N_11910,N_10038,N_10538);
and U11911 (N_11911,N_10979,N_10326);
xnor U11912 (N_11912,N_10516,N_10008);
and U11913 (N_11913,N_10540,N_10518);
xor U11914 (N_11914,N_10070,N_10549);
nor U11915 (N_11915,N_10855,N_10687);
nor U11916 (N_11916,N_10823,N_10194);
or U11917 (N_11917,N_10349,N_10666);
nand U11918 (N_11918,N_10087,N_10702);
nand U11919 (N_11919,N_10660,N_10163);
or U11920 (N_11920,N_10471,N_10033);
and U11921 (N_11921,N_10857,N_10854);
or U11922 (N_11922,N_10721,N_10928);
or U11923 (N_11923,N_10537,N_10683);
nor U11924 (N_11924,N_10514,N_10575);
nor U11925 (N_11925,N_10496,N_10264);
or U11926 (N_11926,N_10056,N_10980);
nand U11927 (N_11927,N_10659,N_10813);
or U11928 (N_11928,N_10157,N_10261);
nor U11929 (N_11929,N_10547,N_10582);
nand U11930 (N_11930,N_10610,N_10818);
and U11931 (N_11931,N_10214,N_10197);
nor U11932 (N_11932,N_10282,N_10039);
nand U11933 (N_11933,N_10541,N_10052);
nor U11934 (N_11934,N_10400,N_10398);
or U11935 (N_11935,N_10237,N_10832);
nor U11936 (N_11936,N_10838,N_10270);
and U11937 (N_11937,N_10875,N_10810);
and U11938 (N_11938,N_10757,N_10911);
or U11939 (N_11939,N_10795,N_10393);
nor U11940 (N_11940,N_10163,N_10759);
nand U11941 (N_11941,N_10769,N_10912);
and U11942 (N_11942,N_10584,N_10840);
xor U11943 (N_11943,N_10549,N_10466);
or U11944 (N_11944,N_10231,N_10623);
nor U11945 (N_11945,N_10809,N_10264);
nand U11946 (N_11946,N_10711,N_10614);
and U11947 (N_11947,N_10562,N_10864);
nand U11948 (N_11948,N_10655,N_10589);
nand U11949 (N_11949,N_10621,N_10470);
nor U11950 (N_11950,N_10454,N_10582);
or U11951 (N_11951,N_10169,N_10714);
or U11952 (N_11952,N_10889,N_10983);
and U11953 (N_11953,N_10080,N_10299);
or U11954 (N_11954,N_10098,N_10942);
or U11955 (N_11955,N_10407,N_10213);
or U11956 (N_11956,N_10576,N_10686);
or U11957 (N_11957,N_10725,N_10918);
nand U11958 (N_11958,N_10551,N_10665);
and U11959 (N_11959,N_10256,N_10818);
nand U11960 (N_11960,N_10956,N_10721);
and U11961 (N_11961,N_10970,N_10598);
and U11962 (N_11962,N_10341,N_10715);
nor U11963 (N_11963,N_10307,N_10582);
nor U11964 (N_11964,N_10949,N_10140);
nor U11965 (N_11965,N_10333,N_10554);
nor U11966 (N_11966,N_10100,N_10096);
nand U11967 (N_11967,N_10457,N_10128);
nand U11968 (N_11968,N_10367,N_10958);
nor U11969 (N_11969,N_10214,N_10456);
nand U11970 (N_11970,N_10828,N_10619);
or U11971 (N_11971,N_10253,N_10753);
nor U11972 (N_11972,N_10705,N_10459);
nor U11973 (N_11973,N_10636,N_10466);
nand U11974 (N_11974,N_10415,N_10309);
nand U11975 (N_11975,N_10695,N_10017);
nand U11976 (N_11976,N_10865,N_10180);
or U11977 (N_11977,N_10281,N_10396);
and U11978 (N_11978,N_10047,N_10418);
nand U11979 (N_11979,N_10155,N_10758);
nor U11980 (N_11980,N_10990,N_10252);
xor U11981 (N_11981,N_10824,N_10530);
or U11982 (N_11982,N_10176,N_10212);
or U11983 (N_11983,N_10710,N_10097);
or U11984 (N_11984,N_10315,N_10019);
nand U11985 (N_11985,N_10343,N_10894);
nor U11986 (N_11986,N_10010,N_10397);
nand U11987 (N_11987,N_10977,N_10990);
nor U11988 (N_11988,N_10795,N_10836);
nor U11989 (N_11989,N_10861,N_10183);
xor U11990 (N_11990,N_10598,N_10770);
nand U11991 (N_11991,N_10634,N_10158);
nor U11992 (N_11992,N_10440,N_10739);
nor U11993 (N_11993,N_10401,N_10827);
xor U11994 (N_11994,N_10897,N_10768);
nor U11995 (N_11995,N_10952,N_10430);
and U11996 (N_11996,N_10626,N_10817);
and U11997 (N_11997,N_10893,N_10870);
and U11998 (N_11998,N_10818,N_10079);
or U11999 (N_11999,N_10577,N_10360);
and U12000 (N_12000,N_11234,N_11208);
nor U12001 (N_12001,N_11500,N_11028);
nand U12002 (N_12002,N_11056,N_11720);
and U12003 (N_12003,N_11274,N_11979);
nor U12004 (N_12004,N_11092,N_11792);
and U12005 (N_12005,N_11745,N_11312);
or U12006 (N_12006,N_11818,N_11146);
and U12007 (N_12007,N_11664,N_11088);
and U12008 (N_12008,N_11996,N_11292);
nand U12009 (N_12009,N_11885,N_11364);
nor U12010 (N_12010,N_11330,N_11077);
nor U12011 (N_12011,N_11323,N_11660);
and U12012 (N_12012,N_11412,N_11756);
xor U12013 (N_12013,N_11398,N_11270);
nor U12014 (N_12014,N_11129,N_11573);
and U12015 (N_12015,N_11944,N_11509);
and U12016 (N_12016,N_11755,N_11052);
nor U12017 (N_12017,N_11566,N_11859);
and U12018 (N_12018,N_11237,N_11299);
nor U12019 (N_12019,N_11012,N_11327);
and U12020 (N_12020,N_11909,N_11184);
nor U12021 (N_12021,N_11383,N_11258);
and U12022 (N_12022,N_11157,N_11997);
xor U12023 (N_12023,N_11030,N_11005);
nor U12024 (N_12024,N_11222,N_11071);
xnor U12025 (N_12025,N_11356,N_11122);
and U12026 (N_12026,N_11160,N_11989);
and U12027 (N_12027,N_11911,N_11840);
and U12028 (N_12028,N_11953,N_11582);
xor U12029 (N_12029,N_11809,N_11023);
and U12030 (N_12030,N_11978,N_11605);
or U12031 (N_12031,N_11450,N_11279);
nand U12032 (N_12032,N_11864,N_11226);
or U12033 (N_12033,N_11457,N_11259);
or U12034 (N_12034,N_11073,N_11452);
nand U12035 (N_12035,N_11638,N_11317);
or U12036 (N_12036,N_11860,N_11281);
nor U12037 (N_12037,N_11812,N_11654);
or U12038 (N_12038,N_11882,N_11201);
or U12039 (N_12039,N_11109,N_11333);
nor U12040 (N_12040,N_11959,N_11414);
xor U12041 (N_12041,N_11928,N_11712);
and U12042 (N_12042,N_11851,N_11772);
nand U12043 (N_12043,N_11041,N_11729);
nor U12044 (N_12044,N_11103,N_11665);
nand U12045 (N_12045,N_11766,N_11986);
nand U12046 (N_12046,N_11326,N_11562);
or U12047 (N_12047,N_11114,N_11991);
nand U12048 (N_12048,N_11140,N_11421);
nor U12049 (N_12049,N_11767,N_11229);
or U12050 (N_12050,N_11040,N_11213);
and U12051 (N_12051,N_11010,N_11617);
and U12052 (N_12052,N_11974,N_11190);
and U12053 (N_12053,N_11725,N_11038);
nor U12054 (N_12054,N_11053,N_11607);
or U12055 (N_12055,N_11295,N_11531);
nor U12056 (N_12056,N_11194,N_11915);
nor U12057 (N_12057,N_11872,N_11212);
and U12058 (N_12058,N_11486,N_11446);
nand U12059 (N_12059,N_11940,N_11761);
or U12060 (N_12060,N_11062,N_11185);
nand U12061 (N_12061,N_11415,N_11656);
xnor U12062 (N_12062,N_11692,N_11130);
nand U12063 (N_12063,N_11425,N_11433);
nand U12064 (N_12064,N_11791,N_11522);
and U12065 (N_12065,N_11247,N_11080);
and U12066 (N_12066,N_11925,N_11018);
nand U12067 (N_12067,N_11104,N_11796);
and U12068 (N_12068,N_11847,N_11966);
and U12069 (N_12069,N_11139,N_11085);
or U12070 (N_12070,N_11900,N_11983);
and U12071 (N_12071,N_11307,N_11291);
and U12072 (N_12072,N_11701,N_11963);
nand U12073 (N_12073,N_11008,N_11138);
nand U12074 (N_12074,N_11144,N_11559);
or U12075 (N_12075,N_11225,N_11172);
or U12076 (N_12076,N_11802,N_11586);
nand U12077 (N_12077,N_11227,N_11126);
nand U12078 (N_12078,N_11434,N_11361);
nor U12079 (N_12079,N_11357,N_11055);
or U12080 (N_12080,N_11039,N_11666);
nand U12081 (N_12081,N_11496,N_11703);
nor U12082 (N_12082,N_11804,N_11154);
or U12083 (N_12083,N_11694,N_11454);
and U12084 (N_12084,N_11706,N_11595);
or U12085 (N_12085,N_11598,N_11527);
nand U12086 (N_12086,N_11969,N_11045);
or U12087 (N_12087,N_11111,N_11972);
and U12088 (N_12088,N_11752,N_11964);
or U12089 (N_12089,N_11492,N_11708);
or U12090 (N_12090,N_11485,N_11680);
and U12091 (N_12091,N_11675,N_11843);
nor U12092 (N_12092,N_11118,N_11453);
nor U12093 (N_12093,N_11475,N_11801);
xor U12094 (N_12094,N_11629,N_11494);
or U12095 (N_12095,N_11917,N_11945);
xor U12096 (N_12096,N_11596,N_11868);
or U12097 (N_12097,N_11774,N_11831);
and U12098 (N_12098,N_11856,N_11568);
nand U12099 (N_12099,N_11306,N_11006);
or U12100 (N_12100,N_11798,N_11137);
and U12101 (N_12101,N_11250,N_11193);
nand U12102 (N_12102,N_11423,N_11322);
nor U12103 (N_12103,N_11685,N_11519);
or U12104 (N_12104,N_11866,N_11621);
nor U12105 (N_12105,N_11839,N_11002);
and U12106 (N_12106,N_11921,N_11520);
nor U12107 (N_12107,N_11378,N_11702);
nor U12108 (N_12108,N_11417,N_11204);
and U12109 (N_12109,N_11777,N_11061);
or U12110 (N_12110,N_11123,N_11113);
nor U12111 (N_12111,N_11673,N_11100);
or U12112 (N_12112,N_11059,N_11167);
nor U12113 (N_12113,N_11047,N_11298);
and U12114 (N_12114,N_11913,N_11313);
or U12115 (N_12115,N_11112,N_11683);
nor U12116 (N_12116,N_11633,N_11411);
and U12117 (N_12117,N_11657,N_11624);
and U12118 (N_12118,N_11899,N_11143);
and U12119 (N_12119,N_11719,N_11558);
and U12120 (N_12120,N_11662,N_11120);
and U12121 (N_12121,N_11391,N_11387);
nand U12122 (N_12122,N_11310,N_11439);
and U12123 (N_12123,N_11099,N_11904);
or U12124 (N_12124,N_11700,N_11230);
nor U12125 (N_12125,N_11328,N_11858);
and U12126 (N_12126,N_11611,N_11579);
xnor U12127 (N_12127,N_11108,N_11233);
nand U12128 (N_12128,N_11181,N_11340);
xor U12129 (N_12129,N_11949,N_11263);
nor U12130 (N_12130,N_11783,N_11488);
nor U12131 (N_12131,N_11158,N_11141);
and U12132 (N_12132,N_11764,N_11183);
nand U12133 (N_12133,N_11058,N_11922);
and U12134 (N_12134,N_11553,N_11407);
and U12135 (N_12135,N_11554,N_11821);
and U12136 (N_12136,N_11516,N_11536);
nor U12137 (N_12137,N_11287,N_11739);
or U12138 (N_12138,N_11540,N_11093);
xnor U12139 (N_12139,N_11195,N_11630);
or U12140 (N_12140,N_11031,N_11399);
and U12141 (N_12141,N_11187,N_11360);
nor U12142 (N_12142,N_11395,N_11083);
or U12143 (N_12143,N_11174,N_11724);
or U12144 (N_12144,N_11029,N_11243);
nor U12145 (N_12145,N_11634,N_11737);
and U12146 (N_12146,N_11848,N_11314);
and U12147 (N_12147,N_11127,N_11881);
nor U12148 (N_12148,N_11479,N_11468);
and U12149 (N_12149,N_11884,N_11166);
nand U12150 (N_12150,N_11923,N_11875);
nand U12151 (N_12151,N_11749,N_11861);
nand U12152 (N_12152,N_11197,N_11723);
and U12153 (N_12153,N_11537,N_11511);
xnor U12154 (N_12154,N_11003,N_11982);
nor U12155 (N_12155,N_11602,N_11209);
and U12156 (N_12156,N_11240,N_11691);
or U12157 (N_12157,N_11797,N_11869);
nor U12158 (N_12158,N_11024,N_11939);
and U12159 (N_12159,N_11043,N_11987);
or U12160 (N_12160,N_11781,N_11615);
or U12161 (N_12161,N_11311,N_11060);
or U12162 (N_12162,N_11535,N_11569);
or U12163 (N_12163,N_11455,N_11202);
or U12164 (N_12164,N_11431,N_11710);
nor U12165 (N_12165,N_11348,N_11179);
nand U12166 (N_12166,N_11658,N_11806);
nand U12167 (N_12167,N_11510,N_11156);
or U12168 (N_12168,N_11319,N_11463);
nand U12169 (N_12169,N_11932,N_11929);
nand U12170 (N_12170,N_11625,N_11735);
nand U12171 (N_12171,N_11242,N_11854);
nand U12172 (N_12172,N_11564,N_11897);
and U12173 (N_12173,N_11275,N_11345);
or U12174 (N_12174,N_11013,N_11542);
nor U12175 (N_12175,N_11367,N_11763);
or U12176 (N_12176,N_11918,N_11272);
or U12177 (N_12177,N_11771,N_11693);
or U12178 (N_12178,N_11142,N_11366);
nand U12179 (N_12179,N_11663,N_11075);
xor U12180 (N_12180,N_11171,N_11779);
nor U12181 (N_12181,N_11462,N_11941);
and U12182 (N_12182,N_11355,N_11653);
or U12183 (N_12183,N_11970,N_11117);
nand U12184 (N_12184,N_11416,N_11521);
xnor U12185 (N_12185,N_11121,N_11526);
or U12186 (N_12186,N_11427,N_11042);
and U12187 (N_12187,N_11320,N_11684);
nand U12188 (N_12188,N_11159,N_11614);
xnor U12189 (N_12189,N_11722,N_11449);
nor U12190 (N_12190,N_11440,N_11539);
and U12191 (N_12191,N_11758,N_11682);
or U12192 (N_12192,N_11132,N_11493);
nor U12193 (N_12193,N_11035,N_11017);
or U12194 (N_12194,N_11760,N_11445);
nand U12195 (N_12195,N_11902,N_11943);
nand U12196 (N_12196,N_11740,N_11464);
xnor U12197 (N_12197,N_11089,N_11436);
nor U12198 (N_12198,N_11910,N_11402);
or U12199 (N_12199,N_11645,N_11577);
nand U12200 (N_12200,N_11068,N_11538);
and U12201 (N_12201,N_11955,N_11097);
or U12202 (N_12202,N_11381,N_11776);
nand U12203 (N_12203,N_11962,N_11200);
and U12204 (N_12204,N_11321,N_11473);
and U12205 (N_12205,N_11981,N_11704);
nand U12206 (N_12206,N_11186,N_11343);
nand U12207 (N_12207,N_11273,N_11458);
or U12208 (N_12208,N_11594,N_11618);
or U12209 (N_12209,N_11992,N_11841);
nor U12210 (N_12210,N_11775,N_11380);
xnor U12211 (N_12211,N_11846,N_11616);
and U12212 (N_12212,N_11968,N_11285);
nor U12213 (N_12213,N_11886,N_11971);
nor U12214 (N_12214,N_11529,N_11432);
xnor U12215 (N_12215,N_11613,N_11346);
or U12216 (N_12216,N_11773,N_11480);
nor U12217 (N_12217,N_11958,N_11671);
nor U12218 (N_12218,N_11852,N_11876);
nand U12219 (N_12219,N_11845,N_11246);
or U12220 (N_12220,N_11474,N_11072);
and U12221 (N_12221,N_11032,N_11561);
xor U12222 (N_12222,N_11823,N_11726);
and U12223 (N_12223,N_11189,N_11556);
nor U12224 (N_12224,N_11550,N_11895);
and U12225 (N_12225,N_11507,N_11620);
or U12226 (N_12226,N_11670,N_11857);
nand U12227 (N_12227,N_11107,N_11437);
or U12228 (N_12228,N_11094,N_11268);
xor U12229 (N_12229,N_11257,N_11021);
xor U12230 (N_12230,N_11125,N_11622);
or U12231 (N_12231,N_11495,N_11718);
xor U12232 (N_12232,N_11525,N_11297);
nand U12233 (N_12233,N_11549,N_11078);
nand U12234 (N_12234,N_11919,N_11905);
and U12235 (N_12235,N_11887,N_11467);
xnor U12236 (N_12236,N_11484,N_11736);
nand U12237 (N_12237,N_11309,N_11954);
nand U12238 (N_12238,N_11067,N_11908);
nand U12239 (N_12239,N_11177,N_11027);
or U12240 (N_12240,N_11590,N_11499);
or U12241 (N_12241,N_11588,N_11482);
nand U12242 (N_12242,N_11942,N_11961);
nor U12243 (N_12243,N_11667,N_11935);
or U12244 (N_12244,N_11661,N_11266);
and U12245 (N_12245,N_11920,N_11198);
and U12246 (N_12246,N_11235,N_11221);
or U12247 (N_12247,N_11151,N_11105);
or U12248 (N_12248,N_11228,N_11048);
or U12249 (N_12249,N_11512,N_11603);
nand U12250 (N_12250,N_11570,N_11397);
and U12251 (N_12251,N_11543,N_11822);
and U12252 (N_12252,N_11000,N_11074);
or U12253 (N_12253,N_11734,N_11370);
or U12254 (N_12254,N_11199,N_11359);
or U12255 (N_12255,N_11681,N_11571);
or U12256 (N_12256,N_11081,N_11191);
and U12257 (N_12257,N_11305,N_11517);
xnor U12258 (N_12258,N_11998,N_11049);
and U12259 (N_12259,N_11635,N_11523);
and U12260 (N_12260,N_11632,N_11363);
or U12261 (N_12261,N_11807,N_11051);
and U12262 (N_12262,N_11862,N_11502);
xnor U12263 (N_12263,N_11286,N_11178);
and U12264 (N_12264,N_11651,N_11057);
or U12265 (N_12265,N_11483,N_11557);
and U12266 (N_12266,N_11575,N_11747);
or U12267 (N_12267,N_11769,N_11342);
or U12268 (N_12268,N_11631,N_11254);
nand U12269 (N_12269,N_11255,N_11816);
or U12270 (N_12270,N_11296,N_11688);
and U12271 (N_12271,N_11064,N_11591);
and U12272 (N_12272,N_11789,N_11372);
or U12273 (N_12273,N_11608,N_11394);
or U12274 (N_12274,N_11863,N_11889);
or U12275 (N_12275,N_11820,N_11597);
or U12276 (N_12276,N_11552,N_11985);
nand U12277 (N_12277,N_11231,N_11344);
and U12278 (N_12278,N_11716,N_11612);
and U12279 (N_12279,N_11717,N_11341);
nand U12280 (N_12280,N_11335,N_11388);
and U12281 (N_12281,N_11481,N_11447);
or U12282 (N_12282,N_11528,N_11168);
or U12283 (N_12283,N_11169,N_11379);
nand U12284 (N_12284,N_11293,N_11547);
nor U12285 (N_12285,N_11371,N_11261);
or U12286 (N_12286,N_11995,N_11604);
xor U12287 (N_12287,N_11714,N_11686);
and U12288 (N_12288,N_11162,N_11757);
or U12289 (N_12289,N_11907,N_11659);
or U12290 (N_12290,N_11283,N_11980);
nor U12291 (N_12291,N_11689,N_11390);
nand U12292 (N_12292,N_11422,N_11192);
and U12293 (N_12293,N_11420,N_11046);
and U12294 (N_12294,N_11498,N_11903);
and U12295 (N_12295,N_11696,N_11106);
nor U12296 (N_12296,N_11419,N_11898);
and U12297 (N_12297,N_11084,N_11101);
and U12298 (N_12298,N_11515,N_11785);
nand U12299 (N_12299,N_11351,N_11265);
nor U12300 (N_12300,N_11581,N_11400);
and U12301 (N_12301,N_11838,N_11079);
and U12302 (N_12302,N_11477,N_11731);
nor U12303 (N_12303,N_11303,N_11513);
or U12304 (N_12304,N_11019,N_11891);
xnor U12305 (N_12305,N_11173,N_11377);
and U12306 (N_12306,N_11438,N_11965);
and U12307 (N_12307,N_11606,N_11548);
and U12308 (N_12308,N_11877,N_11946);
or U12309 (N_12309,N_11648,N_11076);
and U12310 (N_12310,N_11894,N_11728);
xnor U12311 (N_12311,N_11063,N_11241);
or U12312 (N_12312,N_11389,N_11832);
and U12313 (N_12313,N_11803,N_11698);
or U12314 (N_12314,N_11033,N_11644);
nand U12315 (N_12315,N_11135,N_11392);
xnor U12316 (N_12316,N_11124,N_11619);
nand U12317 (N_12317,N_11408,N_11679);
and U12318 (N_12318,N_11930,N_11182);
nand U12319 (N_12319,N_11034,N_11282);
nand U12320 (N_12320,N_11800,N_11396);
nand U12321 (N_12321,N_11460,N_11386);
xnor U12322 (N_12322,N_11338,N_11115);
nand U12323 (N_12323,N_11456,N_11461);
and U12324 (N_12324,N_11793,N_11251);
or U12325 (N_12325,N_11782,N_11469);
and U12326 (N_12326,N_11788,N_11136);
or U12327 (N_12327,N_11647,N_11196);
nor U12328 (N_12328,N_11170,N_11677);
or U12329 (N_12329,N_11950,N_11678);
nand U12330 (N_12330,N_11896,N_11478);
nor U12331 (N_12331,N_11880,N_11145);
or U12332 (N_12332,N_11238,N_11623);
nor U12333 (N_12333,N_11410,N_11426);
and U12334 (N_12334,N_11276,N_11655);
and U12335 (N_12335,N_11873,N_11765);
nor U12336 (N_12336,N_11727,N_11879);
nand U12337 (N_12337,N_11505,N_11826);
xor U12338 (N_12338,N_11428,N_11835);
nor U12339 (N_12339,N_11705,N_11837);
xor U12340 (N_12340,N_11459,N_11787);
nand U12341 (N_12341,N_11609,N_11715);
or U12342 (N_12342,N_11834,N_11207);
nand U12343 (N_12343,N_11874,N_11354);
nor U12344 (N_12344,N_11116,N_11811);
nor U12345 (N_12345,N_11646,N_11210);
or U12346 (N_12346,N_11795,N_11487);
nand U12347 (N_12347,N_11352,N_11813);
nand U12348 (N_12348,N_11302,N_11697);
nand U12349 (N_12349,N_11551,N_11278);
or U12350 (N_12350,N_11050,N_11133);
nand U12351 (N_12351,N_11730,N_11339);
nor U12352 (N_12352,N_11912,N_11336);
or U12353 (N_12353,N_11687,N_11574);
nor U12354 (N_12354,N_11376,N_11733);
or U12355 (N_12355,N_11743,N_11814);
nand U12356 (N_12356,N_11674,N_11290);
or U12357 (N_12357,N_11331,N_11096);
nand U12358 (N_12358,N_11260,N_11025);
or U12359 (N_12359,N_11750,N_11610);
xor U12360 (N_12360,N_11690,N_11090);
nor U12361 (N_12361,N_11435,N_11770);
nand U12362 (N_12362,N_11741,N_11709);
nand U12363 (N_12363,N_11871,N_11565);
nand U12364 (N_12364,N_11990,N_11784);
nand U12365 (N_12365,N_11640,N_11914);
nor U12366 (N_12366,N_11842,N_11824);
nand U12367 (N_12367,N_11036,N_11584);
xor U12368 (N_12368,N_11382,N_11707);
or U12369 (N_12369,N_11466,N_11748);
or U12370 (N_12370,N_11444,N_11828);
or U12371 (N_12371,N_11365,N_11065);
nor U12372 (N_12372,N_11218,N_11476);
and U12373 (N_12373,N_11593,N_11546);
nor U12374 (N_12374,N_11936,N_11161);
and U12375 (N_12375,N_11165,N_11927);
and U12376 (N_12376,N_11649,N_11150);
nor U12377 (N_12377,N_11799,N_11870);
or U12378 (N_12378,N_11855,N_11890);
xnor U12379 (N_12379,N_11497,N_11815);
nor U12380 (N_12380,N_11324,N_11180);
nor U12381 (N_12381,N_11626,N_11545);
nor U12382 (N_12382,N_11867,N_11451);
nand U12383 (N_12383,N_11406,N_11711);
nand U12384 (N_12384,N_11530,N_11514);
nor U12385 (N_12385,N_11587,N_11650);
nand U12386 (N_12386,N_11219,N_11128);
or U12387 (N_12387,N_11926,N_11284);
or U12388 (N_12388,N_11470,N_11347);
or U12389 (N_12389,N_11533,N_11636);
xnor U12390 (N_12390,N_11054,N_11424);
or U12391 (N_12391,N_11205,N_11224);
or U12392 (N_12392,N_11110,N_11069);
and U12393 (N_12393,N_11599,N_11931);
or U12394 (N_12394,N_11037,N_11506);
nand U12395 (N_12395,N_11742,N_11206);
xor U12396 (N_12396,N_11011,N_11746);
nor U12397 (N_12397,N_11368,N_11751);
or U12398 (N_12398,N_11153,N_11409);
nor U12399 (N_12399,N_11163,N_11504);
nor U12400 (N_12400,N_11131,N_11264);
nor U12401 (N_12401,N_11014,N_11374);
or U12402 (N_12402,N_11325,N_11541);
nor U12403 (N_12403,N_11288,N_11308);
nand U12404 (N_12404,N_11262,N_11999);
nor U12405 (N_12405,N_11952,N_11016);
nand U12406 (N_12406,N_11768,N_11589);
or U12407 (N_12407,N_11244,N_11350);
and U12408 (N_12408,N_11924,N_11975);
nand U12409 (N_12409,N_11713,N_11892);
and U12410 (N_12410,N_11967,N_11628);
or U12411 (N_12411,N_11300,N_11249);
nor U12412 (N_12412,N_11267,N_11009);
and U12413 (N_12413,N_11066,N_11015);
nand U12414 (N_12414,N_11937,N_11849);
or U12415 (N_12415,N_11534,N_11220);
nand U12416 (N_12416,N_11738,N_11349);
xnor U12417 (N_12417,N_11808,N_11429);
or U12418 (N_12418,N_11256,N_11413);
nand U12419 (N_12419,N_11091,N_11585);
nor U12420 (N_12420,N_11901,N_11836);
nand U12421 (N_12421,N_11087,N_11865);
nand U12422 (N_12422,N_11786,N_11956);
nor U12423 (N_12423,N_11933,N_11362);
or U12424 (N_12424,N_11906,N_11044);
or U12425 (N_12425,N_11393,N_11916);
and U12426 (N_12426,N_11639,N_11984);
and U12427 (N_12427,N_11642,N_11332);
or U12428 (N_12428,N_11252,N_11503);
xor U12429 (N_12429,N_11443,N_11304);
nand U12430 (N_12430,N_11947,N_11373);
nor U12431 (N_12431,N_11810,N_11676);
and U12432 (N_12432,N_11652,N_11794);
nand U12433 (N_12433,N_11501,N_11280);
nand U12434 (N_12434,N_11850,N_11418);
or U12435 (N_12435,N_11833,N_11442);
xor U12436 (N_12436,N_11223,N_11289);
nand U12437 (N_12437,N_11175,N_11819);
or U12438 (N_12438,N_11384,N_11544);
nand U12439 (N_12439,N_11369,N_11576);
nand U12440 (N_12440,N_11236,N_11277);
nor U12441 (N_12441,N_11778,N_11973);
nor U12442 (N_12442,N_11948,N_11938);
and U12443 (N_12443,N_11699,N_11441);
nand U12444 (N_12444,N_11893,N_11883);
and U12445 (N_12445,N_11853,N_11318);
xor U12446 (N_12446,N_11672,N_11215);
xnor U12447 (N_12447,N_11641,N_11994);
nor U12448 (N_12448,N_11600,N_11888);
nor U12449 (N_12449,N_11817,N_11560);
nand U12450 (N_12450,N_11508,N_11405);
and U12451 (N_12451,N_11578,N_11401);
nand U12452 (N_12452,N_11134,N_11721);
or U12453 (N_12453,N_11271,N_11164);
nand U12454 (N_12454,N_11524,N_11188);
nor U12455 (N_12455,N_11334,N_11301);
or U12456 (N_12456,N_11176,N_11098);
and U12457 (N_12457,N_11216,N_11026);
xnor U12458 (N_12458,N_11375,N_11957);
nor U12459 (N_12459,N_11627,N_11214);
and U12460 (N_12460,N_11001,N_11404);
and U12461 (N_12461,N_11465,N_11669);
and U12462 (N_12462,N_11753,N_11358);
nand U12463 (N_12463,N_11004,N_11329);
and U12464 (N_12464,N_11601,N_11472);
nor U12465 (N_12465,N_11239,N_11385);
nand U12466 (N_12466,N_11203,N_11430);
xor U12467 (N_12467,N_11643,N_11825);
nand U12468 (N_12468,N_11353,N_11020);
nor U12469 (N_12469,N_11572,N_11007);
and U12470 (N_12470,N_11294,N_11518);
xnor U12471 (N_12471,N_11082,N_11637);
nand U12472 (N_12472,N_11448,N_11934);
or U12473 (N_12473,N_11976,N_11403);
or U12474 (N_12474,N_11232,N_11759);
or U12475 (N_12475,N_11951,N_11248);
nand U12476 (N_12476,N_11829,N_11253);
xnor U12477 (N_12477,N_11668,N_11583);
nor U12478 (N_12478,N_11211,N_11316);
or U12479 (N_12479,N_11490,N_11532);
nor U12480 (N_12480,N_11155,N_11315);
xnor U12481 (N_12481,N_11780,N_11086);
xor U12482 (N_12482,N_11337,N_11269);
nand U12483 (N_12483,N_11471,N_11555);
xor U12484 (N_12484,N_11070,N_11762);
xor U12485 (N_12485,N_11827,N_11491);
nor U12486 (N_12486,N_11489,N_11790);
or U12487 (N_12487,N_11695,N_11960);
nor U12488 (N_12488,N_11148,N_11563);
and U12489 (N_12489,N_11022,N_11095);
nand U12490 (N_12490,N_11744,N_11102);
xor U12491 (N_12491,N_11149,N_11592);
nand U12492 (N_12492,N_11988,N_11844);
and U12493 (N_12493,N_11830,N_11993);
xor U12494 (N_12494,N_11878,N_11732);
and U12495 (N_12495,N_11217,N_11567);
nand U12496 (N_12496,N_11754,N_11152);
nand U12497 (N_12497,N_11580,N_11119);
or U12498 (N_12498,N_11147,N_11977);
nor U12499 (N_12499,N_11805,N_11245);
or U12500 (N_12500,N_11160,N_11973);
and U12501 (N_12501,N_11553,N_11916);
or U12502 (N_12502,N_11599,N_11132);
nor U12503 (N_12503,N_11751,N_11268);
nand U12504 (N_12504,N_11999,N_11383);
and U12505 (N_12505,N_11414,N_11670);
or U12506 (N_12506,N_11840,N_11883);
or U12507 (N_12507,N_11656,N_11741);
nor U12508 (N_12508,N_11577,N_11638);
nand U12509 (N_12509,N_11493,N_11637);
and U12510 (N_12510,N_11437,N_11365);
or U12511 (N_12511,N_11671,N_11227);
nand U12512 (N_12512,N_11589,N_11501);
and U12513 (N_12513,N_11182,N_11065);
nor U12514 (N_12514,N_11292,N_11706);
and U12515 (N_12515,N_11089,N_11217);
and U12516 (N_12516,N_11819,N_11245);
nand U12517 (N_12517,N_11021,N_11977);
or U12518 (N_12518,N_11496,N_11638);
nor U12519 (N_12519,N_11312,N_11383);
or U12520 (N_12520,N_11659,N_11861);
nand U12521 (N_12521,N_11620,N_11218);
or U12522 (N_12522,N_11897,N_11759);
xor U12523 (N_12523,N_11728,N_11345);
xnor U12524 (N_12524,N_11436,N_11602);
or U12525 (N_12525,N_11445,N_11914);
or U12526 (N_12526,N_11154,N_11386);
or U12527 (N_12527,N_11951,N_11151);
nand U12528 (N_12528,N_11120,N_11937);
nand U12529 (N_12529,N_11276,N_11216);
or U12530 (N_12530,N_11722,N_11992);
and U12531 (N_12531,N_11899,N_11432);
or U12532 (N_12532,N_11822,N_11491);
xor U12533 (N_12533,N_11678,N_11390);
or U12534 (N_12534,N_11576,N_11614);
and U12535 (N_12535,N_11138,N_11428);
or U12536 (N_12536,N_11205,N_11056);
or U12537 (N_12537,N_11282,N_11445);
nor U12538 (N_12538,N_11153,N_11859);
and U12539 (N_12539,N_11558,N_11271);
and U12540 (N_12540,N_11931,N_11809);
and U12541 (N_12541,N_11149,N_11300);
nor U12542 (N_12542,N_11068,N_11223);
or U12543 (N_12543,N_11245,N_11239);
and U12544 (N_12544,N_11584,N_11714);
nor U12545 (N_12545,N_11165,N_11678);
nor U12546 (N_12546,N_11463,N_11004);
xor U12547 (N_12547,N_11212,N_11947);
or U12548 (N_12548,N_11847,N_11597);
nand U12549 (N_12549,N_11890,N_11129);
nor U12550 (N_12550,N_11827,N_11829);
and U12551 (N_12551,N_11425,N_11272);
or U12552 (N_12552,N_11329,N_11413);
or U12553 (N_12553,N_11317,N_11949);
or U12554 (N_12554,N_11932,N_11996);
nand U12555 (N_12555,N_11713,N_11187);
nor U12556 (N_12556,N_11907,N_11354);
nand U12557 (N_12557,N_11415,N_11312);
nor U12558 (N_12558,N_11410,N_11539);
nand U12559 (N_12559,N_11876,N_11820);
nand U12560 (N_12560,N_11698,N_11581);
xor U12561 (N_12561,N_11034,N_11656);
nand U12562 (N_12562,N_11838,N_11747);
xnor U12563 (N_12563,N_11503,N_11678);
nor U12564 (N_12564,N_11877,N_11645);
or U12565 (N_12565,N_11990,N_11472);
nand U12566 (N_12566,N_11923,N_11602);
nand U12567 (N_12567,N_11058,N_11348);
and U12568 (N_12568,N_11573,N_11189);
xor U12569 (N_12569,N_11049,N_11746);
nand U12570 (N_12570,N_11173,N_11858);
nand U12571 (N_12571,N_11096,N_11988);
nand U12572 (N_12572,N_11784,N_11234);
and U12573 (N_12573,N_11776,N_11989);
nand U12574 (N_12574,N_11842,N_11096);
nor U12575 (N_12575,N_11472,N_11597);
or U12576 (N_12576,N_11080,N_11103);
nor U12577 (N_12577,N_11255,N_11340);
xnor U12578 (N_12578,N_11552,N_11264);
nor U12579 (N_12579,N_11797,N_11862);
xor U12580 (N_12580,N_11947,N_11282);
xor U12581 (N_12581,N_11704,N_11871);
xnor U12582 (N_12582,N_11060,N_11495);
and U12583 (N_12583,N_11672,N_11538);
and U12584 (N_12584,N_11084,N_11636);
xnor U12585 (N_12585,N_11616,N_11189);
nor U12586 (N_12586,N_11571,N_11708);
and U12587 (N_12587,N_11283,N_11888);
nor U12588 (N_12588,N_11845,N_11979);
and U12589 (N_12589,N_11313,N_11826);
xnor U12590 (N_12590,N_11676,N_11469);
or U12591 (N_12591,N_11798,N_11060);
and U12592 (N_12592,N_11633,N_11387);
nand U12593 (N_12593,N_11123,N_11265);
nor U12594 (N_12594,N_11595,N_11624);
or U12595 (N_12595,N_11090,N_11620);
or U12596 (N_12596,N_11706,N_11331);
xnor U12597 (N_12597,N_11056,N_11894);
nand U12598 (N_12598,N_11457,N_11541);
and U12599 (N_12599,N_11368,N_11448);
or U12600 (N_12600,N_11934,N_11526);
and U12601 (N_12601,N_11804,N_11278);
nand U12602 (N_12602,N_11425,N_11414);
nand U12603 (N_12603,N_11117,N_11941);
nor U12604 (N_12604,N_11855,N_11387);
xor U12605 (N_12605,N_11942,N_11799);
nor U12606 (N_12606,N_11475,N_11421);
xor U12607 (N_12607,N_11665,N_11400);
xnor U12608 (N_12608,N_11507,N_11398);
or U12609 (N_12609,N_11166,N_11953);
nor U12610 (N_12610,N_11385,N_11880);
nor U12611 (N_12611,N_11539,N_11126);
nand U12612 (N_12612,N_11408,N_11842);
nor U12613 (N_12613,N_11085,N_11595);
and U12614 (N_12614,N_11379,N_11700);
and U12615 (N_12615,N_11761,N_11667);
xnor U12616 (N_12616,N_11170,N_11448);
or U12617 (N_12617,N_11140,N_11852);
xnor U12618 (N_12618,N_11859,N_11092);
and U12619 (N_12619,N_11733,N_11230);
or U12620 (N_12620,N_11140,N_11516);
or U12621 (N_12621,N_11247,N_11430);
or U12622 (N_12622,N_11275,N_11608);
and U12623 (N_12623,N_11260,N_11115);
nor U12624 (N_12624,N_11099,N_11868);
nor U12625 (N_12625,N_11529,N_11290);
or U12626 (N_12626,N_11036,N_11130);
or U12627 (N_12627,N_11268,N_11063);
nor U12628 (N_12628,N_11762,N_11502);
nor U12629 (N_12629,N_11949,N_11260);
nor U12630 (N_12630,N_11010,N_11994);
and U12631 (N_12631,N_11024,N_11318);
and U12632 (N_12632,N_11518,N_11390);
and U12633 (N_12633,N_11992,N_11496);
or U12634 (N_12634,N_11110,N_11408);
nor U12635 (N_12635,N_11156,N_11885);
nor U12636 (N_12636,N_11999,N_11295);
nand U12637 (N_12637,N_11508,N_11916);
xnor U12638 (N_12638,N_11664,N_11069);
nand U12639 (N_12639,N_11460,N_11189);
nand U12640 (N_12640,N_11826,N_11688);
or U12641 (N_12641,N_11132,N_11631);
and U12642 (N_12642,N_11870,N_11428);
xor U12643 (N_12643,N_11570,N_11807);
nor U12644 (N_12644,N_11216,N_11620);
nor U12645 (N_12645,N_11710,N_11344);
and U12646 (N_12646,N_11547,N_11577);
and U12647 (N_12647,N_11174,N_11545);
and U12648 (N_12648,N_11842,N_11513);
and U12649 (N_12649,N_11046,N_11499);
nor U12650 (N_12650,N_11713,N_11847);
nand U12651 (N_12651,N_11817,N_11441);
and U12652 (N_12652,N_11624,N_11883);
nand U12653 (N_12653,N_11038,N_11228);
nand U12654 (N_12654,N_11792,N_11367);
nand U12655 (N_12655,N_11328,N_11311);
nand U12656 (N_12656,N_11676,N_11038);
nor U12657 (N_12657,N_11390,N_11986);
nor U12658 (N_12658,N_11395,N_11209);
nor U12659 (N_12659,N_11500,N_11376);
nor U12660 (N_12660,N_11212,N_11754);
or U12661 (N_12661,N_11868,N_11419);
or U12662 (N_12662,N_11690,N_11790);
nand U12663 (N_12663,N_11999,N_11587);
and U12664 (N_12664,N_11409,N_11615);
nor U12665 (N_12665,N_11157,N_11013);
or U12666 (N_12666,N_11143,N_11392);
or U12667 (N_12667,N_11083,N_11768);
nand U12668 (N_12668,N_11650,N_11814);
and U12669 (N_12669,N_11036,N_11910);
and U12670 (N_12670,N_11583,N_11144);
or U12671 (N_12671,N_11325,N_11995);
and U12672 (N_12672,N_11873,N_11736);
nand U12673 (N_12673,N_11351,N_11906);
nand U12674 (N_12674,N_11555,N_11805);
nor U12675 (N_12675,N_11822,N_11788);
and U12676 (N_12676,N_11086,N_11831);
nand U12677 (N_12677,N_11877,N_11363);
nor U12678 (N_12678,N_11715,N_11515);
nor U12679 (N_12679,N_11688,N_11168);
nor U12680 (N_12680,N_11403,N_11811);
nor U12681 (N_12681,N_11259,N_11825);
nor U12682 (N_12682,N_11183,N_11924);
xor U12683 (N_12683,N_11081,N_11350);
and U12684 (N_12684,N_11503,N_11090);
and U12685 (N_12685,N_11288,N_11838);
nand U12686 (N_12686,N_11187,N_11529);
or U12687 (N_12687,N_11783,N_11577);
nor U12688 (N_12688,N_11747,N_11782);
or U12689 (N_12689,N_11522,N_11653);
nand U12690 (N_12690,N_11146,N_11986);
and U12691 (N_12691,N_11588,N_11289);
or U12692 (N_12692,N_11503,N_11743);
nand U12693 (N_12693,N_11599,N_11731);
and U12694 (N_12694,N_11330,N_11010);
nand U12695 (N_12695,N_11074,N_11789);
nand U12696 (N_12696,N_11743,N_11368);
and U12697 (N_12697,N_11041,N_11518);
or U12698 (N_12698,N_11846,N_11394);
xnor U12699 (N_12699,N_11473,N_11219);
xor U12700 (N_12700,N_11679,N_11152);
or U12701 (N_12701,N_11099,N_11137);
or U12702 (N_12702,N_11479,N_11902);
xnor U12703 (N_12703,N_11233,N_11850);
or U12704 (N_12704,N_11600,N_11746);
and U12705 (N_12705,N_11203,N_11774);
xnor U12706 (N_12706,N_11823,N_11531);
and U12707 (N_12707,N_11061,N_11934);
nor U12708 (N_12708,N_11564,N_11706);
nor U12709 (N_12709,N_11038,N_11662);
or U12710 (N_12710,N_11099,N_11455);
nand U12711 (N_12711,N_11744,N_11226);
or U12712 (N_12712,N_11639,N_11930);
nand U12713 (N_12713,N_11964,N_11356);
and U12714 (N_12714,N_11029,N_11157);
or U12715 (N_12715,N_11836,N_11670);
or U12716 (N_12716,N_11288,N_11701);
nor U12717 (N_12717,N_11111,N_11713);
nor U12718 (N_12718,N_11771,N_11661);
xnor U12719 (N_12719,N_11782,N_11587);
and U12720 (N_12720,N_11825,N_11762);
and U12721 (N_12721,N_11346,N_11268);
nand U12722 (N_12722,N_11643,N_11281);
or U12723 (N_12723,N_11903,N_11186);
or U12724 (N_12724,N_11453,N_11261);
and U12725 (N_12725,N_11354,N_11964);
nand U12726 (N_12726,N_11228,N_11489);
nor U12727 (N_12727,N_11182,N_11335);
or U12728 (N_12728,N_11337,N_11411);
nand U12729 (N_12729,N_11930,N_11132);
nor U12730 (N_12730,N_11938,N_11858);
nor U12731 (N_12731,N_11757,N_11441);
or U12732 (N_12732,N_11045,N_11895);
nand U12733 (N_12733,N_11005,N_11236);
and U12734 (N_12734,N_11488,N_11417);
nor U12735 (N_12735,N_11500,N_11705);
and U12736 (N_12736,N_11666,N_11195);
nand U12737 (N_12737,N_11900,N_11274);
or U12738 (N_12738,N_11845,N_11743);
and U12739 (N_12739,N_11370,N_11020);
nor U12740 (N_12740,N_11582,N_11086);
and U12741 (N_12741,N_11473,N_11833);
or U12742 (N_12742,N_11249,N_11060);
or U12743 (N_12743,N_11291,N_11198);
or U12744 (N_12744,N_11020,N_11758);
and U12745 (N_12745,N_11943,N_11255);
or U12746 (N_12746,N_11367,N_11850);
nor U12747 (N_12747,N_11579,N_11460);
and U12748 (N_12748,N_11543,N_11773);
nor U12749 (N_12749,N_11818,N_11561);
and U12750 (N_12750,N_11827,N_11667);
xnor U12751 (N_12751,N_11615,N_11296);
or U12752 (N_12752,N_11841,N_11475);
or U12753 (N_12753,N_11741,N_11347);
nor U12754 (N_12754,N_11181,N_11753);
or U12755 (N_12755,N_11967,N_11893);
or U12756 (N_12756,N_11880,N_11397);
nor U12757 (N_12757,N_11878,N_11624);
and U12758 (N_12758,N_11918,N_11479);
nand U12759 (N_12759,N_11000,N_11970);
nor U12760 (N_12760,N_11959,N_11325);
and U12761 (N_12761,N_11976,N_11781);
or U12762 (N_12762,N_11398,N_11255);
nor U12763 (N_12763,N_11140,N_11386);
nor U12764 (N_12764,N_11367,N_11580);
or U12765 (N_12765,N_11792,N_11719);
nand U12766 (N_12766,N_11296,N_11761);
nor U12767 (N_12767,N_11862,N_11908);
xnor U12768 (N_12768,N_11391,N_11602);
nor U12769 (N_12769,N_11478,N_11840);
nor U12770 (N_12770,N_11416,N_11793);
and U12771 (N_12771,N_11316,N_11422);
or U12772 (N_12772,N_11154,N_11823);
and U12773 (N_12773,N_11161,N_11191);
nand U12774 (N_12774,N_11077,N_11505);
nor U12775 (N_12775,N_11531,N_11879);
or U12776 (N_12776,N_11621,N_11611);
nand U12777 (N_12777,N_11915,N_11582);
nor U12778 (N_12778,N_11288,N_11704);
nor U12779 (N_12779,N_11878,N_11119);
and U12780 (N_12780,N_11393,N_11260);
xnor U12781 (N_12781,N_11801,N_11028);
nor U12782 (N_12782,N_11900,N_11472);
or U12783 (N_12783,N_11084,N_11791);
or U12784 (N_12784,N_11626,N_11787);
and U12785 (N_12785,N_11490,N_11936);
or U12786 (N_12786,N_11346,N_11142);
or U12787 (N_12787,N_11292,N_11340);
or U12788 (N_12788,N_11570,N_11911);
xnor U12789 (N_12789,N_11717,N_11458);
nand U12790 (N_12790,N_11217,N_11066);
and U12791 (N_12791,N_11080,N_11438);
and U12792 (N_12792,N_11504,N_11354);
or U12793 (N_12793,N_11174,N_11454);
xnor U12794 (N_12794,N_11689,N_11936);
nand U12795 (N_12795,N_11609,N_11401);
and U12796 (N_12796,N_11582,N_11159);
or U12797 (N_12797,N_11824,N_11938);
and U12798 (N_12798,N_11220,N_11516);
xnor U12799 (N_12799,N_11380,N_11958);
nor U12800 (N_12800,N_11922,N_11728);
nand U12801 (N_12801,N_11111,N_11989);
or U12802 (N_12802,N_11127,N_11313);
xor U12803 (N_12803,N_11911,N_11306);
and U12804 (N_12804,N_11918,N_11211);
or U12805 (N_12805,N_11212,N_11018);
nor U12806 (N_12806,N_11378,N_11915);
xnor U12807 (N_12807,N_11615,N_11618);
nor U12808 (N_12808,N_11572,N_11756);
nor U12809 (N_12809,N_11940,N_11909);
or U12810 (N_12810,N_11128,N_11791);
and U12811 (N_12811,N_11178,N_11462);
and U12812 (N_12812,N_11936,N_11258);
nor U12813 (N_12813,N_11442,N_11080);
and U12814 (N_12814,N_11319,N_11373);
nand U12815 (N_12815,N_11061,N_11786);
and U12816 (N_12816,N_11771,N_11729);
or U12817 (N_12817,N_11627,N_11357);
nand U12818 (N_12818,N_11612,N_11634);
nand U12819 (N_12819,N_11757,N_11431);
or U12820 (N_12820,N_11058,N_11274);
nor U12821 (N_12821,N_11922,N_11046);
xor U12822 (N_12822,N_11031,N_11145);
nand U12823 (N_12823,N_11609,N_11664);
nor U12824 (N_12824,N_11926,N_11013);
nor U12825 (N_12825,N_11424,N_11465);
or U12826 (N_12826,N_11515,N_11916);
and U12827 (N_12827,N_11850,N_11343);
xnor U12828 (N_12828,N_11956,N_11789);
nand U12829 (N_12829,N_11185,N_11082);
nand U12830 (N_12830,N_11422,N_11551);
and U12831 (N_12831,N_11658,N_11107);
and U12832 (N_12832,N_11984,N_11082);
nand U12833 (N_12833,N_11316,N_11024);
or U12834 (N_12834,N_11566,N_11118);
xnor U12835 (N_12835,N_11415,N_11875);
nor U12836 (N_12836,N_11702,N_11516);
or U12837 (N_12837,N_11299,N_11604);
or U12838 (N_12838,N_11408,N_11317);
or U12839 (N_12839,N_11894,N_11179);
nor U12840 (N_12840,N_11913,N_11653);
nor U12841 (N_12841,N_11093,N_11714);
nand U12842 (N_12842,N_11468,N_11935);
nand U12843 (N_12843,N_11121,N_11426);
nor U12844 (N_12844,N_11442,N_11624);
nor U12845 (N_12845,N_11081,N_11021);
nor U12846 (N_12846,N_11931,N_11765);
nand U12847 (N_12847,N_11334,N_11550);
and U12848 (N_12848,N_11186,N_11491);
nand U12849 (N_12849,N_11562,N_11035);
nand U12850 (N_12850,N_11353,N_11266);
and U12851 (N_12851,N_11628,N_11959);
and U12852 (N_12852,N_11422,N_11717);
or U12853 (N_12853,N_11843,N_11797);
or U12854 (N_12854,N_11962,N_11095);
and U12855 (N_12855,N_11455,N_11173);
or U12856 (N_12856,N_11889,N_11065);
nand U12857 (N_12857,N_11255,N_11060);
or U12858 (N_12858,N_11067,N_11885);
nor U12859 (N_12859,N_11836,N_11469);
xor U12860 (N_12860,N_11182,N_11428);
and U12861 (N_12861,N_11035,N_11204);
xor U12862 (N_12862,N_11947,N_11800);
or U12863 (N_12863,N_11058,N_11152);
xnor U12864 (N_12864,N_11512,N_11893);
xor U12865 (N_12865,N_11805,N_11700);
or U12866 (N_12866,N_11209,N_11477);
or U12867 (N_12867,N_11766,N_11943);
nor U12868 (N_12868,N_11566,N_11025);
or U12869 (N_12869,N_11718,N_11351);
and U12870 (N_12870,N_11387,N_11061);
and U12871 (N_12871,N_11223,N_11436);
and U12872 (N_12872,N_11799,N_11647);
or U12873 (N_12873,N_11028,N_11851);
nor U12874 (N_12874,N_11510,N_11669);
xor U12875 (N_12875,N_11344,N_11889);
xor U12876 (N_12876,N_11179,N_11291);
and U12877 (N_12877,N_11410,N_11556);
or U12878 (N_12878,N_11978,N_11935);
or U12879 (N_12879,N_11179,N_11410);
nor U12880 (N_12880,N_11979,N_11364);
or U12881 (N_12881,N_11392,N_11251);
or U12882 (N_12882,N_11251,N_11862);
nand U12883 (N_12883,N_11809,N_11194);
nand U12884 (N_12884,N_11460,N_11764);
or U12885 (N_12885,N_11073,N_11301);
and U12886 (N_12886,N_11864,N_11699);
nor U12887 (N_12887,N_11866,N_11833);
and U12888 (N_12888,N_11680,N_11951);
and U12889 (N_12889,N_11424,N_11275);
nand U12890 (N_12890,N_11932,N_11692);
nand U12891 (N_12891,N_11925,N_11158);
and U12892 (N_12892,N_11126,N_11172);
nor U12893 (N_12893,N_11588,N_11410);
or U12894 (N_12894,N_11089,N_11434);
nand U12895 (N_12895,N_11986,N_11386);
or U12896 (N_12896,N_11065,N_11333);
xor U12897 (N_12897,N_11907,N_11290);
or U12898 (N_12898,N_11956,N_11062);
and U12899 (N_12899,N_11883,N_11516);
or U12900 (N_12900,N_11411,N_11966);
xnor U12901 (N_12901,N_11742,N_11745);
nor U12902 (N_12902,N_11000,N_11934);
nand U12903 (N_12903,N_11265,N_11142);
and U12904 (N_12904,N_11656,N_11851);
or U12905 (N_12905,N_11824,N_11032);
nand U12906 (N_12906,N_11615,N_11408);
or U12907 (N_12907,N_11122,N_11089);
and U12908 (N_12908,N_11548,N_11576);
nor U12909 (N_12909,N_11981,N_11113);
nor U12910 (N_12910,N_11709,N_11316);
and U12911 (N_12911,N_11459,N_11769);
nand U12912 (N_12912,N_11739,N_11641);
and U12913 (N_12913,N_11112,N_11745);
and U12914 (N_12914,N_11158,N_11873);
or U12915 (N_12915,N_11945,N_11372);
nand U12916 (N_12916,N_11087,N_11950);
and U12917 (N_12917,N_11945,N_11723);
xnor U12918 (N_12918,N_11910,N_11309);
xor U12919 (N_12919,N_11586,N_11877);
nor U12920 (N_12920,N_11128,N_11089);
and U12921 (N_12921,N_11051,N_11657);
and U12922 (N_12922,N_11104,N_11969);
nor U12923 (N_12923,N_11837,N_11482);
and U12924 (N_12924,N_11672,N_11163);
nor U12925 (N_12925,N_11313,N_11373);
or U12926 (N_12926,N_11348,N_11595);
nand U12927 (N_12927,N_11126,N_11312);
or U12928 (N_12928,N_11342,N_11446);
xnor U12929 (N_12929,N_11497,N_11663);
or U12930 (N_12930,N_11347,N_11327);
nand U12931 (N_12931,N_11656,N_11165);
nand U12932 (N_12932,N_11648,N_11138);
xor U12933 (N_12933,N_11883,N_11475);
or U12934 (N_12934,N_11735,N_11910);
nand U12935 (N_12935,N_11988,N_11235);
or U12936 (N_12936,N_11023,N_11721);
and U12937 (N_12937,N_11216,N_11440);
or U12938 (N_12938,N_11627,N_11863);
and U12939 (N_12939,N_11743,N_11313);
nand U12940 (N_12940,N_11598,N_11278);
nand U12941 (N_12941,N_11767,N_11216);
nand U12942 (N_12942,N_11437,N_11900);
nor U12943 (N_12943,N_11654,N_11264);
and U12944 (N_12944,N_11712,N_11719);
and U12945 (N_12945,N_11855,N_11841);
or U12946 (N_12946,N_11383,N_11413);
xor U12947 (N_12947,N_11822,N_11719);
nor U12948 (N_12948,N_11671,N_11041);
and U12949 (N_12949,N_11734,N_11913);
nor U12950 (N_12950,N_11440,N_11283);
and U12951 (N_12951,N_11565,N_11859);
or U12952 (N_12952,N_11767,N_11185);
or U12953 (N_12953,N_11609,N_11794);
and U12954 (N_12954,N_11955,N_11846);
nor U12955 (N_12955,N_11637,N_11365);
or U12956 (N_12956,N_11563,N_11470);
nand U12957 (N_12957,N_11853,N_11276);
nor U12958 (N_12958,N_11809,N_11748);
and U12959 (N_12959,N_11479,N_11448);
or U12960 (N_12960,N_11088,N_11004);
nor U12961 (N_12961,N_11782,N_11044);
and U12962 (N_12962,N_11111,N_11303);
and U12963 (N_12963,N_11319,N_11630);
nand U12964 (N_12964,N_11617,N_11968);
or U12965 (N_12965,N_11171,N_11595);
nand U12966 (N_12966,N_11470,N_11397);
and U12967 (N_12967,N_11344,N_11773);
xor U12968 (N_12968,N_11262,N_11098);
and U12969 (N_12969,N_11330,N_11087);
and U12970 (N_12970,N_11123,N_11752);
xor U12971 (N_12971,N_11817,N_11367);
or U12972 (N_12972,N_11397,N_11080);
nand U12973 (N_12973,N_11660,N_11593);
nor U12974 (N_12974,N_11024,N_11227);
nand U12975 (N_12975,N_11490,N_11127);
or U12976 (N_12976,N_11128,N_11245);
nor U12977 (N_12977,N_11429,N_11534);
and U12978 (N_12978,N_11999,N_11237);
and U12979 (N_12979,N_11285,N_11133);
nand U12980 (N_12980,N_11761,N_11731);
nor U12981 (N_12981,N_11593,N_11995);
or U12982 (N_12982,N_11405,N_11251);
or U12983 (N_12983,N_11569,N_11062);
nor U12984 (N_12984,N_11177,N_11732);
or U12985 (N_12985,N_11414,N_11119);
or U12986 (N_12986,N_11558,N_11784);
nor U12987 (N_12987,N_11312,N_11286);
or U12988 (N_12988,N_11536,N_11160);
nor U12989 (N_12989,N_11193,N_11430);
and U12990 (N_12990,N_11095,N_11894);
nor U12991 (N_12991,N_11481,N_11008);
nor U12992 (N_12992,N_11775,N_11596);
xnor U12993 (N_12993,N_11457,N_11786);
xnor U12994 (N_12994,N_11647,N_11612);
nand U12995 (N_12995,N_11453,N_11777);
nand U12996 (N_12996,N_11097,N_11848);
nand U12997 (N_12997,N_11699,N_11509);
nand U12998 (N_12998,N_11447,N_11388);
and U12999 (N_12999,N_11812,N_11567);
and U13000 (N_13000,N_12187,N_12495);
and U13001 (N_13001,N_12227,N_12288);
nor U13002 (N_13002,N_12353,N_12253);
or U13003 (N_13003,N_12304,N_12399);
nand U13004 (N_13004,N_12238,N_12844);
nand U13005 (N_13005,N_12568,N_12015);
nand U13006 (N_13006,N_12664,N_12791);
and U13007 (N_13007,N_12979,N_12872);
and U13008 (N_13008,N_12051,N_12684);
nand U13009 (N_13009,N_12333,N_12340);
nor U13010 (N_13010,N_12052,N_12858);
nand U13011 (N_13011,N_12726,N_12958);
xnor U13012 (N_13012,N_12870,N_12005);
xnor U13013 (N_13013,N_12910,N_12632);
nor U13014 (N_13014,N_12907,N_12072);
nand U13015 (N_13015,N_12433,N_12714);
and U13016 (N_13016,N_12836,N_12258);
or U13017 (N_13017,N_12670,N_12554);
nand U13018 (N_13018,N_12219,N_12257);
nor U13019 (N_13019,N_12633,N_12742);
nand U13020 (N_13020,N_12502,N_12161);
nand U13021 (N_13021,N_12044,N_12553);
and U13022 (N_13022,N_12600,N_12056);
nand U13023 (N_13023,N_12454,N_12816);
nand U13024 (N_13024,N_12375,N_12681);
or U13025 (N_13025,N_12099,N_12203);
nand U13026 (N_13026,N_12496,N_12416);
or U13027 (N_13027,N_12316,N_12149);
or U13028 (N_13028,N_12107,N_12384);
nor U13029 (N_13029,N_12699,N_12050);
nand U13030 (N_13030,N_12271,N_12727);
nor U13031 (N_13031,N_12901,N_12960);
and U13032 (N_13032,N_12508,N_12482);
and U13033 (N_13033,N_12248,N_12711);
nor U13034 (N_13034,N_12693,N_12522);
and U13035 (N_13035,N_12669,N_12178);
or U13036 (N_13036,N_12543,N_12045);
and U13037 (N_13037,N_12725,N_12467);
or U13038 (N_13038,N_12860,N_12087);
and U13039 (N_13039,N_12940,N_12041);
and U13040 (N_13040,N_12426,N_12499);
nor U13041 (N_13041,N_12010,N_12127);
or U13042 (N_13042,N_12710,N_12410);
nor U13043 (N_13043,N_12446,N_12067);
nand U13044 (N_13044,N_12878,N_12953);
and U13045 (N_13045,N_12401,N_12436);
nand U13046 (N_13046,N_12671,N_12829);
or U13047 (N_13047,N_12284,N_12898);
nand U13048 (N_13048,N_12552,N_12945);
xor U13049 (N_13049,N_12623,N_12466);
nor U13050 (N_13050,N_12130,N_12046);
nor U13051 (N_13051,N_12705,N_12639);
or U13052 (N_13052,N_12515,N_12166);
nand U13053 (N_13053,N_12473,N_12272);
nor U13054 (N_13054,N_12477,N_12925);
or U13055 (N_13055,N_12199,N_12246);
and U13056 (N_13056,N_12438,N_12922);
and U13057 (N_13057,N_12776,N_12141);
and U13058 (N_13058,N_12027,N_12255);
nor U13059 (N_13059,N_12692,N_12789);
nor U13060 (N_13060,N_12819,N_12704);
nand U13061 (N_13061,N_12479,N_12345);
and U13062 (N_13062,N_12205,N_12174);
and U13063 (N_13063,N_12407,N_12905);
and U13064 (N_13064,N_12900,N_12531);
and U13065 (N_13065,N_12882,N_12969);
nor U13066 (N_13066,N_12212,N_12064);
and U13067 (N_13067,N_12920,N_12579);
nor U13068 (N_13068,N_12456,N_12625);
and U13069 (N_13069,N_12190,N_12786);
and U13070 (N_13070,N_12757,N_12621);
nand U13071 (N_13071,N_12852,N_12546);
nor U13072 (N_13072,N_12790,N_12525);
nor U13073 (N_13073,N_12817,N_12528);
nor U13074 (N_13074,N_12465,N_12128);
or U13075 (N_13075,N_12042,N_12291);
xor U13076 (N_13076,N_12468,N_12570);
nor U13077 (N_13077,N_12631,N_12730);
or U13078 (N_13078,N_12023,N_12311);
nor U13079 (N_13079,N_12832,N_12105);
or U13080 (N_13080,N_12779,N_12302);
xor U13081 (N_13081,N_12748,N_12142);
nor U13082 (N_13082,N_12124,N_12767);
or U13083 (N_13083,N_12307,N_12551);
nor U13084 (N_13084,N_12285,N_12521);
nand U13085 (N_13085,N_12497,N_12157);
or U13086 (N_13086,N_12108,N_12722);
nor U13087 (N_13087,N_12924,N_12651);
xnor U13088 (N_13088,N_12873,N_12923);
nor U13089 (N_13089,N_12662,N_12047);
nor U13090 (N_13090,N_12063,N_12918);
or U13091 (N_13091,N_12618,N_12169);
nand U13092 (N_13092,N_12950,N_12524);
nand U13093 (N_13093,N_12626,N_12665);
and U13094 (N_13094,N_12392,N_12787);
nor U13095 (N_13095,N_12777,N_12721);
nand U13096 (N_13096,N_12491,N_12912);
or U13097 (N_13097,N_12752,N_12661);
or U13098 (N_13098,N_12598,N_12961);
or U13099 (N_13099,N_12332,N_12514);
and U13100 (N_13100,N_12241,N_12480);
nand U13101 (N_13101,N_12887,N_12507);
or U13102 (N_13102,N_12509,N_12442);
or U13103 (N_13103,N_12987,N_12697);
nor U13104 (N_13104,N_12996,N_12782);
nand U13105 (N_13105,N_12739,N_12354);
or U13106 (N_13106,N_12372,N_12327);
nor U13107 (N_13107,N_12755,N_12619);
and U13108 (N_13108,N_12716,N_12040);
and U13109 (N_13109,N_12139,N_12440);
nor U13110 (N_13110,N_12298,N_12013);
or U13111 (N_13111,N_12245,N_12098);
and U13112 (N_13112,N_12445,N_12305);
nor U13113 (N_13113,N_12695,N_12158);
xnor U13114 (N_13114,N_12523,N_12562);
nor U13115 (N_13115,N_12628,N_12207);
nor U13116 (N_13116,N_12059,N_12415);
nand U13117 (N_13117,N_12113,N_12053);
or U13118 (N_13118,N_12388,N_12629);
and U13119 (N_13119,N_12864,N_12679);
xnor U13120 (N_13120,N_12537,N_12191);
and U13121 (N_13121,N_12949,N_12989);
nand U13122 (N_13122,N_12983,N_12718);
and U13123 (N_13123,N_12772,N_12688);
or U13124 (N_13124,N_12432,N_12137);
nand U13125 (N_13125,N_12549,N_12380);
nor U13126 (N_13126,N_12602,N_12492);
nor U13127 (N_13127,N_12303,N_12608);
xor U13128 (N_13128,N_12261,N_12797);
nand U13129 (N_13129,N_12642,N_12186);
nor U13130 (N_13130,N_12657,N_12247);
nand U13131 (N_13131,N_12076,N_12250);
or U13132 (N_13132,N_12315,N_12706);
and U13133 (N_13133,N_12453,N_12656);
nor U13134 (N_13134,N_12096,N_12545);
or U13135 (N_13135,N_12418,N_12588);
and U13136 (N_13136,N_12249,N_12361);
nor U13137 (N_13137,N_12982,N_12812);
nor U13138 (N_13138,N_12532,N_12323);
nand U13139 (N_13139,N_12820,N_12260);
nor U13140 (N_13140,N_12999,N_12017);
and U13141 (N_13141,N_12848,N_12377);
nor U13142 (N_13142,N_12559,N_12796);
or U13143 (N_13143,N_12390,N_12992);
nor U13144 (N_13144,N_12609,N_12743);
or U13145 (N_13145,N_12172,N_12421);
and U13146 (N_13146,N_12188,N_12037);
nor U13147 (N_13147,N_12935,N_12338);
nand U13148 (N_13148,N_12685,N_12703);
nand U13149 (N_13149,N_12266,N_12165);
or U13150 (N_13150,N_12022,N_12262);
and U13151 (N_13151,N_12863,N_12004);
or U13152 (N_13152,N_12610,N_12753);
or U13153 (N_13153,N_12118,N_12398);
nand U13154 (N_13154,N_12798,N_12036);
nor U13155 (N_13155,N_12318,N_12897);
nor U13156 (N_13156,N_12917,N_12823);
and U13157 (N_13157,N_12673,N_12460);
nand U13158 (N_13158,N_12694,N_12210);
and U13159 (N_13159,N_12228,N_12264);
nor U13160 (N_13160,N_12648,N_12014);
nand U13161 (N_13161,N_12846,N_12385);
or U13162 (N_13162,N_12234,N_12397);
and U13163 (N_13163,N_12117,N_12556);
xor U13164 (N_13164,N_12908,N_12675);
nand U13165 (N_13165,N_12993,N_12696);
nand U13166 (N_13166,N_12963,N_12955);
or U13167 (N_13167,N_12344,N_12198);
and U13168 (N_13168,N_12254,N_12206);
xor U13169 (N_13169,N_12538,N_12075);
and U13170 (N_13170,N_12484,N_12069);
and U13171 (N_13171,N_12707,N_12874);
and U13172 (N_13172,N_12313,N_12194);
nor U13173 (N_13173,N_12712,N_12932);
or U13174 (N_13174,N_12400,N_12270);
nand U13175 (N_13175,N_12571,N_12815);
or U13176 (N_13176,N_12283,N_12849);
nor U13177 (N_13177,N_12810,N_12183);
or U13178 (N_13178,N_12309,N_12273);
nand U13179 (N_13179,N_12857,N_12282);
nor U13180 (N_13180,N_12801,N_12404);
nor U13181 (N_13181,N_12594,N_12181);
or U13182 (N_13182,N_12599,N_12913);
or U13183 (N_13183,N_12342,N_12991);
nand U13184 (N_13184,N_12434,N_12483);
nand U13185 (N_13185,N_12214,N_12615);
or U13186 (N_13186,N_12737,N_12038);
or U13187 (N_13187,N_12474,N_12411);
and U13188 (N_13188,N_12109,N_12176);
or U13189 (N_13189,N_12966,N_12448);
nand U13190 (N_13190,N_12487,N_12222);
nand U13191 (N_13191,N_12121,N_12175);
and U13192 (N_13192,N_12463,N_12869);
nand U13193 (N_13193,N_12855,N_12567);
nor U13194 (N_13194,N_12605,N_12564);
and U13195 (N_13195,N_12529,N_12114);
or U13196 (N_13196,N_12833,N_12321);
or U13197 (N_13197,N_12211,N_12256);
and U13198 (N_13198,N_12363,N_12825);
and U13199 (N_13199,N_12083,N_12702);
and U13200 (N_13200,N_12209,N_12906);
xor U13201 (N_13201,N_12613,N_12091);
and U13202 (N_13202,N_12640,N_12731);
nor U13203 (N_13203,N_12837,N_12417);
nand U13204 (N_13204,N_12563,N_12217);
nand U13205 (N_13205,N_12814,N_12152);
or U13206 (N_13206,N_12242,N_12676);
and U13207 (N_13207,N_12638,N_12319);
or U13208 (N_13208,N_12542,N_12896);
nand U13209 (N_13209,N_12019,N_12429);
nand U13210 (N_13210,N_12376,N_12252);
nor U13211 (N_13211,N_12539,N_12308);
nor U13212 (N_13212,N_12971,N_12208);
and U13213 (N_13213,N_12572,N_12503);
and U13214 (N_13214,N_12799,N_12856);
and U13215 (N_13215,N_12589,N_12422);
nand U13216 (N_13216,N_12151,N_12182);
or U13217 (N_13217,N_12895,N_12348);
or U13218 (N_13218,N_12978,N_12011);
xnor U13219 (N_13219,N_12795,N_12455);
nand U13220 (N_13220,N_12775,N_12140);
nor U13221 (N_13221,N_12170,N_12359);
nor U13222 (N_13222,N_12667,N_12173);
nor U13223 (N_13223,N_12061,N_12343);
nor U13224 (N_13224,N_12754,N_12143);
or U13225 (N_13225,N_12634,N_12092);
nor U13226 (N_13226,N_12736,N_12202);
and U13227 (N_13227,N_12746,N_12367);
xor U13228 (N_13228,N_12698,N_12070);
and U13229 (N_13229,N_12469,N_12781);
xnor U13230 (N_13230,N_12513,N_12942);
nand U13231 (N_13231,N_12148,N_12948);
nor U13232 (N_13232,N_12947,N_12557);
and U13233 (N_13233,N_12998,N_12094);
nor U13234 (N_13234,N_12120,N_12106);
and U13235 (N_13235,N_12095,N_12592);
and U13236 (N_13236,N_12396,N_12678);
nor U13237 (N_13237,N_12000,N_12723);
or U13238 (N_13238,N_12437,N_12603);
and U13239 (N_13239,N_12994,N_12216);
nand U13240 (N_13240,N_12689,N_12079);
nor U13241 (N_13241,N_12624,N_12197);
and U13242 (N_13242,N_12735,N_12885);
nand U13243 (N_13243,N_12180,N_12881);
nand U13244 (N_13244,N_12902,N_12290);
and U13245 (N_13245,N_12876,N_12773);
nand U13246 (N_13246,N_12066,N_12007);
nor U13247 (N_13247,N_12459,N_12065);
xor U13248 (N_13248,N_12530,N_12792);
or U13249 (N_13249,N_12936,N_12793);
nor U13250 (N_13250,N_12035,N_12871);
nand U13251 (N_13251,N_12766,N_12462);
or U13252 (N_13252,N_12774,N_12221);
or U13253 (N_13253,N_12803,N_12494);
or U13254 (N_13254,N_12709,N_12831);
nor U13255 (N_13255,N_12974,N_12604);
and U13256 (N_13256,N_12297,N_12607);
or U13257 (N_13257,N_12805,N_12593);
nor U13258 (N_13258,N_12393,N_12566);
nor U13259 (N_13259,N_12850,N_12826);
nor U13260 (N_13260,N_12237,N_12511);
nor U13261 (N_13261,N_12813,N_12759);
nand U13262 (N_13262,N_12548,N_12637);
and U13263 (N_13263,N_12547,N_12403);
and U13264 (N_13264,N_12541,N_12420);
xnor U13265 (N_13265,N_12841,N_12189);
xor U13266 (N_13266,N_12500,N_12928);
and U13267 (N_13267,N_12365,N_12575);
nor U13268 (N_13268,N_12439,N_12893);
xor U13269 (N_13269,N_12488,N_12478);
xnor U13270 (N_13270,N_12569,N_12449);
xor U13271 (N_13271,N_12682,N_12006);
and U13272 (N_13272,N_12761,N_12374);
or U13273 (N_13273,N_12658,N_12030);
nand U13274 (N_13274,N_12171,N_12464);
nand U13275 (N_13275,N_12879,N_12962);
xnor U13276 (N_13276,N_12904,N_12251);
and U13277 (N_13277,N_12104,N_12026);
or U13278 (N_13278,N_12110,N_12576);
xor U13279 (N_13279,N_12389,N_12144);
nor U13280 (N_13280,N_12715,N_12690);
nand U13281 (N_13281,N_12235,N_12101);
nor U13282 (N_13282,N_12341,N_12233);
or U13283 (N_13283,N_12031,N_12926);
nor U13284 (N_13284,N_12423,N_12585);
or U13285 (N_13285,N_12164,N_12506);
xnor U13286 (N_13286,N_12074,N_12977);
and U13287 (N_13287,N_12984,N_12859);
and U13288 (N_13288,N_12891,N_12163);
or U13289 (N_13289,N_12630,N_12424);
nand U13290 (N_13290,N_12830,N_12965);
nor U13291 (N_13291,N_12352,N_12744);
nand U13292 (N_13292,N_12560,N_12314);
and U13293 (N_13293,N_12934,N_12299);
nand U13294 (N_13294,N_12154,N_12324);
nand U13295 (N_13295,N_12583,N_12058);
and U13296 (N_13296,N_12601,N_12929);
nor U13297 (N_13297,N_12783,N_12584);
or U13298 (N_13298,N_12890,N_12225);
nand U13299 (N_13299,N_12077,N_12339);
or U13300 (N_13300,N_12750,N_12724);
and U13301 (N_13301,N_12627,N_12756);
nor U13302 (N_13302,N_12865,N_12230);
nand U13303 (N_13303,N_12636,N_12889);
nor U13304 (N_13304,N_12822,N_12741);
nor U13305 (N_13305,N_12119,N_12071);
nor U13306 (N_13306,N_12847,N_12195);
xnor U13307 (N_13307,N_12867,N_12485);
or U13308 (N_13308,N_12135,N_12024);
nand U13309 (N_13309,N_12168,N_12880);
or U13310 (N_13310,N_12443,N_12884);
or U13311 (N_13311,N_12921,N_12738);
or U13312 (N_13312,N_12360,N_12103);
nor U13313 (N_13313,N_12888,N_12807);
nor U13314 (N_13314,N_12719,N_12294);
or U13315 (N_13315,N_12177,N_12957);
xnor U13316 (N_13316,N_12780,N_12854);
or U13317 (N_13317,N_12419,N_12806);
nand U13318 (N_13318,N_12328,N_12371);
nand U13319 (N_13319,N_12020,N_12193);
nor U13320 (N_13320,N_12581,N_12184);
xnor U13321 (N_13321,N_12268,N_12663);
and U13322 (N_13322,N_12580,N_12201);
or U13323 (N_13323,N_12534,N_12116);
nand U13324 (N_13324,N_12018,N_12431);
nand U13325 (N_13325,N_12461,N_12391);
nand U13326 (N_13326,N_12808,N_12196);
and U13327 (N_13327,N_12862,N_12842);
and U13328 (N_13328,N_12160,N_12062);
and U13329 (N_13329,N_12931,N_12972);
nor U13330 (N_13330,N_12911,N_12645);
nor U13331 (N_13331,N_12526,N_12281);
xnor U13332 (N_13332,N_12244,N_12312);
nor U13333 (N_13333,N_12951,N_12100);
nor U13334 (N_13334,N_12717,N_12090);
nand U13335 (N_13335,N_12734,N_12012);
or U13336 (N_13336,N_12335,N_12520);
and U13337 (N_13337,N_12555,N_12561);
and U13338 (N_13338,N_12591,N_12112);
xor U13339 (N_13339,N_12330,N_12747);
nor U13340 (N_13340,N_12668,N_12296);
nand U13341 (N_13341,N_12350,N_12387);
xnor U13342 (N_13342,N_12596,N_12574);
and U13343 (N_13343,N_12544,N_12068);
nand U13344 (N_13344,N_12125,N_12278);
nand U13345 (N_13345,N_12078,N_12956);
xor U13346 (N_13346,N_12644,N_12954);
nor U13347 (N_13347,N_12927,N_12686);
nor U13348 (N_13348,N_12851,N_12622);
and U13349 (N_13349,N_12519,N_12666);
and U13350 (N_13350,N_12381,N_12995);
nor U13351 (N_13351,N_12489,N_12336);
or U13352 (N_13352,N_12606,N_12232);
nand U13353 (N_13353,N_12729,N_12586);
nand U13354 (N_13354,N_12276,N_12740);
and U13355 (N_13355,N_12617,N_12952);
nand U13356 (N_13356,N_12370,N_12728);
or U13357 (N_13357,N_12827,N_12368);
or U13358 (N_13358,N_12840,N_12732);
and U13359 (N_13359,N_12086,N_12029);
or U13360 (N_13360,N_12226,N_12301);
nor U13361 (N_13361,N_12768,N_12771);
or U13362 (N_13362,N_12239,N_12647);
nand U13363 (N_13363,N_12973,N_12909);
or U13364 (N_13364,N_12369,N_12941);
or U13365 (N_13365,N_12213,N_12408);
and U13366 (N_13366,N_12649,N_12981);
or U13367 (N_13367,N_12131,N_12153);
nor U13368 (N_13368,N_12259,N_12620);
and U13369 (N_13369,N_12654,N_12573);
xnor U13370 (N_13370,N_12527,N_12025);
nor U13371 (N_13371,N_12073,N_12414);
nand U13372 (N_13372,N_12457,N_12204);
or U13373 (N_13373,N_12821,N_12413);
xor U13374 (N_13374,N_12039,N_12471);
nand U13375 (N_13375,N_12358,N_12937);
and U13376 (N_13376,N_12292,N_12395);
nor U13377 (N_13377,N_12486,N_12223);
nor U13378 (N_13378,N_12587,N_12021);
or U13379 (N_13379,N_12828,N_12049);
or U13380 (N_13380,N_12997,N_12224);
xor U13381 (N_13381,N_12938,N_12914);
and U13382 (N_13382,N_12265,N_12122);
and U13383 (N_13383,N_12765,N_12286);
nor U13384 (N_13384,N_12231,N_12818);
xor U13385 (N_13385,N_12749,N_12334);
nor U13386 (N_13386,N_12470,N_12967);
nor U13387 (N_13387,N_12536,N_12428);
xnor U13388 (N_13388,N_12458,N_12452);
nand U13389 (N_13389,N_12655,N_12970);
or U13390 (N_13390,N_12293,N_12762);
nand U13391 (N_13391,N_12412,N_12032);
nor U13392 (N_13392,N_12824,N_12578);
xnor U13393 (N_13393,N_12009,N_12317);
or U13394 (N_13394,N_12975,N_12677);
nand U13395 (N_13395,N_12001,N_12356);
nand U13396 (N_13396,N_12476,N_12512);
or U13397 (N_13397,N_12156,N_12274);
and U13398 (N_13398,N_12691,N_12349);
nand U13399 (N_13399,N_12295,N_12751);
nand U13400 (N_13400,N_12081,N_12660);
nor U13401 (N_13401,N_12720,N_12764);
nand U13402 (N_13402,N_12451,N_12944);
xnor U13403 (N_13403,N_12322,N_12763);
and U13404 (N_13404,N_12351,N_12883);
and U13405 (N_13405,N_12145,N_12788);
or U13406 (N_13406,N_12337,N_12394);
or U13407 (N_13407,N_12435,N_12287);
or U13408 (N_13408,N_12346,N_12835);
xnor U13409 (N_13409,N_12409,N_12614);
and U13410 (N_13410,N_12533,N_12861);
or U13411 (N_13411,N_12147,N_12980);
xnor U13412 (N_13412,N_12016,N_12565);
xnor U13413 (N_13413,N_12868,N_12427);
or U13414 (N_13414,N_12155,N_12845);
nand U13415 (N_13415,N_12939,N_12843);
nor U13416 (N_13416,N_12085,N_12472);
nor U13417 (N_13417,N_12916,N_12635);
and U13418 (N_13418,N_12279,N_12577);
and U13419 (N_13419,N_12138,N_12760);
xnor U13420 (N_13420,N_12672,N_12280);
or U13421 (N_13421,N_12386,N_12192);
or U13422 (N_13422,N_12802,N_12490);
xor U13423 (N_13423,N_12986,N_12150);
and U13424 (N_13424,N_12357,N_12839);
or U13425 (N_13425,N_12976,N_12892);
or U13426 (N_13426,N_12383,N_12243);
nor U13427 (N_13427,N_12811,N_12088);
nor U13428 (N_13428,N_12269,N_12126);
and U13429 (N_13429,N_12263,N_12641);
nor U13430 (N_13430,N_12134,N_12054);
nand U13431 (N_13431,N_12043,N_12425);
and U13432 (N_13432,N_12111,N_12946);
nand U13433 (N_13433,N_12060,N_12866);
nand U13434 (N_13434,N_12405,N_12028);
nand U13435 (N_13435,N_12379,N_12650);
and U13436 (N_13436,N_12200,N_12590);
or U13437 (N_13437,N_12877,N_12875);
xor U13438 (N_13438,N_12329,N_12289);
and U13439 (N_13439,N_12652,N_12700);
or U13440 (N_13440,N_12535,N_12612);
nand U13441 (N_13441,N_12988,N_12008);
nand U13442 (N_13442,N_12115,N_12550);
nand U13443 (N_13443,N_12785,N_12943);
and U13444 (N_13444,N_12300,N_12708);
nand U13445 (N_13445,N_12162,N_12236);
and U13446 (N_13446,N_12364,N_12758);
nand U13447 (N_13447,N_12277,N_12838);
nand U13448 (N_13448,N_12097,N_12683);
and U13449 (N_13449,N_12701,N_12441);
or U13450 (N_13450,N_12220,N_12450);
nand U13451 (N_13451,N_12930,N_12504);
nor U13452 (N_13452,N_12516,N_12990);
or U13453 (N_13453,N_12136,N_12320);
nor U13454 (N_13454,N_12804,N_12123);
and U13455 (N_13455,N_12964,N_12084);
xor U13456 (N_13456,N_12687,N_12362);
or U13457 (N_13457,N_12853,N_12582);
nand U13458 (N_13458,N_12406,N_12055);
nor U13459 (N_13459,N_12809,N_12903);
and U13460 (N_13460,N_12218,N_12326);
nand U13461 (N_13461,N_12674,N_12745);
nor U13462 (N_13462,N_12331,N_12048);
nor U13463 (N_13463,N_12784,N_12475);
nand U13464 (N_13464,N_12034,N_12057);
xor U13465 (N_13465,N_12933,N_12985);
nand U13466 (N_13466,N_12325,N_12894);
and U13467 (N_13467,N_12102,N_12033);
nor U13468 (N_13468,N_12680,N_12132);
nor U13469 (N_13469,N_12505,N_12402);
or U13470 (N_13470,N_12778,N_12659);
nand U13471 (N_13471,N_12378,N_12267);
or U13472 (N_13472,N_12713,N_12834);
nand U13473 (N_13473,N_12501,N_12646);
and U13474 (N_13474,N_12133,N_12616);
xor U13475 (N_13475,N_12179,N_12518);
nor U13476 (N_13476,N_12366,N_12899);
nand U13477 (N_13477,N_12229,N_12481);
nor U13478 (N_13478,N_12306,N_12093);
and U13479 (N_13479,N_12373,N_12240);
nor U13480 (N_13480,N_12444,N_12959);
and U13481 (N_13481,N_12968,N_12643);
or U13482 (N_13482,N_12540,N_12447);
nor U13483 (N_13483,N_12510,N_12919);
nand U13484 (N_13484,N_12347,N_12915);
and U13485 (N_13485,N_12498,N_12002);
nor U13486 (N_13486,N_12653,N_12275);
or U13487 (N_13487,N_12129,N_12185);
and U13488 (N_13488,N_12493,N_12430);
nor U13489 (N_13489,N_12800,N_12310);
nor U13490 (N_13490,N_12769,N_12517);
nand U13491 (N_13491,N_12595,N_12003);
and U13492 (N_13492,N_12080,N_12382);
or U13493 (N_13493,N_12215,N_12794);
or U13494 (N_13494,N_12167,N_12611);
or U13495 (N_13495,N_12597,N_12886);
or U13496 (N_13496,N_12733,N_12146);
or U13497 (N_13497,N_12089,N_12558);
and U13498 (N_13498,N_12082,N_12770);
nor U13499 (N_13499,N_12355,N_12159);
nor U13500 (N_13500,N_12940,N_12945);
and U13501 (N_13501,N_12145,N_12408);
or U13502 (N_13502,N_12484,N_12293);
nor U13503 (N_13503,N_12852,N_12853);
or U13504 (N_13504,N_12504,N_12365);
and U13505 (N_13505,N_12566,N_12062);
xor U13506 (N_13506,N_12767,N_12872);
nand U13507 (N_13507,N_12309,N_12531);
nand U13508 (N_13508,N_12161,N_12349);
xor U13509 (N_13509,N_12145,N_12473);
and U13510 (N_13510,N_12786,N_12125);
nand U13511 (N_13511,N_12002,N_12542);
nand U13512 (N_13512,N_12810,N_12977);
nand U13513 (N_13513,N_12134,N_12567);
nand U13514 (N_13514,N_12528,N_12902);
or U13515 (N_13515,N_12507,N_12735);
nor U13516 (N_13516,N_12800,N_12491);
or U13517 (N_13517,N_12068,N_12827);
nor U13518 (N_13518,N_12562,N_12065);
or U13519 (N_13519,N_12630,N_12827);
xnor U13520 (N_13520,N_12951,N_12084);
nand U13521 (N_13521,N_12937,N_12605);
or U13522 (N_13522,N_12819,N_12912);
and U13523 (N_13523,N_12279,N_12587);
or U13524 (N_13524,N_12036,N_12777);
nand U13525 (N_13525,N_12383,N_12100);
nand U13526 (N_13526,N_12744,N_12638);
xnor U13527 (N_13527,N_12381,N_12778);
and U13528 (N_13528,N_12439,N_12187);
xor U13529 (N_13529,N_12330,N_12926);
nand U13530 (N_13530,N_12061,N_12370);
and U13531 (N_13531,N_12654,N_12261);
nor U13532 (N_13532,N_12479,N_12107);
xnor U13533 (N_13533,N_12572,N_12926);
nor U13534 (N_13534,N_12131,N_12315);
or U13535 (N_13535,N_12530,N_12894);
nand U13536 (N_13536,N_12958,N_12596);
nand U13537 (N_13537,N_12324,N_12456);
nor U13538 (N_13538,N_12571,N_12703);
and U13539 (N_13539,N_12489,N_12268);
nand U13540 (N_13540,N_12318,N_12425);
xor U13541 (N_13541,N_12883,N_12424);
or U13542 (N_13542,N_12897,N_12488);
nand U13543 (N_13543,N_12738,N_12424);
or U13544 (N_13544,N_12209,N_12318);
or U13545 (N_13545,N_12971,N_12824);
nand U13546 (N_13546,N_12153,N_12738);
nand U13547 (N_13547,N_12307,N_12509);
nor U13548 (N_13548,N_12660,N_12553);
nor U13549 (N_13549,N_12001,N_12581);
xor U13550 (N_13550,N_12373,N_12526);
and U13551 (N_13551,N_12103,N_12730);
or U13552 (N_13552,N_12611,N_12776);
xor U13553 (N_13553,N_12184,N_12020);
nand U13554 (N_13554,N_12383,N_12440);
nor U13555 (N_13555,N_12809,N_12612);
or U13556 (N_13556,N_12569,N_12929);
nand U13557 (N_13557,N_12282,N_12173);
nor U13558 (N_13558,N_12621,N_12633);
xor U13559 (N_13559,N_12449,N_12981);
nor U13560 (N_13560,N_12978,N_12081);
xnor U13561 (N_13561,N_12046,N_12468);
nor U13562 (N_13562,N_12369,N_12646);
or U13563 (N_13563,N_12408,N_12588);
and U13564 (N_13564,N_12461,N_12026);
nor U13565 (N_13565,N_12803,N_12774);
nor U13566 (N_13566,N_12229,N_12068);
nor U13567 (N_13567,N_12728,N_12627);
xnor U13568 (N_13568,N_12727,N_12525);
nand U13569 (N_13569,N_12954,N_12270);
nor U13570 (N_13570,N_12179,N_12188);
nand U13571 (N_13571,N_12859,N_12605);
nand U13572 (N_13572,N_12698,N_12269);
xor U13573 (N_13573,N_12361,N_12267);
nand U13574 (N_13574,N_12894,N_12058);
or U13575 (N_13575,N_12843,N_12600);
nor U13576 (N_13576,N_12379,N_12178);
or U13577 (N_13577,N_12476,N_12430);
xnor U13578 (N_13578,N_12779,N_12077);
or U13579 (N_13579,N_12285,N_12248);
nor U13580 (N_13580,N_12536,N_12026);
and U13581 (N_13581,N_12487,N_12896);
and U13582 (N_13582,N_12528,N_12931);
or U13583 (N_13583,N_12455,N_12778);
nand U13584 (N_13584,N_12360,N_12266);
nor U13585 (N_13585,N_12364,N_12883);
and U13586 (N_13586,N_12794,N_12242);
nand U13587 (N_13587,N_12666,N_12811);
and U13588 (N_13588,N_12651,N_12635);
and U13589 (N_13589,N_12794,N_12921);
xor U13590 (N_13590,N_12090,N_12851);
or U13591 (N_13591,N_12441,N_12410);
or U13592 (N_13592,N_12833,N_12604);
nor U13593 (N_13593,N_12682,N_12829);
nand U13594 (N_13594,N_12056,N_12599);
and U13595 (N_13595,N_12401,N_12092);
or U13596 (N_13596,N_12294,N_12055);
and U13597 (N_13597,N_12131,N_12486);
xnor U13598 (N_13598,N_12517,N_12284);
nand U13599 (N_13599,N_12579,N_12552);
nand U13600 (N_13600,N_12713,N_12734);
nand U13601 (N_13601,N_12408,N_12433);
nand U13602 (N_13602,N_12729,N_12927);
nand U13603 (N_13603,N_12540,N_12983);
xnor U13604 (N_13604,N_12787,N_12961);
nand U13605 (N_13605,N_12287,N_12994);
nand U13606 (N_13606,N_12595,N_12441);
and U13607 (N_13607,N_12646,N_12290);
and U13608 (N_13608,N_12689,N_12983);
nor U13609 (N_13609,N_12188,N_12814);
nand U13610 (N_13610,N_12515,N_12829);
and U13611 (N_13611,N_12211,N_12395);
or U13612 (N_13612,N_12780,N_12656);
nor U13613 (N_13613,N_12436,N_12586);
nand U13614 (N_13614,N_12266,N_12483);
nand U13615 (N_13615,N_12127,N_12458);
nor U13616 (N_13616,N_12675,N_12339);
nand U13617 (N_13617,N_12016,N_12156);
nor U13618 (N_13618,N_12040,N_12627);
xnor U13619 (N_13619,N_12827,N_12889);
or U13620 (N_13620,N_12384,N_12193);
nor U13621 (N_13621,N_12380,N_12106);
and U13622 (N_13622,N_12530,N_12080);
nand U13623 (N_13623,N_12167,N_12594);
and U13624 (N_13624,N_12413,N_12253);
nor U13625 (N_13625,N_12275,N_12671);
and U13626 (N_13626,N_12751,N_12475);
and U13627 (N_13627,N_12258,N_12699);
nand U13628 (N_13628,N_12150,N_12867);
nor U13629 (N_13629,N_12287,N_12175);
and U13630 (N_13630,N_12645,N_12870);
nand U13631 (N_13631,N_12739,N_12672);
or U13632 (N_13632,N_12218,N_12706);
or U13633 (N_13633,N_12915,N_12527);
and U13634 (N_13634,N_12958,N_12443);
nor U13635 (N_13635,N_12565,N_12075);
and U13636 (N_13636,N_12236,N_12649);
xnor U13637 (N_13637,N_12436,N_12091);
and U13638 (N_13638,N_12895,N_12652);
or U13639 (N_13639,N_12324,N_12058);
and U13640 (N_13640,N_12861,N_12918);
nand U13641 (N_13641,N_12131,N_12830);
nor U13642 (N_13642,N_12288,N_12890);
nor U13643 (N_13643,N_12468,N_12936);
nand U13644 (N_13644,N_12944,N_12466);
xor U13645 (N_13645,N_12729,N_12080);
xnor U13646 (N_13646,N_12246,N_12425);
nor U13647 (N_13647,N_12567,N_12447);
nand U13648 (N_13648,N_12561,N_12922);
and U13649 (N_13649,N_12641,N_12260);
nor U13650 (N_13650,N_12158,N_12643);
and U13651 (N_13651,N_12668,N_12579);
nor U13652 (N_13652,N_12185,N_12499);
nand U13653 (N_13653,N_12557,N_12482);
and U13654 (N_13654,N_12467,N_12061);
and U13655 (N_13655,N_12801,N_12836);
xor U13656 (N_13656,N_12746,N_12321);
or U13657 (N_13657,N_12804,N_12909);
nand U13658 (N_13658,N_12013,N_12881);
or U13659 (N_13659,N_12084,N_12370);
or U13660 (N_13660,N_12089,N_12840);
nand U13661 (N_13661,N_12638,N_12277);
nand U13662 (N_13662,N_12388,N_12249);
or U13663 (N_13663,N_12701,N_12455);
or U13664 (N_13664,N_12184,N_12941);
and U13665 (N_13665,N_12144,N_12494);
and U13666 (N_13666,N_12918,N_12113);
or U13667 (N_13667,N_12987,N_12656);
and U13668 (N_13668,N_12316,N_12463);
nand U13669 (N_13669,N_12231,N_12023);
xnor U13670 (N_13670,N_12388,N_12857);
nor U13671 (N_13671,N_12581,N_12732);
or U13672 (N_13672,N_12220,N_12049);
or U13673 (N_13673,N_12583,N_12283);
or U13674 (N_13674,N_12747,N_12974);
nand U13675 (N_13675,N_12442,N_12577);
and U13676 (N_13676,N_12514,N_12539);
nor U13677 (N_13677,N_12118,N_12422);
and U13678 (N_13678,N_12160,N_12882);
xnor U13679 (N_13679,N_12757,N_12239);
nand U13680 (N_13680,N_12408,N_12015);
xnor U13681 (N_13681,N_12994,N_12793);
nor U13682 (N_13682,N_12674,N_12646);
or U13683 (N_13683,N_12763,N_12369);
xor U13684 (N_13684,N_12305,N_12442);
and U13685 (N_13685,N_12422,N_12890);
and U13686 (N_13686,N_12117,N_12461);
nor U13687 (N_13687,N_12048,N_12286);
nor U13688 (N_13688,N_12583,N_12750);
nand U13689 (N_13689,N_12214,N_12763);
nor U13690 (N_13690,N_12818,N_12900);
or U13691 (N_13691,N_12066,N_12314);
nand U13692 (N_13692,N_12073,N_12772);
or U13693 (N_13693,N_12470,N_12040);
nand U13694 (N_13694,N_12392,N_12195);
nor U13695 (N_13695,N_12474,N_12970);
xor U13696 (N_13696,N_12674,N_12129);
xnor U13697 (N_13697,N_12519,N_12267);
or U13698 (N_13698,N_12371,N_12835);
nand U13699 (N_13699,N_12521,N_12478);
nor U13700 (N_13700,N_12357,N_12068);
nor U13701 (N_13701,N_12200,N_12122);
nand U13702 (N_13702,N_12289,N_12125);
and U13703 (N_13703,N_12192,N_12199);
xor U13704 (N_13704,N_12873,N_12427);
nor U13705 (N_13705,N_12674,N_12657);
nand U13706 (N_13706,N_12787,N_12080);
and U13707 (N_13707,N_12105,N_12249);
and U13708 (N_13708,N_12811,N_12968);
nand U13709 (N_13709,N_12966,N_12112);
or U13710 (N_13710,N_12056,N_12962);
xnor U13711 (N_13711,N_12129,N_12508);
nor U13712 (N_13712,N_12460,N_12418);
nor U13713 (N_13713,N_12836,N_12701);
nand U13714 (N_13714,N_12959,N_12674);
xor U13715 (N_13715,N_12043,N_12018);
nor U13716 (N_13716,N_12705,N_12355);
xor U13717 (N_13717,N_12171,N_12045);
and U13718 (N_13718,N_12354,N_12749);
xor U13719 (N_13719,N_12094,N_12521);
nand U13720 (N_13720,N_12278,N_12482);
nor U13721 (N_13721,N_12565,N_12930);
and U13722 (N_13722,N_12591,N_12811);
nor U13723 (N_13723,N_12128,N_12422);
nor U13724 (N_13724,N_12786,N_12508);
or U13725 (N_13725,N_12106,N_12890);
or U13726 (N_13726,N_12408,N_12017);
xor U13727 (N_13727,N_12322,N_12465);
xor U13728 (N_13728,N_12399,N_12515);
and U13729 (N_13729,N_12480,N_12411);
nor U13730 (N_13730,N_12332,N_12866);
nand U13731 (N_13731,N_12450,N_12615);
or U13732 (N_13732,N_12972,N_12839);
nor U13733 (N_13733,N_12369,N_12094);
nor U13734 (N_13734,N_12909,N_12277);
or U13735 (N_13735,N_12551,N_12170);
and U13736 (N_13736,N_12398,N_12651);
nand U13737 (N_13737,N_12288,N_12934);
nand U13738 (N_13738,N_12234,N_12969);
xor U13739 (N_13739,N_12090,N_12367);
nor U13740 (N_13740,N_12635,N_12634);
nor U13741 (N_13741,N_12541,N_12417);
nor U13742 (N_13742,N_12570,N_12467);
nor U13743 (N_13743,N_12053,N_12614);
and U13744 (N_13744,N_12862,N_12843);
nand U13745 (N_13745,N_12003,N_12714);
nand U13746 (N_13746,N_12171,N_12911);
nand U13747 (N_13747,N_12528,N_12690);
xor U13748 (N_13748,N_12200,N_12378);
or U13749 (N_13749,N_12885,N_12398);
or U13750 (N_13750,N_12010,N_12805);
or U13751 (N_13751,N_12477,N_12681);
nand U13752 (N_13752,N_12182,N_12423);
nor U13753 (N_13753,N_12466,N_12213);
and U13754 (N_13754,N_12240,N_12148);
nor U13755 (N_13755,N_12718,N_12247);
nand U13756 (N_13756,N_12912,N_12301);
xnor U13757 (N_13757,N_12108,N_12414);
xor U13758 (N_13758,N_12976,N_12246);
nor U13759 (N_13759,N_12718,N_12269);
nor U13760 (N_13760,N_12836,N_12363);
nand U13761 (N_13761,N_12643,N_12188);
nand U13762 (N_13762,N_12213,N_12557);
nand U13763 (N_13763,N_12083,N_12524);
xnor U13764 (N_13764,N_12952,N_12738);
nand U13765 (N_13765,N_12577,N_12112);
nor U13766 (N_13766,N_12467,N_12044);
nor U13767 (N_13767,N_12803,N_12718);
nor U13768 (N_13768,N_12178,N_12103);
and U13769 (N_13769,N_12169,N_12291);
and U13770 (N_13770,N_12043,N_12437);
and U13771 (N_13771,N_12837,N_12456);
nand U13772 (N_13772,N_12873,N_12397);
nor U13773 (N_13773,N_12000,N_12064);
nor U13774 (N_13774,N_12517,N_12873);
nor U13775 (N_13775,N_12011,N_12186);
xor U13776 (N_13776,N_12282,N_12647);
nand U13777 (N_13777,N_12457,N_12576);
xnor U13778 (N_13778,N_12782,N_12551);
nand U13779 (N_13779,N_12950,N_12660);
nor U13780 (N_13780,N_12230,N_12773);
and U13781 (N_13781,N_12177,N_12338);
nand U13782 (N_13782,N_12661,N_12415);
and U13783 (N_13783,N_12102,N_12661);
xnor U13784 (N_13784,N_12375,N_12054);
nand U13785 (N_13785,N_12964,N_12074);
nor U13786 (N_13786,N_12183,N_12531);
or U13787 (N_13787,N_12715,N_12779);
nand U13788 (N_13788,N_12503,N_12181);
nand U13789 (N_13789,N_12917,N_12208);
or U13790 (N_13790,N_12039,N_12837);
or U13791 (N_13791,N_12214,N_12679);
and U13792 (N_13792,N_12923,N_12173);
or U13793 (N_13793,N_12131,N_12529);
nor U13794 (N_13794,N_12686,N_12150);
or U13795 (N_13795,N_12243,N_12109);
or U13796 (N_13796,N_12047,N_12789);
or U13797 (N_13797,N_12634,N_12981);
and U13798 (N_13798,N_12420,N_12492);
and U13799 (N_13799,N_12942,N_12566);
and U13800 (N_13800,N_12733,N_12565);
nand U13801 (N_13801,N_12553,N_12954);
nand U13802 (N_13802,N_12036,N_12160);
or U13803 (N_13803,N_12816,N_12367);
nand U13804 (N_13804,N_12511,N_12480);
nand U13805 (N_13805,N_12141,N_12589);
and U13806 (N_13806,N_12184,N_12073);
and U13807 (N_13807,N_12855,N_12305);
nand U13808 (N_13808,N_12104,N_12515);
xnor U13809 (N_13809,N_12578,N_12996);
and U13810 (N_13810,N_12873,N_12931);
or U13811 (N_13811,N_12878,N_12451);
and U13812 (N_13812,N_12920,N_12433);
nor U13813 (N_13813,N_12860,N_12223);
nand U13814 (N_13814,N_12794,N_12930);
or U13815 (N_13815,N_12134,N_12241);
nor U13816 (N_13816,N_12459,N_12193);
xnor U13817 (N_13817,N_12637,N_12216);
xnor U13818 (N_13818,N_12804,N_12697);
or U13819 (N_13819,N_12364,N_12966);
or U13820 (N_13820,N_12084,N_12065);
nor U13821 (N_13821,N_12040,N_12629);
or U13822 (N_13822,N_12996,N_12282);
and U13823 (N_13823,N_12612,N_12058);
and U13824 (N_13824,N_12334,N_12498);
or U13825 (N_13825,N_12024,N_12241);
and U13826 (N_13826,N_12737,N_12048);
xor U13827 (N_13827,N_12258,N_12036);
nor U13828 (N_13828,N_12408,N_12661);
nand U13829 (N_13829,N_12813,N_12507);
nor U13830 (N_13830,N_12688,N_12484);
nand U13831 (N_13831,N_12075,N_12086);
nand U13832 (N_13832,N_12657,N_12334);
nor U13833 (N_13833,N_12280,N_12041);
or U13834 (N_13834,N_12248,N_12550);
or U13835 (N_13835,N_12092,N_12770);
or U13836 (N_13836,N_12864,N_12694);
and U13837 (N_13837,N_12914,N_12297);
and U13838 (N_13838,N_12160,N_12173);
nand U13839 (N_13839,N_12848,N_12847);
or U13840 (N_13840,N_12284,N_12348);
or U13841 (N_13841,N_12277,N_12779);
nor U13842 (N_13842,N_12835,N_12121);
nand U13843 (N_13843,N_12349,N_12148);
nand U13844 (N_13844,N_12295,N_12707);
nor U13845 (N_13845,N_12448,N_12780);
nor U13846 (N_13846,N_12781,N_12873);
and U13847 (N_13847,N_12869,N_12611);
xor U13848 (N_13848,N_12052,N_12150);
or U13849 (N_13849,N_12236,N_12496);
nand U13850 (N_13850,N_12835,N_12857);
nor U13851 (N_13851,N_12597,N_12084);
nor U13852 (N_13852,N_12624,N_12417);
or U13853 (N_13853,N_12518,N_12326);
or U13854 (N_13854,N_12928,N_12893);
nand U13855 (N_13855,N_12082,N_12501);
nor U13856 (N_13856,N_12610,N_12848);
xor U13857 (N_13857,N_12552,N_12391);
nand U13858 (N_13858,N_12802,N_12748);
or U13859 (N_13859,N_12817,N_12151);
or U13860 (N_13860,N_12194,N_12622);
and U13861 (N_13861,N_12205,N_12151);
or U13862 (N_13862,N_12375,N_12523);
nand U13863 (N_13863,N_12585,N_12369);
and U13864 (N_13864,N_12583,N_12692);
or U13865 (N_13865,N_12100,N_12632);
nand U13866 (N_13866,N_12443,N_12478);
xnor U13867 (N_13867,N_12965,N_12142);
nor U13868 (N_13868,N_12780,N_12733);
nand U13869 (N_13869,N_12194,N_12148);
nand U13870 (N_13870,N_12853,N_12061);
and U13871 (N_13871,N_12089,N_12145);
or U13872 (N_13872,N_12075,N_12522);
nor U13873 (N_13873,N_12832,N_12688);
or U13874 (N_13874,N_12924,N_12407);
and U13875 (N_13875,N_12401,N_12462);
or U13876 (N_13876,N_12548,N_12451);
and U13877 (N_13877,N_12414,N_12743);
nand U13878 (N_13878,N_12858,N_12871);
nor U13879 (N_13879,N_12340,N_12579);
or U13880 (N_13880,N_12777,N_12882);
nor U13881 (N_13881,N_12448,N_12476);
nand U13882 (N_13882,N_12878,N_12350);
nand U13883 (N_13883,N_12893,N_12021);
nand U13884 (N_13884,N_12753,N_12174);
and U13885 (N_13885,N_12237,N_12172);
nor U13886 (N_13886,N_12230,N_12765);
nand U13887 (N_13887,N_12407,N_12697);
or U13888 (N_13888,N_12834,N_12040);
nor U13889 (N_13889,N_12207,N_12624);
nand U13890 (N_13890,N_12165,N_12313);
xor U13891 (N_13891,N_12996,N_12719);
nand U13892 (N_13892,N_12567,N_12497);
and U13893 (N_13893,N_12056,N_12716);
nand U13894 (N_13894,N_12796,N_12613);
or U13895 (N_13895,N_12985,N_12972);
or U13896 (N_13896,N_12625,N_12275);
or U13897 (N_13897,N_12832,N_12837);
nor U13898 (N_13898,N_12799,N_12906);
nand U13899 (N_13899,N_12184,N_12095);
and U13900 (N_13900,N_12630,N_12446);
nor U13901 (N_13901,N_12002,N_12016);
or U13902 (N_13902,N_12559,N_12720);
nor U13903 (N_13903,N_12394,N_12673);
xnor U13904 (N_13904,N_12657,N_12862);
nand U13905 (N_13905,N_12253,N_12473);
nand U13906 (N_13906,N_12503,N_12683);
or U13907 (N_13907,N_12961,N_12716);
nor U13908 (N_13908,N_12227,N_12072);
nand U13909 (N_13909,N_12621,N_12701);
or U13910 (N_13910,N_12959,N_12201);
nand U13911 (N_13911,N_12313,N_12955);
or U13912 (N_13912,N_12314,N_12640);
or U13913 (N_13913,N_12947,N_12432);
nor U13914 (N_13914,N_12609,N_12213);
xor U13915 (N_13915,N_12516,N_12822);
and U13916 (N_13916,N_12270,N_12441);
or U13917 (N_13917,N_12971,N_12098);
or U13918 (N_13918,N_12907,N_12700);
nand U13919 (N_13919,N_12337,N_12939);
or U13920 (N_13920,N_12449,N_12620);
or U13921 (N_13921,N_12540,N_12952);
or U13922 (N_13922,N_12319,N_12991);
or U13923 (N_13923,N_12779,N_12088);
xnor U13924 (N_13924,N_12278,N_12024);
nand U13925 (N_13925,N_12170,N_12436);
xnor U13926 (N_13926,N_12484,N_12333);
and U13927 (N_13927,N_12288,N_12034);
and U13928 (N_13928,N_12516,N_12345);
xnor U13929 (N_13929,N_12099,N_12143);
xor U13930 (N_13930,N_12913,N_12851);
and U13931 (N_13931,N_12117,N_12850);
or U13932 (N_13932,N_12571,N_12959);
and U13933 (N_13933,N_12120,N_12743);
nand U13934 (N_13934,N_12464,N_12439);
and U13935 (N_13935,N_12987,N_12031);
xnor U13936 (N_13936,N_12332,N_12480);
nor U13937 (N_13937,N_12636,N_12066);
nand U13938 (N_13938,N_12730,N_12479);
nor U13939 (N_13939,N_12088,N_12025);
or U13940 (N_13940,N_12691,N_12794);
or U13941 (N_13941,N_12836,N_12966);
and U13942 (N_13942,N_12821,N_12546);
and U13943 (N_13943,N_12854,N_12980);
nor U13944 (N_13944,N_12907,N_12224);
or U13945 (N_13945,N_12139,N_12076);
xnor U13946 (N_13946,N_12108,N_12390);
nor U13947 (N_13947,N_12483,N_12548);
nand U13948 (N_13948,N_12323,N_12231);
or U13949 (N_13949,N_12462,N_12310);
xor U13950 (N_13950,N_12674,N_12162);
xor U13951 (N_13951,N_12021,N_12920);
nand U13952 (N_13952,N_12062,N_12491);
and U13953 (N_13953,N_12184,N_12092);
nor U13954 (N_13954,N_12481,N_12887);
or U13955 (N_13955,N_12055,N_12247);
and U13956 (N_13956,N_12565,N_12478);
nand U13957 (N_13957,N_12029,N_12758);
or U13958 (N_13958,N_12520,N_12856);
nor U13959 (N_13959,N_12561,N_12078);
nor U13960 (N_13960,N_12582,N_12694);
or U13961 (N_13961,N_12742,N_12600);
or U13962 (N_13962,N_12536,N_12665);
nor U13963 (N_13963,N_12655,N_12562);
nor U13964 (N_13964,N_12799,N_12544);
xnor U13965 (N_13965,N_12003,N_12720);
nor U13966 (N_13966,N_12096,N_12119);
nor U13967 (N_13967,N_12443,N_12495);
and U13968 (N_13968,N_12361,N_12405);
xor U13969 (N_13969,N_12472,N_12415);
or U13970 (N_13970,N_12189,N_12724);
xor U13971 (N_13971,N_12896,N_12095);
nand U13972 (N_13972,N_12527,N_12697);
nor U13973 (N_13973,N_12873,N_12529);
and U13974 (N_13974,N_12323,N_12102);
nor U13975 (N_13975,N_12465,N_12983);
nand U13976 (N_13976,N_12719,N_12689);
nor U13977 (N_13977,N_12130,N_12580);
xnor U13978 (N_13978,N_12514,N_12477);
nor U13979 (N_13979,N_12098,N_12743);
and U13980 (N_13980,N_12081,N_12203);
and U13981 (N_13981,N_12797,N_12517);
and U13982 (N_13982,N_12381,N_12907);
or U13983 (N_13983,N_12047,N_12126);
xor U13984 (N_13984,N_12371,N_12433);
xor U13985 (N_13985,N_12740,N_12736);
nor U13986 (N_13986,N_12043,N_12190);
nor U13987 (N_13987,N_12663,N_12209);
and U13988 (N_13988,N_12449,N_12939);
xor U13989 (N_13989,N_12409,N_12953);
and U13990 (N_13990,N_12529,N_12142);
nor U13991 (N_13991,N_12901,N_12127);
and U13992 (N_13992,N_12752,N_12520);
nand U13993 (N_13993,N_12481,N_12336);
and U13994 (N_13994,N_12975,N_12946);
nand U13995 (N_13995,N_12862,N_12648);
xnor U13996 (N_13996,N_12791,N_12087);
nand U13997 (N_13997,N_12807,N_12584);
and U13998 (N_13998,N_12325,N_12965);
or U13999 (N_13999,N_12610,N_12853);
nor U14000 (N_14000,N_13724,N_13624);
xnor U14001 (N_14001,N_13030,N_13980);
nor U14002 (N_14002,N_13756,N_13375);
or U14003 (N_14003,N_13012,N_13549);
nor U14004 (N_14004,N_13665,N_13363);
nand U14005 (N_14005,N_13746,N_13581);
xnor U14006 (N_14006,N_13370,N_13646);
xnor U14007 (N_14007,N_13951,N_13804);
nand U14008 (N_14008,N_13047,N_13409);
or U14009 (N_14009,N_13236,N_13537);
nand U14010 (N_14010,N_13222,N_13832);
nor U14011 (N_14011,N_13253,N_13502);
or U14012 (N_14012,N_13563,N_13616);
nand U14013 (N_14013,N_13512,N_13632);
or U14014 (N_14014,N_13949,N_13550);
nor U14015 (N_14015,N_13493,N_13490);
nand U14016 (N_14016,N_13190,N_13544);
xnor U14017 (N_14017,N_13655,N_13643);
or U14018 (N_14018,N_13462,N_13240);
nor U14019 (N_14019,N_13191,N_13780);
and U14020 (N_14020,N_13471,N_13040);
or U14021 (N_14021,N_13694,N_13141);
nor U14022 (N_14022,N_13171,N_13451);
or U14023 (N_14023,N_13510,N_13132);
nand U14024 (N_14024,N_13459,N_13991);
or U14025 (N_14025,N_13196,N_13662);
and U14026 (N_14026,N_13175,N_13960);
or U14027 (N_14027,N_13970,N_13206);
or U14028 (N_14028,N_13693,N_13754);
and U14029 (N_14029,N_13975,N_13997);
nor U14030 (N_14030,N_13433,N_13388);
nand U14031 (N_14031,N_13577,N_13984);
nand U14032 (N_14032,N_13144,N_13416);
or U14033 (N_14033,N_13091,N_13114);
xor U14034 (N_14034,N_13080,N_13189);
nand U14035 (N_14035,N_13653,N_13257);
nand U14036 (N_14036,N_13648,N_13509);
or U14037 (N_14037,N_13677,N_13159);
nand U14038 (N_14038,N_13521,N_13306);
nand U14039 (N_14039,N_13546,N_13172);
and U14040 (N_14040,N_13015,N_13339);
nand U14041 (N_14041,N_13365,N_13186);
nor U14042 (N_14042,N_13018,N_13052);
nor U14043 (N_14043,N_13942,N_13274);
or U14044 (N_14044,N_13783,N_13859);
nand U14045 (N_14045,N_13219,N_13249);
nor U14046 (N_14046,N_13481,N_13461);
nand U14047 (N_14047,N_13226,N_13237);
nor U14048 (N_14048,N_13188,N_13273);
xor U14049 (N_14049,N_13759,N_13953);
and U14050 (N_14050,N_13848,N_13491);
nand U14051 (N_14051,N_13928,N_13800);
nor U14052 (N_14052,N_13495,N_13183);
and U14053 (N_14053,N_13663,N_13088);
and U14054 (N_14054,N_13879,N_13619);
nand U14055 (N_14055,N_13011,N_13041);
or U14056 (N_14056,N_13305,N_13115);
and U14057 (N_14057,N_13883,N_13831);
and U14058 (N_14058,N_13538,N_13340);
nor U14059 (N_14059,N_13452,N_13393);
nand U14060 (N_14060,N_13634,N_13788);
and U14061 (N_14061,N_13841,N_13422);
nor U14062 (N_14062,N_13193,N_13642);
and U14063 (N_14063,N_13977,N_13966);
nor U14064 (N_14064,N_13534,N_13728);
or U14065 (N_14065,N_13936,N_13212);
and U14066 (N_14066,N_13364,N_13057);
nand U14067 (N_14067,N_13152,N_13398);
nor U14068 (N_14068,N_13153,N_13664);
nor U14069 (N_14069,N_13245,N_13808);
nor U14070 (N_14070,N_13711,N_13683);
or U14071 (N_14071,N_13582,N_13947);
or U14072 (N_14072,N_13164,N_13307);
or U14073 (N_14073,N_13629,N_13707);
nor U14074 (N_14074,N_13496,N_13044);
nand U14075 (N_14075,N_13527,N_13081);
and U14076 (N_14076,N_13691,N_13372);
xor U14077 (N_14077,N_13448,N_13368);
and U14078 (N_14078,N_13916,N_13034);
nand U14079 (N_14079,N_13813,N_13633);
nand U14080 (N_14080,N_13134,N_13874);
nand U14081 (N_14081,N_13014,N_13116);
xnor U14082 (N_14082,N_13126,N_13921);
nand U14083 (N_14083,N_13476,N_13926);
xor U14084 (N_14084,N_13466,N_13743);
and U14085 (N_14085,N_13732,N_13553);
and U14086 (N_14086,N_13096,N_13666);
nand U14087 (N_14087,N_13238,N_13342);
and U14088 (N_14088,N_13024,N_13397);
xor U14089 (N_14089,N_13199,N_13559);
or U14090 (N_14090,N_13726,N_13233);
nor U14091 (N_14091,N_13501,N_13678);
nor U14092 (N_14092,N_13705,N_13809);
and U14093 (N_14093,N_13596,N_13676);
and U14094 (N_14094,N_13149,N_13647);
and U14095 (N_14095,N_13661,N_13252);
nand U14096 (N_14096,N_13635,N_13455);
nand U14097 (N_14097,N_13837,N_13794);
nor U14098 (N_14098,N_13264,N_13009);
or U14099 (N_14099,N_13300,N_13346);
and U14100 (N_14100,N_13280,N_13505);
and U14101 (N_14101,N_13427,N_13042);
and U14102 (N_14102,N_13875,N_13934);
nor U14103 (N_14103,N_13922,N_13757);
and U14104 (N_14104,N_13344,N_13295);
nor U14105 (N_14105,N_13519,N_13299);
nor U14106 (N_14106,N_13860,N_13479);
nor U14107 (N_14107,N_13962,N_13389);
xnor U14108 (N_14108,N_13426,N_13310);
nor U14109 (N_14109,N_13939,N_13197);
nand U14110 (N_14110,N_13535,N_13680);
and U14111 (N_14111,N_13465,N_13271);
nor U14112 (N_14112,N_13444,N_13328);
nor U14113 (N_14113,N_13350,N_13688);
nand U14114 (N_14114,N_13355,N_13296);
and U14115 (N_14115,N_13434,N_13863);
and U14116 (N_14116,N_13637,N_13708);
or U14117 (N_14117,N_13309,N_13901);
and U14118 (N_14118,N_13784,N_13628);
or U14119 (N_14119,N_13781,N_13805);
or U14120 (N_14120,N_13806,N_13399);
and U14121 (N_14121,N_13109,N_13076);
xor U14122 (N_14122,N_13354,N_13558);
or U14123 (N_14123,N_13303,N_13500);
and U14124 (N_14124,N_13971,N_13716);
nor U14125 (N_14125,N_13774,N_13838);
and U14126 (N_14126,N_13564,N_13626);
nand U14127 (N_14127,N_13897,N_13998);
nor U14128 (N_14128,N_13820,N_13542);
nor U14129 (N_14129,N_13259,N_13819);
xor U14130 (N_14130,N_13325,N_13792);
nand U14131 (N_14131,N_13378,N_13656);
nand U14132 (N_14132,N_13557,N_13570);
or U14133 (N_14133,N_13105,N_13737);
and U14134 (N_14134,N_13367,N_13021);
nor U14135 (N_14135,N_13963,N_13529);
xnor U14136 (N_14136,N_13752,N_13767);
nand U14137 (N_14137,N_13652,N_13288);
xor U14138 (N_14138,N_13727,N_13994);
nand U14139 (N_14139,N_13078,N_13441);
nor U14140 (N_14140,N_13170,N_13488);
or U14141 (N_14141,N_13195,N_13506);
and U14142 (N_14142,N_13486,N_13585);
xnor U14143 (N_14143,N_13074,N_13405);
or U14144 (N_14144,N_13996,N_13508);
xor U14145 (N_14145,N_13337,N_13002);
or U14146 (N_14146,N_13571,N_13326);
nor U14147 (N_14147,N_13704,N_13321);
nand U14148 (N_14148,N_13540,N_13979);
or U14149 (N_14149,N_13825,N_13920);
or U14150 (N_14150,N_13083,N_13391);
and U14151 (N_14151,N_13120,N_13896);
and U14152 (N_14152,N_13541,N_13404);
nand U14153 (N_14153,N_13595,N_13227);
or U14154 (N_14154,N_13122,N_13379);
and U14155 (N_14155,N_13061,N_13513);
or U14156 (N_14156,N_13394,N_13343);
or U14157 (N_14157,N_13981,N_13467);
or U14158 (N_14158,N_13039,N_13889);
nand U14159 (N_14159,N_13686,N_13142);
and U14160 (N_14160,N_13167,N_13959);
nor U14161 (N_14161,N_13477,N_13782);
nand U14162 (N_14162,N_13871,N_13133);
xor U14163 (N_14163,N_13045,N_13004);
or U14164 (N_14164,N_13617,N_13881);
and U14165 (N_14165,N_13613,N_13673);
xnor U14166 (N_14166,N_13130,N_13762);
nand U14167 (N_14167,N_13766,N_13531);
or U14168 (N_14168,N_13318,N_13265);
nor U14169 (N_14169,N_13995,N_13161);
xnor U14170 (N_14170,N_13761,N_13507);
or U14171 (N_14171,N_13698,N_13866);
and U14172 (N_14172,N_13160,N_13103);
or U14173 (N_14173,N_13539,N_13763);
and U14174 (N_14174,N_13194,N_13868);
nand U14175 (N_14175,N_13100,N_13352);
nor U14176 (N_14176,N_13695,N_13670);
and U14177 (N_14177,N_13400,N_13740);
or U14178 (N_14178,N_13445,N_13154);
xor U14179 (N_14179,N_13843,N_13948);
and U14180 (N_14180,N_13200,N_13880);
or U14181 (N_14181,N_13447,N_13087);
nand U14182 (N_14182,N_13353,N_13438);
and U14183 (N_14183,N_13023,N_13861);
and U14184 (N_14184,N_13700,N_13483);
or U14185 (N_14185,N_13138,N_13381);
xor U14186 (N_14186,N_13803,N_13791);
nand U14187 (N_14187,N_13168,N_13623);
and U14188 (N_14188,N_13776,N_13954);
nand U14189 (N_14189,N_13988,N_13904);
nand U14190 (N_14190,N_13812,N_13575);
or U14191 (N_14191,N_13330,N_13218);
nor U14192 (N_14192,N_13873,N_13086);
or U14193 (N_14193,N_13258,N_13940);
and U14194 (N_14194,N_13056,N_13079);
nor U14195 (N_14195,N_13213,N_13048);
xor U14196 (N_14196,N_13514,N_13899);
nor U14197 (N_14197,N_13840,N_13703);
nor U14198 (N_14198,N_13877,N_13935);
and U14199 (N_14199,N_13450,N_13392);
xnor U14200 (N_14200,N_13058,N_13025);
or U14201 (N_14201,N_13232,N_13870);
and U14202 (N_14202,N_13589,N_13692);
nor U14203 (N_14203,N_13059,N_13900);
nand U14204 (N_14204,N_13890,N_13341);
or U14205 (N_14205,N_13473,N_13031);
nor U14206 (N_14206,N_13649,N_13972);
or U14207 (N_14207,N_13147,N_13923);
nor U14208 (N_14208,N_13854,N_13659);
nor U14209 (N_14209,N_13256,N_13129);
or U14210 (N_14210,N_13440,N_13464);
and U14211 (N_14211,N_13672,N_13121);
and U14212 (N_14212,N_13143,N_13658);
nor U14213 (N_14213,N_13718,N_13978);
nor U14214 (N_14214,N_13135,N_13796);
and U14215 (N_14215,N_13383,N_13119);
or U14216 (N_14216,N_13106,N_13064);
nor U14217 (N_14217,N_13001,N_13669);
nor U14218 (N_14218,N_13424,N_13811);
or U14219 (N_14219,N_13583,N_13586);
and U14220 (N_14220,N_13801,N_13362);
and U14221 (N_14221,N_13552,N_13822);
and U14222 (N_14222,N_13764,N_13660);
xor U14223 (N_14223,N_13329,N_13099);
and U14224 (N_14224,N_13667,N_13419);
nand U14225 (N_14225,N_13580,N_13855);
and U14226 (N_14226,N_13414,N_13373);
nand U14227 (N_14227,N_13876,N_13888);
nand U14228 (N_14228,N_13579,N_13145);
and U14229 (N_14229,N_13914,N_13443);
and U14230 (N_14230,N_13173,N_13773);
and U14231 (N_14231,N_13210,N_13554);
nor U14232 (N_14232,N_13903,N_13421);
and U14233 (N_14233,N_13208,N_13894);
and U14234 (N_14234,N_13182,N_13192);
or U14235 (N_14235,N_13163,N_13517);
xnor U14236 (N_14236,N_13753,N_13205);
xor U14237 (N_14237,N_13261,N_13906);
xor U14238 (N_14238,N_13687,N_13290);
xnor U14239 (N_14239,N_13730,N_13180);
xnor U14240 (N_14240,N_13815,N_13853);
and U14241 (N_14241,N_13036,N_13937);
or U14242 (N_14242,N_13260,N_13912);
nor U14243 (N_14243,N_13610,N_13231);
or U14244 (N_14244,N_13140,N_13911);
and U14245 (N_14245,N_13892,N_13316);
and U14246 (N_14246,N_13032,N_13003);
or U14247 (N_14247,N_13826,N_13184);
or U14248 (N_14248,N_13098,N_13107);
and U14249 (N_14249,N_13591,N_13857);
xor U14250 (N_14250,N_13242,N_13956);
nand U14251 (N_14251,N_13204,N_13244);
xnor U14252 (N_14252,N_13964,N_13640);
or U14253 (N_14253,N_13834,N_13987);
xor U14254 (N_14254,N_13967,N_13915);
and U14255 (N_14255,N_13384,N_13779);
or U14256 (N_14256,N_13177,N_13789);
or U14257 (N_14257,N_13602,N_13331);
nand U14258 (N_14258,N_13136,N_13387);
nor U14259 (N_14259,N_13046,N_13395);
and U14260 (N_14260,N_13515,N_13010);
nor U14261 (N_14261,N_13584,N_13844);
or U14262 (N_14262,N_13179,N_13124);
nor U14263 (N_14263,N_13351,N_13470);
nand U14264 (N_14264,N_13055,N_13930);
and U14265 (N_14265,N_13597,N_13101);
or U14266 (N_14266,N_13682,N_13230);
or U14267 (N_14267,N_13035,N_13576);
or U14268 (N_14268,N_13484,N_13733);
or U14269 (N_14269,N_13775,N_13603);
nor U14270 (N_14270,N_13385,N_13590);
or U14271 (N_14271,N_13952,N_13442);
nand U14272 (N_14272,N_13093,N_13068);
xnor U14273 (N_14273,N_13038,N_13458);
nand U14274 (N_14274,N_13498,N_13319);
and U14275 (N_14275,N_13282,N_13286);
nand U14276 (N_14276,N_13945,N_13714);
nand U14277 (N_14277,N_13713,N_13333);
or U14278 (N_14278,N_13958,N_13839);
nand U14279 (N_14279,N_13221,N_13262);
and U14280 (N_14280,N_13181,N_13250);
nand U14281 (N_14281,N_13469,N_13216);
nand U14282 (N_14282,N_13578,N_13263);
nand U14283 (N_14283,N_13220,N_13723);
or U14284 (N_14284,N_13816,N_13943);
or U14285 (N_14285,N_13178,N_13070);
or U14286 (N_14286,N_13000,N_13090);
and U14287 (N_14287,N_13835,N_13402);
and U14288 (N_14288,N_13908,N_13715);
xnor U14289 (N_14289,N_13437,N_13974);
and U14290 (N_14290,N_13066,N_13525);
or U14291 (N_14291,N_13986,N_13569);
nor U14292 (N_14292,N_13089,N_13008);
nand U14293 (N_14293,N_13411,N_13065);
xnor U14294 (N_14294,N_13335,N_13396);
and U14295 (N_14295,N_13403,N_13818);
nand U14296 (N_14296,N_13289,N_13872);
and U14297 (N_14297,N_13156,N_13551);
or U14298 (N_14298,N_13965,N_13255);
and U14299 (N_14299,N_13702,N_13611);
nand U14300 (N_14300,N_13618,N_13829);
and U14301 (N_14301,N_13174,N_13311);
nand U14302 (N_14302,N_13157,N_13671);
or U14303 (N_14303,N_13545,N_13478);
or U14304 (N_14304,N_13504,N_13037);
or U14305 (N_14305,N_13919,N_13574);
nand U14306 (N_14306,N_13865,N_13533);
and U14307 (N_14307,N_13146,N_13360);
nand U14308 (N_14308,N_13334,N_13439);
nand U14309 (N_14309,N_13281,N_13750);
nor U14310 (N_14310,N_13347,N_13650);
or U14311 (N_14311,N_13668,N_13689);
and U14312 (N_14312,N_13374,N_13925);
or U14313 (N_14313,N_13494,N_13909);
and U14314 (N_14314,N_13587,N_13814);
nand U14315 (N_14315,N_13968,N_13690);
nand U14316 (N_14316,N_13717,N_13770);
nand U14317 (N_14317,N_13830,N_13701);
xnor U14318 (N_14318,N_13913,N_13786);
nand U14319 (N_14319,N_13969,N_13797);
nor U14320 (N_14320,N_13085,N_13884);
nor U14321 (N_14321,N_13612,N_13847);
and U14322 (N_14322,N_13769,N_13741);
nand U14323 (N_14323,N_13802,N_13377);
nand U14324 (N_14324,N_13270,N_13312);
nand U14325 (N_14325,N_13893,N_13429);
or U14326 (N_14326,N_13069,N_13446);
or U14327 (N_14327,N_13294,N_13102);
nor U14328 (N_14328,N_13856,N_13125);
or U14329 (N_14329,N_13567,N_13721);
or U14330 (N_14330,N_13606,N_13412);
nor U14331 (N_14331,N_13833,N_13645);
or U14332 (N_14332,N_13449,N_13543);
nand U14333 (N_14333,N_13071,N_13565);
nor U14334 (N_14334,N_13845,N_13005);
xor U14335 (N_14335,N_13760,N_13675);
nor U14336 (N_14336,N_13739,N_13836);
nand U14337 (N_14337,N_13744,N_13927);
nor U14338 (N_14338,N_13123,N_13150);
nor U14339 (N_14339,N_13572,N_13104);
xor U14340 (N_14340,N_13878,N_13828);
and U14341 (N_14341,N_13735,N_13749);
or U14342 (N_14342,N_13654,N_13139);
nor U14343 (N_14343,N_13275,N_13778);
and U14344 (N_14344,N_13277,N_13850);
and U14345 (N_14345,N_13094,N_13198);
and U14346 (N_14346,N_13285,N_13607);
and U14347 (N_14347,N_13075,N_13625);
and U14348 (N_14348,N_13072,N_13622);
and U14349 (N_14349,N_13931,N_13428);
nor U14350 (N_14350,N_13291,N_13401);
nor U14351 (N_14351,N_13224,N_13082);
or U14352 (N_14352,N_13308,N_13530);
nand U14353 (N_14353,N_13166,N_13386);
nor U14354 (N_14354,N_13187,N_13598);
nor U14355 (N_14355,N_13961,N_13097);
nor U14356 (N_14356,N_13851,N_13348);
nor U14357 (N_14357,N_13938,N_13006);
and U14358 (N_14358,N_13063,N_13241);
xor U14359 (N_14359,N_13371,N_13176);
and U14360 (N_14360,N_13022,N_13933);
or U14361 (N_14361,N_13751,N_13929);
nand U14362 (N_14362,N_13799,N_13456);
nor U14363 (N_14363,N_13720,N_13638);
nand U14364 (N_14364,N_13485,N_13482);
nand U14365 (N_14365,N_13536,N_13468);
or U14366 (N_14366,N_13073,N_13910);
and U14367 (N_14367,N_13408,N_13887);
nand U14368 (N_14368,N_13999,N_13361);
or U14369 (N_14369,N_13731,N_13284);
or U14370 (N_14370,N_13382,N_13357);
or U14371 (N_14371,N_13017,N_13453);
nand U14372 (N_14372,N_13054,N_13725);
nor U14373 (N_14373,N_13019,N_13084);
and U14374 (N_14374,N_13787,N_13932);
and U14375 (N_14375,N_13941,N_13425);
or U14376 (N_14376,N_13983,N_13269);
and U14377 (N_14377,N_13415,N_13641);
nor U14378 (N_14378,N_13092,N_13033);
nor U14379 (N_14379,N_13918,N_13293);
nand U14380 (N_14380,N_13674,N_13165);
nand U14381 (N_14381,N_13267,N_13982);
or U14382 (N_14382,N_13706,N_13390);
nand U14383 (N_14383,N_13685,N_13007);
and U14384 (N_14384,N_13821,N_13679);
nand U14385 (N_14385,N_13867,N_13407);
and U14386 (N_14386,N_13547,N_13020);
or U14387 (N_14387,N_13601,N_13474);
or U14388 (N_14388,N_13118,N_13765);
nand U14389 (N_14389,N_13487,N_13946);
or U14390 (N_14390,N_13522,N_13560);
nor U14391 (N_14391,N_13338,N_13526);
nor U14392 (N_14392,N_13768,N_13302);
nand U14393 (N_14393,N_13413,N_13060);
or U14394 (N_14394,N_13279,N_13620);
nor U14395 (N_14395,N_13214,N_13566);
and U14396 (N_14396,N_13247,N_13957);
or U14397 (N_14397,N_13110,N_13593);
nor U14398 (N_14398,N_13272,N_13862);
or U14399 (N_14399,N_13235,N_13511);
nand U14400 (N_14400,N_13380,N_13636);
or U14401 (N_14401,N_13710,N_13317);
or U14402 (N_14402,N_13532,N_13651);
nand U14403 (N_14403,N_13223,N_13320);
nor U14404 (N_14404,N_13148,N_13738);
nand U14405 (N_14405,N_13882,N_13327);
or U14406 (N_14406,N_13292,N_13457);
xor U14407 (N_14407,N_13127,N_13117);
nor U14408 (N_14408,N_13588,N_13864);
or U14409 (N_14409,N_13627,N_13217);
nor U14410 (N_14410,N_13699,N_13062);
xor U14411 (N_14411,N_13229,N_13823);
and U14412 (N_14412,N_13817,N_13907);
nor U14413 (N_14413,N_13684,N_13842);
or U14414 (N_14414,N_13599,N_13431);
nor U14415 (N_14415,N_13053,N_13810);
nand U14416 (N_14416,N_13898,N_13324);
or U14417 (N_14417,N_13067,N_13917);
nor U14418 (N_14418,N_13356,N_13499);
xor U14419 (N_14419,N_13518,N_13993);
and U14420 (N_14420,N_13793,N_13131);
nor U14421 (N_14421,N_13795,N_13436);
nor U14422 (N_14422,N_13709,N_13243);
or U14423 (N_14423,N_13742,N_13950);
xnor U14424 (N_14424,N_13475,N_13137);
nor U14425 (N_14425,N_13614,N_13523);
or U14426 (N_14426,N_13824,N_13609);
and U14427 (N_14427,N_13480,N_13418);
and U14428 (N_14428,N_13314,N_13990);
nand U14429 (N_14429,N_13358,N_13417);
nand U14430 (N_14430,N_13029,N_13359);
nor U14431 (N_14431,N_13266,N_13251);
nor U14432 (N_14432,N_13605,N_13283);
xnor U14433 (N_14433,N_13049,N_13028);
or U14434 (N_14434,N_13209,N_13631);
and U14435 (N_14435,N_13524,N_13254);
xor U14436 (N_14436,N_13016,N_13077);
or U14437 (N_14437,N_13248,N_13155);
or U14438 (N_14438,N_13313,N_13315);
nor U14439 (N_14439,N_13472,N_13298);
nor U14440 (N_14440,N_13322,N_13207);
nand U14441 (N_14441,N_13798,N_13228);
or U14442 (N_14442,N_13944,N_13777);
nand U14443 (N_14443,N_13734,N_13556);
nor U14444 (N_14444,N_13846,N_13600);
nand U14445 (N_14445,N_13169,N_13332);
or U14446 (N_14446,N_13050,N_13376);
nand U14447 (N_14447,N_13516,N_13410);
and U14448 (N_14448,N_13736,N_13454);
and U14449 (N_14449,N_13608,N_13573);
and U14450 (N_14450,N_13246,N_13051);
nand U14451 (N_14451,N_13158,N_13722);
xor U14452 (N_14452,N_13973,N_13748);
and U14453 (N_14453,N_13604,N_13423);
nand U14454 (N_14454,N_13108,N_13712);
nand U14455 (N_14455,N_13304,N_13460);
nand U14456 (N_14456,N_13592,N_13095);
or U14457 (N_14457,N_13827,N_13548);
nor U14458 (N_14458,N_13852,N_13349);
or U14459 (N_14459,N_13492,N_13162);
nor U14460 (N_14460,N_13503,N_13406);
nor U14461 (N_14461,N_13772,N_13211);
or U14462 (N_14462,N_13790,N_13201);
nor U14463 (N_14463,N_13639,N_13043);
or U14464 (N_14464,N_13621,N_13268);
or U14465 (N_14465,N_13785,N_13902);
nor U14466 (N_14466,N_13336,N_13955);
nor U14467 (N_14467,N_13430,N_13215);
nand U14468 (N_14468,N_13027,N_13594);
nand U14469 (N_14469,N_13992,N_13432);
or U14470 (N_14470,N_13807,N_13644);
nand U14471 (N_14471,N_13528,N_13323);
nand U14472 (N_14472,N_13151,N_13112);
nand U14473 (N_14473,N_13435,N_13562);
nor U14474 (N_14474,N_13234,N_13976);
nor U14475 (N_14475,N_13719,N_13924);
nand U14476 (N_14476,N_13420,N_13369);
xnor U14477 (N_14477,N_13697,N_13849);
and U14478 (N_14478,N_13745,N_13287);
nand U14479 (N_14479,N_13497,N_13891);
and U14480 (N_14480,N_13520,N_13203);
and U14481 (N_14481,N_13366,N_13905);
nand U14482 (N_14482,N_13276,N_13895);
nand U14483 (N_14483,N_13185,N_13128);
or U14484 (N_14484,N_13561,N_13568);
nand U14485 (N_14485,N_13278,N_13555);
nor U14486 (N_14486,N_13111,N_13345);
or U14487 (N_14487,N_13113,N_13729);
or U14488 (N_14488,N_13869,N_13463);
xor U14489 (N_14489,N_13013,N_13858);
nand U14490 (N_14490,N_13630,N_13615);
and U14491 (N_14491,N_13297,N_13696);
nor U14492 (N_14492,N_13771,N_13885);
xor U14493 (N_14493,N_13301,N_13681);
nand U14494 (N_14494,N_13225,N_13755);
nand U14495 (N_14495,N_13026,N_13985);
xor U14496 (N_14496,N_13657,N_13747);
xor U14497 (N_14497,N_13489,N_13758);
or U14498 (N_14498,N_13202,N_13989);
nor U14499 (N_14499,N_13239,N_13886);
xor U14500 (N_14500,N_13190,N_13916);
or U14501 (N_14501,N_13099,N_13814);
nor U14502 (N_14502,N_13338,N_13398);
nor U14503 (N_14503,N_13992,N_13525);
nand U14504 (N_14504,N_13782,N_13714);
or U14505 (N_14505,N_13278,N_13438);
or U14506 (N_14506,N_13577,N_13839);
and U14507 (N_14507,N_13004,N_13332);
xnor U14508 (N_14508,N_13886,N_13541);
nand U14509 (N_14509,N_13136,N_13700);
and U14510 (N_14510,N_13222,N_13456);
nand U14511 (N_14511,N_13671,N_13652);
nand U14512 (N_14512,N_13333,N_13258);
and U14513 (N_14513,N_13627,N_13503);
and U14514 (N_14514,N_13020,N_13919);
nand U14515 (N_14515,N_13948,N_13258);
nand U14516 (N_14516,N_13679,N_13043);
and U14517 (N_14517,N_13716,N_13264);
and U14518 (N_14518,N_13485,N_13895);
and U14519 (N_14519,N_13572,N_13735);
and U14520 (N_14520,N_13400,N_13167);
xnor U14521 (N_14521,N_13339,N_13499);
and U14522 (N_14522,N_13732,N_13646);
nor U14523 (N_14523,N_13800,N_13072);
nand U14524 (N_14524,N_13145,N_13273);
nand U14525 (N_14525,N_13309,N_13526);
and U14526 (N_14526,N_13670,N_13966);
nor U14527 (N_14527,N_13563,N_13588);
and U14528 (N_14528,N_13848,N_13564);
nand U14529 (N_14529,N_13901,N_13574);
or U14530 (N_14530,N_13076,N_13390);
xor U14531 (N_14531,N_13952,N_13509);
or U14532 (N_14532,N_13614,N_13586);
and U14533 (N_14533,N_13379,N_13167);
or U14534 (N_14534,N_13907,N_13279);
and U14535 (N_14535,N_13661,N_13081);
or U14536 (N_14536,N_13802,N_13139);
nand U14537 (N_14537,N_13134,N_13614);
and U14538 (N_14538,N_13889,N_13855);
or U14539 (N_14539,N_13557,N_13563);
nand U14540 (N_14540,N_13919,N_13738);
and U14541 (N_14541,N_13554,N_13266);
or U14542 (N_14542,N_13011,N_13577);
and U14543 (N_14543,N_13309,N_13318);
and U14544 (N_14544,N_13330,N_13283);
nor U14545 (N_14545,N_13586,N_13467);
nand U14546 (N_14546,N_13201,N_13464);
or U14547 (N_14547,N_13402,N_13194);
or U14548 (N_14548,N_13766,N_13392);
nand U14549 (N_14549,N_13390,N_13350);
nand U14550 (N_14550,N_13474,N_13043);
nand U14551 (N_14551,N_13948,N_13561);
and U14552 (N_14552,N_13077,N_13984);
or U14553 (N_14553,N_13249,N_13528);
or U14554 (N_14554,N_13675,N_13111);
or U14555 (N_14555,N_13055,N_13528);
nor U14556 (N_14556,N_13496,N_13881);
nand U14557 (N_14557,N_13405,N_13295);
nand U14558 (N_14558,N_13123,N_13042);
and U14559 (N_14559,N_13835,N_13414);
and U14560 (N_14560,N_13107,N_13855);
and U14561 (N_14561,N_13958,N_13908);
xnor U14562 (N_14562,N_13284,N_13422);
and U14563 (N_14563,N_13469,N_13875);
and U14564 (N_14564,N_13069,N_13382);
or U14565 (N_14565,N_13886,N_13340);
nand U14566 (N_14566,N_13483,N_13024);
nand U14567 (N_14567,N_13829,N_13002);
xnor U14568 (N_14568,N_13889,N_13662);
or U14569 (N_14569,N_13408,N_13213);
nand U14570 (N_14570,N_13274,N_13987);
xor U14571 (N_14571,N_13618,N_13741);
and U14572 (N_14572,N_13930,N_13379);
xnor U14573 (N_14573,N_13269,N_13800);
or U14574 (N_14574,N_13758,N_13834);
and U14575 (N_14575,N_13582,N_13457);
xor U14576 (N_14576,N_13888,N_13725);
xor U14577 (N_14577,N_13191,N_13771);
nor U14578 (N_14578,N_13899,N_13613);
xnor U14579 (N_14579,N_13349,N_13725);
nand U14580 (N_14580,N_13601,N_13699);
xnor U14581 (N_14581,N_13457,N_13991);
or U14582 (N_14582,N_13625,N_13177);
and U14583 (N_14583,N_13487,N_13540);
or U14584 (N_14584,N_13026,N_13273);
or U14585 (N_14585,N_13193,N_13479);
or U14586 (N_14586,N_13041,N_13739);
nor U14587 (N_14587,N_13984,N_13224);
nor U14588 (N_14588,N_13264,N_13216);
nor U14589 (N_14589,N_13226,N_13461);
and U14590 (N_14590,N_13837,N_13405);
nand U14591 (N_14591,N_13457,N_13116);
xnor U14592 (N_14592,N_13882,N_13392);
or U14593 (N_14593,N_13407,N_13972);
or U14594 (N_14594,N_13845,N_13976);
xor U14595 (N_14595,N_13827,N_13743);
xnor U14596 (N_14596,N_13117,N_13327);
nand U14597 (N_14597,N_13891,N_13628);
or U14598 (N_14598,N_13587,N_13164);
nand U14599 (N_14599,N_13850,N_13112);
or U14600 (N_14600,N_13283,N_13146);
nand U14601 (N_14601,N_13433,N_13495);
nor U14602 (N_14602,N_13346,N_13654);
xnor U14603 (N_14603,N_13713,N_13460);
and U14604 (N_14604,N_13025,N_13796);
nand U14605 (N_14605,N_13833,N_13228);
and U14606 (N_14606,N_13312,N_13153);
xnor U14607 (N_14607,N_13398,N_13794);
and U14608 (N_14608,N_13219,N_13288);
nand U14609 (N_14609,N_13337,N_13560);
nor U14610 (N_14610,N_13258,N_13849);
and U14611 (N_14611,N_13750,N_13508);
or U14612 (N_14612,N_13046,N_13204);
nor U14613 (N_14613,N_13165,N_13925);
and U14614 (N_14614,N_13257,N_13442);
nor U14615 (N_14615,N_13376,N_13415);
and U14616 (N_14616,N_13367,N_13846);
nor U14617 (N_14617,N_13982,N_13501);
and U14618 (N_14618,N_13869,N_13057);
and U14619 (N_14619,N_13194,N_13800);
or U14620 (N_14620,N_13565,N_13497);
nor U14621 (N_14621,N_13058,N_13759);
nand U14622 (N_14622,N_13601,N_13484);
nand U14623 (N_14623,N_13392,N_13659);
and U14624 (N_14624,N_13053,N_13803);
nor U14625 (N_14625,N_13714,N_13169);
nand U14626 (N_14626,N_13168,N_13883);
or U14627 (N_14627,N_13625,N_13044);
nor U14628 (N_14628,N_13166,N_13066);
xor U14629 (N_14629,N_13893,N_13851);
nand U14630 (N_14630,N_13630,N_13652);
or U14631 (N_14631,N_13685,N_13849);
or U14632 (N_14632,N_13480,N_13356);
nand U14633 (N_14633,N_13604,N_13179);
xor U14634 (N_14634,N_13793,N_13674);
or U14635 (N_14635,N_13379,N_13552);
nand U14636 (N_14636,N_13215,N_13241);
nand U14637 (N_14637,N_13004,N_13584);
and U14638 (N_14638,N_13025,N_13663);
nor U14639 (N_14639,N_13978,N_13783);
or U14640 (N_14640,N_13299,N_13389);
xnor U14641 (N_14641,N_13596,N_13644);
nand U14642 (N_14642,N_13132,N_13566);
and U14643 (N_14643,N_13823,N_13406);
nand U14644 (N_14644,N_13974,N_13210);
xor U14645 (N_14645,N_13324,N_13329);
nor U14646 (N_14646,N_13792,N_13726);
nor U14647 (N_14647,N_13798,N_13005);
and U14648 (N_14648,N_13823,N_13616);
nand U14649 (N_14649,N_13513,N_13963);
or U14650 (N_14650,N_13682,N_13512);
or U14651 (N_14651,N_13069,N_13120);
and U14652 (N_14652,N_13946,N_13313);
or U14653 (N_14653,N_13484,N_13452);
and U14654 (N_14654,N_13488,N_13857);
nor U14655 (N_14655,N_13116,N_13580);
nor U14656 (N_14656,N_13311,N_13502);
nor U14657 (N_14657,N_13120,N_13067);
or U14658 (N_14658,N_13426,N_13512);
xnor U14659 (N_14659,N_13496,N_13933);
nor U14660 (N_14660,N_13297,N_13982);
nand U14661 (N_14661,N_13108,N_13756);
and U14662 (N_14662,N_13215,N_13107);
and U14663 (N_14663,N_13883,N_13680);
xor U14664 (N_14664,N_13097,N_13601);
nor U14665 (N_14665,N_13228,N_13132);
and U14666 (N_14666,N_13149,N_13151);
and U14667 (N_14667,N_13832,N_13891);
nor U14668 (N_14668,N_13127,N_13597);
nand U14669 (N_14669,N_13585,N_13586);
nand U14670 (N_14670,N_13832,N_13282);
nor U14671 (N_14671,N_13453,N_13862);
and U14672 (N_14672,N_13324,N_13777);
xor U14673 (N_14673,N_13827,N_13305);
xor U14674 (N_14674,N_13494,N_13700);
or U14675 (N_14675,N_13892,N_13979);
nor U14676 (N_14676,N_13934,N_13315);
or U14677 (N_14677,N_13656,N_13948);
or U14678 (N_14678,N_13956,N_13801);
and U14679 (N_14679,N_13920,N_13610);
and U14680 (N_14680,N_13869,N_13832);
and U14681 (N_14681,N_13615,N_13076);
nand U14682 (N_14682,N_13019,N_13618);
and U14683 (N_14683,N_13955,N_13626);
or U14684 (N_14684,N_13152,N_13536);
and U14685 (N_14685,N_13661,N_13785);
nand U14686 (N_14686,N_13550,N_13689);
xnor U14687 (N_14687,N_13825,N_13913);
nand U14688 (N_14688,N_13300,N_13421);
or U14689 (N_14689,N_13661,N_13228);
nor U14690 (N_14690,N_13439,N_13597);
or U14691 (N_14691,N_13252,N_13895);
and U14692 (N_14692,N_13240,N_13092);
xnor U14693 (N_14693,N_13572,N_13184);
nand U14694 (N_14694,N_13402,N_13492);
nand U14695 (N_14695,N_13369,N_13668);
nand U14696 (N_14696,N_13623,N_13810);
nand U14697 (N_14697,N_13030,N_13874);
xnor U14698 (N_14698,N_13618,N_13359);
nor U14699 (N_14699,N_13505,N_13292);
and U14700 (N_14700,N_13962,N_13627);
nand U14701 (N_14701,N_13237,N_13413);
nand U14702 (N_14702,N_13680,N_13763);
nand U14703 (N_14703,N_13089,N_13190);
and U14704 (N_14704,N_13313,N_13637);
nor U14705 (N_14705,N_13908,N_13829);
nand U14706 (N_14706,N_13895,N_13726);
or U14707 (N_14707,N_13534,N_13066);
or U14708 (N_14708,N_13467,N_13289);
and U14709 (N_14709,N_13199,N_13158);
nand U14710 (N_14710,N_13729,N_13963);
and U14711 (N_14711,N_13612,N_13969);
nor U14712 (N_14712,N_13994,N_13880);
xor U14713 (N_14713,N_13308,N_13681);
nand U14714 (N_14714,N_13150,N_13770);
nand U14715 (N_14715,N_13590,N_13589);
nor U14716 (N_14716,N_13774,N_13018);
and U14717 (N_14717,N_13050,N_13238);
or U14718 (N_14718,N_13956,N_13542);
and U14719 (N_14719,N_13451,N_13174);
and U14720 (N_14720,N_13709,N_13653);
or U14721 (N_14721,N_13432,N_13821);
nand U14722 (N_14722,N_13136,N_13732);
xor U14723 (N_14723,N_13880,N_13333);
nor U14724 (N_14724,N_13182,N_13355);
and U14725 (N_14725,N_13206,N_13876);
nand U14726 (N_14726,N_13152,N_13283);
xor U14727 (N_14727,N_13082,N_13860);
nand U14728 (N_14728,N_13845,N_13632);
nor U14729 (N_14729,N_13438,N_13886);
xnor U14730 (N_14730,N_13281,N_13713);
or U14731 (N_14731,N_13494,N_13702);
and U14732 (N_14732,N_13852,N_13033);
nor U14733 (N_14733,N_13469,N_13745);
nor U14734 (N_14734,N_13355,N_13524);
or U14735 (N_14735,N_13672,N_13282);
nand U14736 (N_14736,N_13929,N_13437);
and U14737 (N_14737,N_13610,N_13345);
nor U14738 (N_14738,N_13631,N_13131);
or U14739 (N_14739,N_13702,N_13710);
and U14740 (N_14740,N_13458,N_13883);
nor U14741 (N_14741,N_13478,N_13083);
or U14742 (N_14742,N_13381,N_13666);
and U14743 (N_14743,N_13149,N_13410);
nand U14744 (N_14744,N_13965,N_13516);
nand U14745 (N_14745,N_13042,N_13607);
nor U14746 (N_14746,N_13069,N_13044);
nor U14747 (N_14747,N_13385,N_13929);
or U14748 (N_14748,N_13343,N_13159);
and U14749 (N_14749,N_13107,N_13902);
and U14750 (N_14750,N_13874,N_13890);
nand U14751 (N_14751,N_13665,N_13289);
or U14752 (N_14752,N_13751,N_13573);
nor U14753 (N_14753,N_13981,N_13419);
xnor U14754 (N_14754,N_13445,N_13407);
nand U14755 (N_14755,N_13771,N_13070);
or U14756 (N_14756,N_13992,N_13976);
nor U14757 (N_14757,N_13459,N_13043);
nand U14758 (N_14758,N_13091,N_13445);
nand U14759 (N_14759,N_13206,N_13372);
or U14760 (N_14760,N_13612,N_13825);
nand U14761 (N_14761,N_13049,N_13504);
xnor U14762 (N_14762,N_13076,N_13965);
nand U14763 (N_14763,N_13382,N_13786);
xor U14764 (N_14764,N_13058,N_13360);
and U14765 (N_14765,N_13765,N_13315);
and U14766 (N_14766,N_13242,N_13730);
nor U14767 (N_14767,N_13476,N_13552);
nor U14768 (N_14768,N_13995,N_13578);
nand U14769 (N_14769,N_13051,N_13060);
nor U14770 (N_14770,N_13851,N_13850);
xnor U14771 (N_14771,N_13718,N_13287);
and U14772 (N_14772,N_13873,N_13442);
nor U14773 (N_14773,N_13640,N_13007);
xor U14774 (N_14774,N_13425,N_13170);
xor U14775 (N_14775,N_13079,N_13202);
nor U14776 (N_14776,N_13783,N_13906);
nand U14777 (N_14777,N_13576,N_13434);
nand U14778 (N_14778,N_13600,N_13498);
nand U14779 (N_14779,N_13808,N_13360);
and U14780 (N_14780,N_13177,N_13872);
xor U14781 (N_14781,N_13999,N_13851);
nand U14782 (N_14782,N_13733,N_13027);
nor U14783 (N_14783,N_13123,N_13867);
nand U14784 (N_14784,N_13821,N_13175);
xor U14785 (N_14785,N_13562,N_13400);
nor U14786 (N_14786,N_13878,N_13166);
and U14787 (N_14787,N_13846,N_13719);
xor U14788 (N_14788,N_13671,N_13073);
xnor U14789 (N_14789,N_13574,N_13216);
and U14790 (N_14790,N_13722,N_13067);
nor U14791 (N_14791,N_13583,N_13632);
xnor U14792 (N_14792,N_13555,N_13251);
xnor U14793 (N_14793,N_13829,N_13898);
and U14794 (N_14794,N_13972,N_13343);
nor U14795 (N_14795,N_13214,N_13294);
nand U14796 (N_14796,N_13166,N_13945);
xnor U14797 (N_14797,N_13072,N_13728);
or U14798 (N_14798,N_13272,N_13433);
nand U14799 (N_14799,N_13371,N_13478);
or U14800 (N_14800,N_13818,N_13160);
or U14801 (N_14801,N_13328,N_13724);
nand U14802 (N_14802,N_13942,N_13857);
xor U14803 (N_14803,N_13919,N_13829);
or U14804 (N_14804,N_13098,N_13134);
and U14805 (N_14805,N_13589,N_13381);
and U14806 (N_14806,N_13195,N_13458);
or U14807 (N_14807,N_13335,N_13880);
or U14808 (N_14808,N_13862,N_13208);
nand U14809 (N_14809,N_13228,N_13024);
nor U14810 (N_14810,N_13980,N_13573);
nand U14811 (N_14811,N_13759,N_13532);
xnor U14812 (N_14812,N_13772,N_13485);
nand U14813 (N_14813,N_13988,N_13532);
or U14814 (N_14814,N_13619,N_13743);
xor U14815 (N_14815,N_13109,N_13428);
and U14816 (N_14816,N_13027,N_13677);
and U14817 (N_14817,N_13422,N_13106);
xor U14818 (N_14818,N_13591,N_13499);
xnor U14819 (N_14819,N_13649,N_13641);
nor U14820 (N_14820,N_13866,N_13808);
or U14821 (N_14821,N_13167,N_13958);
nor U14822 (N_14822,N_13182,N_13433);
nand U14823 (N_14823,N_13824,N_13727);
nand U14824 (N_14824,N_13155,N_13093);
or U14825 (N_14825,N_13259,N_13019);
or U14826 (N_14826,N_13759,N_13952);
nor U14827 (N_14827,N_13057,N_13182);
and U14828 (N_14828,N_13878,N_13531);
and U14829 (N_14829,N_13432,N_13161);
nand U14830 (N_14830,N_13485,N_13177);
and U14831 (N_14831,N_13134,N_13596);
or U14832 (N_14832,N_13732,N_13740);
xor U14833 (N_14833,N_13303,N_13526);
or U14834 (N_14834,N_13292,N_13189);
nand U14835 (N_14835,N_13135,N_13663);
or U14836 (N_14836,N_13516,N_13003);
xor U14837 (N_14837,N_13110,N_13616);
or U14838 (N_14838,N_13031,N_13225);
or U14839 (N_14839,N_13600,N_13475);
or U14840 (N_14840,N_13215,N_13523);
nand U14841 (N_14841,N_13088,N_13843);
and U14842 (N_14842,N_13475,N_13879);
nand U14843 (N_14843,N_13943,N_13948);
and U14844 (N_14844,N_13163,N_13168);
nor U14845 (N_14845,N_13997,N_13732);
nand U14846 (N_14846,N_13236,N_13234);
and U14847 (N_14847,N_13606,N_13881);
nor U14848 (N_14848,N_13739,N_13461);
or U14849 (N_14849,N_13569,N_13474);
nor U14850 (N_14850,N_13103,N_13507);
and U14851 (N_14851,N_13627,N_13328);
and U14852 (N_14852,N_13485,N_13120);
or U14853 (N_14853,N_13479,N_13695);
and U14854 (N_14854,N_13555,N_13704);
or U14855 (N_14855,N_13485,N_13034);
nor U14856 (N_14856,N_13949,N_13766);
nand U14857 (N_14857,N_13701,N_13618);
or U14858 (N_14858,N_13487,N_13351);
or U14859 (N_14859,N_13500,N_13111);
nand U14860 (N_14860,N_13994,N_13384);
xor U14861 (N_14861,N_13157,N_13554);
nand U14862 (N_14862,N_13475,N_13576);
nor U14863 (N_14863,N_13353,N_13639);
nand U14864 (N_14864,N_13970,N_13040);
xor U14865 (N_14865,N_13534,N_13835);
nand U14866 (N_14866,N_13551,N_13144);
nor U14867 (N_14867,N_13015,N_13155);
nor U14868 (N_14868,N_13204,N_13088);
nand U14869 (N_14869,N_13314,N_13022);
and U14870 (N_14870,N_13283,N_13891);
or U14871 (N_14871,N_13783,N_13565);
and U14872 (N_14872,N_13308,N_13730);
nand U14873 (N_14873,N_13189,N_13220);
xor U14874 (N_14874,N_13069,N_13894);
nor U14875 (N_14875,N_13203,N_13853);
and U14876 (N_14876,N_13644,N_13548);
nor U14877 (N_14877,N_13472,N_13335);
and U14878 (N_14878,N_13356,N_13706);
or U14879 (N_14879,N_13073,N_13807);
nand U14880 (N_14880,N_13614,N_13169);
or U14881 (N_14881,N_13922,N_13818);
and U14882 (N_14882,N_13522,N_13078);
nor U14883 (N_14883,N_13266,N_13924);
and U14884 (N_14884,N_13977,N_13923);
nor U14885 (N_14885,N_13758,N_13442);
or U14886 (N_14886,N_13531,N_13416);
and U14887 (N_14887,N_13447,N_13769);
and U14888 (N_14888,N_13257,N_13352);
or U14889 (N_14889,N_13388,N_13622);
nand U14890 (N_14890,N_13455,N_13029);
and U14891 (N_14891,N_13207,N_13796);
nor U14892 (N_14892,N_13710,N_13910);
and U14893 (N_14893,N_13097,N_13805);
nor U14894 (N_14894,N_13652,N_13627);
nor U14895 (N_14895,N_13817,N_13025);
and U14896 (N_14896,N_13724,N_13623);
nand U14897 (N_14897,N_13683,N_13230);
or U14898 (N_14898,N_13861,N_13766);
or U14899 (N_14899,N_13297,N_13922);
and U14900 (N_14900,N_13595,N_13214);
xnor U14901 (N_14901,N_13762,N_13842);
nor U14902 (N_14902,N_13092,N_13458);
nor U14903 (N_14903,N_13116,N_13509);
nor U14904 (N_14904,N_13366,N_13533);
nor U14905 (N_14905,N_13572,N_13093);
and U14906 (N_14906,N_13672,N_13353);
or U14907 (N_14907,N_13127,N_13759);
nor U14908 (N_14908,N_13918,N_13163);
nor U14909 (N_14909,N_13086,N_13415);
and U14910 (N_14910,N_13833,N_13247);
and U14911 (N_14911,N_13837,N_13860);
nor U14912 (N_14912,N_13093,N_13932);
nand U14913 (N_14913,N_13776,N_13779);
nand U14914 (N_14914,N_13930,N_13829);
or U14915 (N_14915,N_13720,N_13718);
nor U14916 (N_14916,N_13171,N_13005);
or U14917 (N_14917,N_13084,N_13446);
and U14918 (N_14918,N_13550,N_13323);
nor U14919 (N_14919,N_13485,N_13009);
nor U14920 (N_14920,N_13886,N_13197);
xor U14921 (N_14921,N_13819,N_13611);
and U14922 (N_14922,N_13928,N_13612);
and U14923 (N_14923,N_13876,N_13462);
nor U14924 (N_14924,N_13829,N_13026);
nor U14925 (N_14925,N_13109,N_13487);
nand U14926 (N_14926,N_13271,N_13805);
and U14927 (N_14927,N_13815,N_13148);
or U14928 (N_14928,N_13468,N_13264);
xor U14929 (N_14929,N_13658,N_13413);
or U14930 (N_14930,N_13002,N_13904);
xnor U14931 (N_14931,N_13789,N_13197);
and U14932 (N_14932,N_13409,N_13993);
nor U14933 (N_14933,N_13206,N_13133);
nand U14934 (N_14934,N_13157,N_13617);
nand U14935 (N_14935,N_13096,N_13061);
nor U14936 (N_14936,N_13802,N_13540);
and U14937 (N_14937,N_13106,N_13380);
or U14938 (N_14938,N_13337,N_13223);
or U14939 (N_14939,N_13549,N_13693);
nor U14940 (N_14940,N_13286,N_13181);
nand U14941 (N_14941,N_13900,N_13689);
nand U14942 (N_14942,N_13623,N_13491);
nor U14943 (N_14943,N_13047,N_13641);
or U14944 (N_14944,N_13438,N_13554);
nor U14945 (N_14945,N_13803,N_13048);
nor U14946 (N_14946,N_13728,N_13834);
and U14947 (N_14947,N_13915,N_13519);
or U14948 (N_14948,N_13639,N_13785);
nand U14949 (N_14949,N_13266,N_13021);
nor U14950 (N_14950,N_13882,N_13726);
and U14951 (N_14951,N_13227,N_13922);
nand U14952 (N_14952,N_13111,N_13832);
nor U14953 (N_14953,N_13402,N_13210);
nand U14954 (N_14954,N_13820,N_13706);
xnor U14955 (N_14955,N_13519,N_13175);
and U14956 (N_14956,N_13955,N_13509);
xnor U14957 (N_14957,N_13966,N_13691);
or U14958 (N_14958,N_13285,N_13618);
nor U14959 (N_14959,N_13587,N_13432);
or U14960 (N_14960,N_13308,N_13989);
and U14961 (N_14961,N_13309,N_13236);
or U14962 (N_14962,N_13808,N_13532);
nor U14963 (N_14963,N_13077,N_13826);
and U14964 (N_14964,N_13882,N_13431);
and U14965 (N_14965,N_13065,N_13213);
nor U14966 (N_14966,N_13107,N_13708);
or U14967 (N_14967,N_13292,N_13320);
nor U14968 (N_14968,N_13108,N_13151);
or U14969 (N_14969,N_13437,N_13659);
nor U14970 (N_14970,N_13366,N_13890);
nand U14971 (N_14971,N_13385,N_13643);
or U14972 (N_14972,N_13391,N_13424);
nand U14973 (N_14973,N_13922,N_13365);
and U14974 (N_14974,N_13995,N_13075);
nand U14975 (N_14975,N_13511,N_13823);
xor U14976 (N_14976,N_13585,N_13169);
and U14977 (N_14977,N_13947,N_13306);
nor U14978 (N_14978,N_13684,N_13401);
nor U14979 (N_14979,N_13420,N_13424);
and U14980 (N_14980,N_13184,N_13224);
and U14981 (N_14981,N_13855,N_13742);
nand U14982 (N_14982,N_13222,N_13779);
nor U14983 (N_14983,N_13153,N_13532);
or U14984 (N_14984,N_13820,N_13225);
or U14985 (N_14985,N_13270,N_13580);
xnor U14986 (N_14986,N_13460,N_13472);
nand U14987 (N_14987,N_13089,N_13294);
or U14988 (N_14988,N_13591,N_13080);
and U14989 (N_14989,N_13503,N_13021);
and U14990 (N_14990,N_13646,N_13225);
nand U14991 (N_14991,N_13048,N_13043);
nor U14992 (N_14992,N_13350,N_13913);
nand U14993 (N_14993,N_13915,N_13326);
nand U14994 (N_14994,N_13121,N_13534);
and U14995 (N_14995,N_13282,N_13668);
nor U14996 (N_14996,N_13690,N_13600);
and U14997 (N_14997,N_13401,N_13932);
nor U14998 (N_14998,N_13642,N_13927);
nor U14999 (N_14999,N_13090,N_13929);
nand UO_0 (O_0,N_14613,N_14024);
or UO_1 (O_1,N_14140,N_14513);
xor UO_2 (O_2,N_14167,N_14102);
nand UO_3 (O_3,N_14837,N_14303);
nand UO_4 (O_4,N_14236,N_14659);
nor UO_5 (O_5,N_14630,N_14302);
nor UO_6 (O_6,N_14903,N_14571);
or UO_7 (O_7,N_14436,N_14652);
and UO_8 (O_8,N_14979,N_14769);
or UO_9 (O_9,N_14395,N_14737);
or UO_10 (O_10,N_14381,N_14095);
nor UO_11 (O_11,N_14676,N_14271);
or UO_12 (O_12,N_14727,N_14614);
nor UO_13 (O_13,N_14075,N_14404);
nand UO_14 (O_14,N_14914,N_14782);
and UO_15 (O_15,N_14699,N_14774);
nor UO_16 (O_16,N_14124,N_14161);
nand UO_17 (O_17,N_14537,N_14834);
and UO_18 (O_18,N_14215,N_14087);
or UO_19 (O_19,N_14157,N_14940);
and UO_20 (O_20,N_14870,N_14094);
or UO_21 (O_21,N_14581,N_14410);
or UO_22 (O_22,N_14309,N_14246);
nand UO_23 (O_23,N_14068,N_14627);
nor UO_24 (O_24,N_14883,N_14665);
or UO_25 (O_25,N_14781,N_14437);
nor UO_26 (O_26,N_14120,N_14864);
nand UO_27 (O_27,N_14162,N_14447);
nor UO_28 (O_28,N_14748,N_14625);
nand UO_29 (O_29,N_14229,N_14304);
nor UO_30 (O_30,N_14424,N_14214);
or UO_31 (O_31,N_14143,N_14399);
and UO_32 (O_32,N_14792,N_14487);
nor UO_33 (O_33,N_14108,N_14929);
and UO_34 (O_34,N_14560,N_14921);
nor UO_35 (O_35,N_14975,N_14474);
and UO_36 (O_36,N_14242,N_14556);
or UO_37 (O_37,N_14319,N_14298);
nor UO_38 (O_38,N_14517,N_14357);
or UO_39 (O_39,N_14709,N_14023);
and UO_40 (O_40,N_14502,N_14086);
nand UO_41 (O_41,N_14322,N_14606);
and UO_42 (O_42,N_14189,N_14332);
nor UO_43 (O_43,N_14127,N_14377);
or UO_44 (O_44,N_14547,N_14478);
and UO_45 (O_45,N_14635,N_14551);
and UO_46 (O_46,N_14380,N_14412);
nand UO_47 (O_47,N_14053,N_14706);
nand UO_48 (O_48,N_14969,N_14186);
nand UO_49 (O_49,N_14582,N_14018);
nand UO_50 (O_50,N_14958,N_14907);
nand UO_51 (O_51,N_14790,N_14240);
nand UO_52 (O_52,N_14360,N_14476);
nand UO_53 (O_53,N_14388,N_14374);
or UO_54 (O_54,N_14937,N_14521);
or UO_55 (O_55,N_14378,N_14671);
nor UO_56 (O_56,N_14558,N_14961);
and UO_57 (O_57,N_14924,N_14664);
or UO_58 (O_58,N_14421,N_14029);
and UO_59 (O_59,N_14799,N_14464);
and UO_60 (O_60,N_14829,N_14997);
or UO_61 (O_61,N_14225,N_14529);
nand UO_62 (O_62,N_14310,N_14758);
nor UO_63 (O_63,N_14454,N_14411);
nor UO_64 (O_64,N_14221,N_14123);
nand UO_65 (O_65,N_14099,N_14599);
nor UO_66 (O_66,N_14072,N_14836);
or UO_67 (O_67,N_14314,N_14052);
nor UO_68 (O_68,N_14469,N_14237);
nor UO_69 (O_69,N_14500,N_14512);
nand UO_70 (O_70,N_14909,N_14065);
nor UO_71 (O_71,N_14020,N_14441);
and UO_72 (O_72,N_14701,N_14363);
nor UO_73 (O_73,N_14337,N_14753);
xor UO_74 (O_74,N_14180,N_14058);
and UO_75 (O_75,N_14900,N_14384);
or UO_76 (O_76,N_14771,N_14735);
and UO_77 (O_77,N_14467,N_14848);
xnor UO_78 (O_78,N_14603,N_14498);
xnor UO_79 (O_79,N_14700,N_14037);
or UO_80 (O_80,N_14455,N_14986);
or UO_81 (O_81,N_14504,N_14187);
or UO_82 (O_82,N_14823,N_14389);
or UO_83 (O_83,N_14165,N_14861);
nor UO_84 (O_84,N_14150,N_14159);
nand UO_85 (O_85,N_14543,N_14015);
xnor UO_86 (O_86,N_14062,N_14256);
nand UO_87 (O_87,N_14845,N_14146);
or UO_88 (O_88,N_14433,N_14089);
and UO_89 (O_89,N_14001,N_14561);
and UO_90 (O_90,N_14098,N_14260);
or UO_91 (O_91,N_14922,N_14335);
nand UO_92 (O_92,N_14448,N_14041);
nor UO_93 (O_93,N_14249,N_14695);
and UO_94 (O_94,N_14207,N_14947);
nand UO_95 (O_95,N_14341,N_14925);
or UO_96 (O_96,N_14767,N_14873);
or UO_97 (O_97,N_14876,N_14773);
and UO_98 (O_98,N_14682,N_14672);
nand UO_99 (O_99,N_14675,N_14830);
and UO_100 (O_100,N_14141,N_14882);
nor UO_101 (O_101,N_14879,N_14716);
nand UO_102 (O_102,N_14253,N_14283);
nand UO_103 (O_103,N_14164,N_14546);
and UO_104 (O_104,N_14756,N_14567);
and UO_105 (O_105,N_14850,N_14577);
or UO_106 (O_106,N_14480,N_14393);
or UO_107 (O_107,N_14936,N_14601);
nor UO_108 (O_108,N_14645,N_14524);
nand UO_109 (O_109,N_14134,N_14745);
or UO_110 (O_110,N_14609,N_14431);
and UO_111 (O_111,N_14730,N_14515);
or UO_112 (O_112,N_14422,N_14438);
or UO_113 (O_113,N_14895,N_14465);
xnor UO_114 (O_114,N_14807,N_14538);
nand UO_115 (O_115,N_14586,N_14295);
or UO_116 (O_116,N_14373,N_14083);
nor UO_117 (O_117,N_14550,N_14638);
nand UO_118 (O_118,N_14181,N_14928);
or UO_119 (O_119,N_14359,N_14149);
nor UO_120 (O_120,N_14854,N_14640);
or UO_121 (O_121,N_14163,N_14276);
nand UO_122 (O_122,N_14982,N_14172);
or UO_123 (O_123,N_14797,N_14043);
and UO_124 (O_124,N_14840,N_14235);
xor UO_125 (O_125,N_14579,N_14796);
and UO_126 (O_126,N_14416,N_14967);
or UO_127 (O_127,N_14770,N_14604);
or UO_128 (O_128,N_14950,N_14628);
xor UO_129 (O_129,N_14230,N_14270);
nor UO_130 (O_130,N_14791,N_14398);
nand UO_131 (O_131,N_14691,N_14281);
nand UO_132 (O_132,N_14642,N_14336);
and UO_133 (O_133,N_14911,N_14046);
or UO_134 (O_134,N_14492,N_14009);
or UO_135 (O_135,N_14852,N_14832);
nor UO_136 (O_136,N_14152,N_14254);
nor UO_137 (O_137,N_14918,N_14494);
nand UO_138 (O_138,N_14194,N_14689);
xor UO_139 (O_139,N_14503,N_14472);
nand UO_140 (O_140,N_14802,N_14554);
and UO_141 (O_141,N_14949,N_14425);
and UO_142 (O_142,N_14044,N_14368);
or UO_143 (O_143,N_14347,N_14875);
xnor UO_144 (O_144,N_14200,N_14430);
or UO_145 (O_145,N_14833,N_14592);
xor UO_146 (O_146,N_14803,N_14632);
or UO_147 (O_147,N_14618,N_14477);
and UO_148 (O_148,N_14941,N_14865);
nand UO_149 (O_149,N_14012,N_14506);
nor UO_150 (O_150,N_14564,N_14060);
xor UO_151 (O_151,N_14468,N_14419);
nor UO_152 (O_152,N_14261,N_14764);
nor UO_153 (O_153,N_14725,N_14344);
or UO_154 (O_154,N_14429,N_14305);
or UO_155 (O_155,N_14541,N_14483);
or UO_156 (O_156,N_14598,N_14247);
nand UO_157 (O_157,N_14401,N_14135);
and UO_158 (O_158,N_14884,N_14788);
and UO_159 (O_159,N_14209,N_14809);
or UO_160 (O_160,N_14101,N_14473);
and UO_161 (O_161,N_14106,N_14100);
nor UO_162 (O_162,N_14731,N_14435);
nand UO_163 (O_163,N_14703,N_14973);
or UO_164 (O_164,N_14039,N_14501);
nand UO_165 (O_165,N_14996,N_14348);
nand UO_166 (O_166,N_14536,N_14461);
and UO_167 (O_167,N_14655,N_14821);
or UO_168 (O_168,N_14905,N_14712);
and UO_169 (O_169,N_14623,N_14596);
and UO_170 (O_170,N_14131,N_14128);
and UO_171 (O_171,N_14456,N_14828);
and UO_172 (O_172,N_14277,N_14103);
and UO_173 (O_173,N_14514,N_14813);
nand UO_174 (O_174,N_14499,N_14413);
and UO_175 (O_175,N_14130,N_14148);
or UO_176 (O_176,N_14216,N_14654);
or UO_177 (O_177,N_14219,N_14831);
and UO_178 (O_178,N_14602,N_14000);
or UO_179 (O_179,N_14780,N_14213);
or UO_180 (O_180,N_14077,N_14228);
or UO_181 (O_181,N_14858,N_14853);
nand UO_182 (O_182,N_14508,N_14061);
nand UO_183 (O_183,N_14051,N_14226);
and UO_184 (O_184,N_14463,N_14066);
nor UO_185 (O_185,N_14375,N_14734);
or UO_186 (O_186,N_14010,N_14370);
nand UO_187 (O_187,N_14278,N_14316);
or UO_188 (O_188,N_14129,N_14170);
or UO_189 (O_189,N_14785,N_14805);
nor UO_190 (O_190,N_14174,N_14339);
nor UO_191 (O_191,N_14810,N_14290);
or UO_192 (O_192,N_14003,N_14379);
and UO_193 (O_193,N_14588,N_14679);
or UO_194 (O_194,N_14743,N_14386);
or UO_195 (O_195,N_14005,N_14136);
nor UO_196 (O_196,N_14451,N_14585);
and UO_197 (O_197,N_14594,N_14400);
xor UO_198 (O_198,N_14205,N_14442);
nand UO_199 (O_199,N_14568,N_14783);
nand UO_200 (O_200,N_14917,N_14634);
nor UO_201 (O_201,N_14479,N_14739);
and UO_202 (O_202,N_14491,N_14485);
nand UO_203 (O_203,N_14522,N_14651);
nand UO_204 (O_204,N_14184,N_14202);
or UO_205 (O_205,N_14307,N_14637);
xnor UO_206 (O_206,N_14763,N_14825);
nand UO_207 (O_207,N_14067,N_14275);
nand UO_208 (O_208,N_14574,N_14816);
nand UO_209 (O_209,N_14239,N_14292);
and UO_210 (O_210,N_14778,N_14656);
and UO_211 (O_211,N_14391,N_14624);
nand UO_212 (O_212,N_14121,N_14443);
and UO_213 (O_213,N_14999,N_14284);
and UO_214 (O_214,N_14583,N_14683);
and UO_215 (O_215,N_14251,N_14680);
nand UO_216 (O_216,N_14263,N_14231);
xor UO_217 (O_217,N_14318,N_14266);
nor UO_218 (O_218,N_14084,N_14877);
xnor UO_219 (O_219,N_14173,N_14971);
nor UO_220 (O_220,N_14153,N_14880);
and UO_221 (O_221,N_14484,N_14233);
or UO_222 (O_222,N_14063,N_14607);
nor UO_223 (O_223,N_14686,N_14608);
nor UO_224 (O_224,N_14578,N_14203);
xor UO_225 (O_225,N_14262,N_14033);
xnor UO_226 (O_226,N_14432,N_14715);
nor UO_227 (O_227,N_14736,N_14926);
nand UO_228 (O_228,N_14533,N_14022);
and UO_229 (O_229,N_14587,N_14862);
nor UO_230 (O_230,N_14320,N_14252);
or UO_231 (O_231,N_14509,N_14078);
nand UO_232 (O_232,N_14976,N_14188);
nand UO_233 (O_233,N_14641,N_14273);
nand UO_234 (O_234,N_14315,N_14396);
nor UO_235 (O_235,N_14698,N_14025);
or UO_236 (O_236,N_14299,N_14201);
xor UO_237 (O_237,N_14939,N_14994);
and UO_238 (O_238,N_14409,N_14932);
nor UO_239 (O_239,N_14032,N_14555);
nand UO_240 (O_240,N_14620,N_14017);
xor UO_241 (O_241,N_14705,N_14049);
nor UO_242 (O_242,N_14789,N_14800);
nand UO_243 (O_243,N_14376,N_14662);
or UO_244 (O_244,N_14863,N_14684);
or UO_245 (O_245,N_14050,N_14394);
xnor UO_246 (O_246,N_14096,N_14144);
nor UO_247 (O_247,N_14460,N_14542);
or UO_248 (O_248,N_14415,N_14245);
or UO_249 (O_249,N_14064,N_14570);
or UO_250 (O_250,N_14697,N_14666);
xor UO_251 (O_251,N_14372,N_14718);
nand UO_252 (O_252,N_14387,N_14330);
nand UO_253 (O_253,N_14747,N_14449);
or UO_254 (O_254,N_14016,N_14989);
and UO_255 (O_255,N_14338,N_14346);
nand UO_256 (O_256,N_14227,N_14944);
and UO_257 (O_257,N_14563,N_14343);
or UO_258 (O_258,N_14274,N_14311);
and UO_259 (O_259,N_14211,N_14943);
nor UO_260 (O_260,N_14324,N_14857);
or UO_261 (O_261,N_14729,N_14667);
and UO_262 (O_262,N_14351,N_14107);
or UO_263 (O_263,N_14297,N_14647);
and UO_264 (O_264,N_14321,N_14927);
xor UO_265 (O_265,N_14768,N_14220);
and UO_266 (O_266,N_14369,N_14912);
or UO_267 (O_267,N_14931,N_14964);
nor UO_268 (O_268,N_14361,N_14794);
nor UO_269 (O_269,N_14968,N_14553);
or UO_270 (O_270,N_14294,N_14125);
xnor UO_271 (O_271,N_14080,N_14983);
nand UO_272 (O_272,N_14855,N_14471);
or UO_273 (O_273,N_14616,N_14030);
nand UO_274 (O_274,N_14291,N_14019);
and UO_275 (O_275,N_14045,N_14113);
nor UO_276 (O_276,N_14817,N_14988);
and UO_277 (O_277,N_14722,N_14754);
and UO_278 (O_278,N_14728,N_14629);
or UO_279 (O_279,N_14757,N_14403);
or UO_280 (O_280,N_14779,N_14566);
nand UO_281 (O_281,N_14279,N_14866);
nand UO_282 (O_282,N_14523,N_14268);
nand UO_283 (O_283,N_14908,N_14349);
and UO_284 (O_284,N_14688,N_14289);
nand UO_285 (O_285,N_14147,N_14804);
or UO_286 (O_286,N_14074,N_14511);
or UO_287 (O_287,N_14933,N_14660);
or UO_288 (O_288,N_14327,N_14674);
nor UO_289 (O_289,N_14693,N_14902);
nand UO_290 (O_290,N_14385,N_14462);
xnor UO_291 (O_291,N_14137,N_14955);
nor UO_292 (O_292,N_14356,N_14114);
nand UO_293 (O_293,N_14977,N_14923);
nor UO_294 (O_294,N_14364,N_14827);
and UO_295 (O_295,N_14946,N_14169);
nand UO_296 (O_296,N_14942,N_14985);
nand UO_297 (O_297,N_14844,N_14034);
nand UO_298 (O_298,N_14992,N_14450);
nand UO_299 (O_299,N_14573,N_14871);
xor UO_300 (O_300,N_14822,N_14481);
xor UO_301 (O_301,N_14459,N_14612);
and UO_302 (O_302,N_14591,N_14076);
nand UO_303 (O_303,N_14259,N_14160);
xor UO_304 (O_304,N_14138,N_14913);
nor UO_305 (O_305,N_14183,N_14258);
or UO_306 (O_306,N_14264,N_14085);
and UO_307 (O_307,N_14826,N_14520);
or UO_308 (O_308,N_14584,N_14562);
or UO_309 (O_309,N_14595,N_14819);
nand UO_310 (O_310,N_14525,N_14057);
nor UO_311 (O_311,N_14678,N_14255);
nand UO_312 (O_312,N_14945,N_14109);
nand UO_313 (O_313,N_14742,N_14286);
and UO_314 (O_314,N_14856,N_14453);
and UO_315 (O_315,N_14593,N_14663);
nor UO_316 (O_316,N_14177,N_14151);
or UO_317 (O_317,N_14991,N_14518);
nand UO_318 (O_318,N_14091,N_14119);
nand UO_319 (O_319,N_14489,N_14887);
nor UO_320 (O_320,N_14726,N_14013);
nand UO_321 (O_321,N_14285,N_14760);
nor UO_322 (O_322,N_14708,N_14176);
xor UO_323 (O_323,N_14457,N_14673);
nor UO_324 (O_324,N_14766,N_14071);
and UO_325 (O_325,N_14073,N_14510);
nand UO_326 (O_326,N_14014,N_14496);
nand UO_327 (O_327,N_14420,N_14869);
nand UO_328 (O_328,N_14527,N_14539);
or UO_329 (O_329,N_14648,N_14957);
nand UO_330 (O_330,N_14210,N_14371);
and UO_331 (O_331,N_14191,N_14702);
xnor UO_332 (O_332,N_14244,N_14952);
and UO_333 (O_333,N_14843,N_14007);
nand UO_334 (O_334,N_14193,N_14079);
nand UO_335 (O_335,N_14962,N_14801);
nand UO_336 (O_336,N_14313,N_14427);
xnor UO_337 (O_337,N_14890,N_14744);
and UO_338 (O_338,N_14116,N_14133);
or UO_339 (O_339,N_14793,N_14897);
xnor UO_340 (O_340,N_14681,N_14250);
or UO_341 (O_341,N_14751,N_14565);
or UO_342 (O_342,N_14860,N_14185);
xnor UO_343 (O_343,N_14423,N_14426);
nand UO_344 (O_344,N_14323,N_14519);
nor UO_345 (O_345,N_14732,N_14657);
nor UO_346 (O_346,N_14987,N_14362);
and UO_347 (O_347,N_14885,N_14301);
and UO_348 (O_348,N_14892,N_14910);
nand UO_349 (O_349,N_14434,N_14741);
nor UO_350 (O_350,N_14904,N_14685);
or UO_351 (O_351,N_14199,N_14998);
and UO_352 (O_352,N_14569,N_14776);
nor UO_353 (O_353,N_14296,N_14026);
nand UO_354 (O_354,N_14198,N_14047);
nor UO_355 (O_355,N_14960,N_14719);
xor UO_356 (O_356,N_14325,N_14340);
xor UO_357 (O_357,N_14740,N_14267);
or UO_358 (O_358,N_14786,N_14197);
xnor UO_359 (O_359,N_14145,N_14995);
or UO_360 (O_360,N_14218,N_14488);
nand UO_361 (O_361,N_14406,N_14366);
nor UO_362 (O_362,N_14179,N_14636);
and UO_363 (O_363,N_14054,N_14507);
nand UO_364 (O_364,N_14466,N_14963);
xor UO_365 (O_365,N_14755,N_14906);
nand UO_366 (O_366,N_14707,N_14031);
and UO_367 (O_367,N_14241,N_14710);
nand UO_368 (O_368,N_14894,N_14600);
nor UO_369 (O_369,N_14008,N_14493);
nor UO_370 (O_370,N_14806,N_14670);
or UO_371 (O_371,N_14749,N_14970);
or UO_372 (O_372,N_14530,N_14649);
nand UO_373 (O_373,N_14090,N_14408);
and UO_374 (O_374,N_14956,N_14446);
nand UO_375 (O_375,N_14444,N_14717);
xnor UO_376 (O_376,N_14516,N_14617);
or UO_377 (O_377,N_14280,N_14540);
nand UO_378 (O_378,N_14893,N_14312);
nand UO_379 (O_379,N_14117,N_14040);
xnor UO_380 (O_380,N_14872,N_14661);
nand UO_381 (O_381,N_14818,N_14650);
nand UO_382 (O_382,N_14690,N_14287);
nor UO_383 (O_383,N_14972,N_14953);
nor UO_384 (O_384,N_14548,N_14795);
and UO_385 (O_385,N_14981,N_14397);
nand UO_386 (O_386,N_14759,N_14723);
xor UO_387 (O_387,N_14223,N_14544);
nor UO_388 (O_388,N_14293,N_14610);
and UO_389 (O_389,N_14938,N_14458);
nor UO_390 (O_390,N_14535,N_14392);
or UO_391 (O_391,N_14093,N_14824);
nand UO_392 (O_392,N_14166,N_14713);
nor UO_393 (O_393,N_14204,N_14300);
nor UO_394 (O_394,N_14317,N_14633);
or UO_395 (O_395,N_14445,N_14639);
or UO_396 (O_396,N_14104,N_14993);
nor UO_397 (O_397,N_14653,N_14417);
or UO_398 (O_398,N_14784,N_14486);
and UO_399 (O_399,N_14965,N_14452);
or UO_400 (O_400,N_14954,N_14677);
and UO_401 (O_401,N_14234,N_14405);
and UO_402 (O_402,N_14990,N_14238);
xor UO_403 (O_403,N_14733,N_14935);
and UO_404 (O_404,N_14118,N_14122);
and UO_405 (O_405,N_14257,N_14390);
nor UO_406 (O_406,N_14605,N_14414);
nor UO_407 (O_407,N_14126,N_14889);
nand UO_408 (O_408,N_14358,N_14021);
nor UO_409 (O_409,N_14721,N_14557);
xnor UO_410 (O_410,N_14222,N_14232);
or UO_411 (O_411,N_14978,N_14055);
and UO_412 (O_412,N_14048,N_14798);
nor UO_413 (O_413,N_14308,N_14811);
or UO_414 (O_414,N_14916,N_14915);
nor UO_415 (O_415,N_14808,N_14168);
nor UO_416 (O_416,N_14692,N_14192);
nor UO_417 (O_417,N_14777,N_14886);
nor UO_418 (O_418,N_14342,N_14011);
nand UO_419 (O_419,N_14006,N_14178);
nand UO_420 (O_420,N_14765,N_14888);
nand UO_421 (O_421,N_14714,N_14272);
nand UO_422 (O_422,N_14407,N_14081);
and UO_423 (O_423,N_14966,N_14545);
and UO_424 (O_424,N_14038,N_14331);
nor UO_425 (O_425,N_14746,N_14752);
and UO_426 (O_426,N_14775,N_14035);
or UO_427 (O_427,N_14212,N_14814);
nor UO_428 (O_428,N_14646,N_14835);
or UO_429 (O_429,N_14838,N_14028);
nor UO_430 (O_430,N_14867,N_14004);
nor UO_431 (O_431,N_14899,N_14132);
nor UO_432 (O_432,N_14559,N_14352);
nor UO_433 (O_433,N_14110,N_14528);
nand UO_434 (O_434,N_14490,N_14626);
xor UO_435 (O_435,N_14590,N_14248);
nand UO_436 (O_436,N_14575,N_14851);
nand UO_437 (O_437,N_14382,N_14353);
and UO_438 (O_438,N_14846,N_14439);
nand UO_439 (O_439,N_14097,N_14355);
nand UO_440 (O_440,N_14552,N_14919);
nand UO_441 (O_441,N_14156,N_14333);
nor UO_442 (O_442,N_14984,N_14580);
or UO_443 (O_443,N_14328,N_14027);
nor UO_444 (O_444,N_14859,N_14669);
nor UO_445 (O_445,N_14772,N_14470);
or UO_446 (O_446,N_14898,N_14190);
nor UO_447 (O_447,N_14059,N_14505);
xnor UO_448 (O_448,N_14111,N_14951);
and UO_449 (O_449,N_14724,N_14497);
nor UO_450 (O_450,N_14154,N_14265);
nand UO_451 (O_451,N_14182,N_14694);
or UO_452 (O_452,N_14622,N_14847);
xnor UO_453 (O_453,N_14345,N_14841);
nand UO_454 (O_454,N_14839,N_14820);
and UO_455 (O_455,N_14326,N_14367);
or UO_456 (O_456,N_14224,N_14644);
or UO_457 (O_457,N_14115,N_14112);
nor UO_458 (O_458,N_14597,N_14139);
xnor UO_459 (O_459,N_14534,N_14056);
xor UO_460 (O_460,N_14668,N_14762);
nor UO_461 (O_461,N_14750,N_14365);
or UO_462 (O_462,N_14495,N_14930);
nand UO_463 (O_463,N_14383,N_14842);
and UO_464 (O_464,N_14980,N_14868);
xor UO_465 (O_465,N_14531,N_14155);
nor UO_466 (O_466,N_14878,N_14269);
xnor UO_467 (O_467,N_14069,N_14288);
or UO_468 (O_468,N_14206,N_14329);
and UO_469 (O_469,N_14482,N_14959);
nand UO_470 (O_470,N_14175,N_14619);
nor UO_471 (O_471,N_14402,N_14704);
or UO_472 (O_472,N_14948,N_14621);
nand UO_473 (O_473,N_14428,N_14440);
nor UO_474 (O_474,N_14643,N_14874);
nand UO_475 (O_475,N_14881,N_14815);
nor UO_476 (O_476,N_14088,N_14526);
or UO_477 (O_477,N_14896,N_14070);
nand UO_478 (O_478,N_14092,N_14738);
and UO_479 (O_479,N_14195,N_14572);
or UO_480 (O_480,N_14217,N_14934);
or UO_481 (O_481,N_14082,N_14171);
or UO_482 (O_482,N_14787,N_14761);
nor UO_483 (O_483,N_14354,N_14532);
nor UO_484 (O_484,N_14475,N_14658);
nor UO_485 (O_485,N_14036,N_14576);
or UO_486 (O_486,N_14549,N_14350);
nor UO_487 (O_487,N_14042,N_14282);
and UO_488 (O_488,N_14812,N_14720);
nand UO_489 (O_489,N_14418,N_14002);
and UO_490 (O_490,N_14696,N_14142);
nand UO_491 (O_491,N_14334,N_14920);
nand UO_492 (O_492,N_14243,N_14974);
or UO_493 (O_493,N_14891,N_14901);
xor UO_494 (O_494,N_14306,N_14711);
nand UO_495 (O_495,N_14849,N_14631);
xnor UO_496 (O_496,N_14208,N_14615);
nor UO_497 (O_497,N_14105,N_14589);
and UO_498 (O_498,N_14158,N_14611);
and UO_499 (O_499,N_14687,N_14196);
and UO_500 (O_500,N_14291,N_14871);
nand UO_501 (O_501,N_14682,N_14254);
or UO_502 (O_502,N_14187,N_14845);
and UO_503 (O_503,N_14407,N_14892);
or UO_504 (O_504,N_14572,N_14092);
and UO_505 (O_505,N_14004,N_14632);
or UO_506 (O_506,N_14431,N_14850);
nor UO_507 (O_507,N_14136,N_14789);
and UO_508 (O_508,N_14372,N_14643);
and UO_509 (O_509,N_14309,N_14063);
or UO_510 (O_510,N_14533,N_14480);
nor UO_511 (O_511,N_14530,N_14515);
nand UO_512 (O_512,N_14830,N_14768);
or UO_513 (O_513,N_14927,N_14191);
and UO_514 (O_514,N_14905,N_14766);
and UO_515 (O_515,N_14750,N_14896);
or UO_516 (O_516,N_14934,N_14057);
and UO_517 (O_517,N_14002,N_14087);
nand UO_518 (O_518,N_14906,N_14492);
nor UO_519 (O_519,N_14699,N_14294);
or UO_520 (O_520,N_14758,N_14948);
nand UO_521 (O_521,N_14927,N_14793);
or UO_522 (O_522,N_14166,N_14016);
and UO_523 (O_523,N_14686,N_14822);
or UO_524 (O_524,N_14108,N_14389);
or UO_525 (O_525,N_14303,N_14857);
nand UO_526 (O_526,N_14338,N_14925);
and UO_527 (O_527,N_14903,N_14033);
nand UO_528 (O_528,N_14872,N_14154);
or UO_529 (O_529,N_14748,N_14605);
xnor UO_530 (O_530,N_14901,N_14295);
nand UO_531 (O_531,N_14866,N_14448);
nand UO_532 (O_532,N_14723,N_14815);
and UO_533 (O_533,N_14324,N_14440);
nor UO_534 (O_534,N_14238,N_14605);
and UO_535 (O_535,N_14361,N_14872);
nand UO_536 (O_536,N_14707,N_14914);
or UO_537 (O_537,N_14921,N_14791);
and UO_538 (O_538,N_14331,N_14143);
nand UO_539 (O_539,N_14004,N_14935);
nand UO_540 (O_540,N_14635,N_14861);
or UO_541 (O_541,N_14641,N_14326);
and UO_542 (O_542,N_14773,N_14624);
nor UO_543 (O_543,N_14657,N_14351);
nor UO_544 (O_544,N_14537,N_14626);
or UO_545 (O_545,N_14589,N_14009);
xnor UO_546 (O_546,N_14615,N_14123);
or UO_547 (O_547,N_14453,N_14801);
nand UO_548 (O_548,N_14134,N_14940);
xnor UO_549 (O_549,N_14145,N_14376);
or UO_550 (O_550,N_14735,N_14753);
and UO_551 (O_551,N_14460,N_14897);
and UO_552 (O_552,N_14419,N_14665);
nand UO_553 (O_553,N_14874,N_14199);
or UO_554 (O_554,N_14165,N_14605);
or UO_555 (O_555,N_14790,N_14583);
and UO_556 (O_556,N_14116,N_14613);
and UO_557 (O_557,N_14255,N_14431);
nand UO_558 (O_558,N_14425,N_14054);
nor UO_559 (O_559,N_14888,N_14736);
or UO_560 (O_560,N_14795,N_14547);
xnor UO_561 (O_561,N_14682,N_14267);
xor UO_562 (O_562,N_14624,N_14293);
nor UO_563 (O_563,N_14160,N_14876);
and UO_564 (O_564,N_14611,N_14974);
and UO_565 (O_565,N_14580,N_14325);
nor UO_566 (O_566,N_14749,N_14808);
nor UO_567 (O_567,N_14330,N_14103);
or UO_568 (O_568,N_14492,N_14780);
or UO_569 (O_569,N_14863,N_14605);
or UO_570 (O_570,N_14146,N_14691);
xnor UO_571 (O_571,N_14091,N_14084);
and UO_572 (O_572,N_14682,N_14474);
nor UO_573 (O_573,N_14371,N_14946);
and UO_574 (O_574,N_14380,N_14395);
and UO_575 (O_575,N_14706,N_14515);
nand UO_576 (O_576,N_14623,N_14180);
nand UO_577 (O_577,N_14046,N_14904);
and UO_578 (O_578,N_14990,N_14709);
and UO_579 (O_579,N_14467,N_14383);
and UO_580 (O_580,N_14657,N_14745);
xor UO_581 (O_581,N_14367,N_14841);
nand UO_582 (O_582,N_14874,N_14500);
nand UO_583 (O_583,N_14160,N_14627);
nand UO_584 (O_584,N_14528,N_14669);
xnor UO_585 (O_585,N_14465,N_14952);
or UO_586 (O_586,N_14607,N_14343);
or UO_587 (O_587,N_14850,N_14666);
nor UO_588 (O_588,N_14272,N_14859);
nor UO_589 (O_589,N_14427,N_14815);
xor UO_590 (O_590,N_14520,N_14719);
nand UO_591 (O_591,N_14000,N_14381);
nand UO_592 (O_592,N_14128,N_14660);
xor UO_593 (O_593,N_14997,N_14356);
nor UO_594 (O_594,N_14860,N_14341);
nand UO_595 (O_595,N_14158,N_14770);
nor UO_596 (O_596,N_14895,N_14778);
nand UO_597 (O_597,N_14601,N_14465);
or UO_598 (O_598,N_14304,N_14227);
nor UO_599 (O_599,N_14071,N_14756);
nand UO_600 (O_600,N_14306,N_14912);
nor UO_601 (O_601,N_14477,N_14847);
nand UO_602 (O_602,N_14749,N_14246);
or UO_603 (O_603,N_14578,N_14103);
or UO_604 (O_604,N_14764,N_14852);
nand UO_605 (O_605,N_14585,N_14710);
nor UO_606 (O_606,N_14263,N_14645);
nand UO_607 (O_607,N_14635,N_14426);
nor UO_608 (O_608,N_14280,N_14859);
nor UO_609 (O_609,N_14149,N_14022);
nor UO_610 (O_610,N_14229,N_14864);
and UO_611 (O_611,N_14376,N_14419);
and UO_612 (O_612,N_14561,N_14906);
and UO_613 (O_613,N_14400,N_14221);
nor UO_614 (O_614,N_14097,N_14705);
nor UO_615 (O_615,N_14680,N_14305);
nand UO_616 (O_616,N_14388,N_14296);
nor UO_617 (O_617,N_14660,N_14657);
nor UO_618 (O_618,N_14293,N_14548);
and UO_619 (O_619,N_14484,N_14290);
or UO_620 (O_620,N_14256,N_14101);
or UO_621 (O_621,N_14658,N_14306);
and UO_622 (O_622,N_14014,N_14133);
or UO_623 (O_623,N_14193,N_14890);
and UO_624 (O_624,N_14967,N_14361);
nand UO_625 (O_625,N_14670,N_14553);
or UO_626 (O_626,N_14617,N_14445);
and UO_627 (O_627,N_14527,N_14774);
and UO_628 (O_628,N_14457,N_14487);
nand UO_629 (O_629,N_14190,N_14348);
nor UO_630 (O_630,N_14283,N_14365);
or UO_631 (O_631,N_14477,N_14589);
xnor UO_632 (O_632,N_14700,N_14549);
nor UO_633 (O_633,N_14377,N_14842);
and UO_634 (O_634,N_14559,N_14857);
or UO_635 (O_635,N_14093,N_14452);
nand UO_636 (O_636,N_14515,N_14631);
and UO_637 (O_637,N_14010,N_14277);
nor UO_638 (O_638,N_14982,N_14346);
and UO_639 (O_639,N_14935,N_14401);
nand UO_640 (O_640,N_14788,N_14686);
nor UO_641 (O_641,N_14305,N_14126);
nor UO_642 (O_642,N_14208,N_14796);
nand UO_643 (O_643,N_14888,N_14605);
or UO_644 (O_644,N_14527,N_14773);
nor UO_645 (O_645,N_14371,N_14150);
or UO_646 (O_646,N_14148,N_14555);
and UO_647 (O_647,N_14727,N_14398);
and UO_648 (O_648,N_14592,N_14816);
xor UO_649 (O_649,N_14860,N_14360);
nor UO_650 (O_650,N_14039,N_14087);
nor UO_651 (O_651,N_14972,N_14735);
nor UO_652 (O_652,N_14504,N_14746);
and UO_653 (O_653,N_14096,N_14677);
nand UO_654 (O_654,N_14697,N_14274);
and UO_655 (O_655,N_14580,N_14112);
nor UO_656 (O_656,N_14956,N_14197);
and UO_657 (O_657,N_14257,N_14242);
xnor UO_658 (O_658,N_14821,N_14548);
nand UO_659 (O_659,N_14496,N_14137);
or UO_660 (O_660,N_14490,N_14374);
nand UO_661 (O_661,N_14358,N_14463);
or UO_662 (O_662,N_14450,N_14697);
nand UO_663 (O_663,N_14940,N_14102);
nand UO_664 (O_664,N_14560,N_14282);
and UO_665 (O_665,N_14199,N_14506);
or UO_666 (O_666,N_14602,N_14191);
or UO_667 (O_667,N_14383,N_14579);
and UO_668 (O_668,N_14132,N_14028);
nor UO_669 (O_669,N_14723,N_14674);
nor UO_670 (O_670,N_14262,N_14672);
nand UO_671 (O_671,N_14382,N_14076);
and UO_672 (O_672,N_14436,N_14477);
and UO_673 (O_673,N_14721,N_14391);
or UO_674 (O_674,N_14150,N_14798);
and UO_675 (O_675,N_14199,N_14849);
xnor UO_676 (O_676,N_14385,N_14729);
nor UO_677 (O_677,N_14834,N_14899);
xnor UO_678 (O_678,N_14536,N_14340);
nand UO_679 (O_679,N_14482,N_14104);
nand UO_680 (O_680,N_14520,N_14649);
nor UO_681 (O_681,N_14792,N_14847);
nor UO_682 (O_682,N_14137,N_14657);
and UO_683 (O_683,N_14493,N_14380);
or UO_684 (O_684,N_14423,N_14547);
nor UO_685 (O_685,N_14372,N_14778);
nand UO_686 (O_686,N_14964,N_14820);
nand UO_687 (O_687,N_14962,N_14109);
nor UO_688 (O_688,N_14552,N_14039);
or UO_689 (O_689,N_14190,N_14822);
nand UO_690 (O_690,N_14543,N_14934);
or UO_691 (O_691,N_14954,N_14774);
nand UO_692 (O_692,N_14830,N_14248);
nand UO_693 (O_693,N_14458,N_14088);
and UO_694 (O_694,N_14344,N_14696);
nor UO_695 (O_695,N_14847,N_14497);
and UO_696 (O_696,N_14494,N_14825);
or UO_697 (O_697,N_14311,N_14360);
nand UO_698 (O_698,N_14623,N_14961);
nor UO_699 (O_699,N_14172,N_14074);
or UO_700 (O_700,N_14480,N_14527);
and UO_701 (O_701,N_14537,N_14906);
or UO_702 (O_702,N_14697,N_14209);
and UO_703 (O_703,N_14967,N_14961);
or UO_704 (O_704,N_14567,N_14508);
and UO_705 (O_705,N_14323,N_14165);
xor UO_706 (O_706,N_14850,N_14891);
nand UO_707 (O_707,N_14865,N_14175);
nor UO_708 (O_708,N_14403,N_14357);
or UO_709 (O_709,N_14497,N_14305);
and UO_710 (O_710,N_14518,N_14446);
and UO_711 (O_711,N_14314,N_14181);
nand UO_712 (O_712,N_14906,N_14982);
nor UO_713 (O_713,N_14686,N_14102);
nand UO_714 (O_714,N_14138,N_14922);
and UO_715 (O_715,N_14648,N_14398);
and UO_716 (O_716,N_14891,N_14647);
or UO_717 (O_717,N_14850,N_14634);
and UO_718 (O_718,N_14627,N_14355);
xnor UO_719 (O_719,N_14945,N_14241);
or UO_720 (O_720,N_14110,N_14136);
or UO_721 (O_721,N_14367,N_14001);
and UO_722 (O_722,N_14415,N_14971);
and UO_723 (O_723,N_14131,N_14603);
or UO_724 (O_724,N_14111,N_14875);
nand UO_725 (O_725,N_14879,N_14275);
or UO_726 (O_726,N_14789,N_14766);
and UO_727 (O_727,N_14133,N_14887);
nor UO_728 (O_728,N_14960,N_14565);
nor UO_729 (O_729,N_14879,N_14775);
and UO_730 (O_730,N_14851,N_14017);
and UO_731 (O_731,N_14739,N_14708);
nor UO_732 (O_732,N_14525,N_14254);
xnor UO_733 (O_733,N_14711,N_14133);
and UO_734 (O_734,N_14103,N_14548);
nand UO_735 (O_735,N_14404,N_14566);
or UO_736 (O_736,N_14552,N_14816);
xnor UO_737 (O_737,N_14437,N_14471);
nor UO_738 (O_738,N_14581,N_14635);
nand UO_739 (O_739,N_14340,N_14472);
nor UO_740 (O_740,N_14997,N_14354);
or UO_741 (O_741,N_14030,N_14773);
and UO_742 (O_742,N_14113,N_14698);
nand UO_743 (O_743,N_14354,N_14138);
or UO_744 (O_744,N_14094,N_14782);
or UO_745 (O_745,N_14930,N_14426);
and UO_746 (O_746,N_14778,N_14436);
nand UO_747 (O_747,N_14086,N_14808);
or UO_748 (O_748,N_14046,N_14179);
and UO_749 (O_749,N_14525,N_14711);
and UO_750 (O_750,N_14226,N_14179);
xor UO_751 (O_751,N_14559,N_14396);
or UO_752 (O_752,N_14292,N_14342);
xnor UO_753 (O_753,N_14136,N_14287);
nor UO_754 (O_754,N_14893,N_14220);
xor UO_755 (O_755,N_14548,N_14386);
and UO_756 (O_756,N_14567,N_14410);
nand UO_757 (O_757,N_14506,N_14848);
nor UO_758 (O_758,N_14013,N_14660);
or UO_759 (O_759,N_14483,N_14939);
and UO_760 (O_760,N_14060,N_14512);
nand UO_761 (O_761,N_14853,N_14772);
or UO_762 (O_762,N_14405,N_14978);
and UO_763 (O_763,N_14827,N_14851);
nor UO_764 (O_764,N_14378,N_14301);
and UO_765 (O_765,N_14564,N_14809);
nor UO_766 (O_766,N_14834,N_14137);
nor UO_767 (O_767,N_14338,N_14129);
xor UO_768 (O_768,N_14460,N_14949);
or UO_769 (O_769,N_14151,N_14869);
or UO_770 (O_770,N_14883,N_14500);
nand UO_771 (O_771,N_14154,N_14400);
nand UO_772 (O_772,N_14627,N_14827);
nor UO_773 (O_773,N_14008,N_14025);
nand UO_774 (O_774,N_14888,N_14509);
xnor UO_775 (O_775,N_14855,N_14038);
or UO_776 (O_776,N_14304,N_14786);
nor UO_777 (O_777,N_14247,N_14451);
nand UO_778 (O_778,N_14330,N_14879);
nand UO_779 (O_779,N_14509,N_14512);
and UO_780 (O_780,N_14264,N_14985);
and UO_781 (O_781,N_14398,N_14350);
and UO_782 (O_782,N_14934,N_14688);
or UO_783 (O_783,N_14429,N_14464);
and UO_784 (O_784,N_14167,N_14357);
nor UO_785 (O_785,N_14525,N_14003);
or UO_786 (O_786,N_14772,N_14510);
or UO_787 (O_787,N_14668,N_14480);
nor UO_788 (O_788,N_14866,N_14655);
nand UO_789 (O_789,N_14531,N_14221);
or UO_790 (O_790,N_14760,N_14442);
or UO_791 (O_791,N_14116,N_14429);
nand UO_792 (O_792,N_14357,N_14224);
nand UO_793 (O_793,N_14605,N_14398);
nor UO_794 (O_794,N_14751,N_14657);
or UO_795 (O_795,N_14567,N_14660);
and UO_796 (O_796,N_14109,N_14654);
xnor UO_797 (O_797,N_14844,N_14367);
xnor UO_798 (O_798,N_14961,N_14199);
and UO_799 (O_799,N_14611,N_14536);
nand UO_800 (O_800,N_14518,N_14964);
and UO_801 (O_801,N_14791,N_14374);
nor UO_802 (O_802,N_14168,N_14179);
or UO_803 (O_803,N_14014,N_14570);
nand UO_804 (O_804,N_14500,N_14663);
nand UO_805 (O_805,N_14849,N_14541);
xor UO_806 (O_806,N_14152,N_14931);
and UO_807 (O_807,N_14531,N_14797);
nor UO_808 (O_808,N_14786,N_14939);
and UO_809 (O_809,N_14666,N_14842);
xor UO_810 (O_810,N_14204,N_14429);
nand UO_811 (O_811,N_14481,N_14333);
nand UO_812 (O_812,N_14082,N_14102);
nand UO_813 (O_813,N_14534,N_14375);
nand UO_814 (O_814,N_14358,N_14329);
nand UO_815 (O_815,N_14411,N_14794);
and UO_816 (O_816,N_14695,N_14848);
or UO_817 (O_817,N_14822,N_14203);
and UO_818 (O_818,N_14510,N_14050);
xnor UO_819 (O_819,N_14239,N_14245);
or UO_820 (O_820,N_14371,N_14362);
nor UO_821 (O_821,N_14163,N_14731);
nor UO_822 (O_822,N_14834,N_14408);
xnor UO_823 (O_823,N_14160,N_14678);
and UO_824 (O_824,N_14991,N_14010);
xor UO_825 (O_825,N_14847,N_14285);
xnor UO_826 (O_826,N_14169,N_14588);
or UO_827 (O_827,N_14780,N_14879);
and UO_828 (O_828,N_14895,N_14674);
or UO_829 (O_829,N_14115,N_14949);
nand UO_830 (O_830,N_14539,N_14833);
and UO_831 (O_831,N_14622,N_14629);
or UO_832 (O_832,N_14166,N_14841);
nor UO_833 (O_833,N_14885,N_14166);
or UO_834 (O_834,N_14831,N_14900);
or UO_835 (O_835,N_14959,N_14086);
nor UO_836 (O_836,N_14038,N_14492);
nor UO_837 (O_837,N_14401,N_14315);
and UO_838 (O_838,N_14495,N_14072);
nor UO_839 (O_839,N_14297,N_14861);
xor UO_840 (O_840,N_14232,N_14108);
nand UO_841 (O_841,N_14371,N_14836);
nor UO_842 (O_842,N_14528,N_14729);
nor UO_843 (O_843,N_14947,N_14044);
nor UO_844 (O_844,N_14577,N_14748);
nand UO_845 (O_845,N_14933,N_14571);
nand UO_846 (O_846,N_14136,N_14285);
and UO_847 (O_847,N_14904,N_14896);
and UO_848 (O_848,N_14391,N_14574);
nor UO_849 (O_849,N_14391,N_14872);
nand UO_850 (O_850,N_14668,N_14942);
or UO_851 (O_851,N_14354,N_14541);
or UO_852 (O_852,N_14416,N_14749);
or UO_853 (O_853,N_14843,N_14615);
or UO_854 (O_854,N_14474,N_14127);
and UO_855 (O_855,N_14968,N_14056);
nand UO_856 (O_856,N_14844,N_14068);
nand UO_857 (O_857,N_14884,N_14165);
nand UO_858 (O_858,N_14871,N_14638);
and UO_859 (O_859,N_14958,N_14707);
nor UO_860 (O_860,N_14776,N_14945);
xor UO_861 (O_861,N_14690,N_14063);
or UO_862 (O_862,N_14472,N_14237);
or UO_863 (O_863,N_14304,N_14355);
nand UO_864 (O_864,N_14557,N_14277);
nand UO_865 (O_865,N_14226,N_14216);
nand UO_866 (O_866,N_14811,N_14489);
xnor UO_867 (O_867,N_14835,N_14955);
and UO_868 (O_868,N_14280,N_14238);
nand UO_869 (O_869,N_14827,N_14184);
nor UO_870 (O_870,N_14436,N_14096);
or UO_871 (O_871,N_14139,N_14274);
xor UO_872 (O_872,N_14487,N_14281);
nor UO_873 (O_873,N_14108,N_14625);
and UO_874 (O_874,N_14903,N_14036);
nor UO_875 (O_875,N_14066,N_14710);
nand UO_876 (O_876,N_14896,N_14305);
nand UO_877 (O_877,N_14786,N_14144);
nor UO_878 (O_878,N_14601,N_14060);
xor UO_879 (O_879,N_14796,N_14106);
or UO_880 (O_880,N_14109,N_14498);
xor UO_881 (O_881,N_14915,N_14121);
nand UO_882 (O_882,N_14377,N_14236);
nand UO_883 (O_883,N_14031,N_14056);
nand UO_884 (O_884,N_14405,N_14638);
nor UO_885 (O_885,N_14770,N_14617);
and UO_886 (O_886,N_14265,N_14454);
nand UO_887 (O_887,N_14434,N_14150);
and UO_888 (O_888,N_14017,N_14567);
nand UO_889 (O_889,N_14561,N_14268);
or UO_890 (O_890,N_14554,N_14341);
nand UO_891 (O_891,N_14818,N_14106);
nand UO_892 (O_892,N_14214,N_14334);
xnor UO_893 (O_893,N_14283,N_14529);
or UO_894 (O_894,N_14809,N_14163);
nand UO_895 (O_895,N_14598,N_14602);
nor UO_896 (O_896,N_14117,N_14932);
nor UO_897 (O_897,N_14259,N_14079);
and UO_898 (O_898,N_14031,N_14152);
nor UO_899 (O_899,N_14723,N_14315);
and UO_900 (O_900,N_14433,N_14191);
or UO_901 (O_901,N_14022,N_14226);
nor UO_902 (O_902,N_14124,N_14982);
nor UO_903 (O_903,N_14673,N_14377);
nand UO_904 (O_904,N_14386,N_14704);
and UO_905 (O_905,N_14503,N_14757);
xor UO_906 (O_906,N_14383,N_14286);
and UO_907 (O_907,N_14784,N_14764);
nand UO_908 (O_908,N_14694,N_14210);
nor UO_909 (O_909,N_14611,N_14947);
nor UO_910 (O_910,N_14073,N_14798);
nor UO_911 (O_911,N_14516,N_14327);
nor UO_912 (O_912,N_14250,N_14756);
or UO_913 (O_913,N_14341,N_14084);
or UO_914 (O_914,N_14247,N_14510);
or UO_915 (O_915,N_14630,N_14788);
or UO_916 (O_916,N_14338,N_14449);
nand UO_917 (O_917,N_14321,N_14929);
xnor UO_918 (O_918,N_14535,N_14195);
and UO_919 (O_919,N_14447,N_14544);
or UO_920 (O_920,N_14274,N_14082);
nand UO_921 (O_921,N_14639,N_14265);
or UO_922 (O_922,N_14521,N_14539);
or UO_923 (O_923,N_14682,N_14473);
or UO_924 (O_924,N_14344,N_14074);
and UO_925 (O_925,N_14235,N_14619);
nand UO_926 (O_926,N_14539,N_14337);
or UO_927 (O_927,N_14332,N_14196);
or UO_928 (O_928,N_14878,N_14284);
xnor UO_929 (O_929,N_14123,N_14929);
nand UO_930 (O_930,N_14197,N_14798);
and UO_931 (O_931,N_14326,N_14339);
or UO_932 (O_932,N_14858,N_14969);
and UO_933 (O_933,N_14655,N_14189);
or UO_934 (O_934,N_14720,N_14223);
nor UO_935 (O_935,N_14341,N_14520);
xor UO_936 (O_936,N_14027,N_14870);
or UO_937 (O_937,N_14071,N_14280);
xnor UO_938 (O_938,N_14410,N_14962);
or UO_939 (O_939,N_14127,N_14131);
nor UO_940 (O_940,N_14039,N_14881);
nor UO_941 (O_941,N_14278,N_14966);
or UO_942 (O_942,N_14456,N_14850);
or UO_943 (O_943,N_14377,N_14883);
nand UO_944 (O_944,N_14127,N_14863);
or UO_945 (O_945,N_14175,N_14575);
xor UO_946 (O_946,N_14182,N_14686);
nor UO_947 (O_947,N_14706,N_14676);
or UO_948 (O_948,N_14755,N_14457);
nor UO_949 (O_949,N_14588,N_14148);
or UO_950 (O_950,N_14411,N_14101);
nand UO_951 (O_951,N_14707,N_14141);
or UO_952 (O_952,N_14214,N_14862);
nor UO_953 (O_953,N_14195,N_14461);
xor UO_954 (O_954,N_14691,N_14553);
nand UO_955 (O_955,N_14584,N_14343);
nand UO_956 (O_956,N_14609,N_14158);
and UO_957 (O_957,N_14690,N_14222);
nor UO_958 (O_958,N_14929,N_14490);
and UO_959 (O_959,N_14346,N_14890);
nor UO_960 (O_960,N_14329,N_14018);
nor UO_961 (O_961,N_14417,N_14755);
nand UO_962 (O_962,N_14660,N_14640);
and UO_963 (O_963,N_14777,N_14212);
nor UO_964 (O_964,N_14295,N_14167);
xor UO_965 (O_965,N_14757,N_14580);
nor UO_966 (O_966,N_14479,N_14738);
or UO_967 (O_967,N_14383,N_14313);
and UO_968 (O_968,N_14475,N_14071);
and UO_969 (O_969,N_14845,N_14765);
nor UO_970 (O_970,N_14112,N_14988);
nand UO_971 (O_971,N_14841,N_14872);
xor UO_972 (O_972,N_14708,N_14951);
and UO_973 (O_973,N_14457,N_14015);
xor UO_974 (O_974,N_14832,N_14160);
or UO_975 (O_975,N_14646,N_14195);
or UO_976 (O_976,N_14573,N_14125);
or UO_977 (O_977,N_14212,N_14813);
nor UO_978 (O_978,N_14891,N_14028);
nor UO_979 (O_979,N_14040,N_14921);
nand UO_980 (O_980,N_14489,N_14171);
and UO_981 (O_981,N_14931,N_14409);
nor UO_982 (O_982,N_14586,N_14271);
nor UO_983 (O_983,N_14227,N_14731);
nor UO_984 (O_984,N_14785,N_14472);
and UO_985 (O_985,N_14334,N_14137);
nor UO_986 (O_986,N_14496,N_14691);
nand UO_987 (O_987,N_14424,N_14271);
nand UO_988 (O_988,N_14131,N_14072);
nand UO_989 (O_989,N_14923,N_14764);
or UO_990 (O_990,N_14332,N_14452);
nand UO_991 (O_991,N_14778,N_14716);
and UO_992 (O_992,N_14449,N_14879);
nand UO_993 (O_993,N_14380,N_14663);
or UO_994 (O_994,N_14537,N_14127);
nor UO_995 (O_995,N_14104,N_14633);
nor UO_996 (O_996,N_14524,N_14009);
and UO_997 (O_997,N_14187,N_14662);
and UO_998 (O_998,N_14252,N_14630);
and UO_999 (O_999,N_14340,N_14517);
nor UO_1000 (O_1000,N_14922,N_14879);
xnor UO_1001 (O_1001,N_14699,N_14107);
nand UO_1002 (O_1002,N_14141,N_14389);
nand UO_1003 (O_1003,N_14475,N_14558);
or UO_1004 (O_1004,N_14932,N_14010);
or UO_1005 (O_1005,N_14952,N_14293);
nor UO_1006 (O_1006,N_14288,N_14213);
xnor UO_1007 (O_1007,N_14248,N_14806);
nor UO_1008 (O_1008,N_14661,N_14300);
and UO_1009 (O_1009,N_14319,N_14961);
and UO_1010 (O_1010,N_14222,N_14015);
or UO_1011 (O_1011,N_14380,N_14675);
nand UO_1012 (O_1012,N_14388,N_14282);
and UO_1013 (O_1013,N_14520,N_14709);
or UO_1014 (O_1014,N_14864,N_14014);
nand UO_1015 (O_1015,N_14477,N_14388);
or UO_1016 (O_1016,N_14171,N_14275);
and UO_1017 (O_1017,N_14307,N_14186);
nor UO_1018 (O_1018,N_14450,N_14617);
or UO_1019 (O_1019,N_14323,N_14963);
or UO_1020 (O_1020,N_14585,N_14162);
and UO_1021 (O_1021,N_14719,N_14241);
nor UO_1022 (O_1022,N_14079,N_14206);
and UO_1023 (O_1023,N_14318,N_14271);
or UO_1024 (O_1024,N_14286,N_14639);
nor UO_1025 (O_1025,N_14445,N_14222);
or UO_1026 (O_1026,N_14902,N_14398);
nor UO_1027 (O_1027,N_14329,N_14084);
or UO_1028 (O_1028,N_14170,N_14227);
nor UO_1029 (O_1029,N_14272,N_14321);
or UO_1030 (O_1030,N_14952,N_14030);
or UO_1031 (O_1031,N_14184,N_14460);
nand UO_1032 (O_1032,N_14959,N_14600);
or UO_1033 (O_1033,N_14578,N_14732);
nor UO_1034 (O_1034,N_14476,N_14297);
and UO_1035 (O_1035,N_14066,N_14361);
and UO_1036 (O_1036,N_14799,N_14886);
nor UO_1037 (O_1037,N_14621,N_14310);
nor UO_1038 (O_1038,N_14254,N_14336);
or UO_1039 (O_1039,N_14617,N_14937);
nand UO_1040 (O_1040,N_14390,N_14309);
nand UO_1041 (O_1041,N_14449,N_14770);
or UO_1042 (O_1042,N_14397,N_14181);
and UO_1043 (O_1043,N_14273,N_14046);
or UO_1044 (O_1044,N_14090,N_14202);
nor UO_1045 (O_1045,N_14981,N_14085);
nor UO_1046 (O_1046,N_14504,N_14252);
nor UO_1047 (O_1047,N_14632,N_14196);
or UO_1048 (O_1048,N_14000,N_14239);
or UO_1049 (O_1049,N_14258,N_14959);
and UO_1050 (O_1050,N_14969,N_14320);
or UO_1051 (O_1051,N_14140,N_14179);
or UO_1052 (O_1052,N_14545,N_14871);
and UO_1053 (O_1053,N_14127,N_14910);
nor UO_1054 (O_1054,N_14621,N_14569);
and UO_1055 (O_1055,N_14055,N_14334);
nor UO_1056 (O_1056,N_14323,N_14518);
nor UO_1057 (O_1057,N_14033,N_14964);
nor UO_1058 (O_1058,N_14652,N_14545);
or UO_1059 (O_1059,N_14600,N_14379);
and UO_1060 (O_1060,N_14135,N_14329);
xnor UO_1061 (O_1061,N_14599,N_14090);
xor UO_1062 (O_1062,N_14083,N_14288);
or UO_1063 (O_1063,N_14248,N_14142);
and UO_1064 (O_1064,N_14195,N_14701);
or UO_1065 (O_1065,N_14439,N_14689);
or UO_1066 (O_1066,N_14176,N_14074);
nor UO_1067 (O_1067,N_14432,N_14725);
nand UO_1068 (O_1068,N_14097,N_14431);
or UO_1069 (O_1069,N_14815,N_14639);
or UO_1070 (O_1070,N_14389,N_14366);
or UO_1071 (O_1071,N_14874,N_14312);
nor UO_1072 (O_1072,N_14339,N_14486);
nor UO_1073 (O_1073,N_14565,N_14522);
and UO_1074 (O_1074,N_14564,N_14689);
nand UO_1075 (O_1075,N_14222,N_14500);
nor UO_1076 (O_1076,N_14008,N_14099);
xnor UO_1077 (O_1077,N_14942,N_14339);
xor UO_1078 (O_1078,N_14682,N_14913);
and UO_1079 (O_1079,N_14218,N_14870);
nand UO_1080 (O_1080,N_14073,N_14809);
and UO_1081 (O_1081,N_14953,N_14328);
nand UO_1082 (O_1082,N_14326,N_14855);
nand UO_1083 (O_1083,N_14600,N_14988);
or UO_1084 (O_1084,N_14855,N_14987);
and UO_1085 (O_1085,N_14930,N_14176);
xor UO_1086 (O_1086,N_14823,N_14544);
and UO_1087 (O_1087,N_14261,N_14205);
nand UO_1088 (O_1088,N_14154,N_14838);
and UO_1089 (O_1089,N_14636,N_14820);
nand UO_1090 (O_1090,N_14971,N_14800);
or UO_1091 (O_1091,N_14167,N_14264);
nand UO_1092 (O_1092,N_14722,N_14906);
nor UO_1093 (O_1093,N_14586,N_14803);
nand UO_1094 (O_1094,N_14661,N_14761);
and UO_1095 (O_1095,N_14918,N_14158);
and UO_1096 (O_1096,N_14325,N_14303);
nor UO_1097 (O_1097,N_14805,N_14245);
or UO_1098 (O_1098,N_14547,N_14078);
xor UO_1099 (O_1099,N_14515,N_14406);
nor UO_1100 (O_1100,N_14331,N_14126);
nor UO_1101 (O_1101,N_14777,N_14309);
or UO_1102 (O_1102,N_14166,N_14596);
nor UO_1103 (O_1103,N_14051,N_14590);
and UO_1104 (O_1104,N_14216,N_14741);
and UO_1105 (O_1105,N_14559,N_14941);
nand UO_1106 (O_1106,N_14023,N_14296);
or UO_1107 (O_1107,N_14853,N_14926);
nand UO_1108 (O_1108,N_14157,N_14928);
nor UO_1109 (O_1109,N_14706,N_14374);
or UO_1110 (O_1110,N_14698,N_14562);
nand UO_1111 (O_1111,N_14243,N_14662);
nand UO_1112 (O_1112,N_14309,N_14339);
xnor UO_1113 (O_1113,N_14565,N_14072);
or UO_1114 (O_1114,N_14555,N_14428);
nand UO_1115 (O_1115,N_14821,N_14449);
nor UO_1116 (O_1116,N_14027,N_14408);
or UO_1117 (O_1117,N_14419,N_14554);
nor UO_1118 (O_1118,N_14212,N_14931);
nor UO_1119 (O_1119,N_14999,N_14241);
nand UO_1120 (O_1120,N_14080,N_14672);
and UO_1121 (O_1121,N_14040,N_14957);
or UO_1122 (O_1122,N_14377,N_14973);
nor UO_1123 (O_1123,N_14963,N_14369);
nand UO_1124 (O_1124,N_14192,N_14306);
nand UO_1125 (O_1125,N_14466,N_14693);
nor UO_1126 (O_1126,N_14315,N_14157);
or UO_1127 (O_1127,N_14736,N_14564);
nor UO_1128 (O_1128,N_14162,N_14606);
nand UO_1129 (O_1129,N_14199,N_14160);
nand UO_1130 (O_1130,N_14301,N_14268);
and UO_1131 (O_1131,N_14027,N_14472);
xor UO_1132 (O_1132,N_14306,N_14883);
or UO_1133 (O_1133,N_14106,N_14651);
nor UO_1134 (O_1134,N_14423,N_14372);
xor UO_1135 (O_1135,N_14604,N_14479);
nand UO_1136 (O_1136,N_14749,N_14333);
nand UO_1137 (O_1137,N_14570,N_14488);
or UO_1138 (O_1138,N_14917,N_14133);
or UO_1139 (O_1139,N_14751,N_14467);
and UO_1140 (O_1140,N_14540,N_14710);
or UO_1141 (O_1141,N_14643,N_14697);
xnor UO_1142 (O_1142,N_14622,N_14828);
or UO_1143 (O_1143,N_14667,N_14039);
nand UO_1144 (O_1144,N_14977,N_14144);
nor UO_1145 (O_1145,N_14401,N_14062);
nand UO_1146 (O_1146,N_14623,N_14711);
nor UO_1147 (O_1147,N_14197,N_14334);
nor UO_1148 (O_1148,N_14962,N_14692);
and UO_1149 (O_1149,N_14193,N_14113);
nor UO_1150 (O_1150,N_14170,N_14070);
and UO_1151 (O_1151,N_14981,N_14611);
or UO_1152 (O_1152,N_14866,N_14508);
nand UO_1153 (O_1153,N_14711,N_14157);
or UO_1154 (O_1154,N_14968,N_14969);
and UO_1155 (O_1155,N_14446,N_14540);
nand UO_1156 (O_1156,N_14587,N_14472);
or UO_1157 (O_1157,N_14195,N_14074);
nand UO_1158 (O_1158,N_14558,N_14878);
nand UO_1159 (O_1159,N_14715,N_14514);
nand UO_1160 (O_1160,N_14276,N_14499);
nand UO_1161 (O_1161,N_14089,N_14417);
and UO_1162 (O_1162,N_14220,N_14865);
nor UO_1163 (O_1163,N_14592,N_14657);
nand UO_1164 (O_1164,N_14052,N_14404);
nand UO_1165 (O_1165,N_14850,N_14214);
and UO_1166 (O_1166,N_14149,N_14787);
and UO_1167 (O_1167,N_14340,N_14947);
or UO_1168 (O_1168,N_14748,N_14559);
nor UO_1169 (O_1169,N_14356,N_14813);
nand UO_1170 (O_1170,N_14082,N_14255);
and UO_1171 (O_1171,N_14484,N_14316);
or UO_1172 (O_1172,N_14972,N_14095);
or UO_1173 (O_1173,N_14974,N_14819);
and UO_1174 (O_1174,N_14865,N_14856);
nand UO_1175 (O_1175,N_14839,N_14597);
nor UO_1176 (O_1176,N_14543,N_14816);
and UO_1177 (O_1177,N_14222,N_14253);
nand UO_1178 (O_1178,N_14049,N_14313);
nand UO_1179 (O_1179,N_14620,N_14373);
nand UO_1180 (O_1180,N_14047,N_14731);
or UO_1181 (O_1181,N_14479,N_14246);
nand UO_1182 (O_1182,N_14510,N_14928);
xor UO_1183 (O_1183,N_14061,N_14661);
or UO_1184 (O_1184,N_14155,N_14336);
and UO_1185 (O_1185,N_14969,N_14334);
nand UO_1186 (O_1186,N_14301,N_14234);
nor UO_1187 (O_1187,N_14163,N_14892);
nor UO_1188 (O_1188,N_14344,N_14989);
nand UO_1189 (O_1189,N_14652,N_14170);
or UO_1190 (O_1190,N_14939,N_14745);
or UO_1191 (O_1191,N_14232,N_14224);
and UO_1192 (O_1192,N_14506,N_14788);
nand UO_1193 (O_1193,N_14768,N_14716);
nand UO_1194 (O_1194,N_14242,N_14682);
xor UO_1195 (O_1195,N_14493,N_14313);
or UO_1196 (O_1196,N_14331,N_14111);
nand UO_1197 (O_1197,N_14065,N_14611);
xor UO_1198 (O_1198,N_14820,N_14036);
and UO_1199 (O_1199,N_14521,N_14010);
and UO_1200 (O_1200,N_14541,N_14219);
xor UO_1201 (O_1201,N_14608,N_14585);
nand UO_1202 (O_1202,N_14197,N_14962);
or UO_1203 (O_1203,N_14272,N_14818);
and UO_1204 (O_1204,N_14863,N_14482);
nor UO_1205 (O_1205,N_14538,N_14355);
or UO_1206 (O_1206,N_14648,N_14460);
and UO_1207 (O_1207,N_14452,N_14325);
or UO_1208 (O_1208,N_14975,N_14891);
or UO_1209 (O_1209,N_14509,N_14167);
nand UO_1210 (O_1210,N_14829,N_14209);
nor UO_1211 (O_1211,N_14416,N_14856);
and UO_1212 (O_1212,N_14497,N_14576);
and UO_1213 (O_1213,N_14391,N_14401);
nand UO_1214 (O_1214,N_14034,N_14788);
nor UO_1215 (O_1215,N_14093,N_14578);
and UO_1216 (O_1216,N_14618,N_14817);
or UO_1217 (O_1217,N_14109,N_14075);
and UO_1218 (O_1218,N_14340,N_14294);
nor UO_1219 (O_1219,N_14864,N_14782);
xnor UO_1220 (O_1220,N_14429,N_14361);
nor UO_1221 (O_1221,N_14517,N_14121);
or UO_1222 (O_1222,N_14298,N_14245);
nor UO_1223 (O_1223,N_14692,N_14415);
or UO_1224 (O_1224,N_14433,N_14289);
nor UO_1225 (O_1225,N_14331,N_14815);
and UO_1226 (O_1226,N_14410,N_14385);
xnor UO_1227 (O_1227,N_14767,N_14127);
or UO_1228 (O_1228,N_14806,N_14750);
nor UO_1229 (O_1229,N_14462,N_14625);
or UO_1230 (O_1230,N_14907,N_14884);
or UO_1231 (O_1231,N_14931,N_14738);
and UO_1232 (O_1232,N_14559,N_14358);
nor UO_1233 (O_1233,N_14281,N_14689);
or UO_1234 (O_1234,N_14505,N_14552);
nor UO_1235 (O_1235,N_14423,N_14091);
nand UO_1236 (O_1236,N_14537,N_14230);
nand UO_1237 (O_1237,N_14623,N_14677);
xnor UO_1238 (O_1238,N_14460,N_14659);
and UO_1239 (O_1239,N_14115,N_14774);
or UO_1240 (O_1240,N_14475,N_14913);
nand UO_1241 (O_1241,N_14470,N_14453);
and UO_1242 (O_1242,N_14857,N_14734);
and UO_1243 (O_1243,N_14165,N_14538);
and UO_1244 (O_1244,N_14375,N_14625);
or UO_1245 (O_1245,N_14683,N_14258);
nand UO_1246 (O_1246,N_14943,N_14981);
nand UO_1247 (O_1247,N_14159,N_14826);
nor UO_1248 (O_1248,N_14389,N_14066);
xnor UO_1249 (O_1249,N_14911,N_14885);
xor UO_1250 (O_1250,N_14770,N_14484);
nand UO_1251 (O_1251,N_14911,N_14192);
nor UO_1252 (O_1252,N_14756,N_14840);
or UO_1253 (O_1253,N_14718,N_14490);
nand UO_1254 (O_1254,N_14091,N_14470);
and UO_1255 (O_1255,N_14418,N_14388);
nand UO_1256 (O_1256,N_14510,N_14407);
nor UO_1257 (O_1257,N_14813,N_14267);
or UO_1258 (O_1258,N_14926,N_14016);
xnor UO_1259 (O_1259,N_14855,N_14963);
or UO_1260 (O_1260,N_14894,N_14396);
nand UO_1261 (O_1261,N_14870,N_14415);
nand UO_1262 (O_1262,N_14545,N_14281);
xor UO_1263 (O_1263,N_14550,N_14697);
nor UO_1264 (O_1264,N_14463,N_14508);
nand UO_1265 (O_1265,N_14299,N_14626);
nand UO_1266 (O_1266,N_14174,N_14781);
or UO_1267 (O_1267,N_14975,N_14187);
nor UO_1268 (O_1268,N_14629,N_14670);
or UO_1269 (O_1269,N_14801,N_14467);
and UO_1270 (O_1270,N_14616,N_14433);
or UO_1271 (O_1271,N_14749,N_14360);
nand UO_1272 (O_1272,N_14190,N_14674);
nand UO_1273 (O_1273,N_14569,N_14561);
nor UO_1274 (O_1274,N_14590,N_14762);
and UO_1275 (O_1275,N_14196,N_14579);
and UO_1276 (O_1276,N_14213,N_14122);
or UO_1277 (O_1277,N_14291,N_14817);
and UO_1278 (O_1278,N_14780,N_14185);
nand UO_1279 (O_1279,N_14074,N_14834);
and UO_1280 (O_1280,N_14027,N_14043);
nor UO_1281 (O_1281,N_14899,N_14172);
nand UO_1282 (O_1282,N_14936,N_14958);
nor UO_1283 (O_1283,N_14507,N_14052);
nand UO_1284 (O_1284,N_14097,N_14414);
nor UO_1285 (O_1285,N_14273,N_14150);
nand UO_1286 (O_1286,N_14909,N_14390);
nor UO_1287 (O_1287,N_14586,N_14976);
and UO_1288 (O_1288,N_14470,N_14682);
nand UO_1289 (O_1289,N_14968,N_14171);
nor UO_1290 (O_1290,N_14011,N_14719);
nand UO_1291 (O_1291,N_14664,N_14747);
nand UO_1292 (O_1292,N_14577,N_14674);
xnor UO_1293 (O_1293,N_14691,N_14100);
nor UO_1294 (O_1294,N_14558,N_14849);
nor UO_1295 (O_1295,N_14642,N_14393);
nand UO_1296 (O_1296,N_14992,N_14486);
nand UO_1297 (O_1297,N_14585,N_14485);
nor UO_1298 (O_1298,N_14661,N_14906);
nand UO_1299 (O_1299,N_14036,N_14706);
nand UO_1300 (O_1300,N_14748,N_14220);
xor UO_1301 (O_1301,N_14068,N_14927);
nor UO_1302 (O_1302,N_14298,N_14304);
nand UO_1303 (O_1303,N_14742,N_14957);
nand UO_1304 (O_1304,N_14308,N_14869);
or UO_1305 (O_1305,N_14328,N_14562);
or UO_1306 (O_1306,N_14924,N_14617);
and UO_1307 (O_1307,N_14512,N_14231);
nor UO_1308 (O_1308,N_14953,N_14878);
and UO_1309 (O_1309,N_14519,N_14587);
and UO_1310 (O_1310,N_14141,N_14709);
xnor UO_1311 (O_1311,N_14449,N_14907);
nand UO_1312 (O_1312,N_14375,N_14219);
or UO_1313 (O_1313,N_14453,N_14522);
xor UO_1314 (O_1314,N_14863,N_14200);
xnor UO_1315 (O_1315,N_14073,N_14560);
and UO_1316 (O_1316,N_14914,N_14992);
nor UO_1317 (O_1317,N_14930,N_14394);
nand UO_1318 (O_1318,N_14133,N_14751);
or UO_1319 (O_1319,N_14811,N_14449);
and UO_1320 (O_1320,N_14537,N_14158);
or UO_1321 (O_1321,N_14619,N_14477);
nor UO_1322 (O_1322,N_14644,N_14656);
nand UO_1323 (O_1323,N_14745,N_14828);
and UO_1324 (O_1324,N_14556,N_14010);
or UO_1325 (O_1325,N_14244,N_14193);
nand UO_1326 (O_1326,N_14933,N_14542);
nand UO_1327 (O_1327,N_14552,N_14720);
nand UO_1328 (O_1328,N_14716,N_14481);
nand UO_1329 (O_1329,N_14221,N_14325);
nand UO_1330 (O_1330,N_14609,N_14218);
nand UO_1331 (O_1331,N_14981,N_14791);
and UO_1332 (O_1332,N_14544,N_14638);
nand UO_1333 (O_1333,N_14448,N_14337);
nor UO_1334 (O_1334,N_14449,N_14665);
nand UO_1335 (O_1335,N_14093,N_14911);
or UO_1336 (O_1336,N_14501,N_14851);
nor UO_1337 (O_1337,N_14491,N_14133);
nand UO_1338 (O_1338,N_14125,N_14448);
and UO_1339 (O_1339,N_14743,N_14467);
or UO_1340 (O_1340,N_14212,N_14615);
and UO_1341 (O_1341,N_14184,N_14899);
or UO_1342 (O_1342,N_14985,N_14839);
or UO_1343 (O_1343,N_14279,N_14177);
nor UO_1344 (O_1344,N_14411,N_14455);
nand UO_1345 (O_1345,N_14556,N_14883);
and UO_1346 (O_1346,N_14878,N_14223);
and UO_1347 (O_1347,N_14917,N_14117);
nand UO_1348 (O_1348,N_14675,N_14207);
or UO_1349 (O_1349,N_14503,N_14532);
nand UO_1350 (O_1350,N_14778,N_14983);
nand UO_1351 (O_1351,N_14731,N_14653);
xnor UO_1352 (O_1352,N_14148,N_14270);
or UO_1353 (O_1353,N_14376,N_14108);
and UO_1354 (O_1354,N_14434,N_14993);
and UO_1355 (O_1355,N_14610,N_14829);
nor UO_1356 (O_1356,N_14411,N_14406);
nor UO_1357 (O_1357,N_14554,N_14619);
nor UO_1358 (O_1358,N_14000,N_14485);
xor UO_1359 (O_1359,N_14053,N_14608);
xor UO_1360 (O_1360,N_14684,N_14107);
nor UO_1361 (O_1361,N_14403,N_14217);
or UO_1362 (O_1362,N_14849,N_14726);
and UO_1363 (O_1363,N_14731,N_14404);
nand UO_1364 (O_1364,N_14733,N_14522);
or UO_1365 (O_1365,N_14572,N_14706);
nand UO_1366 (O_1366,N_14086,N_14919);
or UO_1367 (O_1367,N_14755,N_14695);
or UO_1368 (O_1368,N_14794,N_14308);
nor UO_1369 (O_1369,N_14979,N_14033);
or UO_1370 (O_1370,N_14117,N_14078);
xnor UO_1371 (O_1371,N_14821,N_14547);
or UO_1372 (O_1372,N_14322,N_14729);
and UO_1373 (O_1373,N_14537,N_14305);
nor UO_1374 (O_1374,N_14431,N_14102);
nor UO_1375 (O_1375,N_14281,N_14560);
and UO_1376 (O_1376,N_14333,N_14766);
and UO_1377 (O_1377,N_14324,N_14614);
or UO_1378 (O_1378,N_14729,N_14960);
and UO_1379 (O_1379,N_14565,N_14843);
nor UO_1380 (O_1380,N_14290,N_14518);
and UO_1381 (O_1381,N_14787,N_14242);
xor UO_1382 (O_1382,N_14786,N_14866);
xnor UO_1383 (O_1383,N_14445,N_14303);
nor UO_1384 (O_1384,N_14407,N_14024);
nand UO_1385 (O_1385,N_14934,N_14459);
xnor UO_1386 (O_1386,N_14753,N_14125);
xor UO_1387 (O_1387,N_14900,N_14939);
and UO_1388 (O_1388,N_14183,N_14266);
nor UO_1389 (O_1389,N_14853,N_14268);
or UO_1390 (O_1390,N_14370,N_14816);
xnor UO_1391 (O_1391,N_14940,N_14335);
nand UO_1392 (O_1392,N_14195,N_14913);
nor UO_1393 (O_1393,N_14586,N_14428);
nand UO_1394 (O_1394,N_14030,N_14053);
or UO_1395 (O_1395,N_14230,N_14081);
xnor UO_1396 (O_1396,N_14288,N_14564);
and UO_1397 (O_1397,N_14701,N_14308);
nor UO_1398 (O_1398,N_14590,N_14275);
and UO_1399 (O_1399,N_14603,N_14324);
or UO_1400 (O_1400,N_14391,N_14639);
or UO_1401 (O_1401,N_14170,N_14835);
nand UO_1402 (O_1402,N_14309,N_14580);
or UO_1403 (O_1403,N_14982,N_14602);
and UO_1404 (O_1404,N_14410,N_14837);
nor UO_1405 (O_1405,N_14111,N_14936);
xor UO_1406 (O_1406,N_14898,N_14407);
nor UO_1407 (O_1407,N_14523,N_14891);
nand UO_1408 (O_1408,N_14440,N_14918);
or UO_1409 (O_1409,N_14315,N_14891);
or UO_1410 (O_1410,N_14883,N_14630);
nor UO_1411 (O_1411,N_14074,N_14389);
nor UO_1412 (O_1412,N_14755,N_14812);
or UO_1413 (O_1413,N_14095,N_14067);
nor UO_1414 (O_1414,N_14147,N_14612);
nand UO_1415 (O_1415,N_14027,N_14357);
or UO_1416 (O_1416,N_14279,N_14962);
and UO_1417 (O_1417,N_14114,N_14081);
and UO_1418 (O_1418,N_14629,N_14598);
and UO_1419 (O_1419,N_14343,N_14471);
nand UO_1420 (O_1420,N_14739,N_14760);
nand UO_1421 (O_1421,N_14269,N_14883);
and UO_1422 (O_1422,N_14811,N_14154);
nor UO_1423 (O_1423,N_14665,N_14475);
nor UO_1424 (O_1424,N_14833,N_14879);
xor UO_1425 (O_1425,N_14247,N_14886);
nor UO_1426 (O_1426,N_14434,N_14531);
nor UO_1427 (O_1427,N_14651,N_14569);
and UO_1428 (O_1428,N_14243,N_14320);
nand UO_1429 (O_1429,N_14339,N_14023);
or UO_1430 (O_1430,N_14015,N_14712);
xnor UO_1431 (O_1431,N_14271,N_14932);
or UO_1432 (O_1432,N_14728,N_14766);
and UO_1433 (O_1433,N_14867,N_14116);
and UO_1434 (O_1434,N_14128,N_14391);
nand UO_1435 (O_1435,N_14103,N_14519);
or UO_1436 (O_1436,N_14234,N_14103);
nor UO_1437 (O_1437,N_14596,N_14893);
and UO_1438 (O_1438,N_14385,N_14576);
or UO_1439 (O_1439,N_14511,N_14561);
nor UO_1440 (O_1440,N_14908,N_14329);
nor UO_1441 (O_1441,N_14323,N_14089);
and UO_1442 (O_1442,N_14987,N_14954);
xnor UO_1443 (O_1443,N_14908,N_14966);
or UO_1444 (O_1444,N_14913,N_14982);
and UO_1445 (O_1445,N_14282,N_14067);
nand UO_1446 (O_1446,N_14058,N_14605);
or UO_1447 (O_1447,N_14993,N_14842);
or UO_1448 (O_1448,N_14112,N_14329);
nor UO_1449 (O_1449,N_14368,N_14955);
nand UO_1450 (O_1450,N_14940,N_14018);
and UO_1451 (O_1451,N_14587,N_14155);
nor UO_1452 (O_1452,N_14481,N_14670);
nand UO_1453 (O_1453,N_14037,N_14376);
nand UO_1454 (O_1454,N_14073,N_14453);
nor UO_1455 (O_1455,N_14934,N_14127);
or UO_1456 (O_1456,N_14330,N_14789);
nor UO_1457 (O_1457,N_14847,N_14978);
nand UO_1458 (O_1458,N_14723,N_14553);
nand UO_1459 (O_1459,N_14802,N_14388);
nand UO_1460 (O_1460,N_14874,N_14014);
xor UO_1461 (O_1461,N_14632,N_14814);
nor UO_1462 (O_1462,N_14212,N_14471);
or UO_1463 (O_1463,N_14534,N_14071);
or UO_1464 (O_1464,N_14397,N_14984);
nand UO_1465 (O_1465,N_14216,N_14637);
nor UO_1466 (O_1466,N_14180,N_14716);
nor UO_1467 (O_1467,N_14758,N_14089);
xor UO_1468 (O_1468,N_14741,N_14988);
nor UO_1469 (O_1469,N_14230,N_14581);
nand UO_1470 (O_1470,N_14102,N_14575);
or UO_1471 (O_1471,N_14642,N_14389);
or UO_1472 (O_1472,N_14481,N_14694);
nor UO_1473 (O_1473,N_14948,N_14918);
xnor UO_1474 (O_1474,N_14944,N_14012);
or UO_1475 (O_1475,N_14329,N_14327);
nor UO_1476 (O_1476,N_14524,N_14372);
and UO_1477 (O_1477,N_14150,N_14554);
nand UO_1478 (O_1478,N_14803,N_14523);
nand UO_1479 (O_1479,N_14551,N_14190);
nor UO_1480 (O_1480,N_14228,N_14660);
or UO_1481 (O_1481,N_14573,N_14144);
nand UO_1482 (O_1482,N_14440,N_14526);
xnor UO_1483 (O_1483,N_14728,N_14757);
or UO_1484 (O_1484,N_14881,N_14794);
xor UO_1485 (O_1485,N_14962,N_14012);
nand UO_1486 (O_1486,N_14379,N_14936);
and UO_1487 (O_1487,N_14072,N_14725);
and UO_1488 (O_1488,N_14535,N_14940);
or UO_1489 (O_1489,N_14317,N_14308);
or UO_1490 (O_1490,N_14325,N_14777);
and UO_1491 (O_1491,N_14939,N_14461);
and UO_1492 (O_1492,N_14824,N_14081);
xor UO_1493 (O_1493,N_14148,N_14646);
and UO_1494 (O_1494,N_14326,N_14710);
nor UO_1495 (O_1495,N_14366,N_14051);
nor UO_1496 (O_1496,N_14250,N_14910);
xor UO_1497 (O_1497,N_14651,N_14256);
or UO_1498 (O_1498,N_14407,N_14149);
nand UO_1499 (O_1499,N_14238,N_14964);
or UO_1500 (O_1500,N_14609,N_14979);
or UO_1501 (O_1501,N_14563,N_14683);
nand UO_1502 (O_1502,N_14522,N_14977);
or UO_1503 (O_1503,N_14472,N_14193);
and UO_1504 (O_1504,N_14422,N_14599);
xor UO_1505 (O_1505,N_14232,N_14457);
nand UO_1506 (O_1506,N_14311,N_14940);
and UO_1507 (O_1507,N_14874,N_14138);
or UO_1508 (O_1508,N_14325,N_14282);
nor UO_1509 (O_1509,N_14338,N_14140);
nor UO_1510 (O_1510,N_14593,N_14672);
nand UO_1511 (O_1511,N_14391,N_14263);
nand UO_1512 (O_1512,N_14356,N_14068);
and UO_1513 (O_1513,N_14518,N_14933);
and UO_1514 (O_1514,N_14820,N_14735);
or UO_1515 (O_1515,N_14101,N_14192);
or UO_1516 (O_1516,N_14456,N_14181);
nor UO_1517 (O_1517,N_14696,N_14505);
and UO_1518 (O_1518,N_14431,N_14837);
nor UO_1519 (O_1519,N_14446,N_14830);
nor UO_1520 (O_1520,N_14248,N_14555);
nand UO_1521 (O_1521,N_14036,N_14448);
and UO_1522 (O_1522,N_14065,N_14963);
nand UO_1523 (O_1523,N_14403,N_14654);
nand UO_1524 (O_1524,N_14657,N_14970);
nor UO_1525 (O_1525,N_14641,N_14193);
nor UO_1526 (O_1526,N_14206,N_14939);
nor UO_1527 (O_1527,N_14245,N_14648);
nor UO_1528 (O_1528,N_14787,N_14012);
nor UO_1529 (O_1529,N_14592,N_14332);
or UO_1530 (O_1530,N_14143,N_14586);
xnor UO_1531 (O_1531,N_14924,N_14773);
and UO_1532 (O_1532,N_14440,N_14129);
nand UO_1533 (O_1533,N_14886,N_14828);
nand UO_1534 (O_1534,N_14857,N_14932);
nand UO_1535 (O_1535,N_14357,N_14283);
xor UO_1536 (O_1536,N_14540,N_14878);
nand UO_1537 (O_1537,N_14175,N_14197);
and UO_1538 (O_1538,N_14830,N_14339);
nand UO_1539 (O_1539,N_14913,N_14789);
or UO_1540 (O_1540,N_14365,N_14262);
nor UO_1541 (O_1541,N_14602,N_14716);
xnor UO_1542 (O_1542,N_14575,N_14512);
and UO_1543 (O_1543,N_14325,N_14057);
and UO_1544 (O_1544,N_14460,N_14870);
and UO_1545 (O_1545,N_14953,N_14058);
nor UO_1546 (O_1546,N_14734,N_14557);
nand UO_1547 (O_1547,N_14635,N_14451);
and UO_1548 (O_1548,N_14473,N_14102);
and UO_1549 (O_1549,N_14644,N_14139);
and UO_1550 (O_1550,N_14523,N_14153);
nand UO_1551 (O_1551,N_14840,N_14782);
nor UO_1552 (O_1552,N_14915,N_14292);
nor UO_1553 (O_1553,N_14182,N_14189);
and UO_1554 (O_1554,N_14096,N_14272);
xor UO_1555 (O_1555,N_14920,N_14371);
or UO_1556 (O_1556,N_14921,N_14665);
xnor UO_1557 (O_1557,N_14500,N_14490);
nand UO_1558 (O_1558,N_14374,N_14879);
nor UO_1559 (O_1559,N_14097,N_14693);
nor UO_1560 (O_1560,N_14110,N_14447);
nor UO_1561 (O_1561,N_14215,N_14031);
and UO_1562 (O_1562,N_14757,N_14746);
nor UO_1563 (O_1563,N_14935,N_14952);
nand UO_1564 (O_1564,N_14080,N_14801);
or UO_1565 (O_1565,N_14299,N_14950);
or UO_1566 (O_1566,N_14628,N_14254);
and UO_1567 (O_1567,N_14662,N_14078);
nand UO_1568 (O_1568,N_14386,N_14440);
and UO_1569 (O_1569,N_14073,N_14455);
xnor UO_1570 (O_1570,N_14589,N_14102);
and UO_1571 (O_1571,N_14884,N_14294);
nand UO_1572 (O_1572,N_14571,N_14159);
xor UO_1573 (O_1573,N_14109,N_14472);
nor UO_1574 (O_1574,N_14167,N_14289);
nor UO_1575 (O_1575,N_14243,N_14966);
and UO_1576 (O_1576,N_14541,N_14797);
nor UO_1577 (O_1577,N_14044,N_14383);
or UO_1578 (O_1578,N_14561,N_14941);
nand UO_1579 (O_1579,N_14787,N_14023);
nor UO_1580 (O_1580,N_14395,N_14475);
or UO_1581 (O_1581,N_14401,N_14553);
nand UO_1582 (O_1582,N_14525,N_14273);
or UO_1583 (O_1583,N_14881,N_14393);
nand UO_1584 (O_1584,N_14417,N_14630);
nor UO_1585 (O_1585,N_14797,N_14550);
nor UO_1586 (O_1586,N_14888,N_14302);
nor UO_1587 (O_1587,N_14809,N_14674);
nand UO_1588 (O_1588,N_14074,N_14911);
nor UO_1589 (O_1589,N_14737,N_14740);
nand UO_1590 (O_1590,N_14937,N_14492);
and UO_1591 (O_1591,N_14332,N_14411);
nand UO_1592 (O_1592,N_14083,N_14384);
and UO_1593 (O_1593,N_14077,N_14577);
or UO_1594 (O_1594,N_14963,N_14893);
and UO_1595 (O_1595,N_14140,N_14714);
or UO_1596 (O_1596,N_14476,N_14718);
nor UO_1597 (O_1597,N_14661,N_14411);
xnor UO_1598 (O_1598,N_14895,N_14786);
nand UO_1599 (O_1599,N_14071,N_14222);
or UO_1600 (O_1600,N_14890,N_14982);
or UO_1601 (O_1601,N_14981,N_14422);
nand UO_1602 (O_1602,N_14815,N_14140);
nand UO_1603 (O_1603,N_14349,N_14365);
and UO_1604 (O_1604,N_14421,N_14949);
or UO_1605 (O_1605,N_14827,N_14206);
nor UO_1606 (O_1606,N_14194,N_14894);
and UO_1607 (O_1607,N_14688,N_14503);
nand UO_1608 (O_1608,N_14619,N_14656);
nand UO_1609 (O_1609,N_14516,N_14901);
nand UO_1610 (O_1610,N_14258,N_14666);
nand UO_1611 (O_1611,N_14112,N_14187);
and UO_1612 (O_1612,N_14799,N_14237);
or UO_1613 (O_1613,N_14105,N_14178);
xnor UO_1614 (O_1614,N_14583,N_14184);
nor UO_1615 (O_1615,N_14453,N_14812);
or UO_1616 (O_1616,N_14760,N_14527);
nor UO_1617 (O_1617,N_14699,N_14247);
or UO_1618 (O_1618,N_14739,N_14006);
or UO_1619 (O_1619,N_14022,N_14783);
or UO_1620 (O_1620,N_14655,N_14065);
and UO_1621 (O_1621,N_14014,N_14125);
and UO_1622 (O_1622,N_14970,N_14117);
or UO_1623 (O_1623,N_14412,N_14734);
or UO_1624 (O_1624,N_14884,N_14820);
or UO_1625 (O_1625,N_14108,N_14531);
nand UO_1626 (O_1626,N_14137,N_14735);
nor UO_1627 (O_1627,N_14210,N_14144);
nor UO_1628 (O_1628,N_14079,N_14347);
or UO_1629 (O_1629,N_14399,N_14398);
and UO_1630 (O_1630,N_14266,N_14448);
and UO_1631 (O_1631,N_14993,N_14535);
and UO_1632 (O_1632,N_14510,N_14498);
nor UO_1633 (O_1633,N_14186,N_14122);
nor UO_1634 (O_1634,N_14295,N_14941);
and UO_1635 (O_1635,N_14929,N_14280);
and UO_1636 (O_1636,N_14975,N_14154);
and UO_1637 (O_1637,N_14193,N_14213);
and UO_1638 (O_1638,N_14616,N_14701);
and UO_1639 (O_1639,N_14613,N_14541);
or UO_1640 (O_1640,N_14758,N_14129);
or UO_1641 (O_1641,N_14415,N_14996);
nand UO_1642 (O_1642,N_14462,N_14363);
nand UO_1643 (O_1643,N_14890,N_14115);
nand UO_1644 (O_1644,N_14251,N_14930);
and UO_1645 (O_1645,N_14940,N_14845);
nor UO_1646 (O_1646,N_14500,N_14416);
or UO_1647 (O_1647,N_14445,N_14790);
nor UO_1648 (O_1648,N_14616,N_14865);
and UO_1649 (O_1649,N_14872,N_14879);
nor UO_1650 (O_1650,N_14461,N_14189);
and UO_1651 (O_1651,N_14671,N_14119);
nor UO_1652 (O_1652,N_14801,N_14128);
or UO_1653 (O_1653,N_14917,N_14283);
or UO_1654 (O_1654,N_14182,N_14427);
nand UO_1655 (O_1655,N_14134,N_14267);
or UO_1656 (O_1656,N_14157,N_14581);
xor UO_1657 (O_1657,N_14471,N_14605);
or UO_1658 (O_1658,N_14921,N_14324);
and UO_1659 (O_1659,N_14995,N_14721);
or UO_1660 (O_1660,N_14850,N_14444);
xnor UO_1661 (O_1661,N_14145,N_14373);
xor UO_1662 (O_1662,N_14322,N_14825);
nor UO_1663 (O_1663,N_14431,N_14500);
nor UO_1664 (O_1664,N_14240,N_14620);
or UO_1665 (O_1665,N_14687,N_14529);
and UO_1666 (O_1666,N_14507,N_14360);
nand UO_1667 (O_1667,N_14730,N_14309);
or UO_1668 (O_1668,N_14455,N_14719);
nor UO_1669 (O_1669,N_14503,N_14602);
nor UO_1670 (O_1670,N_14965,N_14589);
nand UO_1671 (O_1671,N_14368,N_14615);
and UO_1672 (O_1672,N_14929,N_14137);
or UO_1673 (O_1673,N_14574,N_14729);
or UO_1674 (O_1674,N_14294,N_14917);
or UO_1675 (O_1675,N_14045,N_14891);
or UO_1676 (O_1676,N_14369,N_14526);
and UO_1677 (O_1677,N_14372,N_14320);
and UO_1678 (O_1678,N_14153,N_14892);
nand UO_1679 (O_1679,N_14006,N_14067);
nor UO_1680 (O_1680,N_14926,N_14635);
and UO_1681 (O_1681,N_14152,N_14135);
or UO_1682 (O_1682,N_14525,N_14008);
and UO_1683 (O_1683,N_14992,N_14511);
nor UO_1684 (O_1684,N_14793,N_14686);
nand UO_1685 (O_1685,N_14647,N_14539);
nand UO_1686 (O_1686,N_14601,N_14271);
nor UO_1687 (O_1687,N_14721,N_14236);
or UO_1688 (O_1688,N_14334,N_14022);
or UO_1689 (O_1689,N_14893,N_14525);
nand UO_1690 (O_1690,N_14369,N_14847);
nor UO_1691 (O_1691,N_14115,N_14655);
or UO_1692 (O_1692,N_14753,N_14778);
nand UO_1693 (O_1693,N_14776,N_14075);
nor UO_1694 (O_1694,N_14569,N_14527);
nor UO_1695 (O_1695,N_14911,N_14841);
and UO_1696 (O_1696,N_14218,N_14317);
or UO_1697 (O_1697,N_14262,N_14487);
nand UO_1698 (O_1698,N_14768,N_14788);
xor UO_1699 (O_1699,N_14029,N_14985);
nand UO_1700 (O_1700,N_14233,N_14410);
and UO_1701 (O_1701,N_14195,N_14612);
nor UO_1702 (O_1702,N_14859,N_14972);
xor UO_1703 (O_1703,N_14311,N_14378);
or UO_1704 (O_1704,N_14776,N_14544);
nand UO_1705 (O_1705,N_14686,N_14886);
nor UO_1706 (O_1706,N_14537,N_14304);
nand UO_1707 (O_1707,N_14057,N_14736);
xor UO_1708 (O_1708,N_14224,N_14998);
nand UO_1709 (O_1709,N_14372,N_14910);
xnor UO_1710 (O_1710,N_14765,N_14659);
and UO_1711 (O_1711,N_14488,N_14569);
nor UO_1712 (O_1712,N_14796,N_14382);
or UO_1713 (O_1713,N_14572,N_14040);
xnor UO_1714 (O_1714,N_14514,N_14012);
nand UO_1715 (O_1715,N_14803,N_14365);
nand UO_1716 (O_1716,N_14544,N_14378);
nand UO_1717 (O_1717,N_14834,N_14138);
nor UO_1718 (O_1718,N_14147,N_14889);
nand UO_1719 (O_1719,N_14233,N_14803);
or UO_1720 (O_1720,N_14510,N_14260);
and UO_1721 (O_1721,N_14481,N_14311);
nor UO_1722 (O_1722,N_14710,N_14155);
and UO_1723 (O_1723,N_14590,N_14011);
or UO_1724 (O_1724,N_14595,N_14070);
nand UO_1725 (O_1725,N_14926,N_14806);
or UO_1726 (O_1726,N_14273,N_14357);
nor UO_1727 (O_1727,N_14984,N_14908);
and UO_1728 (O_1728,N_14994,N_14034);
nor UO_1729 (O_1729,N_14992,N_14110);
or UO_1730 (O_1730,N_14641,N_14523);
and UO_1731 (O_1731,N_14856,N_14251);
or UO_1732 (O_1732,N_14682,N_14239);
nand UO_1733 (O_1733,N_14245,N_14424);
or UO_1734 (O_1734,N_14791,N_14109);
nand UO_1735 (O_1735,N_14324,N_14276);
nand UO_1736 (O_1736,N_14495,N_14677);
nor UO_1737 (O_1737,N_14694,N_14100);
xor UO_1738 (O_1738,N_14023,N_14866);
and UO_1739 (O_1739,N_14793,N_14220);
and UO_1740 (O_1740,N_14764,N_14607);
nor UO_1741 (O_1741,N_14282,N_14506);
and UO_1742 (O_1742,N_14413,N_14868);
nand UO_1743 (O_1743,N_14875,N_14180);
or UO_1744 (O_1744,N_14176,N_14761);
nand UO_1745 (O_1745,N_14483,N_14288);
or UO_1746 (O_1746,N_14260,N_14308);
nor UO_1747 (O_1747,N_14132,N_14007);
or UO_1748 (O_1748,N_14485,N_14789);
nor UO_1749 (O_1749,N_14784,N_14697);
and UO_1750 (O_1750,N_14217,N_14813);
and UO_1751 (O_1751,N_14638,N_14719);
nor UO_1752 (O_1752,N_14816,N_14138);
nand UO_1753 (O_1753,N_14050,N_14054);
nor UO_1754 (O_1754,N_14578,N_14435);
and UO_1755 (O_1755,N_14280,N_14824);
nor UO_1756 (O_1756,N_14681,N_14657);
nand UO_1757 (O_1757,N_14494,N_14194);
xor UO_1758 (O_1758,N_14425,N_14631);
nor UO_1759 (O_1759,N_14065,N_14603);
or UO_1760 (O_1760,N_14451,N_14893);
nand UO_1761 (O_1761,N_14832,N_14307);
and UO_1762 (O_1762,N_14169,N_14112);
nor UO_1763 (O_1763,N_14469,N_14675);
nor UO_1764 (O_1764,N_14219,N_14618);
and UO_1765 (O_1765,N_14099,N_14741);
nand UO_1766 (O_1766,N_14026,N_14987);
nor UO_1767 (O_1767,N_14332,N_14207);
or UO_1768 (O_1768,N_14923,N_14688);
nor UO_1769 (O_1769,N_14492,N_14402);
nand UO_1770 (O_1770,N_14087,N_14916);
nand UO_1771 (O_1771,N_14362,N_14654);
nor UO_1772 (O_1772,N_14970,N_14283);
nor UO_1773 (O_1773,N_14910,N_14126);
and UO_1774 (O_1774,N_14586,N_14649);
or UO_1775 (O_1775,N_14151,N_14225);
nand UO_1776 (O_1776,N_14827,N_14769);
xor UO_1777 (O_1777,N_14573,N_14668);
or UO_1778 (O_1778,N_14700,N_14129);
or UO_1779 (O_1779,N_14870,N_14616);
xnor UO_1780 (O_1780,N_14173,N_14880);
nand UO_1781 (O_1781,N_14641,N_14816);
or UO_1782 (O_1782,N_14031,N_14088);
nor UO_1783 (O_1783,N_14048,N_14824);
nor UO_1784 (O_1784,N_14934,N_14137);
nor UO_1785 (O_1785,N_14240,N_14252);
and UO_1786 (O_1786,N_14118,N_14695);
nand UO_1787 (O_1787,N_14896,N_14339);
nand UO_1788 (O_1788,N_14214,N_14035);
or UO_1789 (O_1789,N_14226,N_14146);
or UO_1790 (O_1790,N_14780,N_14983);
or UO_1791 (O_1791,N_14700,N_14191);
and UO_1792 (O_1792,N_14346,N_14507);
or UO_1793 (O_1793,N_14935,N_14789);
xor UO_1794 (O_1794,N_14374,N_14226);
nor UO_1795 (O_1795,N_14198,N_14494);
nand UO_1796 (O_1796,N_14905,N_14979);
and UO_1797 (O_1797,N_14086,N_14746);
or UO_1798 (O_1798,N_14449,N_14928);
or UO_1799 (O_1799,N_14201,N_14680);
nand UO_1800 (O_1800,N_14131,N_14313);
nand UO_1801 (O_1801,N_14241,N_14573);
nand UO_1802 (O_1802,N_14553,N_14211);
xnor UO_1803 (O_1803,N_14364,N_14599);
nor UO_1804 (O_1804,N_14094,N_14152);
or UO_1805 (O_1805,N_14132,N_14298);
or UO_1806 (O_1806,N_14136,N_14777);
nor UO_1807 (O_1807,N_14219,N_14200);
or UO_1808 (O_1808,N_14713,N_14456);
nor UO_1809 (O_1809,N_14601,N_14082);
xnor UO_1810 (O_1810,N_14489,N_14306);
xnor UO_1811 (O_1811,N_14175,N_14887);
and UO_1812 (O_1812,N_14601,N_14182);
or UO_1813 (O_1813,N_14623,N_14101);
or UO_1814 (O_1814,N_14926,N_14516);
nand UO_1815 (O_1815,N_14984,N_14301);
nand UO_1816 (O_1816,N_14692,N_14713);
nand UO_1817 (O_1817,N_14399,N_14370);
nor UO_1818 (O_1818,N_14646,N_14898);
nor UO_1819 (O_1819,N_14496,N_14296);
or UO_1820 (O_1820,N_14013,N_14711);
or UO_1821 (O_1821,N_14388,N_14238);
and UO_1822 (O_1822,N_14383,N_14256);
and UO_1823 (O_1823,N_14801,N_14629);
nand UO_1824 (O_1824,N_14937,N_14827);
or UO_1825 (O_1825,N_14268,N_14643);
nand UO_1826 (O_1826,N_14109,N_14084);
or UO_1827 (O_1827,N_14030,N_14882);
or UO_1828 (O_1828,N_14352,N_14446);
or UO_1829 (O_1829,N_14154,N_14921);
and UO_1830 (O_1830,N_14812,N_14928);
nand UO_1831 (O_1831,N_14840,N_14604);
or UO_1832 (O_1832,N_14212,N_14911);
nand UO_1833 (O_1833,N_14095,N_14914);
nor UO_1834 (O_1834,N_14883,N_14275);
nor UO_1835 (O_1835,N_14415,N_14263);
and UO_1836 (O_1836,N_14409,N_14659);
and UO_1837 (O_1837,N_14579,N_14956);
nor UO_1838 (O_1838,N_14614,N_14609);
or UO_1839 (O_1839,N_14770,N_14395);
nand UO_1840 (O_1840,N_14510,N_14657);
nor UO_1841 (O_1841,N_14490,N_14580);
and UO_1842 (O_1842,N_14145,N_14906);
xor UO_1843 (O_1843,N_14572,N_14294);
xor UO_1844 (O_1844,N_14195,N_14336);
xor UO_1845 (O_1845,N_14878,N_14402);
and UO_1846 (O_1846,N_14210,N_14551);
and UO_1847 (O_1847,N_14140,N_14355);
nor UO_1848 (O_1848,N_14365,N_14440);
nor UO_1849 (O_1849,N_14103,N_14857);
and UO_1850 (O_1850,N_14529,N_14833);
nand UO_1851 (O_1851,N_14456,N_14081);
xor UO_1852 (O_1852,N_14850,N_14755);
or UO_1853 (O_1853,N_14271,N_14032);
or UO_1854 (O_1854,N_14817,N_14641);
nand UO_1855 (O_1855,N_14054,N_14253);
nand UO_1856 (O_1856,N_14100,N_14910);
nor UO_1857 (O_1857,N_14590,N_14038);
nand UO_1858 (O_1858,N_14437,N_14342);
or UO_1859 (O_1859,N_14686,N_14089);
and UO_1860 (O_1860,N_14984,N_14632);
nand UO_1861 (O_1861,N_14549,N_14606);
xnor UO_1862 (O_1862,N_14171,N_14962);
and UO_1863 (O_1863,N_14284,N_14980);
xor UO_1864 (O_1864,N_14573,N_14945);
or UO_1865 (O_1865,N_14804,N_14404);
or UO_1866 (O_1866,N_14947,N_14913);
or UO_1867 (O_1867,N_14931,N_14308);
nor UO_1868 (O_1868,N_14704,N_14641);
nand UO_1869 (O_1869,N_14203,N_14005);
xor UO_1870 (O_1870,N_14262,N_14333);
and UO_1871 (O_1871,N_14344,N_14419);
and UO_1872 (O_1872,N_14996,N_14552);
nand UO_1873 (O_1873,N_14379,N_14890);
or UO_1874 (O_1874,N_14515,N_14174);
nand UO_1875 (O_1875,N_14451,N_14866);
nor UO_1876 (O_1876,N_14340,N_14665);
nor UO_1877 (O_1877,N_14923,N_14362);
or UO_1878 (O_1878,N_14983,N_14745);
and UO_1879 (O_1879,N_14244,N_14397);
or UO_1880 (O_1880,N_14630,N_14565);
nor UO_1881 (O_1881,N_14074,N_14904);
nand UO_1882 (O_1882,N_14277,N_14732);
and UO_1883 (O_1883,N_14588,N_14365);
or UO_1884 (O_1884,N_14383,N_14581);
and UO_1885 (O_1885,N_14045,N_14657);
or UO_1886 (O_1886,N_14098,N_14174);
xor UO_1887 (O_1887,N_14830,N_14751);
and UO_1888 (O_1888,N_14563,N_14243);
or UO_1889 (O_1889,N_14505,N_14963);
or UO_1890 (O_1890,N_14320,N_14048);
and UO_1891 (O_1891,N_14669,N_14679);
nor UO_1892 (O_1892,N_14302,N_14502);
nand UO_1893 (O_1893,N_14540,N_14424);
and UO_1894 (O_1894,N_14127,N_14121);
nand UO_1895 (O_1895,N_14826,N_14244);
nand UO_1896 (O_1896,N_14801,N_14123);
or UO_1897 (O_1897,N_14250,N_14524);
nor UO_1898 (O_1898,N_14961,N_14919);
nor UO_1899 (O_1899,N_14684,N_14923);
or UO_1900 (O_1900,N_14168,N_14596);
nand UO_1901 (O_1901,N_14648,N_14390);
nand UO_1902 (O_1902,N_14817,N_14624);
or UO_1903 (O_1903,N_14773,N_14236);
nor UO_1904 (O_1904,N_14545,N_14950);
nor UO_1905 (O_1905,N_14703,N_14552);
xnor UO_1906 (O_1906,N_14559,N_14368);
and UO_1907 (O_1907,N_14270,N_14294);
nor UO_1908 (O_1908,N_14709,N_14232);
xor UO_1909 (O_1909,N_14881,N_14209);
and UO_1910 (O_1910,N_14951,N_14431);
nand UO_1911 (O_1911,N_14841,N_14652);
and UO_1912 (O_1912,N_14469,N_14714);
or UO_1913 (O_1913,N_14931,N_14191);
nand UO_1914 (O_1914,N_14124,N_14932);
nand UO_1915 (O_1915,N_14042,N_14022);
and UO_1916 (O_1916,N_14564,N_14744);
and UO_1917 (O_1917,N_14060,N_14173);
or UO_1918 (O_1918,N_14993,N_14355);
xnor UO_1919 (O_1919,N_14017,N_14335);
nor UO_1920 (O_1920,N_14148,N_14417);
and UO_1921 (O_1921,N_14608,N_14830);
or UO_1922 (O_1922,N_14068,N_14162);
xor UO_1923 (O_1923,N_14325,N_14160);
or UO_1924 (O_1924,N_14732,N_14133);
and UO_1925 (O_1925,N_14752,N_14819);
nand UO_1926 (O_1926,N_14671,N_14238);
and UO_1927 (O_1927,N_14268,N_14796);
nand UO_1928 (O_1928,N_14418,N_14045);
nand UO_1929 (O_1929,N_14185,N_14896);
xor UO_1930 (O_1930,N_14619,N_14534);
nand UO_1931 (O_1931,N_14335,N_14373);
or UO_1932 (O_1932,N_14482,N_14400);
nor UO_1933 (O_1933,N_14158,N_14818);
nor UO_1934 (O_1934,N_14408,N_14478);
or UO_1935 (O_1935,N_14272,N_14796);
or UO_1936 (O_1936,N_14400,N_14575);
nand UO_1937 (O_1937,N_14557,N_14964);
nor UO_1938 (O_1938,N_14839,N_14947);
nor UO_1939 (O_1939,N_14408,N_14093);
xor UO_1940 (O_1940,N_14628,N_14796);
or UO_1941 (O_1941,N_14420,N_14345);
or UO_1942 (O_1942,N_14534,N_14417);
nand UO_1943 (O_1943,N_14091,N_14615);
or UO_1944 (O_1944,N_14380,N_14622);
or UO_1945 (O_1945,N_14736,N_14067);
nor UO_1946 (O_1946,N_14537,N_14969);
nor UO_1947 (O_1947,N_14655,N_14077);
and UO_1948 (O_1948,N_14788,N_14024);
nand UO_1949 (O_1949,N_14982,N_14551);
and UO_1950 (O_1950,N_14730,N_14738);
nand UO_1951 (O_1951,N_14497,N_14120);
or UO_1952 (O_1952,N_14931,N_14813);
nand UO_1953 (O_1953,N_14579,N_14927);
xor UO_1954 (O_1954,N_14246,N_14084);
xnor UO_1955 (O_1955,N_14238,N_14857);
nand UO_1956 (O_1956,N_14191,N_14875);
nand UO_1957 (O_1957,N_14818,N_14782);
nand UO_1958 (O_1958,N_14731,N_14847);
or UO_1959 (O_1959,N_14540,N_14806);
nand UO_1960 (O_1960,N_14112,N_14934);
nor UO_1961 (O_1961,N_14016,N_14872);
and UO_1962 (O_1962,N_14239,N_14473);
nor UO_1963 (O_1963,N_14575,N_14022);
nor UO_1964 (O_1964,N_14570,N_14818);
nor UO_1965 (O_1965,N_14825,N_14558);
nor UO_1966 (O_1966,N_14994,N_14158);
nand UO_1967 (O_1967,N_14386,N_14780);
or UO_1968 (O_1968,N_14553,N_14704);
nand UO_1969 (O_1969,N_14482,N_14106);
nor UO_1970 (O_1970,N_14653,N_14895);
nand UO_1971 (O_1971,N_14249,N_14730);
or UO_1972 (O_1972,N_14180,N_14789);
or UO_1973 (O_1973,N_14268,N_14672);
nand UO_1974 (O_1974,N_14101,N_14189);
or UO_1975 (O_1975,N_14654,N_14795);
or UO_1976 (O_1976,N_14479,N_14124);
and UO_1977 (O_1977,N_14570,N_14536);
nand UO_1978 (O_1978,N_14060,N_14820);
nand UO_1979 (O_1979,N_14327,N_14349);
nor UO_1980 (O_1980,N_14267,N_14426);
or UO_1981 (O_1981,N_14783,N_14130);
or UO_1982 (O_1982,N_14491,N_14920);
nand UO_1983 (O_1983,N_14978,N_14177);
and UO_1984 (O_1984,N_14113,N_14198);
nand UO_1985 (O_1985,N_14012,N_14792);
nor UO_1986 (O_1986,N_14668,N_14429);
nor UO_1987 (O_1987,N_14849,N_14489);
and UO_1988 (O_1988,N_14686,N_14671);
xnor UO_1989 (O_1989,N_14081,N_14561);
nor UO_1990 (O_1990,N_14985,N_14709);
nand UO_1991 (O_1991,N_14353,N_14485);
and UO_1992 (O_1992,N_14941,N_14053);
and UO_1993 (O_1993,N_14102,N_14417);
nor UO_1994 (O_1994,N_14960,N_14971);
nor UO_1995 (O_1995,N_14778,N_14502);
nor UO_1996 (O_1996,N_14864,N_14910);
nand UO_1997 (O_1997,N_14304,N_14790);
or UO_1998 (O_1998,N_14269,N_14045);
or UO_1999 (O_1999,N_14839,N_14103);
endmodule