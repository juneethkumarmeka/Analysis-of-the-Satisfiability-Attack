module basic_1000_10000_1500_4_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_782,In_176);
nand U1 (N_1,In_913,In_644);
and U2 (N_2,In_490,In_69);
nor U3 (N_3,In_338,In_511);
nand U4 (N_4,In_67,In_964);
nand U5 (N_5,In_992,In_610);
xor U6 (N_6,In_130,In_263);
nor U7 (N_7,In_286,In_862);
and U8 (N_8,In_800,In_932);
and U9 (N_9,In_354,In_600);
or U10 (N_10,In_816,In_659);
nor U11 (N_11,In_984,In_189);
nand U12 (N_12,In_145,In_47);
and U13 (N_13,In_438,In_572);
nor U14 (N_14,In_366,In_753);
and U15 (N_15,In_966,In_520);
nand U16 (N_16,In_685,In_714);
and U17 (N_17,In_805,In_298);
nand U18 (N_18,In_336,In_818);
nor U19 (N_19,In_206,In_751);
or U20 (N_20,In_726,In_17);
nand U21 (N_21,In_920,In_792);
nor U22 (N_22,In_916,In_537);
nor U23 (N_23,In_914,In_849);
or U24 (N_24,In_759,In_367);
or U25 (N_25,In_215,In_907);
or U26 (N_26,In_895,In_549);
and U27 (N_27,In_426,In_306);
nand U28 (N_28,In_276,In_404);
or U29 (N_29,In_140,In_789);
and U30 (N_30,In_975,In_936);
nor U31 (N_31,In_742,In_584);
or U32 (N_32,In_281,In_668);
and U33 (N_33,In_847,In_703);
and U34 (N_34,In_326,In_793);
and U35 (N_35,In_479,In_182);
or U36 (N_36,In_798,In_749);
xnor U37 (N_37,In_178,In_831);
and U38 (N_38,In_157,In_557);
nand U39 (N_39,In_829,In_440);
nand U40 (N_40,In_663,In_465);
and U41 (N_41,In_952,In_794);
nand U42 (N_42,In_321,In_629);
xor U43 (N_43,In_409,In_347);
nor U44 (N_44,In_233,In_962);
xor U45 (N_45,In_525,In_294);
or U46 (N_46,In_459,In_686);
or U47 (N_47,In_590,In_718);
and U48 (N_48,In_729,In_344);
nor U49 (N_49,In_78,In_356);
nor U50 (N_50,In_894,In_692);
or U51 (N_51,In_133,In_124);
nor U52 (N_52,In_425,In_160);
nand U53 (N_53,In_716,In_758);
nand U54 (N_54,In_407,In_436);
xor U55 (N_55,In_222,In_1);
and U56 (N_56,In_402,In_599);
xor U57 (N_57,In_823,In_117);
or U58 (N_58,In_987,In_672);
or U59 (N_59,In_583,In_710);
nor U60 (N_60,In_740,In_784);
nand U61 (N_61,In_587,In_567);
nor U62 (N_62,In_540,In_223);
nand U63 (N_63,In_555,In_566);
nor U64 (N_64,In_134,In_531);
nand U65 (N_65,In_314,In_589);
or U66 (N_66,In_18,In_494);
or U67 (N_67,In_447,In_395);
and U68 (N_68,In_397,In_528);
and U69 (N_69,In_99,In_614);
nand U70 (N_70,In_605,In_35);
or U71 (N_71,In_981,In_89);
nor U72 (N_72,In_899,In_448);
nor U73 (N_73,In_217,In_743);
and U74 (N_74,In_131,In_435);
nor U75 (N_75,In_876,In_390);
xor U76 (N_76,In_503,In_717);
and U77 (N_77,In_299,In_437);
or U78 (N_78,In_150,In_116);
or U79 (N_79,In_658,In_989);
and U80 (N_80,In_346,In_575);
and U81 (N_81,In_288,In_512);
and U82 (N_82,In_776,In_954);
and U83 (N_83,In_603,In_677);
and U84 (N_84,In_342,In_577);
nand U85 (N_85,In_161,In_240);
nor U86 (N_86,In_495,In_999);
nor U87 (N_87,In_12,In_845);
and U88 (N_88,In_15,In_735);
nand U89 (N_89,In_467,In_271);
or U90 (N_90,In_678,In_400);
or U91 (N_91,In_484,In_897);
xnor U92 (N_92,In_868,In_655);
nor U93 (N_93,In_227,In_543);
xnor U94 (N_94,In_834,In_188);
and U95 (N_95,In_126,In_98);
nand U96 (N_96,In_372,In_391);
nor U97 (N_97,In_348,In_880);
and U98 (N_98,In_754,In_451);
or U99 (N_99,In_660,In_921);
and U100 (N_100,In_934,In_41);
nand U101 (N_101,In_747,In_592);
nor U102 (N_102,In_807,In_838);
nor U103 (N_103,In_682,In_825);
nand U104 (N_104,In_602,In_449);
nand U105 (N_105,In_226,In_68);
xnor U106 (N_106,In_890,In_96);
and U107 (N_107,In_691,In_656);
or U108 (N_108,In_959,In_303);
and U109 (N_109,In_997,In_33);
nand U110 (N_110,In_219,In_679);
nor U111 (N_111,In_305,In_87);
or U112 (N_112,In_995,In_381);
xor U113 (N_113,In_302,In_159);
and U114 (N_114,In_637,In_115);
or U115 (N_115,In_273,In_983);
or U116 (N_116,In_455,In_2);
xnor U117 (N_117,In_486,In_766);
and U118 (N_118,In_25,In_576);
and U119 (N_119,In_214,In_120);
or U120 (N_120,In_196,In_421);
and U121 (N_121,In_260,In_42);
nor U122 (N_122,In_405,In_351);
and U123 (N_123,In_205,In_547);
nor U124 (N_124,In_380,In_257);
nand U125 (N_125,In_166,In_34);
and U126 (N_126,In_990,In_957);
nor U127 (N_127,In_413,In_284);
or U128 (N_128,In_396,In_700);
xor U129 (N_129,In_951,In_653);
or U130 (N_130,In_852,In_173);
nand U131 (N_131,In_755,In_993);
xnor U132 (N_132,In_593,In_739);
and U133 (N_133,In_869,In_77);
and U134 (N_134,In_345,In_97);
and U135 (N_135,In_171,In_596);
or U136 (N_136,In_536,In_974);
or U137 (N_137,In_522,In_300);
or U138 (N_138,In_184,In_725);
nor U139 (N_139,In_778,In_621);
and U140 (N_140,In_406,In_569);
or U141 (N_141,In_953,In_343);
nand U142 (N_142,In_943,In_103);
nand U143 (N_143,In_362,In_665);
nor U144 (N_144,In_927,In_195);
and U145 (N_145,In_243,In_462);
or U146 (N_146,In_330,In_86);
xor U147 (N_147,In_79,In_732);
xor U148 (N_148,In_388,In_606);
nand U149 (N_149,In_563,In_272);
or U150 (N_150,In_901,In_363);
nor U151 (N_151,In_369,In_349);
nor U152 (N_152,In_669,In_529);
nand U153 (N_153,In_118,In_382);
or U154 (N_154,In_452,In_822);
and U155 (N_155,In_379,In_239);
nand U156 (N_156,In_72,In_411);
and U157 (N_157,In_872,In_969);
nor U158 (N_158,In_616,In_197);
nand U159 (N_159,In_560,In_285);
nor U160 (N_160,In_82,In_374);
nor U161 (N_161,In_521,In_533);
nand U162 (N_162,In_724,In_450);
nor U163 (N_163,In_859,In_247);
nand U164 (N_164,In_339,In_323);
xnor U165 (N_165,In_552,In_481);
nor U166 (N_166,In_752,In_194);
or U167 (N_167,In_733,In_961);
nand U168 (N_168,In_444,In_358);
and U169 (N_169,In_854,In_52);
nand U170 (N_170,In_101,In_551);
xnor U171 (N_171,In_307,In_688);
or U172 (N_172,In_996,In_918);
nor U173 (N_173,In_162,In_279);
or U174 (N_174,In_891,In_698);
or U175 (N_175,In_635,In_169);
nand U176 (N_176,In_625,In_799);
nor U177 (N_177,In_628,In_333);
nand U178 (N_178,In_75,In_797);
nor U179 (N_179,In_327,In_43);
nor U180 (N_180,In_213,In_866);
nor U181 (N_181,In_627,In_251);
nor U182 (N_182,In_846,In_645);
and U183 (N_183,In_378,In_445);
xnor U184 (N_184,In_721,In_772);
nand U185 (N_185,In_295,In_225);
nor U186 (N_186,In_648,In_485);
or U187 (N_187,In_304,In_147);
and U188 (N_188,In_168,In_745);
or U189 (N_189,In_428,In_837);
nand U190 (N_190,In_882,In_22);
nor U191 (N_191,In_228,In_982);
nor U192 (N_192,In_308,In_550);
xor U193 (N_193,In_473,In_221);
and U194 (N_194,In_177,In_142);
or U195 (N_195,In_764,In_201);
nand U196 (N_196,In_938,In_350);
nor U197 (N_197,In_736,In_256);
nor U198 (N_198,In_209,In_453);
or U199 (N_199,In_242,In_611);
or U200 (N_200,In_274,In_49);
nand U201 (N_201,In_814,In_102);
nand U202 (N_202,In_879,In_657);
nor U203 (N_203,In_715,In_108);
or U204 (N_204,In_808,In_675);
nor U205 (N_205,In_942,In_492);
nor U206 (N_206,In_4,In_624);
nand U207 (N_207,In_867,In_463);
nor U208 (N_208,In_670,In_788);
or U209 (N_209,In_368,In_496);
nor U210 (N_210,In_387,In_640);
nand U211 (N_211,In_722,In_945);
nor U212 (N_212,In_191,In_950);
nand U213 (N_213,In_20,In_626);
or U214 (N_214,In_187,In_297);
nand U215 (N_215,In_579,In_73);
nor U216 (N_216,In_539,In_335);
or U217 (N_217,In_478,In_850);
and U218 (N_218,In_61,In_609);
nand U219 (N_219,In_141,In_940);
nand U220 (N_220,In_430,In_355);
or U221 (N_221,In_801,In_154);
nor U222 (N_222,In_59,In_865);
nand U223 (N_223,In_802,In_234);
and U224 (N_224,In_519,In_693);
and U225 (N_225,In_554,In_958);
xor U226 (N_226,In_332,In_873);
or U227 (N_227,In_482,In_418);
or U228 (N_228,In_694,In_229);
nor U229 (N_229,In_826,In_3);
and U230 (N_230,In_331,In_727);
or U231 (N_231,In_235,In_506);
and U232 (N_232,In_84,In_199);
nor U233 (N_233,In_896,In_8);
nor U234 (N_234,In_230,In_538);
or U235 (N_235,In_40,In_746);
nor U236 (N_236,In_965,In_948);
nor U237 (N_237,In_517,In_95);
xor U238 (N_238,In_900,In_530);
and U239 (N_239,In_713,In_483);
nor U240 (N_240,In_967,In_524);
nand U241 (N_241,In_149,In_877);
or U242 (N_242,In_887,In_32);
and U243 (N_243,In_119,In_851);
or U244 (N_244,In_631,In_647);
xnor U245 (N_245,In_5,In_991);
xor U246 (N_246,In_132,In_777);
or U247 (N_247,In_970,In_804);
or U248 (N_248,In_458,In_341);
nor U249 (N_249,In_289,In_889);
and U250 (N_250,In_128,In_246);
or U251 (N_251,In_269,In_19);
nand U252 (N_252,In_828,In_526);
nor U253 (N_253,In_16,In_139);
or U254 (N_254,In_787,In_283);
and U255 (N_255,In_121,In_109);
nor U256 (N_256,In_947,In_734);
nand U257 (N_257,In_412,In_919);
or U258 (N_258,In_471,In_137);
and U259 (N_259,In_666,In_662);
or U260 (N_260,In_280,In_401);
xnor U261 (N_261,In_158,In_56);
nor U262 (N_262,In_598,In_44);
xor U263 (N_263,In_472,In_10);
and U264 (N_264,In_886,In_90);
or U265 (N_265,In_972,In_296);
and U266 (N_266,In_844,In_237);
and U267 (N_267,In_697,In_744);
nor U268 (N_268,In_930,In_45);
or U269 (N_269,In_783,In_265);
nor U270 (N_270,In_671,In_29);
nand U271 (N_271,In_773,In_893);
xnor U272 (N_272,In_100,In_245);
and U273 (N_273,In_820,In_489);
nor U274 (N_274,In_85,In_291);
or U275 (N_275,In_619,In_443);
nor U276 (N_276,In_155,In_542);
and U277 (N_277,In_170,In_594);
or U278 (N_278,In_70,In_864);
or U279 (N_279,In_313,In_595);
nand U280 (N_280,In_705,In_558);
and U281 (N_281,In_803,In_293);
or U282 (N_282,In_48,In_192);
and U283 (N_283,In_216,In_586);
nand U284 (N_284,In_578,In_500);
and U285 (N_285,In_446,In_937);
and U286 (N_286,In_384,In_518);
nor U287 (N_287,In_875,In_433);
and U288 (N_288,In_534,In_750);
nor U289 (N_289,In_352,In_960);
xor U290 (N_290,In_241,In_708);
or U291 (N_291,In_701,In_357);
or U292 (N_292,In_232,In_819);
xnor U293 (N_293,In_224,In_806);
nand U294 (N_294,In_810,In_203);
nand U295 (N_295,In_337,In_0);
nor U296 (N_296,In_261,In_884);
nand U297 (N_297,In_253,In_264);
and U298 (N_298,In_856,In_135);
or U299 (N_299,In_687,In_591);
and U300 (N_300,In_353,In_39);
nand U301 (N_301,In_316,In_270);
nand U302 (N_302,In_27,In_419);
and U303 (N_303,In_902,In_699);
and U304 (N_304,In_979,In_870);
nand U305 (N_305,In_383,In_218);
xnor U306 (N_306,In_198,In_153);
nor U307 (N_307,In_516,In_46);
nand U308 (N_308,In_986,In_977);
nor U309 (N_309,In_988,In_23);
nor U310 (N_310,In_770,In_944);
and U311 (N_311,In_786,In_65);
nor U312 (N_312,In_664,In_290);
nand U313 (N_313,In_815,In_62);
nand U314 (N_314,In_597,In_607);
or U315 (N_315,In_277,In_994);
and U316 (N_316,In_207,In_985);
nor U317 (N_317,In_620,In_633);
and U318 (N_318,In_174,In_92);
and U319 (N_319,In_532,In_31);
xor U320 (N_320,In_709,In_535);
nand U321 (N_321,In_165,In_112);
xnor U322 (N_322,In_429,In_623);
nand U323 (N_323,In_202,In_386);
nand U324 (N_324,In_53,In_748);
and U325 (N_325,In_762,In_559);
nand U326 (N_326,In_11,In_278);
nand U327 (N_327,In_695,In_334);
nor U328 (N_328,In_564,In_50);
nor U329 (N_329,In_612,In_585);
and U330 (N_330,In_683,In_464);
nor U331 (N_331,In_910,In_978);
or U332 (N_332,In_136,In_220);
nor U333 (N_333,In_842,In_545);
nand U334 (N_334,In_172,In_185);
or U335 (N_335,In_457,In_561);
nand U336 (N_336,In_491,In_501);
nand U337 (N_337,In_676,In_649);
and U338 (N_338,In_833,In_630);
nand U339 (N_339,In_292,In_817);
or U340 (N_340,In_888,In_681);
or U341 (N_341,In_863,In_375);
or U342 (N_342,In_474,In_615);
or U343 (N_343,In_156,In_774);
nand U344 (N_344,In_915,In_779);
and U345 (N_345,In_325,In_638);
nand U346 (N_346,In_573,In_146);
or U347 (N_347,In_925,In_652);
nand U348 (N_348,In_427,In_38);
nand U349 (N_349,In_238,In_812);
and U350 (N_350,In_392,In_871);
or U351 (N_351,In_841,In_832);
nor U352 (N_352,In_371,In_127);
nand U353 (N_353,In_365,In_809);
nor U354 (N_354,In_582,In_416);
and U355 (N_355,In_393,In_874);
nor U356 (N_356,In_946,In_843);
nand U357 (N_357,In_499,In_939);
or U358 (N_358,In_36,In_81);
nand U359 (N_359,In_507,In_439);
and U360 (N_360,In_26,In_570);
nand U361 (N_361,In_180,In_608);
or U362 (N_362,In_175,In_152);
nor U363 (N_363,In_674,In_909);
or U364 (N_364,In_760,In_505);
nand U365 (N_365,In_861,In_183);
and U366 (N_366,In_267,In_309);
or U367 (N_367,In_642,In_475);
nor U368 (N_368,In_763,In_122);
and U369 (N_369,In_824,In_431);
nand U370 (N_370,In_636,In_312);
and U371 (N_371,In_768,In_556);
nand U372 (N_372,In_480,In_493);
nand U373 (N_373,In_14,In_696);
nand U374 (N_374,In_827,In_317);
nand U375 (N_375,In_604,In_310);
or U376 (N_376,In_254,In_167);
and U377 (N_377,In_477,In_148);
and U378 (N_378,In_37,In_468);
nand U379 (N_379,In_830,In_193);
or U380 (N_380,In_905,In_144);
and U381 (N_381,In_422,In_704);
and U382 (N_382,In_821,In_973);
nand U383 (N_383,In_104,In_963);
nor U384 (N_384,In_424,In_76);
and U385 (N_385,In_923,In_769);
xor U386 (N_386,In_340,In_641);
nand U387 (N_387,In_883,In_720);
and U388 (N_388,In_860,In_211);
nand U389 (N_389,In_487,In_903);
nand U390 (N_390,In_855,In_858);
and U391 (N_391,In_376,In_706);
or U392 (N_392,In_723,In_403);
nor U393 (N_393,In_58,In_83);
and U394 (N_394,In_885,In_30);
and U395 (N_395,In_684,In_780);
or U396 (N_396,In_622,In_498);
xor U397 (N_397,In_998,In_651);
nand U398 (N_398,In_208,In_730);
xnor U399 (N_399,In_574,In_527);
or U400 (N_400,In_661,In_931);
and U401 (N_401,In_839,In_926);
nor U402 (N_402,In_282,In_795);
and U403 (N_403,In_7,In_200);
or U404 (N_404,In_775,In_151);
or U405 (N_405,In_301,In_581);
or U406 (N_406,In_790,In_370);
nand U407 (N_407,In_466,In_924);
and U408 (N_408,In_255,In_568);
nand U409 (N_409,In_731,In_143);
xor U410 (N_410,In_508,In_711);
or U411 (N_411,In_66,In_588);
nand U412 (N_412,In_80,In_667);
nand U413 (N_413,In_728,In_911);
or U414 (N_414,In_21,In_617);
or U415 (N_415,In_24,In_250);
nand U416 (N_416,In_249,In_968);
nand U417 (N_417,In_510,In_571);
nand U418 (N_418,In_781,In_138);
and U419 (N_419,In_580,In_259);
nand U420 (N_420,In_553,In_107);
nand U421 (N_421,In_497,In_315);
and U422 (N_422,In_707,In_377);
nor U423 (N_423,In_976,In_476);
nor U424 (N_424,In_523,In_917);
nand U425 (N_425,In_423,In_385);
or U426 (N_426,In_761,In_318);
xnor U427 (N_427,In_892,In_231);
or U428 (N_428,In_935,In_544);
nand U429 (N_429,In_949,In_509);
xor U430 (N_430,In_324,In_361);
and U431 (N_431,In_634,In_88);
or U432 (N_432,In_181,In_771);
or U433 (N_433,In_971,In_359);
and U434 (N_434,In_513,In_712);
or U435 (N_435,In_129,In_114);
xor U436 (N_436,In_757,In_414);
nand U437 (N_437,In_63,In_646);
nand U438 (N_438,In_456,In_6);
or U439 (N_439,In_319,In_163);
and U440 (N_440,In_853,In_410);
nand U441 (N_441,In_904,In_650);
nand U442 (N_442,In_373,In_941);
nand U443 (N_443,In_186,In_125);
and U444 (N_444,In_791,In_565);
nor U445 (N_445,In_548,In_461);
nand U446 (N_446,In_248,In_955);
and U447 (N_447,In_13,In_111);
or U448 (N_448,In_737,In_618);
and U449 (N_449,In_639,In_204);
nor U450 (N_450,In_980,In_113);
and U451 (N_451,In_906,In_94);
and U452 (N_452,In_460,In_546);
and U453 (N_453,In_74,In_767);
or U454 (N_454,In_389,In_928);
or U455 (N_455,In_908,In_51);
or U456 (N_456,In_441,In_123);
nor U457 (N_457,In_244,In_702);
nand U458 (N_458,In_929,In_654);
or U459 (N_459,In_262,In_57);
and U460 (N_460,In_601,In_110);
and U461 (N_461,In_328,In_813);
and U462 (N_462,In_541,In_398);
and U463 (N_463,In_454,In_210);
and U464 (N_464,In_179,In_311);
or U465 (N_465,In_756,In_933);
nor U466 (N_466,In_266,In_322);
or U467 (N_467,In_690,In_765);
nand U468 (N_468,In_399,In_673);
xnor U469 (N_469,In_470,In_434);
or U470 (N_470,In_785,In_898);
or U471 (N_471,In_680,In_912);
nor U472 (N_472,In_835,In_836);
and U473 (N_473,In_54,In_275);
nor U474 (N_474,In_55,In_738);
or U475 (N_475,In_848,In_420);
xnor U476 (N_476,In_504,In_287);
and U477 (N_477,In_258,In_469);
xor U478 (N_478,In_922,In_91);
nand U479 (N_479,In_881,In_956);
or U480 (N_480,In_106,In_502);
or U481 (N_481,In_796,In_60);
nand U482 (N_482,In_857,In_632);
nor U483 (N_483,In_515,In_878);
and U484 (N_484,In_252,In_719);
or U485 (N_485,In_105,In_442);
nor U486 (N_486,In_613,In_236);
or U487 (N_487,In_190,In_432);
nor U488 (N_488,In_811,In_562);
nand U489 (N_489,In_514,In_320);
and U490 (N_490,In_408,In_364);
xnor U491 (N_491,In_9,In_741);
and U492 (N_492,In_394,In_488);
nor U493 (N_493,In_689,In_64);
xnor U494 (N_494,In_28,In_417);
nor U495 (N_495,In_329,In_415);
xor U496 (N_496,In_71,In_360);
and U497 (N_497,In_840,In_212);
or U498 (N_498,In_93,In_268);
nand U499 (N_499,In_643,In_164);
nand U500 (N_500,In_38,In_25);
xor U501 (N_501,In_879,In_383);
nor U502 (N_502,In_665,In_135);
and U503 (N_503,In_721,In_361);
or U504 (N_504,In_113,In_850);
nand U505 (N_505,In_117,In_322);
nor U506 (N_506,In_174,In_984);
xnor U507 (N_507,In_942,In_425);
and U508 (N_508,In_105,In_571);
nor U509 (N_509,In_53,In_264);
nand U510 (N_510,In_938,In_701);
or U511 (N_511,In_342,In_934);
nand U512 (N_512,In_598,In_845);
or U513 (N_513,In_565,In_16);
nand U514 (N_514,In_72,In_0);
nand U515 (N_515,In_823,In_347);
or U516 (N_516,In_11,In_577);
and U517 (N_517,In_22,In_351);
and U518 (N_518,In_482,In_771);
xnor U519 (N_519,In_569,In_150);
and U520 (N_520,In_792,In_166);
nor U521 (N_521,In_632,In_507);
and U522 (N_522,In_134,In_874);
nand U523 (N_523,In_273,In_675);
nand U524 (N_524,In_655,In_45);
nor U525 (N_525,In_749,In_535);
and U526 (N_526,In_941,In_312);
or U527 (N_527,In_947,In_855);
nor U528 (N_528,In_470,In_515);
nand U529 (N_529,In_724,In_721);
nor U530 (N_530,In_984,In_663);
xnor U531 (N_531,In_974,In_957);
and U532 (N_532,In_434,In_534);
and U533 (N_533,In_999,In_694);
xnor U534 (N_534,In_776,In_104);
nand U535 (N_535,In_828,In_662);
or U536 (N_536,In_334,In_999);
and U537 (N_537,In_700,In_226);
and U538 (N_538,In_93,In_549);
nor U539 (N_539,In_139,In_95);
nor U540 (N_540,In_885,In_983);
xnor U541 (N_541,In_22,In_318);
nor U542 (N_542,In_418,In_792);
nand U543 (N_543,In_957,In_333);
nand U544 (N_544,In_140,In_529);
nor U545 (N_545,In_174,In_882);
or U546 (N_546,In_136,In_98);
nor U547 (N_547,In_881,In_632);
nor U548 (N_548,In_413,In_670);
and U549 (N_549,In_740,In_451);
and U550 (N_550,In_378,In_154);
or U551 (N_551,In_380,In_970);
or U552 (N_552,In_824,In_168);
xor U553 (N_553,In_344,In_886);
nor U554 (N_554,In_762,In_734);
nor U555 (N_555,In_559,In_924);
nand U556 (N_556,In_529,In_974);
xnor U557 (N_557,In_46,In_786);
nor U558 (N_558,In_726,In_755);
and U559 (N_559,In_490,In_551);
xor U560 (N_560,In_865,In_414);
or U561 (N_561,In_999,In_521);
nor U562 (N_562,In_265,In_988);
and U563 (N_563,In_872,In_723);
nand U564 (N_564,In_386,In_727);
nand U565 (N_565,In_406,In_630);
and U566 (N_566,In_940,In_821);
or U567 (N_567,In_306,In_204);
or U568 (N_568,In_610,In_42);
nor U569 (N_569,In_118,In_651);
nand U570 (N_570,In_512,In_613);
nand U571 (N_571,In_159,In_207);
or U572 (N_572,In_509,In_363);
xnor U573 (N_573,In_834,In_454);
and U574 (N_574,In_635,In_568);
and U575 (N_575,In_759,In_627);
nand U576 (N_576,In_350,In_907);
and U577 (N_577,In_668,In_661);
nor U578 (N_578,In_393,In_714);
and U579 (N_579,In_72,In_533);
nand U580 (N_580,In_66,In_8);
or U581 (N_581,In_16,In_812);
nand U582 (N_582,In_511,In_777);
nand U583 (N_583,In_931,In_112);
or U584 (N_584,In_96,In_865);
nor U585 (N_585,In_480,In_531);
nor U586 (N_586,In_185,In_90);
nor U587 (N_587,In_292,In_90);
nor U588 (N_588,In_524,In_61);
nor U589 (N_589,In_726,In_475);
or U590 (N_590,In_566,In_633);
or U591 (N_591,In_817,In_236);
and U592 (N_592,In_442,In_752);
and U593 (N_593,In_843,In_450);
or U594 (N_594,In_567,In_746);
nand U595 (N_595,In_801,In_331);
nor U596 (N_596,In_380,In_491);
nor U597 (N_597,In_36,In_942);
and U598 (N_598,In_714,In_595);
nand U599 (N_599,In_189,In_943);
nor U600 (N_600,In_674,In_35);
or U601 (N_601,In_880,In_228);
and U602 (N_602,In_85,In_427);
nand U603 (N_603,In_954,In_596);
nand U604 (N_604,In_539,In_889);
and U605 (N_605,In_589,In_558);
nand U606 (N_606,In_439,In_119);
or U607 (N_607,In_395,In_892);
xnor U608 (N_608,In_54,In_488);
xor U609 (N_609,In_74,In_24);
nand U610 (N_610,In_665,In_589);
nand U611 (N_611,In_278,In_958);
xnor U612 (N_612,In_83,In_762);
or U613 (N_613,In_886,In_142);
nor U614 (N_614,In_645,In_489);
xnor U615 (N_615,In_586,In_725);
xnor U616 (N_616,In_908,In_793);
nand U617 (N_617,In_906,In_723);
nand U618 (N_618,In_530,In_301);
nor U619 (N_619,In_927,In_216);
and U620 (N_620,In_249,In_524);
xnor U621 (N_621,In_126,In_577);
and U622 (N_622,In_380,In_348);
or U623 (N_623,In_883,In_240);
xnor U624 (N_624,In_89,In_691);
or U625 (N_625,In_514,In_20);
and U626 (N_626,In_348,In_846);
and U627 (N_627,In_407,In_241);
nor U628 (N_628,In_932,In_881);
and U629 (N_629,In_920,In_710);
and U630 (N_630,In_56,In_883);
nor U631 (N_631,In_739,In_871);
nor U632 (N_632,In_576,In_821);
nand U633 (N_633,In_543,In_817);
nand U634 (N_634,In_862,In_904);
and U635 (N_635,In_187,In_333);
or U636 (N_636,In_829,In_341);
or U637 (N_637,In_78,In_966);
nor U638 (N_638,In_852,In_649);
and U639 (N_639,In_794,In_570);
or U640 (N_640,In_229,In_138);
or U641 (N_641,In_844,In_258);
nand U642 (N_642,In_112,In_612);
nor U643 (N_643,In_816,In_730);
nor U644 (N_644,In_703,In_981);
nand U645 (N_645,In_737,In_297);
nand U646 (N_646,In_363,In_285);
nand U647 (N_647,In_312,In_824);
or U648 (N_648,In_975,In_801);
nor U649 (N_649,In_919,In_472);
nand U650 (N_650,In_534,In_89);
or U651 (N_651,In_283,In_100);
nor U652 (N_652,In_184,In_803);
xnor U653 (N_653,In_638,In_342);
nor U654 (N_654,In_68,In_161);
and U655 (N_655,In_289,In_237);
nor U656 (N_656,In_653,In_914);
or U657 (N_657,In_904,In_735);
and U658 (N_658,In_291,In_318);
xnor U659 (N_659,In_923,In_142);
xnor U660 (N_660,In_806,In_962);
and U661 (N_661,In_398,In_829);
nand U662 (N_662,In_536,In_642);
or U663 (N_663,In_830,In_859);
nand U664 (N_664,In_813,In_186);
nand U665 (N_665,In_455,In_747);
nor U666 (N_666,In_0,In_647);
xor U667 (N_667,In_111,In_199);
and U668 (N_668,In_558,In_948);
or U669 (N_669,In_79,In_293);
nand U670 (N_670,In_185,In_910);
or U671 (N_671,In_282,In_526);
nor U672 (N_672,In_254,In_280);
and U673 (N_673,In_180,In_995);
xor U674 (N_674,In_503,In_136);
nand U675 (N_675,In_598,In_521);
xnor U676 (N_676,In_868,In_17);
and U677 (N_677,In_220,In_223);
and U678 (N_678,In_701,In_756);
nor U679 (N_679,In_487,In_361);
nor U680 (N_680,In_757,In_872);
nor U681 (N_681,In_353,In_800);
or U682 (N_682,In_848,In_237);
and U683 (N_683,In_46,In_384);
nand U684 (N_684,In_704,In_51);
nand U685 (N_685,In_454,In_378);
nand U686 (N_686,In_919,In_927);
and U687 (N_687,In_843,In_822);
nor U688 (N_688,In_317,In_208);
nor U689 (N_689,In_200,In_804);
nand U690 (N_690,In_542,In_186);
and U691 (N_691,In_268,In_21);
nor U692 (N_692,In_125,In_49);
or U693 (N_693,In_437,In_296);
nor U694 (N_694,In_14,In_304);
nand U695 (N_695,In_255,In_125);
nor U696 (N_696,In_342,In_389);
nor U697 (N_697,In_151,In_352);
xnor U698 (N_698,In_256,In_348);
or U699 (N_699,In_955,In_452);
nor U700 (N_700,In_482,In_779);
and U701 (N_701,In_946,In_377);
nor U702 (N_702,In_650,In_670);
and U703 (N_703,In_389,In_230);
or U704 (N_704,In_706,In_922);
nor U705 (N_705,In_809,In_700);
and U706 (N_706,In_402,In_192);
nand U707 (N_707,In_567,In_982);
xnor U708 (N_708,In_833,In_70);
nor U709 (N_709,In_309,In_727);
and U710 (N_710,In_785,In_35);
nand U711 (N_711,In_755,In_248);
nand U712 (N_712,In_615,In_627);
nor U713 (N_713,In_880,In_159);
xor U714 (N_714,In_864,In_443);
or U715 (N_715,In_151,In_896);
and U716 (N_716,In_222,In_15);
or U717 (N_717,In_915,In_24);
nor U718 (N_718,In_986,In_268);
or U719 (N_719,In_839,In_364);
and U720 (N_720,In_800,In_102);
nor U721 (N_721,In_66,In_946);
nand U722 (N_722,In_858,In_732);
and U723 (N_723,In_635,In_238);
nand U724 (N_724,In_831,In_361);
nand U725 (N_725,In_683,In_8);
and U726 (N_726,In_4,In_592);
or U727 (N_727,In_227,In_784);
nor U728 (N_728,In_797,In_199);
nand U729 (N_729,In_650,In_787);
or U730 (N_730,In_706,In_715);
and U731 (N_731,In_694,In_582);
or U732 (N_732,In_389,In_237);
nor U733 (N_733,In_780,In_555);
nand U734 (N_734,In_273,In_304);
or U735 (N_735,In_216,In_58);
or U736 (N_736,In_571,In_36);
and U737 (N_737,In_929,In_867);
nand U738 (N_738,In_447,In_209);
nor U739 (N_739,In_850,In_783);
or U740 (N_740,In_575,In_62);
nor U741 (N_741,In_51,In_290);
nor U742 (N_742,In_373,In_671);
nand U743 (N_743,In_691,In_441);
nand U744 (N_744,In_15,In_765);
nand U745 (N_745,In_957,In_637);
nor U746 (N_746,In_848,In_890);
and U747 (N_747,In_907,In_999);
or U748 (N_748,In_350,In_764);
nor U749 (N_749,In_901,In_292);
xor U750 (N_750,In_393,In_542);
and U751 (N_751,In_670,In_993);
or U752 (N_752,In_62,In_677);
nor U753 (N_753,In_345,In_538);
xnor U754 (N_754,In_38,In_279);
or U755 (N_755,In_491,In_588);
nand U756 (N_756,In_27,In_436);
nor U757 (N_757,In_506,In_385);
or U758 (N_758,In_744,In_198);
nor U759 (N_759,In_392,In_895);
nor U760 (N_760,In_807,In_581);
nor U761 (N_761,In_844,In_554);
nand U762 (N_762,In_489,In_14);
or U763 (N_763,In_446,In_601);
nand U764 (N_764,In_341,In_793);
and U765 (N_765,In_0,In_942);
and U766 (N_766,In_82,In_970);
nand U767 (N_767,In_478,In_819);
nor U768 (N_768,In_326,In_773);
or U769 (N_769,In_391,In_359);
or U770 (N_770,In_869,In_87);
nand U771 (N_771,In_873,In_104);
and U772 (N_772,In_939,In_891);
xnor U773 (N_773,In_79,In_859);
or U774 (N_774,In_39,In_89);
and U775 (N_775,In_545,In_801);
nor U776 (N_776,In_626,In_256);
or U777 (N_777,In_762,In_516);
or U778 (N_778,In_561,In_729);
nor U779 (N_779,In_582,In_246);
nand U780 (N_780,In_34,In_919);
nand U781 (N_781,In_592,In_290);
nor U782 (N_782,In_75,In_343);
nand U783 (N_783,In_514,In_426);
xnor U784 (N_784,In_321,In_471);
nand U785 (N_785,In_614,In_985);
or U786 (N_786,In_316,In_676);
nor U787 (N_787,In_799,In_207);
and U788 (N_788,In_803,In_876);
nor U789 (N_789,In_836,In_93);
nor U790 (N_790,In_716,In_887);
or U791 (N_791,In_983,In_620);
nand U792 (N_792,In_743,In_93);
nand U793 (N_793,In_904,In_377);
nor U794 (N_794,In_885,In_152);
nor U795 (N_795,In_870,In_923);
and U796 (N_796,In_496,In_40);
or U797 (N_797,In_895,In_132);
or U798 (N_798,In_565,In_275);
nand U799 (N_799,In_54,In_360);
and U800 (N_800,In_492,In_624);
nand U801 (N_801,In_754,In_70);
nor U802 (N_802,In_448,In_390);
nand U803 (N_803,In_428,In_641);
nand U804 (N_804,In_140,In_320);
nand U805 (N_805,In_313,In_41);
xnor U806 (N_806,In_405,In_280);
or U807 (N_807,In_203,In_300);
nor U808 (N_808,In_672,In_479);
or U809 (N_809,In_623,In_448);
and U810 (N_810,In_100,In_531);
and U811 (N_811,In_434,In_33);
nand U812 (N_812,In_48,In_253);
nand U813 (N_813,In_338,In_162);
xor U814 (N_814,In_123,In_349);
and U815 (N_815,In_256,In_895);
or U816 (N_816,In_851,In_70);
nand U817 (N_817,In_464,In_215);
nor U818 (N_818,In_403,In_568);
and U819 (N_819,In_155,In_667);
nand U820 (N_820,In_149,In_426);
xor U821 (N_821,In_940,In_418);
nand U822 (N_822,In_650,In_61);
xor U823 (N_823,In_704,In_726);
or U824 (N_824,In_621,In_134);
and U825 (N_825,In_664,In_865);
or U826 (N_826,In_164,In_244);
xnor U827 (N_827,In_672,In_571);
or U828 (N_828,In_748,In_667);
nor U829 (N_829,In_787,In_577);
and U830 (N_830,In_887,In_670);
or U831 (N_831,In_920,In_905);
and U832 (N_832,In_757,In_900);
and U833 (N_833,In_969,In_64);
and U834 (N_834,In_409,In_427);
nand U835 (N_835,In_171,In_83);
nor U836 (N_836,In_394,In_37);
nand U837 (N_837,In_312,In_311);
or U838 (N_838,In_193,In_218);
or U839 (N_839,In_764,In_486);
and U840 (N_840,In_983,In_471);
xnor U841 (N_841,In_345,In_826);
or U842 (N_842,In_916,In_842);
or U843 (N_843,In_21,In_981);
and U844 (N_844,In_979,In_157);
and U845 (N_845,In_880,In_314);
nor U846 (N_846,In_440,In_989);
nor U847 (N_847,In_796,In_115);
nor U848 (N_848,In_585,In_968);
or U849 (N_849,In_508,In_573);
and U850 (N_850,In_136,In_80);
and U851 (N_851,In_923,In_59);
nand U852 (N_852,In_862,In_659);
nand U853 (N_853,In_893,In_329);
or U854 (N_854,In_634,In_242);
and U855 (N_855,In_42,In_355);
nor U856 (N_856,In_849,In_122);
and U857 (N_857,In_691,In_598);
nand U858 (N_858,In_546,In_827);
nor U859 (N_859,In_70,In_604);
and U860 (N_860,In_585,In_271);
and U861 (N_861,In_251,In_914);
xor U862 (N_862,In_96,In_736);
or U863 (N_863,In_413,In_199);
or U864 (N_864,In_952,In_791);
and U865 (N_865,In_479,In_611);
or U866 (N_866,In_156,In_848);
or U867 (N_867,In_241,In_237);
or U868 (N_868,In_973,In_512);
nand U869 (N_869,In_348,In_971);
nor U870 (N_870,In_187,In_789);
or U871 (N_871,In_978,In_271);
xnor U872 (N_872,In_886,In_902);
xnor U873 (N_873,In_547,In_484);
nor U874 (N_874,In_957,In_810);
nand U875 (N_875,In_562,In_843);
nand U876 (N_876,In_260,In_413);
or U877 (N_877,In_849,In_560);
nor U878 (N_878,In_943,In_396);
nand U879 (N_879,In_741,In_363);
xor U880 (N_880,In_119,In_345);
or U881 (N_881,In_604,In_984);
and U882 (N_882,In_513,In_802);
nor U883 (N_883,In_236,In_862);
nor U884 (N_884,In_319,In_11);
or U885 (N_885,In_115,In_343);
and U886 (N_886,In_693,In_35);
nor U887 (N_887,In_526,In_26);
or U888 (N_888,In_757,In_570);
nand U889 (N_889,In_650,In_857);
nand U890 (N_890,In_933,In_139);
nand U891 (N_891,In_956,In_318);
nor U892 (N_892,In_788,In_391);
or U893 (N_893,In_320,In_846);
or U894 (N_894,In_383,In_870);
nor U895 (N_895,In_966,In_996);
or U896 (N_896,In_253,In_298);
nand U897 (N_897,In_426,In_812);
nand U898 (N_898,In_982,In_432);
nor U899 (N_899,In_270,In_466);
nand U900 (N_900,In_996,In_896);
nand U901 (N_901,In_275,In_455);
nand U902 (N_902,In_779,In_651);
nand U903 (N_903,In_888,In_575);
and U904 (N_904,In_981,In_979);
nand U905 (N_905,In_141,In_690);
or U906 (N_906,In_2,In_907);
or U907 (N_907,In_610,In_793);
or U908 (N_908,In_751,In_587);
nand U909 (N_909,In_840,In_433);
and U910 (N_910,In_693,In_967);
or U911 (N_911,In_474,In_918);
and U912 (N_912,In_844,In_392);
nor U913 (N_913,In_318,In_808);
or U914 (N_914,In_461,In_37);
nand U915 (N_915,In_718,In_446);
or U916 (N_916,In_55,In_877);
nor U917 (N_917,In_100,In_215);
or U918 (N_918,In_842,In_26);
nand U919 (N_919,In_545,In_747);
nand U920 (N_920,In_956,In_37);
nand U921 (N_921,In_517,In_153);
or U922 (N_922,In_159,In_933);
or U923 (N_923,In_954,In_680);
or U924 (N_924,In_655,In_915);
or U925 (N_925,In_66,In_510);
and U926 (N_926,In_481,In_546);
nor U927 (N_927,In_27,In_444);
nor U928 (N_928,In_762,In_358);
nand U929 (N_929,In_108,In_795);
or U930 (N_930,In_730,In_55);
xor U931 (N_931,In_392,In_729);
or U932 (N_932,In_893,In_185);
nand U933 (N_933,In_201,In_841);
and U934 (N_934,In_723,In_287);
and U935 (N_935,In_814,In_992);
and U936 (N_936,In_889,In_712);
and U937 (N_937,In_23,In_198);
nand U938 (N_938,In_585,In_776);
nor U939 (N_939,In_286,In_603);
nor U940 (N_940,In_214,In_607);
nor U941 (N_941,In_889,In_135);
nor U942 (N_942,In_854,In_206);
nor U943 (N_943,In_644,In_609);
or U944 (N_944,In_300,In_970);
and U945 (N_945,In_10,In_39);
nor U946 (N_946,In_18,In_252);
and U947 (N_947,In_183,In_56);
nand U948 (N_948,In_711,In_519);
nor U949 (N_949,In_718,In_656);
and U950 (N_950,In_339,In_903);
nand U951 (N_951,In_31,In_295);
and U952 (N_952,In_900,In_478);
nor U953 (N_953,In_771,In_137);
nor U954 (N_954,In_213,In_385);
or U955 (N_955,In_397,In_548);
nor U956 (N_956,In_682,In_899);
or U957 (N_957,In_496,In_304);
and U958 (N_958,In_403,In_14);
nor U959 (N_959,In_435,In_540);
nor U960 (N_960,In_605,In_932);
nor U961 (N_961,In_221,In_868);
nor U962 (N_962,In_435,In_309);
xor U963 (N_963,In_165,In_436);
or U964 (N_964,In_132,In_542);
nand U965 (N_965,In_261,In_551);
nand U966 (N_966,In_59,In_67);
or U967 (N_967,In_192,In_579);
or U968 (N_968,In_373,In_480);
xor U969 (N_969,In_420,In_299);
or U970 (N_970,In_299,In_646);
nor U971 (N_971,In_503,In_905);
and U972 (N_972,In_718,In_386);
or U973 (N_973,In_529,In_170);
or U974 (N_974,In_447,In_897);
nor U975 (N_975,In_824,In_689);
or U976 (N_976,In_636,In_97);
nor U977 (N_977,In_989,In_789);
nor U978 (N_978,In_512,In_337);
and U979 (N_979,In_998,In_388);
and U980 (N_980,In_875,In_387);
and U981 (N_981,In_83,In_154);
nor U982 (N_982,In_935,In_110);
and U983 (N_983,In_536,In_961);
nand U984 (N_984,In_885,In_496);
nand U985 (N_985,In_244,In_792);
nor U986 (N_986,In_723,In_767);
nor U987 (N_987,In_914,In_793);
and U988 (N_988,In_472,In_107);
and U989 (N_989,In_650,In_465);
and U990 (N_990,In_514,In_79);
and U991 (N_991,In_307,In_710);
nand U992 (N_992,In_500,In_965);
and U993 (N_993,In_341,In_35);
nand U994 (N_994,In_635,In_342);
nand U995 (N_995,In_235,In_419);
nor U996 (N_996,In_108,In_192);
nor U997 (N_997,In_983,In_545);
and U998 (N_998,In_549,In_701);
nor U999 (N_999,In_155,In_701);
nor U1000 (N_1000,In_926,In_165);
and U1001 (N_1001,In_748,In_25);
nand U1002 (N_1002,In_978,In_357);
nand U1003 (N_1003,In_909,In_794);
nor U1004 (N_1004,In_888,In_830);
nor U1005 (N_1005,In_216,In_25);
or U1006 (N_1006,In_354,In_185);
xnor U1007 (N_1007,In_342,In_321);
and U1008 (N_1008,In_351,In_933);
or U1009 (N_1009,In_178,In_853);
or U1010 (N_1010,In_534,In_970);
or U1011 (N_1011,In_181,In_150);
and U1012 (N_1012,In_83,In_458);
nand U1013 (N_1013,In_725,In_377);
or U1014 (N_1014,In_435,In_469);
nand U1015 (N_1015,In_123,In_510);
or U1016 (N_1016,In_379,In_879);
or U1017 (N_1017,In_765,In_251);
or U1018 (N_1018,In_671,In_303);
and U1019 (N_1019,In_680,In_51);
or U1020 (N_1020,In_805,In_831);
xnor U1021 (N_1021,In_1,In_267);
and U1022 (N_1022,In_174,In_722);
nor U1023 (N_1023,In_548,In_497);
nand U1024 (N_1024,In_86,In_230);
nor U1025 (N_1025,In_893,In_595);
xnor U1026 (N_1026,In_970,In_4);
or U1027 (N_1027,In_376,In_995);
nor U1028 (N_1028,In_534,In_11);
and U1029 (N_1029,In_122,In_142);
nor U1030 (N_1030,In_201,In_995);
xnor U1031 (N_1031,In_679,In_997);
xor U1032 (N_1032,In_195,In_394);
nand U1033 (N_1033,In_812,In_136);
nand U1034 (N_1034,In_184,In_228);
nor U1035 (N_1035,In_311,In_680);
or U1036 (N_1036,In_802,In_820);
and U1037 (N_1037,In_745,In_56);
nor U1038 (N_1038,In_749,In_928);
nand U1039 (N_1039,In_427,In_834);
and U1040 (N_1040,In_9,In_438);
nand U1041 (N_1041,In_354,In_38);
nor U1042 (N_1042,In_912,In_919);
or U1043 (N_1043,In_241,In_423);
or U1044 (N_1044,In_97,In_465);
or U1045 (N_1045,In_268,In_121);
or U1046 (N_1046,In_830,In_21);
and U1047 (N_1047,In_631,In_236);
or U1048 (N_1048,In_349,In_974);
and U1049 (N_1049,In_494,In_399);
nor U1050 (N_1050,In_375,In_93);
nand U1051 (N_1051,In_100,In_149);
or U1052 (N_1052,In_808,In_168);
or U1053 (N_1053,In_699,In_372);
or U1054 (N_1054,In_180,In_417);
and U1055 (N_1055,In_502,In_49);
nand U1056 (N_1056,In_70,In_368);
and U1057 (N_1057,In_566,In_613);
and U1058 (N_1058,In_38,In_342);
xnor U1059 (N_1059,In_827,In_361);
and U1060 (N_1060,In_679,In_274);
nor U1061 (N_1061,In_927,In_299);
xor U1062 (N_1062,In_658,In_450);
nor U1063 (N_1063,In_27,In_498);
nand U1064 (N_1064,In_147,In_733);
or U1065 (N_1065,In_221,In_226);
or U1066 (N_1066,In_820,In_690);
nand U1067 (N_1067,In_90,In_484);
nor U1068 (N_1068,In_230,In_853);
nor U1069 (N_1069,In_628,In_564);
or U1070 (N_1070,In_984,In_239);
or U1071 (N_1071,In_526,In_753);
and U1072 (N_1072,In_284,In_973);
nor U1073 (N_1073,In_831,In_618);
or U1074 (N_1074,In_10,In_458);
or U1075 (N_1075,In_613,In_75);
and U1076 (N_1076,In_443,In_183);
or U1077 (N_1077,In_213,In_834);
nand U1078 (N_1078,In_772,In_764);
and U1079 (N_1079,In_864,In_859);
nor U1080 (N_1080,In_733,In_589);
or U1081 (N_1081,In_370,In_174);
and U1082 (N_1082,In_57,In_613);
nand U1083 (N_1083,In_766,In_924);
or U1084 (N_1084,In_255,In_521);
xnor U1085 (N_1085,In_295,In_419);
nor U1086 (N_1086,In_647,In_544);
nor U1087 (N_1087,In_886,In_168);
and U1088 (N_1088,In_46,In_885);
xnor U1089 (N_1089,In_739,In_966);
nor U1090 (N_1090,In_507,In_2);
and U1091 (N_1091,In_402,In_564);
and U1092 (N_1092,In_971,In_323);
nor U1093 (N_1093,In_903,In_587);
and U1094 (N_1094,In_420,In_520);
or U1095 (N_1095,In_949,In_278);
or U1096 (N_1096,In_927,In_199);
or U1097 (N_1097,In_386,In_601);
nand U1098 (N_1098,In_646,In_554);
nor U1099 (N_1099,In_955,In_352);
nand U1100 (N_1100,In_416,In_550);
or U1101 (N_1101,In_969,In_949);
nand U1102 (N_1102,In_502,In_947);
nand U1103 (N_1103,In_261,In_7);
nor U1104 (N_1104,In_63,In_711);
or U1105 (N_1105,In_627,In_123);
or U1106 (N_1106,In_158,In_201);
or U1107 (N_1107,In_242,In_298);
nand U1108 (N_1108,In_363,In_535);
nand U1109 (N_1109,In_952,In_893);
or U1110 (N_1110,In_247,In_64);
nand U1111 (N_1111,In_746,In_526);
and U1112 (N_1112,In_814,In_122);
nor U1113 (N_1113,In_544,In_828);
nand U1114 (N_1114,In_789,In_776);
nand U1115 (N_1115,In_274,In_393);
nor U1116 (N_1116,In_827,In_243);
and U1117 (N_1117,In_819,In_954);
nor U1118 (N_1118,In_410,In_475);
or U1119 (N_1119,In_495,In_829);
nor U1120 (N_1120,In_449,In_543);
nand U1121 (N_1121,In_536,In_888);
and U1122 (N_1122,In_274,In_423);
nor U1123 (N_1123,In_404,In_231);
or U1124 (N_1124,In_844,In_214);
nand U1125 (N_1125,In_842,In_890);
nor U1126 (N_1126,In_482,In_927);
or U1127 (N_1127,In_559,In_423);
nand U1128 (N_1128,In_458,In_567);
or U1129 (N_1129,In_861,In_449);
nand U1130 (N_1130,In_831,In_741);
or U1131 (N_1131,In_516,In_717);
or U1132 (N_1132,In_790,In_777);
and U1133 (N_1133,In_912,In_402);
nand U1134 (N_1134,In_120,In_193);
nand U1135 (N_1135,In_571,In_400);
nor U1136 (N_1136,In_981,In_623);
or U1137 (N_1137,In_343,In_807);
nand U1138 (N_1138,In_623,In_963);
and U1139 (N_1139,In_753,In_847);
or U1140 (N_1140,In_208,In_424);
nand U1141 (N_1141,In_570,In_921);
and U1142 (N_1142,In_154,In_993);
xnor U1143 (N_1143,In_956,In_909);
and U1144 (N_1144,In_151,In_570);
nand U1145 (N_1145,In_557,In_856);
nand U1146 (N_1146,In_726,In_466);
and U1147 (N_1147,In_577,In_370);
xor U1148 (N_1148,In_991,In_58);
nor U1149 (N_1149,In_227,In_428);
and U1150 (N_1150,In_903,In_677);
nor U1151 (N_1151,In_868,In_762);
or U1152 (N_1152,In_942,In_162);
xor U1153 (N_1153,In_533,In_837);
nand U1154 (N_1154,In_8,In_420);
nand U1155 (N_1155,In_280,In_607);
nand U1156 (N_1156,In_326,In_116);
nor U1157 (N_1157,In_808,In_660);
nand U1158 (N_1158,In_886,In_505);
or U1159 (N_1159,In_152,In_564);
or U1160 (N_1160,In_467,In_912);
and U1161 (N_1161,In_304,In_377);
and U1162 (N_1162,In_155,In_578);
nor U1163 (N_1163,In_556,In_305);
or U1164 (N_1164,In_166,In_636);
nor U1165 (N_1165,In_777,In_7);
nand U1166 (N_1166,In_155,In_99);
nand U1167 (N_1167,In_204,In_490);
xnor U1168 (N_1168,In_803,In_468);
and U1169 (N_1169,In_575,In_618);
and U1170 (N_1170,In_99,In_769);
nor U1171 (N_1171,In_993,In_324);
or U1172 (N_1172,In_472,In_743);
nand U1173 (N_1173,In_431,In_333);
nand U1174 (N_1174,In_370,In_392);
nand U1175 (N_1175,In_652,In_795);
nand U1176 (N_1176,In_955,In_982);
nor U1177 (N_1177,In_229,In_134);
nand U1178 (N_1178,In_86,In_68);
nand U1179 (N_1179,In_692,In_66);
and U1180 (N_1180,In_244,In_715);
or U1181 (N_1181,In_112,In_908);
nand U1182 (N_1182,In_292,In_99);
or U1183 (N_1183,In_525,In_833);
and U1184 (N_1184,In_407,In_448);
nand U1185 (N_1185,In_235,In_925);
nor U1186 (N_1186,In_779,In_62);
or U1187 (N_1187,In_209,In_650);
and U1188 (N_1188,In_124,In_137);
xor U1189 (N_1189,In_669,In_701);
and U1190 (N_1190,In_523,In_835);
or U1191 (N_1191,In_217,In_565);
nor U1192 (N_1192,In_609,In_607);
xor U1193 (N_1193,In_628,In_704);
and U1194 (N_1194,In_127,In_939);
nand U1195 (N_1195,In_295,In_827);
and U1196 (N_1196,In_479,In_765);
nand U1197 (N_1197,In_71,In_108);
and U1198 (N_1198,In_206,In_783);
nor U1199 (N_1199,In_90,In_610);
nor U1200 (N_1200,In_335,In_682);
or U1201 (N_1201,In_631,In_242);
nor U1202 (N_1202,In_776,In_406);
nor U1203 (N_1203,In_636,In_179);
or U1204 (N_1204,In_960,In_611);
xor U1205 (N_1205,In_527,In_591);
nand U1206 (N_1206,In_151,In_310);
nor U1207 (N_1207,In_445,In_330);
nand U1208 (N_1208,In_509,In_909);
nand U1209 (N_1209,In_204,In_643);
nor U1210 (N_1210,In_149,In_863);
or U1211 (N_1211,In_524,In_282);
or U1212 (N_1212,In_27,In_420);
or U1213 (N_1213,In_438,In_970);
or U1214 (N_1214,In_625,In_209);
nand U1215 (N_1215,In_628,In_567);
and U1216 (N_1216,In_697,In_905);
nor U1217 (N_1217,In_938,In_76);
nor U1218 (N_1218,In_7,In_272);
or U1219 (N_1219,In_559,In_966);
nand U1220 (N_1220,In_901,In_52);
or U1221 (N_1221,In_628,In_917);
nor U1222 (N_1222,In_29,In_783);
nor U1223 (N_1223,In_57,In_424);
or U1224 (N_1224,In_398,In_210);
nand U1225 (N_1225,In_621,In_815);
and U1226 (N_1226,In_368,In_753);
or U1227 (N_1227,In_59,In_538);
and U1228 (N_1228,In_815,In_295);
nor U1229 (N_1229,In_279,In_55);
nor U1230 (N_1230,In_553,In_370);
nor U1231 (N_1231,In_550,In_407);
or U1232 (N_1232,In_379,In_722);
or U1233 (N_1233,In_887,In_240);
nand U1234 (N_1234,In_811,In_679);
and U1235 (N_1235,In_46,In_379);
nand U1236 (N_1236,In_57,In_645);
or U1237 (N_1237,In_795,In_800);
and U1238 (N_1238,In_625,In_630);
xor U1239 (N_1239,In_370,In_574);
nand U1240 (N_1240,In_720,In_27);
nor U1241 (N_1241,In_804,In_361);
nor U1242 (N_1242,In_103,In_618);
and U1243 (N_1243,In_589,In_365);
nand U1244 (N_1244,In_350,In_120);
and U1245 (N_1245,In_684,In_334);
or U1246 (N_1246,In_345,In_251);
nand U1247 (N_1247,In_211,In_278);
xor U1248 (N_1248,In_355,In_465);
nor U1249 (N_1249,In_940,In_21);
or U1250 (N_1250,In_706,In_624);
nand U1251 (N_1251,In_345,In_562);
nor U1252 (N_1252,In_419,In_154);
xor U1253 (N_1253,In_561,In_393);
nand U1254 (N_1254,In_259,In_631);
nand U1255 (N_1255,In_877,In_484);
and U1256 (N_1256,In_576,In_843);
or U1257 (N_1257,In_867,In_343);
xnor U1258 (N_1258,In_700,In_57);
and U1259 (N_1259,In_380,In_992);
nor U1260 (N_1260,In_447,In_280);
nand U1261 (N_1261,In_886,In_562);
or U1262 (N_1262,In_893,In_241);
nor U1263 (N_1263,In_673,In_761);
and U1264 (N_1264,In_993,In_772);
and U1265 (N_1265,In_628,In_107);
or U1266 (N_1266,In_326,In_201);
xor U1267 (N_1267,In_498,In_752);
nand U1268 (N_1268,In_260,In_778);
xnor U1269 (N_1269,In_19,In_610);
nand U1270 (N_1270,In_494,In_168);
nand U1271 (N_1271,In_824,In_218);
nand U1272 (N_1272,In_299,In_756);
or U1273 (N_1273,In_51,In_222);
nand U1274 (N_1274,In_994,In_468);
nand U1275 (N_1275,In_983,In_623);
nor U1276 (N_1276,In_445,In_287);
nand U1277 (N_1277,In_64,In_646);
nor U1278 (N_1278,In_600,In_257);
and U1279 (N_1279,In_396,In_331);
nor U1280 (N_1280,In_647,In_678);
nand U1281 (N_1281,In_470,In_79);
nor U1282 (N_1282,In_808,In_355);
xnor U1283 (N_1283,In_579,In_376);
and U1284 (N_1284,In_170,In_17);
or U1285 (N_1285,In_348,In_781);
or U1286 (N_1286,In_376,In_162);
nand U1287 (N_1287,In_334,In_836);
and U1288 (N_1288,In_204,In_163);
and U1289 (N_1289,In_306,In_310);
or U1290 (N_1290,In_550,In_488);
nor U1291 (N_1291,In_54,In_576);
nor U1292 (N_1292,In_754,In_646);
or U1293 (N_1293,In_396,In_723);
xnor U1294 (N_1294,In_772,In_173);
xnor U1295 (N_1295,In_358,In_822);
and U1296 (N_1296,In_927,In_761);
and U1297 (N_1297,In_350,In_484);
nor U1298 (N_1298,In_546,In_643);
and U1299 (N_1299,In_167,In_416);
nor U1300 (N_1300,In_519,In_773);
nand U1301 (N_1301,In_199,In_91);
and U1302 (N_1302,In_606,In_167);
or U1303 (N_1303,In_748,In_463);
nor U1304 (N_1304,In_393,In_860);
or U1305 (N_1305,In_168,In_816);
nand U1306 (N_1306,In_487,In_832);
xnor U1307 (N_1307,In_135,In_537);
nand U1308 (N_1308,In_85,In_643);
nor U1309 (N_1309,In_382,In_884);
and U1310 (N_1310,In_501,In_184);
nand U1311 (N_1311,In_952,In_517);
xor U1312 (N_1312,In_18,In_978);
or U1313 (N_1313,In_855,In_868);
nand U1314 (N_1314,In_141,In_895);
nand U1315 (N_1315,In_575,In_517);
and U1316 (N_1316,In_725,In_842);
nor U1317 (N_1317,In_769,In_663);
or U1318 (N_1318,In_995,In_167);
and U1319 (N_1319,In_13,In_771);
and U1320 (N_1320,In_569,In_377);
nor U1321 (N_1321,In_663,In_468);
or U1322 (N_1322,In_85,In_206);
nor U1323 (N_1323,In_588,In_702);
and U1324 (N_1324,In_573,In_848);
or U1325 (N_1325,In_647,In_375);
nor U1326 (N_1326,In_834,In_738);
nand U1327 (N_1327,In_514,In_83);
and U1328 (N_1328,In_343,In_805);
and U1329 (N_1329,In_858,In_492);
nand U1330 (N_1330,In_761,In_59);
nand U1331 (N_1331,In_947,In_903);
or U1332 (N_1332,In_234,In_138);
nor U1333 (N_1333,In_371,In_29);
nand U1334 (N_1334,In_296,In_562);
and U1335 (N_1335,In_263,In_229);
nor U1336 (N_1336,In_890,In_67);
and U1337 (N_1337,In_756,In_714);
nand U1338 (N_1338,In_247,In_394);
xnor U1339 (N_1339,In_76,In_239);
or U1340 (N_1340,In_873,In_856);
nor U1341 (N_1341,In_747,In_711);
nor U1342 (N_1342,In_798,In_878);
or U1343 (N_1343,In_53,In_612);
or U1344 (N_1344,In_56,In_127);
nor U1345 (N_1345,In_42,In_528);
nand U1346 (N_1346,In_378,In_853);
or U1347 (N_1347,In_645,In_434);
and U1348 (N_1348,In_292,In_272);
nand U1349 (N_1349,In_81,In_401);
nand U1350 (N_1350,In_497,In_221);
or U1351 (N_1351,In_619,In_316);
or U1352 (N_1352,In_193,In_159);
xnor U1353 (N_1353,In_426,In_209);
or U1354 (N_1354,In_228,In_113);
nand U1355 (N_1355,In_390,In_121);
and U1356 (N_1356,In_927,In_406);
and U1357 (N_1357,In_348,In_937);
nand U1358 (N_1358,In_32,In_586);
nor U1359 (N_1359,In_76,In_932);
and U1360 (N_1360,In_868,In_264);
or U1361 (N_1361,In_132,In_650);
nor U1362 (N_1362,In_126,In_340);
or U1363 (N_1363,In_143,In_677);
and U1364 (N_1364,In_89,In_583);
and U1365 (N_1365,In_709,In_787);
and U1366 (N_1366,In_306,In_965);
nor U1367 (N_1367,In_178,In_35);
and U1368 (N_1368,In_435,In_341);
and U1369 (N_1369,In_66,In_738);
and U1370 (N_1370,In_190,In_426);
and U1371 (N_1371,In_75,In_809);
or U1372 (N_1372,In_523,In_607);
nor U1373 (N_1373,In_806,In_135);
or U1374 (N_1374,In_450,In_322);
and U1375 (N_1375,In_650,In_25);
and U1376 (N_1376,In_275,In_941);
nor U1377 (N_1377,In_779,In_642);
xnor U1378 (N_1378,In_986,In_761);
and U1379 (N_1379,In_972,In_287);
nor U1380 (N_1380,In_412,In_854);
nor U1381 (N_1381,In_43,In_292);
nand U1382 (N_1382,In_662,In_466);
nor U1383 (N_1383,In_597,In_164);
nand U1384 (N_1384,In_823,In_225);
nor U1385 (N_1385,In_362,In_975);
nand U1386 (N_1386,In_666,In_959);
or U1387 (N_1387,In_273,In_560);
or U1388 (N_1388,In_376,In_763);
nor U1389 (N_1389,In_147,In_441);
and U1390 (N_1390,In_220,In_705);
nand U1391 (N_1391,In_797,In_89);
nand U1392 (N_1392,In_150,In_637);
nand U1393 (N_1393,In_753,In_178);
or U1394 (N_1394,In_258,In_165);
and U1395 (N_1395,In_494,In_247);
nand U1396 (N_1396,In_518,In_28);
and U1397 (N_1397,In_490,In_574);
nor U1398 (N_1398,In_994,In_769);
nand U1399 (N_1399,In_291,In_712);
and U1400 (N_1400,In_195,In_181);
or U1401 (N_1401,In_239,In_74);
and U1402 (N_1402,In_59,In_920);
or U1403 (N_1403,In_842,In_776);
nand U1404 (N_1404,In_962,In_859);
nor U1405 (N_1405,In_812,In_692);
nand U1406 (N_1406,In_468,In_219);
and U1407 (N_1407,In_715,In_707);
and U1408 (N_1408,In_701,In_134);
nor U1409 (N_1409,In_789,In_919);
nor U1410 (N_1410,In_602,In_130);
or U1411 (N_1411,In_197,In_160);
or U1412 (N_1412,In_357,In_321);
and U1413 (N_1413,In_976,In_680);
and U1414 (N_1414,In_261,In_896);
nor U1415 (N_1415,In_563,In_917);
nor U1416 (N_1416,In_817,In_349);
or U1417 (N_1417,In_657,In_60);
nand U1418 (N_1418,In_49,In_434);
or U1419 (N_1419,In_931,In_511);
nor U1420 (N_1420,In_788,In_467);
xor U1421 (N_1421,In_978,In_332);
xor U1422 (N_1422,In_833,In_505);
xor U1423 (N_1423,In_361,In_997);
or U1424 (N_1424,In_422,In_625);
nand U1425 (N_1425,In_259,In_579);
nand U1426 (N_1426,In_986,In_558);
or U1427 (N_1427,In_340,In_160);
xnor U1428 (N_1428,In_433,In_118);
nand U1429 (N_1429,In_773,In_500);
or U1430 (N_1430,In_70,In_18);
and U1431 (N_1431,In_372,In_158);
and U1432 (N_1432,In_11,In_42);
nor U1433 (N_1433,In_652,In_235);
or U1434 (N_1434,In_917,In_99);
nor U1435 (N_1435,In_632,In_613);
nor U1436 (N_1436,In_507,In_210);
nand U1437 (N_1437,In_303,In_510);
and U1438 (N_1438,In_512,In_353);
or U1439 (N_1439,In_895,In_811);
and U1440 (N_1440,In_948,In_477);
and U1441 (N_1441,In_564,In_478);
xor U1442 (N_1442,In_161,In_594);
nor U1443 (N_1443,In_934,In_592);
nor U1444 (N_1444,In_468,In_606);
nor U1445 (N_1445,In_270,In_705);
nand U1446 (N_1446,In_557,In_191);
and U1447 (N_1447,In_470,In_97);
xor U1448 (N_1448,In_835,In_809);
nand U1449 (N_1449,In_498,In_648);
and U1450 (N_1450,In_722,In_40);
nor U1451 (N_1451,In_688,In_359);
xnor U1452 (N_1452,In_507,In_97);
xnor U1453 (N_1453,In_27,In_761);
nor U1454 (N_1454,In_840,In_970);
nor U1455 (N_1455,In_239,In_603);
nand U1456 (N_1456,In_27,In_695);
nor U1457 (N_1457,In_78,In_492);
nor U1458 (N_1458,In_953,In_264);
or U1459 (N_1459,In_506,In_860);
and U1460 (N_1460,In_401,In_866);
nor U1461 (N_1461,In_131,In_926);
nor U1462 (N_1462,In_38,In_177);
or U1463 (N_1463,In_69,In_702);
nand U1464 (N_1464,In_342,In_100);
nand U1465 (N_1465,In_572,In_925);
nor U1466 (N_1466,In_107,In_581);
nand U1467 (N_1467,In_159,In_423);
nand U1468 (N_1468,In_11,In_834);
xor U1469 (N_1469,In_332,In_792);
nand U1470 (N_1470,In_800,In_976);
nor U1471 (N_1471,In_64,In_406);
and U1472 (N_1472,In_719,In_305);
and U1473 (N_1473,In_581,In_907);
nand U1474 (N_1474,In_629,In_899);
xnor U1475 (N_1475,In_450,In_164);
nor U1476 (N_1476,In_886,In_125);
nor U1477 (N_1477,In_732,In_908);
nor U1478 (N_1478,In_569,In_253);
xor U1479 (N_1479,In_530,In_451);
and U1480 (N_1480,In_156,In_296);
nand U1481 (N_1481,In_325,In_988);
xnor U1482 (N_1482,In_921,In_435);
nor U1483 (N_1483,In_707,In_994);
and U1484 (N_1484,In_531,In_185);
nand U1485 (N_1485,In_597,In_861);
nand U1486 (N_1486,In_867,In_202);
and U1487 (N_1487,In_592,In_286);
nand U1488 (N_1488,In_139,In_397);
nor U1489 (N_1489,In_234,In_509);
and U1490 (N_1490,In_445,In_503);
xor U1491 (N_1491,In_890,In_522);
or U1492 (N_1492,In_841,In_322);
nand U1493 (N_1493,In_548,In_513);
xor U1494 (N_1494,In_534,In_381);
or U1495 (N_1495,In_292,In_152);
nand U1496 (N_1496,In_704,In_533);
and U1497 (N_1497,In_327,In_901);
or U1498 (N_1498,In_426,In_453);
or U1499 (N_1499,In_522,In_365);
nor U1500 (N_1500,In_68,In_167);
or U1501 (N_1501,In_655,In_961);
nand U1502 (N_1502,In_940,In_596);
and U1503 (N_1503,In_104,In_448);
nor U1504 (N_1504,In_212,In_983);
and U1505 (N_1505,In_485,In_489);
nor U1506 (N_1506,In_481,In_970);
nand U1507 (N_1507,In_949,In_484);
nand U1508 (N_1508,In_775,In_15);
xnor U1509 (N_1509,In_600,In_754);
nand U1510 (N_1510,In_58,In_776);
xnor U1511 (N_1511,In_894,In_571);
nor U1512 (N_1512,In_520,In_946);
and U1513 (N_1513,In_190,In_446);
nand U1514 (N_1514,In_747,In_618);
and U1515 (N_1515,In_841,In_571);
nor U1516 (N_1516,In_808,In_451);
xnor U1517 (N_1517,In_319,In_512);
or U1518 (N_1518,In_49,In_784);
nor U1519 (N_1519,In_54,In_229);
nand U1520 (N_1520,In_938,In_544);
or U1521 (N_1521,In_794,In_332);
and U1522 (N_1522,In_640,In_527);
xnor U1523 (N_1523,In_366,In_36);
xnor U1524 (N_1524,In_961,In_563);
and U1525 (N_1525,In_839,In_153);
and U1526 (N_1526,In_383,In_547);
or U1527 (N_1527,In_367,In_217);
nand U1528 (N_1528,In_58,In_751);
or U1529 (N_1529,In_337,In_331);
or U1530 (N_1530,In_753,In_316);
nand U1531 (N_1531,In_592,In_677);
nor U1532 (N_1532,In_404,In_110);
and U1533 (N_1533,In_891,In_364);
and U1534 (N_1534,In_739,In_0);
and U1535 (N_1535,In_532,In_470);
nor U1536 (N_1536,In_890,In_943);
nand U1537 (N_1537,In_281,In_474);
or U1538 (N_1538,In_903,In_75);
nand U1539 (N_1539,In_987,In_290);
nand U1540 (N_1540,In_700,In_618);
and U1541 (N_1541,In_567,In_128);
or U1542 (N_1542,In_705,In_361);
nand U1543 (N_1543,In_962,In_924);
or U1544 (N_1544,In_574,In_70);
and U1545 (N_1545,In_866,In_374);
nand U1546 (N_1546,In_397,In_541);
nand U1547 (N_1547,In_128,In_97);
nand U1548 (N_1548,In_151,In_589);
nor U1549 (N_1549,In_256,In_798);
nor U1550 (N_1550,In_39,In_467);
and U1551 (N_1551,In_704,In_469);
nand U1552 (N_1552,In_996,In_225);
xor U1553 (N_1553,In_670,In_898);
or U1554 (N_1554,In_489,In_207);
nor U1555 (N_1555,In_451,In_158);
and U1556 (N_1556,In_813,In_911);
and U1557 (N_1557,In_634,In_877);
and U1558 (N_1558,In_793,In_654);
nand U1559 (N_1559,In_125,In_355);
or U1560 (N_1560,In_764,In_966);
and U1561 (N_1561,In_878,In_870);
or U1562 (N_1562,In_980,In_66);
nand U1563 (N_1563,In_397,In_557);
and U1564 (N_1564,In_116,In_534);
nand U1565 (N_1565,In_708,In_213);
or U1566 (N_1566,In_768,In_761);
or U1567 (N_1567,In_319,In_156);
and U1568 (N_1568,In_465,In_955);
or U1569 (N_1569,In_399,In_133);
xor U1570 (N_1570,In_150,In_96);
or U1571 (N_1571,In_803,In_894);
and U1572 (N_1572,In_555,In_614);
nor U1573 (N_1573,In_754,In_694);
nand U1574 (N_1574,In_732,In_849);
xnor U1575 (N_1575,In_822,In_496);
nand U1576 (N_1576,In_946,In_914);
nand U1577 (N_1577,In_809,In_763);
nor U1578 (N_1578,In_407,In_861);
xnor U1579 (N_1579,In_440,In_233);
and U1580 (N_1580,In_521,In_340);
and U1581 (N_1581,In_757,In_840);
or U1582 (N_1582,In_539,In_430);
or U1583 (N_1583,In_418,In_824);
or U1584 (N_1584,In_20,In_922);
and U1585 (N_1585,In_395,In_505);
nand U1586 (N_1586,In_219,In_349);
xor U1587 (N_1587,In_784,In_127);
nand U1588 (N_1588,In_820,In_567);
and U1589 (N_1589,In_828,In_924);
or U1590 (N_1590,In_218,In_653);
and U1591 (N_1591,In_431,In_192);
and U1592 (N_1592,In_507,In_972);
nor U1593 (N_1593,In_354,In_514);
nand U1594 (N_1594,In_157,In_64);
and U1595 (N_1595,In_262,In_578);
or U1596 (N_1596,In_506,In_702);
nor U1597 (N_1597,In_757,In_92);
nor U1598 (N_1598,In_421,In_138);
and U1599 (N_1599,In_142,In_674);
nor U1600 (N_1600,In_250,In_137);
or U1601 (N_1601,In_380,In_948);
and U1602 (N_1602,In_327,In_942);
or U1603 (N_1603,In_499,In_346);
xor U1604 (N_1604,In_614,In_668);
and U1605 (N_1605,In_511,In_438);
nand U1606 (N_1606,In_374,In_735);
nand U1607 (N_1607,In_408,In_579);
and U1608 (N_1608,In_612,In_392);
nand U1609 (N_1609,In_956,In_999);
or U1610 (N_1610,In_149,In_260);
and U1611 (N_1611,In_473,In_412);
nand U1612 (N_1612,In_538,In_67);
and U1613 (N_1613,In_683,In_830);
or U1614 (N_1614,In_375,In_954);
nor U1615 (N_1615,In_902,In_813);
or U1616 (N_1616,In_744,In_925);
and U1617 (N_1617,In_574,In_786);
and U1618 (N_1618,In_886,In_825);
or U1619 (N_1619,In_471,In_937);
or U1620 (N_1620,In_269,In_376);
or U1621 (N_1621,In_714,In_752);
and U1622 (N_1622,In_788,In_577);
and U1623 (N_1623,In_902,In_82);
nand U1624 (N_1624,In_458,In_37);
and U1625 (N_1625,In_833,In_353);
nor U1626 (N_1626,In_516,In_362);
xnor U1627 (N_1627,In_172,In_745);
nor U1628 (N_1628,In_93,In_345);
nand U1629 (N_1629,In_298,In_909);
and U1630 (N_1630,In_478,In_135);
nand U1631 (N_1631,In_318,In_47);
nand U1632 (N_1632,In_754,In_222);
nand U1633 (N_1633,In_3,In_486);
nand U1634 (N_1634,In_919,In_51);
nand U1635 (N_1635,In_788,In_256);
nand U1636 (N_1636,In_507,In_394);
nand U1637 (N_1637,In_387,In_653);
nand U1638 (N_1638,In_67,In_886);
and U1639 (N_1639,In_495,In_169);
or U1640 (N_1640,In_654,In_605);
nand U1641 (N_1641,In_475,In_351);
or U1642 (N_1642,In_437,In_632);
or U1643 (N_1643,In_447,In_984);
or U1644 (N_1644,In_675,In_236);
nand U1645 (N_1645,In_21,In_843);
xnor U1646 (N_1646,In_916,In_829);
or U1647 (N_1647,In_766,In_263);
nor U1648 (N_1648,In_425,In_183);
nand U1649 (N_1649,In_316,In_314);
nand U1650 (N_1650,In_219,In_348);
or U1651 (N_1651,In_91,In_822);
and U1652 (N_1652,In_826,In_442);
nand U1653 (N_1653,In_123,In_842);
or U1654 (N_1654,In_576,In_813);
nand U1655 (N_1655,In_609,In_360);
and U1656 (N_1656,In_636,In_921);
or U1657 (N_1657,In_490,In_219);
or U1658 (N_1658,In_573,In_640);
nand U1659 (N_1659,In_865,In_151);
nor U1660 (N_1660,In_972,In_824);
xnor U1661 (N_1661,In_666,In_151);
nand U1662 (N_1662,In_926,In_936);
nor U1663 (N_1663,In_105,In_162);
nand U1664 (N_1664,In_208,In_919);
nand U1665 (N_1665,In_620,In_825);
nand U1666 (N_1666,In_26,In_447);
nor U1667 (N_1667,In_554,In_461);
or U1668 (N_1668,In_716,In_834);
nor U1669 (N_1669,In_385,In_370);
xor U1670 (N_1670,In_406,In_503);
or U1671 (N_1671,In_8,In_448);
nor U1672 (N_1672,In_584,In_45);
nand U1673 (N_1673,In_579,In_961);
and U1674 (N_1674,In_39,In_54);
nor U1675 (N_1675,In_556,In_268);
and U1676 (N_1676,In_977,In_336);
nand U1677 (N_1677,In_227,In_932);
nand U1678 (N_1678,In_346,In_190);
nand U1679 (N_1679,In_422,In_973);
nor U1680 (N_1680,In_485,In_121);
nor U1681 (N_1681,In_280,In_507);
and U1682 (N_1682,In_839,In_398);
nor U1683 (N_1683,In_703,In_274);
nor U1684 (N_1684,In_472,In_502);
or U1685 (N_1685,In_278,In_260);
and U1686 (N_1686,In_347,In_128);
and U1687 (N_1687,In_198,In_133);
or U1688 (N_1688,In_171,In_501);
or U1689 (N_1689,In_582,In_600);
nand U1690 (N_1690,In_82,In_939);
nand U1691 (N_1691,In_436,In_470);
and U1692 (N_1692,In_313,In_773);
or U1693 (N_1693,In_162,In_326);
nor U1694 (N_1694,In_810,In_67);
xnor U1695 (N_1695,In_141,In_885);
nand U1696 (N_1696,In_295,In_672);
or U1697 (N_1697,In_99,In_379);
nand U1698 (N_1698,In_123,In_326);
nor U1699 (N_1699,In_901,In_716);
and U1700 (N_1700,In_987,In_876);
or U1701 (N_1701,In_927,In_549);
nand U1702 (N_1702,In_616,In_761);
nand U1703 (N_1703,In_206,In_253);
xnor U1704 (N_1704,In_446,In_263);
or U1705 (N_1705,In_103,In_900);
or U1706 (N_1706,In_865,In_836);
or U1707 (N_1707,In_280,In_692);
or U1708 (N_1708,In_801,In_413);
or U1709 (N_1709,In_50,In_355);
or U1710 (N_1710,In_334,In_431);
and U1711 (N_1711,In_413,In_262);
and U1712 (N_1712,In_427,In_828);
nand U1713 (N_1713,In_89,In_321);
xnor U1714 (N_1714,In_948,In_659);
nor U1715 (N_1715,In_447,In_126);
nand U1716 (N_1716,In_448,In_461);
xor U1717 (N_1717,In_312,In_687);
xnor U1718 (N_1718,In_887,In_874);
nand U1719 (N_1719,In_692,In_203);
or U1720 (N_1720,In_170,In_378);
nor U1721 (N_1721,In_196,In_570);
xor U1722 (N_1722,In_810,In_400);
or U1723 (N_1723,In_847,In_569);
or U1724 (N_1724,In_548,In_44);
nor U1725 (N_1725,In_602,In_190);
nand U1726 (N_1726,In_165,In_898);
or U1727 (N_1727,In_794,In_765);
xor U1728 (N_1728,In_826,In_675);
xor U1729 (N_1729,In_208,In_661);
nand U1730 (N_1730,In_899,In_623);
and U1731 (N_1731,In_95,In_487);
or U1732 (N_1732,In_837,In_508);
nor U1733 (N_1733,In_508,In_149);
or U1734 (N_1734,In_610,In_605);
nor U1735 (N_1735,In_508,In_48);
xnor U1736 (N_1736,In_457,In_878);
nand U1737 (N_1737,In_241,In_991);
nor U1738 (N_1738,In_262,In_907);
and U1739 (N_1739,In_579,In_418);
or U1740 (N_1740,In_823,In_233);
and U1741 (N_1741,In_27,In_627);
and U1742 (N_1742,In_624,In_521);
and U1743 (N_1743,In_910,In_914);
nor U1744 (N_1744,In_609,In_430);
nor U1745 (N_1745,In_95,In_106);
xor U1746 (N_1746,In_269,In_403);
and U1747 (N_1747,In_100,In_781);
nand U1748 (N_1748,In_566,In_772);
nand U1749 (N_1749,In_322,In_449);
or U1750 (N_1750,In_386,In_299);
nor U1751 (N_1751,In_925,In_383);
xor U1752 (N_1752,In_173,In_869);
and U1753 (N_1753,In_624,In_491);
nand U1754 (N_1754,In_275,In_977);
nor U1755 (N_1755,In_155,In_904);
and U1756 (N_1756,In_542,In_630);
nand U1757 (N_1757,In_16,In_133);
xnor U1758 (N_1758,In_122,In_778);
or U1759 (N_1759,In_834,In_346);
nor U1760 (N_1760,In_652,In_846);
nand U1761 (N_1761,In_842,In_697);
nor U1762 (N_1762,In_204,In_900);
and U1763 (N_1763,In_925,In_900);
or U1764 (N_1764,In_330,In_270);
xnor U1765 (N_1765,In_850,In_650);
nor U1766 (N_1766,In_239,In_461);
and U1767 (N_1767,In_406,In_431);
nor U1768 (N_1768,In_480,In_822);
nor U1769 (N_1769,In_745,In_382);
xor U1770 (N_1770,In_231,In_979);
xor U1771 (N_1771,In_89,In_471);
and U1772 (N_1772,In_991,In_324);
or U1773 (N_1773,In_228,In_537);
xnor U1774 (N_1774,In_609,In_254);
nor U1775 (N_1775,In_104,In_819);
nor U1776 (N_1776,In_822,In_64);
nor U1777 (N_1777,In_25,In_2);
and U1778 (N_1778,In_257,In_209);
nor U1779 (N_1779,In_364,In_114);
nor U1780 (N_1780,In_113,In_805);
nor U1781 (N_1781,In_769,In_471);
or U1782 (N_1782,In_172,In_493);
or U1783 (N_1783,In_568,In_804);
and U1784 (N_1784,In_101,In_593);
nand U1785 (N_1785,In_594,In_513);
or U1786 (N_1786,In_328,In_961);
or U1787 (N_1787,In_766,In_884);
nand U1788 (N_1788,In_909,In_150);
nor U1789 (N_1789,In_927,In_396);
and U1790 (N_1790,In_161,In_563);
nand U1791 (N_1791,In_178,In_738);
nand U1792 (N_1792,In_618,In_953);
nand U1793 (N_1793,In_814,In_820);
nor U1794 (N_1794,In_194,In_966);
nand U1795 (N_1795,In_33,In_554);
and U1796 (N_1796,In_852,In_230);
xnor U1797 (N_1797,In_293,In_649);
xnor U1798 (N_1798,In_54,In_205);
and U1799 (N_1799,In_696,In_326);
and U1800 (N_1800,In_521,In_993);
and U1801 (N_1801,In_832,In_300);
nor U1802 (N_1802,In_715,In_780);
or U1803 (N_1803,In_153,In_844);
nor U1804 (N_1804,In_655,In_204);
nor U1805 (N_1805,In_242,In_725);
nor U1806 (N_1806,In_496,In_786);
nor U1807 (N_1807,In_599,In_593);
xor U1808 (N_1808,In_696,In_889);
nor U1809 (N_1809,In_445,In_35);
and U1810 (N_1810,In_921,In_931);
nor U1811 (N_1811,In_226,In_330);
or U1812 (N_1812,In_755,In_826);
or U1813 (N_1813,In_871,In_395);
or U1814 (N_1814,In_75,In_864);
nor U1815 (N_1815,In_296,In_103);
xnor U1816 (N_1816,In_22,In_689);
nand U1817 (N_1817,In_847,In_790);
and U1818 (N_1818,In_849,In_593);
nor U1819 (N_1819,In_950,In_218);
or U1820 (N_1820,In_117,In_373);
nor U1821 (N_1821,In_478,In_106);
and U1822 (N_1822,In_418,In_776);
or U1823 (N_1823,In_170,In_65);
xnor U1824 (N_1824,In_858,In_184);
or U1825 (N_1825,In_765,In_792);
nand U1826 (N_1826,In_137,In_398);
and U1827 (N_1827,In_300,In_802);
nand U1828 (N_1828,In_192,In_569);
nor U1829 (N_1829,In_156,In_25);
or U1830 (N_1830,In_719,In_396);
nand U1831 (N_1831,In_853,In_367);
nand U1832 (N_1832,In_532,In_324);
or U1833 (N_1833,In_563,In_637);
xor U1834 (N_1834,In_612,In_720);
xor U1835 (N_1835,In_638,In_105);
and U1836 (N_1836,In_194,In_856);
nor U1837 (N_1837,In_666,In_425);
xor U1838 (N_1838,In_773,In_910);
or U1839 (N_1839,In_900,In_579);
and U1840 (N_1840,In_127,In_212);
and U1841 (N_1841,In_488,In_281);
and U1842 (N_1842,In_79,In_52);
nand U1843 (N_1843,In_577,In_638);
nor U1844 (N_1844,In_55,In_751);
nor U1845 (N_1845,In_112,In_287);
xor U1846 (N_1846,In_492,In_147);
nand U1847 (N_1847,In_347,In_863);
or U1848 (N_1848,In_751,In_394);
nor U1849 (N_1849,In_940,In_30);
nor U1850 (N_1850,In_274,In_33);
and U1851 (N_1851,In_247,In_502);
or U1852 (N_1852,In_610,In_560);
and U1853 (N_1853,In_578,In_115);
and U1854 (N_1854,In_169,In_809);
nor U1855 (N_1855,In_632,In_826);
and U1856 (N_1856,In_497,In_185);
nor U1857 (N_1857,In_666,In_300);
nand U1858 (N_1858,In_371,In_772);
nand U1859 (N_1859,In_608,In_987);
nor U1860 (N_1860,In_41,In_964);
xor U1861 (N_1861,In_812,In_287);
nor U1862 (N_1862,In_103,In_49);
or U1863 (N_1863,In_441,In_471);
nand U1864 (N_1864,In_496,In_585);
xnor U1865 (N_1865,In_356,In_577);
nor U1866 (N_1866,In_783,In_901);
nand U1867 (N_1867,In_188,In_520);
nor U1868 (N_1868,In_773,In_908);
and U1869 (N_1869,In_412,In_287);
nor U1870 (N_1870,In_676,In_710);
nor U1871 (N_1871,In_676,In_562);
nand U1872 (N_1872,In_483,In_855);
and U1873 (N_1873,In_104,In_537);
xnor U1874 (N_1874,In_380,In_398);
or U1875 (N_1875,In_682,In_291);
nor U1876 (N_1876,In_712,In_311);
and U1877 (N_1877,In_327,In_819);
nor U1878 (N_1878,In_103,In_911);
and U1879 (N_1879,In_860,In_408);
xnor U1880 (N_1880,In_337,In_303);
nor U1881 (N_1881,In_134,In_983);
or U1882 (N_1882,In_406,In_992);
or U1883 (N_1883,In_262,In_506);
and U1884 (N_1884,In_914,In_385);
nand U1885 (N_1885,In_308,In_93);
and U1886 (N_1886,In_290,In_80);
xor U1887 (N_1887,In_767,In_36);
or U1888 (N_1888,In_117,In_392);
and U1889 (N_1889,In_384,In_421);
nand U1890 (N_1890,In_523,In_313);
or U1891 (N_1891,In_815,In_309);
xor U1892 (N_1892,In_186,In_921);
nor U1893 (N_1893,In_280,In_604);
nor U1894 (N_1894,In_425,In_490);
nor U1895 (N_1895,In_228,In_299);
or U1896 (N_1896,In_951,In_13);
xor U1897 (N_1897,In_626,In_189);
and U1898 (N_1898,In_118,In_530);
and U1899 (N_1899,In_771,In_650);
nand U1900 (N_1900,In_559,In_683);
xor U1901 (N_1901,In_142,In_499);
nand U1902 (N_1902,In_475,In_882);
nor U1903 (N_1903,In_195,In_68);
nand U1904 (N_1904,In_138,In_993);
and U1905 (N_1905,In_636,In_811);
and U1906 (N_1906,In_151,In_693);
xnor U1907 (N_1907,In_523,In_333);
nand U1908 (N_1908,In_97,In_365);
and U1909 (N_1909,In_889,In_171);
and U1910 (N_1910,In_398,In_770);
nand U1911 (N_1911,In_438,In_319);
and U1912 (N_1912,In_930,In_253);
and U1913 (N_1913,In_632,In_474);
xor U1914 (N_1914,In_291,In_599);
or U1915 (N_1915,In_698,In_331);
nand U1916 (N_1916,In_378,In_656);
or U1917 (N_1917,In_275,In_584);
or U1918 (N_1918,In_154,In_176);
nand U1919 (N_1919,In_239,In_463);
nand U1920 (N_1920,In_14,In_285);
and U1921 (N_1921,In_941,In_370);
xnor U1922 (N_1922,In_233,In_169);
or U1923 (N_1923,In_54,In_514);
nor U1924 (N_1924,In_95,In_731);
or U1925 (N_1925,In_292,In_92);
xor U1926 (N_1926,In_205,In_572);
and U1927 (N_1927,In_265,In_50);
nand U1928 (N_1928,In_231,In_467);
nor U1929 (N_1929,In_374,In_222);
or U1930 (N_1930,In_154,In_953);
nor U1931 (N_1931,In_432,In_283);
nor U1932 (N_1932,In_500,In_587);
nor U1933 (N_1933,In_361,In_49);
or U1934 (N_1934,In_803,In_886);
nor U1935 (N_1935,In_172,In_914);
and U1936 (N_1936,In_3,In_608);
or U1937 (N_1937,In_445,In_926);
or U1938 (N_1938,In_303,In_928);
xor U1939 (N_1939,In_960,In_277);
or U1940 (N_1940,In_516,In_657);
and U1941 (N_1941,In_31,In_60);
xnor U1942 (N_1942,In_217,In_63);
nor U1943 (N_1943,In_88,In_706);
and U1944 (N_1944,In_926,In_188);
or U1945 (N_1945,In_960,In_329);
nand U1946 (N_1946,In_618,In_929);
nand U1947 (N_1947,In_157,In_382);
nor U1948 (N_1948,In_265,In_261);
nand U1949 (N_1949,In_355,In_503);
or U1950 (N_1950,In_914,In_912);
nand U1951 (N_1951,In_432,In_530);
nand U1952 (N_1952,In_880,In_615);
nor U1953 (N_1953,In_829,In_981);
and U1954 (N_1954,In_991,In_239);
nor U1955 (N_1955,In_891,In_256);
nor U1956 (N_1956,In_786,In_140);
nand U1957 (N_1957,In_139,In_177);
or U1958 (N_1958,In_621,In_230);
nand U1959 (N_1959,In_318,In_237);
nand U1960 (N_1960,In_732,In_367);
xor U1961 (N_1961,In_349,In_965);
or U1962 (N_1962,In_336,In_758);
and U1963 (N_1963,In_370,In_64);
and U1964 (N_1964,In_731,In_282);
nand U1965 (N_1965,In_686,In_993);
nand U1966 (N_1966,In_643,In_753);
nand U1967 (N_1967,In_314,In_897);
and U1968 (N_1968,In_146,In_117);
nor U1969 (N_1969,In_946,In_262);
or U1970 (N_1970,In_63,In_587);
xor U1971 (N_1971,In_815,In_919);
and U1972 (N_1972,In_194,In_982);
xnor U1973 (N_1973,In_275,In_71);
xor U1974 (N_1974,In_913,In_899);
and U1975 (N_1975,In_714,In_147);
or U1976 (N_1976,In_452,In_670);
nand U1977 (N_1977,In_962,In_964);
nor U1978 (N_1978,In_550,In_288);
nand U1979 (N_1979,In_119,In_352);
and U1980 (N_1980,In_717,In_874);
or U1981 (N_1981,In_552,In_533);
and U1982 (N_1982,In_892,In_829);
or U1983 (N_1983,In_932,In_58);
nand U1984 (N_1984,In_716,In_373);
xor U1985 (N_1985,In_886,In_144);
nor U1986 (N_1986,In_377,In_971);
and U1987 (N_1987,In_492,In_25);
xor U1988 (N_1988,In_706,In_572);
nand U1989 (N_1989,In_683,In_733);
nand U1990 (N_1990,In_851,In_256);
nand U1991 (N_1991,In_618,In_556);
nor U1992 (N_1992,In_965,In_651);
and U1993 (N_1993,In_629,In_618);
or U1994 (N_1994,In_670,In_528);
nand U1995 (N_1995,In_326,In_749);
nand U1996 (N_1996,In_107,In_805);
nor U1997 (N_1997,In_593,In_33);
nand U1998 (N_1998,In_973,In_834);
xnor U1999 (N_1999,In_525,In_520);
xor U2000 (N_2000,In_90,In_957);
and U2001 (N_2001,In_253,In_212);
xor U2002 (N_2002,In_658,In_224);
xnor U2003 (N_2003,In_712,In_121);
and U2004 (N_2004,In_652,In_952);
nand U2005 (N_2005,In_570,In_63);
or U2006 (N_2006,In_10,In_254);
nor U2007 (N_2007,In_106,In_776);
and U2008 (N_2008,In_984,In_241);
nand U2009 (N_2009,In_629,In_709);
nor U2010 (N_2010,In_543,In_126);
xnor U2011 (N_2011,In_227,In_221);
or U2012 (N_2012,In_100,In_357);
nand U2013 (N_2013,In_69,In_711);
nor U2014 (N_2014,In_148,In_246);
nor U2015 (N_2015,In_786,In_429);
xor U2016 (N_2016,In_138,In_956);
xor U2017 (N_2017,In_725,In_848);
nand U2018 (N_2018,In_160,In_404);
and U2019 (N_2019,In_299,In_866);
nand U2020 (N_2020,In_51,In_520);
or U2021 (N_2021,In_816,In_221);
or U2022 (N_2022,In_201,In_488);
or U2023 (N_2023,In_540,In_410);
nor U2024 (N_2024,In_722,In_879);
xor U2025 (N_2025,In_884,In_444);
and U2026 (N_2026,In_756,In_879);
and U2027 (N_2027,In_619,In_905);
xor U2028 (N_2028,In_630,In_460);
nor U2029 (N_2029,In_198,In_328);
and U2030 (N_2030,In_356,In_265);
and U2031 (N_2031,In_403,In_227);
nand U2032 (N_2032,In_997,In_123);
or U2033 (N_2033,In_608,In_731);
and U2034 (N_2034,In_132,In_367);
or U2035 (N_2035,In_430,In_471);
nor U2036 (N_2036,In_183,In_100);
nor U2037 (N_2037,In_114,In_639);
nand U2038 (N_2038,In_920,In_407);
and U2039 (N_2039,In_952,In_743);
xnor U2040 (N_2040,In_472,In_111);
nand U2041 (N_2041,In_436,In_125);
and U2042 (N_2042,In_349,In_9);
xnor U2043 (N_2043,In_426,In_179);
nand U2044 (N_2044,In_174,In_417);
xor U2045 (N_2045,In_268,In_616);
nor U2046 (N_2046,In_789,In_111);
nand U2047 (N_2047,In_153,In_828);
or U2048 (N_2048,In_186,In_765);
nand U2049 (N_2049,In_934,In_176);
nand U2050 (N_2050,In_554,In_305);
and U2051 (N_2051,In_74,In_79);
and U2052 (N_2052,In_536,In_555);
or U2053 (N_2053,In_270,In_414);
and U2054 (N_2054,In_329,In_410);
and U2055 (N_2055,In_359,In_657);
and U2056 (N_2056,In_961,In_900);
nand U2057 (N_2057,In_752,In_905);
and U2058 (N_2058,In_716,In_506);
nor U2059 (N_2059,In_154,In_394);
nand U2060 (N_2060,In_160,In_313);
and U2061 (N_2061,In_118,In_970);
or U2062 (N_2062,In_468,In_27);
nor U2063 (N_2063,In_913,In_6);
and U2064 (N_2064,In_448,In_349);
nand U2065 (N_2065,In_874,In_871);
nand U2066 (N_2066,In_160,In_895);
or U2067 (N_2067,In_878,In_199);
or U2068 (N_2068,In_107,In_634);
and U2069 (N_2069,In_625,In_208);
nand U2070 (N_2070,In_740,In_845);
and U2071 (N_2071,In_171,In_629);
and U2072 (N_2072,In_438,In_623);
nor U2073 (N_2073,In_1,In_639);
and U2074 (N_2074,In_249,In_820);
nand U2075 (N_2075,In_819,In_575);
nand U2076 (N_2076,In_614,In_204);
or U2077 (N_2077,In_956,In_273);
and U2078 (N_2078,In_869,In_340);
nor U2079 (N_2079,In_96,In_385);
and U2080 (N_2080,In_239,In_300);
or U2081 (N_2081,In_541,In_133);
xnor U2082 (N_2082,In_986,In_842);
and U2083 (N_2083,In_78,In_875);
and U2084 (N_2084,In_307,In_116);
and U2085 (N_2085,In_607,In_145);
or U2086 (N_2086,In_518,In_66);
nor U2087 (N_2087,In_150,In_420);
xnor U2088 (N_2088,In_591,In_114);
or U2089 (N_2089,In_22,In_190);
nor U2090 (N_2090,In_161,In_27);
or U2091 (N_2091,In_510,In_503);
nor U2092 (N_2092,In_896,In_69);
or U2093 (N_2093,In_728,In_913);
nor U2094 (N_2094,In_609,In_718);
and U2095 (N_2095,In_189,In_680);
nand U2096 (N_2096,In_991,In_145);
and U2097 (N_2097,In_285,In_902);
nand U2098 (N_2098,In_835,In_59);
and U2099 (N_2099,In_357,In_724);
nand U2100 (N_2100,In_622,In_38);
and U2101 (N_2101,In_785,In_281);
or U2102 (N_2102,In_313,In_781);
nand U2103 (N_2103,In_945,In_691);
xnor U2104 (N_2104,In_919,In_565);
nand U2105 (N_2105,In_119,In_139);
nand U2106 (N_2106,In_543,In_242);
nand U2107 (N_2107,In_741,In_456);
and U2108 (N_2108,In_361,In_636);
or U2109 (N_2109,In_710,In_800);
nor U2110 (N_2110,In_866,In_816);
nor U2111 (N_2111,In_429,In_20);
and U2112 (N_2112,In_757,In_451);
and U2113 (N_2113,In_374,In_871);
nand U2114 (N_2114,In_814,In_323);
and U2115 (N_2115,In_887,In_305);
and U2116 (N_2116,In_989,In_5);
xor U2117 (N_2117,In_915,In_551);
or U2118 (N_2118,In_728,In_951);
nand U2119 (N_2119,In_766,In_186);
nor U2120 (N_2120,In_968,In_611);
and U2121 (N_2121,In_539,In_523);
nand U2122 (N_2122,In_430,In_716);
and U2123 (N_2123,In_85,In_770);
or U2124 (N_2124,In_734,In_300);
nor U2125 (N_2125,In_182,In_365);
nor U2126 (N_2126,In_374,In_16);
xnor U2127 (N_2127,In_595,In_633);
and U2128 (N_2128,In_601,In_146);
and U2129 (N_2129,In_509,In_728);
nand U2130 (N_2130,In_640,In_365);
xor U2131 (N_2131,In_609,In_114);
nor U2132 (N_2132,In_939,In_121);
nor U2133 (N_2133,In_155,In_304);
nand U2134 (N_2134,In_395,In_345);
xnor U2135 (N_2135,In_511,In_680);
nand U2136 (N_2136,In_822,In_588);
or U2137 (N_2137,In_98,In_365);
xnor U2138 (N_2138,In_883,In_1);
nor U2139 (N_2139,In_295,In_456);
xnor U2140 (N_2140,In_227,In_611);
and U2141 (N_2141,In_88,In_477);
xnor U2142 (N_2142,In_779,In_605);
and U2143 (N_2143,In_387,In_218);
and U2144 (N_2144,In_241,In_333);
and U2145 (N_2145,In_645,In_74);
or U2146 (N_2146,In_810,In_679);
or U2147 (N_2147,In_453,In_840);
and U2148 (N_2148,In_343,In_15);
nand U2149 (N_2149,In_486,In_433);
or U2150 (N_2150,In_258,In_727);
and U2151 (N_2151,In_938,In_398);
nor U2152 (N_2152,In_963,In_258);
and U2153 (N_2153,In_810,In_175);
and U2154 (N_2154,In_897,In_325);
or U2155 (N_2155,In_454,In_648);
nor U2156 (N_2156,In_456,In_617);
or U2157 (N_2157,In_422,In_758);
nand U2158 (N_2158,In_861,In_146);
and U2159 (N_2159,In_19,In_604);
and U2160 (N_2160,In_338,In_281);
and U2161 (N_2161,In_15,In_405);
xnor U2162 (N_2162,In_278,In_546);
nand U2163 (N_2163,In_38,In_998);
nor U2164 (N_2164,In_181,In_810);
or U2165 (N_2165,In_928,In_989);
xor U2166 (N_2166,In_372,In_448);
and U2167 (N_2167,In_628,In_697);
nor U2168 (N_2168,In_284,In_81);
nor U2169 (N_2169,In_163,In_791);
xnor U2170 (N_2170,In_380,In_892);
or U2171 (N_2171,In_708,In_474);
or U2172 (N_2172,In_130,In_878);
nand U2173 (N_2173,In_207,In_695);
and U2174 (N_2174,In_770,In_832);
nor U2175 (N_2175,In_814,In_341);
or U2176 (N_2176,In_326,In_949);
or U2177 (N_2177,In_658,In_349);
and U2178 (N_2178,In_878,In_623);
and U2179 (N_2179,In_404,In_941);
or U2180 (N_2180,In_709,In_311);
or U2181 (N_2181,In_558,In_397);
nand U2182 (N_2182,In_687,In_529);
or U2183 (N_2183,In_522,In_775);
nor U2184 (N_2184,In_195,In_751);
xor U2185 (N_2185,In_139,In_822);
xor U2186 (N_2186,In_254,In_374);
or U2187 (N_2187,In_992,In_402);
nor U2188 (N_2188,In_81,In_767);
and U2189 (N_2189,In_580,In_725);
and U2190 (N_2190,In_31,In_511);
and U2191 (N_2191,In_810,In_518);
or U2192 (N_2192,In_209,In_289);
xnor U2193 (N_2193,In_953,In_599);
xor U2194 (N_2194,In_408,In_628);
and U2195 (N_2195,In_401,In_345);
or U2196 (N_2196,In_930,In_262);
or U2197 (N_2197,In_252,In_189);
nand U2198 (N_2198,In_615,In_519);
and U2199 (N_2199,In_343,In_636);
or U2200 (N_2200,In_367,In_325);
or U2201 (N_2201,In_306,In_746);
nand U2202 (N_2202,In_660,In_586);
nor U2203 (N_2203,In_269,In_119);
nor U2204 (N_2204,In_560,In_153);
nand U2205 (N_2205,In_991,In_644);
or U2206 (N_2206,In_619,In_41);
xor U2207 (N_2207,In_69,In_871);
xnor U2208 (N_2208,In_556,In_534);
xnor U2209 (N_2209,In_592,In_382);
nor U2210 (N_2210,In_167,In_697);
xnor U2211 (N_2211,In_290,In_154);
nor U2212 (N_2212,In_539,In_526);
and U2213 (N_2213,In_8,In_804);
or U2214 (N_2214,In_873,In_70);
and U2215 (N_2215,In_704,In_328);
and U2216 (N_2216,In_976,In_475);
nand U2217 (N_2217,In_72,In_400);
nand U2218 (N_2218,In_874,In_658);
xnor U2219 (N_2219,In_674,In_987);
nand U2220 (N_2220,In_48,In_350);
and U2221 (N_2221,In_71,In_217);
xnor U2222 (N_2222,In_900,In_403);
nor U2223 (N_2223,In_67,In_712);
xnor U2224 (N_2224,In_766,In_588);
and U2225 (N_2225,In_953,In_281);
and U2226 (N_2226,In_182,In_602);
nor U2227 (N_2227,In_489,In_723);
nor U2228 (N_2228,In_949,In_339);
and U2229 (N_2229,In_112,In_456);
nor U2230 (N_2230,In_500,In_919);
or U2231 (N_2231,In_387,In_597);
nor U2232 (N_2232,In_429,In_369);
and U2233 (N_2233,In_298,In_138);
nand U2234 (N_2234,In_213,In_977);
nor U2235 (N_2235,In_406,In_748);
nand U2236 (N_2236,In_588,In_620);
nand U2237 (N_2237,In_827,In_286);
nor U2238 (N_2238,In_766,In_240);
nor U2239 (N_2239,In_765,In_227);
nand U2240 (N_2240,In_926,In_860);
nor U2241 (N_2241,In_296,In_866);
or U2242 (N_2242,In_389,In_926);
or U2243 (N_2243,In_264,In_48);
nand U2244 (N_2244,In_142,In_578);
nand U2245 (N_2245,In_678,In_786);
nand U2246 (N_2246,In_555,In_52);
nor U2247 (N_2247,In_725,In_974);
and U2248 (N_2248,In_824,In_27);
or U2249 (N_2249,In_522,In_659);
or U2250 (N_2250,In_881,In_570);
nor U2251 (N_2251,In_296,In_978);
xor U2252 (N_2252,In_233,In_665);
nand U2253 (N_2253,In_816,In_780);
or U2254 (N_2254,In_359,In_52);
xnor U2255 (N_2255,In_818,In_684);
nand U2256 (N_2256,In_338,In_649);
or U2257 (N_2257,In_217,In_966);
nand U2258 (N_2258,In_190,In_154);
nor U2259 (N_2259,In_842,In_571);
nor U2260 (N_2260,In_318,In_845);
nor U2261 (N_2261,In_497,In_494);
and U2262 (N_2262,In_242,In_133);
nand U2263 (N_2263,In_625,In_282);
nor U2264 (N_2264,In_739,In_177);
nand U2265 (N_2265,In_638,In_804);
or U2266 (N_2266,In_228,In_344);
and U2267 (N_2267,In_564,In_2);
nand U2268 (N_2268,In_973,In_757);
xor U2269 (N_2269,In_608,In_286);
nor U2270 (N_2270,In_769,In_518);
or U2271 (N_2271,In_461,In_167);
or U2272 (N_2272,In_24,In_219);
nor U2273 (N_2273,In_284,In_947);
xor U2274 (N_2274,In_887,In_546);
and U2275 (N_2275,In_72,In_852);
nand U2276 (N_2276,In_62,In_238);
nand U2277 (N_2277,In_238,In_249);
or U2278 (N_2278,In_667,In_629);
xnor U2279 (N_2279,In_730,In_724);
nor U2280 (N_2280,In_770,In_732);
xor U2281 (N_2281,In_991,In_894);
or U2282 (N_2282,In_925,In_248);
nand U2283 (N_2283,In_222,In_919);
and U2284 (N_2284,In_961,In_155);
nand U2285 (N_2285,In_68,In_820);
xnor U2286 (N_2286,In_28,In_985);
or U2287 (N_2287,In_143,In_206);
and U2288 (N_2288,In_715,In_206);
or U2289 (N_2289,In_598,In_206);
nor U2290 (N_2290,In_712,In_320);
nor U2291 (N_2291,In_728,In_347);
nor U2292 (N_2292,In_717,In_949);
xor U2293 (N_2293,In_667,In_766);
nand U2294 (N_2294,In_521,In_747);
nor U2295 (N_2295,In_193,In_770);
or U2296 (N_2296,In_829,In_949);
or U2297 (N_2297,In_936,In_400);
nor U2298 (N_2298,In_152,In_794);
and U2299 (N_2299,In_34,In_279);
and U2300 (N_2300,In_63,In_371);
nand U2301 (N_2301,In_913,In_477);
and U2302 (N_2302,In_794,In_123);
and U2303 (N_2303,In_918,In_674);
and U2304 (N_2304,In_594,In_415);
nand U2305 (N_2305,In_662,In_35);
nand U2306 (N_2306,In_406,In_354);
or U2307 (N_2307,In_529,In_372);
nand U2308 (N_2308,In_85,In_3);
or U2309 (N_2309,In_264,In_518);
and U2310 (N_2310,In_370,In_932);
and U2311 (N_2311,In_695,In_771);
and U2312 (N_2312,In_66,In_53);
nor U2313 (N_2313,In_260,In_261);
nand U2314 (N_2314,In_775,In_898);
nand U2315 (N_2315,In_432,In_794);
xnor U2316 (N_2316,In_872,In_314);
or U2317 (N_2317,In_697,In_391);
nor U2318 (N_2318,In_537,In_850);
or U2319 (N_2319,In_402,In_244);
nor U2320 (N_2320,In_459,In_485);
xnor U2321 (N_2321,In_19,In_80);
nand U2322 (N_2322,In_156,In_273);
nand U2323 (N_2323,In_555,In_380);
nor U2324 (N_2324,In_489,In_452);
nor U2325 (N_2325,In_174,In_403);
nand U2326 (N_2326,In_282,In_429);
nand U2327 (N_2327,In_265,In_60);
or U2328 (N_2328,In_134,In_938);
xor U2329 (N_2329,In_520,In_619);
or U2330 (N_2330,In_436,In_825);
nor U2331 (N_2331,In_892,In_387);
nor U2332 (N_2332,In_64,In_900);
nand U2333 (N_2333,In_631,In_147);
nand U2334 (N_2334,In_630,In_832);
or U2335 (N_2335,In_990,In_397);
nor U2336 (N_2336,In_39,In_949);
and U2337 (N_2337,In_209,In_557);
and U2338 (N_2338,In_979,In_227);
or U2339 (N_2339,In_279,In_821);
nand U2340 (N_2340,In_746,In_826);
and U2341 (N_2341,In_382,In_375);
and U2342 (N_2342,In_482,In_541);
nor U2343 (N_2343,In_748,In_517);
and U2344 (N_2344,In_645,In_250);
nor U2345 (N_2345,In_860,In_685);
nand U2346 (N_2346,In_316,In_610);
nor U2347 (N_2347,In_777,In_236);
or U2348 (N_2348,In_690,In_56);
nor U2349 (N_2349,In_162,In_206);
and U2350 (N_2350,In_89,In_44);
nand U2351 (N_2351,In_997,In_933);
xnor U2352 (N_2352,In_98,In_58);
and U2353 (N_2353,In_190,In_326);
xnor U2354 (N_2354,In_767,In_637);
xnor U2355 (N_2355,In_53,In_147);
and U2356 (N_2356,In_835,In_70);
xnor U2357 (N_2357,In_495,In_344);
and U2358 (N_2358,In_993,In_914);
nor U2359 (N_2359,In_212,In_673);
nor U2360 (N_2360,In_386,In_272);
nor U2361 (N_2361,In_769,In_436);
or U2362 (N_2362,In_335,In_711);
nor U2363 (N_2363,In_628,In_382);
or U2364 (N_2364,In_807,In_142);
or U2365 (N_2365,In_825,In_951);
nand U2366 (N_2366,In_915,In_998);
or U2367 (N_2367,In_869,In_559);
and U2368 (N_2368,In_568,In_850);
nor U2369 (N_2369,In_541,In_339);
and U2370 (N_2370,In_465,In_542);
nor U2371 (N_2371,In_695,In_708);
and U2372 (N_2372,In_178,In_603);
nand U2373 (N_2373,In_949,In_396);
xnor U2374 (N_2374,In_757,In_419);
nor U2375 (N_2375,In_151,In_772);
nand U2376 (N_2376,In_945,In_317);
xor U2377 (N_2377,In_387,In_492);
nand U2378 (N_2378,In_420,In_377);
nand U2379 (N_2379,In_894,In_675);
nor U2380 (N_2380,In_288,In_793);
nand U2381 (N_2381,In_919,In_326);
or U2382 (N_2382,In_255,In_335);
nor U2383 (N_2383,In_706,In_38);
nor U2384 (N_2384,In_892,In_172);
or U2385 (N_2385,In_463,In_616);
xnor U2386 (N_2386,In_861,In_719);
or U2387 (N_2387,In_508,In_211);
and U2388 (N_2388,In_598,In_980);
or U2389 (N_2389,In_919,In_699);
xnor U2390 (N_2390,In_804,In_303);
nand U2391 (N_2391,In_390,In_671);
xor U2392 (N_2392,In_934,In_972);
nand U2393 (N_2393,In_317,In_75);
and U2394 (N_2394,In_268,In_463);
or U2395 (N_2395,In_300,In_814);
or U2396 (N_2396,In_103,In_977);
or U2397 (N_2397,In_699,In_704);
or U2398 (N_2398,In_716,In_860);
xor U2399 (N_2399,In_654,In_403);
and U2400 (N_2400,In_707,In_167);
nand U2401 (N_2401,In_686,In_35);
and U2402 (N_2402,In_282,In_712);
or U2403 (N_2403,In_663,In_936);
xor U2404 (N_2404,In_440,In_61);
or U2405 (N_2405,In_301,In_278);
and U2406 (N_2406,In_243,In_99);
nand U2407 (N_2407,In_922,In_348);
and U2408 (N_2408,In_559,In_388);
xnor U2409 (N_2409,In_331,In_729);
nor U2410 (N_2410,In_317,In_239);
xor U2411 (N_2411,In_996,In_816);
and U2412 (N_2412,In_783,In_360);
nor U2413 (N_2413,In_703,In_790);
or U2414 (N_2414,In_741,In_977);
or U2415 (N_2415,In_519,In_944);
nand U2416 (N_2416,In_394,In_124);
and U2417 (N_2417,In_294,In_261);
nor U2418 (N_2418,In_576,In_16);
nor U2419 (N_2419,In_356,In_140);
nor U2420 (N_2420,In_176,In_277);
and U2421 (N_2421,In_844,In_384);
nand U2422 (N_2422,In_403,In_590);
nand U2423 (N_2423,In_128,In_571);
and U2424 (N_2424,In_890,In_359);
nor U2425 (N_2425,In_528,In_808);
and U2426 (N_2426,In_570,In_358);
and U2427 (N_2427,In_948,In_957);
or U2428 (N_2428,In_194,In_461);
nand U2429 (N_2429,In_590,In_456);
or U2430 (N_2430,In_354,In_896);
or U2431 (N_2431,In_761,In_185);
nor U2432 (N_2432,In_335,In_846);
and U2433 (N_2433,In_263,In_183);
and U2434 (N_2434,In_633,In_878);
nand U2435 (N_2435,In_70,In_56);
or U2436 (N_2436,In_693,In_764);
or U2437 (N_2437,In_103,In_77);
or U2438 (N_2438,In_963,In_804);
and U2439 (N_2439,In_190,In_508);
nor U2440 (N_2440,In_353,In_733);
nand U2441 (N_2441,In_449,In_833);
xor U2442 (N_2442,In_460,In_440);
nor U2443 (N_2443,In_736,In_34);
xnor U2444 (N_2444,In_566,In_796);
nand U2445 (N_2445,In_471,In_514);
and U2446 (N_2446,In_973,In_127);
or U2447 (N_2447,In_640,In_235);
nand U2448 (N_2448,In_52,In_783);
nand U2449 (N_2449,In_670,In_608);
and U2450 (N_2450,In_948,In_375);
or U2451 (N_2451,In_990,In_582);
and U2452 (N_2452,In_87,In_528);
nand U2453 (N_2453,In_77,In_740);
nand U2454 (N_2454,In_346,In_748);
nor U2455 (N_2455,In_79,In_76);
nand U2456 (N_2456,In_524,In_843);
or U2457 (N_2457,In_120,In_331);
and U2458 (N_2458,In_866,In_227);
nand U2459 (N_2459,In_628,In_483);
nor U2460 (N_2460,In_326,In_516);
nand U2461 (N_2461,In_110,In_762);
nand U2462 (N_2462,In_776,In_680);
nor U2463 (N_2463,In_594,In_522);
or U2464 (N_2464,In_966,In_422);
and U2465 (N_2465,In_346,In_246);
or U2466 (N_2466,In_191,In_1);
nand U2467 (N_2467,In_767,In_160);
nor U2468 (N_2468,In_799,In_457);
nand U2469 (N_2469,In_864,In_806);
nor U2470 (N_2470,In_766,In_832);
nor U2471 (N_2471,In_766,In_326);
nor U2472 (N_2472,In_918,In_407);
or U2473 (N_2473,In_612,In_238);
or U2474 (N_2474,In_802,In_107);
nor U2475 (N_2475,In_927,In_147);
and U2476 (N_2476,In_746,In_849);
nand U2477 (N_2477,In_481,In_878);
and U2478 (N_2478,In_280,In_431);
or U2479 (N_2479,In_862,In_455);
or U2480 (N_2480,In_480,In_172);
and U2481 (N_2481,In_965,In_229);
and U2482 (N_2482,In_711,In_332);
and U2483 (N_2483,In_208,In_238);
nor U2484 (N_2484,In_59,In_561);
or U2485 (N_2485,In_767,In_317);
or U2486 (N_2486,In_55,In_160);
and U2487 (N_2487,In_983,In_706);
nand U2488 (N_2488,In_75,In_754);
nor U2489 (N_2489,In_534,In_397);
nand U2490 (N_2490,In_384,In_120);
and U2491 (N_2491,In_520,In_578);
nand U2492 (N_2492,In_190,In_940);
nor U2493 (N_2493,In_254,In_516);
nand U2494 (N_2494,In_179,In_327);
nor U2495 (N_2495,In_600,In_928);
nand U2496 (N_2496,In_460,In_747);
nand U2497 (N_2497,In_106,In_395);
or U2498 (N_2498,In_10,In_563);
nand U2499 (N_2499,In_545,In_529);
nand U2500 (N_2500,N_1962,N_2284);
or U2501 (N_2501,N_2041,N_1993);
or U2502 (N_2502,N_702,N_659);
and U2503 (N_2503,N_312,N_822);
and U2504 (N_2504,N_1749,N_598);
nand U2505 (N_2505,N_43,N_1335);
xnor U2506 (N_2506,N_483,N_1442);
and U2507 (N_2507,N_70,N_678);
nand U2508 (N_2508,N_237,N_1847);
nor U2509 (N_2509,N_132,N_2055);
nand U2510 (N_2510,N_1271,N_1114);
and U2511 (N_2511,N_1493,N_75);
or U2512 (N_2512,N_665,N_161);
nand U2513 (N_2513,N_1126,N_464);
xnor U2514 (N_2514,N_2173,N_478);
xor U2515 (N_2515,N_1416,N_113);
and U2516 (N_2516,N_1183,N_1156);
and U2517 (N_2517,N_916,N_325);
or U2518 (N_2518,N_2171,N_1265);
nand U2519 (N_2519,N_1655,N_109);
nor U2520 (N_2520,N_418,N_1365);
nand U2521 (N_2521,N_2147,N_837);
nand U2522 (N_2522,N_842,N_502);
and U2523 (N_2523,N_1235,N_2403);
and U2524 (N_2524,N_972,N_1176);
nor U2525 (N_2525,N_2118,N_596);
nor U2526 (N_2526,N_376,N_891);
nor U2527 (N_2527,N_1476,N_744);
or U2528 (N_2528,N_2373,N_384);
or U2529 (N_2529,N_581,N_2050);
or U2530 (N_2530,N_2148,N_1836);
nor U2531 (N_2531,N_371,N_492);
or U2532 (N_2532,N_396,N_434);
and U2533 (N_2533,N_949,N_560);
and U2534 (N_2534,N_348,N_1578);
or U2535 (N_2535,N_305,N_1044);
nand U2536 (N_2536,N_441,N_353);
or U2537 (N_2537,N_2441,N_1141);
nand U2538 (N_2538,N_1826,N_1672);
nor U2539 (N_2539,N_2290,N_858);
or U2540 (N_2540,N_673,N_482);
or U2541 (N_2541,N_936,N_2064);
nor U2542 (N_2542,N_1394,N_76);
or U2543 (N_2543,N_2166,N_2392);
or U2544 (N_2544,N_701,N_760);
nor U2545 (N_2545,N_1827,N_68);
or U2546 (N_2546,N_2297,N_2233);
nand U2547 (N_2547,N_1653,N_1911);
nor U2548 (N_2548,N_2440,N_1157);
nand U2549 (N_2549,N_2389,N_1703);
nand U2550 (N_2550,N_2397,N_1293);
or U2551 (N_2551,N_1298,N_2030);
nand U2552 (N_2552,N_1279,N_92);
nor U2553 (N_2553,N_223,N_2028);
nor U2554 (N_2554,N_643,N_863);
and U2555 (N_2555,N_2438,N_2198);
and U2556 (N_2556,N_1031,N_1459);
nand U2557 (N_2557,N_1694,N_617);
or U2558 (N_2558,N_2323,N_1783);
or U2559 (N_2559,N_272,N_2033);
nand U2560 (N_2560,N_463,N_2398);
and U2561 (N_2561,N_1452,N_279);
or U2562 (N_2562,N_1479,N_1385);
xnor U2563 (N_2563,N_465,N_1172);
xnor U2564 (N_2564,N_1532,N_394);
nand U2565 (N_2565,N_77,N_933);
xor U2566 (N_2566,N_1419,N_895);
or U2567 (N_2567,N_939,N_1789);
nand U2568 (N_2568,N_715,N_439);
and U2569 (N_2569,N_1978,N_1399);
and U2570 (N_2570,N_606,N_1292);
nand U2571 (N_2571,N_74,N_423);
or U2572 (N_2572,N_1494,N_117);
or U2573 (N_2573,N_763,N_1460);
nand U2574 (N_2574,N_1805,N_2481);
xnor U2575 (N_2575,N_214,N_1546);
and U2576 (N_2576,N_513,N_183);
nand U2577 (N_2577,N_1750,N_1935);
and U2578 (N_2578,N_694,N_341);
nand U2579 (N_2579,N_1919,N_1237);
or U2580 (N_2580,N_1066,N_1926);
or U2581 (N_2581,N_998,N_1830);
or U2582 (N_2582,N_444,N_1143);
nor U2583 (N_2583,N_1297,N_1304);
nor U2584 (N_2584,N_1633,N_707);
and U2585 (N_2585,N_335,N_339);
and U2586 (N_2586,N_2218,N_892);
or U2587 (N_2587,N_1753,N_1153);
nand U2588 (N_2588,N_767,N_1545);
xor U2589 (N_2589,N_2220,N_1272);
nand U2590 (N_2590,N_125,N_968);
or U2591 (N_2591,N_170,N_2150);
nor U2592 (N_2592,N_2329,N_169);
or U2593 (N_2593,N_1051,N_1523);
nor U2594 (N_2594,N_53,N_1988);
or U2595 (N_2595,N_2486,N_1191);
and U2596 (N_2596,N_1357,N_1547);
or U2597 (N_2597,N_1923,N_81);
and U2598 (N_2598,N_752,N_738);
nor U2599 (N_2599,N_918,N_1280);
nand U2600 (N_2600,N_794,N_898);
nand U2601 (N_2601,N_664,N_594);
nand U2602 (N_2602,N_628,N_85);
xnor U2603 (N_2603,N_346,N_299);
or U2604 (N_2604,N_1027,N_2449);
nor U2605 (N_2605,N_593,N_1870);
nand U2606 (N_2606,N_605,N_804);
nand U2607 (N_2607,N_1517,N_386);
nand U2608 (N_2608,N_1282,N_2022);
and U2609 (N_2609,N_1039,N_2263);
or U2610 (N_2610,N_2360,N_369);
and U2611 (N_2611,N_682,N_407);
and U2612 (N_2612,N_2324,N_798);
nand U2613 (N_2613,N_1758,N_637);
nor U2614 (N_2614,N_1806,N_2090);
or U2615 (N_2615,N_1192,N_385);
nand U2616 (N_2616,N_978,N_654);
nor U2617 (N_2617,N_2453,N_2425);
and U2618 (N_2618,N_362,N_149);
and U2619 (N_2619,N_881,N_2145);
or U2620 (N_2620,N_83,N_2071);
or U2621 (N_2621,N_1884,N_1702);
nor U2622 (N_2622,N_1996,N_921);
and U2623 (N_2623,N_2303,N_818);
nand U2624 (N_2624,N_2488,N_2119);
nand U2625 (N_2625,N_160,N_1573);
nor U2626 (N_2626,N_1195,N_914);
nand U2627 (N_2627,N_2436,N_1595);
and U2628 (N_2628,N_449,N_90);
or U2629 (N_2629,N_1364,N_1409);
nand U2630 (N_2630,N_1150,N_2244);
nor U2631 (N_2631,N_505,N_1200);
nand U2632 (N_2632,N_34,N_189);
nand U2633 (N_2633,N_1255,N_995);
or U2634 (N_2634,N_2154,N_685);
and U2635 (N_2635,N_496,N_1437);
nor U2636 (N_2636,N_1418,N_994);
xor U2637 (N_2637,N_271,N_247);
or U2638 (N_2638,N_1915,N_719);
nor U2639 (N_2639,N_1128,N_1270);
nor U2640 (N_2640,N_336,N_996);
nand U2641 (N_2641,N_2428,N_1345);
and U2642 (N_2642,N_1554,N_2343);
nand U2643 (N_2643,N_352,N_535);
and U2644 (N_2644,N_1916,N_1893);
nor U2645 (N_2645,N_1859,N_1053);
nand U2646 (N_2646,N_1116,N_118);
xnor U2647 (N_2647,N_1047,N_656);
and U2648 (N_2648,N_2252,N_790);
xnor U2649 (N_2649,N_556,N_37);
or U2650 (N_2650,N_1086,N_1690);
and U2651 (N_2651,N_1036,N_2376);
nor U2652 (N_2652,N_1751,N_1107);
or U2653 (N_2653,N_1638,N_1226);
nand U2654 (N_2654,N_1092,N_1151);
or U2655 (N_2655,N_1930,N_350);
nor U2656 (N_2656,N_1186,N_2188);
or U2657 (N_2657,N_86,N_2142);
nand U2658 (N_2658,N_44,N_539);
and U2659 (N_2659,N_736,N_1995);
nor U2660 (N_2660,N_850,N_35);
nor U2661 (N_2661,N_2182,N_937);
or U2662 (N_2662,N_1076,N_140);
nand U2663 (N_2663,N_1012,N_1465);
xnor U2664 (N_2664,N_433,N_1225);
or U2665 (N_2665,N_2298,N_1468);
and U2666 (N_2666,N_1303,N_1987);
and U2667 (N_2667,N_1363,N_946);
and U2668 (N_2668,N_2306,N_1649);
xor U2669 (N_2669,N_1563,N_262);
and U2670 (N_2670,N_1008,N_1273);
nand U2671 (N_2671,N_1918,N_2085);
nor U2672 (N_2672,N_1743,N_1078);
nand U2673 (N_2673,N_1193,N_1770);
nand U2674 (N_2674,N_1097,N_40);
nor U2675 (N_2675,N_15,N_1056);
nor U2676 (N_2676,N_256,N_1887);
nor U2677 (N_2677,N_1982,N_2247);
nor U2678 (N_2678,N_1881,N_458);
nand U2679 (N_2679,N_1854,N_2065);
nor U2680 (N_2680,N_0,N_101);
nor U2681 (N_2681,N_2472,N_2045);
xnor U2682 (N_2682,N_1949,N_651);
and U2683 (N_2683,N_401,N_1050);
and U2684 (N_2684,N_1689,N_1388);
nand U2685 (N_2685,N_116,N_301);
xnor U2686 (N_2686,N_2248,N_2219);
nor U2687 (N_2687,N_564,N_2206);
nor U2688 (N_2688,N_2086,N_134);
nand U2689 (N_2689,N_126,N_1171);
or U2690 (N_2690,N_1332,N_1106);
or U2691 (N_2691,N_668,N_1615);
nor U2692 (N_2692,N_1984,N_249);
and U2693 (N_2693,N_1792,N_1041);
and U2694 (N_2694,N_1851,N_1257);
or U2695 (N_2695,N_32,N_609);
nor U2696 (N_2696,N_203,N_1070);
nor U2697 (N_2697,N_506,N_42);
xnor U2698 (N_2698,N_1212,N_139);
and U2699 (N_2699,N_1467,N_1161);
or U2700 (N_2700,N_1669,N_1367);
or U2701 (N_2701,N_1801,N_819);
nand U2702 (N_2702,N_1797,N_2245);
nand U2703 (N_2703,N_1897,N_1920);
and U2704 (N_2704,N_2098,N_313);
xnor U2705 (N_2705,N_620,N_985);
nor U2706 (N_2706,N_1372,N_1478);
nor U2707 (N_2707,N_2266,N_1360);
and U2708 (N_2708,N_1351,N_532);
and U2709 (N_2709,N_1855,N_530);
nor U2710 (N_2710,N_991,N_1811);
and U2711 (N_2711,N_1045,N_445);
nand U2712 (N_2712,N_1540,N_1456);
or U2713 (N_2713,N_337,N_2460);
or U2714 (N_2714,N_1739,N_759);
nor U2715 (N_2715,N_811,N_275);
nand U2716 (N_2716,N_1175,N_1163);
nand U2717 (N_2717,N_1137,N_2051);
nand U2718 (N_2718,N_2092,N_851);
or U2719 (N_2719,N_2137,N_2399);
and U2720 (N_2720,N_2358,N_1625);
and U2721 (N_2721,N_2474,N_2074);
nor U2722 (N_2722,N_768,N_860);
or U2723 (N_2723,N_1818,N_864);
xnor U2724 (N_2724,N_849,N_1230);
or U2725 (N_2725,N_457,N_263);
or U2726 (N_2726,N_296,N_357);
nand U2727 (N_2727,N_1671,N_2240);
nand U2728 (N_2728,N_1502,N_468);
xor U2729 (N_2729,N_26,N_1768);
xor U2730 (N_2730,N_1565,N_1073);
or U2731 (N_2731,N_2169,N_60);
and U2732 (N_2732,N_1636,N_431);
or U2733 (N_2733,N_1829,N_615);
nor U2734 (N_2734,N_1715,N_1986);
nor U2735 (N_2735,N_2463,N_1274);
nand U2736 (N_2736,N_2280,N_2008);
or U2737 (N_2737,N_2040,N_2190);
nand U2738 (N_2738,N_283,N_861);
and U2739 (N_2739,N_372,N_1773);
and U2740 (N_2740,N_577,N_655);
and U2741 (N_2741,N_2186,N_1350);
nand U2742 (N_2742,N_460,N_574);
nor U2743 (N_2743,N_1515,N_2369);
and U2744 (N_2744,N_1673,N_640);
and U2745 (N_2745,N_1555,N_1333);
or U2746 (N_2746,N_1403,N_2404);
and U2747 (N_2747,N_1950,N_1311);
or U2748 (N_2748,N_1602,N_1069);
nand U2749 (N_2749,N_1646,N_195);
or U2750 (N_2750,N_1947,N_805);
nor U2751 (N_2751,N_1119,N_2108);
or U2752 (N_2752,N_408,N_876);
nand U2753 (N_2753,N_1981,N_650);
nor U2754 (N_2754,N_31,N_135);
nand U2755 (N_2755,N_2493,N_52);
or U2756 (N_2756,N_2288,N_1927);
nor U2757 (N_2757,N_1975,N_45);
xor U2758 (N_2758,N_1324,N_316);
or U2759 (N_2759,N_2151,N_938);
or U2760 (N_2760,N_1810,N_2371);
nor U2761 (N_2761,N_1666,N_289);
nand U2762 (N_2762,N_1170,N_1943);
or U2763 (N_2763,N_568,N_2357);
nor U2764 (N_2764,N_2391,N_603);
and U2765 (N_2765,N_1965,N_1214);
and U2766 (N_2766,N_2320,N_1104);
nand U2767 (N_2767,N_2423,N_1992);
xnor U2768 (N_2768,N_228,N_330);
nand U2769 (N_2769,N_2014,N_1411);
xor U2770 (N_2770,N_634,N_2383);
and U2771 (N_2771,N_291,N_2189);
nor U2772 (N_2772,N_2468,N_1980);
and U2773 (N_2773,N_1264,N_1075);
nand U2774 (N_2774,N_1256,N_1501);
nor U2775 (N_2775,N_803,N_575);
or U2776 (N_2776,N_2331,N_879);
or U2777 (N_2777,N_927,N_1509);
nor U2778 (N_2778,N_1135,N_1908);
or U2779 (N_2779,N_997,N_2279);
or U2780 (N_2780,N_493,N_1809);
nor U2781 (N_2781,N_602,N_309);
and U2782 (N_2782,N_147,N_729);
or U2783 (N_2783,N_753,N_834);
xnor U2784 (N_2784,N_1706,N_1679);
and U2785 (N_2785,N_2123,N_2380);
and U2786 (N_2786,N_447,N_41);
nor U2787 (N_2787,N_2,N_1708);
nand U2788 (N_2788,N_2334,N_795);
nor U2789 (N_2789,N_2333,N_221);
nor U2790 (N_2790,N_2448,N_1910);
nand U2791 (N_2791,N_636,N_725);
nor U2792 (N_2792,N_1952,N_479);
or U2793 (N_2793,N_558,N_1948);
xnor U2794 (N_2794,N_287,N_1060);
nand U2795 (N_2795,N_839,N_2260);
and U2796 (N_2796,N_2039,N_1368);
nand U2797 (N_2797,N_2078,N_382);
and U2798 (N_2798,N_315,N_1366);
nor U2799 (N_2799,N_1654,N_1017);
nand U2800 (N_2800,N_345,N_1296);
and U2801 (N_2801,N_627,N_1334);
nor U2802 (N_2802,N_1722,N_2350);
nor U2803 (N_2803,N_711,N_1590);
and U2804 (N_2804,N_2196,N_207);
and U2805 (N_2805,N_1342,N_286);
nand U2806 (N_2806,N_708,N_2439);
nor U2807 (N_2807,N_424,N_1823);
or U2808 (N_2808,N_1660,N_2070);
and U2809 (N_2809,N_2381,N_1937);
nand U2810 (N_2810,N_219,N_781);
nand U2811 (N_2811,N_2200,N_1022);
and U2812 (N_2812,N_1958,N_1656);
and U2813 (N_2813,N_1187,N_1648);
or U2814 (N_2814,N_800,N_1251);
or U2815 (N_2815,N_1833,N_802);
nor U2816 (N_2816,N_1727,N_661);
nor U2817 (N_2817,N_856,N_2272);
xnor U2818 (N_2818,N_1815,N_1754);
xnor U2819 (N_2819,N_1011,N_419);
nor U2820 (N_2820,N_1824,N_1560);
or U2821 (N_2821,N_1283,N_1744);
xnor U2822 (N_2822,N_190,N_658);
nor U2823 (N_2823,N_801,N_2158);
or U2824 (N_2824,N_1432,N_2434);
nor U2825 (N_2825,N_2094,N_2253);
or U2826 (N_2826,N_1068,N_243);
and U2827 (N_2827,N_1637,N_2255);
nand U2828 (N_2828,N_578,N_751);
nand U2829 (N_2829,N_1470,N_512);
and U2830 (N_2830,N_1131,N_1985);
or U2831 (N_2831,N_80,N_956);
nand U2832 (N_2832,N_425,N_785);
nor U2833 (N_2833,N_1471,N_1871);
and U2834 (N_2834,N_123,N_2146);
nand U2835 (N_2835,N_1601,N_1164);
and U2836 (N_2836,N_18,N_409);
nand U2837 (N_2837,N_1144,N_2413);
or U2838 (N_2838,N_1215,N_1307);
and U2839 (N_2839,N_186,N_2048);
or U2840 (N_2840,N_1775,N_1598);
or U2841 (N_2841,N_200,N_1699);
nor U2842 (N_2842,N_776,N_1341);
and U2843 (N_2843,N_1719,N_897);
xor U2844 (N_2844,N_2304,N_25);
and U2845 (N_2845,N_2372,N_495);
or U2846 (N_2846,N_2273,N_1604);
or U2847 (N_2847,N_239,N_2204);
nand U2848 (N_2848,N_1499,N_727);
nor U2849 (N_2849,N_66,N_142);
nor U2850 (N_2850,N_1804,N_1302);
nand U2851 (N_2851,N_1267,N_9);
nand U2852 (N_2852,N_1043,N_1288);
nor U2853 (N_2853,N_1899,N_2328);
nand U2854 (N_2854,N_1441,N_2484);
and U2855 (N_2855,N_2429,N_206);
or U2856 (N_2856,N_905,N_824);
nor U2857 (N_2857,N_2215,N_1430);
and U2858 (N_2858,N_1379,N_649);
or U2859 (N_2859,N_240,N_601);
and U2860 (N_2860,N_2003,N_473);
nor U2861 (N_2861,N_1780,N_197);
and U2862 (N_2862,N_1704,N_2442);
or U2863 (N_2863,N_2079,N_900);
and U2864 (N_2864,N_588,N_2164);
nand U2865 (N_2865,N_2465,N_2282);
or U2866 (N_2866,N_706,N_1166);
xnor U2867 (N_2867,N_2370,N_1177);
and U2868 (N_2868,N_1874,N_499);
or U2869 (N_2869,N_2197,N_276);
nor U2870 (N_2870,N_1108,N_1663);
or U2871 (N_2871,N_1301,N_527);
nor U2872 (N_2872,N_2302,N_306);
and U2873 (N_2873,N_1179,N_2013);
or U2874 (N_2874,N_961,N_1317);
nor U2875 (N_2875,N_1084,N_1490);
nor U2876 (N_2876,N_2444,N_1817);
and U2877 (N_2877,N_779,N_1433);
or U2878 (N_2878,N_762,N_1312);
nor U2879 (N_2879,N_973,N_1393);
nand U2880 (N_2880,N_127,N_467);
nand U2881 (N_2881,N_1426,N_778);
nand U2882 (N_2882,N_1574,N_1322);
and U2883 (N_2883,N_2222,N_943);
xor U2884 (N_2884,N_1480,N_748);
or U2885 (N_2885,N_882,N_456);
xnor U2886 (N_2886,N_1767,N_156);
nor U2887 (N_2887,N_2120,N_347);
nor U2888 (N_2888,N_1392,N_2162);
and U2889 (N_2889,N_1380,N_2101);
nand U2890 (N_2890,N_1489,N_2419);
nor U2891 (N_2891,N_1165,N_1510);
nand U2892 (N_2892,N_222,N_378);
and U2893 (N_2893,N_2479,N_1194);
or U2894 (N_2894,N_2455,N_1856);
nor U2895 (N_2895,N_2378,N_2499);
nand U2896 (N_2896,N_469,N_2281);
nor U2897 (N_2897,N_630,N_526);
and U2898 (N_2898,N_2365,N_590);
xor U2899 (N_2899,N_1895,N_1289);
nor U2900 (N_2900,N_1087,N_393);
nor U2901 (N_2901,N_1306,N_387);
and U2902 (N_2902,N_524,N_1321);
nand U2903 (N_2903,N_130,N_1032);
or U2904 (N_2904,N_1410,N_2192);
nand U2905 (N_2905,N_545,N_1009);
or U2906 (N_2906,N_202,N_2308);
nand U2907 (N_2907,N_522,N_2049);
nor U2908 (N_2908,N_1015,N_1627);
or U2909 (N_2909,N_884,N_924);
and U2910 (N_2910,N_1863,N_355);
and U2911 (N_2911,N_106,N_926);
nand U2912 (N_2912,N_213,N_2062);
nand U2913 (N_2913,N_979,N_1683);
and U2914 (N_2914,N_911,N_1922);
and U2915 (N_2915,N_944,N_461);
and U2916 (N_2916,N_910,N_1029);
xor U2917 (N_2917,N_1759,N_831);
or U2918 (N_2918,N_2312,N_1640);
nor U2919 (N_2919,N_1945,N_2344);
nor U2920 (N_2920,N_740,N_501);
and U2921 (N_2921,N_1630,N_1026);
nand U2922 (N_2922,N_1586,N_880);
and U2923 (N_2923,N_2470,N_1239);
or U2924 (N_2924,N_2337,N_1966);
nand U2925 (N_2925,N_1771,N_342);
and U2926 (N_2926,N_2491,N_1583);
nor U2927 (N_2927,N_1798,N_508);
nor U2928 (N_2928,N_807,N_1575);
nor U2929 (N_2929,N_2433,N_769);
or U2930 (N_2930,N_1048,N_328);
or U2931 (N_2931,N_1852,N_919);
nand U2932 (N_2932,N_1198,N_2335);
and U2933 (N_2933,N_1216,N_2316);
nor U2934 (N_2934,N_1866,N_148);
xor U2935 (N_2935,N_1406,N_1956);
and U2936 (N_2936,N_294,N_913);
or U2937 (N_2937,N_1756,N_755);
nand U2938 (N_2938,N_254,N_1422);
xnor U2939 (N_2939,N_8,N_533);
nor U2940 (N_2940,N_400,N_1772);
or U2941 (N_2941,N_611,N_2268);
nor U2942 (N_2942,N_2338,N_232);
nor U2943 (N_2943,N_138,N_1831);
xor U2944 (N_2944,N_278,N_826);
nand U2945 (N_2945,N_1932,N_1111);
and U2946 (N_2946,N_1925,N_1951);
nand U2947 (N_2947,N_308,N_497);
and U2948 (N_2948,N_923,N_1764);
nor U2949 (N_2949,N_626,N_209);
nand U2950 (N_2950,N_36,N_1603);
or U2951 (N_2951,N_1858,N_1080);
nor U2952 (N_2952,N_2012,N_11);
or U2953 (N_2953,N_1760,N_510);
or U2954 (N_2954,N_2223,N_1446);
nor U2955 (N_2955,N_2485,N_1300);
and U2956 (N_2956,N_1243,N_635);
nand U2957 (N_2957,N_297,N_1375);
and U2958 (N_2958,N_1142,N_561);
and U2959 (N_2959,N_1954,N_370);
or U2960 (N_2960,N_1784,N_1556);
nand U2961 (N_2961,N_1623,N_1145);
or U2962 (N_2962,N_1199,N_573);
and U2963 (N_2963,N_1796,N_367);
or U2964 (N_2964,N_1055,N_761);
or U2965 (N_2965,N_2430,N_1917);
nor U2966 (N_2966,N_295,N_1358);
or U2967 (N_2967,N_1482,N_515);
or U2968 (N_2968,N_1588,N_1967);
or U2969 (N_2969,N_2226,N_1572);
nor U2970 (N_2970,N_2227,N_877);
and U2971 (N_2971,N_1415,N_1533);
or U2972 (N_2972,N_1761,N_546);
and U2973 (N_2973,N_525,N_2379);
or U2974 (N_2974,N_1308,N_1979);
xnor U2975 (N_2975,N_288,N_737);
and U2976 (N_2976,N_1969,N_173);
nand U2977 (N_2977,N_982,N_1207);
or U2978 (N_2978,N_318,N_1258);
nor U2979 (N_2979,N_1331,N_720);
or U2980 (N_2980,N_1310,N_146);
and U2981 (N_2981,N_2053,N_716);
and U2982 (N_2982,N_1440,N_2242);
nor U2983 (N_2983,N_1353,N_1019);
or U2984 (N_2984,N_16,N_1386);
and U2985 (N_2985,N_1990,N_300);
nand U2986 (N_2986,N_144,N_374);
nor U2987 (N_2987,N_30,N_1326);
nor U2988 (N_2988,N_1946,N_572);
nor U2989 (N_2989,N_380,N_260);
xor U2990 (N_2990,N_1412,N_1983);
nand U2991 (N_2991,N_307,N_912);
and U2992 (N_2992,N_413,N_1449);
and U2993 (N_2993,N_1034,N_2224);
or U2994 (N_2994,N_621,N_1261);
nor U2995 (N_2995,N_2031,N_1685);
nand U2996 (N_2996,N_88,N_405);
nor U2997 (N_2997,N_1619,N_1294);
nand U2998 (N_2998,N_329,N_1535);
nor U2999 (N_2999,N_1718,N_1072);
or U3000 (N_3000,N_1250,N_1733);
nand U3001 (N_3001,N_554,N_2327);
and U3002 (N_3002,N_1472,N_1731);
or U3003 (N_3003,N_1645,N_1561);
nor U3004 (N_3004,N_2249,N_717);
and U3005 (N_3005,N_710,N_451);
nor U3006 (N_3006,N_2394,N_504);
nand U3007 (N_3007,N_1204,N_1748);
nor U3008 (N_3008,N_854,N_2042);
nor U3009 (N_3009,N_290,N_730);
nand U3010 (N_3010,N_2246,N_2126);
xor U3011 (N_3011,N_1263,N_1240);
and U3012 (N_3012,N_1832,N_1550);
or U3013 (N_3013,N_1890,N_2270);
and U3014 (N_3014,N_1680,N_181);
and U3015 (N_3015,N_2144,N_810);
nand U3016 (N_3016,N_2210,N_2077);
xor U3017 (N_3017,N_2374,N_521);
xor U3018 (N_3018,N_2482,N_959);
or U3019 (N_3019,N_191,N_100);
and U3020 (N_3020,N_217,N_2157);
nor U3021 (N_3021,N_792,N_1323);
and U3022 (N_3022,N_1488,N_322);
nor U3023 (N_3023,N_1695,N_267);
nand U3024 (N_3024,N_893,N_1955);
nor U3025 (N_3025,N_1387,N_793);
or U3026 (N_3026,N_1071,N_1732);
or U3027 (N_3027,N_582,N_1989);
nor U3028 (N_3028,N_1693,N_2417);
and U3029 (N_3029,N_1089,N_242);
and U3030 (N_3030,N_193,N_820);
xor U3031 (N_3031,N_580,N_462);
nor U3032 (N_3032,N_332,N_1609);
and U3033 (N_3033,N_2239,N_366);
or U3034 (N_3034,N_1181,N_164);
nand U3035 (N_3035,N_2149,N_1543);
or U3036 (N_3036,N_1115,N_365);
and U3037 (N_3037,N_71,N_1664);
nand U3038 (N_3038,N_269,N_1425);
xnor U3039 (N_3039,N_1617,N_1447);
nor U3040 (N_3040,N_907,N_666);
nand U3041 (N_3041,N_1524,N_2393);
nor U3042 (N_3042,N_1936,N_872);
nand U3043 (N_3043,N_403,N_2489);
and U3044 (N_3044,N_487,N_845);
xnor U3045 (N_3045,N_1971,N_1241);
nor U3046 (N_3046,N_1994,N_1841);
nor U3047 (N_3047,N_1000,N_503);
nand U3048 (N_3048,N_2277,N_1495);
nor U3049 (N_3049,N_1374,N_364);
nor U3050 (N_3050,N_1612,N_266);
and U3051 (N_3051,N_268,N_1928);
nor U3052 (N_3052,N_592,N_1867);
and U3053 (N_3053,N_2167,N_1558);
nand U3054 (N_3054,N_2382,N_1778);
nor U3055 (N_3055,N_1132,N_2083);
xor U3056 (N_3056,N_1455,N_746);
and U3057 (N_3057,N_844,N_1058);
or U3058 (N_3058,N_1716,N_1837);
and U3059 (N_3059,N_1242,N_653);
and U3060 (N_3060,N_1325,N_2080);
nand U3061 (N_3061,N_426,N_102);
nor U3062 (N_3062,N_1892,N_1390);
nor U3063 (N_3063,N_1794,N_1620);
and U3064 (N_3064,N_2205,N_1913);
nor U3065 (N_3065,N_848,N_2134);
nand U3066 (N_3066,N_326,N_2293);
and U3067 (N_3067,N_1024,N_1082);
nand U3068 (N_3068,N_619,N_2309);
nor U3069 (N_3069,N_2212,N_1668);
and U3070 (N_3070,N_1921,N_2258);
nand U3071 (N_3071,N_2473,N_772);
nand U3072 (N_3072,N_2229,N_2267);
xnor U3073 (N_3073,N_2035,N_1081);
nand U3074 (N_3074,N_1551,N_1781);
or U3075 (N_3075,N_391,N_2096);
or U3076 (N_3076,N_1266,N_1201);
nand U3077 (N_3077,N_338,N_528);
or U3078 (N_3078,N_2109,N_865);
or U3079 (N_3079,N_2466,N_1621);
and U3080 (N_3080,N_1020,N_2140);
nand U3081 (N_3081,N_452,N_2179);
nand U3082 (N_3082,N_1063,N_1850);
nor U3083 (N_3083,N_1205,N_111);
or U3084 (N_3084,N_1231,N_1407);
xor U3085 (N_3085,N_885,N_1876);
or U3086 (N_3086,N_2483,N_1028);
or U3087 (N_3087,N_1428,N_311);
or U3088 (N_3088,N_1894,N_1121);
nor U3089 (N_3089,N_836,N_360);
nor U3090 (N_3090,N_1228,N_2208);
xnor U3091 (N_3091,N_1227,N_696);
and U3092 (N_3092,N_607,N_2418);
and U3093 (N_3093,N_1587,N_108);
or U3094 (N_3094,N_1938,N_2002);
or U3095 (N_3095,N_1464,N_199);
nor U3096 (N_3096,N_1315,N_2015);
and U3097 (N_3097,N_1802,N_543);
or U3098 (N_3098,N_1652,N_814);
nor U3099 (N_3099,N_852,N_2122);
nor U3100 (N_3100,N_1688,N_95);
and U3101 (N_3101,N_523,N_2217);
nor U3102 (N_3102,N_6,N_1762);
or U3103 (N_3103,N_691,N_1738);
or U3104 (N_3104,N_2221,N_1347);
or U3105 (N_3105,N_1101,N_789);
nand U3106 (N_3106,N_1429,N_414);
nand U3107 (N_3107,N_1674,N_1662);
or U3108 (N_3108,N_816,N_1217);
or U3109 (N_3109,N_1597,N_2004);
and U3110 (N_3110,N_1040,N_808);
nand U3111 (N_3111,N_1846,N_2351);
nor U3112 (N_3112,N_103,N_773);
xor U3113 (N_3113,N_1065,N_1641);
nand U3114 (N_3114,N_771,N_1549);
nor U3115 (N_3115,N_868,N_1210);
nand U3116 (N_3116,N_205,N_319);
xnor U3117 (N_3117,N_612,N_1492);
or U3118 (N_3118,N_1496,N_579);
and U3119 (N_3119,N_2230,N_17);
or U3120 (N_3120,N_1378,N_1904);
or U3121 (N_3121,N_964,N_420);
nand U3122 (N_3122,N_1795,N_1548);
nand U3123 (N_3123,N_934,N_2464);
and U3124 (N_3124,N_1125,N_1860);
or U3125 (N_3125,N_2076,N_1628);
nand U3126 (N_3126,N_1421,N_450);
or U3127 (N_3127,N_2424,N_2091);
or U3128 (N_3128,N_618,N_1377);
and U3129 (N_3129,N_641,N_1202);
nor U3130 (N_3130,N_1234,N_344);
or U3131 (N_3131,N_1381,N_2456);
nand U3132 (N_3132,N_1105,N_1373);
nor U3133 (N_3133,N_1180,N_1741);
xor U3134 (N_3134,N_1178,N_110);
nand U3135 (N_3135,N_486,N_1057);
or U3136 (N_3136,N_459,N_2475);
and U3137 (N_3137,N_1404,N_343);
or U3138 (N_3138,N_1878,N_1585);
or U3139 (N_3139,N_1445,N_1238);
nand U3140 (N_3140,N_4,N_2361);
and U3141 (N_3141,N_2467,N_1140);
nand U3142 (N_3142,N_2353,N_692);
or U3143 (N_3143,N_2203,N_211);
nor U3144 (N_3144,N_1697,N_1912);
or U3145 (N_3145,N_1277,N_743);
and U3146 (N_3146,N_987,N_99);
nor U3147 (N_3147,N_1891,N_2276);
nand U3148 (N_3148,N_2063,N_2170);
and U3149 (N_3149,N_2143,N_1724);
or U3150 (N_3150,N_1352,N_733);
and U3151 (N_3151,N_697,N_1534);
and U3152 (N_3152,N_2011,N_591);
and U3153 (N_3153,N_1021,N_1085);
nor U3154 (N_3154,N_1591,N_498);
nor U3155 (N_3155,N_657,N_166);
xnor U3156 (N_3156,N_2432,N_1395);
nand U3157 (N_3157,N_1939,N_1539);
and U3158 (N_3158,N_2087,N_2032);
and U3159 (N_3159,N_1343,N_951);
nor U3160 (N_3160,N_780,N_2478);
nor U3161 (N_3161,N_73,N_115);
nand U3162 (N_3162,N_1531,N_406);
nor U3163 (N_3163,N_1552,N_224);
nor U3164 (N_3164,N_122,N_2201);
and U3165 (N_3165,N_2232,N_79);
or U3166 (N_3166,N_965,N_684);
or U3167 (N_3167,N_1461,N_1035);
or U3168 (N_3168,N_1711,N_153);
nor U3169 (N_3169,N_1864,N_667);
and U3170 (N_3170,N_1370,N_2207);
xor U3171 (N_3171,N_1808,N_2278);
or U3172 (N_3172,N_131,N_732);
nor U3173 (N_3173,N_1707,N_1218);
or U3174 (N_3174,N_2451,N_2416);
or U3175 (N_3175,N_2415,N_185);
nor U3176 (N_3176,N_119,N_2131);
and U3177 (N_3177,N_2057,N_1635);
or U3178 (N_3178,N_813,N_1536);
nand U3179 (N_3179,N_970,N_1576);
nand U3180 (N_3180,N_604,N_2125);
nor U3181 (N_3181,N_2250,N_1963);
nand U3182 (N_3182,N_1618,N_2480);
nand U3183 (N_3183,N_1873,N_687);
xor U3184 (N_3184,N_2461,N_2155);
nor U3185 (N_3185,N_1338,N_756);
and U3186 (N_3186,N_990,N_229);
and U3187 (N_3187,N_1843,N_971);
nand U3188 (N_3188,N_797,N_323);
or U3189 (N_3189,N_1340,N_1220);
and U3190 (N_3190,N_1844,N_1188);
or U3191 (N_3191,N_1091,N_1877);
or U3192 (N_3192,N_1328,N_988);
nand U3193 (N_3193,N_2025,N_883);
nand U3194 (N_3194,N_114,N_2251);
and U3195 (N_3195,N_2363,N_977);
nand U3196 (N_3196,N_866,N_1776);
nand U3197 (N_3197,N_1745,N_838);
nand U3198 (N_3198,N_734,N_33);
nor U3199 (N_3199,N_906,N_2112);
and U3200 (N_3200,N_1582,N_2160);
or U3201 (N_3201,N_133,N_1570);
or U3202 (N_3202,N_1095,N_1742);
nor U3203 (N_3203,N_2168,N_599);
and U3204 (N_3204,N_1670,N_1098);
and U3205 (N_3205,N_2177,N_2257);
xnor U3206 (N_3206,N_63,N_782);
xor U3207 (N_3207,N_832,N_1903);
and U3208 (N_3208,N_1530,N_1610);
and U3209 (N_3209,N_2082,N_544);
or U3210 (N_3210,N_1431,N_2307);
nand U3211 (N_3211,N_392,N_538);
and U3212 (N_3212,N_698,N_304);
nor U3213 (N_3213,N_963,N_51);
nor U3214 (N_3214,N_1752,N_175);
or U3215 (N_3215,N_476,N_1889);
and U3216 (N_3216,N_96,N_171);
and U3217 (N_3217,N_786,N_1713);
and U3218 (N_3218,N_1608,N_1278);
or U3219 (N_3219,N_62,N_1348);
or U3220 (N_3220,N_932,N_775);
nand U3221 (N_3221,N_1730,N_1173);
nand U3222 (N_3222,N_1337,N_629);
nor U3223 (N_3223,N_432,N_261);
or U3224 (N_3224,N_1147,N_1998);
and U3225 (N_3225,N_680,N_1541);
nor U3226 (N_3226,N_1835,N_652);
or U3227 (N_3227,N_520,N_174);
nand U3228 (N_3228,N_676,N_843);
or U3229 (N_3229,N_1622,N_537);
xor U3230 (N_3230,N_2301,N_2005);
nor U3231 (N_3231,N_314,N_1313);
nand U3232 (N_3232,N_1828,N_2006);
nor U3233 (N_3233,N_1589,N_98);
or U3234 (N_3234,N_728,N_2023);
or U3235 (N_3235,N_1133,N_796);
or U3236 (N_3236,N_583,N_516);
xnor U3237 (N_3237,N_1475,N_2052);
or U3238 (N_3238,N_847,N_280);
nor U3239 (N_3239,N_745,N_2400);
nor U3240 (N_3240,N_600,N_2422);
and U3241 (N_3241,N_2390,N_1206);
or U3242 (N_3242,N_1944,N_1514);
nor U3243 (N_3243,N_1497,N_331);
nor U3244 (N_3244,N_1037,N_1138);
nand U3245 (N_3245,N_1074,N_1010);
or U3246 (N_3246,N_1700,N_1765);
nor U3247 (N_3247,N_741,N_2097);
or U3248 (N_3248,N_340,N_1162);
nand U3249 (N_3249,N_69,N_1016);
and U3250 (N_3250,N_1469,N_2326);
and U3251 (N_3251,N_187,N_489);
or U3252 (N_3252,N_1196,N_1146);
and U3253 (N_3253,N_1281,N_689);
and U3254 (N_3254,N_1224,N_1149);
or U3255 (N_3255,N_2214,N_1408);
nor U3256 (N_3256,N_216,N_2172);
or U3257 (N_3257,N_894,N_1320);
and U3258 (N_3258,N_112,N_1498);
or U3259 (N_3259,N_999,N_2066);
or U3260 (N_3260,N_1571,N_723);
nor U3261 (N_3261,N_2121,N_1276);
nand U3262 (N_3262,N_47,N_46);
nor U3263 (N_3263,N_2235,N_2490);
nor U3264 (N_3264,N_1684,N_150);
and U3265 (N_3265,N_1687,N_1972);
or U3266 (N_3266,N_1568,N_1814);
xor U3267 (N_3267,N_265,N_1940);
xor U3268 (N_3268,N_1042,N_1580);
or U3269 (N_3269,N_2426,N_1124);
and U3270 (N_3270,N_1825,N_2044);
and U3271 (N_3271,N_674,N_1003);
and U3272 (N_3272,N_1769,N_1339);
nor U3273 (N_3273,N_2089,N_700);
nor U3274 (N_3274,N_569,N_917);
and U3275 (N_3275,N_1397,N_2305);
or U3276 (N_3276,N_124,N_1168);
and U3277 (N_3277,N_2265,N_770);
xor U3278 (N_3278,N_1061,N_1025);
or U3279 (N_3279,N_250,N_1839);
nor U3280 (N_3280,N_2354,N_563);
xnor U3281 (N_3281,N_1599,N_1682);
nand U3282 (N_3282,N_178,N_2262);
nand U3283 (N_3283,N_143,N_302);
and U3284 (N_3284,N_1254,N_7);
xnor U3285 (N_3285,N_1152,N_1139);
and U3286 (N_3286,N_953,N_2018);
or U3287 (N_3287,N_2346,N_1644);
and U3288 (N_3288,N_2184,N_3);
nand U3289 (N_3289,N_1500,N_1675);
and U3290 (N_3290,N_2180,N_368);
and U3291 (N_3291,N_1710,N_1520);
or U3292 (N_3292,N_1507,N_1361);
nor U3293 (N_3293,N_2259,N_1537);
and U3294 (N_3294,N_28,N_472);
and U3295 (N_3295,N_20,N_1600);
xnor U3296 (N_3296,N_1450,N_2336);
nor U3297 (N_3297,N_1544,N_1513);
nand U3298 (N_3298,N_947,N_589);
nor U3299 (N_3299,N_948,N_241);
nand U3300 (N_3300,N_567,N_2081);
or U3301 (N_3301,N_1840,N_1639);
and U3302 (N_3302,N_1626,N_1616);
and U3303 (N_3303,N_210,N_438);
or U3304 (N_3304,N_1799,N_390);
xor U3305 (N_3305,N_470,N_258);
and U3306 (N_3306,N_540,N_454);
nand U3307 (N_3307,N_105,N_2105);
and U3308 (N_3308,N_960,N_2100);
and U3309 (N_3309,N_282,N_1737);
or U3310 (N_3310,N_1,N_2310);
or U3311 (N_3311,N_1355,N_1245);
or U3312 (N_3312,N_2443,N_2311);
nor U3313 (N_3313,N_152,N_91);
nor U3314 (N_3314,N_2183,N_871);
nor U3315 (N_3315,N_1942,N_1260);
nor U3316 (N_3316,N_681,N_1803);
nor U3317 (N_3317,N_608,N_2202);
or U3318 (N_3318,N_1508,N_2342);
and U3319 (N_3319,N_1820,N_484);
nand U3320 (N_3320,N_163,N_1167);
xnor U3321 (N_3321,N_1857,N_557);
or U3322 (N_3322,N_552,N_1088);
nand U3323 (N_3323,N_541,N_1376);
or U3324 (N_3324,N_1007,N_162);
and U3325 (N_3325,N_253,N_2292);
nand U3326 (N_3326,N_2347,N_1439);
or U3327 (N_3327,N_298,N_356);
nand U3328 (N_3328,N_1970,N_638);
nand U3329 (N_3329,N_324,N_576);
nand U3330 (N_3330,N_859,N_889);
and U3331 (N_3331,N_777,N_993);
nand U3332 (N_3332,N_167,N_587);
nor U3333 (N_3333,N_531,N_1330);
nor U3334 (N_3334,N_1046,N_61);
and U3335 (N_3335,N_1869,N_176);
xnor U3336 (N_3336,N_2213,N_2352);
nor U3337 (N_3337,N_1632,N_1853);
xnor U3338 (N_3338,N_1849,N_2340);
and U3339 (N_3339,N_89,N_1606);
or U3340 (N_3340,N_2275,N_2236);
xnor U3341 (N_3341,N_915,N_1605);
xor U3342 (N_3342,N_644,N_1117);
and U3343 (N_3343,N_2068,N_1902);
and U3344 (N_3344,N_1102,N_1295);
xor U3345 (N_3345,N_264,N_477);
nor U3346 (N_3346,N_2036,N_507);
xnor U3347 (N_3347,N_1714,N_2385);
xor U3348 (N_3348,N_1709,N_2296);
nand U3349 (N_3349,N_1221,N_1821);
nor U3350 (N_3350,N_1286,N_549);
and U3351 (N_3351,N_2457,N_1766);
or U3352 (N_3352,N_2414,N_2356);
or U3353 (N_3353,N_992,N_10);
nor U3354 (N_3354,N_1400,N_829);
or U3355 (N_3355,N_2067,N_1968);
nor U3356 (N_3356,N_422,N_500);
and U3357 (N_3357,N_981,N_754);
and U3358 (N_3358,N_2152,N_2034);
nor U3359 (N_3359,N_1006,N_766);
nand U3360 (N_3360,N_1991,N_1934);
or U3361 (N_3361,N_904,N_749);
and U3362 (N_3362,N_1567,N_1249);
nor U3363 (N_3363,N_184,N_886);
nor U3364 (N_3364,N_787,N_235);
or U3365 (N_3365,N_1729,N_1607);
nand U3366 (N_3366,N_1518,N_1747);
and U3367 (N_3367,N_2359,N_899);
or U3368 (N_3368,N_1883,N_1233);
nor U3369 (N_3369,N_446,N_1592);
nor U3370 (N_3370,N_2104,N_373);
and U3371 (N_3371,N_248,N_1049);
or U3372 (N_3372,N_1405,N_595);
nand U3373 (N_3373,N_1880,N_67);
and U3374 (N_3374,N_281,N_448);
nor U3375 (N_3375,N_204,N_2027);
or U3376 (N_3376,N_2492,N_584);
nand U3377 (N_3377,N_1005,N_349);
nor U3378 (N_3378,N_1977,N_1882);
xnor U3379 (N_3379,N_1905,N_1787);
xnor U3380 (N_3380,N_1236,N_547);
nor U3381 (N_3381,N_957,N_662);
or U3382 (N_3382,N_2093,N_2387);
nor U3383 (N_3383,N_2176,N_867);
xor U3384 (N_3384,N_1451,N_375);
or U3385 (N_3385,N_389,N_1557);
or U3386 (N_3386,N_519,N_1705);
or U3387 (N_3387,N_2175,N_1594);
or U3388 (N_3388,N_2061,N_610);
nor U3389 (N_3389,N_1093,N_1110);
nand U3390 (N_3390,N_485,N_2450);
or U3391 (N_3391,N_1961,N_1208);
nor U3392 (N_3392,N_415,N_709);
xor U3393 (N_3393,N_1062,N_774);
xnor U3394 (N_3394,N_428,N_54);
and U3395 (N_3395,N_158,N_817);
and U3396 (N_3396,N_1678,N_2110);
nand U3397 (N_3397,N_1865,N_1077);
nand U3398 (N_3398,N_559,N_1562);
and U3399 (N_3399,N_455,N_255);
and U3400 (N_3400,N_1782,N_1845);
nand U3401 (N_3401,N_1122,N_827);
nor U3402 (N_3402,N_2195,N_1435);
nand U3403 (N_3403,N_1577,N_2411);
nor U3404 (N_3404,N_2209,N_2314);
nand U3405 (N_3405,N_293,N_929);
nor U3406 (N_3406,N_2075,N_2437);
nor U3407 (N_3407,N_1677,N_2362);
and U3408 (N_3408,N_1346,N_548);
nand U3409 (N_3409,N_1686,N_1349);
or U3410 (N_3410,N_2286,N_215);
and U3411 (N_3411,N_648,N_1389);
and U3412 (N_3412,N_1290,N_958);
nand U3413 (N_3413,N_1420,N_1542);
and U3414 (N_3414,N_220,N_835);
nand U3415 (N_3415,N_1896,N_257);
or U3416 (N_3416,N_398,N_1013);
or U3417 (N_3417,N_50,N_1336);
and U3418 (N_3418,N_1484,N_429);
or U3419 (N_3419,N_1129,N_2459);
nor U3420 (N_3420,N_930,N_334);
or U3421 (N_3421,N_65,N_677);
and U3422 (N_3422,N_2001,N_1222);
nand U3423 (N_3423,N_955,N_1504);
nor U3424 (N_3424,N_2401,N_969);
or U3425 (N_3425,N_1209,N_2124);
or U3426 (N_3426,N_2386,N_230);
nor U3427 (N_3427,N_2287,N_1816);
or U3428 (N_3428,N_1099,N_1736);
nand U3429 (N_3429,N_1030,N_120);
and U3430 (N_3430,N_72,N_1941);
nor U3431 (N_3431,N_878,N_379);
and U3432 (N_3432,N_1083,N_2375);
or U3433 (N_3433,N_1190,N_2116);
and U3434 (N_3434,N_2127,N_1356);
xnor U3435 (N_3435,N_2128,N_1774);
or U3436 (N_3436,N_1933,N_453);
or U3437 (N_3437,N_1463,N_2103);
or U3438 (N_3438,N_2254,N_1692);
xnor U3439 (N_3439,N_1566,N_2447);
nand U3440 (N_3440,N_1485,N_285);
nor U3441 (N_3441,N_2017,N_1100);
nand U3442 (N_3442,N_359,N_1757);
nor U3443 (N_3443,N_5,N_1134);
xor U3444 (N_3444,N_1481,N_954);
nand U3445 (N_3445,N_1486,N_410);
xnor U3446 (N_3446,N_1454,N_1519);
or U3447 (N_3447,N_2368,N_2130);
xnor U3448 (N_3448,N_179,N_1309);
nand U3449 (N_3449,N_1299,N_2410);
or U3450 (N_3450,N_1726,N_481);
and U3451 (N_3451,N_2291,N_1812);
nand U3452 (N_3452,N_2107,N_855);
nand U3453 (N_3453,N_177,N_1136);
or U3454 (N_3454,N_2193,N_2129);
or U3455 (N_3455,N_1785,N_238);
xnor U3456 (N_3456,N_1344,N_683);
or U3457 (N_3457,N_758,N_2138);
or U3458 (N_3458,N_1901,N_815);
nor U3459 (N_3459,N_679,N_1203);
nand U3460 (N_3460,N_2495,N_1090);
and U3461 (N_3461,N_1800,N_2496);
nand U3462 (N_3462,N_597,N_529);
nand U3463 (N_3463,N_1155,N_1974);
or U3464 (N_3464,N_1959,N_421);
nor U3465 (N_3465,N_1462,N_252);
or U3466 (N_3466,N_1734,N_862);
and U3467 (N_3467,N_59,N_920);
or U3468 (N_3468,N_14,N_231);
nand U3469 (N_3469,N_2238,N_1120);
nor U3470 (N_3470,N_1052,N_1529);
nand U3471 (N_3471,N_1316,N_1613);
or U3472 (N_3472,N_2243,N_1647);
and U3473 (N_3473,N_1130,N_1973);
and U3474 (N_3474,N_1807,N_225);
nor U3475 (N_3475,N_1038,N_2072);
and U3476 (N_3476,N_1651,N_491);
nand U3477 (N_3477,N_570,N_416);
and U3478 (N_3478,N_1721,N_647);
nand U3479 (N_3479,N_412,N_129);
nor U3480 (N_3480,N_922,N_218);
xor U3481 (N_3481,N_208,N_693);
or U3482 (N_3482,N_2132,N_1174);
nand U3483 (N_3483,N_704,N_1314);
and U3484 (N_3484,N_2133,N_2234);
and U3485 (N_3485,N_857,N_1650);
nand U3486 (N_3486,N_277,N_2161);
nor U3487 (N_3487,N_1957,N_404);
nor U3488 (N_3488,N_212,N_84);
xor U3489 (N_3489,N_1285,N_436);
nor U3490 (N_3490,N_1148,N_901);
or U3491 (N_3491,N_1868,N_440);
and U3492 (N_3492,N_292,N_731);
or U3493 (N_3493,N_1318,N_2228);
xor U3494 (N_3494,N_226,N_2322);
and U3495 (N_3495,N_1907,N_1158);
and U3496 (N_3496,N_551,N_1383);
and U3497 (N_3497,N_2056,N_1611);
or U3498 (N_3498,N_427,N_251);
xnor U3499 (N_3499,N_1813,N_742);
nand U3500 (N_3500,N_1252,N_534);
nand U3501 (N_3501,N_1213,N_1521);
nor U3502 (N_3502,N_1819,N_870);
nand U3503 (N_3503,N_1861,N_82);
nor U3504 (N_3504,N_2231,N_361);
and U3505 (N_3505,N_182,N_397);
nand U3506 (N_3506,N_1777,N_1477);
xnor U3507 (N_3507,N_671,N_1763);
xor U3508 (N_3508,N_1960,N_155);
nor U3509 (N_3509,N_739,N_1838);
nand U3510 (N_3510,N_2405,N_614);
and U3511 (N_3511,N_690,N_784);
or U3512 (N_3512,N_57,N_2261);
nor U3513 (N_3513,N_165,N_151);
or U3514 (N_3514,N_1154,N_940);
and U3515 (N_3515,N_869,N_511);
or U3516 (N_3516,N_1253,N_2318);
xor U3517 (N_3517,N_2099,N_2454);
or U3518 (N_3518,N_2476,N_1079);
nand U3519 (N_3519,N_1999,N_1886);
xor U3520 (N_3520,N_358,N_1898);
xor U3521 (N_3521,N_925,N_1436);
or U3522 (N_3522,N_354,N_196);
or U3523 (N_3523,N_714,N_2315);
and U3524 (N_3524,N_87,N_2384);
nor U3525 (N_3525,N_2194,N_157);
or U3526 (N_3526,N_669,N_2237);
nand U3527 (N_3527,N_2285,N_1438);
and U3528 (N_3528,N_2317,N_1790);
or U3529 (N_3529,N_1698,N_1755);
or U3530 (N_3530,N_488,N_989);
xor U3531 (N_3531,N_55,N_1291);
nand U3532 (N_3532,N_1189,N_321);
nand U3533 (N_3533,N_509,N_874);
and U3534 (N_3534,N_1631,N_395);
nor U3535 (N_3535,N_1466,N_631);
nor U3536 (N_3536,N_1329,N_381);
nand U3537 (N_3537,N_2396,N_1362);
nor U3538 (N_3538,N_104,N_2349);
or U3539 (N_3539,N_726,N_2084);
or U3540 (N_3540,N_686,N_2289);
nor U3541 (N_3541,N_402,N_757);
and U3542 (N_3542,N_1665,N_270);
nand U3543 (N_3543,N_984,N_22);
nor U3544 (N_3544,N_2037,N_1676);
and U3545 (N_3545,N_712,N_1287);
or U3546 (N_3546,N_201,N_2054);
and U3547 (N_3547,N_1275,N_1503);
xor U3548 (N_3548,N_1246,N_1696);
nor U3549 (N_3549,N_2156,N_812);
and U3550 (N_3550,N_1740,N_1123);
nor U3551 (N_3551,N_1402,N_639);
nand U3552 (N_3552,N_1417,N_2477);
nor U3553 (N_3553,N_514,N_672);
nor U3554 (N_3554,N_1169,N_2321);
or U3555 (N_3555,N_2024,N_1746);
or U3556 (N_3556,N_1924,N_1384);
and U3557 (N_3557,N_435,N_1423);
and U3558 (N_3558,N_718,N_2106);
nand U3559 (N_3559,N_490,N_783);
and U3560 (N_3560,N_1511,N_2114);
nor U3561 (N_3561,N_2199,N_908);
or U3562 (N_3562,N_168,N_2377);
xnor U3563 (N_3563,N_688,N_1284);
nor U3564 (N_3564,N_1004,N_2355);
xor U3565 (N_3565,N_1848,N_2136);
or U3566 (N_3566,N_1094,N_1862);
nand U3567 (N_3567,N_1900,N_2299);
nor U3568 (N_3568,N_2000,N_136);
or U3569 (N_3569,N_986,N_1427);
nand U3570 (N_3570,N_1396,N_2174);
nand U3571 (N_3571,N_983,N_2366);
nor U3572 (N_3572,N_236,N_1018);
or U3573 (N_3573,N_351,N_259);
and U3574 (N_3574,N_555,N_1914);
or U3575 (N_3575,N_623,N_2191);
xor U3576 (N_3576,N_1382,N_310);
nand U3577 (N_3577,N_660,N_2060);
nand U3578 (N_3578,N_317,N_2348);
and U3579 (N_3579,N_245,N_1834);
and U3580 (N_3580,N_1064,N_586);
and U3581 (N_3581,N_646,N_887);
nand U3582 (N_3582,N_1444,N_107);
and U3583 (N_3583,N_750,N_1458);
nand U3584 (N_3584,N_1527,N_1872);
and U3585 (N_3585,N_2409,N_1931);
nand U3586 (N_3586,N_466,N_2026);
nand U3587 (N_3587,N_2216,N_399);
nand U3588 (N_3588,N_2020,N_2016);
nand U3589 (N_3589,N_474,N_2187);
or U3590 (N_3590,N_1885,N_430);
nor U3591 (N_3591,N_2241,N_1491);
nand U3592 (N_3592,N_39,N_2181);
and U3593 (N_3593,N_1434,N_1701);
xnor U3594 (N_3594,N_1788,N_1185);
nor U3595 (N_3595,N_1659,N_49);
or U3596 (N_3596,N_853,N_830);
or U3597 (N_3597,N_2211,N_2007);
or U3598 (N_3598,N_1569,N_198);
nor U3599 (N_3599,N_571,N_94);
xor U3600 (N_3600,N_622,N_2427);
nor U3601 (N_3601,N_333,N_442);
and U3602 (N_3602,N_2332,N_553);
nor U3603 (N_3603,N_809,N_1997);
nor U3604 (N_3604,N_517,N_2043);
nand U3605 (N_3605,N_699,N_13);
nor U3606 (N_3606,N_1369,N_2283);
nand U3607 (N_3607,N_2019,N_1786);
and U3608 (N_3608,N_38,N_645);
nor U3609 (N_3609,N_873,N_2294);
nand U3610 (N_3610,N_1182,N_833);
nor U3611 (N_3611,N_1842,N_27);
xnor U3612 (N_3612,N_2088,N_2102);
or U3613 (N_3613,N_2395,N_2269);
or U3614 (N_3614,N_2111,N_2487);
nor U3615 (N_3615,N_1642,N_2339);
nand U3616 (N_3616,N_550,N_941);
xor U3617 (N_3617,N_2010,N_1691);
nand U3618 (N_3618,N_159,N_180);
or U3619 (N_3619,N_383,N_1953);
or U3620 (N_3620,N_928,N_137);
and U3621 (N_3621,N_192,N_320);
and U3622 (N_3622,N_1067,N_975);
nor U3623 (N_3623,N_1596,N_1443);
and U3624 (N_3624,N_1424,N_903);
nor U3625 (N_3625,N_1197,N_2185);
and U3626 (N_3626,N_2159,N_1059);
or U3627 (N_3627,N_1453,N_2469);
nand U3628 (N_3628,N_1584,N_1512);
nand U3629 (N_3629,N_2225,N_2029);
or U3630 (N_3630,N_1909,N_1879);
nand U3631 (N_3631,N_1579,N_613);
xor U3632 (N_3632,N_1160,N_1725);
nor U3633 (N_3633,N_2153,N_56);
xnor U3634 (N_3634,N_722,N_585);
or U3635 (N_3635,N_616,N_821);
nor U3636 (N_3636,N_1624,N_2445);
xor U3637 (N_3637,N_1822,N_2264);
nand U3638 (N_3638,N_1118,N_1268);
nand U3639 (N_3639,N_1657,N_2313);
or U3640 (N_3640,N_735,N_2038);
nand U3641 (N_3641,N_2178,N_2497);
nand U3642 (N_3642,N_1413,N_2271);
or U3643 (N_3643,N_1559,N_1244);
nand U3644 (N_3644,N_1033,N_2113);
and U3645 (N_3645,N_2435,N_724);
xor U3646 (N_3646,N_234,N_980);
and U3647 (N_3647,N_443,N_950);
or U3648 (N_3648,N_625,N_1735);
nor U3649 (N_3649,N_1305,N_1109);
or U3650 (N_3650,N_536,N_942);
and U3651 (N_3651,N_97,N_791);
and U3652 (N_3652,N_1112,N_1593);
nand U3653 (N_3653,N_388,N_675);
nor U3654 (N_3654,N_154,N_19);
nor U3655 (N_3655,N_1014,N_841);
or U3656 (N_3656,N_2141,N_1906);
xor U3657 (N_3657,N_976,N_2274);
nor U3658 (N_3658,N_1525,N_2073);
nand U3659 (N_3659,N_2364,N_1681);
nand U3660 (N_3660,N_2069,N_1614);
or U3661 (N_3661,N_1096,N_2319);
xor U3662 (N_3662,N_2458,N_695);
nand U3663 (N_3663,N_494,N_1487);
and U3664 (N_3664,N_1401,N_1474);
or U3665 (N_3665,N_633,N_1875);
or U3666 (N_3666,N_480,N_1629);
or U3667 (N_3667,N_2367,N_765);
and U3668 (N_3668,N_713,N_2406);
nand U3669 (N_3669,N_2135,N_2446);
and U3670 (N_3670,N_2330,N_2462);
nor U3671 (N_3671,N_966,N_93);
or U3672 (N_3672,N_705,N_2407);
nand U3673 (N_3673,N_1223,N_2256);
or U3674 (N_3674,N_1054,N_2046);
nand U3675 (N_3675,N_670,N_721);
nor U3676 (N_3676,N_1359,N_2412);
nand U3677 (N_3677,N_12,N_1354);
nand U3678 (N_3678,N_747,N_1516);
nand U3679 (N_3679,N_2009,N_2059);
nor U3680 (N_3680,N_1720,N_1248);
and U3681 (N_3681,N_1103,N_1229);
nand U3682 (N_3682,N_2498,N_1219);
and U3683 (N_3683,N_1184,N_1634);
nand U3684 (N_3684,N_121,N_1269);
nor U3685 (N_3685,N_890,N_273);
nand U3686 (N_3686,N_962,N_1506);
and U3687 (N_3687,N_566,N_1791);
and U3688 (N_3688,N_1259,N_377);
and U3689 (N_3689,N_471,N_227);
and U3690 (N_3690,N_1528,N_1793);
nor U3691 (N_3691,N_1522,N_974);
nand U3692 (N_3692,N_244,N_145);
or U3693 (N_3693,N_952,N_141);
or U3694 (N_3694,N_1159,N_29);
nor U3695 (N_3695,N_1001,N_2115);
and U3696 (N_3696,N_475,N_2452);
nor U3697 (N_3697,N_1483,N_967);
and U3698 (N_3698,N_1581,N_703);
or U3699 (N_3699,N_1023,N_2047);
nor U3700 (N_3700,N_1113,N_788);
nand U3701 (N_3701,N_2165,N_1526);
nor U3702 (N_3702,N_2021,N_840);
nand U3703 (N_3703,N_2295,N_1553);
or U3704 (N_3704,N_128,N_274);
or U3705 (N_3705,N_58,N_1723);
and U3706 (N_3706,N_1643,N_624);
and U3707 (N_3707,N_888,N_188);
or U3708 (N_3708,N_2420,N_2431);
and U3709 (N_3709,N_194,N_2341);
and U3710 (N_3710,N_1728,N_828);
nor U3711 (N_3711,N_2471,N_2139);
and U3712 (N_3712,N_2163,N_24);
or U3713 (N_3713,N_1505,N_437);
nand U3714 (N_3714,N_21,N_902);
nor U3715 (N_3715,N_2325,N_1779);
nand U3716 (N_3716,N_1473,N_172);
nor U3717 (N_3717,N_1319,N_2402);
and U3718 (N_3718,N_2300,N_303);
nor U3719 (N_3719,N_806,N_2408);
nor U3720 (N_3720,N_1211,N_2095);
nand U3721 (N_3721,N_411,N_2058);
and U3722 (N_3722,N_1564,N_1661);
or U3723 (N_3723,N_1976,N_48);
or U3724 (N_3724,N_823,N_2388);
and U3725 (N_3725,N_2117,N_799);
nand U3726 (N_3726,N_909,N_363);
nand U3727 (N_3727,N_1371,N_2494);
nor U3728 (N_3728,N_1888,N_1247);
nor U3729 (N_3729,N_233,N_875);
nand U3730 (N_3730,N_417,N_1667);
nor U3731 (N_3731,N_1457,N_78);
and U3732 (N_3732,N_542,N_1127);
nand U3733 (N_3733,N_896,N_764);
nand U3734 (N_3734,N_1327,N_945);
nand U3735 (N_3735,N_846,N_284);
nand U3736 (N_3736,N_1448,N_2345);
or U3737 (N_3737,N_642,N_1232);
nand U3738 (N_3738,N_1658,N_562);
and U3739 (N_3739,N_1712,N_825);
xnor U3740 (N_3740,N_1391,N_518);
xnor U3741 (N_3741,N_1964,N_1929);
nand U3742 (N_3742,N_2421,N_1262);
or U3743 (N_3743,N_565,N_663);
nor U3744 (N_3744,N_632,N_327);
nor U3745 (N_3745,N_246,N_1414);
nor U3746 (N_3746,N_1717,N_64);
xor U3747 (N_3747,N_1398,N_931);
nor U3748 (N_3748,N_1538,N_935);
xnor U3749 (N_3749,N_23,N_1002);
and U3750 (N_3750,N_894,N_1499);
xor U3751 (N_3751,N_983,N_278);
nor U3752 (N_3752,N_1423,N_1864);
nor U3753 (N_3753,N_1050,N_831);
and U3754 (N_3754,N_2263,N_912);
xnor U3755 (N_3755,N_1175,N_405);
nand U3756 (N_3756,N_2425,N_561);
nand U3757 (N_3757,N_773,N_432);
and U3758 (N_3758,N_249,N_1654);
or U3759 (N_3759,N_709,N_1943);
nand U3760 (N_3760,N_1923,N_450);
nand U3761 (N_3761,N_2031,N_2160);
or U3762 (N_3762,N_1960,N_1972);
nand U3763 (N_3763,N_807,N_1223);
nor U3764 (N_3764,N_1533,N_488);
or U3765 (N_3765,N_1437,N_210);
and U3766 (N_3766,N_438,N_2268);
xnor U3767 (N_3767,N_2208,N_2234);
or U3768 (N_3768,N_1225,N_1710);
nor U3769 (N_3769,N_1524,N_618);
xnor U3770 (N_3770,N_509,N_2051);
nor U3771 (N_3771,N_1572,N_1707);
and U3772 (N_3772,N_2010,N_1621);
nand U3773 (N_3773,N_1497,N_56);
nor U3774 (N_3774,N_148,N_235);
nand U3775 (N_3775,N_2130,N_1674);
or U3776 (N_3776,N_19,N_1927);
nor U3777 (N_3777,N_2161,N_459);
nand U3778 (N_3778,N_1969,N_613);
nand U3779 (N_3779,N_2452,N_386);
and U3780 (N_3780,N_1483,N_1506);
or U3781 (N_3781,N_981,N_924);
xor U3782 (N_3782,N_513,N_1175);
xnor U3783 (N_3783,N_2005,N_261);
or U3784 (N_3784,N_265,N_2162);
and U3785 (N_3785,N_2152,N_2081);
nand U3786 (N_3786,N_1829,N_1190);
xor U3787 (N_3787,N_770,N_2355);
xor U3788 (N_3788,N_2031,N_2063);
nand U3789 (N_3789,N_68,N_2258);
xnor U3790 (N_3790,N_622,N_2113);
and U3791 (N_3791,N_1819,N_2167);
nand U3792 (N_3792,N_919,N_469);
or U3793 (N_3793,N_1628,N_1066);
and U3794 (N_3794,N_1370,N_2041);
nor U3795 (N_3795,N_1432,N_670);
xnor U3796 (N_3796,N_2086,N_807);
nor U3797 (N_3797,N_269,N_2314);
or U3798 (N_3798,N_366,N_2072);
nand U3799 (N_3799,N_2092,N_1814);
or U3800 (N_3800,N_2224,N_1112);
nor U3801 (N_3801,N_1955,N_1803);
and U3802 (N_3802,N_2224,N_203);
nor U3803 (N_3803,N_355,N_769);
and U3804 (N_3804,N_1389,N_1616);
or U3805 (N_3805,N_1985,N_499);
or U3806 (N_3806,N_2133,N_1885);
or U3807 (N_3807,N_1855,N_74);
nand U3808 (N_3808,N_230,N_1047);
or U3809 (N_3809,N_1566,N_2486);
or U3810 (N_3810,N_930,N_1026);
nor U3811 (N_3811,N_1668,N_520);
nand U3812 (N_3812,N_2327,N_1704);
and U3813 (N_3813,N_1494,N_677);
xor U3814 (N_3814,N_1412,N_398);
or U3815 (N_3815,N_2433,N_1090);
xnor U3816 (N_3816,N_1819,N_40);
xor U3817 (N_3817,N_2093,N_1969);
nand U3818 (N_3818,N_86,N_1348);
or U3819 (N_3819,N_81,N_1940);
and U3820 (N_3820,N_2302,N_1988);
nand U3821 (N_3821,N_2369,N_1218);
or U3822 (N_3822,N_2454,N_2371);
and U3823 (N_3823,N_2369,N_966);
xnor U3824 (N_3824,N_2021,N_1728);
nor U3825 (N_3825,N_681,N_927);
or U3826 (N_3826,N_2074,N_507);
or U3827 (N_3827,N_2374,N_274);
nand U3828 (N_3828,N_1522,N_1591);
and U3829 (N_3829,N_2177,N_1065);
xnor U3830 (N_3830,N_1107,N_1856);
nand U3831 (N_3831,N_1953,N_2334);
nor U3832 (N_3832,N_285,N_1376);
nand U3833 (N_3833,N_743,N_136);
nor U3834 (N_3834,N_765,N_2413);
and U3835 (N_3835,N_2193,N_906);
nand U3836 (N_3836,N_2206,N_1449);
xor U3837 (N_3837,N_150,N_441);
or U3838 (N_3838,N_482,N_1599);
nor U3839 (N_3839,N_1088,N_708);
and U3840 (N_3840,N_99,N_2294);
nor U3841 (N_3841,N_448,N_1769);
nand U3842 (N_3842,N_1669,N_449);
or U3843 (N_3843,N_566,N_74);
nor U3844 (N_3844,N_523,N_328);
and U3845 (N_3845,N_2096,N_2164);
and U3846 (N_3846,N_68,N_717);
nor U3847 (N_3847,N_1316,N_1690);
or U3848 (N_3848,N_1450,N_2390);
nand U3849 (N_3849,N_1667,N_94);
and U3850 (N_3850,N_2008,N_1205);
and U3851 (N_3851,N_898,N_1775);
or U3852 (N_3852,N_1804,N_789);
or U3853 (N_3853,N_1825,N_2029);
nand U3854 (N_3854,N_895,N_1976);
nand U3855 (N_3855,N_1772,N_987);
nor U3856 (N_3856,N_1886,N_2419);
nand U3857 (N_3857,N_945,N_1857);
nor U3858 (N_3858,N_47,N_1461);
and U3859 (N_3859,N_656,N_966);
or U3860 (N_3860,N_1329,N_2493);
nand U3861 (N_3861,N_2387,N_218);
nand U3862 (N_3862,N_2193,N_1030);
and U3863 (N_3863,N_1961,N_985);
nor U3864 (N_3864,N_2034,N_2069);
or U3865 (N_3865,N_1982,N_92);
nand U3866 (N_3866,N_1044,N_316);
and U3867 (N_3867,N_1943,N_722);
nor U3868 (N_3868,N_755,N_2006);
xor U3869 (N_3869,N_1222,N_407);
and U3870 (N_3870,N_358,N_1810);
nor U3871 (N_3871,N_1662,N_2379);
nor U3872 (N_3872,N_1225,N_391);
nand U3873 (N_3873,N_215,N_1200);
nand U3874 (N_3874,N_631,N_2363);
xor U3875 (N_3875,N_753,N_2326);
xor U3876 (N_3876,N_1126,N_2413);
nand U3877 (N_3877,N_1695,N_919);
or U3878 (N_3878,N_2148,N_2476);
or U3879 (N_3879,N_763,N_165);
nand U3880 (N_3880,N_2395,N_1872);
nor U3881 (N_3881,N_1828,N_189);
nand U3882 (N_3882,N_346,N_1495);
xor U3883 (N_3883,N_196,N_95);
nor U3884 (N_3884,N_1976,N_1099);
nor U3885 (N_3885,N_1584,N_610);
nand U3886 (N_3886,N_617,N_1647);
or U3887 (N_3887,N_1948,N_540);
and U3888 (N_3888,N_657,N_147);
nand U3889 (N_3889,N_1767,N_2237);
nor U3890 (N_3890,N_107,N_1017);
and U3891 (N_3891,N_1633,N_28);
or U3892 (N_3892,N_1692,N_1565);
nor U3893 (N_3893,N_713,N_32);
and U3894 (N_3894,N_1227,N_655);
nor U3895 (N_3895,N_1581,N_286);
nand U3896 (N_3896,N_171,N_145);
or U3897 (N_3897,N_408,N_1383);
or U3898 (N_3898,N_1346,N_2280);
nor U3899 (N_3899,N_1160,N_1581);
or U3900 (N_3900,N_2456,N_305);
and U3901 (N_3901,N_1965,N_1747);
or U3902 (N_3902,N_2108,N_566);
and U3903 (N_3903,N_353,N_1163);
and U3904 (N_3904,N_377,N_1552);
nand U3905 (N_3905,N_1673,N_2497);
and U3906 (N_3906,N_691,N_509);
and U3907 (N_3907,N_1563,N_952);
or U3908 (N_3908,N_1176,N_1284);
nor U3909 (N_3909,N_2276,N_1617);
nand U3910 (N_3910,N_100,N_2494);
or U3911 (N_3911,N_1019,N_2015);
xnor U3912 (N_3912,N_1811,N_804);
or U3913 (N_3913,N_2175,N_2345);
nor U3914 (N_3914,N_248,N_1985);
nor U3915 (N_3915,N_818,N_2295);
nand U3916 (N_3916,N_1824,N_2057);
and U3917 (N_3917,N_196,N_346);
or U3918 (N_3918,N_2037,N_1504);
or U3919 (N_3919,N_1171,N_1829);
or U3920 (N_3920,N_2029,N_1144);
nand U3921 (N_3921,N_1440,N_773);
or U3922 (N_3922,N_2442,N_1007);
and U3923 (N_3923,N_1636,N_1080);
and U3924 (N_3924,N_194,N_1959);
nand U3925 (N_3925,N_1716,N_1711);
nand U3926 (N_3926,N_2394,N_279);
and U3927 (N_3927,N_1720,N_831);
nor U3928 (N_3928,N_2062,N_200);
or U3929 (N_3929,N_463,N_615);
nand U3930 (N_3930,N_278,N_1552);
or U3931 (N_3931,N_1144,N_406);
nor U3932 (N_3932,N_2466,N_1837);
nand U3933 (N_3933,N_2130,N_1908);
nor U3934 (N_3934,N_223,N_2424);
and U3935 (N_3935,N_1342,N_2148);
and U3936 (N_3936,N_649,N_1741);
nand U3937 (N_3937,N_2325,N_2181);
nand U3938 (N_3938,N_551,N_203);
or U3939 (N_3939,N_2048,N_1916);
or U3940 (N_3940,N_1891,N_822);
or U3941 (N_3941,N_2037,N_333);
and U3942 (N_3942,N_1365,N_1910);
or U3943 (N_3943,N_594,N_1585);
and U3944 (N_3944,N_255,N_166);
or U3945 (N_3945,N_191,N_674);
nand U3946 (N_3946,N_283,N_1715);
nor U3947 (N_3947,N_676,N_652);
xor U3948 (N_3948,N_151,N_1871);
nor U3949 (N_3949,N_596,N_1897);
and U3950 (N_3950,N_1836,N_2101);
and U3951 (N_3951,N_2117,N_211);
nand U3952 (N_3952,N_464,N_1768);
or U3953 (N_3953,N_2257,N_95);
and U3954 (N_3954,N_571,N_941);
or U3955 (N_3955,N_572,N_2282);
nor U3956 (N_3956,N_1147,N_2206);
or U3957 (N_3957,N_6,N_2194);
nand U3958 (N_3958,N_1813,N_1871);
xnor U3959 (N_3959,N_1624,N_1519);
nor U3960 (N_3960,N_2289,N_2322);
nor U3961 (N_3961,N_1781,N_1685);
nor U3962 (N_3962,N_1524,N_298);
or U3963 (N_3963,N_2168,N_171);
nor U3964 (N_3964,N_928,N_2264);
nor U3965 (N_3965,N_1667,N_1991);
nand U3966 (N_3966,N_1158,N_187);
nand U3967 (N_3967,N_2309,N_1024);
xor U3968 (N_3968,N_931,N_172);
nor U3969 (N_3969,N_316,N_1619);
nor U3970 (N_3970,N_48,N_1886);
nand U3971 (N_3971,N_403,N_1408);
nand U3972 (N_3972,N_1684,N_2495);
or U3973 (N_3973,N_1412,N_1523);
and U3974 (N_3974,N_34,N_529);
or U3975 (N_3975,N_448,N_2160);
and U3976 (N_3976,N_1578,N_1838);
nand U3977 (N_3977,N_515,N_1754);
nand U3978 (N_3978,N_2378,N_807);
and U3979 (N_3979,N_690,N_1741);
nor U3980 (N_3980,N_720,N_2457);
nand U3981 (N_3981,N_209,N_1773);
or U3982 (N_3982,N_542,N_494);
nand U3983 (N_3983,N_1519,N_776);
and U3984 (N_3984,N_1781,N_2109);
nand U3985 (N_3985,N_2274,N_1944);
nand U3986 (N_3986,N_742,N_1329);
nand U3987 (N_3987,N_2218,N_1879);
and U3988 (N_3988,N_667,N_1333);
or U3989 (N_3989,N_887,N_346);
nand U3990 (N_3990,N_459,N_381);
nor U3991 (N_3991,N_1284,N_159);
and U3992 (N_3992,N_1931,N_1197);
nand U3993 (N_3993,N_1422,N_773);
and U3994 (N_3994,N_157,N_1385);
nor U3995 (N_3995,N_2079,N_649);
or U3996 (N_3996,N_720,N_2227);
xnor U3997 (N_3997,N_1799,N_1466);
and U3998 (N_3998,N_624,N_1467);
or U3999 (N_3999,N_1797,N_607);
nor U4000 (N_4000,N_1172,N_479);
and U4001 (N_4001,N_1054,N_1710);
nand U4002 (N_4002,N_366,N_1008);
xnor U4003 (N_4003,N_2032,N_548);
and U4004 (N_4004,N_1711,N_279);
and U4005 (N_4005,N_62,N_1313);
nor U4006 (N_4006,N_1387,N_937);
or U4007 (N_4007,N_339,N_1207);
nor U4008 (N_4008,N_1990,N_2127);
nand U4009 (N_4009,N_2166,N_2451);
and U4010 (N_4010,N_286,N_2022);
nor U4011 (N_4011,N_2373,N_397);
or U4012 (N_4012,N_223,N_1216);
and U4013 (N_4013,N_1195,N_1633);
nand U4014 (N_4014,N_1063,N_411);
nand U4015 (N_4015,N_673,N_1207);
or U4016 (N_4016,N_47,N_662);
and U4017 (N_4017,N_1304,N_1948);
xor U4018 (N_4018,N_2033,N_288);
or U4019 (N_4019,N_1268,N_2451);
nor U4020 (N_4020,N_814,N_1617);
nor U4021 (N_4021,N_80,N_1376);
and U4022 (N_4022,N_2339,N_1394);
nand U4023 (N_4023,N_105,N_332);
nor U4024 (N_4024,N_1417,N_1500);
or U4025 (N_4025,N_709,N_59);
and U4026 (N_4026,N_62,N_2379);
or U4027 (N_4027,N_2288,N_2245);
nand U4028 (N_4028,N_1986,N_1028);
nor U4029 (N_4029,N_1102,N_185);
nor U4030 (N_4030,N_1060,N_1768);
or U4031 (N_4031,N_890,N_1195);
nor U4032 (N_4032,N_594,N_1526);
nor U4033 (N_4033,N_261,N_2290);
and U4034 (N_4034,N_1475,N_1304);
xor U4035 (N_4035,N_2489,N_447);
nand U4036 (N_4036,N_1630,N_377);
and U4037 (N_4037,N_383,N_1913);
nor U4038 (N_4038,N_1308,N_71);
or U4039 (N_4039,N_1456,N_2367);
or U4040 (N_4040,N_1838,N_1484);
nor U4041 (N_4041,N_1865,N_979);
and U4042 (N_4042,N_1336,N_1085);
nor U4043 (N_4043,N_462,N_1431);
and U4044 (N_4044,N_979,N_1710);
xor U4045 (N_4045,N_246,N_420);
or U4046 (N_4046,N_1163,N_1537);
and U4047 (N_4047,N_84,N_1411);
nand U4048 (N_4048,N_287,N_2413);
xnor U4049 (N_4049,N_1061,N_437);
nor U4050 (N_4050,N_637,N_1090);
xor U4051 (N_4051,N_61,N_174);
nor U4052 (N_4052,N_2254,N_816);
nor U4053 (N_4053,N_153,N_2360);
and U4054 (N_4054,N_2169,N_1189);
or U4055 (N_4055,N_364,N_1082);
nand U4056 (N_4056,N_900,N_29);
nor U4057 (N_4057,N_1846,N_1171);
nor U4058 (N_4058,N_2406,N_1209);
nor U4059 (N_4059,N_478,N_758);
nor U4060 (N_4060,N_1462,N_1609);
or U4061 (N_4061,N_450,N_1482);
or U4062 (N_4062,N_936,N_1714);
xnor U4063 (N_4063,N_985,N_470);
xor U4064 (N_4064,N_1520,N_548);
nor U4065 (N_4065,N_554,N_630);
or U4066 (N_4066,N_2222,N_2460);
and U4067 (N_4067,N_126,N_122);
nand U4068 (N_4068,N_1975,N_1115);
and U4069 (N_4069,N_5,N_2096);
and U4070 (N_4070,N_186,N_222);
nand U4071 (N_4071,N_1495,N_1324);
and U4072 (N_4072,N_1556,N_778);
nand U4073 (N_4073,N_2281,N_1476);
or U4074 (N_4074,N_651,N_1324);
nor U4075 (N_4075,N_2435,N_2114);
or U4076 (N_4076,N_480,N_1578);
xnor U4077 (N_4077,N_2423,N_1337);
xnor U4078 (N_4078,N_381,N_298);
or U4079 (N_4079,N_1345,N_1263);
nor U4080 (N_4080,N_2464,N_823);
or U4081 (N_4081,N_595,N_1795);
or U4082 (N_4082,N_1721,N_1640);
and U4083 (N_4083,N_1991,N_1259);
nor U4084 (N_4084,N_1911,N_49);
and U4085 (N_4085,N_1306,N_2183);
and U4086 (N_4086,N_57,N_2479);
nand U4087 (N_4087,N_79,N_1789);
and U4088 (N_4088,N_681,N_1828);
nand U4089 (N_4089,N_991,N_83);
xor U4090 (N_4090,N_1119,N_1359);
and U4091 (N_4091,N_1951,N_2272);
nor U4092 (N_4092,N_1054,N_1137);
or U4093 (N_4093,N_1897,N_825);
or U4094 (N_4094,N_1214,N_2420);
nand U4095 (N_4095,N_1029,N_758);
or U4096 (N_4096,N_1110,N_437);
and U4097 (N_4097,N_648,N_657);
and U4098 (N_4098,N_522,N_1762);
nor U4099 (N_4099,N_1434,N_1757);
or U4100 (N_4100,N_1716,N_1634);
nand U4101 (N_4101,N_913,N_2361);
nor U4102 (N_4102,N_1809,N_118);
and U4103 (N_4103,N_761,N_2200);
nand U4104 (N_4104,N_544,N_1729);
nand U4105 (N_4105,N_658,N_218);
and U4106 (N_4106,N_347,N_864);
nand U4107 (N_4107,N_1223,N_356);
nand U4108 (N_4108,N_1248,N_567);
nor U4109 (N_4109,N_1781,N_204);
or U4110 (N_4110,N_1912,N_1269);
or U4111 (N_4111,N_926,N_126);
nor U4112 (N_4112,N_56,N_1292);
or U4113 (N_4113,N_1227,N_2255);
nor U4114 (N_4114,N_2488,N_729);
nand U4115 (N_4115,N_1083,N_729);
or U4116 (N_4116,N_1647,N_2312);
nor U4117 (N_4117,N_1878,N_1449);
nor U4118 (N_4118,N_1509,N_611);
nor U4119 (N_4119,N_983,N_2291);
or U4120 (N_4120,N_1535,N_627);
or U4121 (N_4121,N_1590,N_1921);
or U4122 (N_4122,N_1590,N_1612);
nor U4123 (N_4123,N_1594,N_616);
or U4124 (N_4124,N_948,N_456);
nor U4125 (N_4125,N_2218,N_1547);
nand U4126 (N_4126,N_723,N_1687);
nand U4127 (N_4127,N_189,N_1831);
or U4128 (N_4128,N_280,N_1312);
xnor U4129 (N_4129,N_1233,N_1665);
nand U4130 (N_4130,N_2285,N_568);
or U4131 (N_4131,N_1623,N_2451);
xnor U4132 (N_4132,N_740,N_52);
or U4133 (N_4133,N_883,N_2108);
nor U4134 (N_4134,N_1371,N_1966);
nand U4135 (N_4135,N_2352,N_932);
nor U4136 (N_4136,N_2291,N_2108);
nor U4137 (N_4137,N_1697,N_1521);
and U4138 (N_4138,N_2178,N_449);
nor U4139 (N_4139,N_1804,N_347);
xor U4140 (N_4140,N_2209,N_546);
nand U4141 (N_4141,N_643,N_1188);
xnor U4142 (N_4142,N_2471,N_2304);
nor U4143 (N_4143,N_1023,N_29);
nor U4144 (N_4144,N_1701,N_190);
nor U4145 (N_4145,N_2073,N_310);
nand U4146 (N_4146,N_1734,N_2424);
or U4147 (N_4147,N_1502,N_111);
or U4148 (N_4148,N_2442,N_2285);
and U4149 (N_4149,N_683,N_1959);
nor U4150 (N_4150,N_2415,N_341);
or U4151 (N_4151,N_310,N_21);
nand U4152 (N_4152,N_336,N_1185);
and U4153 (N_4153,N_1795,N_1097);
nand U4154 (N_4154,N_2150,N_1843);
or U4155 (N_4155,N_1745,N_855);
xor U4156 (N_4156,N_203,N_1653);
and U4157 (N_4157,N_2256,N_759);
or U4158 (N_4158,N_751,N_1130);
nand U4159 (N_4159,N_1893,N_415);
nand U4160 (N_4160,N_1196,N_517);
nor U4161 (N_4161,N_1453,N_2030);
or U4162 (N_4162,N_1904,N_1447);
and U4163 (N_4163,N_1655,N_2254);
or U4164 (N_4164,N_2231,N_2446);
and U4165 (N_4165,N_2227,N_1182);
xnor U4166 (N_4166,N_1888,N_1963);
and U4167 (N_4167,N_364,N_307);
and U4168 (N_4168,N_381,N_2235);
and U4169 (N_4169,N_1179,N_1226);
and U4170 (N_4170,N_1097,N_1227);
nand U4171 (N_4171,N_2498,N_709);
or U4172 (N_4172,N_1259,N_2350);
xnor U4173 (N_4173,N_134,N_1219);
nor U4174 (N_4174,N_2221,N_339);
or U4175 (N_4175,N_1760,N_8);
nor U4176 (N_4176,N_1127,N_1046);
or U4177 (N_4177,N_1593,N_143);
nor U4178 (N_4178,N_1249,N_1775);
xor U4179 (N_4179,N_1263,N_292);
or U4180 (N_4180,N_1610,N_1309);
nor U4181 (N_4181,N_13,N_1217);
or U4182 (N_4182,N_1044,N_1740);
and U4183 (N_4183,N_1644,N_2216);
and U4184 (N_4184,N_1169,N_35);
or U4185 (N_4185,N_107,N_570);
nor U4186 (N_4186,N_232,N_656);
nand U4187 (N_4187,N_1011,N_691);
or U4188 (N_4188,N_1568,N_1313);
nor U4189 (N_4189,N_239,N_1980);
nor U4190 (N_4190,N_157,N_2284);
nor U4191 (N_4191,N_688,N_846);
and U4192 (N_4192,N_795,N_201);
and U4193 (N_4193,N_1292,N_930);
nor U4194 (N_4194,N_707,N_885);
nor U4195 (N_4195,N_1873,N_1353);
or U4196 (N_4196,N_1337,N_1346);
nor U4197 (N_4197,N_632,N_24);
or U4198 (N_4198,N_1184,N_122);
nor U4199 (N_4199,N_438,N_923);
or U4200 (N_4200,N_388,N_1383);
nand U4201 (N_4201,N_1770,N_371);
nand U4202 (N_4202,N_1137,N_2353);
or U4203 (N_4203,N_1325,N_1132);
nand U4204 (N_4204,N_47,N_171);
nor U4205 (N_4205,N_2348,N_2301);
or U4206 (N_4206,N_668,N_987);
nor U4207 (N_4207,N_1914,N_271);
nand U4208 (N_4208,N_1569,N_1677);
and U4209 (N_4209,N_1225,N_622);
nor U4210 (N_4210,N_452,N_753);
and U4211 (N_4211,N_2068,N_613);
or U4212 (N_4212,N_2428,N_1508);
and U4213 (N_4213,N_1505,N_665);
xnor U4214 (N_4214,N_1019,N_76);
xnor U4215 (N_4215,N_628,N_2039);
nor U4216 (N_4216,N_1919,N_2449);
nand U4217 (N_4217,N_2474,N_939);
and U4218 (N_4218,N_2134,N_1073);
and U4219 (N_4219,N_1639,N_1852);
and U4220 (N_4220,N_18,N_1071);
nand U4221 (N_4221,N_754,N_2040);
and U4222 (N_4222,N_1814,N_2488);
or U4223 (N_4223,N_1152,N_547);
and U4224 (N_4224,N_1421,N_482);
xnor U4225 (N_4225,N_465,N_1197);
nand U4226 (N_4226,N_2449,N_1767);
nand U4227 (N_4227,N_568,N_1306);
and U4228 (N_4228,N_1526,N_588);
or U4229 (N_4229,N_1804,N_1292);
or U4230 (N_4230,N_694,N_1944);
nor U4231 (N_4231,N_69,N_1994);
nand U4232 (N_4232,N_657,N_1990);
nand U4233 (N_4233,N_689,N_931);
nand U4234 (N_4234,N_1967,N_1209);
nand U4235 (N_4235,N_1082,N_1499);
nand U4236 (N_4236,N_47,N_302);
or U4237 (N_4237,N_159,N_380);
and U4238 (N_4238,N_750,N_2297);
nor U4239 (N_4239,N_429,N_2265);
and U4240 (N_4240,N_919,N_2186);
xnor U4241 (N_4241,N_886,N_1249);
nor U4242 (N_4242,N_1998,N_2424);
nor U4243 (N_4243,N_1571,N_678);
and U4244 (N_4244,N_801,N_779);
nor U4245 (N_4245,N_1988,N_933);
and U4246 (N_4246,N_2287,N_1834);
nand U4247 (N_4247,N_2395,N_1550);
and U4248 (N_4248,N_1649,N_619);
nand U4249 (N_4249,N_1488,N_1696);
nor U4250 (N_4250,N_1789,N_1595);
nor U4251 (N_4251,N_2315,N_1529);
nand U4252 (N_4252,N_1345,N_2392);
or U4253 (N_4253,N_1578,N_779);
and U4254 (N_4254,N_552,N_1077);
nor U4255 (N_4255,N_790,N_148);
xnor U4256 (N_4256,N_1939,N_1659);
and U4257 (N_4257,N_2203,N_2452);
or U4258 (N_4258,N_1634,N_1457);
and U4259 (N_4259,N_1728,N_1450);
and U4260 (N_4260,N_1005,N_1203);
or U4261 (N_4261,N_922,N_1083);
nor U4262 (N_4262,N_1822,N_2058);
nor U4263 (N_4263,N_992,N_2239);
or U4264 (N_4264,N_1248,N_592);
or U4265 (N_4265,N_370,N_1062);
and U4266 (N_4266,N_3,N_98);
or U4267 (N_4267,N_1704,N_196);
nand U4268 (N_4268,N_1642,N_1460);
nor U4269 (N_4269,N_1665,N_1094);
nand U4270 (N_4270,N_2241,N_2087);
xor U4271 (N_4271,N_400,N_270);
and U4272 (N_4272,N_1127,N_1113);
nand U4273 (N_4273,N_375,N_2396);
and U4274 (N_4274,N_971,N_334);
nand U4275 (N_4275,N_1939,N_761);
and U4276 (N_4276,N_851,N_979);
nand U4277 (N_4277,N_1599,N_761);
and U4278 (N_4278,N_1015,N_147);
or U4279 (N_4279,N_98,N_776);
and U4280 (N_4280,N_361,N_2198);
nor U4281 (N_4281,N_302,N_1213);
or U4282 (N_4282,N_1173,N_848);
nand U4283 (N_4283,N_2112,N_502);
and U4284 (N_4284,N_665,N_627);
and U4285 (N_4285,N_620,N_1417);
xnor U4286 (N_4286,N_1949,N_1039);
nor U4287 (N_4287,N_36,N_1689);
nor U4288 (N_4288,N_1202,N_2070);
nand U4289 (N_4289,N_449,N_84);
or U4290 (N_4290,N_1354,N_525);
and U4291 (N_4291,N_135,N_267);
nand U4292 (N_4292,N_591,N_602);
nor U4293 (N_4293,N_2428,N_1968);
or U4294 (N_4294,N_1042,N_155);
nand U4295 (N_4295,N_1730,N_2093);
or U4296 (N_4296,N_836,N_1040);
nand U4297 (N_4297,N_2121,N_1593);
xor U4298 (N_4298,N_1712,N_41);
nand U4299 (N_4299,N_823,N_1428);
and U4300 (N_4300,N_1842,N_174);
nand U4301 (N_4301,N_945,N_2177);
nand U4302 (N_4302,N_132,N_708);
nand U4303 (N_4303,N_732,N_2034);
nor U4304 (N_4304,N_2176,N_285);
and U4305 (N_4305,N_2080,N_2140);
xor U4306 (N_4306,N_925,N_535);
and U4307 (N_4307,N_2365,N_1105);
xnor U4308 (N_4308,N_1677,N_2181);
nand U4309 (N_4309,N_2258,N_958);
or U4310 (N_4310,N_2409,N_1803);
nand U4311 (N_4311,N_1320,N_585);
nor U4312 (N_4312,N_1199,N_540);
and U4313 (N_4313,N_1812,N_1423);
and U4314 (N_4314,N_2405,N_742);
nand U4315 (N_4315,N_935,N_1474);
nor U4316 (N_4316,N_1137,N_1315);
or U4317 (N_4317,N_104,N_21);
and U4318 (N_4318,N_1693,N_1157);
nand U4319 (N_4319,N_164,N_1650);
nor U4320 (N_4320,N_2374,N_465);
and U4321 (N_4321,N_2201,N_2042);
and U4322 (N_4322,N_2148,N_1965);
or U4323 (N_4323,N_497,N_599);
or U4324 (N_4324,N_1377,N_64);
xnor U4325 (N_4325,N_1241,N_1148);
or U4326 (N_4326,N_792,N_2181);
or U4327 (N_4327,N_2002,N_1374);
nor U4328 (N_4328,N_1400,N_1527);
and U4329 (N_4329,N_1911,N_2263);
and U4330 (N_4330,N_1305,N_788);
and U4331 (N_4331,N_2257,N_376);
nor U4332 (N_4332,N_1634,N_80);
and U4333 (N_4333,N_2390,N_1945);
xnor U4334 (N_4334,N_1373,N_2438);
or U4335 (N_4335,N_1628,N_246);
nand U4336 (N_4336,N_2046,N_497);
xnor U4337 (N_4337,N_479,N_450);
or U4338 (N_4338,N_661,N_833);
xnor U4339 (N_4339,N_748,N_1627);
and U4340 (N_4340,N_598,N_1118);
or U4341 (N_4341,N_2092,N_154);
nand U4342 (N_4342,N_2483,N_1821);
nand U4343 (N_4343,N_757,N_1462);
and U4344 (N_4344,N_243,N_563);
nand U4345 (N_4345,N_1042,N_1765);
nor U4346 (N_4346,N_15,N_1344);
and U4347 (N_4347,N_416,N_1883);
nand U4348 (N_4348,N_589,N_212);
and U4349 (N_4349,N_974,N_484);
or U4350 (N_4350,N_1776,N_2087);
or U4351 (N_4351,N_876,N_905);
and U4352 (N_4352,N_2108,N_767);
and U4353 (N_4353,N_1691,N_242);
and U4354 (N_4354,N_1193,N_2343);
and U4355 (N_4355,N_1379,N_860);
and U4356 (N_4356,N_519,N_306);
nor U4357 (N_4357,N_430,N_1558);
or U4358 (N_4358,N_1682,N_1330);
xnor U4359 (N_4359,N_760,N_2431);
or U4360 (N_4360,N_2008,N_1050);
nand U4361 (N_4361,N_917,N_171);
and U4362 (N_4362,N_1532,N_9);
and U4363 (N_4363,N_1596,N_1724);
nor U4364 (N_4364,N_523,N_1095);
or U4365 (N_4365,N_1552,N_466);
and U4366 (N_4366,N_685,N_552);
or U4367 (N_4367,N_1828,N_1267);
or U4368 (N_4368,N_1814,N_1400);
nand U4369 (N_4369,N_979,N_688);
nand U4370 (N_4370,N_1219,N_1659);
or U4371 (N_4371,N_2305,N_2477);
and U4372 (N_4372,N_562,N_717);
and U4373 (N_4373,N_208,N_1429);
and U4374 (N_4374,N_1604,N_1052);
nand U4375 (N_4375,N_646,N_1088);
and U4376 (N_4376,N_1437,N_1274);
or U4377 (N_4377,N_2049,N_728);
nand U4378 (N_4378,N_1144,N_1627);
and U4379 (N_4379,N_911,N_230);
and U4380 (N_4380,N_777,N_1473);
nand U4381 (N_4381,N_25,N_32);
and U4382 (N_4382,N_1092,N_1670);
nand U4383 (N_4383,N_1700,N_658);
xor U4384 (N_4384,N_1448,N_1580);
nand U4385 (N_4385,N_1868,N_645);
nor U4386 (N_4386,N_1570,N_2408);
nor U4387 (N_4387,N_543,N_363);
nor U4388 (N_4388,N_335,N_491);
or U4389 (N_4389,N_1476,N_424);
and U4390 (N_4390,N_657,N_485);
nand U4391 (N_4391,N_1630,N_2238);
nand U4392 (N_4392,N_1818,N_820);
and U4393 (N_4393,N_4,N_2495);
and U4394 (N_4394,N_705,N_590);
or U4395 (N_4395,N_855,N_2383);
or U4396 (N_4396,N_1591,N_2243);
or U4397 (N_4397,N_2450,N_1293);
nor U4398 (N_4398,N_212,N_706);
or U4399 (N_4399,N_84,N_1819);
or U4400 (N_4400,N_1447,N_1062);
nand U4401 (N_4401,N_663,N_216);
or U4402 (N_4402,N_2479,N_910);
nand U4403 (N_4403,N_577,N_565);
and U4404 (N_4404,N_2220,N_1608);
or U4405 (N_4405,N_1184,N_1180);
xnor U4406 (N_4406,N_24,N_933);
nand U4407 (N_4407,N_821,N_2247);
or U4408 (N_4408,N_1304,N_688);
or U4409 (N_4409,N_1328,N_1005);
nor U4410 (N_4410,N_2427,N_1913);
or U4411 (N_4411,N_399,N_2360);
nor U4412 (N_4412,N_1173,N_1010);
nor U4413 (N_4413,N_2349,N_1187);
nor U4414 (N_4414,N_1787,N_2224);
nand U4415 (N_4415,N_325,N_1881);
or U4416 (N_4416,N_324,N_1220);
nor U4417 (N_4417,N_1225,N_1726);
and U4418 (N_4418,N_2313,N_1244);
nor U4419 (N_4419,N_52,N_999);
nand U4420 (N_4420,N_2077,N_1743);
nand U4421 (N_4421,N_1138,N_17);
nor U4422 (N_4422,N_387,N_1938);
nand U4423 (N_4423,N_1596,N_2246);
nand U4424 (N_4424,N_37,N_817);
and U4425 (N_4425,N_1796,N_747);
and U4426 (N_4426,N_2166,N_1430);
or U4427 (N_4427,N_328,N_604);
or U4428 (N_4428,N_69,N_1562);
nor U4429 (N_4429,N_1763,N_1008);
nand U4430 (N_4430,N_2480,N_151);
or U4431 (N_4431,N_80,N_22);
nor U4432 (N_4432,N_1508,N_2412);
or U4433 (N_4433,N_1230,N_1695);
or U4434 (N_4434,N_594,N_48);
or U4435 (N_4435,N_150,N_281);
and U4436 (N_4436,N_1723,N_1311);
nand U4437 (N_4437,N_1988,N_737);
nor U4438 (N_4438,N_885,N_1165);
xnor U4439 (N_4439,N_1348,N_1318);
xor U4440 (N_4440,N_2017,N_936);
and U4441 (N_4441,N_1783,N_280);
nor U4442 (N_4442,N_850,N_2302);
nor U4443 (N_4443,N_167,N_1911);
and U4444 (N_4444,N_901,N_2375);
nor U4445 (N_4445,N_815,N_2249);
nor U4446 (N_4446,N_251,N_299);
nand U4447 (N_4447,N_2485,N_1126);
nand U4448 (N_4448,N_1729,N_597);
and U4449 (N_4449,N_523,N_2411);
nand U4450 (N_4450,N_1693,N_1190);
xor U4451 (N_4451,N_2421,N_1194);
nor U4452 (N_4452,N_327,N_1694);
or U4453 (N_4453,N_756,N_1952);
nand U4454 (N_4454,N_335,N_1757);
nand U4455 (N_4455,N_562,N_2060);
or U4456 (N_4456,N_2453,N_397);
and U4457 (N_4457,N_171,N_228);
and U4458 (N_4458,N_1166,N_169);
or U4459 (N_4459,N_321,N_1732);
or U4460 (N_4460,N_1243,N_433);
or U4461 (N_4461,N_323,N_1774);
nand U4462 (N_4462,N_2495,N_1519);
or U4463 (N_4463,N_1916,N_16);
and U4464 (N_4464,N_1145,N_1356);
nand U4465 (N_4465,N_27,N_2443);
and U4466 (N_4466,N_689,N_1175);
or U4467 (N_4467,N_1267,N_853);
xnor U4468 (N_4468,N_891,N_2370);
and U4469 (N_4469,N_1573,N_2311);
nor U4470 (N_4470,N_13,N_2377);
and U4471 (N_4471,N_1957,N_154);
or U4472 (N_4472,N_706,N_2088);
or U4473 (N_4473,N_1153,N_562);
or U4474 (N_4474,N_223,N_1172);
xor U4475 (N_4475,N_1325,N_1260);
nor U4476 (N_4476,N_1210,N_2278);
xor U4477 (N_4477,N_299,N_2153);
xor U4478 (N_4478,N_1247,N_389);
or U4479 (N_4479,N_1932,N_2262);
and U4480 (N_4480,N_1820,N_1314);
and U4481 (N_4481,N_1045,N_567);
nor U4482 (N_4482,N_2230,N_1719);
or U4483 (N_4483,N_1221,N_448);
and U4484 (N_4484,N_1004,N_287);
and U4485 (N_4485,N_1770,N_646);
nand U4486 (N_4486,N_405,N_1739);
xnor U4487 (N_4487,N_68,N_253);
nor U4488 (N_4488,N_959,N_1328);
nor U4489 (N_4489,N_689,N_2006);
and U4490 (N_4490,N_112,N_1815);
nand U4491 (N_4491,N_813,N_2063);
nand U4492 (N_4492,N_2469,N_128);
or U4493 (N_4493,N_1981,N_1438);
and U4494 (N_4494,N_1799,N_124);
or U4495 (N_4495,N_2381,N_1201);
or U4496 (N_4496,N_223,N_1365);
xnor U4497 (N_4497,N_2092,N_963);
nand U4498 (N_4498,N_2274,N_896);
nand U4499 (N_4499,N_1552,N_1748);
or U4500 (N_4500,N_791,N_1170);
xor U4501 (N_4501,N_1765,N_231);
or U4502 (N_4502,N_1038,N_1087);
xor U4503 (N_4503,N_1001,N_1529);
or U4504 (N_4504,N_390,N_2275);
and U4505 (N_4505,N_395,N_1821);
nor U4506 (N_4506,N_2035,N_435);
nor U4507 (N_4507,N_1031,N_1368);
nor U4508 (N_4508,N_2169,N_2411);
and U4509 (N_4509,N_695,N_161);
nand U4510 (N_4510,N_2477,N_1443);
or U4511 (N_4511,N_1224,N_1487);
nor U4512 (N_4512,N_1765,N_1523);
and U4513 (N_4513,N_1669,N_187);
and U4514 (N_4514,N_1267,N_1570);
nand U4515 (N_4515,N_2426,N_2107);
or U4516 (N_4516,N_717,N_879);
or U4517 (N_4517,N_1487,N_1500);
and U4518 (N_4518,N_2307,N_2489);
or U4519 (N_4519,N_573,N_107);
nand U4520 (N_4520,N_2321,N_1638);
nor U4521 (N_4521,N_1585,N_58);
or U4522 (N_4522,N_2356,N_827);
nor U4523 (N_4523,N_535,N_2247);
or U4524 (N_4524,N_2130,N_474);
nand U4525 (N_4525,N_1020,N_6);
and U4526 (N_4526,N_284,N_154);
and U4527 (N_4527,N_1465,N_409);
nand U4528 (N_4528,N_2225,N_1032);
nor U4529 (N_4529,N_397,N_1652);
xor U4530 (N_4530,N_22,N_801);
nand U4531 (N_4531,N_1636,N_2097);
nor U4532 (N_4532,N_1472,N_1163);
and U4533 (N_4533,N_1276,N_568);
xor U4534 (N_4534,N_77,N_1184);
nand U4535 (N_4535,N_2215,N_881);
or U4536 (N_4536,N_1641,N_75);
and U4537 (N_4537,N_1390,N_2429);
xor U4538 (N_4538,N_1461,N_1426);
and U4539 (N_4539,N_413,N_1678);
nor U4540 (N_4540,N_826,N_2025);
and U4541 (N_4541,N_1737,N_1139);
nor U4542 (N_4542,N_336,N_1302);
xnor U4543 (N_4543,N_2341,N_966);
and U4544 (N_4544,N_224,N_1376);
nor U4545 (N_4545,N_2399,N_950);
nor U4546 (N_4546,N_1749,N_2479);
and U4547 (N_4547,N_139,N_1919);
nor U4548 (N_4548,N_1892,N_697);
and U4549 (N_4549,N_492,N_1301);
nand U4550 (N_4550,N_306,N_1571);
nand U4551 (N_4551,N_783,N_2024);
nand U4552 (N_4552,N_338,N_2312);
or U4553 (N_4553,N_1903,N_53);
nor U4554 (N_4554,N_2007,N_144);
or U4555 (N_4555,N_2125,N_1819);
and U4556 (N_4556,N_2451,N_142);
nand U4557 (N_4557,N_235,N_465);
and U4558 (N_4558,N_1497,N_2164);
nand U4559 (N_4559,N_825,N_398);
or U4560 (N_4560,N_212,N_936);
nand U4561 (N_4561,N_730,N_960);
or U4562 (N_4562,N_2144,N_226);
and U4563 (N_4563,N_73,N_2027);
nor U4564 (N_4564,N_621,N_1930);
nor U4565 (N_4565,N_228,N_1026);
nand U4566 (N_4566,N_2468,N_679);
or U4567 (N_4567,N_736,N_1425);
nor U4568 (N_4568,N_1130,N_1112);
nand U4569 (N_4569,N_749,N_309);
nand U4570 (N_4570,N_584,N_2289);
nand U4571 (N_4571,N_775,N_1821);
nor U4572 (N_4572,N_968,N_41);
nand U4573 (N_4573,N_2390,N_1773);
nand U4574 (N_4574,N_1631,N_2009);
nor U4575 (N_4575,N_1874,N_259);
and U4576 (N_4576,N_2002,N_1246);
nor U4577 (N_4577,N_2240,N_773);
nor U4578 (N_4578,N_903,N_1060);
xnor U4579 (N_4579,N_774,N_833);
and U4580 (N_4580,N_182,N_358);
and U4581 (N_4581,N_1979,N_2295);
nor U4582 (N_4582,N_2075,N_609);
nand U4583 (N_4583,N_1351,N_680);
or U4584 (N_4584,N_1668,N_1147);
nor U4585 (N_4585,N_2343,N_1039);
nand U4586 (N_4586,N_792,N_1351);
nand U4587 (N_4587,N_485,N_2376);
and U4588 (N_4588,N_1766,N_336);
and U4589 (N_4589,N_1071,N_1487);
nand U4590 (N_4590,N_1231,N_786);
and U4591 (N_4591,N_537,N_1154);
nand U4592 (N_4592,N_2411,N_370);
nand U4593 (N_4593,N_2410,N_898);
or U4594 (N_4594,N_1782,N_353);
or U4595 (N_4595,N_633,N_1183);
or U4596 (N_4596,N_812,N_2032);
nand U4597 (N_4597,N_914,N_1861);
and U4598 (N_4598,N_858,N_1394);
or U4599 (N_4599,N_496,N_2029);
nor U4600 (N_4600,N_694,N_2221);
nand U4601 (N_4601,N_1641,N_1100);
nor U4602 (N_4602,N_1642,N_664);
and U4603 (N_4603,N_1677,N_655);
nand U4604 (N_4604,N_1872,N_401);
and U4605 (N_4605,N_282,N_1310);
or U4606 (N_4606,N_1864,N_1090);
nor U4607 (N_4607,N_1223,N_731);
or U4608 (N_4608,N_2033,N_1487);
or U4609 (N_4609,N_2405,N_810);
nor U4610 (N_4610,N_301,N_2418);
nor U4611 (N_4611,N_380,N_1444);
nand U4612 (N_4612,N_957,N_1491);
or U4613 (N_4613,N_1741,N_864);
or U4614 (N_4614,N_15,N_492);
nor U4615 (N_4615,N_1579,N_57);
and U4616 (N_4616,N_900,N_286);
nand U4617 (N_4617,N_1859,N_1439);
or U4618 (N_4618,N_1318,N_1638);
nor U4619 (N_4619,N_900,N_730);
xor U4620 (N_4620,N_1549,N_1329);
nor U4621 (N_4621,N_1415,N_204);
nand U4622 (N_4622,N_659,N_2410);
nor U4623 (N_4623,N_507,N_1045);
nor U4624 (N_4624,N_1954,N_1238);
nor U4625 (N_4625,N_2030,N_536);
nand U4626 (N_4626,N_1829,N_1761);
nand U4627 (N_4627,N_1958,N_1574);
and U4628 (N_4628,N_102,N_138);
xor U4629 (N_4629,N_1188,N_2273);
and U4630 (N_4630,N_2493,N_1729);
nand U4631 (N_4631,N_1224,N_1735);
nor U4632 (N_4632,N_242,N_1934);
and U4633 (N_4633,N_475,N_1718);
nor U4634 (N_4634,N_2138,N_867);
or U4635 (N_4635,N_2493,N_249);
nand U4636 (N_4636,N_92,N_1490);
or U4637 (N_4637,N_85,N_2009);
nand U4638 (N_4638,N_1425,N_895);
nor U4639 (N_4639,N_2064,N_1542);
xor U4640 (N_4640,N_353,N_835);
nor U4641 (N_4641,N_2256,N_2030);
nor U4642 (N_4642,N_2217,N_728);
or U4643 (N_4643,N_38,N_483);
xnor U4644 (N_4644,N_305,N_407);
nand U4645 (N_4645,N_1463,N_2198);
and U4646 (N_4646,N_2318,N_218);
or U4647 (N_4647,N_375,N_941);
nor U4648 (N_4648,N_1806,N_1863);
xnor U4649 (N_4649,N_706,N_496);
and U4650 (N_4650,N_2117,N_1088);
and U4651 (N_4651,N_558,N_1446);
nand U4652 (N_4652,N_1193,N_118);
nor U4653 (N_4653,N_2124,N_13);
nand U4654 (N_4654,N_1399,N_357);
nand U4655 (N_4655,N_671,N_360);
or U4656 (N_4656,N_1346,N_629);
nand U4657 (N_4657,N_1720,N_1469);
nand U4658 (N_4658,N_1956,N_44);
and U4659 (N_4659,N_663,N_934);
and U4660 (N_4660,N_1902,N_2307);
nor U4661 (N_4661,N_2490,N_2179);
or U4662 (N_4662,N_1751,N_2444);
nor U4663 (N_4663,N_267,N_1064);
xor U4664 (N_4664,N_876,N_88);
or U4665 (N_4665,N_1760,N_1222);
nand U4666 (N_4666,N_506,N_1762);
nor U4667 (N_4667,N_2043,N_2119);
xor U4668 (N_4668,N_1508,N_411);
or U4669 (N_4669,N_839,N_148);
and U4670 (N_4670,N_799,N_1335);
or U4671 (N_4671,N_926,N_67);
or U4672 (N_4672,N_640,N_2311);
xor U4673 (N_4673,N_2123,N_1078);
nor U4674 (N_4674,N_1138,N_1880);
nand U4675 (N_4675,N_1996,N_220);
nor U4676 (N_4676,N_788,N_469);
nand U4677 (N_4677,N_211,N_780);
nor U4678 (N_4678,N_2114,N_294);
nor U4679 (N_4679,N_1646,N_1878);
and U4680 (N_4680,N_2394,N_1349);
xor U4681 (N_4681,N_1846,N_1328);
or U4682 (N_4682,N_2056,N_285);
or U4683 (N_4683,N_1139,N_444);
or U4684 (N_4684,N_1378,N_291);
xnor U4685 (N_4685,N_1041,N_816);
and U4686 (N_4686,N_93,N_261);
or U4687 (N_4687,N_406,N_1924);
or U4688 (N_4688,N_331,N_43);
nand U4689 (N_4689,N_314,N_836);
and U4690 (N_4690,N_1919,N_481);
and U4691 (N_4691,N_1448,N_382);
or U4692 (N_4692,N_1757,N_2324);
nor U4693 (N_4693,N_2304,N_130);
and U4694 (N_4694,N_755,N_2384);
xnor U4695 (N_4695,N_251,N_2276);
and U4696 (N_4696,N_1703,N_497);
nor U4697 (N_4697,N_1987,N_54);
or U4698 (N_4698,N_2148,N_1040);
xnor U4699 (N_4699,N_1469,N_1124);
and U4700 (N_4700,N_1342,N_1664);
nor U4701 (N_4701,N_557,N_234);
xor U4702 (N_4702,N_484,N_2293);
xor U4703 (N_4703,N_1762,N_1861);
nand U4704 (N_4704,N_778,N_627);
nand U4705 (N_4705,N_2317,N_909);
and U4706 (N_4706,N_988,N_2201);
nor U4707 (N_4707,N_473,N_708);
nor U4708 (N_4708,N_1397,N_1009);
and U4709 (N_4709,N_2352,N_395);
nor U4710 (N_4710,N_940,N_2287);
xor U4711 (N_4711,N_536,N_111);
xor U4712 (N_4712,N_2232,N_2142);
nand U4713 (N_4713,N_1261,N_616);
and U4714 (N_4714,N_1252,N_1372);
and U4715 (N_4715,N_2244,N_173);
nand U4716 (N_4716,N_1168,N_1894);
and U4717 (N_4717,N_1532,N_133);
xor U4718 (N_4718,N_1699,N_947);
nand U4719 (N_4719,N_1039,N_2203);
and U4720 (N_4720,N_1672,N_1319);
nor U4721 (N_4721,N_750,N_1031);
or U4722 (N_4722,N_1180,N_642);
nand U4723 (N_4723,N_192,N_2172);
xor U4724 (N_4724,N_351,N_1217);
or U4725 (N_4725,N_143,N_554);
nor U4726 (N_4726,N_1381,N_429);
and U4727 (N_4727,N_372,N_1584);
and U4728 (N_4728,N_435,N_2319);
nand U4729 (N_4729,N_614,N_1511);
xnor U4730 (N_4730,N_1630,N_2338);
nor U4731 (N_4731,N_69,N_1401);
nor U4732 (N_4732,N_332,N_640);
and U4733 (N_4733,N_1829,N_824);
nand U4734 (N_4734,N_1378,N_920);
nand U4735 (N_4735,N_733,N_261);
or U4736 (N_4736,N_1246,N_2464);
nor U4737 (N_4737,N_1507,N_613);
nand U4738 (N_4738,N_1629,N_60);
and U4739 (N_4739,N_218,N_1190);
nand U4740 (N_4740,N_1408,N_1726);
or U4741 (N_4741,N_2456,N_1706);
xnor U4742 (N_4742,N_738,N_1840);
or U4743 (N_4743,N_2320,N_2299);
and U4744 (N_4744,N_984,N_1034);
nor U4745 (N_4745,N_2210,N_1783);
and U4746 (N_4746,N_2388,N_1990);
nor U4747 (N_4747,N_1048,N_1530);
xnor U4748 (N_4748,N_372,N_2361);
nor U4749 (N_4749,N_1663,N_645);
or U4750 (N_4750,N_2089,N_1906);
nand U4751 (N_4751,N_338,N_1649);
nand U4752 (N_4752,N_1430,N_76);
nand U4753 (N_4753,N_2090,N_600);
xor U4754 (N_4754,N_363,N_1574);
nor U4755 (N_4755,N_2426,N_657);
xor U4756 (N_4756,N_2284,N_2489);
xnor U4757 (N_4757,N_236,N_2042);
nand U4758 (N_4758,N_716,N_156);
and U4759 (N_4759,N_864,N_86);
nand U4760 (N_4760,N_2201,N_2224);
nor U4761 (N_4761,N_86,N_1441);
or U4762 (N_4762,N_607,N_1750);
xor U4763 (N_4763,N_533,N_1676);
nand U4764 (N_4764,N_1959,N_183);
and U4765 (N_4765,N_427,N_1129);
or U4766 (N_4766,N_50,N_1547);
nand U4767 (N_4767,N_365,N_2242);
and U4768 (N_4768,N_1430,N_210);
nand U4769 (N_4769,N_142,N_226);
nand U4770 (N_4770,N_808,N_1446);
and U4771 (N_4771,N_141,N_2000);
nand U4772 (N_4772,N_2009,N_1026);
and U4773 (N_4773,N_302,N_1221);
or U4774 (N_4774,N_1981,N_49);
or U4775 (N_4775,N_851,N_296);
nor U4776 (N_4776,N_2172,N_1539);
nor U4777 (N_4777,N_1224,N_1120);
xor U4778 (N_4778,N_551,N_1705);
or U4779 (N_4779,N_654,N_114);
and U4780 (N_4780,N_1909,N_744);
or U4781 (N_4781,N_2395,N_2092);
or U4782 (N_4782,N_1053,N_1508);
nor U4783 (N_4783,N_492,N_992);
nor U4784 (N_4784,N_900,N_2396);
nand U4785 (N_4785,N_892,N_1052);
xor U4786 (N_4786,N_997,N_2347);
and U4787 (N_4787,N_674,N_1419);
or U4788 (N_4788,N_1896,N_1487);
nor U4789 (N_4789,N_1058,N_2300);
or U4790 (N_4790,N_624,N_542);
or U4791 (N_4791,N_1209,N_1465);
or U4792 (N_4792,N_1150,N_2161);
nand U4793 (N_4793,N_166,N_2421);
xnor U4794 (N_4794,N_1320,N_1283);
or U4795 (N_4795,N_115,N_177);
and U4796 (N_4796,N_1979,N_2474);
and U4797 (N_4797,N_523,N_2360);
nor U4798 (N_4798,N_963,N_874);
or U4799 (N_4799,N_1233,N_868);
or U4800 (N_4800,N_1013,N_1376);
and U4801 (N_4801,N_1119,N_413);
and U4802 (N_4802,N_582,N_1318);
or U4803 (N_4803,N_1716,N_874);
or U4804 (N_4804,N_2017,N_111);
nor U4805 (N_4805,N_353,N_1380);
or U4806 (N_4806,N_2482,N_1551);
or U4807 (N_4807,N_249,N_1003);
nand U4808 (N_4808,N_1958,N_1547);
nand U4809 (N_4809,N_1279,N_2066);
nor U4810 (N_4810,N_639,N_1317);
xor U4811 (N_4811,N_2158,N_2374);
nand U4812 (N_4812,N_110,N_1981);
nor U4813 (N_4813,N_2217,N_180);
and U4814 (N_4814,N_2199,N_1583);
or U4815 (N_4815,N_2100,N_2473);
nor U4816 (N_4816,N_32,N_1401);
nor U4817 (N_4817,N_696,N_1430);
and U4818 (N_4818,N_2279,N_1574);
and U4819 (N_4819,N_792,N_655);
or U4820 (N_4820,N_2157,N_415);
and U4821 (N_4821,N_101,N_2134);
or U4822 (N_4822,N_1113,N_1915);
and U4823 (N_4823,N_287,N_121);
nand U4824 (N_4824,N_3,N_183);
nor U4825 (N_4825,N_1380,N_2430);
or U4826 (N_4826,N_2103,N_2355);
nor U4827 (N_4827,N_2487,N_1497);
nand U4828 (N_4828,N_504,N_258);
nor U4829 (N_4829,N_279,N_510);
nand U4830 (N_4830,N_2036,N_1791);
and U4831 (N_4831,N_1195,N_1358);
nand U4832 (N_4832,N_1568,N_1673);
xnor U4833 (N_4833,N_256,N_738);
xor U4834 (N_4834,N_1972,N_217);
nor U4835 (N_4835,N_906,N_550);
and U4836 (N_4836,N_1713,N_569);
nor U4837 (N_4837,N_565,N_569);
xnor U4838 (N_4838,N_74,N_1200);
or U4839 (N_4839,N_704,N_1107);
and U4840 (N_4840,N_2269,N_2347);
and U4841 (N_4841,N_674,N_301);
nor U4842 (N_4842,N_1152,N_1202);
nor U4843 (N_4843,N_360,N_2099);
or U4844 (N_4844,N_2231,N_1336);
and U4845 (N_4845,N_1877,N_2400);
and U4846 (N_4846,N_1847,N_1412);
nand U4847 (N_4847,N_1500,N_2190);
or U4848 (N_4848,N_986,N_1033);
or U4849 (N_4849,N_460,N_572);
and U4850 (N_4850,N_1451,N_292);
or U4851 (N_4851,N_302,N_757);
and U4852 (N_4852,N_531,N_2489);
or U4853 (N_4853,N_1936,N_1630);
and U4854 (N_4854,N_870,N_22);
and U4855 (N_4855,N_350,N_1621);
and U4856 (N_4856,N_270,N_560);
and U4857 (N_4857,N_2344,N_629);
or U4858 (N_4858,N_1280,N_407);
xnor U4859 (N_4859,N_483,N_1202);
nor U4860 (N_4860,N_1887,N_1259);
and U4861 (N_4861,N_1496,N_592);
and U4862 (N_4862,N_341,N_606);
nor U4863 (N_4863,N_1027,N_1822);
nor U4864 (N_4864,N_549,N_425);
nand U4865 (N_4865,N_824,N_1052);
or U4866 (N_4866,N_2240,N_1431);
nor U4867 (N_4867,N_1687,N_741);
nand U4868 (N_4868,N_1709,N_820);
nand U4869 (N_4869,N_1976,N_1592);
or U4870 (N_4870,N_1003,N_1719);
xor U4871 (N_4871,N_305,N_2330);
nand U4872 (N_4872,N_539,N_1034);
xor U4873 (N_4873,N_1090,N_568);
and U4874 (N_4874,N_1586,N_2269);
xnor U4875 (N_4875,N_1509,N_522);
nor U4876 (N_4876,N_626,N_1853);
xor U4877 (N_4877,N_72,N_2410);
nand U4878 (N_4878,N_2447,N_1287);
nor U4879 (N_4879,N_458,N_454);
and U4880 (N_4880,N_1134,N_282);
nand U4881 (N_4881,N_1722,N_507);
nor U4882 (N_4882,N_84,N_1559);
nor U4883 (N_4883,N_2130,N_191);
nor U4884 (N_4884,N_507,N_1389);
and U4885 (N_4885,N_1287,N_1352);
or U4886 (N_4886,N_2162,N_112);
or U4887 (N_4887,N_2019,N_2464);
nand U4888 (N_4888,N_593,N_1722);
and U4889 (N_4889,N_2076,N_1225);
xnor U4890 (N_4890,N_1732,N_1098);
nand U4891 (N_4891,N_1759,N_1813);
or U4892 (N_4892,N_1357,N_2312);
and U4893 (N_4893,N_750,N_2094);
nand U4894 (N_4894,N_2482,N_568);
or U4895 (N_4895,N_1929,N_2121);
or U4896 (N_4896,N_899,N_2463);
nor U4897 (N_4897,N_780,N_368);
and U4898 (N_4898,N_1630,N_1816);
nor U4899 (N_4899,N_548,N_1495);
nor U4900 (N_4900,N_1604,N_1754);
and U4901 (N_4901,N_1867,N_1461);
xnor U4902 (N_4902,N_1780,N_1557);
and U4903 (N_4903,N_937,N_684);
nand U4904 (N_4904,N_120,N_543);
or U4905 (N_4905,N_515,N_149);
nor U4906 (N_4906,N_1005,N_1469);
nor U4907 (N_4907,N_820,N_1480);
nor U4908 (N_4908,N_922,N_1720);
nand U4909 (N_4909,N_196,N_2289);
nor U4910 (N_4910,N_328,N_1609);
nand U4911 (N_4911,N_2089,N_710);
nand U4912 (N_4912,N_2331,N_1065);
and U4913 (N_4913,N_1941,N_1208);
nand U4914 (N_4914,N_2201,N_16);
and U4915 (N_4915,N_197,N_775);
xnor U4916 (N_4916,N_293,N_2129);
xnor U4917 (N_4917,N_203,N_1196);
or U4918 (N_4918,N_2410,N_1212);
nor U4919 (N_4919,N_776,N_65);
nand U4920 (N_4920,N_2239,N_2218);
nand U4921 (N_4921,N_59,N_1493);
xnor U4922 (N_4922,N_2350,N_2067);
and U4923 (N_4923,N_2035,N_642);
and U4924 (N_4924,N_2157,N_754);
nand U4925 (N_4925,N_2050,N_1673);
and U4926 (N_4926,N_1758,N_317);
nor U4927 (N_4927,N_1555,N_1954);
and U4928 (N_4928,N_1207,N_489);
or U4929 (N_4929,N_1407,N_618);
or U4930 (N_4930,N_504,N_95);
nand U4931 (N_4931,N_1682,N_1538);
nor U4932 (N_4932,N_110,N_1307);
nand U4933 (N_4933,N_1335,N_544);
and U4934 (N_4934,N_2356,N_1928);
or U4935 (N_4935,N_1489,N_2126);
and U4936 (N_4936,N_1265,N_1579);
nand U4937 (N_4937,N_55,N_686);
and U4938 (N_4938,N_1054,N_1835);
nand U4939 (N_4939,N_1514,N_269);
and U4940 (N_4940,N_1321,N_2275);
and U4941 (N_4941,N_1355,N_589);
or U4942 (N_4942,N_677,N_1139);
nand U4943 (N_4943,N_1552,N_2026);
xor U4944 (N_4944,N_691,N_1549);
or U4945 (N_4945,N_844,N_960);
xnor U4946 (N_4946,N_789,N_339);
xor U4947 (N_4947,N_1291,N_25);
or U4948 (N_4948,N_2304,N_2135);
nor U4949 (N_4949,N_1084,N_1670);
and U4950 (N_4950,N_714,N_1321);
or U4951 (N_4951,N_1301,N_1961);
xor U4952 (N_4952,N_1837,N_1223);
or U4953 (N_4953,N_794,N_630);
or U4954 (N_4954,N_785,N_272);
nor U4955 (N_4955,N_69,N_1576);
nand U4956 (N_4956,N_2037,N_1865);
nor U4957 (N_4957,N_1795,N_248);
or U4958 (N_4958,N_630,N_1900);
or U4959 (N_4959,N_898,N_933);
nand U4960 (N_4960,N_2416,N_710);
nand U4961 (N_4961,N_133,N_1161);
or U4962 (N_4962,N_854,N_1646);
or U4963 (N_4963,N_921,N_1549);
nand U4964 (N_4964,N_1229,N_418);
nand U4965 (N_4965,N_1848,N_1981);
and U4966 (N_4966,N_1066,N_1220);
or U4967 (N_4967,N_498,N_2414);
nor U4968 (N_4968,N_15,N_502);
nand U4969 (N_4969,N_2178,N_9);
or U4970 (N_4970,N_1449,N_2158);
and U4971 (N_4971,N_122,N_1375);
and U4972 (N_4972,N_666,N_64);
nand U4973 (N_4973,N_2492,N_609);
nand U4974 (N_4974,N_2025,N_512);
or U4975 (N_4975,N_579,N_1664);
or U4976 (N_4976,N_881,N_1744);
or U4977 (N_4977,N_647,N_1478);
nand U4978 (N_4978,N_1420,N_1998);
and U4979 (N_4979,N_1824,N_236);
xor U4980 (N_4980,N_1958,N_2222);
xor U4981 (N_4981,N_1155,N_1460);
or U4982 (N_4982,N_669,N_817);
and U4983 (N_4983,N_1405,N_1098);
nand U4984 (N_4984,N_764,N_756);
nand U4985 (N_4985,N_1451,N_325);
and U4986 (N_4986,N_1342,N_1375);
or U4987 (N_4987,N_318,N_842);
xor U4988 (N_4988,N_263,N_321);
or U4989 (N_4989,N_113,N_743);
or U4990 (N_4990,N_2182,N_1026);
or U4991 (N_4991,N_2057,N_464);
nand U4992 (N_4992,N_1041,N_1404);
and U4993 (N_4993,N_1838,N_919);
and U4994 (N_4994,N_1937,N_1590);
or U4995 (N_4995,N_247,N_948);
nor U4996 (N_4996,N_181,N_1903);
nand U4997 (N_4997,N_1261,N_1919);
and U4998 (N_4998,N_2422,N_1999);
nor U4999 (N_4999,N_958,N_1199);
or U5000 (N_5000,N_3651,N_3333);
nor U5001 (N_5001,N_4046,N_3457);
nor U5002 (N_5002,N_4562,N_4846);
xor U5003 (N_5003,N_3421,N_3143);
or U5004 (N_5004,N_4711,N_3385);
nor U5005 (N_5005,N_4309,N_4844);
xor U5006 (N_5006,N_4585,N_4918);
nand U5007 (N_5007,N_4950,N_4411);
nor U5008 (N_5008,N_4869,N_3928);
xnor U5009 (N_5009,N_4390,N_2926);
nand U5010 (N_5010,N_3717,N_4089);
or U5011 (N_5011,N_3970,N_3334);
nand U5012 (N_5012,N_2870,N_4777);
nor U5013 (N_5013,N_3695,N_4349);
or U5014 (N_5014,N_3559,N_3590);
or U5015 (N_5015,N_4468,N_4454);
nand U5016 (N_5016,N_3686,N_3829);
or U5017 (N_5017,N_4868,N_3026);
nand U5018 (N_5018,N_3544,N_3068);
xor U5019 (N_5019,N_4507,N_2877);
or U5020 (N_5020,N_4009,N_4624);
nand U5021 (N_5021,N_3029,N_2673);
nand U5022 (N_5022,N_4016,N_3360);
and U5023 (N_5023,N_3800,N_2928);
or U5024 (N_5024,N_3512,N_3546);
or U5025 (N_5025,N_3934,N_4266);
or U5026 (N_5026,N_4200,N_3950);
and U5027 (N_5027,N_4901,N_4516);
and U5028 (N_5028,N_4322,N_3203);
nor U5029 (N_5029,N_3035,N_4775);
nand U5030 (N_5030,N_3424,N_3657);
and U5031 (N_5031,N_2572,N_4884);
nor U5032 (N_5032,N_3084,N_4938);
and U5033 (N_5033,N_3428,N_4772);
nor U5034 (N_5034,N_3151,N_4874);
or U5035 (N_5035,N_4958,N_3471);
or U5036 (N_5036,N_2895,N_2545);
nor U5037 (N_5037,N_3407,N_4651);
or U5038 (N_5038,N_3045,N_4972);
or U5039 (N_5039,N_3230,N_2754);
nand U5040 (N_5040,N_4665,N_3804);
nand U5041 (N_5041,N_2610,N_3850);
or U5042 (N_5042,N_4098,N_2621);
and U5043 (N_5043,N_4133,N_4378);
and U5044 (N_5044,N_2938,N_4000);
and U5045 (N_5045,N_4925,N_3410);
nor U5046 (N_5046,N_2683,N_2562);
nand U5047 (N_5047,N_4881,N_4426);
or U5048 (N_5048,N_3898,N_3274);
nand U5049 (N_5049,N_2514,N_4629);
nand U5050 (N_5050,N_3117,N_4243);
nand U5051 (N_5051,N_4337,N_3614);
or U5052 (N_5052,N_2645,N_3925);
nand U5053 (N_5053,N_2910,N_4823);
nor U5054 (N_5054,N_3320,N_3364);
nor U5055 (N_5055,N_2540,N_3915);
and U5056 (N_5056,N_4916,N_3005);
nor U5057 (N_5057,N_2639,N_2699);
nor U5058 (N_5058,N_4939,N_4835);
nor U5059 (N_5059,N_3636,N_4499);
and U5060 (N_5060,N_4091,N_3622);
nand U5061 (N_5061,N_2724,N_4843);
and U5062 (N_5062,N_2833,N_2966);
and U5063 (N_5063,N_4635,N_4371);
or U5064 (N_5064,N_4857,N_4415);
and U5065 (N_5065,N_3818,N_3705);
nor U5066 (N_5066,N_4431,N_4077);
nor U5067 (N_5067,N_4804,N_4928);
or U5068 (N_5068,N_3855,N_4943);
and U5069 (N_5069,N_3841,N_4376);
and U5070 (N_5070,N_4080,N_3699);
nor U5071 (N_5071,N_4936,N_3535);
nand U5072 (N_5072,N_2842,N_3191);
and U5073 (N_5073,N_2764,N_4787);
nand U5074 (N_5074,N_2618,N_2819);
nand U5075 (N_5075,N_4970,N_4304);
and U5076 (N_5076,N_3980,N_4754);
or U5077 (N_5077,N_4441,N_4050);
nor U5078 (N_5078,N_2729,N_2635);
nand U5079 (N_5079,N_3213,N_3234);
and U5080 (N_5080,N_4439,N_3924);
nand U5081 (N_5081,N_3401,N_4265);
nor U5082 (N_5082,N_3777,N_4871);
or U5083 (N_5083,N_3399,N_4842);
nor U5084 (N_5084,N_2971,N_3408);
or U5085 (N_5085,N_3397,N_2711);
and U5086 (N_5086,N_2933,N_3779);
nor U5087 (N_5087,N_4234,N_4527);
nor U5088 (N_5088,N_3135,N_3157);
nor U5089 (N_5089,N_4433,N_2919);
and U5090 (N_5090,N_3437,N_3991);
nand U5091 (N_5091,N_4708,N_3724);
and U5092 (N_5092,N_4087,N_4644);
and U5093 (N_5093,N_3888,N_4501);
xnor U5094 (N_5094,N_3957,N_4677);
xor U5095 (N_5095,N_4386,N_2553);
nand U5096 (N_5096,N_4953,N_4668);
xor U5097 (N_5097,N_3171,N_2978);
or U5098 (N_5098,N_2896,N_4765);
and U5099 (N_5099,N_3944,N_4097);
xor U5100 (N_5100,N_2583,N_3581);
and U5101 (N_5101,N_3530,N_3478);
and U5102 (N_5102,N_2801,N_2828);
nand U5103 (N_5103,N_4167,N_2740);
or U5104 (N_5104,N_4774,N_3186);
or U5105 (N_5105,N_2948,N_2998);
or U5106 (N_5106,N_3498,N_2722);
and U5107 (N_5107,N_4258,N_3048);
or U5108 (N_5108,N_4510,N_3264);
or U5109 (N_5109,N_3880,N_4450);
xnor U5110 (N_5110,N_3570,N_4839);
and U5111 (N_5111,N_4028,N_2759);
or U5112 (N_5112,N_2875,N_4191);
nor U5113 (N_5113,N_3795,N_3731);
nand U5114 (N_5114,N_4422,N_3612);
xnor U5115 (N_5115,N_3433,N_3150);
or U5116 (N_5116,N_4180,N_3525);
xor U5117 (N_5117,N_2911,N_4546);
nand U5118 (N_5118,N_3484,N_3147);
and U5119 (N_5119,N_4382,N_4241);
nor U5120 (N_5120,N_3069,N_4989);
nor U5121 (N_5121,N_3932,N_2761);
and U5122 (N_5122,N_3582,N_3736);
and U5123 (N_5123,N_4333,N_4713);
nand U5124 (N_5124,N_3403,N_4866);
and U5125 (N_5125,N_4902,N_2524);
and U5126 (N_5126,N_2560,N_3776);
and U5127 (N_5127,N_4566,N_2602);
or U5128 (N_5128,N_3825,N_2772);
and U5129 (N_5129,N_3439,N_4075);
and U5130 (N_5130,N_4800,N_3466);
and U5131 (N_5131,N_3485,N_4538);
or U5132 (N_5132,N_2899,N_2892);
or U5133 (N_5133,N_3893,N_4025);
or U5134 (N_5134,N_2791,N_3609);
nor U5135 (N_5135,N_4654,N_4303);
or U5136 (N_5136,N_3543,N_3493);
nor U5137 (N_5137,N_2682,N_3761);
nor U5138 (N_5138,N_4421,N_4791);
and U5139 (N_5139,N_4622,N_2613);
nor U5140 (N_5140,N_4963,N_2665);
or U5141 (N_5141,N_4617,N_4803);
nand U5142 (N_5142,N_4306,N_4325);
and U5143 (N_5143,N_4008,N_3221);
xor U5144 (N_5144,N_2605,N_3383);
and U5145 (N_5145,N_4537,N_4455);
and U5146 (N_5146,N_4771,N_2537);
and U5147 (N_5147,N_4412,N_4590);
or U5148 (N_5148,N_4108,N_4400);
or U5149 (N_5149,N_3946,N_2717);
nor U5150 (N_5150,N_3853,N_2719);
and U5151 (N_5151,N_2557,N_4014);
xor U5152 (N_5152,N_2686,N_4512);
nor U5153 (N_5153,N_4825,N_3159);
xor U5154 (N_5154,N_4039,N_4559);
or U5155 (N_5155,N_4619,N_4892);
and U5156 (N_5156,N_3895,N_2783);
nor U5157 (N_5157,N_4710,N_4814);
nor U5158 (N_5158,N_3820,N_4033);
nand U5159 (N_5159,N_4305,N_3345);
nor U5160 (N_5160,N_4345,N_3844);
and U5161 (N_5161,N_2871,N_2932);
xor U5162 (N_5162,N_3205,N_4608);
nand U5163 (N_5163,N_4886,N_3426);
nor U5164 (N_5164,N_4784,N_3375);
nand U5165 (N_5165,N_3577,N_3318);
nand U5166 (N_5166,N_4885,N_4639);
nand U5167 (N_5167,N_2677,N_3951);
or U5168 (N_5168,N_3311,N_3630);
nor U5169 (N_5169,N_3256,N_2579);
nand U5170 (N_5170,N_4905,N_3259);
nand U5171 (N_5171,N_3587,N_3303);
and U5172 (N_5172,N_2632,N_4976);
and U5173 (N_5173,N_4796,N_3227);
or U5174 (N_5174,N_4385,N_3859);
nor U5175 (N_5175,N_4658,N_3286);
nor U5176 (N_5176,N_4142,N_3109);
nand U5177 (N_5177,N_3769,N_3835);
and U5178 (N_5178,N_2817,N_3631);
and U5179 (N_5179,N_4145,N_2771);
nor U5180 (N_5180,N_4579,N_4863);
nand U5181 (N_5181,N_4352,N_4383);
nor U5182 (N_5182,N_3642,N_4096);
nand U5183 (N_5183,N_3142,N_2561);
or U5184 (N_5184,N_2917,N_3955);
or U5185 (N_5185,N_4432,N_2853);
xor U5186 (N_5186,N_4270,N_3673);
nor U5187 (N_5187,N_3066,N_2977);
or U5188 (N_5188,N_4340,N_4286);
xnor U5189 (N_5189,N_4144,N_2789);
or U5190 (N_5190,N_2884,N_3499);
nand U5191 (N_5191,N_4474,N_4214);
and U5192 (N_5192,N_4808,N_3353);
and U5193 (N_5193,N_3575,N_3672);
or U5194 (N_5194,N_4114,N_3542);
nand U5195 (N_5195,N_4111,N_4427);
or U5196 (N_5196,N_4914,N_3237);
nand U5197 (N_5197,N_3658,N_2799);
or U5198 (N_5198,N_4120,N_2504);
nor U5199 (N_5199,N_3821,N_3112);
xnor U5200 (N_5200,N_4969,N_4170);
xnor U5201 (N_5201,N_2947,N_3700);
nor U5202 (N_5202,N_3899,N_4079);
or U5203 (N_5203,N_3819,N_4653);
and U5204 (N_5204,N_3046,N_4947);
or U5205 (N_5205,N_2972,N_3669);
nand U5206 (N_5206,N_3156,N_3453);
and U5207 (N_5207,N_3146,N_4567);
and U5208 (N_5208,N_3101,N_3121);
and U5209 (N_5209,N_4504,N_4154);
nor U5210 (N_5210,N_3462,N_4946);
and U5211 (N_5211,N_3794,N_3200);
xnor U5212 (N_5212,N_4311,N_4209);
nand U5213 (N_5213,N_2784,N_3172);
or U5214 (N_5214,N_3624,N_3459);
and U5215 (N_5215,N_3852,N_4931);
nor U5216 (N_5216,N_4864,N_4380);
nand U5217 (N_5217,N_3976,N_4374);
nand U5218 (N_5218,N_3877,N_3185);
or U5219 (N_5219,N_2873,N_3770);
nor U5220 (N_5220,N_4147,N_3414);
and U5221 (N_5221,N_3192,N_3929);
nand U5222 (N_5222,N_4794,N_4563);
xnor U5223 (N_5223,N_4093,N_2694);
and U5224 (N_5224,N_3762,N_3655);
nor U5225 (N_5225,N_3640,N_3248);
nor U5226 (N_5226,N_2860,N_3404);
xnor U5227 (N_5227,N_4656,N_4263);
nor U5228 (N_5228,N_2646,N_4148);
xor U5229 (N_5229,N_3718,N_4109);
and U5230 (N_5230,N_3436,N_4485);
nand U5231 (N_5231,N_4910,N_4235);
nor U5232 (N_5232,N_3774,N_4778);
and U5233 (N_5233,N_2953,N_4528);
xnor U5234 (N_5234,N_2538,N_3273);
and U5235 (N_5235,N_4381,N_4712);
xor U5236 (N_5236,N_4059,N_3197);
nand U5237 (N_5237,N_3400,N_4420);
or U5238 (N_5238,N_3638,N_3782);
nor U5239 (N_5239,N_3301,N_4460);
nand U5240 (N_5240,N_4944,N_3801);
nor U5241 (N_5241,N_3552,N_4188);
xnor U5242 (N_5242,N_4113,N_2924);
or U5243 (N_5243,N_4288,N_4475);
xnor U5244 (N_5244,N_2575,N_3492);
nand U5245 (N_5245,N_3793,N_4466);
nand U5246 (N_5246,N_2564,N_3506);
and U5247 (N_5247,N_2937,N_2643);
nand U5248 (N_5248,N_4082,N_4092);
nand U5249 (N_5249,N_4321,N_4802);
and U5250 (N_5250,N_2957,N_4599);
nand U5251 (N_5251,N_3441,N_3519);
or U5252 (N_5252,N_4893,N_3323);
nor U5253 (N_5253,N_4756,N_3927);
nand U5254 (N_5254,N_4078,N_3534);
or U5255 (N_5255,N_3677,N_2940);
nor U5256 (N_5256,N_4999,N_3827);
and U5257 (N_5257,N_3602,N_4663);
nor U5258 (N_5258,N_3584,N_4903);
nand U5259 (N_5259,N_3966,N_4026);
nor U5260 (N_5260,N_2970,N_4519);
or U5261 (N_5261,N_4573,N_4671);
nor U5262 (N_5262,N_3984,N_4511);
or U5263 (N_5263,N_4965,N_4094);
or U5264 (N_5264,N_4535,N_3707);
xor U5265 (N_5265,N_2531,N_2725);
nor U5266 (N_5266,N_2727,N_2865);
nand U5267 (N_5267,N_3971,N_3565);
or U5268 (N_5268,N_2925,N_2747);
and U5269 (N_5269,N_2834,N_2796);
xor U5270 (N_5270,N_2787,N_4291);
nand U5271 (N_5271,N_3742,N_4469);
and U5272 (N_5272,N_4012,N_4126);
nor U5273 (N_5273,N_4399,N_4967);
and U5274 (N_5274,N_3016,N_3784);
nand U5275 (N_5275,N_3632,N_3646);
nor U5276 (N_5276,N_3785,N_3247);
nor U5277 (N_5277,N_3983,N_2608);
and U5278 (N_5278,N_4642,N_4542);
xor U5279 (N_5279,N_2768,N_2567);
or U5280 (N_5280,N_4926,N_2521);
or U5281 (N_5281,N_4506,N_2659);
nand U5282 (N_5282,N_3743,N_4860);
and U5283 (N_5283,N_4490,N_4733);
nor U5284 (N_5284,N_4156,N_4621);
nand U5285 (N_5285,N_4201,N_3733);
nand U5286 (N_5286,N_4586,N_4995);
nor U5287 (N_5287,N_3253,N_4979);
nor U5288 (N_5288,N_4312,N_2958);
nand U5289 (N_5289,N_3716,N_4202);
nor U5290 (N_5290,N_4837,N_4011);
nor U5291 (N_5291,N_3154,N_3729);
or U5292 (N_5292,N_4690,N_4701);
nand U5293 (N_5293,N_4678,N_3219);
and U5294 (N_5294,N_3365,N_4865);
xnor U5295 (N_5295,N_4888,N_2611);
xor U5296 (N_5296,N_3475,N_3326);
nand U5297 (N_5297,N_3442,N_3232);
and U5298 (N_5298,N_4206,N_3900);
nand U5299 (N_5299,N_2775,N_2532);
or U5300 (N_5300,N_4254,N_4081);
nor U5301 (N_5301,N_4323,N_4006);
nor U5302 (N_5302,N_4205,N_3910);
or U5303 (N_5303,N_3596,N_3148);
or U5304 (N_5304,N_4673,N_3454);
or U5305 (N_5305,N_4363,N_4521);
or U5306 (N_5306,N_3313,N_4676);
nand U5307 (N_5307,N_2617,N_3920);
xor U5308 (N_5308,N_4744,N_3430);
and U5309 (N_5309,N_3759,N_4149);
xnor U5310 (N_5310,N_4034,N_3260);
nand U5311 (N_5311,N_4375,N_3134);
and U5312 (N_5312,N_2695,N_2507);
nor U5313 (N_5313,N_3509,N_3997);
or U5314 (N_5314,N_3124,N_2951);
xor U5315 (N_5315,N_4102,N_4410);
and U5316 (N_5316,N_2590,N_3017);
nor U5317 (N_5317,N_4010,N_2546);
nand U5318 (N_5318,N_2806,N_2704);
and U5319 (N_5319,N_3494,N_2949);
or U5320 (N_5320,N_2767,N_3141);
nand U5321 (N_5321,N_3398,N_4799);
or U5322 (N_5322,N_4699,N_4020);
nor U5323 (N_5323,N_3078,N_3711);
xnor U5324 (N_5324,N_2793,N_4334);
and U5325 (N_5325,N_4623,N_3495);
nand U5326 (N_5326,N_3238,N_4829);
or U5327 (N_5327,N_3905,N_4135);
nor U5328 (N_5328,N_4734,N_4072);
nor U5329 (N_5329,N_3958,N_4841);
xnor U5330 (N_5330,N_4341,N_4290);
nor U5331 (N_5331,N_4786,N_2558);
xnor U5332 (N_5332,N_2968,N_4130);
nand U5333 (N_5333,N_3090,N_2522);
nand U5334 (N_5334,N_3336,N_2890);
and U5335 (N_5335,N_2751,N_2520);
or U5336 (N_5336,N_2755,N_3158);
nand U5337 (N_5337,N_2660,N_3889);
or U5338 (N_5338,N_4347,N_2519);
nor U5339 (N_5339,N_2689,N_3972);
or U5340 (N_5340,N_4740,N_3790);
nor U5341 (N_5341,N_3954,N_2889);
nand U5342 (N_5342,N_3993,N_3805);
nand U5343 (N_5343,N_4704,N_4223);
or U5344 (N_5344,N_3826,N_4486);
nor U5345 (N_5345,N_4463,N_3223);
nor U5346 (N_5346,N_3050,N_2541);
nor U5347 (N_5347,N_4143,N_4489);
or U5348 (N_5348,N_2855,N_3131);
or U5349 (N_5349,N_2581,N_3222);
nand U5350 (N_5350,N_3366,N_3515);
xor U5351 (N_5351,N_3487,N_3254);
nand U5352 (N_5352,N_4549,N_4358);
xor U5353 (N_5353,N_2996,N_2526);
or U5354 (N_5354,N_2941,N_3110);
or U5355 (N_5355,N_3797,N_3434);
or U5356 (N_5356,N_4880,N_4032);
or U5357 (N_5357,N_4998,N_3873);
nand U5358 (N_5358,N_3680,N_4178);
or U5359 (N_5359,N_3178,N_3276);
xor U5360 (N_5360,N_4879,N_3257);
nand U5361 (N_5361,N_4123,N_4187);
nor U5362 (N_5362,N_4416,N_2511);
and U5363 (N_5363,N_4913,N_2624);
nand U5364 (N_5364,N_3338,N_2628);
nand U5365 (N_5365,N_4759,N_3295);
nand U5366 (N_5366,N_4895,N_3176);
and U5367 (N_5367,N_3059,N_3604);
nor U5368 (N_5368,N_4850,N_4346);
or U5369 (N_5369,N_2987,N_2650);
nor U5370 (N_5370,N_2509,N_3754);
and U5371 (N_5371,N_4933,N_3942);
and U5372 (N_5372,N_3479,N_3560);
and U5373 (N_5373,N_4483,N_4184);
nand U5374 (N_5374,N_3569,N_3714);
and U5375 (N_5375,N_3752,N_3181);
or U5376 (N_5376,N_3740,N_4961);
or U5377 (N_5377,N_4199,N_4021);
nor U5378 (N_5378,N_3860,N_3637);
nand U5379 (N_5379,N_3449,N_2837);
nand U5380 (N_5380,N_4652,N_4056);
nor U5381 (N_5381,N_3753,N_2534);
or U5382 (N_5382,N_3396,N_2942);
or U5383 (N_5383,N_4981,N_3628);
nor U5384 (N_5384,N_3662,N_4480);
nor U5385 (N_5385,N_3550,N_3362);
or U5386 (N_5386,N_3173,N_3335);
or U5387 (N_5387,N_3874,N_2742);
and U5388 (N_5388,N_3576,N_3974);
xor U5389 (N_5389,N_4366,N_4132);
nor U5390 (N_5390,N_4887,N_3981);
xnor U5391 (N_5391,N_4153,N_2915);
nor U5392 (N_5392,N_3262,N_3593);
nor U5393 (N_5393,N_3079,N_3890);
and U5394 (N_5394,N_3568,N_3541);
nand U5395 (N_5395,N_4987,N_2706);
and U5396 (N_5396,N_4508,N_4447);
and U5397 (N_5397,N_4851,N_4398);
nand U5398 (N_5398,N_2914,N_4196);
nor U5399 (N_5399,N_3216,N_4137);
nor U5400 (N_5400,N_3242,N_4449);
nand U5401 (N_5401,N_4182,N_4788);
nand U5402 (N_5402,N_4458,N_3869);
nor U5403 (N_5403,N_4437,N_4686);
and U5404 (N_5404,N_4604,N_4878);
nand U5405 (N_5405,N_4634,N_4588);
nor U5406 (N_5406,N_4577,N_2832);
nor U5407 (N_5407,N_3763,N_4747);
or U5408 (N_5408,N_3463,N_4237);
nor U5409 (N_5409,N_2908,N_4095);
nor U5410 (N_5410,N_4236,N_4282);
xor U5411 (N_5411,N_3432,N_3020);
xnor U5412 (N_5412,N_2840,N_4581);
nor U5413 (N_5413,N_2597,N_3160);
nor U5414 (N_5414,N_3300,N_4707);
and U5415 (N_5415,N_4018,N_2991);
nand U5416 (N_5416,N_4889,N_4780);
nand U5417 (N_5417,N_4986,N_2636);
or U5418 (N_5418,N_4146,N_4664);
nor U5419 (N_5419,N_2735,N_3083);
nor U5420 (N_5420,N_3663,N_4662);
nor U5421 (N_5421,N_4929,N_4361);
and U5422 (N_5422,N_3374,N_4273);
nand U5423 (N_5423,N_3133,N_4299);
and U5424 (N_5424,N_4732,N_4877);
nand U5425 (N_5425,N_3088,N_4225);
nor U5426 (N_5426,N_4934,N_3634);
or U5427 (N_5427,N_4891,N_3412);
and U5428 (N_5428,N_2863,N_2529);
and U5429 (N_5429,N_4849,N_3698);
and U5430 (N_5430,N_4105,N_3049);
nand U5431 (N_5431,N_3988,N_3817);
nor U5432 (N_5432,N_3583,N_4620);
nor U5433 (N_5433,N_4308,N_3644);
or U5434 (N_5434,N_3545,N_3709);
nor U5435 (N_5435,N_4957,N_4425);
xor U5436 (N_5436,N_4536,N_3025);
and U5437 (N_5437,N_2739,N_4365);
and U5438 (N_5438,N_4601,N_4189);
and U5439 (N_5439,N_4436,N_3706);
or U5440 (N_5440,N_3526,N_3588);
nor U5441 (N_5441,N_3182,N_2843);
or U5442 (N_5442,N_3708,N_2571);
nand U5443 (N_5443,N_4831,N_3688);
or U5444 (N_5444,N_2765,N_4391);
nor U5445 (N_5445,N_3574,N_2599);
and U5446 (N_5446,N_4730,N_4388);
or U5447 (N_5447,N_3091,N_3660);
xnor U5448 (N_5448,N_2716,N_2703);
and U5449 (N_5449,N_4945,N_2777);
or U5450 (N_5450,N_2838,N_4280);
or U5451 (N_5451,N_4495,N_4743);
or U5452 (N_5452,N_4948,N_3551);
or U5453 (N_5453,N_3845,N_2993);
nor U5454 (N_5454,N_4140,N_3690);
and U5455 (N_5455,N_3977,N_2912);
nor U5456 (N_5456,N_2651,N_4515);
and U5457 (N_5457,N_4792,N_4429);
or U5458 (N_5458,N_3828,N_2693);
or U5459 (N_5459,N_4768,N_4328);
nor U5460 (N_5460,N_3358,N_2634);
nor U5461 (N_5461,N_3780,N_3803);
nand U5462 (N_5462,N_3591,N_3833);
or U5463 (N_5463,N_3447,N_3299);
and U5464 (N_5464,N_3746,N_3390);
or U5465 (N_5465,N_4830,N_4240);
xor U5466 (N_5466,N_3979,N_3039);
or U5467 (N_5467,N_2672,N_2866);
nor U5468 (N_5468,N_4257,N_4524);
or U5469 (N_5469,N_4127,N_2633);
or U5470 (N_5470,N_4749,N_3936);
and U5471 (N_5471,N_2615,N_4338);
nand U5472 (N_5472,N_4007,N_4221);
nor U5473 (N_5473,N_3015,N_3246);
nand U5474 (N_5474,N_3347,N_4339);
nand U5475 (N_5475,N_3193,N_4023);
or U5476 (N_5476,N_4529,N_4174);
and U5477 (N_5477,N_2829,N_4279);
and U5478 (N_5478,N_4591,N_4824);
nand U5479 (N_5479,N_4044,N_3962);
nand U5480 (N_5480,N_2578,N_4071);
nand U5481 (N_5481,N_3194,N_3665);
and U5482 (N_5482,N_2861,N_4683);
and U5483 (N_5483,N_3667,N_4319);
or U5484 (N_5484,N_4310,N_3085);
nor U5485 (N_5485,N_2800,N_3639);
nor U5486 (N_5486,N_3382,N_4828);
and U5487 (N_5487,N_3118,N_4525);
and U5488 (N_5488,N_2654,N_2879);
and U5489 (N_5489,N_4053,N_4692);
nand U5490 (N_5490,N_3305,N_4232);
nor U5491 (N_5491,N_2516,N_4125);
or U5492 (N_5492,N_2967,N_4509);
nand U5493 (N_5493,N_3747,N_3792);
or U5494 (N_5494,N_3876,N_2781);
nand U5495 (N_5495,N_4875,N_4723);
nand U5496 (N_5496,N_4779,N_2535);
nor U5497 (N_5497,N_4335,N_2685);
or U5498 (N_5498,N_4896,N_3608);
and U5499 (N_5499,N_3419,N_3990);
nand U5500 (N_5500,N_3255,N_3174);
nand U5501 (N_5501,N_3995,N_2746);
and U5502 (N_5502,N_4065,N_2625);
nor U5503 (N_5503,N_4069,N_2988);
and U5504 (N_5504,N_4548,N_3813);
and U5505 (N_5505,N_3867,N_2588);
and U5506 (N_5506,N_3011,N_4575);
nor U5507 (N_5507,N_2700,N_3537);
xnor U5508 (N_5508,N_3019,N_3082);
nand U5509 (N_5509,N_3621,N_3031);
and U5510 (N_5510,N_2807,N_3540);
or U5511 (N_5511,N_4002,N_4716);
nand U5512 (N_5512,N_3389,N_3138);
nand U5513 (N_5513,N_3728,N_3571);
nand U5514 (N_5514,N_4870,N_3008);
nor U5515 (N_5515,N_2502,N_4742);
or U5516 (N_5516,N_2503,N_3796);
nor U5517 (N_5517,N_4327,N_3913);
nand U5518 (N_5518,N_2778,N_2670);
or U5519 (N_5519,N_3573,N_4909);
nand U5520 (N_5520,N_4853,N_3982);
nand U5521 (N_5521,N_2543,N_4259);
nor U5522 (N_5522,N_3661,N_2726);
or U5523 (N_5523,N_3947,N_2612);
and U5524 (N_5524,N_4674,N_3994);
and U5525 (N_5525,N_3184,N_2849);
and U5526 (N_5526,N_4370,N_4104);
xor U5527 (N_5527,N_3594,N_4186);
or U5528 (N_5528,N_3164,N_3380);
nand U5529 (N_5529,N_4856,N_3987);
nand U5530 (N_5530,N_4594,N_3822);
and U5531 (N_5531,N_2642,N_3938);
nand U5532 (N_5532,N_2687,N_4244);
and U5533 (N_5533,N_4171,N_2681);
or U5534 (N_5534,N_2517,N_3922);
nor U5535 (N_5535,N_3270,N_3070);
nand U5536 (N_5536,N_4767,N_4387);
or U5537 (N_5537,N_4066,N_3750);
xnor U5538 (N_5538,N_3676,N_4598);
and U5539 (N_5539,N_4960,N_4217);
nor U5540 (N_5540,N_4457,N_3616);
nor U5541 (N_5541,N_4074,N_3799);
nor U5542 (N_5542,N_3814,N_3952);
nor U5543 (N_5543,N_4956,N_2878);
nor U5544 (N_5544,N_2851,N_2823);
and U5545 (N_5545,N_3169,N_3963);
nand U5546 (N_5546,N_4100,N_3018);
nand U5547 (N_5547,N_4561,N_3309);
nand U5548 (N_5548,N_2986,N_3502);
or U5549 (N_5549,N_3882,N_2974);
nand U5550 (N_5550,N_4247,N_2850);
nand U5551 (N_5551,N_4988,N_4090);
or U5552 (N_5552,N_3370,N_4605);
nor U5553 (N_5553,N_2826,N_4776);
nand U5554 (N_5554,N_3119,N_4136);
nand U5555 (N_5555,N_4041,N_3038);
nor U5556 (N_5556,N_3357,N_3749);
or U5557 (N_5557,N_3100,N_4057);
or U5558 (N_5558,N_4239,N_4359);
nor U5559 (N_5559,N_2512,N_4165);
nor U5560 (N_5560,N_3330,N_2566);
and U5561 (N_5561,N_3563,N_2525);
nor U5562 (N_5562,N_4602,N_3477);
and U5563 (N_5563,N_4118,N_4966);
and U5564 (N_5564,N_4717,N_4099);
nor U5565 (N_5565,N_2528,N_2769);
nor U5566 (N_5566,N_2518,N_4351);
or U5567 (N_5567,N_4763,N_3218);
nor U5568 (N_5568,N_4637,N_3298);
or U5569 (N_5569,N_2607,N_4500);
nor U5570 (N_5570,N_3126,N_4445);
nand U5571 (N_5571,N_4724,N_3209);
or U5572 (N_5572,N_4295,N_3355);
and U5573 (N_5573,N_4547,N_2965);
nor U5574 (N_5574,N_4070,N_3975);
nand U5575 (N_5575,N_4596,N_2696);
or U5576 (N_5576,N_4294,N_4344);
or U5577 (N_5577,N_3332,N_3562);
and U5578 (N_5578,N_4818,N_2669);
nand U5579 (N_5579,N_4467,N_3180);
nand U5580 (N_5580,N_3871,N_3052);
nand U5581 (N_5581,N_3179,N_4532);
xnor U5582 (N_5582,N_2811,N_4811);
nand U5583 (N_5583,N_4405,N_2565);
xor U5584 (N_5584,N_2959,N_4316);
nand U5585 (N_5585,N_2818,N_4158);
or U5586 (N_5586,N_3294,N_4764);
nand U5587 (N_5587,N_4190,N_3539);
or U5588 (N_5588,N_3252,N_3415);
or U5589 (N_5589,N_4700,N_3317);
nand U5590 (N_5590,N_4694,N_2720);
and U5591 (N_5591,N_3271,N_2662);
and U5592 (N_5592,N_3099,N_2510);
or U5593 (N_5593,N_3229,N_4194);
nand U5594 (N_5594,N_4603,N_2620);
and U5595 (N_5595,N_3586,N_4177);
nand U5596 (N_5596,N_4503,N_4922);
or U5597 (N_5597,N_4715,N_2710);
nand U5598 (N_5598,N_3547,N_2582);
nor U5599 (N_5599,N_4657,N_2601);
or U5600 (N_5600,N_4397,N_4377);
or U5601 (N_5601,N_4954,N_3128);
nor U5602 (N_5602,N_3842,N_3863);
xor U5603 (N_5603,N_2556,N_4085);
xnor U5604 (N_5604,N_4583,N_3467);
nand U5605 (N_5605,N_3786,N_3903);
nand U5606 (N_5606,N_3054,N_4720);
or U5607 (N_5607,N_3346,N_4773);
or U5608 (N_5608,N_3445,N_4298);
and U5609 (N_5609,N_4633,N_2846);
nor U5610 (N_5610,N_4452,N_4448);
nor U5611 (N_5611,N_4753,N_3891);
nand U5612 (N_5612,N_4278,N_3372);
nor U5613 (N_5613,N_3491,N_4611);
nand U5614 (N_5614,N_2559,N_3775);
nor U5615 (N_5615,N_2712,N_3520);
nor U5616 (N_5616,N_3130,N_3812);
and U5617 (N_5617,N_3472,N_3549);
nor U5618 (N_5618,N_3137,N_3697);
or U5619 (N_5619,N_3514,N_3263);
and U5620 (N_5620,N_4962,N_3043);
nor U5621 (N_5621,N_4613,N_4248);
nand U5622 (N_5622,N_3967,N_3765);
and U5623 (N_5623,N_3369,N_4213);
nand U5624 (N_5624,N_3363,N_2982);
nor U5625 (N_5625,N_4899,N_4703);
nor U5626 (N_5626,N_3379,N_3340);
nor U5627 (N_5627,N_3339,N_2891);
nor U5628 (N_5628,N_4353,N_4628);
xnor U5629 (N_5629,N_2956,N_3014);
nor U5630 (N_5630,N_3719,N_2623);
and U5631 (N_5631,N_4434,N_3939);
and U5632 (N_5632,N_4872,N_4616);
or U5633 (N_5633,N_4894,N_4595);
xor U5634 (N_5634,N_4971,N_2805);
nor U5635 (N_5635,N_2939,N_3120);
nand U5636 (N_5636,N_4882,N_4840);
or U5637 (N_5637,N_3122,N_4540);
or U5638 (N_5638,N_3884,N_3196);
nand U5639 (N_5639,N_4526,N_2737);
and U5640 (N_5640,N_2595,N_2678);
or U5641 (N_5641,N_3042,N_4721);
nor U5642 (N_5642,N_2779,N_3376);
nor U5643 (N_5643,N_3766,N_4451);
nor U5644 (N_5644,N_4024,N_3236);
xnor U5645 (N_5645,N_4183,N_3411);
nand U5646 (N_5646,N_3647,N_4131);
or U5647 (N_5647,N_3883,N_4367);
and U5648 (N_5648,N_3107,N_3480);
or U5649 (N_5649,N_2973,N_3650);
xor U5650 (N_5650,N_2797,N_3585);
nand U5651 (N_5651,N_3165,N_3064);
nand U5652 (N_5652,N_3155,N_3715);
and U5653 (N_5653,N_3764,N_3033);
or U5654 (N_5654,N_4252,N_3072);
nor U5655 (N_5655,N_2952,N_4419);
nand U5656 (N_5656,N_3595,N_3189);
xnor U5657 (N_5657,N_4920,N_4181);
or U5658 (N_5658,N_4618,N_3808);
and U5659 (N_5659,N_3351,N_4645);
or U5660 (N_5660,N_3034,N_4275);
and U5661 (N_5661,N_3489,N_4912);
xnor U5662 (N_5662,N_3948,N_3075);
nor U5663 (N_5663,N_2714,N_4973);
and U5664 (N_5664,N_4481,N_2547);
nor U5665 (N_5665,N_2795,N_3003);
nand U5666 (N_5666,N_4330,N_2774);
nand U5667 (N_5667,N_3738,N_3843);
or U5668 (N_5668,N_4300,N_4042);
nor U5669 (N_5669,N_2897,N_2598);
nor U5670 (N_5670,N_2640,N_3104);
xnor U5671 (N_5671,N_3002,N_4937);
and U5672 (N_5672,N_4578,N_2585);
nor U5673 (N_5673,N_4543,N_3831);
or U5674 (N_5674,N_2905,N_3001);
nor U5675 (N_5675,N_4470,N_4264);
or U5676 (N_5676,N_4175,N_2707);
nor U5677 (N_5677,N_4406,N_4318);
and U5678 (N_5678,N_4836,N_3956);
or U5679 (N_5679,N_3327,N_3522);
xnor U5680 (N_5680,N_4822,N_4758);
and U5681 (N_5681,N_4783,N_4952);
nor U5682 (N_5682,N_4977,N_3249);
or U5683 (N_5683,N_3422,N_4428);
xnor U5684 (N_5684,N_4782,N_3840);
nand U5685 (N_5685,N_3720,N_4687);
and U5686 (N_5686,N_4348,N_3513);
nor U5687 (N_5687,N_2616,N_4393);
nor U5688 (N_5688,N_4906,N_2921);
xor U5689 (N_5689,N_3998,N_4128);
and U5690 (N_5690,N_4974,N_3461);
and U5691 (N_5691,N_2936,N_4795);
xnor U5692 (N_5692,N_4013,N_3325);
nor U5693 (N_5693,N_3554,N_3352);
and U5694 (N_5694,N_3116,N_2657);
nand U5695 (N_5695,N_3734,N_3607);
nand U5696 (N_5696,N_4520,N_4997);
or U5697 (N_5697,N_2697,N_2929);
xnor U5698 (N_5698,N_4185,N_4762);
or U5699 (N_5699,N_3190,N_3329);
or U5700 (N_5700,N_4203,N_4169);
or U5701 (N_5701,N_3744,N_2869);
xnor U5702 (N_5702,N_3261,N_4867);
or U5703 (N_5703,N_4417,N_4727);
xnor U5704 (N_5704,N_4459,N_4443);
nand U5705 (N_5705,N_2820,N_3578);
nand U5706 (N_5706,N_4534,N_4584);
nor U5707 (N_5707,N_4904,N_2709);
xnor U5708 (N_5708,N_2653,N_3163);
and U5709 (N_5709,N_4336,N_4462);
xnor U5710 (N_5710,N_3284,N_2955);
or U5711 (N_5711,N_3751,N_2845);
or U5712 (N_5712,N_2705,N_3041);
nor U5713 (N_5713,N_2506,N_3354);
nor U5714 (N_5714,N_3028,N_3275);
nor U5715 (N_5715,N_3906,N_3732);
nand U5716 (N_5716,N_4556,N_4372);
and U5717 (N_5717,N_3755,N_3969);
xor U5718 (N_5718,N_2515,N_3548);
nor U5719 (N_5719,N_4978,N_2857);
and U5720 (N_5720,N_3307,N_4086);
or U5721 (N_5721,N_4413,N_4845);
nand U5722 (N_5722,N_3470,N_2816);
or U5723 (N_5723,N_4496,N_3296);
or U5724 (N_5724,N_2901,N_4819);
and U5725 (N_5725,N_2731,N_3931);
xnor U5726 (N_5726,N_3251,N_2867);
and U5727 (N_5727,N_2713,N_2904);
nand U5728 (N_5728,N_4408,N_4052);
nor U5729 (N_5729,N_3281,N_3894);
xor U5730 (N_5730,N_2920,N_3076);
and U5731 (N_5731,N_2728,N_3044);
nor U5732 (N_5732,N_3611,N_2773);
and U5733 (N_5733,N_2852,N_3023);
or U5734 (N_5734,N_2647,N_4324);
nand U5735 (N_5735,N_3071,N_2663);
and U5736 (N_5736,N_4394,N_3823);
nand U5737 (N_5737,N_3321,N_2821);
nor U5738 (N_5738,N_3006,N_4479);
and U5739 (N_5739,N_3964,N_3907);
nand U5740 (N_5740,N_4919,N_4283);
nor U5741 (N_5741,N_3892,N_2859);
nor U5742 (N_5742,N_4968,N_3508);
nand U5743 (N_5743,N_3310,N_3862);
nand U5744 (N_5744,N_3132,N_4630);
nor U5745 (N_5745,N_4688,N_3712);
nand U5746 (N_5746,N_3177,N_2770);
and U5747 (N_5747,N_4900,N_3599);
nand U5748 (N_5748,N_4150,N_2563);
nand U5749 (N_5749,N_3341,N_4552);
nor U5750 (N_5750,N_4354,N_3211);
nand U5751 (N_5751,N_3210,N_3788);
xor U5752 (N_5752,N_3854,N_4017);
or U5753 (N_5753,N_4569,N_2893);
or U5754 (N_5754,N_2814,N_3872);
and U5755 (N_5755,N_3279,N_3413);
nor U5756 (N_5756,N_3077,N_4151);
and U5757 (N_5757,N_4679,N_3342);
nand U5758 (N_5758,N_3469,N_3022);
nor U5759 (N_5759,N_3392,N_3241);
and U5760 (N_5760,N_4990,N_4313);
nor U5761 (N_5761,N_3532,N_4163);
or U5762 (N_5762,N_3277,N_3600);
or U5763 (N_5763,N_3361,N_3713);
nor U5764 (N_5764,N_2785,N_4464);
nor U5765 (N_5765,N_4862,N_3204);
nor U5766 (N_5766,N_2981,N_4287);
nand U5767 (N_5767,N_3108,N_3605);
and U5768 (N_5768,N_4964,N_2907);
nor U5769 (N_5769,N_3693,N_2741);
xnor U5770 (N_5770,N_3555,N_2963);
and U5771 (N_5771,N_4907,N_3272);
nor U5772 (N_5772,N_2989,N_2584);
or U5773 (N_5773,N_4915,N_3687);
nor U5774 (N_5774,N_4195,N_4238);
nor U5775 (N_5775,N_3316,N_2533);
and U5776 (N_5776,N_2803,N_3721);
and U5777 (N_5777,N_3378,N_4781);
nor U5778 (N_5778,N_4650,N_4531);
and U5779 (N_5779,N_3098,N_2690);
or U5780 (N_5780,N_2790,N_4760);
nor U5781 (N_5781,N_3288,N_4766);
and U5782 (N_5782,N_4806,N_3664);
nor U5783 (N_5783,N_4858,N_3306);
nor U5784 (N_5784,N_4827,N_3468);
nand U5785 (N_5785,N_3789,N_4297);
xor U5786 (N_5786,N_2753,N_4917);
nor U5787 (N_5787,N_2985,N_2631);
or U5788 (N_5788,N_3235,N_4211);
nor U5789 (N_5789,N_4859,N_3096);
and U5790 (N_5790,N_4539,N_4389);
xor U5791 (N_5791,N_4941,N_4402);
nand U5792 (N_5792,N_3032,N_3518);
nand U5793 (N_5793,N_3553,N_4714);
xor U5794 (N_5794,N_3087,N_3809);
and U5795 (N_5795,N_3450,N_3510);
nand U5796 (N_5796,N_2692,N_2591);
nor U5797 (N_5797,N_2702,N_3727);
or U5798 (N_5798,N_2606,N_2794);
nor U5799 (N_5799,N_4949,N_4554);
or U5800 (N_5800,N_3908,N_3161);
or U5801 (N_5801,N_4444,N_3013);
nor U5802 (N_5802,N_4627,N_2822);
and U5803 (N_5803,N_4261,N_4615);
or U5804 (N_5804,N_4484,N_4373);
and U5805 (N_5805,N_2600,N_3878);
nand U5806 (N_5806,N_2882,N_3897);
nand U5807 (N_5807,N_3322,N_4494);
nor U5808 (N_5808,N_4357,N_2630);
and U5809 (N_5809,N_4268,N_2614);
nand U5810 (N_5810,N_3405,N_4051);
nor U5811 (N_5811,N_4116,N_2782);
and U5812 (N_5812,N_2763,N_4737);
nand U5813 (N_5813,N_3293,N_4659);
nand U5814 (N_5814,N_3062,N_3524);
or U5815 (N_5815,N_4326,N_4138);
nor U5816 (N_5816,N_4685,N_2626);
nand U5817 (N_5817,N_2666,N_4614);
or U5818 (N_5818,N_4826,N_2592);
nor U5819 (N_5819,N_4625,N_2715);
nor U5820 (N_5820,N_4129,N_2990);
nor U5821 (N_5821,N_3726,N_2523);
or U5822 (N_5822,N_2809,N_3435);
nand U5823 (N_5823,N_4438,N_4368);
nand U5824 (N_5824,N_3940,N_3166);
nand U5825 (N_5825,N_2549,N_4418);
and U5826 (N_5826,N_2500,N_4255);
and U5827 (N_5827,N_3250,N_2847);
nand U5828 (N_5828,N_4112,N_3289);
and U5829 (N_5829,N_4682,N_4745);
nand U5830 (N_5830,N_3094,N_4612);
xnor U5831 (N_5831,N_4329,N_4932);
nor U5832 (N_5832,N_3037,N_4019);
or U5833 (N_5833,N_4107,N_2802);
and U5834 (N_5834,N_4160,N_4350);
and U5835 (N_5835,N_4161,N_3381);
nor U5836 (N_5836,N_2732,N_3679);
nor U5837 (N_5837,N_2652,N_4269);
or U5838 (N_5838,N_2688,N_2999);
nor U5839 (N_5839,N_3208,N_3802);
or U5840 (N_5840,N_2776,N_3722);
nand U5841 (N_5841,N_3668,N_3105);
nand U5842 (N_5842,N_4121,N_4084);
nand U5843 (N_5843,N_4649,N_3528);
and U5844 (N_5844,N_4655,N_4722);
nor U5845 (N_5845,N_2609,N_3425);
and U5846 (N_5846,N_3024,N_4456);
or U5847 (N_5847,N_3737,N_4582);
or U5848 (N_5848,N_3626,N_2723);
or U5849 (N_5849,N_2835,N_3916);
and U5850 (N_5850,N_2501,N_4576);
xor U5851 (N_5851,N_4572,N_3885);
and U5852 (N_5852,N_3065,N_4083);
and U5853 (N_5853,N_2733,N_4277);
nor U5854 (N_5854,N_2596,N_3312);
and U5855 (N_5855,N_4229,N_4571);
nor U5856 (N_5856,N_3304,N_3739);
nand U5857 (N_5857,N_4797,N_4392);
or U5858 (N_5858,N_4689,N_2954);
or U5859 (N_5859,N_4477,N_4015);
nor U5860 (N_5860,N_3058,N_4164);
nand U5861 (N_5861,N_3455,N_3114);
nand U5862 (N_5862,N_2661,N_4043);
nor U5863 (N_5863,N_3992,N_2810);
and U5864 (N_5864,N_4276,N_2736);
or U5865 (N_5865,N_3217,N_4725);
nand U5866 (N_5866,N_2995,N_4256);
xnor U5867 (N_5867,N_3618,N_4284);
and U5868 (N_5868,N_2544,N_2916);
xor U5869 (N_5869,N_3183,N_3760);
or U5870 (N_5870,N_4362,N_3127);
and U5871 (N_5871,N_3538,N_3056);
or U5872 (N_5872,N_4807,N_3864);
xnor U5873 (N_5873,N_2786,N_4088);
or U5874 (N_5874,N_2886,N_4472);
and U5875 (N_5875,N_3702,N_4424);
nand U5876 (N_5876,N_3517,N_3027);
or U5877 (N_5877,N_2752,N_3511);
and U5878 (N_5878,N_2593,N_2603);
nand U5879 (N_5879,N_3989,N_2701);
nand U5880 (N_5880,N_4073,N_4592);
or U5881 (N_5881,N_3917,N_4801);
nand U5882 (N_5882,N_3051,N_2676);
and U5883 (N_5883,N_3961,N_3265);
nor U5884 (N_5884,N_4314,N_4719);
nand U5885 (N_5885,N_3268,N_3666);
and U5886 (N_5886,N_3648,N_3589);
xor U5887 (N_5887,N_4838,N_2738);
nor U5888 (N_5888,N_4212,N_2674);
nand U5889 (N_5889,N_3757,N_2527);
and U5890 (N_5890,N_3000,N_3643);
and U5891 (N_5891,N_3483,N_3671);
or U5892 (N_5892,N_4471,N_3781);
or U5893 (N_5893,N_4911,N_3060);
or U5894 (N_5894,N_3215,N_4514);
nand U5895 (N_5895,N_3745,N_2983);
or U5896 (N_5896,N_4001,N_4285);
and U5897 (N_5897,N_3710,N_4667);
or U5898 (N_5898,N_4553,N_3896);
nor U5899 (N_5899,N_2836,N_4746);
or U5900 (N_5900,N_4606,N_3092);
nor U5901 (N_5901,N_4317,N_2918);
nor U5902 (N_5902,N_4698,N_4565);
nand U5903 (N_5903,N_2505,N_4923);
nand U5904 (N_5904,N_4218,N_2887);
or U5905 (N_5905,N_3199,N_3402);
nand U5906 (N_5906,N_3440,N_4741);
nand U5907 (N_5907,N_3999,N_4924);
or U5908 (N_5908,N_3865,N_2594);
nor U5909 (N_5909,N_3834,N_3933);
nand U5910 (N_5910,N_4873,N_4593);
and U5911 (N_5911,N_4267,N_2856);
nand U5912 (N_5912,N_2749,N_3278);
xor U5913 (N_5913,N_3606,N_3280);
or U5914 (N_5914,N_3089,N_2542);
nand U5915 (N_5915,N_2744,N_3097);
or U5916 (N_5916,N_3689,N_4793);
or U5917 (N_5917,N_2975,N_3086);
xnor U5918 (N_5918,N_2858,N_4478);
nand U5919 (N_5919,N_4557,N_4231);
xnor U5920 (N_5920,N_4360,N_4834);
xor U5921 (N_5921,N_3149,N_3610);
nand U5922 (N_5922,N_4253,N_4064);
or U5923 (N_5923,N_2839,N_3613);
nand U5924 (N_5924,N_3057,N_4049);
or U5925 (N_5925,N_3615,N_2760);
xnor U5926 (N_5926,N_3870,N_3848);
or U5927 (N_5927,N_2894,N_4736);
nand U5928 (N_5928,N_2927,N_4482);
nand U5929 (N_5929,N_3503,N_3314);
or U5930 (N_5930,N_4320,N_4040);
and U5931 (N_5931,N_2576,N_3030);
nand U5932 (N_5932,N_2874,N_3266);
or U5933 (N_5933,N_3395,N_4192);
nor U5934 (N_5934,N_3115,N_4982);
and U5935 (N_5935,N_4435,N_2698);
or U5936 (N_5936,N_2868,N_3021);
xnor U5937 (N_5937,N_4648,N_2881);
or U5938 (N_5938,N_2548,N_4522);
nand U5939 (N_5939,N_3959,N_4631);
xor U5940 (N_5940,N_4453,N_3965);
nand U5941 (N_5941,N_4993,N_3393);
xnor U5942 (N_5942,N_2552,N_3914);
nor U5943 (N_5943,N_3978,N_4820);
nand U5944 (N_5944,N_4735,N_3556);
nor U5945 (N_5945,N_3394,N_4681);
nand U5946 (N_5946,N_4216,N_4728);
xor U5947 (N_5947,N_4029,N_3331);
xnor U5948 (N_5948,N_3771,N_4307);
and U5949 (N_5949,N_3641,N_3201);
or U5950 (N_5950,N_3773,N_3839);
nand U5951 (N_5951,N_3536,N_2730);
nand U5952 (N_5952,N_4980,N_3488);
nor U5953 (N_5953,N_2945,N_4935);
or U5954 (N_5954,N_4570,N_2830);
and U5955 (N_5955,N_2854,N_4292);
nor U5956 (N_5956,N_3973,N_4414);
or U5957 (N_5957,N_3603,N_3681);
or U5958 (N_5958,N_4560,N_4751);
or U5959 (N_5959,N_4488,N_2675);
and U5960 (N_5960,N_4693,N_4106);
nand U5961 (N_5961,N_3810,N_4661);
or U5962 (N_5962,N_4260,N_3206);
nand U5963 (N_5963,N_3356,N_2798);
xnor U5964 (N_5964,N_4991,N_2864);
and U5965 (N_5965,N_3111,N_3291);
and U5966 (N_5966,N_3996,N_3446);
and U5967 (N_5967,N_3287,N_2979);
nand U5968 (N_5968,N_2758,N_4855);
nor U5969 (N_5969,N_4731,N_2944);
nand U5970 (N_5970,N_4027,N_3911);
nor U5971 (N_5971,N_4031,N_2656);
xnor U5972 (N_5972,N_4262,N_2792);
xor U5973 (N_5973,N_3162,N_4172);
nor U5974 (N_5974,N_4152,N_3748);
or U5975 (N_5975,N_4122,N_3496);
or U5976 (N_5976,N_3597,N_3824);
or U5977 (N_5977,N_3598,N_4789);
xnor U5978 (N_5978,N_4530,N_2530);
and U5979 (N_5979,N_2976,N_3943);
nand U5980 (N_5980,N_3619,N_3106);
or U5981 (N_5981,N_3343,N_4067);
nor U5982 (N_5982,N_4058,N_4940);
nor U5983 (N_5983,N_2935,N_3572);
or U5984 (N_5984,N_2580,N_3620);
nor U5985 (N_5985,N_3074,N_2900);
or U5986 (N_5986,N_3798,N_3224);
or U5987 (N_5987,N_2827,N_3416);
or U5988 (N_5988,N_3730,N_4173);
and U5989 (N_5989,N_4364,N_3067);
nor U5990 (N_5990,N_3308,N_3633);
and U5991 (N_5991,N_4407,N_2718);
or U5992 (N_5992,N_2574,N_4641);
nor U5993 (N_5993,N_2750,N_2812);
nor U5994 (N_5994,N_4246,N_4739);
or U5995 (N_5995,N_4395,N_3486);
nor U5996 (N_5996,N_2992,N_4487);
or U5997 (N_5997,N_4545,N_4985);
nor U5998 (N_5998,N_3465,N_3061);
xnor U5999 (N_5999,N_4227,N_2903);
or U6000 (N_6000,N_4647,N_4430);
nand U6001 (N_6001,N_3212,N_3198);
xnor U6002 (N_6002,N_2997,N_4004);
xor U6003 (N_6003,N_3282,N_3629);
nor U6004 (N_6004,N_4646,N_2934);
and U6005 (N_6005,N_2969,N_2684);
nor U6006 (N_6006,N_4233,N_3443);
nand U6007 (N_6007,N_4293,N_3451);
and U6008 (N_6008,N_2813,N_2748);
nand U6009 (N_6009,N_3290,N_2984);
or U6010 (N_6010,N_4640,N_4491);
nand U6011 (N_6011,N_2980,N_4672);
nand U6012 (N_6012,N_4281,N_3909);
or U6013 (N_6013,N_3846,N_3652);
nor U6014 (N_6014,N_3617,N_3521);
and U6015 (N_6015,N_3725,N_4518);
or U6016 (N_6016,N_3501,N_4384);
and U6017 (N_6017,N_3678,N_4550);
and U6018 (N_6018,N_3315,N_4817);
nor U6019 (N_6019,N_3923,N_3902);
nand U6020 (N_6020,N_3531,N_3861);
or U6021 (N_6021,N_3145,N_4168);
and U6022 (N_6022,N_4813,N_2876);
and U6023 (N_6023,N_2824,N_3635);
or U6024 (N_6024,N_4809,N_4134);
nand U6025 (N_6025,N_4983,N_3093);
nor U6026 (N_6026,N_3941,N_4179);
xnor U6027 (N_6027,N_3791,N_4942);
and U6028 (N_6028,N_2946,N_4302);
nor U6029 (N_6029,N_4669,N_4752);
nand U6030 (N_6030,N_4030,N_3319);
and U6031 (N_6031,N_4047,N_3504);
nand U6032 (N_6032,N_2844,N_4798);
or U6033 (N_6033,N_4748,N_4505);
nor U6034 (N_6034,N_4222,N_4473);
or U6035 (N_6035,N_2902,N_4124);
xnor U6036 (N_6036,N_4289,N_4442);
or U6037 (N_6037,N_3348,N_4226);
xor U6038 (N_6038,N_4228,N_4600);
nand U6039 (N_6039,N_3012,N_3935);
and U6040 (N_6040,N_4587,N_4331);
nand U6041 (N_6041,N_3125,N_2872);
nor U6042 (N_6042,N_3926,N_2638);
xor U6043 (N_6043,N_2587,N_3297);
nand U6044 (N_6044,N_2745,N_2964);
nor U6045 (N_6045,N_3879,N_2962);
nor U6046 (N_6046,N_3625,N_4597);
nand U6047 (N_6047,N_4951,N_3592);
nand U6048 (N_6048,N_3438,N_4876);
and U6049 (N_6049,N_3368,N_3505);
or U6050 (N_6050,N_3564,N_4117);
nand U6051 (N_6051,N_3968,N_4498);
or U6052 (N_6052,N_3388,N_3654);
or U6053 (N_6053,N_4022,N_4230);
nor U6054 (N_6054,N_3649,N_3387);
and U6055 (N_6055,N_2554,N_4003);
nor U6056 (N_6056,N_3811,N_3245);
nor U6057 (N_6057,N_3832,N_4996);
xnor U6058 (N_6058,N_3838,N_2589);
or U6059 (N_6059,N_4626,N_4379);
and U6060 (N_6060,N_3444,N_2885);
nor U6061 (N_6061,N_4533,N_3231);
or U6062 (N_6062,N_4805,N_4497);
or U6063 (N_6063,N_3741,N_2627);
nor U6064 (N_6064,N_4476,N_3464);
nand U6065 (N_6065,N_4198,N_3175);
nor U6066 (N_6066,N_2756,N_4423);
and U6067 (N_6067,N_3815,N_3645);
nor U6068 (N_6068,N_2629,N_3328);
nand U6069 (N_6069,N_2679,N_2913);
and U6070 (N_6070,N_3696,N_3139);
nand U6071 (N_6071,N_3220,N_4061);
or U6072 (N_6072,N_2922,N_4159);
and U6073 (N_6073,N_4558,N_3703);
xor U6074 (N_6074,N_4141,N_4115);
nor U6075 (N_6075,N_4045,N_4908);
nor U6076 (N_6076,N_4219,N_4718);
nand U6077 (N_6077,N_3269,N_4110);
nand U6078 (N_6078,N_3258,N_3226);
and U6079 (N_6079,N_3055,N_3474);
nand U6080 (N_6080,N_2508,N_4890);
or U6081 (N_6081,N_4274,N_4296);
or U6082 (N_6082,N_3685,N_4401);
and U6083 (N_6083,N_2757,N_3207);
nor U6084 (N_6084,N_2880,N_4769);
nand U6085 (N_6085,N_3292,N_4607);
or U6086 (N_6086,N_3007,N_4638);
and U6087 (N_6087,N_2691,N_3901);
nand U6088 (N_6088,N_2637,N_4675);
xnor U6089 (N_6089,N_2658,N_4355);
and U6090 (N_6090,N_3406,N_4155);
nand U6091 (N_6091,N_2668,N_2644);
nand U6092 (N_6092,N_3214,N_3073);
nor U6093 (N_6093,N_3985,N_4176);
nand U6094 (N_6094,N_3168,N_3384);
nand U6095 (N_6095,N_3350,N_3081);
nor U6096 (N_6096,N_4812,N_3095);
nor U6097 (N_6097,N_2655,N_4037);
or U6098 (N_6098,N_4493,N_3123);
nand U6099 (N_6099,N_3337,N_2862);
nand U6100 (N_6100,N_3857,N_4369);
or U6101 (N_6101,N_2888,N_4068);
xor U6102 (N_6102,N_3359,N_3004);
nor U6103 (N_6103,N_3836,N_3113);
or U6104 (N_6104,N_4060,N_4249);
xor U6105 (N_6105,N_2734,N_4544);
xnor U6106 (N_6106,N_2680,N_3807);
and U6107 (N_6107,N_4897,N_4643);
xnor U6108 (N_6108,N_4101,N_3302);
nand U6109 (N_6109,N_2513,N_3858);
and U6110 (N_6110,N_3429,N_2649);
or U6111 (N_6111,N_4702,N_3701);
xor U6112 (N_6112,N_4757,N_3683);
nand U6113 (N_6113,N_3653,N_4036);
nor U6114 (N_6114,N_3187,N_4738);
and U6115 (N_6115,N_2909,N_2883);
nor U6116 (N_6116,N_4204,N_4852);
or U6117 (N_6117,N_3386,N_3875);
and U6118 (N_6118,N_3684,N_2961);
nor U6119 (N_6119,N_3945,N_4119);
or U6120 (N_6120,N_3601,N_3886);
nand U6121 (N_6121,N_3692,N_3391);
nand U6122 (N_6122,N_3144,N_4461);
or U6123 (N_6123,N_3047,N_2664);
or U6124 (N_6124,N_4555,N_4691);
nand U6125 (N_6125,N_2555,N_3458);
and U6126 (N_6126,N_3847,N_4207);
and U6127 (N_6127,N_3567,N_4726);
xnor U6128 (N_6128,N_3768,N_4242);
or U6129 (N_6129,N_4610,N_3919);
and U6130 (N_6130,N_2573,N_3195);
nor U6131 (N_6131,N_4541,N_3921);
xnor U6132 (N_6132,N_3228,N_3772);
nor U6133 (N_6133,N_4959,N_3010);
xor U6134 (N_6134,N_3344,N_3723);
and U6135 (N_6135,N_4580,N_3533);
nor U6136 (N_6136,N_2762,N_4695);
nor U6137 (N_6137,N_4883,N_4245);
nand U6138 (N_6138,N_2804,N_3476);
or U6139 (N_6139,N_3431,N_4251);
nand U6140 (N_6140,N_4898,N_4632);
or U6141 (N_6141,N_3202,N_3140);
nor U6142 (N_6142,N_4005,N_3283);
or U6143 (N_6143,N_3490,N_3529);
or U6144 (N_6144,N_2788,N_3371);
nand U6145 (N_6145,N_2569,N_2619);
or U6146 (N_6146,N_2586,N_4197);
nor U6147 (N_6147,N_3417,N_3460);
and U6148 (N_6148,N_3866,N_3239);
nor U6149 (N_6149,N_3830,N_4210);
or U6150 (N_6150,N_3427,N_3756);
or U6151 (N_6151,N_3557,N_3675);
xnor U6152 (N_6152,N_4103,N_4250);
nor U6153 (N_6153,N_3856,N_3418);
and U6154 (N_6154,N_4166,N_4465);
nor U6155 (N_6155,N_2641,N_4038);
nor U6156 (N_6156,N_4984,N_3849);
and U6157 (N_6157,N_4927,N_4055);
nor U6158 (N_6158,N_2708,N_4994);
or U6159 (N_6159,N_4921,N_3887);
xnor U6160 (N_6160,N_4755,N_3244);
nand U6161 (N_6161,N_4696,N_3912);
or U6162 (N_6162,N_3243,N_2960);
and U6163 (N_6163,N_3240,N_3758);
or U6164 (N_6164,N_2825,N_3816);
nand U6165 (N_6165,N_2923,N_4446);
nor U6166 (N_6166,N_4301,N_3500);
xnor U6167 (N_6167,N_4761,N_3167);
xor U6168 (N_6168,N_4356,N_3881);
and U6169 (N_6169,N_4208,N_3152);
nand U6170 (N_6170,N_2815,N_3778);
and U6171 (N_6171,N_4502,N_4930);
or U6172 (N_6172,N_4847,N_3063);
and U6173 (N_6173,N_4157,N_2550);
xor U6174 (N_6174,N_4770,N_3481);
or U6175 (N_6175,N_2906,N_2570);
or U6176 (N_6176,N_4709,N_3349);
or U6177 (N_6177,N_4332,N_3409);
and U6178 (N_6178,N_2648,N_4162);
nor U6179 (N_6179,N_3986,N_4821);
nand U6180 (N_6180,N_3420,N_3225);
and U6181 (N_6181,N_4666,N_4609);
and U6182 (N_6182,N_3188,N_2841);
xor U6183 (N_6183,N_2721,N_2539);
nor U6184 (N_6184,N_3627,N_3623);
or U6185 (N_6185,N_3837,N_3561);
nor U6186 (N_6186,N_4139,N_2568);
nand U6187 (N_6187,N_4975,N_4215);
nand U6188 (N_6188,N_3767,N_2808);
and U6189 (N_6189,N_3324,N_4785);
and U6190 (N_6190,N_4224,N_3102);
xor U6191 (N_6191,N_3040,N_3136);
nor U6192 (N_6192,N_3918,N_3949);
nand U6193 (N_6193,N_3053,N_3377);
xnor U6194 (N_6194,N_3735,N_2950);
or U6195 (N_6195,N_3233,N_3670);
nor U6196 (N_6196,N_2848,N_3516);
nor U6197 (N_6197,N_3580,N_3009);
and U6198 (N_6198,N_3129,N_3373);
or U6199 (N_6199,N_3456,N_3036);
nor U6200 (N_6200,N_3953,N_2743);
nor U6201 (N_6201,N_4517,N_4193);
and U6202 (N_6202,N_4054,N_4670);
nand U6203 (N_6203,N_4750,N_4992);
and U6204 (N_6204,N_3937,N_4854);
nand U6205 (N_6205,N_4729,N_4048);
nand U6206 (N_6206,N_4861,N_3285);
nand U6207 (N_6207,N_4403,N_3452);
nor U6208 (N_6208,N_4790,N_3482);
nor U6209 (N_6209,N_3787,N_3473);
xnor U6210 (N_6210,N_4523,N_3783);
or U6211 (N_6211,N_3659,N_4342);
nor U6212 (N_6212,N_3497,N_4833);
or U6213 (N_6213,N_3507,N_4706);
xor U6214 (N_6214,N_3527,N_4636);
xor U6215 (N_6215,N_3558,N_2536);
or U6216 (N_6216,N_3080,N_4574);
nor U6217 (N_6217,N_2994,N_3682);
xor U6218 (N_6218,N_4660,N_2930);
or U6219 (N_6219,N_2943,N_3267);
nand U6220 (N_6220,N_4564,N_4815);
nor U6221 (N_6221,N_4705,N_4404);
or U6222 (N_6222,N_4684,N_4063);
nor U6223 (N_6223,N_4062,N_2671);
or U6224 (N_6224,N_3930,N_3806);
nor U6225 (N_6225,N_3851,N_3523);
and U6226 (N_6226,N_3704,N_4832);
nand U6227 (N_6227,N_4680,N_2551);
and U6228 (N_6228,N_4409,N_3448);
nand U6229 (N_6229,N_3694,N_2831);
nand U6230 (N_6230,N_3868,N_3367);
and U6231 (N_6231,N_4589,N_4315);
nand U6232 (N_6232,N_2898,N_3170);
or U6233 (N_6233,N_3691,N_4272);
nand U6234 (N_6234,N_4035,N_4810);
nand U6235 (N_6235,N_2577,N_4955);
or U6236 (N_6236,N_3904,N_2766);
or U6237 (N_6237,N_3960,N_4220);
or U6238 (N_6238,N_3579,N_3423);
nand U6239 (N_6239,N_2622,N_4492);
nand U6240 (N_6240,N_4816,N_4848);
nor U6241 (N_6241,N_4076,N_4697);
or U6242 (N_6242,N_3674,N_4513);
or U6243 (N_6243,N_2780,N_2604);
nand U6244 (N_6244,N_2931,N_3566);
nor U6245 (N_6245,N_3103,N_3656);
and U6246 (N_6246,N_3153,N_4551);
xnor U6247 (N_6247,N_2667,N_4440);
nor U6248 (N_6248,N_4343,N_4568);
and U6249 (N_6249,N_4271,N_4396);
or U6250 (N_6250,N_4356,N_4781);
or U6251 (N_6251,N_3960,N_4342);
nand U6252 (N_6252,N_4333,N_3826);
xnor U6253 (N_6253,N_4797,N_4640);
or U6254 (N_6254,N_3541,N_4317);
or U6255 (N_6255,N_4219,N_3070);
or U6256 (N_6256,N_4349,N_3593);
and U6257 (N_6257,N_3539,N_4458);
nand U6258 (N_6258,N_2768,N_2547);
xnor U6259 (N_6259,N_2657,N_2511);
nor U6260 (N_6260,N_4569,N_2569);
nand U6261 (N_6261,N_3487,N_4591);
nand U6262 (N_6262,N_3055,N_2669);
nor U6263 (N_6263,N_3762,N_3980);
xnor U6264 (N_6264,N_3889,N_3053);
nor U6265 (N_6265,N_3679,N_4280);
and U6266 (N_6266,N_3529,N_3128);
and U6267 (N_6267,N_2543,N_4977);
and U6268 (N_6268,N_3044,N_4275);
or U6269 (N_6269,N_4650,N_2683);
nor U6270 (N_6270,N_3453,N_4688);
nor U6271 (N_6271,N_4852,N_4009);
nor U6272 (N_6272,N_2670,N_2958);
and U6273 (N_6273,N_4227,N_2900);
nor U6274 (N_6274,N_4521,N_3476);
nand U6275 (N_6275,N_3937,N_3909);
or U6276 (N_6276,N_3470,N_2601);
or U6277 (N_6277,N_3319,N_3893);
and U6278 (N_6278,N_2725,N_2539);
nor U6279 (N_6279,N_4996,N_4605);
and U6280 (N_6280,N_4404,N_4333);
nand U6281 (N_6281,N_4227,N_4472);
nor U6282 (N_6282,N_2549,N_4158);
or U6283 (N_6283,N_3235,N_3193);
and U6284 (N_6284,N_3848,N_3224);
or U6285 (N_6285,N_3347,N_2833);
or U6286 (N_6286,N_4494,N_4490);
nand U6287 (N_6287,N_2676,N_2964);
or U6288 (N_6288,N_4505,N_4629);
or U6289 (N_6289,N_4574,N_3339);
nand U6290 (N_6290,N_3996,N_2796);
or U6291 (N_6291,N_3307,N_3806);
nor U6292 (N_6292,N_2915,N_4892);
xor U6293 (N_6293,N_4739,N_2665);
or U6294 (N_6294,N_4180,N_3689);
nor U6295 (N_6295,N_3602,N_3540);
or U6296 (N_6296,N_3618,N_4179);
nand U6297 (N_6297,N_3449,N_3101);
nor U6298 (N_6298,N_2586,N_4099);
xnor U6299 (N_6299,N_2927,N_4529);
and U6300 (N_6300,N_4695,N_2822);
and U6301 (N_6301,N_3257,N_2955);
and U6302 (N_6302,N_4149,N_4025);
or U6303 (N_6303,N_4355,N_4366);
xor U6304 (N_6304,N_4552,N_4565);
or U6305 (N_6305,N_3584,N_3056);
or U6306 (N_6306,N_3615,N_4133);
or U6307 (N_6307,N_4695,N_2833);
nand U6308 (N_6308,N_4342,N_4398);
or U6309 (N_6309,N_2547,N_3525);
or U6310 (N_6310,N_3319,N_4983);
xnor U6311 (N_6311,N_4281,N_3705);
nor U6312 (N_6312,N_4129,N_2767);
and U6313 (N_6313,N_4295,N_4494);
nor U6314 (N_6314,N_3788,N_4836);
nor U6315 (N_6315,N_3892,N_3194);
or U6316 (N_6316,N_2796,N_4191);
nand U6317 (N_6317,N_4661,N_4869);
nand U6318 (N_6318,N_4095,N_4767);
nand U6319 (N_6319,N_2516,N_3583);
or U6320 (N_6320,N_2945,N_2500);
and U6321 (N_6321,N_3550,N_4587);
and U6322 (N_6322,N_3910,N_4726);
and U6323 (N_6323,N_2535,N_3785);
nor U6324 (N_6324,N_3090,N_4598);
and U6325 (N_6325,N_4102,N_3998);
or U6326 (N_6326,N_4860,N_2515);
or U6327 (N_6327,N_2690,N_4750);
and U6328 (N_6328,N_4057,N_2881);
and U6329 (N_6329,N_4973,N_3217);
and U6330 (N_6330,N_3982,N_4531);
or U6331 (N_6331,N_4457,N_3065);
nor U6332 (N_6332,N_2855,N_4569);
nand U6333 (N_6333,N_3438,N_4631);
or U6334 (N_6334,N_3607,N_4574);
or U6335 (N_6335,N_3544,N_2570);
and U6336 (N_6336,N_3120,N_4211);
or U6337 (N_6337,N_4309,N_4183);
xnor U6338 (N_6338,N_4850,N_3155);
nor U6339 (N_6339,N_4468,N_3785);
nor U6340 (N_6340,N_4117,N_3217);
nor U6341 (N_6341,N_3084,N_4011);
and U6342 (N_6342,N_3626,N_4902);
nor U6343 (N_6343,N_3996,N_3763);
nor U6344 (N_6344,N_4116,N_3266);
or U6345 (N_6345,N_4633,N_3883);
nand U6346 (N_6346,N_3485,N_3886);
or U6347 (N_6347,N_2656,N_4995);
and U6348 (N_6348,N_3084,N_4630);
nor U6349 (N_6349,N_4276,N_4407);
or U6350 (N_6350,N_4546,N_3200);
nor U6351 (N_6351,N_3598,N_3245);
and U6352 (N_6352,N_4477,N_2548);
and U6353 (N_6353,N_3942,N_4890);
and U6354 (N_6354,N_3159,N_3324);
nand U6355 (N_6355,N_3439,N_3919);
or U6356 (N_6356,N_3834,N_4935);
xnor U6357 (N_6357,N_4650,N_2893);
nand U6358 (N_6358,N_3195,N_4086);
xor U6359 (N_6359,N_2705,N_3441);
or U6360 (N_6360,N_2999,N_2532);
and U6361 (N_6361,N_2560,N_4619);
and U6362 (N_6362,N_2908,N_4900);
or U6363 (N_6363,N_4377,N_4701);
and U6364 (N_6364,N_3140,N_4132);
nand U6365 (N_6365,N_4793,N_2742);
nor U6366 (N_6366,N_4012,N_4218);
or U6367 (N_6367,N_4280,N_4362);
or U6368 (N_6368,N_3713,N_3240);
nor U6369 (N_6369,N_2814,N_3864);
nor U6370 (N_6370,N_2611,N_2860);
nor U6371 (N_6371,N_3380,N_3081);
and U6372 (N_6372,N_2646,N_3351);
xnor U6373 (N_6373,N_2726,N_3230);
nor U6374 (N_6374,N_2795,N_4087);
or U6375 (N_6375,N_3686,N_2803);
and U6376 (N_6376,N_4432,N_3861);
or U6377 (N_6377,N_4106,N_2822);
or U6378 (N_6378,N_3096,N_3869);
or U6379 (N_6379,N_4828,N_3347);
or U6380 (N_6380,N_2639,N_4683);
nand U6381 (N_6381,N_3125,N_4383);
nor U6382 (N_6382,N_3339,N_2965);
nand U6383 (N_6383,N_2816,N_4082);
and U6384 (N_6384,N_2672,N_3557);
and U6385 (N_6385,N_2556,N_2972);
and U6386 (N_6386,N_3455,N_2734);
nor U6387 (N_6387,N_2778,N_3266);
or U6388 (N_6388,N_4189,N_4383);
and U6389 (N_6389,N_2828,N_3346);
nor U6390 (N_6390,N_3919,N_4300);
and U6391 (N_6391,N_3505,N_3891);
nor U6392 (N_6392,N_3789,N_4591);
or U6393 (N_6393,N_4927,N_3265);
or U6394 (N_6394,N_3372,N_3052);
nand U6395 (N_6395,N_3756,N_4567);
xnor U6396 (N_6396,N_3688,N_4657);
nand U6397 (N_6397,N_4454,N_3913);
or U6398 (N_6398,N_3887,N_4828);
nand U6399 (N_6399,N_2620,N_4035);
and U6400 (N_6400,N_3363,N_4295);
xor U6401 (N_6401,N_4508,N_3978);
and U6402 (N_6402,N_3351,N_2895);
and U6403 (N_6403,N_4409,N_3595);
nor U6404 (N_6404,N_3024,N_4228);
nand U6405 (N_6405,N_3354,N_4635);
or U6406 (N_6406,N_3669,N_3412);
nor U6407 (N_6407,N_4315,N_2790);
nand U6408 (N_6408,N_3322,N_4961);
and U6409 (N_6409,N_2596,N_4036);
nor U6410 (N_6410,N_4618,N_3180);
nand U6411 (N_6411,N_4941,N_2509);
or U6412 (N_6412,N_4785,N_4697);
and U6413 (N_6413,N_4842,N_3524);
nand U6414 (N_6414,N_3959,N_3341);
or U6415 (N_6415,N_3166,N_3311);
xor U6416 (N_6416,N_4001,N_4573);
and U6417 (N_6417,N_4482,N_4329);
and U6418 (N_6418,N_4676,N_3493);
nor U6419 (N_6419,N_4630,N_3523);
nand U6420 (N_6420,N_3712,N_2850);
nand U6421 (N_6421,N_3181,N_4532);
and U6422 (N_6422,N_4224,N_4322);
xor U6423 (N_6423,N_3760,N_3747);
nor U6424 (N_6424,N_3594,N_3596);
nor U6425 (N_6425,N_4819,N_2846);
or U6426 (N_6426,N_3493,N_2531);
nand U6427 (N_6427,N_4838,N_4286);
or U6428 (N_6428,N_2871,N_4489);
nand U6429 (N_6429,N_4359,N_4770);
xnor U6430 (N_6430,N_3150,N_4301);
nand U6431 (N_6431,N_4021,N_3428);
and U6432 (N_6432,N_3529,N_2643);
or U6433 (N_6433,N_4643,N_3443);
nor U6434 (N_6434,N_4214,N_3439);
nand U6435 (N_6435,N_3964,N_2767);
xor U6436 (N_6436,N_2895,N_3459);
nand U6437 (N_6437,N_3093,N_3994);
or U6438 (N_6438,N_4148,N_3269);
nor U6439 (N_6439,N_2832,N_4168);
nor U6440 (N_6440,N_4458,N_3820);
and U6441 (N_6441,N_4753,N_3845);
nor U6442 (N_6442,N_4386,N_4204);
nor U6443 (N_6443,N_3371,N_4689);
nor U6444 (N_6444,N_3571,N_4240);
and U6445 (N_6445,N_4173,N_3590);
and U6446 (N_6446,N_4325,N_2537);
nor U6447 (N_6447,N_4233,N_4417);
and U6448 (N_6448,N_3823,N_4288);
nor U6449 (N_6449,N_4713,N_4457);
or U6450 (N_6450,N_2937,N_3775);
and U6451 (N_6451,N_3937,N_4544);
or U6452 (N_6452,N_4206,N_4948);
nor U6453 (N_6453,N_2994,N_3331);
nor U6454 (N_6454,N_3069,N_4770);
nand U6455 (N_6455,N_2506,N_4293);
nand U6456 (N_6456,N_4901,N_2784);
nand U6457 (N_6457,N_3295,N_4509);
xnor U6458 (N_6458,N_3776,N_4838);
nor U6459 (N_6459,N_3369,N_3281);
and U6460 (N_6460,N_2801,N_3532);
or U6461 (N_6461,N_3192,N_4061);
or U6462 (N_6462,N_3745,N_3928);
xor U6463 (N_6463,N_3495,N_4059);
nand U6464 (N_6464,N_4062,N_3516);
and U6465 (N_6465,N_4369,N_3038);
xnor U6466 (N_6466,N_2531,N_3824);
and U6467 (N_6467,N_3647,N_3447);
and U6468 (N_6468,N_4104,N_3560);
and U6469 (N_6469,N_4452,N_2859);
xnor U6470 (N_6470,N_4641,N_4035);
nand U6471 (N_6471,N_4962,N_2973);
nor U6472 (N_6472,N_2735,N_3496);
xor U6473 (N_6473,N_2886,N_2716);
nor U6474 (N_6474,N_3521,N_3104);
nand U6475 (N_6475,N_3563,N_3366);
nand U6476 (N_6476,N_2899,N_2905);
nand U6477 (N_6477,N_4645,N_3365);
nand U6478 (N_6478,N_2994,N_4174);
or U6479 (N_6479,N_4153,N_3209);
or U6480 (N_6480,N_4957,N_3222);
nand U6481 (N_6481,N_3316,N_3096);
nand U6482 (N_6482,N_3188,N_4934);
nand U6483 (N_6483,N_4367,N_4229);
or U6484 (N_6484,N_2618,N_2854);
or U6485 (N_6485,N_4856,N_4308);
nor U6486 (N_6486,N_4856,N_2683);
or U6487 (N_6487,N_4297,N_4434);
or U6488 (N_6488,N_4210,N_3450);
nor U6489 (N_6489,N_2840,N_3968);
nor U6490 (N_6490,N_2611,N_3175);
or U6491 (N_6491,N_3660,N_4536);
nand U6492 (N_6492,N_4657,N_4241);
and U6493 (N_6493,N_3088,N_4972);
or U6494 (N_6494,N_3698,N_4870);
nand U6495 (N_6495,N_4043,N_2575);
nand U6496 (N_6496,N_3747,N_4464);
and U6497 (N_6497,N_4325,N_4960);
and U6498 (N_6498,N_4570,N_3411);
or U6499 (N_6499,N_3531,N_4654);
nand U6500 (N_6500,N_3373,N_3757);
nor U6501 (N_6501,N_3179,N_3296);
or U6502 (N_6502,N_3669,N_4684);
nor U6503 (N_6503,N_4718,N_3246);
or U6504 (N_6504,N_4038,N_3099);
nor U6505 (N_6505,N_4461,N_3718);
or U6506 (N_6506,N_3948,N_4230);
and U6507 (N_6507,N_3953,N_3534);
or U6508 (N_6508,N_4095,N_4286);
or U6509 (N_6509,N_4847,N_3804);
nand U6510 (N_6510,N_3268,N_3025);
nand U6511 (N_6511,N_3119,N_4434);
or U6512 (N_6512,N_4693,N_3957);
and U6513 (N_6513,N_4989,N_2779);
or U6514 (N_6514,N_2911,N_2586);
or U6515 (N_6515,N_3639,N_3113);
nand U6516 (N_6516,N_4268,N_3185);
and U6517 (N_6517,N_3033,N_4908);
nor U6518 (N_6518,N_4832,N_4224);
or U6519 (N_6519,N_4122,N_4886);
and U6520 (N_6520,N_3712,N_2996);
nand U6521 (N_6521,N_4728,N_4711);
or U6522 (N_6522,N_3149,N_3569);
and U6523 (N_6523,N_4444,N_3085);
and U6524 (N_6524,N_3899,N_4401);
nor U6525 (N_6525,N_3126,N_2973);
nand U6526 (N_6526,N_2908,N_2539);
nor U6527 (N_6527,N_4426,N_4525);
nor U6528 (N_6528,N_3400,N_4779);
nor U6529 (N_6529,N_4913,N_4058);
nand U6530 (N_6530,N_4841,N_4570);
nor U6531 (N_6531,N_4894,N_4461);
nor U6532 (N_6532,N_4358,N_2742);
nand U6533 (N_6533,N_3900,N_3014);
and U6534 (N_6534,N_3395,N_4514);
nand U6535 (N_6535,N_4932,N_4685);
nand U6536 (N_6536,N_4399,N_4028);
nor U6537 (N_6537,N_4893,N_4197);
or U6538 (N_6538,N_3696,N_4796);
and U6539 (N_6539,N_3774,N_4540);
nor U6540 (N_6540,N_4510,N_4876);
and U6541 (N_6541,N_4508,N_4237);
nor U6542 (N_6542,N_3438,N_2757);
or U6543 (N_6543,N_3808,N_3443);
and U6544 (N_6544,N_3976,N_4830);
nand U6545 (N_6545,N_3591,N_4493);
and U6546 (N_6546,N_3404,N_2663);
and U6547 (N_6547,N_4580,N_3340);
or U6548 (N_6548,N_2819,N_3819);
nor U6549 (N_6549,N_4000,N_4701);
xor U6550 (N_6550,N_2957,N_3261);
nand U6551 (N_6551,N_2774,N_4695);
nor U6552 (N_6552,N_4720,N_4140);
nor U6553 (N_6553,N_4486,N_2750);
and U6554 (N_6554,N_3929,N_2691);
nand U6555 (N_6555,N_4233,N_3251);
and U6556 (N_6556,N_4854,N_3867);
nand U6557 (N_6557,N_4069,N_4635);
and U6558 (N_6558,N_4791,N_2654);
nand U6559 (N_6559,N_2969,N_3544);
and U6560 (N_6560,N_2840,N_4724);
nand U6561 (N_6561,N_3927,N_3603);
xnor U6562 (N_6562,N_4518,N_3147);
and U6563 (N_6563,N_4936,N_3728);
or U6564 (N_6564,N_4637,N_4501);
or U6565 (N_6565,N_2959,N_4254);
or U6566 (N_6566,N_4174,N_4560);
and U6567 (N_6567,N_4580,N_3534);
nand U6568 (N_6568,N_4623,N_2887);
and U6569 (N_6569,N_2788,N_4161);
nor U6570 (N_6570,N_4662,N_4671);
nor U6571 (N_6571,N_3928,N_4398);
nand U6572 (N_6572,N_3627,N_4527);
nor U6573 (N_6573,N_3881,N_3541);
xnor U6574 (N_6574,N_4910,N_3957);
nand U6575 (N_6575,N_3780,N_4155);
xor U6576 (N_6576,N_2798,N_3263);
nand U6577 (N_6577,N_3005,N_3524);
nor U6578 (N_6578,N_4685,N_4260);
and U6579 (N_6579,N_3199,N_4947);
or U6580 (N_6580,N_4618,N_4010);
and U6581 (N_6581,N_3381,N_4950);
nor U6582 (N_6582,N_3963,N_4731);
nor U6583 (N_6583,N_2561,N_4116);
nand U6584 (N_6584,N_4762,N_2567);
nand U6585 (N_6585,N_3478,N_3465);
or U6586 (N_6586,N_3472,N_4011);
nor U6587 (N_6587,N_2955,N_4184);
nand U6588 (N_6588,N_3481,N_4453);
nor U6589 (N_6589,N_3995,N_4950);
or U6590 (N_6590,N_4035,N_3239);
and U6591 (N_6591,N_3601,N_2864);
xnor U6592 (N_6592,N_3025,N_3564);
or U6593 (N_6593,N_3362,N_4020);
nand U6594 (N_6594,N_4802,N_4441);
and U6595 (N_6595,N_3151,N_4237);
or U6596 (N_6596,N_4289,N_4714);
nor U6597 (N_6597,N_4779,N_4185);
and U6598 (N_6598,N_3926,N_3782);
or U6599 (N_6599,N_2925,N_4898);
nor U6600 (N_6600,N_2969,N_4741);
or U6601 (N_6601,N_4902,N_4893);
nor U6602 (N_6602,N_2690,N_2900);
and U6603 (N_6603,N_2902,N_4363);
or U6604 (N_6604,N_2688,N_4777);
xnor U6605 (N_6605,N_3270,N_3712);
nor U6606 (N_6606,N_3581,N_4796);
and U6607 (N_6607,N_3503,N_3427);
or U6608 (N_6608,N_3051,N_4549);
nand U6609 (N_6609,N_3943,N_4258);
or U6610 (N_6610,N_4042,N_4959);
nor U6611 (N_6611,N_3769,N_3705);
and U6612 (N_6612,N_4979,N_4707);
nand U6613 (N_6613,N_2893,N_3719);
nand U6614 (N_6614,N_3035,N_2753);
nand U6615 (N_6615,N_3276,N_3406);
or U6616 (N_6616,N_4674,N_2835);
nor U6617 (N_6617,N_2627,N_4919);
nand U6618 (N_6618,N_3142,N_3192);
nor U6619 (N_6619,N_2715,N_2644);
or U6620 (N_6620,N_3835,N_4228);
nand U6621 (N_6621,N_4207,N_4372);
and U6622 (N_6622,N_4195,N_3728);
or U6623 (N_6623,N_4585,N_4908);
xor U6624 (N_6624,N_2527,N_4565);
nor U6625 (N_6625,N_4091,N_3812);
nor U6626 (N_6626,N_4904,N_4623);
nand U6627 (N_6627,N_3352,N_3817);
and U6628 (N_6628,N_4034,N_3191);
or U6629 (N_6629,N_2638,N_3347);
xor U6630 (N_6630,N_3966,N_3909);
nor U6631 (N_6631,N_4717,N_3611);
nand U6632 (N_6632,N_3352,N_3697);
nand U6633 (N_6633,N_2621,N_4260);
xor U6634 (N_6634,N_3413,N_3159);
nand U6635 (N_6635,N_2500,N_2824);
or U6636 (N_6636,N_3193,N_3794);
or U6637 (N_6637,N_3971,N_4627);
or U6638 (N_6638,N_3096,N_4174);
or U6639 (N_6639,N_2985,N_4159);
nand U6640 (N_6640,N_4897,N_3524);
xor U6641 (N_6641,N_3141,N_2811);
nor U6642 (N_6642,N_3456,N_4908);
nor U6643 (N_6643,N_4702,N_4013);
nor U6644 (N_6644,N_2720,N_4758);
nand U6645 (N_6645,N_3653,N_4143);
and U6646 (N_6646,N_3588,N_3561);
nand U6647 (N_6647,N_4670,N_2627);
nand U6648 (N_6648,N_4892,N_4581);
nor U6649 (N_6649,N_4200,N_2703);
nor U6650 (N_6650,N_4957,N_4139);
nand U6651 (N_6651,N_3272,N_3584);
nor U6652 (N_6652,N_3995,N_3127);
nand U6653 (N_6653,N_3256,N_2582);
and U6654 (N_6654,N_4671,N_3764);
or U6655 (N_6655,N_3114,N_2947);
or U6656 (N_6656,N_4094,N_3985);
and U6657 (N_6657,N_2869,N_3747);
or U6658 (N_6658,N_4522,N_4233);
and U6659 (N_6659,N_4031,N_3156);
nand U6660 (N_6660,N_4512,N_3694);
and U6661 (N_6661,N_3440,N_3331);
or U6662 (N_6662,N_3054,N_2992);
or U6663 (N_6663,N_3725,N_2527);
or U6664 (N_6664,N_2736,N_4425);
and U6665 (N_6665,N_4528,N_2779);
and U6666 (N_6666,N_4006,N_3529);
or U6667 (N_6667,N_4175,N_4825);
xnor U6668 (N_6668,N_3505,N_3688);
and U6669 (N_6669,N_4853,N_4143);
or U6670 (N_6670,N_2512,N_4266);
nor U6671 (N_6671,N_4305,N_2597);
nand U6672 (N_6672,N_4677,N_3282);
nor U6673 (N_6673,N_3501,N_2523);
nand U6674 (N_6674,N_4171,N_3290);
and U6675 (N_6675,N_4396,N_3786);
and U6676 (N_6676,N_4339,N_2967);
and U6677 (N_6677,N_3398,N_2860);
or U6678 (N_6678,N_3764,N_4480);
and U6679 (N_6679,N_2676,N_2911);
nand U6680 (N_6680,N_2852,N_2699);
nand U6681 (N_6681,N_2800,N_4855);
nand U6682 (N_6682,N_3034,N_2842);
or U6683 (N_6683,N_4887,N_3447);
nor U6684 (N_6684,N_3604,N_4904);
xor U6685 (N_6685,N_3682,N_3809);
nand U6686 (N_6686,N_3144,N_3955);
nor U6687 (N_6687,N_4131,N_4202);
nand U6688 (N_6688,N_2954,N_3027);
nor U6689 (N_6689,N_2924,N_4557);
or U6690 (N_6690,N_4323,N_4961);
or U6691 (N_6691,N_4754,N_4794);
and U6692 (N_6692,N_2689,N_4340);
nand U6693 (N_6693,N_4318,N_3025);
and U6694 (N_6694,N_2604,N_2503);
nor U6695 (N_6695,N_3528,N_3227);
nor U6696 (N_6696,N_2843,N_2821);
xor U6697 (N_6697,N_4538,N_3198);
or U6698 (N_6698,N_3978,N_4496);
and U6699 (N_6699,N_2501,N_3610);
xnor U6700 (N_6700,N_3537,N_3382);
and U6701 (N_6701,N_3737,N_4761);
nand U6702 (N_6702,N_2589,N_4328);
nor U6703 (N_6703,N_2827,N_2851);
xnor U6704 (N_6704,N_3354,N_3514);
or U6705 (N_6705,N_2719,N_4135);
xnor U6706 (N_6706,N_3546,N_3670);
nand U6707 (N_6707,N_2810,N_3904);
and U6708 (N_6708,N_3513,N_2834);
xor U6709 (N_6709,N_3505,N_2692);
and U6710 (N_6710,N_2582,N_4687);
nor U6711 (N_6711,N_3480,N_2971);
and U6712 (N_6712,N_4103,N_2544);
nand U6713 (N_6713,N_3578,N_4914);
nor U6714 (N_6714,N_2776,N_3032);
or U6715 (N_6715,N_4584,N_3286);
nand U6716 (N_6716,N_4365,N_4626);
and U6717 (N_6717,N_4627,N_2626);
nor U6718 (N_6718,N_3279,N_4837);
nand U6719 (N_6719,N_4202,N_3810);
nand U6720 (N_6720,N_4925,N_4250);
nand U6721 (N_6721,N_2795,N_4641);
nor U6722 (N_6722,N_3513,N_4748);
nand U6723 (N_6723,N_4651,N_4262);
nand U6724 (N_6724,N_2590,N_3071);
nor U6725 (N_6725,N_3425,N_3056);
nor U6726 (N_6726,N_2909,N_4540);
and U6727 (N_6727,N_3880,N_3809);
nand U6728 (N_6728,N_3329,N_2583);
or U6729 (N_6729,N_4678,N_3300);
and U6730 (N_6730,N_4778,N_2749);
nand U6731 (N_6731,N_2887,N_3636);
nor U6732 (N_6732,N_4899,N_3836);
or U6733 (N_6733,N_4831,N_3549);
nor U6734 (N_6734,N_4956,N_2620);
xnor U6735 (N_6735,N_4533,N_3759);
or U6736 (N_6736,N_3321,N_4043);
nor U6737 (N_6737,N_3090,N_4097);
and U6738 (N_6738,N_3683,N_2586);
or U6739 (N_6739,N_3706,N_4667);
and U6740 (N_6740,N_3356,N_3027);
nand U6741 (N_6741,N_3715,N_3964);
and U6742 (N_6742,N_2520,N_4636);
and U6743 (N_6743,N_4912,N_4471);
nand U6744 (N_6744,N_3479,N_4567);
and U6745 (N_6745,N_4863,N_4405);
nand U6746 (N_6746,N_4959,N_2809);
and U6747 (N_6747,N_2716,N_3940);
nor U6748 (N_6748,N_3801,N_3828);
and U6749 (N_6749,N_4373,N_2697);
nand U6750 (N_6750,N_4657,N_4170);
and U6751 (N_6751,N_3530,N_3133);
nor U6752 (N_6752,N_2798,N_2511);
and U6753 (N_6753,N_4692,N_4158);
or U6754 (N_6754,N_3397,N_4850);
nor U6755 (N_6755,N_3038,N_3846);
nand U6756 (N_6756,N_2908,N_4939);
or U6757 (N_6757,N_4564,N_2742);
xnor U6758 (N_6758,N_4761,N_3892);
and U6759 (N_6759,N_4333,N_4914);
nand U6760 (N_6760,N_4136,N_2680);
nor U6761 (N_6761,N_4688,N_4710);
nor U6762 (N_6762,N_4786,N_4725);
nand U6763 (N_6763,N_3758,N_3479);
and U6764 (N_6764,N_4283,N_2579);
nand U6765 (N_6765,N_3769,N_3633);
xor U6766 (N_6766,N_3473,N_3642);
and U6767 (N_6767,N_4273,N_2925);
and U6768 (N_6768,N_4824,N_3144);
nand U6769 (N_6769,N_2615,N_3485);
and U6770 (N_6770,N_2910,N_2666);
nor U6771 (N_6771,N_4513,N_4179);
nand U6772 (N_6772,N_3544,N_4009);
or U6773 (N_6773,N_4977,N_4666);
xnor U6774 (N_6774,N_4432,N_3938);
or U6775 (N_6775,N_4982,N_3317);
or U6776 (N_6776,N_3134,N_2777);
or U6777 (N_6777,N_4953,N_4911);
xor U6778 (N_6778,N_4753,N_3417);
nand U6779 (N_6779,N_4552,N_4387);
nor U6780 (N_6780,N_3337,N_3399);
and U6781 (N_6781,N_3667,N_4093);
nand U6782 (N_6782,N_3289,N_4955);
or U6783 (N_6783,N_4602,N_4834);
nand U6784 (N_6784,N_4931,N_3296);
nand U6785 (N_6785,N_3625,N_2641);
or U6786 (N_6786,N_2529,N_4244);
nand U6787 (N_6787,N_3201,N_4176);
or U6788 (N_6788,N_3533,N_3661);
nor U6789 (N_6789,N_3189,N_4478);
nand U6790 (N_6790,N_4925,N_4655);
nand U6791 (N_6791,N_3308,N_3588);
or U6792 (N_6792,N_3236,N_4351);
or U6793 (N_6793,N_3802,N_3819);
xor U6794 (N_6794,N_4061,N_3568);
or U6795 (N_6795,N_3142,N_4098);
nand U6796 (N_6796,N_3272,N_4881);
nand U6797 (N_6797,N_3566,N_3764);
nand U6798 (N_6798,N_3459,N_4576);
nor U6799 (N_6799,N_3207,N_4580);
and U6800 (N_6800,N_4232,N_3816);
or U6801 (N_6801,N_4133,N_3230);
nand U6802 (N_6802,N_2719,N_3155);
nor U6803 (N_6803,N_3812,N_4130);
or U6804 (N_6804,N_3377,N_4929);
or U6805 (N_6805,N_3292,N_2542);
nand U6806 (N_6806,N_4529,N_4110);
xor U6807 (N_6807,N_3391,N_3629);
xor U6808 (N_6808,N_3122,N_4976);
and U6809 (N_6809,N_4093,N_3586);
nor U6810 (N_6810,N_2599,N_4301);
nand U6811 (N_6811,N_4768,N_3134);
nor U6812 (N_6812,N_4145,N_3233);
and U6813 (N_6813,N_4959,N_4880);
nand U6814 (N_6814,N_3818,N_3741);
nand U6815 (N_6815,N_3528,N_3856);
or U6816 (N_6816,N_4291,N_3360);
nor U6817 (N_6817,N_2916,N_2630);
xor U6818 (N_6818,N_4537,N_4111);
or U6819 (N_6819,N_4997,N_3863);
and U6820 (N_6820,N_3597,N_2956);
nor U6821 (N_6821,N_3319,N_4796);
nand U6822 (N_6822,N_3811,N_3826);
xnor U6823 (N_6823,N_3904,N_2658);
nor U6824 (N_6824,N_2728,N_4942);
nand U6825 (N_6825,N_3308,N_3647);
nor U6826 (N_6826,N_4726,N_3323);
and U6827 (N_6827,N_2777,N_4858);
or U6828 (N_6828,N_3851,N_4394);
or U6829 (N_6829,N_3598,N_4791);
nand U6830 (N_6830,N_4462,N_3681);
nand U6831 (N_6831,N_3525,N_4696);
xnor U6832 (N_6832,N_4582,N_4002);
nand U6833 (N_6833,N_2614,N_4015);
nor U6834 (N_6834,N_4202,N_4649);
or U6835 (N_6835,N_3977,N_3701);
nand U6836 (N_6836,N_4827,N_3653);
nor U6837 (N_6837,N_2686,N_2645);
xor U6838 (N_6838,N_4726,N_4708);
nand U6839 (N_6839,N_3419,N_3247);
nand U6840 (N_6840,N_4711,N_4056);
nand U6841 (N_6841,N_4480,N_4171);
and U6842 (N_6842,N_4581,N_3825);
or U6843 (N_6843,N_2877,N_4007);
nand U6844 (N_6844,N_4896,N_2946);
and U6845 (N_6845,N_3712,N_4824);
nand U6846 (N_6846,N_2522,N_3859);
nand U6847 (N_6847,N_4466,N_4246);
xor U6848 (N_6848,N_3920,N_3955);
and U6849 (N_6849,N_3455,N_4971);
nand U6850 (N_6850,N_4103,N_2951);
or U6851 (N_6851,N_2829,N_4529);
or U6852 (N_6852,N_3622,N_4640);
nor U6853 (N_6853,N_4893,N_3988);
and U6854 (N_6854,N_4395,N_3562);
and U6855 (N_6855,N_4703,N_3198);
nand U6856 (N_6856,N_4449,N_2975);
and U6857 (N_6857,N_4015,N_4451);
xnor U6858 (N_6858,N_3223,N_3359);
nor U6859 (N_6859,N_3374,N_2557);
or U6860 (N_6860,N_3443,N_3260);
and U6861 (N_6861,N_3078,N_3397);
nand U6862 (N_6862,N_4246,N_3214);
nand U6863 (N_6863,N_2567,N_2870);
or U6864 (N_6864,N_4929,N_3757);
or U6865 (N_6865,N_4315,N_4740);
nor U6866 (N_6866,N_2526,N_4648);
or U6867 (N_6867,N_3364,N_2809);
nand U6868 (N_6868,N_3235,N_3874);
or U6869 (N_6869,N_3578,N_3376);
nand U6870 (N_6870,N_4023,N_3746);
and U6871 (N_6871,N_4566,N_4889);
nor U6872 (N_6872,N_3716,N_3087);
nor U6873 (N_6873,N_4263,N_4307);
and U6874 (N_6874,N_3836,N_4433);
or U6875 (N_6875,N_3308,N_3316);
nand U6876 (N_6876,N_2904,N_4925);
nand U6877 (N_6877,N_4274,N_4876);
nor U6878 (N_6878,N_3437,N_3899);
and U6879 (N_6879,N_4760,N_4836);
and U6880 (N_6880,N_4109,N_4574);
and U6881 (N_6881,N_4278,N_4363);
and U6882 (N_6882,N_3948,N_4099);
nor U6883 (N_6883,N_3061,N_3728);
or U6884 (N_6884,N_4420,N_3225);
nor U6885 (N_6885,N_4436,N_3588);
nand U6886 (N_6886,N_4450,N_2709);
nand U6887 (N_6887,N_4034,N_3916);
xnor U6888 (N_6888,N_4302,N_4836);
nand U6889 (N_6889,N_4509,N_3512);
nand U6890 (N_6890,N_4667,N_3561);
and U6891 (N_6891,N_4972,N_3248);
nand U6892 (N_6892,N_4524,N_4904);
or U6893 (N_6893,N_2675,N_2801);
nand U6894 (N_6894,N_4738,N_4918);
nand U6895 (N_6895,N_4134,N_4210);
xor U6896 (N_6896,N_3219,N_3210);
xnor U6897 (N_6897,N_3954,N_3125);
xor U6898 (N_6898,N_3608,N_3796);
and U6899 (N_6899,N_4443,N_3202);
and U6900 (N_6900,N_4922,N_4692);
nor U6901 (N_6901,N_4173,N_2794);
or U6902 (N_6902,N_2990,N_4965);
or U6903 (N_6903,N_4086,N_2620);
nand U6904 (N_6904,N_4587,N_4413);
and U6905 (N_6905,N_3852,N_3354);
or U6906 (N_6906,N_4424,N_4457);
or U6907 (N_6907,N_3437,N_4559);
and U6908 (N_6908,N_4049,N_3106);
xor U6909 (N_6909,N_3752,N_3922);
or U6910 (N_6910,N_4802,N_3267);
and U6911 (N_6911,N_2952,N_3438);
or U6912 (N_6912,N_4082,N_3337);
nor U6913 (N_6913,N_3409,N_3117);
nor U6914 (N_6914,N_4948,N_2775);
or U6915 (N_6915,N_4081,N_2810);
and U6916 (N_6916,N_2954,N_4743);
or U6917 (N_6917,N_4070,N_2657);
xnor U6918 (N_6918,N_4078,N_3720);
nand U6919 (N_6919,N_4466,N_3935);
nor U6920 (N_6920,N_4260,N_2673);
or U6921 (N_6921,N_2665,N_3515);
or U6922 (N_6922,N_4779,N_4372);
and U6923 (N_6923,N_2788,N_4587);
nand U6924 (N_6924,N_4367,N_4158);
nand U6925 (N_6925,N_4878,N_4739);
xor U6926 (N_6926,N_3562,N_4094);
and U6927 (N_6927,N_3454,N_4891);
and U6928 (N_6928,N_2823,N_4570);
nand U6929 (N_6929,N_3144,N_3082);
or U6930 (N_6930,N_3682,N_3606);
nand U6931 (N_6931,N_2724,N_4865);
or U6932 (N_6932,N_3846,N_4861);
or U6933 (N_6933,N_4577,N_2867);
or U6934 (N_6934,N_4992,N_4176);
nand U6935 (N_6935,N_3648,N_4667);
or U6936 (N_6936,N_3869,N_4898);
xor U6937 (N_6937,N_3908,N_4030);
nand U6938 (N_6938,N_4711,N_4404);
nor U6939 (N_6939,N_2876,N_4793);
and U6940 (N_6940,N_3233,N_4713);
xnor U6941 (N_6941,N_4153,N_3065);
nor U6942 (N_6942,N_3623,N_2782);
and U6943 (N_6943,N_4187,N_3662);
and U6944 (N_6944,N_2906,N_4084);
and U6945 (N_6945,N_4145,N_3040);
and U6946 (N_6946,N_2611,N_3908);
nand U6947 (N_6947,N_3690,N_4581);
nor U6948 (N_6948,N_2804,N_3866);
and U6949 (N_6949,N_3927,N_4498);
nor U6950 (N_6950,N_4918,N_2821);
xnor U6951 (N_6951,N_3192,N_4826);
nor U6952 (N_6952,N_4489,N_3571);
or U6953 (N_6953,N_2666,N_4526);
nand U6954 (N_6954,N_4524,N_2559);
nand U6955 (N_6955,N_2874,N_3273);
nand U6956 (N_6956,N_2908,N_4814);
xor U6957 (N_6957,N_4518,N_4154);
or U6958 (N_6958,N_3774,N_3632);
or U6959 (N_6959,N_3404,N_2781);
nor U6960 (N_6960,N_3991,N_3786);
nand U6961 (N_6961,N_4513,N_3402);
xnor U6962 (N_6962,N_3917,N_4804);
and U6963 (N_6963,N_3051,N_2726);
nor U6964 (N_6964,N_4763,N_3194);
and U6965 (N_6965,N_3300,N_2992);
nand U6966 (N_6966,N_3457,N_3235);
or U6967 (N_6967,N_2694,N_3592);
nor U6968 (N_6968,N_3760,N_2968);
nand U6969 (N_6969,N_3839,N_4405);
xnor U6970 (N_6970,N_3453,N_4052);
nand U6971 (N_6971,N_2796,N_4777);
and U6972 (N_6972,N_2864,N_4907);
xnor U6973 (N_6973,N_4554,N_4352);
and U6974 (N_6974,N_4384,N_4283);
nor U6975 (N_6975,N_4225,N_4655);
nor U6976 (N_6976,N_2886,N_3817);
or U6977 (N_6977,N_3910,N_4713);
xor U6978 (N_6978,N_3342,N_3448);
nor U6979 (N_6979,N_3765,N_2552);
or U6980 (N_6980,N_2789,N_4173);
xnor U6981 (N_6981,N_4218,N_2968);
nor U6982 (N_6982,N_3791,N_2512);
and U6983 (N_6983,N_4619,N_3700);
and U6984 (N_6984,N_4288,N_4550);
and U6985 (N_6985,N_2882,N_3978);
and U6986 (N_6986,N_3543,N_3867);
or U6987 (N_6987,N_4699,N_3847);
nand U6988 (N_6988,N_2533,N_3096);
nand U6989 (N_6989,N_4270,N_3520);
and U6990 (N_6990,N_3263,N_4990);
or U6991 (N_6991,N_4291,N_4614);
nand U6992 (N_6992,N_4043,N_4570);
and U6993 (N_6993,N_2839,N_4812);
and U6994 (N_6994,N_3197,N_4521);
and U6995 (N_6995,N_3901,N_3246);
nor U6996 (N_6996,N_4163,N_2980);
nand U6997 (N_6997,N_4018,N_4938);
xor U6998 (N_6998,N_4308,N_3829);
nor U6999 (N_6999,N_2828,N_4945);
and U7000 (N_7000,N_4874,N_2795);
or U7001 (N_7001,N_3533,N_2912);
and U7002 (N_7002,N_3068,N_2530);
nor U7003 (N_7003,N_4653,N_4422);
or U7004 (N_7004,N_3748,N_4041);
nand U7005 (N_7005,N_2659,N_4383);
and U7006 (N_7006,N_4807,N_4313);
nor U7007 (N_7007,N_3435,N_2842);
nand U7008 (N_7008,N_4432,N_3644);
and U7009 (N_7009,N_3631,N_2528);
and U7010 (N_7010,N_4237,N_3954);
or U7011 (N_7011,N_4231,N_2934);
and U7012 (N_7012,N_2900,N_3992);
nor U7013 (N_7013,N_2603,N_2948);
nor U7014 (N_7014,N_3908,N_3936);
and U7015 (N_7015,N_3487,N_3872);
and U7016 (N_7016,N_4226,N_3314);
nor U7017 (N_7017,N_4035,N_4435);
and U7018 (N_7018,N_3261,N_3007);
xnor U7019 (N_7019,N_3718,N_4997);
nor U7020 (N_7020,N_4135,N_4516);
or U7021 (N_7021,N_3774,N_3867);
xor U7022 (N_7022,N_2962,N_4535);
or U7023 (N_7023,N_4038,N_4418);
and U7024 (N_7024,N_2689,N_4685);
or U7025 (N_7025,N_3848,N_2784);
nand U7026 (N_7026,N_2638,N_3715);
or U7027 (N_7027,N_4309,N_4457);
nor U7028 (N_7028,N_3256,N_4021);
or U7029 (N_7029,N_4808,N_2550);
and U7030 (N_7030,N_2796,N_3804);
and U7031 (N_7031,N_3608,N_2970);
nor U7032 (N_7032,N_2935,N_4164);
nand U7033 (N_7033,N_3641,N_3675);
nand U7034 (N_7034,N_3896,N_3161);
nand U7035 (N_7035,N_2861,N_4259);
nor U7036 (N_7036,N_3558,N_3129);
or U7037 (N_7037,N_4991,N_2534);
or U7038 (N_7038,N_2859,N_3528);
xor U7039 (N_7039,N_4778,N_4358);
nor U7040 (N_7040,N_4131,N_4024);
or U7041 (N_7041,N_4977,N_2858);
nor U7042 (N_7042,N_4016,N_3347);
or U7043 (N_7043,N_4276,N_3712);
nand U7044 (N_7044,N_4860,N_4434);
or U7045 (N_7045,N_4505,N_4901);
nand U7046 (N_7046,N_3183,N_4489);
nand U7047 (N_7047,N_4975,N_4123);
or U7048 (N_7048,N_4817,N_2876);
nand U7049 (N_7049,N_3677,N_2995);
or U7050 (N_7050,N_2799,N_4341);
nor U7051 (N_7051,N_3700,N_3719);
and U7052 (N_7052,N_4062,N_3271);
or U7053 (N_7053,N_2704,N_4051);
and U7054 (N_7054,N_3751,N_3323);
or U7055 (N_7055,N_2865,N_3114);
nor U7056 (N_7056,N_3426,N_3036);
and U7057 (N_7057,N_4975,N_3866);
and U7058 (N_7058,N_4587,N_3777);
or U7059 (N_7059,N_3569,N_4498);
or U7060 (N_7060,N_3864,N_3175);
or U7061 (N_7061,N_4098,N_3107);
or U7062 (N_7062,N_2563,N_4396);
nor U7063 (N_7063,N_4230,N_3605);
nor U7064 (N_7064,N_4308,N_4513);
and U7065 (N_7065,N_2553,N_2617);
or U7066 (N_7066,N_2565,N_2796);
or U7067 (N_7067,N_4546,N_3328);
or U7068 (N_7068,N_4296,N_3238);
or U7069 (N_7069,N_3621,N_3478);
nor U7070 (N_7070,N_4935,N_4047);
or U7071 (N_7071,N_3353,N_4184);
nor U7072 (N_7072,N_4966,N_3974);
nor U7073 (N_7073,N_3389,N_3518);
nand U7074 (N_7074,N_3708,N_3334);
nand U7075 (N_7075,N_2948,N_2722);
nand U7076 (N_7076,N_2753,N_2848);
or U7077 (N_7077,N_3116,N_4168);
nor U7078 (N_7078,N_3401,N_4152);
or U7079 (N_7079,N_2718,N_3484);
and U7080 (N_7080,N_2541,N_3492);
or U7081 (N_7081,N_3065,N_4826);
or U7082 (N_7082,N_4161,N_4981);
xor U7083 (N_7083,N_2598,N_3875);
nor U7084 (N_7084,N_2644,N_4923);
xor U7085 (N_7085,N_2903,N_2629);
nor U7086 (N_7086,N_4034,N_4764);
nor U7087 (N_7087,N_4249,N_3334);
or U7088 (N_7088,N_4863,N_2891);
and U7089 (N_7089,N_4754,N_4774);
nand U7090 (N_7090,N_4889,N_4082);
nand U7091 (N_7091,N_3682,N_2961);
nand U7092 (N_7092,N_2642,N_3826);
and U7093 (N_7093,N_3111,N_4084);
nor U7094 (N_7094,N_2533,N_3716);
and U7095 (N_7095,N_4839,N_3951);
nand U7096 (N_7096,N_3916,N_4881);
nor U7097 (N_7097,N_4836,N_4021);
nor U7098 (N_7098,N_4405,N_2886);
xnor U7099 (N_7099,N_2688,N_3261);
nor U7100 (N_7100,N_3904,N_4218);
and U7101 (N_7101,N_4277,N_4663);
or U7102 (N_7102,N_3060,N_3497);
or U7103 (N_7103,N_3788,N_3068);
nor U7104 (N_7104,N_3568,N_3351);
nor U7105 (N_7105,N_3936,N_4977);
nor U7106 (N_7106,N_4006,N_4414);
or U7107 (N_7107,N_4116,N_4552);
nand U7108 (N_7108,N_3941,N_3887);
and U7109 (N_7109,N_3327,N_2686);
nor U7110 (N_7110,N_3024,N_4734);
or U7111 (N_7111,N_2993,N_3959);
and U7112 (N_7112,N_4673,N_4160);
nand U7113 (N_7113,N_3408,N_3572);
nand U7114 (N_7114,N_4284,N_4561);
and U7115 (N_7115,N_2916,N_4397);
nor U7116 (N_7116,N_2825,N_4901);
nand U7117 (N_7117,N_3669,N_2839);
or U7118 (N_7118,N_3012,N_4791);
nand U7119 (N_7119,N_3571,N_4886);
nor U7120 (N_7120,N_3484,N_2770);
nand U7121 (N_7121,N_2736,N_2743);
xnor U7122 (N_7122,N_2735,N_3626);
or U7123 (N_7123,N_4980,N_4692);
nor U7124 (N_7124,N_3218,N_3277);
nor U7125 (N_7125,N_3181,N_3384);
nand U7126 (N_7126,N_4260,N_3435);
xnor U7127 (N_7127,N_3577,N_4214);
nand U7128 (N_7128,N_4589,N_4603);
xor U7129 (N_7129,N_2791,N_3582);
nor U7130 (N_7130,N_4579,N_3568);
nor U7131 (N_7131,N_4265,N_4731);
or U7132 (N_7132,N_3787,N_4459);
nand U7133 (N_7133,N_2890,N_3044);
and U7134 (N_7134,N_4148,N_3125);
and U7135 (N_7135,N_2651,N_3162);
xor U7136 (N_7136,N_2699,N_4915);
xnor U7137 (N_7137,N_4927,N_4818);
or U7138 (N_7138,N_4226,N_2933);
and U7139 (N_7139,N_2553,N_3645);
or U7140 (N_7140,N_2534,N_2869);
or U7141 (N_7141,N_4114,N_3038);
xor U7142 (N_7142,N_3756,N_2655);
and U7143 (N_7143,N_2605,N_4573);
nand U7144 (N_7144,N_2946,N_4347);
nor U7145 (N_7145,N_3298,N_3729);
nand U7146 (N_7146,N_2681,N_2660);
and U7147 (N_7147,N_4079,N_4033);
or U7148 (N_7148,N_3300,N_3762);
or U7149 (N_7149,N_4159,N_2629);
xnor U7150 (N_7150,N_2679,N_3660);
nor U7151 (N_7151,N_4177,N_4966);
nor U7152 (N_7152,N_3816,N_3106);
xnor U7153 (N_7153,N_4940,N_4873);
nand U7154 (N_7154,N_4025,N_4553);
nand U7155 (N_7155,N_4146,N_3182);
nand U7156 (N_7156,N_3413,N_4627);
or U7157 (N_7157,N_4533,N_4637);
or U7158 (N_7158,N_3121,N_3665);
or U7159 (N_7159,N_4842,N_4065);
nor U7160 (N_7160,N_3043,N_4798);
nand U7161 (N_7161,N_3471,N_4403);
xnor U7162 (N_7162,N_3447,N_3802);
xor U7163 (N_7163,N_3782,N_2512);
nand U7164 (N_7164,N_4404,N_4066);
xor U7165 (N_7165,N_3309,N_2624);
or U7166 (N_7166,N_4243,N_2814);
nor U7167 (N_7167,N_3840,N_3197);
or U7168 (N_7168,N_2673,N_3696);
nand U7169 (N_7169,N_4802,N_2689);
xnor U7170 (N_7170,N_2698,N_4959);
nor U7171 (N_7171,N_2741,N_3783);
nor U7172 (N_7172,N_3756,N_4852);
nand U7173 (N_7173,N_4522,N_2527);
nand U7174 (N_7174,N_3140,N_4536);
nor U7175 (N_7175,N_4969,N_3766);
and U7176 (N_7176,N_3066,N_3535);
xor U7177 (N_7177,N_2749,N_4764);
nand U7178 (N_7178,N_3844,N_2845);
or U7179 (N_7179,N_2645,N_4219);
and U7180 (N_7180,N_4243,N_4120);
nand U7181 (N_7181,N_4702,N_2641);
nand U7182 (N_7182,N_2558,N_4164);
or U7183 (N_7183,N_2617,N_4662);
or U7184 (N_7184,N_2526,N_3446);
nand U7185 (N_7185,N_2992,N_4370);
and U7186 (N_7186,N_2578,N_3757);
nor U7187 (N_7187,N_4780,N_4964);
and U7188 (N_7188,N_2647,N_4650);
or U7189 (N_7189,N_3637,N_3544);
and U7190 (N_7190,N_3943,N_2546);
and U7191 (N_7191,N_3205,N_2769);
nand U7192 (N_7192,N_4602,N_2808);
nand U7193 (N_7193,N_4489,N_3562);
nand U7194 (N_7194,N_4119,N_4147);
and U7195 (N_7195,N_3932,N_2566);
or U7196 (N_7196,N_2531,N_3197);
nand U7197 (N_7197,N_4306,N_3631);
and U7198 (N_7198,N_4352,N_4933);
or U7199 (N_7199,N_2693,N_3994);
nand U7200 (N_7200,N_3915,N_2624);
and U7201 (N_7201,N_2973,N_2781);
nor U7202 (N_7202,N_4497,N_3512);
or U7203 (N_7203,N_2592,N_3837);
nand U7204 (N_7204,N_3989,N_3312);
nand U7205 (N_7205,N_2958,N_3495);
or U7206 (N_7206,N_3080,N_4387);
nor U7207 (N_7207,N_4478,N_2615);
nand U7208 (N_7208,N_2884,N_2850);
and U7209 (N_7209,N_4372,N_4413);
nand U7210 (N_7210,N_2638,N_2902);
nand U7211 (N_7211,N_3582,N_2832);
nand U7212 (N_7212,N_3909,N_3307);
nand U7213 (N_7213,N_4585,N_2901);
or U7214 (N_7214,N_4642,N_4028);
and U7215 (N_7215,N_3314,N_4923);
and U7216 (N_7216,N_4480,N_2803);
nor U7217 (N_7217,N_3588,N_2564);
and U7218 (N_7218,N_3535,N_2763);
or U7219 (N_7219,N_4776,N_4721);
or U7220 (N_7220,N_4177,N_2540);
nor U7221 (N_7221,N_4112,N_4130);
or U7222 (N_7222,N_3390,N_3781);
nand U7223 (N_7223,N_4817,N_3908);
or U7224 (N_7224,N_4791,N_3101);
and U7225 (N_7225,N_4185,N_4791);
or U7226 (N_7226,N_4954,N_4656);
or U7227 (N_7227,N_2958,N_2989);
nor U7228 (N_7228,N_4662,N_3868);
and U7229 (N_7229,N_3767,N_2987);
or U7230 (N_7230,N_3684,N_4391);
and U7231 (N_7231,N_4989,N_4787);
and U7232 (N_7232,N_4476,N_4217);
nor U7233 (N_7233,N_4416,N_4445);
xor U7234 (N_7234,N_4423,N_2790);
and U7235 (N_7235,N_2726,N_4830);
or U7236 (N_7236,N_3059,N_3113);
or U7237 (N_7237,N_3007,N_2625);
nand U7238 (N_7238,N_4113,N_2577);
or U7239 (N_7239,N_3368,N_4428);
xor U7240 (N_7240,N_3312,N_3355);
and U7241 (N_7241,N_3490,N_3791);
or U7242 (N_7242,N_4026,N_4913);
xnor U7243 (N_7243,N_3622,N_4291);
nor U7244 (N_7244,N_2843,N_2922);
nor U7245 (N_7245,N_4309,N_3823);
nand U7246 (N_7246,N_4336,N_4185);
nand U7247 (N_7247,N_4044,N_4329);
and U7248 (N_7248,N_4282,N_3480);
nor U7249 (N_7249,N_3582,N_2872);
and U7250 (N_7250,N_2702,N_4838);
nand U7251 (N_7251,N_2669,N_4145);
nand U7252 (N_7252,N_3075,N_2614);
nand U7253 (N_7253,N_4838,N_4568);
or U7254 (N_7254,N_2784,N_2962);
or U7255 (N_7255,N_2596,N_3682);
nand U7256 (N_7256,N_2749,N_4271);
xnor U7257 (N_7257,N_3782,N_3461);
nor U7258 (N_7258,N_3945,N_3278);
and U7259 (N_7259,N_2659,N_2648);
or U7260 (N_7260,N_4629,N_3802);
xnor U7261 (N_7261,N_2848,N_3223);
and U7262 (N_7262,N_4254,N_3490);
and U7263 (N_7263,N_3857,N_3439);
and U7264 (N_7264,N_4921,N_2855);
and U7265 (N_7265,N_2754,N_4708);
nor U7266 (N_7266,N_4776,N_3140);
nor U7267 (N_7267,N_4239,N_4688);
or U7268 (N_7268,N_2923,N_3200);
and U7269 (N_7269,N_4694,N_3775);
nand U7270 (N_7270,N_3286,N_4666);
or U7271 (N_7271,N_4996,N_4482);
nor U7272 (N_7272,N_4895,N_4045);
and U7273 (N_7273,N_3834,N_3352);
or U7274 (N_7274,N_4235,N_4434);
or U7275 (N_7275,N_3856,N_4424);
nor U7276 (N_7276,N_4862,N_3845);
or U7277 (N_7277,N_4101,N_2973);
or U7278 (N_7278,N_2572,N_2670);
or U7279 (N_7279,N_4871,N_4155);
nor U7280 (N_7280,N_4776,N_3671);
and U7281 (N_7281,N_2853,N_4568);
or U7282 (N_7282,N_4663,N_3956);
nand U7283 (N_7283,N_4231,N_3062);
nor U7284 (N_7284,N_3759,N_2857);
nand U7285 (N_7285,N_3878,N_3927);
and U7286 (N_7286,N_2957,N_3113);
and U7287 (N_7287,N_3992,N_3297);
nor U7288 (N_7288,N_3718,N_4961);
nand U7289 (N_7289,N_4593,N_4054);
xor U7290 (N_7290,N_4470,N_4052);
or U7291 (N_7291,N_2977,N_3590);
and U7292 (N_7292,N_3718,N_3325);
nand U7293 (N_7293,N_4948,N_3845);
or U7294 (N_7294,N_3596,N_3497);
nor U7295 (N_7295,N_3619,N_3696);
or U7296 (N_7296,N_3014,N_3584);
and U7297 (N_7297,N_2583,N_2585);
and U7298 (N_7298,N_3674,N_4239);
nor U7299 (N_7299,N_3821,N_2779);
nand U7300 (N_7300,N_3620,N_4267);
nor U7301 (N_7301,N_2648,N_3639);
and U7302 (N_7302,N_3969,N_4629);
xor U7303 (N_7303,N_3851,N_4207);
and U7304 (N_7304,N_3620,N_2524);
nor U7305 (N_7305,N_4645,N_2592);
nor U7306 (N_7306,N_4075,N_3848);
nor U7307 (N_7307,N_3411,N_3739);
nor U7308 (N_7308,N_2923,N_3212);
nor U7309 (N_7309,N_3145,N_4209);
nand U7310 (N_7310,N_4254,N_4497);
xnor U7311 (N_7311,N_3768,N_3042);
nand U7312 (N_7312,N_4503,N_2715);
or U7313 (N_7313,N_3789,N_4220);
and U7314 (N_7314,N_4259,N_4623);
xor U7315 (N_7315,N_4530,N_4389);
nor U7316 (N_7316,N_3675,N_4712);
nand U7317 (N_7317,N_4211,N_3425);
xnor U7318 (N_7318,N_3111,N_3220);
or U7319 (N_7319,N_3333,N_3377);
nand U7320 (N_7320,N_2973,N_2761);
xor U7321 (N_7321,N_3449,N_4965);
nand U7322 (N_7322,N_4091,N_2631);
nor U7323 (N_7323,N_4312,N_2909);
or U7324 (N_7324,N_4579,N_3561);
nand U7325 (N_7325,N_4818,N_4174);
and U7326 (N_7326,N_4123,N_3486);
and U7327 (N_7327,N_3983,N_2892);
nand U7328 (N_7328,N_4011,N_3952);
xor U7329 (N_7329,N_4265,N_3504);
nor U7330 (N_7330,N_4640,N_2886);
nor U7331 (N_7331,N_4299,N_4085);
xor U7332 (N_7332,N_2603,N_3893);
nand U7333 (N_7333,N_4851,N_3818);
or U7334 (N_7334,N_2546,N_4963);
nor U7335 (N_7335,N_3550,N_4204);
or U7336 (N_7336,N_4276,N_2728);
and U7337 (N_7337,N_3498,N_4343);
and U7338 (N_7338,N_3284,N_2936);
nand U7339 (N_7339,N_3105,N_4466);
nand U7340 (N_7340,N_3314,N_4030);
and U7341 (N_7341,N_4096,N_4305);
nand U7342 (N_7342,N_3790,N_4192);
nand U7343 (N_7343,N_4737,N_3354);
xor U7344 (N_7344,N_4067,N_4611);
or U7345 (N_7345,N_3321,N_3029);
or U7346 (N_7346,N_3725,N_3541);
nand U7347 (N_7347,N_3415,N_4059);
nor U7348 (N_7348,N_4911,N_3133);
nor U7349 (N_7349,N_3863,N_4795);
nand U7350 (N_7350,N_3822,N_3381);
or U7351 (N_7351,N_2740,N_4522);
and U7352 (N_7352,N_2928,N_4912);
or U7353 (N_7353,N_3129,N_4285);
and U7354 (N_7354,N_2839,N_3079);
nor U7355 (N_7355,N_4363,N_4079);
nor U7356 (N_7356,N_4441,N_3884);
and U7357 (N_7357,N_3018,N_2794);
xnor U7358 (N_7358,N_3756,N_4783);
nor U7359 (N_7359,N_2821,N_4284);
or U7360 (N_7360,N_4933,N_3545);
and U7361 (N_7361,N_4573,N_3214);
and U7362 (N_7362,N_2530,N_3458);
or U7363 (N_7363,N_3088,N_4420);
and U7364 (N_7364,N_2968,N_3697);
xnor U7365 (N_7365,N_4486,N_2702);
and U7366 (N_7366,N_3234,N_2941);
and U7367 (N_7367,N_4382,N_3532);
nand U7368 (N_7368,N_3340,N_3144);
and U7369 (N_7369,N_4915,N_3876);
and U7370 (N_7370,N_4017,N_2756);
nand U7371 (N_7371,N_4949,N_3002);
nor U7372 (N_7372,N_4960,N_4970);
nor U7373 (N_7373,N_2889,N_4122);
or U7374 (N_7374,N_3588,N_2936);
xor U7375 (N_7375,N_3857,N_4741);
and U7376 (N_7376,N_2890,N_2716);
nand U7377 (N_7377,N_3557,N_4445);
or U7378 (N_7378,N_3945,N_4973);
xnor U7379 (N_7379,N_3713,N_3867);
and U7380 (N_7380,N_3500,N_4796);
nand U7381 (N_7381,N_3321,N_4018);
or U7382 (N_7382,N_2593,N_2550);
nand U7383 (N_7383,N_4067,N_4474);
nand U7384 (N_7384,N_4906,N_4457);
nand U7385 (N_7385,N_4315,N_3641);
nor U7386 (N_7386,N_3110,N_2593);
and U7387 (N_7387,N_4104,N_2815);
xnor U7388 (N_7388,N_2626,N_3832);
and U7389 (N_7389,N_4620,N_3894);
or U7390 (N_7390,N_4967,N_2563);
and U7391 (N_7391,N_4475,N_3823);
nand U7392 (N_7392,N_3628,N_4960);
nor U7393 (N_7393,N_2666,N_2547);
and U7394 (N_7394,N_4053,N_4729);
xnor U7395 (N_7395,N_4390,N_3772);
or U7396 (N_7396,N_3881,N_3492);
nor U7397 (N_7397,N_3528,N_2922);
or U7398 (N_7398,N_4972,N_2683);
nand U7399 (N_7399,N_4190,N_3922);
xnor U7400 (N_7400,N_4816,N_3251);
nand U7401 (N_7401,N_3733,N_4975);
nand U7402 (N_7402,N_3390,N_2776);
or U7403 (N_7403,N_4509,N_2956);
or U7404 (N_7404,N_3003,N_4856);
xor U7405 (N_7405,N_4117,N_3206);
or U7406 (N_7406,N_3027,N_4068);
xnor U7407 (N_7407,N_2578,N_3047);
nor U7408 (N_7408,N_3573,N_3380);
or U7409 (N_7409,N_4061,N_3599);
or U7410 (N_7410,N_4782,N_3984);
nor U7411 (N_7411,N_4518,N_4366);
and U7412 (N_7412,N_4756,N_3811);
xor U7413 (N_7413,N_4603,N_4415);
or U7414 (N_7414,N_2975,N_4367);
nor U7415 (N_7415,N_3005,N_3893);
nand U7416 (N_7416,N_3888,N_2694);
and U7417 (N_7417,N_4279,N_3632);
or U7418 (N_7418,N_4543,N_3484);
or U7419 (N_7419,N_3985,N_2610);
nor U7420 (N_7420,N_3693,N_4063);
xnor U7421 (N_7421,N_2950,N_2806);
nand U7422 (N_7422,N_4203,N_3607);
xor U7423 (N_7423,N_4750,N_3605);
nand U7424 (N_7424,N_4524,N_4119);
and U7425 (N_7425,N_3127,N_4234);
and U7426 (N_7426,N_2708,N_3140);
nor U7427 (N_7427,N_4461,N_2547);
nor U7428 (N_7428,N_3631,N_4318);
or U7429 (N_7429,N_4732,N_4912);
nand U7430 (N_7430,N_3500,N_3516);
or U7431 (N_7431,N_4212,N_4223);
nand U7432 (N_7432,N_4368,N_3217);
and U7433 (N_7433,N_2654,N_3529);
xnor U7434 (N_7434,N_3162,N_4252);
nand U7435 (N_7435,N_4021,N_4986);
or U7436 (N_7436,N_2662,N_4710);
or U7437 (N_7437,N_4184,N_3351);
nor U7438 (N_7438,N_3469,N_4031);
nand U7439 (N_7439,N_4969,N_4930);
or U7440 (N_7440,N_4326,N_4116);
and U7441 (N_7441,N_4452,N_3916);
and U7442 (N_7442,N_2882,N_2682);
xnor U7443 (N_7443,N_4012,N_2835);
and U7444 (N_7444,N_3042,N_4829);
nor U7445 (N_7445,N_4792,N_4820);
nor U7446 (N_7446,N_2915,N_3034);
and U7447 (N_7447,N_4039,N_3907);
or U7448 (N_7448,N_4292,N_2858);
nor U7449 (N_7449,N_3323,N_3296);
nor U7450 (N_7450,N_3575,N_4593);
nor U7451 (N_7451,N_2597,N_3453);
nand U7452 (N_7452,N_2556,N_3637);
or U7453 (N_7453,N_3346,N_2587);
nor U7454 (N_7454,N_3709,N_2884);
xnor U7455 (N_7455,N_3602,N_3732);
and U7456 (N_7456,N_4121,N_4038);
and U7457 (N_7457,N_3907,N_3701);
nand U7458 (N_7458,N_2589,N_4846);
xor U7459 (N_7459,N_3694,N_3820);
nand U7460 (N_7460,N_3381,N_3698);
nand U7461 (N_7461,N_3475,N_3448);
nor U7462 (N_7462,N_2766,N_4296);
nor U7463 (N_7463,N_4055,N_3000);
and U7464 (N_7464,N_3654,N_3709);
nand U7465 (N_7465,N_3908,N_3300);
nand U7466 (N_7466,N_4409,N_2948);
or U7467 (N_7467,N_2579,N_4273);
or U7468 (N_7468,N_2847,N_4017);
nor U7469 (N_7469,N_3740,N_4153);
nand U7470 (N_7470,N_4653,N_3634);
and U7471 (N_7471,N_2910,N_4887);
and U7472 (N_7472,N_4578,N_2724);
nand U7473 (N_7473,N_2876,N_2872);
and U7474 (N_7474,N_4531,N_4443);
nor U7475 (N_7475,N_3272,N_2622);
nand U7476 (N_7476,N_2649,N_4917);
nand U7477 (N_7477,N_4864,N_3046);
nand U7478 (N_7478,N_4429,N_4546);
nand U7479 (N_7479,N_4451,N_3559);
nor U7480 (N_7480,N_3981,N_3311);
nor U7481 (N_7481,N_4637,N_4470);
or U7482 (N_7482,N_3601,N_3788);
or U7483 (N_7483,N_4478,N_3135);
nor U7484 (N_7484,N_3327,N_4852);
and U7485 (N_7485,N_2859,N_2863);
or U7486 (N_7486,N_4611,N_3966);
or U7487 (N_7487,N_4968,N_3438);
xor U7488 (N_7488,N_4480,N_3550);
and U7489 (N_7489,N_3203,N_3244);
nand U7490 (N_7490,N_4195,N_3419);
nor U7491 (N_7491,N_3021,N_3902);
or U7492 (N_7492,N_4547,N_3890);
nand U7493 (N_7493,N_4659,N_3822);
nand U7494 (N_7494,N_4586,N_3812);
nand U7495 (N_7495,N_3511,N_3100);
and U7496 (N_7496,N_3026,N_3523);
nor U7497 (N_7497,N_4240,N_3194);
or U7498 (N_7498,N_4178,N_2542);
or U7499 (N_7499,N_3429,N_4888);
and U7500 (N_7500,N_7477,N_5971);
or U7501 (N_7501,N_5183,N_5484);
or U7502 (N_7502,N_6218,N_6639);
nor U7503 (N_7503,N_7263,N_5406);
nor U7504 (N_7504,N_7415,N_7434);
nor U7505 (N_7505,N_5405,N_5871);
nor U7506 (N_7506,N_5788,N_5664);
xnor U7507 (N_7507,N_7128,N_6682);
xor U7508 (N_7508,N_5457,N_5881);
nor U7509 (N_7509,N_6897,N_5644);
nand U7510 (N_7510,N_7418,N_6717);
and U7511 (N_7511,N_6183,N_5894);
and U7512 (N_7512,N_6012,N_5365);
and U7513 (N_7513,N_7158,N_5371);
xnor U7514 (N_7514,N_5793,N_6339);
nand U7515 (N_7515,N_5532,N_5452);
or U7516 (N_7516,N_5621,N_5366);
nor U7517 (N_7517,N_7412,N_6491);
xnor U7518 (N_7518,N_6790,N_6442);
or U7519 (N_7519,N_6259,N_6818);
nor U7520 (N_7520,N_7453,N_6011);
or U7521 (N_7521,N_6692,N_5542);
and U7522 (N_7522,N_5979,N_7360);
nor U7523 (N_7523,N_7087,N_6546);
nor U7524 (N_7524,N_5562,N_5607);
nand U7525 (N_7525,N_7182,N_6310);
or U7526 (N_7526,N_5787,N_5079);
or U7527 (N_7527,N_7094,N_6593);
xor U7528 (N_7528,N_5159,N_5520);
xnor U7529 (N_7529,N_6410,N_7068);
nand U7530 (N_7530,N_7099,N_5250);
nand U7531 (N_7531,N_6788,N_5011);
nand U7532 (N_7532,N_7344,N_7476);
nor U7533 (N_7533,N_7466,N_5473);
xnor U7534 (N_7534,N_7407,N_6465);
or U7535 (N_7535,N_6726,N_7145);
or U7536 (N_7536,N_7186,N_5505);
xnor U7537 (N_7537,N_5025,N_5261);
xor U7538 (N_7538,N_5047,N_5210);
or U7539 (N_7539,N_7486,N_5102);
nor U7540 (N_7540,N_6062,N_5593);
nand U7541 (N_7541,N_5557,N_7148);
nor U7542 (N_7542,N_6904,N_5627);
nand U7543 (N_7543,N_5746,N_5412);
or U7544 (N_7544,N_7093,N_5563);
xnor U7545 (N_7545,N_6940,N_5437);
nand U7546 (N_7546,N_6802,N_5928);
nand U7547 (N_7547,N_5356,N_5839);
nand U7548 (N_7548,N_7084,N_6283);
xnor U7549 (N_7549,N_6101,N_6582);
or U7550 (N_7550,N_6943,N_6068);
nand U7551 (N_7551,N_6650,N_6051);
nor U7552 (N_7552,N_5551,N_7440);
and U7553 (N_7553,N_6378,N_5554);
nor U7554 (N_7554,N_7107,N_5495);
and U7555 (N_7555,N_7312,N_5483);
or U7556 (N_7556,N_7210,N_6519);
nand U7557 (N_7557,N_5260,N_6120);
and U7558 (N_7558,N_6233,N_7115);
xor U7559 (N_7559,N_5704,N_6347);
or U7560 (N_7560,N_6876,N_6874);
nor U7561 (N_7561,N_6426,N_7484);
nand U7562 (N_7562,N_6178,N_7199);
nor U7563 (N_7563,N_7421,N_6969);
nand U7564 (N_7564,N_6390,N_6646);
nand U7565 (N_7565,N_6782,N_7361);
nor U7566 (N_7566,N_6270,N_7386);
and U7567 (N_7567,N_7005,N_6679);
or U7568 (N_7568,N_5837,N_6321);
nand U7569 (N_7569,N_7159,N_6805);
xor U7570 (N_7570,N_6461,N_6733);
nand U7571 (N_7571,N_5934,N_6439);
nand U7572 (N_7572,N_7037,N_7039);
xor U7573 (N_7573,N_6708,N_5340);
and U7574 (N_7574,N_7358,N_6255);
nor U7575 (N_7575,N_6988,N_6136);
and U7576 (N_7576,N_5286,N_6866);
nor U7577 (N_7577,N_5216,N_6604);
and U7578 (N_7578,N_5058,N_5758);
nand U7579 (N_7579,N_5135,N_7350);
and U7580 (N_7580,N_6325,N_6087);
nand U7581 (N_7581,N_6873,N_5060);
or U7582 (N_7582,N_5416,N_7002);
nand U7583 (N_7583,N_5139,N_6592);
nand U7584 (N_7584,N_7097,N_6365);
and U7585 (N_7585,N_7056,N_5475);
nand U7586 (N_7586,N_7315,N_6205);
nand U7587 (N_7587,N_5622,N_6481);
nor U7588 (N_7588,N_5099,N_5873);
or U7589 (N_7589,N_7130,N_5893);
nor U7590 (N_7590,N_5158,N_7473);
and U7591 (N_7591,N_7262,N_7222);
or U7592 (N_7592,N_5041,N_6318);
nand U7593 (N_7593,N_6272,N_5512);
or U7594 (N_7594,N_6114,N_6375);
xnor U7595 (N_7595,N_5543,N_5635);
xor U7596 (N_7596,N_6888,N_7241);
nor U7597 (N_7597,N_6655,N_5212);
or U7598 (N_7598,N_5978,N_5737);
and U7599 (N_7599,N_6963,N_7025);
nand U7600 (N_7600,N_6337,N_5026);
xor U7601 (N_7601,N_6497,N_6852);
or U7602 (N_7602,N_5461,N_6349);
and U7603 (N_7603,N_6847,N_5775);
and U7604 (N_7604,N_5249,N_5633);
xnor U7605 (N_7605,N_6033,N_5043);
or U7606 (N_7606,N_5790,N_5224);
nor U7607 (N_7607,N_5784,N_5830);
and U7608 (N_7608,N_5929,N_6206);
nor U7609 (N_7609,N_6853,N_6746);
nand U7610 (N_7610,N_5966,N_6532);
nor U7611 (N_7611,N_5377,N_7401);
xnor U7612 (N_7612,N_5391,N_5832);
or U7613 (N_7613,N_5357,N_5811);
or U7614 (N_7614,N_7024,N_7220);
and U7615 (N_7615,N_6602,N_6773);
and U7616 (N_7616,N_6299,N_7328);
or U7617 (N_7617,N_6596,N_6117);
nor U7618 (N_7618,N_5252,N_5151);
nor U7619 (N_7619,N_6258,N_5730);
nand U7620 (N_7620,N_5770,N_5574);
nand U7621 (N_7621,N_5062,N_5676);
or U7622 (N_7622,N_7474,N_6524);
nor U7623 (N_7623,N_5021,N_6486);
xor U7624 (N_7624,N_6251,N_5338);
nor U7625 (N_7625,N_5820,N_6909);
nor U7626 (N_7626,N_5748,N_5480);
nor U7627 (N_7627,N_7051,N_6515);
and U7628 (N_7628,N_5068,N_6413);
nor U7629 (N_7629,N_7032,N_5354);
or U7630 (N_7630,N_6950,N_6577);
xor U7631 (N_7631,N_6621,N_5853);
and U7632 (N_7632,N_6396,N_6828);
nand U7633 (N_7633,N_7425,N_5997);
nor U7634 (N_7634,N_5687,N_7252);
and U7635 (N_7635,N_5383,N_6742);
or U7636 (N_7636,N_6706,N_5118);
or U7637 (N_7637,N_6774,N_6531);
or U7638 (N_7638,N_5465,N_6080);
or U7639 (N_7639,N_7485,N_5258);
nand U7640 (N_7640,N_6077,N_6694);
nand U7641 (N_7641,N_5555,N_5481);
nand U7642 (N_7642,N_6130,N_7430);
nor U7643 (N_7643,N_5828,N_5855);
or U7644 (N_7644,N_5903,N_5314);
nand U7645 (N_7645,N_6228,N_5821);
or U7646 (N_7646,N_7157,N_6883);
or U7647 (N_7647,N_5972,N_7233);
xor U7648 (N_7648,N_6579,N_6766);
or U7649 (N_7649,N_6956,N_7487);
nand U7650 (N_7650,N_7433,N_6690);
nand U7651 (N_7651,N_6118,N_5292);
or U7652 (N_7652,N_6202,N_6970);
nor U7653 (N_7653,N_5439,N_5304);
nor U7654 (N_7654,N_6158,N_5895);
and U7655 (N_7655,N_5991,N_6074);
nand U7656 (N_7656,N_7050,N_6722);
nor U7657 (N_7657,N_6744,N_5612);
nand U7658 (N_7658,N_6350,N_5493);
nor U7659 (N_7659,N_5003,N_6552);
or U7660 (N_7660,N_7392,N_6464);
nor U7661 (N_7661,N_6826,N_6609);
nand U7662 (N_7662,N_6584,N_5231);
nand U7663 (N_7663,N_7388,N_6105);
or U7664 (N_7664,N_6199,N_5975);
and U7665 (N_7665,N_5398,N_6787);
and U7666 (N_7666,N_5333,N_5275);
nor U7667 (N_7667,N_7065,N_6567);
and U7668 (N_7668,N_5606,N_6324);
nor U7669 (N_7669,N_5908,N_5980);
or U7670 (N_7670,N_5950,N_6400);
nand U7671 (N_7671,N_5846,N_5992);
and U7672 (N_7672,N_6835,N_5120);
nand U7673 (N_7673,N_5132,N_7397);
xnor U7674 (N_7674,N_6044,N_5201);
nor U7675 (N_7675,N_5157,N_6658);
or U7676 (N_7676,N_6174,N_6395);
or U7677 (N_7677,N_6222,N_6974);
and U7678 (N_7678,N_6285,N_6588);
and U7679 (N_7679,N_7022,N_7045);
and U7680 (N_7680,N_6132,N_7383);
and U7681 (N_7681,N_6030,N_7150);
or U7682 (N_7682,N_7411,N_5088);
and U7683 (N_7683,N_7490,N_6242);
nor U7684 (N_7684,N_7209,N_5299);
nand U7685 (N_7685,N_5051,N_6751);
nor U7686 (N_7686,N_5358,N_5080);
and U7687 (N_7687,N_5500,N_6081);
or U7688 (N_7688,N_6700,N_7413);
nand U7689 (N_7689,N_7238,N_5022);
and U7690 (N_7690,N_6180,N_7446);
or U7691 (N_7691,N_6487,N_7213);
and U7692 (N_7692,N_6260,N_5032);
and U7693 (N_7693,N_6034,N_5145);
or U7694 (N_7694,N_6121,N_7492);
xnor U7695 (N_7695,N_5152,N_5564);
nor U7696 (N_7696,N_6201,N_6868);
nand U7697 (N_7697,N_5423,N_5293);
nand U7698 (N_7698,N_6143,N_5061);
or U7699 (N_7699,N_5541,N_6411);
nand U7700 (N_7700,N_5812,N_6468);
nand U7701 (N_7701,N_5824,N_6794);
and U7702 (N_7702,N_5727,N_5097);
and U7703 (N_7703,N_5565,N_5795);
and U7704 (N_7704,N_6610,N_5497);
nor U7705 (N_7705,N_6389,N_6110);
and U7706 (N_7706,N_6735,N_6102);
nor U7707 (N_7707,N_6561,N_5107);
nand U7708 (N_7708,N_7147,N_6959);
and U7709 (N_7709,N_7330,N_6470);
and U7710 (N_7710,N_6359,N_5408);
and U7711 (N_7711,N_6098,N_6225);
nor U7712 (N_7712,N_5295,N_6765);
and U7713 (N_7713,N_6368,N_6212);
or U7714 (N_7714,N_6053,N_5754);
nor U7715 (N_7715,N_6998,N_5989);
and U7716 (N_7716,N_6329,N_6428);
nor U7717 (N_7717,N_5174,N_6553);
nor U7718 (N_7718,N_6477,N_7414);
nand U7719 (N_7719,N_5888,N_7160);
or U7720 (N_7720,N_5091,N_5230);
nand U7721 (N_7721,N_5937,N_7038);
nand U7722 (N_7722,N_7390,N_5678);
nor U7723 (N_7723,N_6923,N_6846);
nor U7724 (N_7724,N_7028,N_6691);
or U7725 (N_7725,N_6684,N_5605);
nand U7726 (N_7726,N_7156,N_6328);
nand U7727 (N_7727,N_6387,N_5932);
xnor U7728 (N_7728,N_5350,N_6719);
nand U7729 (N_7729,N_5288,N_6695);
or U7730 (N_7730,N_6887,N_5381);
or U7731 (N_7731,N_5342,N_6469);
and U7732 (N_7732,N_5679,N_6831);
and U7733 (N_7733,N_5947,N_6024);
nand U7734 (N_7734,N_5692,N_6799);
nand U7735 (N_7735,N_6416,N_7498);
or U7736 (N_7736,N_6176,N_6891);
nand U7737 (N_7737,N_6287,N_7030);
and U7738 (N_7738,N_6508,N_6715);
nor U7739 (N_7739,N_6431,N_5889);
and U7740 (N_7740,N_5836,N_7279);
nor U7741 (N_7741,N_5269,N_6987);
or U7742 (N_7742,N_5037,N_5769);
and U7743 (N_7743,N_6376,N_5583);
xor U7744 (N_7744,N_5259,N_5626);
or U7745 (N_7745,N_7172,N_7363);
and U7746 (N_7746,N_5504,N_6560);
nand U7747 (N_7747,N_7482,N_6642);
or U7748 (N_7748,N_5582,N_5104);
nand U7749 (N_7749,N_6947,N_7206);
nand U7750 (N_7750,N_7019,N_6358);
or U7751 (N_7751,N_7137,N_7333);
and U7752 (N_7752,N_7455,N_5789);
nand U7753 (N_7753,N_5432,N_5421);
or U7754 (N_7754,N_6478,N_5267);
nand U7755 (N_7755,N_5890,N_5148);
nor U7756 (N_7756,N_5200,N_7410);
xor U7757 (N_7757,N_7085,N_6342);
nand U7758 (N_7758,N_6764,N_6209);
or U7759 (N_7759,N_7426,N_6574);
nor U7760 (N_7760,N_5345,N_6908);
or U7761 (N_7761,N_5486,N_6374);
or U7762 (N_7762,N_5835,N_5209);
nor U7763 (N_7763,N_7185,N_5388);
and U7764 (N_7764,N_7408,N_5326);
nor U7765 (N_7765,N_5444,N_6274);
nand U7766 (N_7766,N_6433,N_5013);
or U7767 (N_7767,N_5154,N_6076);
nand U7768 (N_7768,N_6443,N_5919);
nand U7769 (N_7769,N_5925,N_7048);
and U7770 (N_7770,N_7323,N_7459);
nor U7771 (N_7771,N_6747,N_5904);
nand U7772 (N_7772,N_7309,N_5144);
and U7773 (N_7773,N_6606,N_6140);
nand U7774 (N_7774,N_5023,N_5066);
xnor U7775 (N_7775,N_5623,N_5017);
or U7776 (N_7776,N_7292,N_6529);
nand U7777 (N_7777,N_6919,N_5175);
and U7778 (N_7778,N_5865,N_7174);
and U7779 (N_7779,N_6814,N_5279);
nand U7780 (N_7780,N_5192,N_5988);
or U7781 (N_7781,N_7378,N_5346);
nor U7782 (N_7782,N_5323,N_5560);
and U7783 (N_7783,N_7140,N_7236);
nor U7784 (N_7784,N_6123,N_6311);
nor U7785 (N_7785,N_5938,N_6902);
nand U7786 (N_7786,N_6598,N_5916);
or U7787 (N_7787,N_7111,N_6775);
nor U7788 (N_7788,N_5092,N_6649);
and U7789 (N_7789,N_5777,N_6677);
or U7790 (N_7790,N_5579,N_5616);
or U7791 (N_7791,N_6388,N_7117);
xor U7792 (N_7792,N_5270,N_6009);
nand U7793 (N_7793,N_5866,N_6944);
and U7794 (N_7794,N_6391,N_6644);
nand U7795 (N_7795,N_6371,N_7235);
nor U7796 (N_7796,N_6289,N_5643);
nor U7797 (N_7797,N_5031,N_6513);
nor U7798 (N_7798,N_5363,N_6097);
nor U7799 (N_7799,N_5352,N_7127);
or U7800 (N_7800,N_6983,N_6405);
or U7801 (N_7801,N_6301,N_7034);
and U7802 (N_7802,N_6126,N_5768);
nand U7803 (N_7803,N_6137,N_7366);
or U7804 (N_7804,N_5734,N_5089);
xor U7805 (N_7805,N_5669,N_5923);
xnor U7806 (N_7806,N_5009,N_6031);
nand U7807 (N_7807,N_5785,N_6793);
xnor U7808 (N_7808,N_5162,N_6162);
or U7809 (N_7809,N_6674,N_6160);
or U7810 (N_7810,N_5983,N_5530);
nand U7811 (N_7811,N_7201,N_6084);
nand U7812 (N_7812,N_5861,N_5180);
nand U7813 (N_7813,N_7198,N_6938);
or U7814 (N_7814,N_5306,N_5113);
xor U7815 (N_7815,N_5732,N_6122);
nor U7816 (N_7816,N_6166,N_6727);
or U7817 (N_7817,N_7188,N_5055);
and U7818 (N_7818,N_7475,N_6641);
xnor U7819 (N_7819,N_6996,N_5915);
xnor U7820 (N_7820,N_5722,N_5321);
nand U7821 (N_7821,N_6952,N_6568);
nor U7822 (N_7822,N_6862,N_6709);
xor U7823 (N_7823,N_6293,N_6770);
nor U7824 (N_7824,N_5545,N_6640);
xor U7825 (N_7825,N_5524,N_5040);
or U7826 (N_7826,N_7000,N_5467);
or U7827 (N_7827,N_6037,N_6666);
and U7828 (N_7828,N_7122,N_6066);
xnor U7829 (N_7829,N_5632,N_6172);
or U7830 (N_7830,N_6955,N_5278);
nand U7831 (N_7831,N_5519,N_6247);
nor U7832 (N_7832,N_6179,N_6454);
nor U7833 (N_7833,N_5984,N_7340);
nand U7834 (N_7834,N_5870,N_6981);
nor U7835 (N_7835,N_5999,N_6984);
nor U7836 (N_7836,N_6762,N_5940);
and U7837 (N_7837,N_5169,N_5459);
and U7838 (N_7838,N_7095,N_6860);
xor U7839 (N_7839,N_5472,N_5792);
and U7840 (N_7840,N_5466,N_7217);
and U7841 (N_7841,N_6131,N_6982);
or U7842 (N_7842,N_7332,N_5651);
xor U7843 (N_7843,N_6334,N_7405);
and U7844 (N_7844,N_7165,N_5624);
nor U7845 (N_7845,N_5375,N_6190);
nor U7846 (N_7846,N_6406,N_6525);
or U7847 (N_7847,N_5711,N_7176);
and U7848 (N_7848,N_6894,N_6834);
nor U7849 (N_7849,N_6925,N_6619);
and U7850 (N_7850,N_6056,N_6444);
nand U7851 (N_7851,N_5313,N_6065);
xor U7852 (N_7852,N_7265,N_6276);
or U7853 (N_7853,N_5911,N_6488);
xor U7854 (N_7854,N_5167,N_6335);
nand U7855 (N_7855,N_6936,N_7371);
and U7856 (N_7856,N_5924,N_7073);
nor U7857 (N_7857,N_6699,N_7288);
or U7858 (N_7858,N_5993,N_6555);
and U7859 (N_7859,N_6346,N_6545);
nor U7860 (N_7860,N_5447,N_5968);
nor U7861 (N_7861,N_5203,N_5712);
xor U7862 (N_7862,N_6718,N_5335);
nand U7863 (N_7863,N_5619,N_6435);
xnor U7864 (N_7864,N_6345,N_5134);
or U7865 (N_7865,N_6587,N_5713);
or U7866 (N_7866,N_6383,N_6502);
and U7867 (N_7867,N_5569,N_6824);
xnor U7868 (N_7868,N_7444,N_5109);
nand U7869 (N_7869,N_5006,N_5182);
and U7870 (N_7870,N_6257,N_7370);
nor U7871 (N_7871,N_6882,N_5397);
nor U7872 (N_7872,N_6784,N_7055);
and U7873 (N_7873,N_7049,N_7373);
or U7874 (N_7874,N_7494,N_7460);
nor U7875 (N_7875,N_5309,N_7003);
or U7876 (N_7876,N_6188,N_6948);
or U7877 (N_7877,N_7356,N_6573);
and U7878 (N_7878,N_5106,N_6939);
nor U7879 (N_7879,N_6341,N_6861);
and U7880 (N_7880,N_6421,N_7403);
or U7881 (N_7881,N_5069,N_6798);
xor U7882 (N_7882,N_5587,N_6119);
or U7883 (N_7883,N_5410,N_5016);
or U7884 (N_7884,N_7479,N_5723);
nor U7885 (N_7885,N_5078,N_5589);
and U7886 (N_7886,N_5816,N_6091);
nand U7887 (N_7887,N_6332,N_7195);
nor U7888 (N_7888,N_5523,N_5553);
nor U7889 (N_7889,N_5905,N_6548);
or U7890 (N_7890,N_7318,N_7074);
nor U7891 (N_7891,N_5096,N_6991);
nand U7892 (N_7892,N_6063,N_5755);
or U7893 (N_7893,N_7106,N_7406);
nor U7894 (N_7894,N_5537,N_6937);
or U7895 (N_7895,N_6778,N_5020);
and U7896 (N_7896,N_5422,N_6189);
nand U7897 (N_7897,N_7493,N_7189);
nor U7898 (N_7898,N_6052,N_5419);
or U7899 (N_7899,N_5232,N_6154);
nor U7900 (N_7900,N_5931,N_5053);
xor U7901 (N_7901,N_6701,N_6271);
and U7902 (N_7902,N_7242,N_5030);
or U7903 (N_7903,N_5456,N_6385);
or U7904 (N_7904,N_5933,N_7221);
and U7905 (N_7905,N_6485,N_6075);
nand U7906 (N_7906,N_7146,N_5747);
xor U7907 (N_7907,N_7230,N_5566);
and U7908 (N_7908,N_5220,N_6711);
xnor U7909 (N_7909,N_5945,N_6683);
nor U7910 (N_7910,N_5625,N_7278);
and U7911 (N_7911,N_5202,N_6792);
nor U7912 (N_7912,N_5875,N_5525);
and U7913 (N_7913,N_7187,N_6246);
nand U7914 (N_7914,N_6195,N_5906);
and U7915 (N_7915,N_7178,N_5477);
or U7916 (N_7916,N_5852,N_6403);
and U7917 (N_7917,N_6038,N_6017);
and U7918 (N_7918,N_5160,N_5415);
or U7919 (N_7919,N_5094,N_7274);
nand U7920 (N_7920,N_6392,N_5897);
nand U7921 (N_7921,N_6356,N_5349);
nand U7922 (N_7922,N_5909,N_5194);
or U7923 (N_7923,N_6005,N_6243);
nand U7924 (N_7924,N_6554,N_5036);
nand U7925 (N_7925,N_6526,N_5280);
and U7926 (N_7926,N_5510,N_7169);
and U7927 (N_7927,N_5018,N_5307);
or U7928 (N_7928,N_6330,N_5329);
nand U7929 (N_7929,N_7175,N_6864);
and U7930 (N_7930,N_7273,N_5764);
nor U7931 (N_7931,N_6369,N_5590);
nor U7932 (N_7932,N_7181,N_5070);
or U7933 (N_7933,N_6463,N_5315);
and U7934 (N_7934,N_6661,N_5050);
nand U7935 (N_7935,N_5900,N_7144);
nor U7936 (N_7936,N_5281,N_5038);
nor U7937 (N_7937,N_6354,N_5806);
or U7938 (N_7938,N_5400,N_6501);
and U7939 (N_7939,N_6856,N_6879);
or U7940 (N_7940,N_5650,N_6550);
and U7941 (N_7941,N_5652,N_6541);
nand U7942 (N_7942,N_5186,N_5516);
or U7943 (N_7943,N_6112,N_7070);
and U7944 (N_7944,N_5600,N_5656);
nor U7945 (N_7945,N_5610,N_5077);
or U7946 (N_7946,N_7064,N_5059);
or U7947 (N_7947,N_6720,N_6924);
or U7948 (N_7948,N_7372,N_5247);
nand U7949 (N_7949,N_7355,N_5885);
nor U7950 (N_7950,N_6379,N_5739);
xor U7951 (N_7951,N_6263,N_7286);
nor U7952 (N_7952,N_7012,N_5319);
and U7953 (N_7953,N_7109,N_5255);
nor U7954 (N_7954,N_6521,N_6838);
nor U7955 (N_7955,N_5659,N_5482);
and U7956 (N_7956,N_6752,N_7452);
nor U7957 (N_7957,N_7325,N_6054);
or U7958 (N_7958,N_5411,N_6971);
nand U7959 (N_7959,N_7125,N_5228);
nand U7960 (N_7960,N_5597,N_6815);
nand U7961 (N_7961,N_5085,N_6945);
nor U7962 (N_7962,N_6801,N_6280);
nand U7963 (N_7963,N_6533,N_7173);
or U7964 (N_7964,N_7123,N_5474);
nand U7965 (N_7965,N_5527,N_6833);
and U7966 (N_7966,N_7326,N_6926);
or U7967 (N_7967,N_5296,N_6922);
and U7968 (N_7968,N_6353,N_5027);
and U7969 (N_7969,N_6322,N_6193);
or U7970 (N_7970,N_6522,N_5233);
xnor U7971 (N_7971,N_6472,N_6331);
nand U7972 (N_7972,N_7257,N_6394);
nand U7973 (N_7973,N_7020,N_6373);
xor U7974 (N_7974,N_5108,N_5362);
nand U7975 (N_7975,N_6039,N_6156);
nor U7976 (N_7976,N_6725,N_6680);
or U7977 (N_7977,N_5353,N_6820);
nor U7978 (N_7978,N_6839,N_5998);
nand U7979 (N_7979,N_5813,N_5334);
xnor U7980 (N_7980,N_6127,N_7054);
and U7981 (N_7981,N_7008,N_5215);
and U7982 (N_7982,N_6608,N_7141);
nor U7983 (N_7983,N_6721,N_5491);
nand U7984 (N_7984,N_5891,N_6500);
and U7985 (N_7985,N_5567,N_5462);
and U7986 (N_7986,N_6419,N_5172);
or U7987 (N_7987,N_6671,N_6370);
or U7988 (N_7988,N_7359,N_6806);
nor U7989 (N_7989,N_6058,N_6138);
and U7990 (N_7990,N_7081,N_5508);
or U7991 (N_7991,N_6363,N_5985);
and U7992 (N_7992,N_6191,N_5742);
xor U7993 (N_7993,N_5434,N_7184);
nand U7994 (N_7994,N_6418,N_7083);
nand U7995 (N_7995,N_7489,N_6015);
or U7996 (N_7996,N_6352,N_5485);
and U7997 (N_7997,N_5318,N_6638);
and U7998 (N_7998,N_6729,N_7052);
nor U7999 (N_7999,N_5170,N_6456);
or U8000 (N_8000,N_7367,N_6106);
and U8001 (N_8001,N_6895,N_5936);
nand U8002 (N_8002,N_5418,N_6633);
nand U8003 (N_8003,N_7416,N_6070);
and U8004 (N_8004,N_7004,N_6253);
nand U8005 (N_8005,N_7409,N_5778);
nand U8006 (N_8006,N_6007,N_5431);
or U8007 (N_8007,N_6576,N_7302);
xor U8008 (N_8008,N_6850,N_6791);
nor U8009 (N_8009,N_5901,N_6103);
and U8010 (N_8010,N_6266,N_5324);
or U8011 (N_8011,N_5517,N_6279);
nand U8012 (N_8012,N_5219,N_5673);
or U8013 (N_8013,N_5862,N_5995);
and U8014 (N_8014,N_7481,N_6064);
or U8015 (N_8015,N_5725,N_5436);
and U8016 (N_8016,N_6543,N_5005);
nor U8017 (N_8017,N_7297,N_5767);
nor U8018 (N_8018,N_6900,N_5445);
or U8019 (N_8019,N_6256,N_6635);
and U8020 (N_8020,N_5166,N_6047);
nand U8021 (N_8021,N_6249,N_5251);
nand U8022 (N_8022,N_6211,N_6230);
nand U8023 (N_8023,N_5399,N_5996);
and U8024 (N_8024,N_5347,N_5283);
xor U8025 (N_8025,N_6600,N_5034);
nand U8026 (N_8026,N_7245,N_5981);
nor U8027 (N_8027,N_6207,N_6819);
nand U8028 (N_8028,N_7454,N_7240);
nor U8029 (N_8029,N_6284,N_5601);
or U8030 (N_8030,N_6286,N_5098);
xor U8031 (N_8031,N_7429,N_5407);
nor U8032 (N_8032,N_5765,N_5187);
and U8033 (N_8033,N_5954,N_5488);
xor U8034 (N_8034,N_5689,N_6905);
or U8035 (N_8035,N_5838,N_5876);
and U8036 (N_8036,N_5124,N_5064);
or U8037 (N_8037,N_5774,N_6504);
and U8038 (N_8038,N_5749,N_5239);
xnor U8039 (N_8039,N_5404,N_6026);
and U8040 (N_8040,N_7301,N_6763);
nand U8041 (N_8041,N_5648,N_6689);
or U8042 (N_8042,N_5805,N_6636);
or U8043 (N_8043,N_6961,N_6264);
nor U8044 (N_8044,N_7192,N_6615);
or U8045 (N_8045,N_6386,N_6223);
nor U8046 (N_8046,N_6150,N_7177);
nor U8047 (N_8047,N_7098,N_5766);
nor U8048 (N_8048,N_6238,N_6498);
nand U8049 (N_8049,N_5243,N_5642);
nor U8050 (N_8050,N_5300,N_6898);
nor U8051 (N_8051,N_5744,N_5463);
or U8052 (N_8052,N_5577,N_5912);
and U8053 (N_8053,N_6046,N_5604);
nor U8054 (N_8054,N_6153,N_5887);
nand U8055 (N_8055,N_6716,N_5277);
or U8056 (N_8056,N_5763,N_7225);
nor U8057 (N_8057,N_7033,N_5552);
and U8058 (N_8058,N_6029,N_6673);
nand U8059 (N_8059,N_7080,N_5959);
nor U8060 (N_8060,N_6273,N_5762);
nor U8061 (N_8061,N_5244,N_5694);
and U8062 (N_8062,N_6186,N_5568);
nor U8063 (N_8063,N_7226,N_6612);
xnor U8064 (N_8064,N_5608,N_5428);
nand U8065 (N_8065,N_7155,N_5443);
nand U8066 (N_8066,N_5561,N_7223);
or U8067 (N_8067,N_5745,N_5207);
or U8068 (N_8068,N_6523,N_7331);
nor U8069 (N_8069,N_6780,N_6441);
xnor U8070 (N_8070,N_6962,N_5798);
and U8071 (N_8071,N_6237,N_6489);
and U8072 (N_8072,N_6965,N_6759);
nand U8073 (N_8073,N_5116,N_5235);
and U8074 (N_8074,N_5921,N_6155);
nor U8075 (N_8075,N_5348,N_5298);
xor U8076 (N_8076,N_7357,N_5044);
nor U8077 (N_8077,N_5425,N_6544);
xnor U8078 (N_8078,N_6366,N_5958);
and U8079 (N_8079,N_5514,N_5653);
nor U8080 (N_8080,N_7171,N_7284);
nand U8081 (N_8081,N_7399,N_5849);
nand U8082 (N_8082,N_6424,N_6096);
or U8083 (N_8083,N_7431,N_7291);
nand U8084 (N_8084,N_5826,N_6845);
or U8085 (N_8085,N_5438,N_6315);
nand U8086 (N_8086,N_6736,N_6306);
and U8087 (N_8087,N_7007,N_5690);
nand U8088 (N_8088,N_7354,N_6645);
nor U8089 (N_8089,N_6250,N_7041);
nor U8090 (N_8090,N_7380,N_6417);
or U8091 (N_8091,N_6298,N_6045);
or U8092 (N_8092,N_6509,N_6147);
and U8093 (N_8093,N_5803,N_7320);
and U8094 (N_8094,N_5442,N_5533);
nor U8095 (N_8095,N_6865,N_6571);
nor U8096 (N_8096,N_6139,N_5639);
nor U8097 (N_8097,N_5378,N_7329);
nand U8098 (N_8098,N_7439,N_7472);
or U8099 (N_8099,N_6482,N_6564);
nand U8100 (N_8100,N_5095,N_6234);
and U8101 (N_8101,N_7462,N_5101);
or U8102 (N_8102,N_6483,N_5580);
or U8103 (N_8103,N_7419,N_6152);
and U8104 (N_8104,N_7365,N_6239);
and U8105 (N_8105,N_6466,N_5355);
and U8106 (N_8106,N_6040,N_7310);
or U8107 (N_8107,N_7076,N_5188);
or U8108 (N_8108,N_7402,N_5128);
and U8109 (N_8109,N_6397,N_6910);
and U8110 (N_8110,N_7134,N_5173);
or U8111 (N_8111,N_5301,N_7483);
xor U8112 (N_8112,N_5864,N_5290);
or U8113 (N_8113,N_7232,N_7143);
or U8114 (N_8114,N_5071,N_5149);
and U8115 (N_8115,N_5655,N_5430);
nand U8116 (N_8116,N_6723,N_6986);
or U8117 (N_8117,N_6412,N_5930);
and U8118 (N_8118,N_6021,N_6113);
nand U8119 (N_8119,N_5282,N_6771);
xnor U8120 (N_8120,N_7069,N_7131);
nand U8121 (N_8121,N_5237,N_6167);
nand U8122 (N_8122,N_6294,N_5658);
and U8123 (N_8123,N_5696,N_5316);
or U8124 (N_8124,N_6623,N_5024);
or U8125 (N_8125,N_6569,N_6927);
and U8126 (N_8126,N_7319,N_5759);
nor U8127 (N_8127,N_6336,N_5654);
or U8128 (N_8128,N_5274,N_5799);
nand U8129 (N_8129,N_5714,N_6929);
nand U8130 (N_8130,N_5303,N_7423);
nor U8131 (N_8131,N_6881,N_7061);
nand U8132 (N_8132,N_5592,N_5122);
and U8133 (N_8133,N_5081,N_5910);
nand U8134 (N_8134,N_6398,N_7264);
nand U8135 (N_8135,N_6618,N_5402);
and U8136 (N_8136,N_5715,N_5364);
and U8137 (N_8137,N_5453,N_5361);
and U8138 (N_8138,N_6681,N_6244);
and U8139 (N_8139,N_6572,N_7465);
nand U8140 (N_8140,N_5208,N_7138);
nand U8141 (N_8141,N_5082,N_7368);
nor U8142 (N_8142,N_5121,N_5424);
or U8143 (N_8143,N_7449,N_5503);
nor U8144 (N_8144,N_5177,N_7112);
nand U8145 (N_8145,N_5140,N_5974);
nand U8146 (N_8146,N_6305,N_7108);
or U8147 (N_8147,N_5773,N_5218);
and U8148 (N_8148,N_5693,N_6932);
or U8149 (N_8149,N_6967,N_5343);
or U8150 (N_8150,N_5728,N_5229);
xnor U8151 (N_8151,N_6652,N_6617);
and U8152 (N_8152,N_5686,N_7227);
and U8153 (N_8153,N_7343,N_5253);
nand U8154 (N_8154,N_7170,N_6148);
and U8155 (N_8155,N_5528,N_5858);
or U8156 (N_8156,N_7254,N_6539);
or U8157 (N_8157,N_5596,N_6093);
or U8158 (N_8158,N_6333,N_5575);
xor U8159 (N_8159,N_6758,N_7258);
nor U8160 (N_8160,N_6078,N_7251);
or U8161 (N_8161,N_7161,N_5441);
nor U8162 (N_8162,N_6855,N_7287);
nand U8163 (N_8163,N_6808,N_6480);
xor U8164 (N_8164,N_6226,N_5147);
nor U8165 (N_8165,N_6267,N_6990);
nor U8166 (N_8166,N_7092,N_5076);
and U8167 (N_8167,N_7334,N_5753);
xor U8168 (N_8168,N_6060,N_6703);
nand U8169 (N_8169,N_6367,N_6614);
nor U8170 (N_8170,N_6807,N_5123);
nand U8171 (N_8171,N_6338,N_6999);
nand U8172 (N_8172,N_6595,N_5957);
nor U8173 (N_8173,N_6023,N_5234);
nand U8174 (N_8174,N_7339,N_7077);
and U8175 (N_8175,N_7324,N_5691);
and U8176 (N_8176,N_6854,N_6144);
nor U8177 (N_8177,N_6453,N_5531);
xnor U8178 (N_8178,N_5193,N_5586);
and U8179 (N_8179,N_6756,N_7015);
nor U8180 (N_8180,N_6008,N_5886);
and U8181 (N_8181,N_6710,N_7247);
nand U8182 (N_8182,N_5196,N_5526);
and U8183 (N_8183,N_5794,N_7432);
nand U8184 (N_8184,N_7029,N_5360);
and U8185 (N_8185,N_5743,N_7001);
nor U8186 (N_8186,N_7266,N_7389);
or U8187 (N_8187,N_6857,N_5289);
or U8188 (N_8188,N_5199,N_6813);
nor U8189 (N_8189,N_7424,N_6810);
or U8190 (N_8190,N_6740,N_7395);
or U8191 (N_8191,N_7103,N_6889);
nor U8192 (N_8192,N_6878,N_6627);
or U8193 (N_8193,N_6559,N_6921);
nand U8194 (N_8194,N_5922,N_6197);
and U8195 (N_8195,N_7194,N_7151);
nand U8196 (N_8196,N_5546,N_7078);
or U8197 (N_8197,N_5489,N_5588);
nand U8198 (N_8198,N_7341,N_5368);
or U8199 (N_8199,N_5529,N_5863);
nor U8200 (N_8200,N_7231,N_5420);
nor U8201 (N_8201,N_7369,N_5409);
nor U8202 (N_8202,N_6302,N_6632);
nor U8203 (N_8203,N_6467,N_6151);
or U8204 (N_8204,N_6240,N_5518);
nand U8205 (N_8205,N_6399,N_6507);
nand U8206 (N_8206,N_5990,N_6743);
xnor U8207 (N_8207,N_5707,N_5522);
xor U8208 (N_8208,N_6979,N_6414);
nor U8209 (N_8209,N_6307,N_5226);
nor U8210 (N_8210,N_5221,N_7322);
nand U8211 (N_8211,N_7491,N_7249);
nand U8212 (N_8212,N_5225,N_6980);
or U8213 (N_8213,N_6171,N_5476);
nand U8214 (N_8214,N_6840,N_5831);
nor U8215 (N_8215,N_6896,N_6953);
xor U8216 (N_8216,N_5584,N_5683);
or U8217 (N_8217,N_5854,N_5513);
nor U8218 (N_8218,N_5322,N_5850);
and U8219 (N_8219,N_6364,N_6997);
or U8220 (N_8220,N_6934,N_6002);
nand U8221 (N_8221,N_7382,N_6558);
or U8222 (N_8222,N_7463,N_6750);
and U8223 (N_8223,N_6479,N_7471);
nand U8224 (N_8224,N_6675,N_5502);
or U8225 (N_8225,N_6432,N_5660);
nor U8226 (N_8226,N_5268,N_6510);
nand U8227 (N_8227,N_7289,N_5750);
nor U8228 (N_8228,N_6812,N_5857);
or U8229 (N_8229,N_5840,N_6978);
nand U8230 (N_8230,N_6004,N_5291);
or U8231 (N_8231,N_6685,N_7035);
and U8232 (N_8232,N_5718,N_6754);
nor U8233 (N_8233,N_7443,N_5920);
and U8234 (N_8234,N_6503,N_5521);
nand U8235 (N_8235,N_5090,N_5636);
or U8236 (N_8236,N_7311,N_5956);
nor U8237 (N_8237,N_7089,N_6591);
and U8238 (N_8238,N_5386,N_5967);
nand U8239 (N_8239,N_5585,N_6935);
and U8240 (N_8240,N_6094,N_5752);
nand U8241 (N_8241,N_5052,N_5287);
nor U8242 (N_8242,N_7277,N_6297);
nor U8243 (N_8243,N_6551,N_7023);
nor U8244 (N_8244,N_5547,N_5851);
nand U8245 (N_8245,N_5771,N_6875);
nand U8246 (N_8246,N_7237,N_5163);
or U8247 (N_8247,N_7229,N_5724);
nor U8248 (N_8248,N_6095,N_5395);
nand U8249 (N_8249,N_6786,N_5982);
xor U8250 (N_8250,N_5164,N_6613);
or U8251 (N_8251,N_5700,N_5131);
nand U8252 (N_8252,N_6800,N_5668);
nor U8253 (N_8253,N_5736,N_6530);
or U8254 (N_8254,N_5918,N_6449);
xor U8255 (N_8255,N_7211,N_6194);
nor U8256 (N_8256,N_6698,N_5074);
and U8257 (N_8257,N_6300,N_7047);
and U8258 (N_8258,N_5136,N_6848);
and U8259 (N_8259,N_5072,N_6916);
nor U8260 (N_8260,N_5550,N_5572);
xor U8261 (N_8261,N_6451,N_5899);
and U8262 (N_8262,N_6995,N_6659);
nand U8263 (N_8263,N_6446,N_5780);
nor U8264 (N_8264,N_6474,N_6964);
nor U8265 (N_8265,N_5227,N_7207);
and U8266 (N_8266,N_6797,N_6484);
nand U8267 (N_8267,N_5369,N_5190);
and U8268 (N_8268,N_5801,N_5661);
and U8269 (N_8269,N_6290,N_7200);
nand U8270 (N_8270,N_6917,N_5100);
nor U8271 (N_8271,N_5191,N_5646);
nand U8272 (N_8272,N_5014,N_7298);
and U8273 (N_8273,N_5786,N_5103);
nor U8274 (N_8274,N_6957,N_6728);
or U8275 (N_8275,N_6538,N_5638);
or U8276 (N_8276,N_6438,N_7377);
and U8277 (N_8277,N_6664,N_5458);
nand U8278 (N_8278,N_6323,N_6662);
nand U8279 (N_8279,N_6867,N_5339);
and U8280 (N_8280,N_6705,N_5702);
nand U8281 (N_8281,N_7391,N_6182);
nor U8282 (N_8282,N_5087,N_6712);
nor U8283 (N_8283,N_7110,N_6676);
or U8284 (N_8284,N_5935,N_5868);
nand U8285 (N_8285,N_7260,N_5137);
nor U8286 (N_8286,N_5454,N_5150);
nand U8287 (N_8287,N_7168,N_6907);
or U8288 (N_8288,N_6562,N_7256);
or U8289 (N_8289,N_7456,N_5682);
nor U8290 (N_8290,N_6304,N_6511);
nand U8291 (N_8291,N_7166,N_7124);
and U8292 (N_8292,N_6265,N_7202);
nand U8293 (N_8293,N_7271,N_5733);
and U8294 (N_8294,N_6288,N_5242);
xor U8295 (N_8295,N_6607,N_6738);
and U8296 (N_8296,N_5130,N_6557);
xnor U8297 (N_8297,N_6415,N_7063);
nand U8298 (N_8298,N_6157,N_5470);
nand U8299 (N_8299,N_5401,N_7290);
and U8300 (N_8300,N_6647,N_6083);
nand U8301 (N_8301,N_6648,N_7299);
or U8302 (N_8302,N_5859,N_5720);
nor U8303 (N_8303,N_6016,N_5845);
and U8304 (N_8304,N_5641,N_5882);
xor U8305 (N_8305,N_6933,N_6817);
xor U8306 (N_8306,N_6877,N_7167);
and U8307 (N_8307,N_7305,N_5663);
nor U8308 (N_8308,N_5238,N_5598);
or U8309 (N_8309,N_6906,N_5305);
and U8310 (N_8310,N_6107,N_6217);
nor U8311 (N_8311,N_6059,N_6816);
nand U8312 (N_8312,N_5819,N_5004);
nor U8313 (N_8313,N_5942,N_7261);
or U8314 (N_8314,N_6252,N_7090);
and U8315 (N_8315,N_7149,N_5331);
nand U8316 (N_8316,N_6380,N_5126);
and U8317 (N_8317,N_5962,N_6372);
nor U8318 (N_8318,N_7269,N_5336);
xnor U8319 (N_8319,N_7121,N_5657);
nand U8320 (N_8320,N_7243,N_6693);
nor U8321 (N_8321,N_5705,N_5847);
xnor U8322 (N_8322,N_5478,N_7387);
or U8323 (N_8323,N_5695,N_6348);
or U8324 (N_8324,N_7384,N_6537);
xor U8325 (N_8325,N_6724,N_5721);
nand U8326 (N_8326,N_5927,N_5223);
nand U8327 (N_8327,N_6145,N_7488);
nand U8328 (N_8328,N_6601,N_6547);
nor U8329 (N_8329,N_7059,N_5468);
xor U8330 (N_8330,N_5028,N_6316);
nand U8331 (N_8331,N_7016,N_6043);
and U8332 (N_8332,N_5083,N_6142);
or U8333 (N_8333,N_5054,N_7120);
nand U8334 (N_8334,N_5084,N_5961);
or U8335 (N_8335,N_7119,N_6384);
xor U8336 (N_8336,N_5902,N_6892);
or U8337 (N_8337,N_7142,N_7129);
nand U8338 (N_8338,N_7393,N_7105);
and U8339 (N_8339,N_6517,N_5818);
nor U8340 (N_8340,N_6804,N_7205);
nand U8341 (N_8341,N_5002,N_7468);
or U8342 (N_8342,N_6913,N_6089);
or U8343 (N_8343,N_6425,N_7057);
nand U8344 (N_8344,N_7480,N_7017);
and U8345 (N_8345,N_5822,N_5571);
and U8346 (N_8346,N_5701,N_5538);
or U8347 (N_8347,N_5241,N_6277);
nor U8348 (N_8348,N_6912,N_6589);
nor U8349 (N_8349,N_6281,N_6050);
and U8350 (N_8350,N_5603,N_5206);
nor U8351 (N_8351,N_6843,N_7104);
nor U8352 (N_8352,N_7218,N_5943);
xor U8353 (N_8353,N_5800,N_7253);
or U8354 (N_8354,N_7248,N_7436);
nand U8355 (N_8355,N_5487,N_6520);
nand U8356 (N_8356,N_6022,N_6823);
xnor U8357 (N_8357,N_5189,N_5256);
nand U8358 (N_8358,N_6629,N_6436);
nand U8359 (N_8359,N_5740,N_7086);
nand U8360 (N_8360,N_6382,N_6317);
nand U8361 (N_8361,N_6518,N_6872);
and U8362 (N_8362,N_5647,N_6493);
and U8363 (N_8363,N_6473,N_5613);
and U8364 (N_8364,N_6181,N_6164);
or U8365 (N_8365,N_6989,N_6975);
xor U8366 (N_8366,N_7031,N_6027);
nor U8367 (N_8367,N_6092,N_5440);
nor U8368 (N_8368,N_5872,N_6796);
nor U8369 (N_8369,N_6458,N_6789);
xnor U8370 (N_8370,N_5195,N_5548);
or U8371 (N_8371,N_7215,N_7133);
nand U8372 (N_8372,N_6170,N_5029);
nor U8373 (N_8373,N_5609,N_6409);
nor U8374 (N_8374,N_5535,N_5370);
nor U8375 (N_8375,N_7272,N_6116);
and U8376 (N_8376,N_5155,N_5977);
or U8377 (N_8377,N_6599,N_6159);
and U8378 (N_8378,N_5117,N_5284);
xnor U8379 (N_8379,N_5848,N_5000);
or U8380 (N_8380,N_6575,N_5302);
nor U8381 (N_8381,N_5198,N_6192);
nand U8382 (N_8382,N_5796,N_7346);
or U8383 (N_8383,N_5595,N_5731);
xnor U8384 (N_8384,N_5540,N_5716);
nand U8385 (N_8385,N_5685,N_5994);
nor U8386 (N_8386,N_5880,N_5662);
nor U8387 (N_8387,N_6656,N_5393);
or U8388 (N_8388,N_7381,N_7259);
and U8389 (N_8389,N_6141,N_6282);
or U8390 (N_8390,N_6018,N_5376);
and U8391 (N_8391,N_5634,N_5614);
nand U8392 (N_8392,N_5165,N_5390);
xnor U8393 (N_8393,N_7018,N_5751);
xnor U8394 (N_8394,N_6309,N_6678);
nand U8395 (N_8395,N_6976,N_7467);
nand U8396 (N_8396,N_7239,N_5973);
nand U8397 (N_8397,N_6781,N_7283);
or U8398 (N_8398,N_5883,N_5620);
or U8399 (N_8399,N_6448,N_5698);
nand U8400 (N_8400,N_5455,N_5896);
or U8401 (N_8401,N_5829,N_6580);
nand U8402 (N_8402,N_6423,N_6404);
and U8403 (N_8403,N_7375,N_6911);
nor U8404 (N_8404,N_5327,N_6447);
nor U8405 (N_8405,N_5761,N_5240);
nor U8406 (N_8406,N_5217,N_7428);
nand U8407 (N_8407,N_6001,N_5257);
or U8408 (N_8408,N_5717,N_6734);
and U8409 (N_8409,N_5631,N_6090);
nand U8410 (N_8410,N_7478,N_7066);
nand U8411 (N_8411,N_5781,N_5581);
or U8412 (N_8412,N_6871,N_7250);
nor U8413 (N_8413,N_6527,N_5332);
or U8414 (N_8414,N_5276,N_7469);
nor U8415 (N_8415,N_6890,N_5591);
and U8416 (N_8416,N_6269,N_5197);
nor U8417 (N_8417,N_6657,N_5374);
or U8418 (N_8418,N_6785,N_5594);
nand U8419 (N_8419,N_5810,N_6115);
or U8420 (N_8420,N_6634,N_5046);
or U8421 (N_8421,N_5776,N_5506);
or U8422 (N_8422,N_7180,N_5960);
nor U8423 (N_8423,N_5048,N_6731);
nand U8424 (N_8424,N_6268,N_6196);
nor U8425 (N_8425,N_5649,N_6941);
nand U8426 (N_8426,N_5615,N_5272);
and U8427 (N_8427,N_7335,N_5337);
nand U8428 (N_8428,N_5825,N_5939);
nor U8429 (N_8429,N_6915,N_6204);
nand U8430 (N_8430,N_5427,N_6825);
nor U8431 (N_8431,N_6697,N_6958);
and U8432 (N_8432,N_5392,N_5618);
or U8433 (N_8433,N_5449,N_5782);
xor U8434 (N_8434,N_7044,N_6061);
nand U8435 (N_8435,N_5884,N_5007);
and U8436 (N_8436,N_6319,N_7244);
nor U8437 (N_8437,N_5955,N_6625);
and U8438 (N_8438,N_7026,N_7114);
nand U8439 (N_8439,N_6184,N_6505);
nor U8440 (N_8440,N_5001,N_5185);
or U8441 (N_8441,N_6236,N_5735);
and U8442 (N_8442,N_6455,N_6000);
or U8443 (N_8443,N_5330,N_7417);
nor U8444 (N_8444,N_6651,N_5133);
nor U8445 (N_8445,N_5490,N_5841);
xor U8446 (N_8446,N_5834,N_6714);
nor U8447 (N_8447,N_6663,N_5063);
nor U8448 (N_8448,N_6777,N_5273);
or U8449 (N_8449,N_5385,N_6111);
xnor U8450 (N_8450,N_6776,N_5110);
or U8451 (N_8451,N_5372,N_7451);
and U8452 (N_8452,N_6434,N_6594);
nand U8453 (N_8453,N_6161,N_7234);
and U8454 (N_8454,N_7385,N_5970);
and U8455 (N_8455,N_5042,N_6631);
xor U8456 (N_8456,N_6930,N_7317);
or U8457 (N_8457,N_6748,N_7027);
and U8458 (N_8458,N_7347,N_6275);
nor U8459 (N_8459,N_7079,N_5065);
xnor U8460 (N_8460,N_6506,N_6471);
and U8461 (N_8461,N_5681,N_6565);
nand U8462 (N_8462,N_7009,N_6556);
nand U8463 (N_8463,N_5448,N_5015);
nand U8464 (N_8464,N_7163,N_5671);
and U8465 (N_8465,N_6668,N_6822);
and U8466 (N_8466,N_5297,N_6704);
and U8467 (N_8467,N_6146,N_6842);
nor U8468 (N_8468,N_6583,N_5558);
or U8469 (N_8469,N_5285,N_6827);
xnor U8470 (N_8470,N_6836,N_7499);
nand U8471 (N_8471,N_6168,N_6175);
nand U8472 (N_8472,N_5127,N_6109);
or U8473 (N_8473,N_6402,N_7196);
or U8474 (N_8474,N_5807,N_6351);
or U8475 (N_8475,N_6585,N_5429);
or U8476 (N_8476,N_7438,N_6811);
nor U8477 (N_8477,N_7275,N_5953);
or U8478 (N_8478,N_6942,N_5057);
nand U8479 (N_8479,N_6643,N_7445);
and U8480 (N_8480,N_7040,N_6198);
or U8481 (N_8481,N_5699,N_6042);
nor U8482 (N_8482,N_5879,N_5019);
and U8483 (N_8483,N_5093,N_6241);
nor U8484 (N_8484,N_5417,N_5213);
or U8485 (N_8485,N_6340,N_6135);
or U8486 (N_8486,N_5012,N_6163);
or U8487 (N_8487,N_6495,N_6994);
and U8488 (N_8488,N_5460,N_6494);
nor U8489 (N_8489,N_6200,N_6667);
or U8490 (N_8490,N_5308,N_6687);
and U8491 (N_8491,N_6753,N_7303);
or U8492 (N_8492,N_7224,N_5389);
or U8493 (N_8493,N_6737,N_7374);
or U8494 (N_8494,N_6928,N_7437);
nand U8495 (N_8495,N_5471,N_7216);
or U8496 (N_8496,N_6457,N_6313);
nand U8497 (N_8497,N_6213,N_5114);
or U8498 (N_8498,N_6124,N_6536);
xor U8499 (N_8499,N_6133,N_6611);
nor U8500 (N_8500,N_6884,N_6540);
nand U8501 (N_8501,N_5168,N_6231);
or U8502 (N_8502,N_6071,N_5779);
nand U8503 (N_8503,N_7100,N_5310);
or U8504 (N_8504,N_6899,N_7270);
or U8505 (N_8505,N_6214,N_6954);
and U8506 (N_8506,N_5791,N_7404);
or U8507 (N_8507,N_6355,N_5511);
or U8508 (N_8508,N_5672,N_5708);
nand U8509 (N_8509,N_5056,N_5204);
or U8510 (N_8510,N_5729,N_5666);
or U8511 (N_8511,N_5869,N_5384);
or U8512 (N_8512,N_5917,N_5709);
or U8513 (N_8513,N_5640,N_5874);
or U8514 (N_8514,N_6173,N_5570);
and U8515 (N_8515,N_6949,N_5507);
or U8516 (N_8516,N_6129,N_6320);
nand U8517 (N_8517,N_5645,N_7307);
nand U8518 (N_8518,N_5738,N_5987);
or U8519 (N_8519,N_6437,N_6057);
nand U8520 (N_8520,N_6262,N_6308);
and U8521 (N_8521,N_6401,N_5963);
or U8522 (N_8522,N_5112,N_6430);
nor U8523 (N_8523,N_7014,N_6535);
nand U8524 (N_8524,N_7191,N_5433);
or U8525 (N_8525,N_6578,N_6327);
xnor U8526 (N_8526,N_5311,N_5033);
nor U8527 (N_8527,N_7364,N_5367);
nor U8528 (N_8528,N_5706,N_6208);
nand U8529 (N_8529,N_5964,N_6972);
xnor U8530 (N_8530,N_5008,N_6261);
and U8531 (N_8531,N_5271,N_7308);
or U8532 (N_8532,N_7267,N_7116);
nor U8533 (N_8533,N_5827,N_6278);
xnor U8534 (N_8534,N_7113,N_5435);
or U8535 (N_8535,N_6010,N_5892);
nor U8536 (N_8536,N_5317,N_7435);
and U8537 (N_8537,N_6903,N_6851);
and U8538 (N_8538,N_7336,N_5756);
and U8539 (N_8539,N_5670,N_5181);
nor U8540 (N_8540,N_6422,N_5726);
nor U8541 (N_8541,N_5263,N_6803);
nor U8542 (N_8542,N_5413,N_6393);
nor U8543 (N_8543,N_6408,N_5667);
xor U8544 (N_8544,N_5464,N_7042);
nor U8545 (N_8545,N_7342,N_7351);
nand U8546 (N_8546,N_5986,N_7293);
xor U8547 (N_8547,N_5246,N_6377);
nor U8548 (N_8548,N_6654,N_6476);
xnor U8549 (N_8549,N_5351,N_6566);
nand U8550 (N_8550,N_5262,N_7228);
nand U8551 (N_8551,N_7152,N_6014);
nand U8552 (N_8552,N_7072,N_5264);
or U8553 (N_8553,N_5184,N_5222);
nand U8554 (N_8554,N_6946,N_6653);
and U8555 (N_8555,N_5630,N_5498);
nand U8556 (N_8556,N_6452,N_5602);
and U8557 (N_8557,N_7348,N_5898);
and U8558 (N_8558,N_6360,N_6125);
nand U8559 (N_8559,N_6450,N_6296);
nand U8560 (N_8560,N_5387,N_5941);
nor U8561 (N_8561,N_6795,N_5951);
or U8562 (N_8562,N_7379,N_7036);
nor U8563 (N_8563,N_6073,N_7306);
nor U8564 (N_8564,N_6528,N_6496);
nor U8565 (N_8565,N_6177,N_5075);
nand U8566 (N_8566,N_5710,N_5817);
and U8567 (N_8567,N_7010,N_5396);
or U8568 (N_8568,N_6049,N_6085);
and U8569 (N_8569,N_6688,N_7316);
nor U8570 (N_8570,N_6886,N_5965);
and U8571 (N_8571,N_5926,N_6210);
nor U8572 (N_8572,N_7396,N_6660);
or U8573 (N_8573,N_7197,N_5067);
and U8574 (N_8574,N_5294,N_5684);
nand U8575 (N_8575,N_5576,N_7164);
or U8576 (N_8576,N_6224,N_6440);
nor U8577 (N_8577,N_6779,N_7295);
nand U8578 (N_8578,N_7464,N_5544);
or U8579 (N_8579,N_5856,N_5814);
nand U8580 (N_8580,N_5573,N_5325);
nand U8581 (N_8581,N_5677,N_6858);
and U8582 (N_8582,N_5878,N_6745);
xor U8583 (N_8583,N_6227,N_6869);
nand U8584 (N_8584,N_7304,N_5952);
and U8585 (N_8585,N_5073,N_6672);
and U8586 (N_8586,N_6702,N_5156);
and U8587 (N_8587,N_7058,N_5860);
or U8588 (N_8588,N_7327,N_6128);
nor U8589 (N_8589,N_6713,N_7376);
nand U8590 (N_8590,N_5617,N_6966);
and U8591 (N_8591,N_7314,N_5515);
and U8592 (N_8592,N_5479,N_7204);
and U8593 (N_8593,N_5142,N_5697);
nand U8594 (N_8594,N_7021,N_7006);
and U8595 (N_8595,N_5969,N_6628);
nand U8596 (N_8596,N_6099,N_5760);
nand U8597 (N_8597,N_5976,N_6992);
xnor U8598 (N_8598,N_6605,N_6427);
and U8599 (N_8599,N_7496,N_6514);
or U8600 (N_8600,N_5674,N_6025);
and U8601 (N_8601,N_6739,N_5105);
and U8602 (N_8602,N_5804,N_7013);
nor U8603 (N_8603,N_6863,N_7337);
xnor U8604 (N_8604,N_6381,N_7219);
and U8605 (N_8605,N_6303,N_5665);
xor U8606 (N_8606,N_6013,N_7101);
nand U8607 (N_8607,N_7208,N_5176);
nand U8608 (N_8608,N_6079,N_5010);
and U8609 (N_8609,N_7062,N_5556);
nand U8610 (N_8610,N_6741,N_6767);
nand U8611 (N_8611,N_6581,N_6006);
nand U8612 (N_8612,N_6475,N_6245);
and U8613 (N_8613,N_5328,N_7338);
and U8614 (N_8614,N_6248,N_7422);
or U8615 (N_8615,N_6901,N_5265);
nand U8616 (N_8616,N_6235,N_6165);
nor U8617 (N_8617,N_5450,N_5115);
nor U8618 (N_8618,N_6032,N_7212);
nand U8619 (N_8619,N_6768,N_7441);
nand U8620 (N_8620,N_7420,N_7139);
nor U8621 (N_8621,N_5783,N_5946);
or U8622 (N_8622,N_7043,N_6849);
and U8623 (N_8623,N_5359,N_7067);
or U8624 (N_8624,N_5797,N_7497);
nand U8625 (N_8625,N_6326,N_7118);
xnor U8626 (N_8626,N_6993,N_7179);
or U8627 (N_8627,N_6232,N_6730);
or U8628 (N_8628,N_5254,N_7281);
and U8629 (N_8629,N_6624,N_7345);
and U8630 (N_8630,N_6041,N_6088);
or U8631 (N_8631,N_6616,N_5141);
xnor U8632 (N_8632,N_7126,N_7300);
or U8633 (N_8633,N_6542,N_5823);
nand U8634 (N_8634,N_6086,N_5809);
or U8635 (N_8635,N_6104,N_5146);
nor U8636 (N_8636,N_7268,N_6362);
nand U8637 (N_8637,N_5914,N_6973);
xor U8638 (N_8638,N_6960,N_7294);
and U8639 (N_8639,N_5772,N_5949);
nand U8640 (N_8640,N_6837,N_6003);
nand U8641 (N_8641,N_5741,N_5844);
or U8642 (N_8642,N_6885,N_6291);
nand U8643 (N_8643,N_6108,N_5578);
nand U8644 (N_8644,N_6314,N_6067);
nand U8645 (N_8645,N_5373,N_6757);
or U8646 (N_8646,N_7442,N_7470);
or U8647 (N_8647,N_5913,N_5539);
nand U8648 (N_8648,N_6512,N_5867);
or U8649 (N_8649,N_6460,N_5877);
xnor U8650 (N_8650,N_6344,N_5045);
or U8651 (N_8651,N_7102,N_6844);
xor U8652 (N_8652,N_6630,N_6931);
nor U8653 (N_8653,N_7088,N_6920);
or U8654 (N_8654,N_7398,N_5035);
or U8655 (N_8655,N_6429,N_5833);
nor U8656 (N_8656,N_5344,N_7400);
or U8657 (N_8657,N_6134,N_5637);
nand U8658 (N_8658,N_7255,N_6985);
nand U8659 (N_8659,N_6082,N_6772);
nand U8660 (N_8660,N_6019,N_6665);
and U8661 (N_8661,N_5403,N_6490);
xnor U8662 (N_8662,N_6597,N_6036);
or U8663 (N_8663,N_6670,N_6570);
xnor U8664 (N_8664,N_7450,N_5236);
nor U8665 (N_8665,N_6221,N_6357);
nor U8666 (N_8666,N_6407,N_5611);
and U8667 (N_8667,N_7321,N_6603);
nand U8668 (N_8668,N_6783,N_5379);
or U8669 (N_8669,N_6620,N_5178);
nand U8670 (N_8670,N_5907,N_6841);
or U8671 (N_8671,N_5948,N_6185);
xnor U8672 (N_8672,N_7461,N_6707);
nor U8673 (N_8673,N_7193,N_7053);
xor U8674 (N_8674,N_6048,N_6870);
and U8675 (N_8675,N_6220,N_6215);
or U8676 (N_8676,N_6590,N_5501);
or U8677 (N_8677,N_5509,N_5266);
or U8678 (N_8678,N_5426,N_7132);
nor U8679 (N_8679,N_5843,N_6516);
and U8680 (N_8680,N_5248,N_7046);
or U8681 (N_8681,N_7082,N_6549);
xnor U8682 (N_8682,N_6203,N_5394);
nor U8683 (N_8683,N_5446,N_7135);
nor U8684 (N_8684,N_7136,N_7190);
and U8685 (N_8685,N_7096,N_7362);
nor U8686 (N_8686,N_5205,N_6420);
nand U8687 (N_8687,N_6821,N_7075);
and U8688 (N_8688,N_5494,N_7203);
or U8689 (N_8689,N_6755,N_5143);
or U8690 (N_8690,N_5211,N_6459);
nor U8691 (N_8691,N_5757,N_6918);
xor U8692 (N_8692,N_6977,N_6809);
nand U8693 (N_8693,N_6292,N_7276);
xor U8694 (N_8694,N_6055,N_6219);
or U8695 (N_8695,N_6534,N_5944);
and U8696 (N_8696,N_6829,N_5129);
or U8697 (N_8697,N_6254,N_5499);
and U8698 (N_8698,N_7349,N_7060);
nor U8699 (N_8699,N_7285,N_6637);
nor U8700 (N_8700,N_5675,N_7282);
and U8701 (N_8701,N_6028,N_5245);
xor U8702 (N_8702,N_6563,N_6669);
xor U8703 (N_8703,N_6492,N_7246);
or U8704 (N_8704,N_6749,N_7457);
or U8705 (N_8705,N_6020,N_7214);
and U8706 (N_8706,N_7162,N_6072);
nor U8707 (N_8707,N_6760,N_5214);
or U8708 (N_8708,N_5138,N_5549);
nor U8709 (N_8709,N_7448,N_6343);
and U8710 (N_8710,N_5414,N_7183);
and U8711 (N_8711,N_7447,N_6761);
xnor U8712 (N_8712,N_5086,N_5599);
or U8713 (N_8713,N_5320,N_7071);
nand U8714 (N_8714,N_5382,N_5380);
nor U8715 (N_8715,N_5703,N_5496);
nand U8716 (N_8716,N_6859,N_5451);
nand U8717 (N_8717,N_7154,N_7495);
nor U8718 (N_8718,N_5161,N_5559);
and U8719 (N_8719,N_7091,N_5680);
nor U8720 (N_8720,N_6361,N_5842);
or U8721 (N_8721,N_7353,N_6445);
nand U8722 (N_8722,N_5629,N_5119);
and U8723 (N_8723,N_5039,N_5802);
and U8724 (N_8724,N_5688,N_7011);
nor U8725 (N_8725,N_6100,N_6832);
and U8726 (N_8726,N_6069,N_5492);
or U8727 (N_8727,N_6686,N_5111);
xor U8728 (N_8728,N_6696,N_7458);
nor U8729 (N_8729,N_7427,N_7296);
xor U8730 (N_8730,N_6169,N_7352);
nand U8731 (N_8731,N_7280,N_6622);
xor U8732 (N_8732,N_6462,N_5808);
nor U8733 (N_8733,N_6035,N_6951);
and U8734 (N_8734,N_6586,N_6312);
nor U8735 (N_8735,N_5815,N_6830);
nor U8736 (N_8736,N_7394,N_5312);
or U8737 (N_8737,N_6914,N_5341);
nor U8738 (N_8738,N_6229,N_6626);
or U8739 (N_8739,N_5719,N_6187);
nand U8740 (N_8740,N_5171,N_5125);
or U8741 (N_8741,N_6880,N_5153);
nor U8742 (N_8742,N_5469,N_5536);
and U8743 (N_8743,N_5534,N_7153);
xnor U8744 (N_8744,N_7313,N_5628);
or U8745 (N_8745,N_6295,N_6968);
nor U8746 (N_8746,N_5179,N_6769);
nand U8747 (N_8747,N_6499,N_6732);
or U8748 (N_8748,N_6149,N_6893);
nand U8749 (N_8749,N_5049,N_6216);
nor U8750 (N_8750,N_6472,N_7184);
nor U8751 (N_8751,N_6866,N_6065);
xnor U8752 (N_8752,N_7231,N_6684);
and U8753 (N_8753,N_6666,N_7388);
and U8754 (N_8754,N_6605,N_5734);
nand U8755 (N_8755,N_5345,N_6131);
or U8756 (N_8756,N_6934,N_5797);
nand U8757 (N_8757,N_6480,N_6434);
nor U8758 (N_8758,N_5488,N_6626);
or U8759 (N_8759,N_5595,N_5490);
or U8760 (N_8760,N_5149,N_7182);
nor U8761 (N_8761,N_6720,N_6628);
or U8762 (N_8762,N_7217,N_5908);
nand U8763 (N_8763,N_6079,N_5204);
nand U8764 (N_8764,N_7376,N_6311);
xnor U8765 (N_8765,N_5422,N_5687);
or U8766 (N_8766,N_5781,N_7176);
or U8767 (N_8767,N_7285,N_5254);
nand U8768 (N_8768,N_6836,N_6252);
and U8769 (N_8769,N_7263,N_5816);
or U8770 (N_8770,N_6509,N_6610);
xnor U8771 (N_8771,N_7383,N_7355);
and U8772 (N_8772,N_6797,N_7312);
or U8773 (N_8773,N_7055,N_7171);
or U8774 (N_8774,N_6213,N_5679);
xnor U8775 (N_8775,N_6473,N_6744);
and U8776 (N_8776,N_6141,N_6788);
nor U8777 (N_8777,N_5097,N_5383);
nand U8778 (N_8778,N_6011,N_6737);
nor U8779 (N_8779,N_6560,N_5670);
and U8780 (N_8780,N_6178,N_6626);
nand U8781 (N_8781,N_6399,N_5467);
xor U8782 (N_8782,N_6151,N_7215);
nor U8783 (N_8783,N_6554,N_6138);
nor U8784 (N_8784,N_6180,N_7094);
nor U8785 (N_8785,N_6307,N_5895);
nand U8786 (N_8786,N_6272,N_5690);
and U8787 (N_8787,N_5516,N_7407);
nand U8788 (N_8788,N_5646,N_7456);
nand U8789 (N_8789,N_7021,N_5215);
and U8790 (N_8790,N_6501,N_5824);
nand U8791 (N_8791,N_6886,N_6379);
or U8792 (N_8792,N_6002,N_5378);
nor U8793 (N_8793,N_5285,N_5465);
and U8794 (N_8794,N_7077,N_6627);
nor U8795 (N_8795,N_7423,N_6228);
or U8796 (N_8796,N_5570,N_7050);
or U8797 (N_8797,N_6919,N_5750);
nor U8798 (N_8798,N_6774,N_6848);
and U8799 (N_8799,N_7037,N_6406);
nor U8800 (N_8800,N_6925,N_6589);
or U8801 (N_8801,N_6777,N_6457);
or U8802 (N_8802,N_6956,N_7166);
nor U8803 (N_8803,N_6757,N_5709);
nor U8804 (N_8804,N_6572,N_5895);
nor U8805 (N_8805,N_7215,N_6599);
and U8806 (N_8806,N_6299,N_5861);
or U8807 (N_8807,N_5837,N_5723);
and U8808 (N_8808,N_7311,N_7257);
or U8809 (N_8809,N_6032,N_5949);
nand U8810 (N_8810,N_5836,N_5658);
nand U8811 (N_8811,N_5623,N_7440);
and U8812 (N_8812,N_5553,N_5944);
xor U8813 (N_8813,N_6825,N_6098);
or U8814 (N_8814,N_6632,N_6056);
or U8815 (N_8815,N_6022,N_5749);
or U8816 (N_8816,N_5296,N_6632);
nor U8817 (N_8817,N_5877,N_6273);
or U8818 (N_8818,N_7471,N_6157);
or U8819 (N_8819,N_5955,N_7467);
nor U8820 (N_8820,N_5026,N_6431);
or U8821 (N_8821,N_6893,N_5286);
xor U8822 (N_8822,N_5770,N_5051);
nand U8823 (N_8823,N_5695,N_7288);
or U8824 (N_8824,N_6559,N_6056);
or U8825 (N_8825,N_6234,N_5212);
and U8826 (N_8826,N_6320,N_6419);
or U8827 (N_8827,N_5865,N_7103);
nor U8828 (N_8828,N_5657,N_5017);
nand U8829 (N_8829,N_6610,N_5287);
or U8830 (N_8830,N_5401,N_7393);
nand U8831 (N_8831,N_6199,N_7317);
nand U8832 (N_8832,N_5182,N_7153);
nand U8833 (N_8833,N_6041,N_7055);
nand U8834 (N_8834,N_5212,N_5793);
nor U8835 (N_8835,N_5131,N_6841);
nor U8836 (N_8836,N_6578,N_7327);
or U8837 (N_8837,N_5525,N_7309);
nor U8838 (N_8838,N_5643,N_7294);
or U8839 (N_8839,N_6400,N_5906);
or U8840 (N_8840,N_7043,N_5038);
nand U8841 (N_8841,N_7067,N_6128);
or U8842 (N_8842,N_5656,N_6768);
xor U8843 (N_8843,N_6760,N_5067);
nor U8844 (N_8844,N_5047,N_5258);
xnor U8845 (N_8845,N_6378,N_7271);
xnor U8846 (N_8846,N_5522,N_6960);
and U8847 (N_8847,N_5714,N_7133);
or U8848 (N_8848,N_6988,N_6093);
and U8849 (N_8849,N_6980,N_6794);
nor U8850 (N_8850,N_5973,N_5531);
nor U8851 (N_8851,N_7112,N_6644);
and U8852 (N_8852,N_7111,N_5120);
and U8853 (N_8853,N_6468,N_7090);
xor U8854 (N_8854,N_7294,N_5278);
or U8855 (N_8855,N_5969,N_6303);
or U8856 (N_8856,N_5171,N_5540);
or U8857 (N_8857,N_6566,N_6726);
nor U8858 (N_8858,N_7409,N_5202);
and U8859 (N_8859,N_5325,N_6432);
or U8860 (N_8860,N_5094,N_6403);
nand U8861 (N_8861,N_7086,N_5892);
nand U8862 (N_8862,N_5066,N_6440);
nand U8863 (N_8863,N_5951,N_7366);
or U8864 (N_8864,N_5750,N_7330);
nand U8865 (N_8865,N_5699,N_7199);
nand U8866 (N_8866,N_6893,N_5722);
and U8867 (N_8867,N_7466,N_5511);
or U8868 (N_8868,N_5485,N_6078);
nand U8869 (N_8869,N_5330,N_7245);
and U8870 (N_8870,N_5641,N_7293);
nand U8871 (N_8871,N_6551,N_7180);
and U8872 (N_8872,N_6166,N_5377);
and U8873 (N_8873,N_5212,N_5944);
nand U8874 (N_8874,N_6908,N_5775);
or U8875 (N_8875,N_5421,N_5128);
or U8876 (N_8876,N_6978,N_5710);
and U8877 (N_8877,N_5822,N_5094);
nand U8878 (N_8878,N_7323,N_5400);
nor U8879 (N_8879,N_5761,N_5053);
or U8880 (N_8880,N_6590,N_6171);
or U8881 (N_8881,N_5831,N_5301);
nand U8882 (N_8882,N_6243,N_5306);
and U8883 (N_8883,N_6132,N_5728);
nand U8884 (N_8884,N_5321,N_5204);
or U8885 (N_8885,N_5135,N_7450);
nand U8886 (N_8886,N_7139,N_5055);
or U8887 (N_8887,N_5713,N_7299);
or U8888 (N_8888,N_6809,N_7123);
and U8889 (N_8889,N_7293,N_5342);
and U8890 (N_8890,N_5630,N_7310);
nand U8891 (N_8891,N_6101,N_6173);
and U8892 (N_8892,N_5777,N_6920);
or U8893 (N_8893,N_6600,N_7135);
nor U8894 (N_8894,N_6682,N_6187);
nor U8895 (N_8895,N_5865,N_6126);
nand U8896 (N_8896,N_7197,N_6727);
nand U8897 (N_8897,N_5540,N_6972);
nand U8898 (N_8898,N_6500,N_6089);
nor U8899 (N_8899,N_5744,N_5292);
or U8900 (N_8900,N_5444,N_5731);
nand U8901 (N_8901,N_6878,N_5303);
or U8902 (N_8902,N_7042,N_5758);
or U8903 (N_8903,N_7373,N_5855);
nand U8904 (N_8904,N_7472,N_5000);
nand U8905 (N_8905,N_5520,N_6734);
nor U8906 (N_8906,N_7282,N_6313);
nand U8907 (N_8907,N_5510,N_7010);
and U8908 (N_8908,N_6226,N_5363);
or U8909 (N_8909,N_6740,N_5984);
nand U8910 (N_8910,N_5590,N_6478);
and U8911 (N_8911,N_7367,N_6914);
and U8912 (N_8912,N_5058,N_5599);
or U8913 (N_8913,N_5184,N_5611);
and U8914 (N_8914,N_5549,N_7273);
nor U8915 (N_8915,N_5158,N_7220);
and U8916 (N_8916,N_5927,N_6639);
nor U8917 (N_8917,N_5022,N_7207);
or U8918 (N_8918,N_7486,N_5746);
or U8919 (N_8919,N_5449,N_5026);
nor U8920 (N_8920,N_7393,N_6193);
and U8921 (N_8921,N_5097,N_6676);
and U8922 (N_8922,N_7397,N_5264);
xor U8923 (N_8923,N_6083,N_5481);
xor U8924 (N_8924,N_5173,N_5181);
and U8925 (N_8925,N_6088,N_5600);
nor U8926 (N_8926,N_5840,N_5224);
xnor U8927 (N_8927,N_5272,N_5831);
nand U8928 (N_8928,N_6377,N_5182);
nor U8929 (N_8929,N_6691,N_5717);
and U8930 (N_8930,N_5850,N_5692);
or U8931 (N_8931,N_5341,N_7285);
nor U8932 (N_8932,N_7187,N_5045);
or U8933 (N_8933,N_5746,N_7342);
or U8934 (N_8934,N_5659,N_5618);
xor U8935 (N_8935,N_7273,N_7301);
nand U8936 (N_8936,N_6165,N_5993);
and U8937 (N_8937,N_6984,N_6197);
nand U8938 (N_8938,N_5576,N_6443);
and U8939 (N_8939,N_7426,N_7135);
and U8940 (N_8940,N_5329,N_6797);
nand U8941 (N_8941,N_6780,N_5518);
nand U8942 (N_8942,N_6505,N_5367);
nor U8943 (N_8943,N_6032,N_7263);
or U8944 (N_8944,N_6685,N_7412);
and U8945 (N_8945,N_7123,N_7296);
or U8946 (N_8946,N_6769,N_5197);
xnor U8947 (N_8947,N_7490,N_6829);
or U8948 (N_8948,N_6080,N_7300);
nand U8949 (N_8949,N_5749,N_5649);
nand U8950 (N_8950,N_6839,N_5369);
nand U8951 (N_8951,N_7222,N_6963);
nor U8952 (N_8952,N_6679,N_7232);
and U8953 (N_8953,N_6406,N_6464);
nor U8954 (N_8954,N_5779,N_6815);
nor U8955 (N_8955,N_5429,N_7293);
or U8956 (N_8956,N_5417,N_6100);
and U8957 (N_8957,N_5156,N_6554);
nand U8958 (N_8958,N_5012,N_6834);
or U8959 (N_8959,N_5830,N_7430);
nor U8960 (N_8960,N_7399,N_6351);
and U8961 (N_8961,N_6309,N_6055);
or U8962 (N_8962,N_7196,N_5763);
or U8963 (N_8963,N_6791,N_6721);
and U8964 (N_8964,N_6247,N_6187);
and U8965 (N_8965,N_5863,N_6435);
xnor U8966 (N_8966,N_6745,N_6318);
xnor U8967 (N_8967,N_5542,N_7019);
nand U8968 (N_8968,N_5206,N_6497);
xnor U8969 (N_8969,N_6171,N_5698);
xnor U8970 (N_8970,N_6702,N_7257);
or U8971 (N_8971,N_7102,N_5084);
and U8972 (N_8972,N_7397,N_5724);
nor U8973 (N_8973,N_6988,N_6030);
xnor U8974 (N_8974,N_5905,N_5925);
and U8975 (N_8975,N_6278,N_6244);
nand U8976 (N_8976,N_5301,N_6925);
or U8977 (N_8977,N_5999,N_5204);
nand U8978 (N_8978,N_6300,N_6804);
xnor U8979 (N_8979,N_7177,N_5525);
and U8980 (N_8980,N_5128,N_6923);
and U8981 (N_8981,N_5481,N_5764);
nand U8982 (N_8982,N_7415,N_6073);
xor U8983 (N_8983,N_5673,N_5769);
nand U8984 (N_8984,N_5075,N_7267);
nor U8985 (N_8985,N_7335,N_5210);
and U8986 (N_8986,N_6776,N_6939);
xnor U8987 (N_8987,N_6538,N_7137);
and U8988 (N_8988,N_5784,N_6170);
nand U8989 (N_8989,N_6315,N_5471);
or U8990 (N_8990,N_7241,N_6687);
or U8991 (N_8991,N_6266,N_5242);
and U8992 (N_8992,N_6223,N_7444);
nor U8993 (N_8993,N_5686,N_6724);
xor U8994 (N_8994,N_6315,N_6198);
nor U8995 (N_8995,N_5447,N_7440);
nand U8996 (N_8996,N_5207,N_5610);
and U8997 (N_8997,N_5396,N_5411);
and U8998 (N_8998,N_6914,N_7314);
or U8999 (N_8999,N_5899,N_5631);
nand U9000 (N_9000,N_5083,N_6517);
nor U9001 (N_9001,N_5388,N_6376);
xnor U9002 (N_9002,N_6098,N_6478);
nand U9003 (N_9003,N_5232,N_5872);
nand U9004 (N_9004,N_6634,N_6912);
nor U9005 (N_9005,N_6877,N_7296);
nor U9006 (N_9006,N_5141,N_7372);
nor U9007 (N_9007,N_7476,N_6636);
or U9008 (N_9008,N_6951,N_6401);
xnor U9009 (N_9009,N_6007,N_6582);
xnor U9010 (N_9010,N_5129,N_6525);
nand U9011 (N_9011,N_5987,N_7323);
or U9012 (N_9012,N_6348,N_6734);
xor U9013 (N_9013,N_5622,N_6085);
nand U9014 (N_9014,N_6253,N_7129);
or U9015 (N_9015,N_5467,N_6059);
and U9016 (N_9016,N_5212,N_6257);
xor U9017 (N_9017,N_6062,N_5982);
nor U9018 (N_9018,N_6938,N_7075);
nand U9019 (N_9019,N_7494,N_6407);
and U9020 (N_9020,N_6577,N_6068);
nor U9021 (N_9021,N_7327,N_7278);
xnor U9022 (N_9022,N_6361,N_5875);
nand U9023 (N_9023,N_6369,N_7023);
nor U9024 (N_9024,N_6754,N_5879);
nand U9025 (N_9025,N_7397,N_5491);
nand U9026 (N_9026,N_5849,N_7449);
xnor U9027 (N_9027,N_5955,N_6739);
nand U9028 (N_9028,N_7065,N_6154);
nor U9029 (N_9029,N_7100,N_6556);
nand U9030 (N_9030,N_5353,N_5292);
and U9031 (N_9031,N_6551,N_5739);
and U9032 (N_9032,N_6628,N_5106);
nand U9033 (N_9033,N_7038,N_5186);
nor U9034 (N_9034,N_5287,N_5409);
xor U9035 (N_9035,N_5347,N_6929);
nand U9036 (N_9036,N_6125,N_7495);
xnor U9037 (N_9037,N_5180,N_5509);
or U9038 (N_9038,N_5361,N_5625);
xnor U9039 (N_9039,N_5371,N_6700);
xor U9040 (N_9040,N_5084,N_7428);
or U9041 (N_9041,N_7344,N_5286);
or U9042 (N_9042,N_5543,N_5335);
and U9043 (N_9043,N_5726,N_7038);
nand U9044 (N_9044,N_7451,N_6997);
nand U9045 (N_9045,N_5711,N_6598);
or U9046 (N_9046,N_6277,N_6292);
and U9047 (N_9047,N_6000,N_5675);
and U9048 (N_9048,N_6735,N_7111);
nor U9049 (N_9049,N_5665,N_5785);
nand U9050 (N_9050,N_7301,N_6258);
and U9051 (N_9051,N_6617,N_5997);
and U9052 (N_9052,N_6184,N_6846);
nor U9053 (N_9053,N_5394,N_6838);
and U9054 (N_9054,N_5832,N_5213);
nor U9055 (N_9055,N_5294,N_6120);
nor U9056 (N_9056,N_7362,N_5832);
or U9057 (N_9057,N_6391,N_6169);
or U9058 (N_9058,N_6717,N_6593);
nand U9059 (N_9059,N_7094,N_6594);
nand U9060 (N_9060,N_5779,N_6784);
and U9061 (N_9061,N_6717,N_5218);
or U9062 (N_9062,N_6303,N_5077);
or U9063 (N_9063,N_6631,N_5564);
nand U9064 (N_9064,N_5486,N_7047);
nor U9065 (N_9065,N_6388,N_6131);
nor U9066 (N_9066,N_6826,N_5077);
or U9067 (N_9067,N_6139,N_7177);
and U9068 (N_9068,N_5112,N_6882);
nor U9069 (N_9069,N_5910,N_5968);
nand U9070 (N_9070,N_6472,N_7109);
or U9071 (N_9071,N_5591,N_5997);
and U9072 (N_9072,N_6683,N_5399);
and U9073 (N_9073,N_7226,N_6456);
xnor U9074 (N_9074,N_6942,N_6604);
or U9075 (N_9075,N_6577,N_6833);
nor U9076 (N_9076,N_5561,N_6615);
nand U9077 (N_9077,N_6139,N_6485);
nor U9078 (N_9078,N_5744,N_6168);
and U9079 (N_9079,N_5658,N_6903);
nand U9080 (N_9080,N_5106,N_6456);
and U9081 (N_9081,N_5180,N_5029);
and U9082 (N_9082,N_6132,N_5760);
nand U9083 (N_9083,N_5134,N_5149);
nor U9084 (N_9084,N_5249,N_7482);
nor U9085 (N_9085,N_5897,N_7116);
or U9086 (N_9086,N_7271,N_5205);
nand U9087 (N_9087,N_6470,N_5215);
or U9088 (N_9088,N_5578,N_7397);
or U9089 (N_9089,N_5441,N_5328);
nand U9090 (N_9090,N_5909,N_6885);
or U9091 (N_9091,N_6042,N_5721);
nand U9092 (N_9092,N_6647,N_6503);
nand U9093 (N_9093,N_7356,N_6958);
nand U9094 (N_9094,N_7062,N_5841);
nor U9095 (N_9095,N_7401,N_5316);
and U9096 (N_9096,N_5482,N_5218);
xor U9097 (N_9097,N_6312,N_6474);
or U9098 (N_9098,N_5475,N_6608);
nor U9099 (N_9099,N_6887,N_6872);
or U9100 (N_9100,N_6710,N_5192);
and U9101 (N_9101,N_6085,N_6951);
or U9102 (N_9102,N_7021,N_7467);
and U9103 (N_9103,N_7374,N_5118);
or U9104 (N_9104,N_6557,N_6524);
nor U9105 (N_9105,N_5022,N_6000);
and U9106 (N_9106,N_5430,N_5727);
and U9107 (N_9107,N_7169,N_5500);
and U9108 (N_9108,N_7241,N_5043);
or U9109 (N_9109,N_5903,N_6961);
nor U9110 (N_9110,N_7432,N_7458);
nand U9111 (N_9111,N_6406,N_7099);
or U9112 (N_9112,N_5130,N_7016);
or U9113 (N_9113,N_6072,N_7314);
or U9114 (N_9114,N_7457,N_5660);
or U9115 (N_9115,N_5021,N_7151);
nor U9116 (N_9116,N_5199,N_6833);
nand U9117 (N_9117,N_7235,N_5691);
or U9118 (N_9118,N_6557,N_7086);
and U9119 (N_9119,N_6403,N_6183);
nand U9120 (N_9120,N_6548,N_5443);
nand U9121 (N_9121,N_7346,N_7421);
and U9122 (N_9122,N_5716,N_5643);
or U9123 (N_9123,N_7404,N_6970);
and U9124 (N_9124,N_5872,N_6076);
nor U9125 (N_9125,N_7010,N_5053);
nor U9126 (N_9126,N_6538,N_5180);
or U9127 (N_9127,N_5422,N_7321);
nor U9128 (N_9128,N_5734,N_6344);
or U9129 (N_9129,N_6549,N_6593);
xor U9130 (N_9130,N_5541,N_5141);
xnor U9131 (N_9131,N_5914,N_5763);
or U9132 (N_9132,N_5496,N_5304);
nand U9133 (N_9133,N_7109,N_5071);
nand U9134 (N_9134,N_5534,N_5987);
nand U9135 (N_9135,N_6482,N_5844);
or U9136 (N_9136,N_7309,N_6236);
nor U9137 (N_9137,N_6650,N_6217);
or U9138 (N_9138,N_6888,N_6260);
nand U9139 (N_9139,N_6710,N_6239);
xnor U9140 (N_9140,N_6740,N_7334);
or U9141 (N_9141,N_5293,N_7443);
nor U9142 (N_9142,N_6098,N_7198);
and U9143 (N_9143,N_6136,N_6503);
and U9144 (N_9144,N_5730,N_7119);
nand U9145 (N_9145,N_5433,N_6610);
nand U9146 (N_9146,N_7118,N_5821);
nor U9147 (N_9147,N_6309,N_6297);
nand U9148 (N_9148,N_6737,N_5964);
nor U9149 (N_9149,N_6926,N_7273);
nor U9150 (N_9150,N_6486,N_6417);
nand U9151 (N_9151,N_6504,N_5288);
or U9152 (N_9152,N_6014,N_6458);
nor U9153 (N_9153,N_5980,N_6686);
or U9154 (N_9154,N_5153,N_5975);
nand U9155 (N_9155,N_6888,N_6886);
and U9156 (N_9156,N_6044,N_5620);
or U9157 (N_9157,N_6526,N_5253);
nor U9158 (N_9158,N_6226,N_6176);
nor U9159 (N_9159,N_7094,N_7314);
nor U9160 (N_9160,N_7007,N_5661);
or U9161 (N_9161,N_7043,N_5132);
xnor U9162 (N_9162,N_5533,N_6654);
or U9163 (N_9163,N_6535,N_5909);
xor U9164 (N_9164,N_7308,N_7021);
nor U9165 (N_9165,N_7396,N_6458);
and U9166 (N_9166,N_6967,N_5108);
and U9167 (N_9167,N_7169,N_5478);
nor U9168 (N_9168,N_5364,N_6132);
and U9169 (N_9169,N_5633,N_6977);
nand U9170 (N_9170,N_5831,N_5392);
or U9171 (N_9171,N_5194,N_6503);
or U9172 (N_9172,N_6721,N_6360);
nor U9173 (N_9173,N_5139,N_6408);
and U9174 (N_9174,N_6428,N_5959);
and U9175 (N_9175,N_5347,N_6833);
xnor U9176 (N_9176,N_6877,N_5008);
nor U9177 (N_9177,N_5917,N_5098);
and U9178 (N_9178,N_6586,N_6398);
nand U9179 (N_9179,N_6962,N_5499);
nand U9180 (N_9180,N_6719,N_6334);
and U9181 (N_9181,N_7467,N_6285);
nor U9182 (N_9182,N_6655,N_5986);
or U9183 (N_9183,N_5731,N_5083);
and U9184 (N_9184,N_6323,N_6750);
and U9185 (N_9185,N_6319,N_5322);
and U9186 (N_9186,N_6106,N_5593);
nand U9187 (N_9187,N_7310,N_6773);
xor U9188 (N_9188,N_5569,N_6122);
or U9189 (N_9189,N_6444,N_7172);
nor U9190 (N_9190,N_6151,N_5253);
and U9191 (N_9191,N_6982,N_5210);
and U9192 (N_9192,N_5043,N_5502);
and U9193 (N_9193,N_6529,N_5569);
or U9194 (N_9194,N_5085,N_5353);
nor U9195 (N_9195,N_5671,N_7079);
xnor U9196 (N_9196,N_6714,N_6793);
and U9197 (N_9197,N_6684,N_6929);
nor U9198 (N_9198,N_6697,N_6365);
nor U9199 (N_9199,N_6242,N_5685);
nand U9200 (N_9200,N_5931,N_6614);
nand U9201 (N_9201,N_5973,N_6066);
and U9202 (N_9202,N_6163,N_6225);
or U9203 (N_9203,N_5443,N_5873);
or U9204 (N_9204,N_7399,N_6828);
and U9205 (N_9205,N_7062,N_5041);
nor U9206 (N_9206,N_5948,N_7078);
nor U9207 (N_9207,N_7178,N_7204);
and U9208 (N_9208,N_7327,N_5679);
or U9209 (N_9209,N_6941,N_7237);
xnor U9210 (N_9210,N_6457,N_7498);
nand U9211 (N_9211,N_6582,N_5749);
xnor U9212 (N_9212,N_5706,N_6329);
nand U9213 (N_9213,N_6908,N_7480);
nor U9214 (N_9214,N_5235,N_6207);
nor U9215 (N_9215,N_5289,N_7408);
nand U9216 (N_9216,N_5088,N_6398);
or U9217 (N_9217,N_7258,N_5984);
nand U9218 (N_9218,N_6909,N_7188);
or U9219 (N_9219,N_5767,N_7123);
nor U9220 (N_9220,N_5798,N_5846);
nand U9221 (N_9221,N_6629,N_6952);
and U9222 (N_9222,N_6527,N_6524);
nor U9223 (N_9223,N_5273,N_5654);
nand U9224 (N_9224,N_5258,N_6901);
nand U9225 (N_9225,N_6678,N_5337);
nor U9226 (N_9226,N_6523,N_5401);
nor U9227 (N_9227,N_6599,N_6569);
and U9228 (N_9228,N_6883,N_6416);
nor U9229 (N_9229,N_5136,N_6835);
xor U9230 (N_9230,N_7393,N_5042);
or U9231 (N_9231,N_5429,N_6546);
nand U9232 (N_9232,N_5172,N_7098);
nand U9233 (N_9233,N_6837,N_5163);
and U9234 (N_9234,N_5731,N_7280);
nand U9235 (N_9235,N_5046,N_6160);
nand U9236 (N_9236,N_6653,N_5609);
or U9237 (N_9237,N_6331,N_5385);
and U9238 (N_9238,N_6059,N_7017);
nand U9239 (N_9239,N_7089,N_5890);
nor U9240 (N_9240,N_7342,N_6417);
nand U9241 (N_9241,N_5451,N_5583);
and U9242 (N_9242,N_5835,N_6575);
and U9243 (N_9243,N_7339,N_5040);
or U9244 (N_9244,N_6898,N_6793);
and U9245 (N_9245,N_5838,N_6056);
or U9246 (N_9246,N_5559,N_6894);
and U9247 (N_9247,N_5223,N_7275);
or U9248 (N_9248,N_5790,N_5771);
and U9249 (N_9249,N_6788,N_6346);
nor U9250 (N_9250,N_5354,N_6598);
or U9251 (N_9251,N_6268,N_5568);
or U9252 (N_9252,N_7154,N_6416);
and U9253 (N_9253,N_6071,N_6825);
nand U9254 (N_9254,N_5118,N_7413);
or U9255 (N_9255,N_5326,N_7277);
and U9256 (N_9256,N_6473,N_7393);
nor U9257 (N_9257,N_7344,N_6221);
nor U9258 (N_9258,N_5633,N_5629);
xnor U9259 (N_9259,N_6355,N_5049);
xnor U9260 (N_9260,N_7021,N_7480);
and U9261 (N_9261,N_7109,N_5672);
and U9262 (N_9262,N_6670,N_7241);
or U9263 (N_9263,N_6152,N_5727);
nor U9264 (N_9264,N_6279,N_5133);
and U9265 (N_9265,N_6058,N_6620);
nand U9266 (N_9266,N_6038,N_6165);
or U9267 (N_9267,N_7464,N_6255);
xor U9268 (N_9268,N_6262,N_6844);
or U9269 (N_9269,N_7055,N_5192);
and U9270 (N_9270,N_5863,N_7220);
or U9271 (N_9271,N_6117,N_5316);
nor U9272 (N_9272,N_6724,N_5230);
or U9273 (N_9273,N_6987,N_5988);
nor U9274 (N_9274,N_5610,N_6400);
and U9275 (N_9275,N_6969,N_5358);
nand U9276 (N_9276,N_5991,N_6498);
and U9277 (N_9277,N_5495,N_5914);
nor U9278 (N_9278,N_5680,N_5016);
or U9279 (N_9279,N_5716,N_6430);
nor U9280 (N_9280,N_6581,N_6854);
and U9281 (N_9281,N_7457,N_5934);
xnor U9282 (N_9282,N_5630,N_7334);
nand U9283 (N_9283,N_6183,N_6915);
nand U9284 (N_9284,N_6811,N_7071);
nand U9285 (N_9285,N_6764,N_6053);
or U9286 (N_9286,N_6905,N_7176);
nor U9287 (N_9287,N_5639,N_7383);
nand U9288 (N_9288,N_7075,N_6918);
and U9289 (N_9289,N_6543,N_5317);
or U9290 (N_9290,N_6782,N_6815);
nand U9291 (N_9291,N_5592,N_6848);
and U9292 (N_9292,N_6131,N_5833);
and U9293 (N_9293,N_6973,N_5054);
or U9294 (N_9294,N_7333,N_5254);
and U9295 (N_9295,N_5812,N_5716);
or U9296 (N_9296,N_6738,N_6284);
xor U9297 (N_9297,N_5055,N_6988);
or U9298 (N_9298,N_5715,N_5770);
and U9299 (N_9299,N_5603,N_7365);
nand U9300 (N_9300,N_6630,N_6362);
nor U9301 (N_9301,N_5523,N_7253);
nand U9302 (N_9302,N_5326,N_5684);
nand U9303 (N_9303,N_6756,N_6878);
nand U9304 (N_9304,N_5098,N_6426);
or U9305 (N_9305,N_6221,N_7200);
nor U9306 (N_9306,N_5949,N_5765);
nand U9307 (N_9307,N_7474,N_6543);
nor U9308 (N_9308,N_5771,N_5157);
or U9309 (N_9309,N_7176,N_7198);
nor U9310 (N_9310,N_7246,N_5958);
nor U9311 (N_9311,N_5121,N_7026);
nand U9312 (N_9312,N_5912,N_5366);
nand U9313 (N_9313,N_6563,N_6966);
and U9314 (N_9314,N_5987,N_6424);
and U9315 (N_9315,N_5350,N_6990);
nand U9316 (N_9316,N_6142,N_5331);
xnor U9317 (N_9317,N_7406,N_6799);
nand U9318 (N_9318,N_5246,N_5746);
and U9319 (N_9319,N_6228,N_5813);
or U9320 (N_9320,N_7227,N_5205);
or U9321 (N_9321,N_7332,N_6580);
nor U9322 (N_9322,N_5855,N_5131);
nand U9323 (N_9323,N_5177,N_7031);
nand U9324 (N_9324,N_5757,N_6912);
and U9325 (N_9325,N_7360,N_5595);
nand U9326 (N_9326,N_7154,N_5985);
nand U9327 (N_9327,N_6130,N_6019);
xnor U9328 (N_9328,N_6072,N_6425);
xor U9329 (N_9329,N_7382,N_6308);
and U9330 (N_9330,N_5570,N_5308);
xnor U9331 (N_9331,N_7325,N_5016);
or U9332 (N_9332,N_6325,N_5308);
and U9333 (N_9333,N_5670,N_6435);
and U9334 (N_9334,N_6939,N_7328);
nand U9335 (N_9335,N_6520,N_5880);
and U9336 (N_9336,N_7224,N_5769);
and U9337 (N_9337,N_5192,N_7171);
nor U9338 (N_9338,N_5700,N_6061);
nand U9339 (N_9339,N_6667,N_7386);
xor U9340 (N_9340,N_5589,N_5114);
nand U9341 (N_9341,N_7138,N_7022);
nor U9342 (N_9342,N_7061,N_7485);
and U9343 (N_9343,N_7400,N_5382);
nor U9344 (N_9344,N_5913,N_5003);
nand U9345 (N_9345,N_5240,N_6558);
and U9346 (N_9346,N_7043,N_5208);
nand U9347 (N_9347,N_5765,N_7067);
and U9348 (N_9348,N_6815,N_7032);
nand U9349 (N_9349,N_5181,N_5830);
or U9350 (N_9350,N_5566,N_5138);
xor U9351 (N_9351,N_5216,N_7130);
nor U9352 (N_9352,N_5082,N_6483);
and U9353 (N_9353,N_6887,N_5440);
nand U9354 (N_9354,N_5085,N_5980);
nand U9355 (N_9355,N_5178,N_6466);
nor U9356 (N_9356,N_5093,N_6692);
and U9357 (N_9357,N_6283,N_7217);
and U9358 (N_9358,N_6855,N_6731);
or U9359 (N_9359,N_5398,N_6415);
or U9360 (N_9360,N_5895,N_7183);
nand U9361 (N_9361,N_7171,N_5647);
nand U9362 (N_9362,N_5036,N_7386);
and U9363 (N_9363,N_6912,N_7036);
nand U9364 (N_9364,N_7002,N_5193);
and U9365 (N_9365,N_6708,N_7269);
nor U9366 (N_9366,N_5715,N_6515);
and U9367 (N_9367,N_7449,N_6741);
nor U9368 (N_9368,N_5756,N_5866);
xor U9369 (N_9369,N_6039,N_7410);
and U9370 (N_9370,N_6215,N_5058);
or U9371 (N_9371,N_6085,N_6375);
nand U9372 (N_9372,N_7200,N_6306);
nand U9373 (N_9373,N_7093,N_5492);
xnor U9374 (N_9374,N_7049,N_5281);
xor U9375 (N_9375,N_5811,N_5933);
or U9376 (N_9376,N_5579,N_5087);
or U9377 (N_9377,N_6724,N_6541);
or U9378 (N_9378,N_6884,N_5997);
nand U9379 (N_9379,N_5066,N_7302);
xnor U9380 (N_9380,N_5158,N_5953);
nand U9381 (N_9381,N_5517,N_5320);
nor U9382 (N_9382,N_5410,N_5312);
and U9383 (N_9383,N_6537,N_7081);
nand U9384 (N_9384,N_6415,N_6885);
or U9385 (N_9385,N_6713,N_5181);
xor U9386 (N_9386,N_6494,N_5217);
and U9387 (N_9387,N_5457,N_7311);
nand U9388 (N_9388,N_5441,N_5476);
and U9389 (N_9389,N_5503,N_6769);
xor U9390 (N_9390,N_5909,N_6373);
or U9391 (N_9391,N_6882,N_7114);
and U9392 (N_9392,N_6637,N_5553);
and U9393 (N_9393,N_6162,N_6485);
or U9394 (N_9394,N_7211,N_5086);
or U9395 (N_9395,N_5195,N_6405);
and U9396 (N_9396,N_6870,N_6291);
nor U9397 (N_9397,N_5370,N_6312);
and U9398 (N_9398,N_6330,N_6017);
and U9399 (N_9399,N_6706,N_5870);
and U9400 (N_9400,N_6490,N_5252);
and U9401 (N_9401,N_5290,N_6483);
and U9402 (N_9402,N_5185,N_6341);
xor U9403 (N_9403,N_6479,N_5061);
nor U9404 (N_9404,N_6257,N_5788);
or U9405 (N_9405,N_5249,N_6444);
or U9406 (N_9406,N_6299,N_7434);
and U9407 (N_9407,N_6916,N_5584);
nor U9408 (N_9408,N_7426,N_5320);
xor U9409 (N_9409,N_5927,N_6698);
nand U9410 (N_9410,N_6181,N_5530);
and U9411 (N_9411,N_6558,N_7292);
nand U9412 (N_9412,N_7195,N_6250);
and U9413 (N_9413,N_6879,N_7127);
nor U9414 (N_9414,N_5251,N_5207);
nor U9415 (N_9415,N_7285,N_7288);
and U9416 (N_9416,N_6807,N_6596);
xor U9417 (N_9417,N_5847,N_5244);
xor U9418 (N_9418,N_5452,N_6862);
nor U9419 (N_9419,N_6538,N_7192);
nor U9420 (N_9420,N_5516,N_6566);
nand U9421 (N_9421,N_5523,N_6066);
and U9422 (N_9422,N_6493,N_5645);
nand U9423 (N_9423,N_5173,N_5423);
xor U9424 (N_9424,N_5902,N_5289);
and U9425 (N_9425,N_5014,N_5818);
and U9426 (N_9426,N_6542,N_5376);
and U9427 (N_9427,N_5929,N_6103);
nand U9428 (N_9428,N_5646,N_7073);
xnor U9429 (N_9429,N_6235,N_6107);
nor U9430 (N_9430,N_6163,N_5459);
or U9431 (N_9431,N_6528,N_6502);
nor U9432 (N_9432,N_7098,N_6347);
xor U9433 (N_9433,N_6357,N_7076);
or U9434 (N_9434,N_5463,N_7479);
xnor U9435 (N_9435,N_6777,N_6641);
or U9436 (N_9436,N_5598,N_5553);
nor U9437 (N_9437,N_6896,N_5711);
and U9438 (N_9438,N_6478,N_5560);
and U9439 (N_9439,N_5868,N_7418);
xnor U9440 (N_9440,N_5390,N_7014);
nor U9441 (N_9441,N_5069,N_6895);
nand U9442 (N_9442,N_5062,N_6718);
and U9443 (N_9443,N_5167,N_7229);
and U9444 (N_9444,N_6700,N_5395);
nor U9445 (N_9445,N_5115,N_6746);
xnor U9446 (N_9446,N_7203,N_6997);
nor U9447 (N_9447,N_5855,N_7053);
or U9448 (N_9448,N_6537,N_5582);
nor U9449 (N_9449,N_6179,N_7141);
or U9450 (N_9450,N_6738,N_7425);
or U9451 (N_9451,N_5437,N_5372);
and U9452 (N_9452,N_6302,N_6929);
or U9453 (N_9453,N_7197,N_5621);
and U9454 (N_9454,N_5498,N_6081);
nand U9455 (N_9455,N_6893,N_6611);
nor U9456 (N_9456,N_7369,N_5603);
or U9457 (N_9457,N_5176,N_5556);
and U9458 (N_9458,N_6139,N_5954);
nor U9459 (N_9459,N_5975,N_6298);
xor U9460 (N_9460,N_6698,N_5758);
xnor U9461 (N_9461,N_5799,N_5475);
nor U9462 (N_9462,N_6928,N_5769);
or U9463 (N_9463,N_5507,N_5631);
nor U9464 (N_9464,N_6681,N_5218);
nor U9465 (N_9465,N_7128,N_5447);
nand U9466 (N_9466,N_7482,N_6102);
xor U9467 (N_9467,N_5454,N_5713);
xor U9468 (N_9468,N_7269,N_7186);
nor U9469 (N_9469,N_7490,N_5539);
nor U9470 (N_9470,N_7012,N_6800);
nand U9471 (N_9471,N_6039,N_5269);
and U9472 (N_9472,N_6437,N_5685);
and U9473 (N_9473,N_5087,N_6238);
nor U9474 (N_9474,N_5969,N_6904);
nand U9475 (N_9475,N_5591,N_7104);
nor U9476 (N_9476,N_7207,N_6469);
nand U9477 (N_9477,N_5687,N_5038);
nor U9478 (N_9478,N_6480,N_7198);
nand U9479 (N_9479,N_6432,N_6993);
nor U9480 (N_9480,N_7436,N_6853);
xor U9481 (N_9481,N_6147,N_6716);
or U9482 (N_9482,N_5923,N_5295);
nor U9483 (N_9483,N_6073,N_5417);
and U9484 (N_9484,N_5138,N_7107);
and U9485 (N_9485,N_7132,N_5472);
nand U9486 (N_9486,N_7137,N_5373);
nor U9487 (N_9487,N_7171,N_5551);
and U9488 (N_9488,N_7468,N_6545);
nor U9489 (N_9489,N_5833,N_6659);
nand U9490 (N_9490,N_6662,N_6596);
nand U9491 (N_9491,N_6112,N_5871);
or U9492 (N_9492,N_5463,N_7084);
nand U9493 (N_9493,N_6977,N_6998);
nand U9494 (N_9494,N_6542,N_6582);
or U9495 (N_9495,N_6698,N_7134);
xor U9496 (N_9496,N_7399,N_5959);
and U9497 (N_9497,N_6827,N_5249);
xnor U9498 (N_9498,N_7038,N_7397);
and U9499 (N_9499,N_7268,N_7423);
nor U9500 (N_9500,N_7037,N_7047);
nor U9501 (N_9501,N_5410,N_7189);
nor U9502 (N_9502,N_5926,N_6533);
nand U9503 (N_9503,N_5616,N_5167);
nor U9504 (N_9504,N_6034,N_5501);
nor U9505 (N_9505,N_5349,N_5209);
or U9506 (N_9506,N_5730,N_5838);
or U9507 (N_9507,N_6756,N_5559);
and U9508 (N_9508,N_5918,N_5964);
nand U9509 (N_9509,N_6643,N_5616);
nand U9510 (N_9510,N_7294,N_5294);
or U9511 (N_9511,N_6691,N_7178);
nor U9512 (N_9512,N_6962,N_6080);
and U9513 (N_9513,N_5977,N_7457);
and U9514 (N_9514,N_5262,N_6986);
or U9515 (N_9515,N_5972,N_7145);
nand U9516 (N_9516,N_5951,N_7413);
nand U9517 (N_9517,N_6727,N_6477);
nand U9518 (N_9518,N_6702,N_6490);
and U9519 (N_9519,N_7308,N_5017);
or U9520 (N_9520,N_7088,N_6091);
nand U9521 (N_9521,N_7072,N_7074);
or U9522 (N_9522,N_6014,N_5478);
nand U9523 (N_9523,N_5288,N_7355);
nand U9524 (N_9524,N_5199,N_6230);
nor U9525 (N_9525,N_5771,N_5904);
nor U9526 (N_9526,N_7114,N_5351);
nor U9527 (N_9527,N_6804,N_7247);
or U9528 (N_9528,N_6729,N_6650);
nor U9529 (N_9529,N_5269,N_7293);
and U9530 (N_9530,N_6458,N_5914);
nor U9531 (N_9531,N_5348,N_5886);
or U9532 (N_9532,N_7139,N_5169);
nand U9533 (N_9533,N_6356,N_5652);
and U9534 (N_9534,N_6208,N_6558);
nor U9535 (N_9535,N_7058,N_6337);
nand U9536 (N_9536,N_5009,N_6417);
and U9537 (N_9537,N_6506,N_7436);
nand U9538 (N_9538,N_5555,N_6852);
xor U9539 (N_9539,N_6228,N_6832);
xnor U9540 (N_9540,N_5586,N_5937);
and U9541 (N_9541,N_6959,N_7454);
xnor U9542 (N_9542,N_5265,N_6507);
nand U9543 (N_9543,N_7382,N_6556);
nand U9544 (N_9544,N_7402,N_6979);
and U9545 (N_9545,N_5673,N_7388);
or U9546 (N_9546,N_6674,N_5812);
and U9547 (N_9547,N_6835,N_5443);
nand U9548 (N_9548,N_6112,N_6044);
nor U9549 (N_9549,N_5840,N_7086);
and U9550 (N_9550,N_6417,N_6222);
nor U9551 (N_9551,N_7412,N_6413);
or U9552 (N_9552,N_6061,N_6267);
xnor U9553 (N_9553,N_7197,N_5226);
xor U9554 (N_9554,N_6839,N_6500);
and U9555 (N_9555,N_7066,N_5015);
or U9556 (N_9556,N_5949,N_5634);
nand U9557 (N_9557,N_5811,N_6771);
or U9558 (N_9558,N_7231,N_5463);
or U9559 (N_9559,N_5601,N_6323);
nor U9560 (N_9560,N_5094,N_5500);
and U9561 (N_9561,N_5744,N_6148);
nand U9562 (N_9562,N_6499,N_7300);
nor U9563 (N_9563,N_5572,N_6146);
nor U9564 (N_9564,N_5120,N_6499);
nor U9565 (N_9565,N_6208,N_6196);
nor U9566 (N_9566,N_6278,N_7473);
xnor U9567 (N_9567,N_5640,N_6255);
nand U9568 (N_9568,N_6527,N_6469);
xor U9569 (N_9569,N_6116,N_6891);
nand U9570 (N_9570,N_5224,N_5205);
nand U9571 (N_9571,N_6785,N_5555);
and U9572 (N_9572,N_6425,N_6311);
and U9573 (N_9573,N_7282,N_6009);
and U9574 (N_9574,N_5508,N_5984);
or U9575 (N_9575,N_5969,N_6554);
nand U9576 (N_9576,N_6639,N_7311);
nor U9577 (N_9577,N_6909,N_5491);
xor U9578 (N_9578,N_7438,N_5180);
nand U9579 (N_9579,N_5596,N_6704);
and U9580 (N_9580,N_7184,N_7402);
nor U9581 (N_9581,N_6838,N_6945);
nand U9582 (N_9582,N_5321,N_6732);
and U9583 (N_9583,N_7450,N_6261);
nor U9584 (N_9584,N_6480,N_5603);
and U9585 (N_9585,N_7291,N_6968);
and U9586 (N_9586,N_6311,N_5230);
or U9587 (N_9587,N_5321,N_5170);
nand U9588 (N_9588,N_7432,N_7240);
and U9589 (N_9589,N_5630,N_5562);
and U9590 (N_9590,N_6870,N_6597);
nor U9591 (N_9591,N_6163,N_5678);
and U9592 (N_9592,N_5034,N_5228);
and U9593 (N_9593,N_5160,N_5942);
nor U9594 (N_9594,N_6797,N_6478);
and U9595 (N_9595,N_7400,N_6823);
nor U9596 (N_9596,N_5587,N_5910);
and U9597 (N_9597,N_5360,N_5030);
nor U9598 (N_9598,N_5955,N_5058);
xor U9599 (N_9599,N_7482,N_6539);
nand U9600 (N_9600,N_5835,N_5416);
or U9601 (N_9601,N_5747,N_6886);
nand U9602 (N_9602,N_7154,N_5664);
nor U9603 (N_9603,N_6871,N_5073);
and U9604 (N_9604,N_6765,N_5184);
nor U9605 (N_9605,N_7235,N_6435);
and U9606 (N_9606,N_6218,N_6307);
nand U9607 (N_9607,N_5389,N_6627);
xor U9608 (N_9608,N_7481,N_6657);
or U9609 (N_9609,N_6718,N_5804);
nand U9610 (N_9610,N_5654,N_5920);
nor U9611 (N_9611,N_5150,N_6640);
nor U9612 (N_9612,N_7404,N_6432);
nand U9613 (N_9613,N_5664,N_5436);
nor U9614 (N_9614,N_5447,N_7302);
nor U9615 (N_9615,N_7048,N_6792);
xnor U9616 (N_9616,N_6486,N_7322);
nor U9617 (N_9617,N_5843,N_6296);
nor U9618 (N_9618,N_7066,N_7424);
nor U9619 (N_9619,N_6294,N_7096);
xor U9620 (N_9620,N_6703,N_5418);
nand U9621 (N_9621,N_6204,N_5887);
nor U9622 (N_9622,N_6955,N_5256);
nand U9623 (N_9623,N_6475,N_6918);
nand U9624 (N_9624,N_6251,N_7002);
and U9625 (N_9625,N_6351,N_6952);
nand U9626 (N_9626,N_6608,N_6664);
and U9627 (N_9627,N_5497,N_5880);
or U9628 (N_9628,N_5124,N_7368);
and U9629 (N_9629,N_5340,N_5150);
or U9630 (N_9630,N_7042,N_7025);
and U9631 (N_9631,N_5390,N_5436);
or U9632 (N_9632,N_6393,N_5729);
xnor U9633 (N_9633,N_6081,N_6274);
nand U9634 (N_9634,N_5387,N_5878);
nor U9635 (N_9635,N_6658,N_7290);
nand U9636 (N_9636,N_5616,N_7445);
nand U9637 (N_9637,N_5427,N_5019);
nor U9638 (N_9638,N_5321,N_7086);
nor U9639 (N_9639,N_7209,N_7459);
xor U9640 (N_9640,N_6026,N_6946);
nand U9641 (N_9641,N_5719,N_6006);
and U9642 (N_9642,N_7106,N_7004);
nand U9643 (N_9643,N_5077,N_5104);
nand U9644 (N_9644,N_5960,N_6768);
and U9645 (N_9645,N_5841,N_6884);
or U9646 (N_9646,N_7183,N_5841);
nand U9647 (N_9647,N_7181,N_5013);
nand U9648 (N_9648,N_5721,N_5891);
and U9649 (N_9649,N_6557,N_6300);
or U9650 (N_9650,N_5137,N_5880);
nor U9651 (N_9651,N_7431,N_6399);
nand U9652 (N_9652,N_7130,N_6554);
and U9653 (N_9653,N_7126,N_5693);
and U9654 (N_9654,N_7365,N_6009);
nand U9655 (N_9655,N_5395,N_5407);
nand U9656 (N_9656,N_7477,N_6121);
or U9657 (N_9657,N_6794,N_6103);
and U9658 (N_9658,N_5667,N_5153);
nor U9659 (N_9659,N_6040,N_6249);
nand U9660 (N_9660,N_6511,N_5374);
nand U9661 (N_9661,N_5823,N_5235);
nand U9662 (N_9662,N_6564,N_7058);
and U9663 (N_9663,N_6948,N_7056);
nor U9664 (N_9664,N_5368,N_5397);
nor U9665 (N_9665,N_6031,N_6223);
nand U9666 (N_9666,N_5450,N_6488);
nor U9667 (N_9667,N_6724,N_6450);
nor U9668 (N_9668,N_6345,N_6995);
nand U9669 (N_9669,N_5981,N_6758);
nand U9670 (N_9670,N_6371,N_6432);
or U9671 (N_9671,N_5147,N_7295);
nor U9672 (N_9672,N_7481,N_5523);
or U9673 (N_9673,N_6650,N_5823);
or U9674 (N_9674,N_6077,N_6957);
and U9675 (N_9675,N_7176,N_6327);
nand U9676 (N_9676,N_7218,N_5327);
and U9677 (N_9677,N_5652,N_6919);
nand U9678 (N_9678,N_6428,N_6302);
nand U9679 (N_9679,N_7006,N_6978);
nand U9680 (N_9680,N_7260,N_7177);
and U9681 (N_9681,N_6394,N_5204);
nor U9682 (N_9682,N_6216,N_6839);
nor U9683 (N_9683,N_6220,N_6019);
or U9684 (N_9684,N_7223,N_5894);
or U9685 (N_9685,N_5209,N_6291);
nor U9686 (N_9686,N_6622,N_6848);
nand U9687 (N_9687,N_5131,N_6208);
and U9688 (N_9688,N_6256,N_7233);
nor U9689 (N_9689,N_5143,N_6717);
or U9690 (N_9690,N_6899,N_7057);
xor U9691 (N_9691,N_6591,N_5834);
and U9692 (N_9692,N_6802,N_5523);
nand U9693 (N_9693,N_7222,N_6956);
or U9694 (N_9694,N_7386,N_6622);
and U9695 (N_9695,N_7338,N_6541);
nand U9696 (N_9696,N_7324,N_5145);
or U9697 (N_9697,N_5259,N_5582);
nor U9698 (N_9698,N_6056,N_6859);
nor U9699 (N_9699,N_5047,N_5269);
and U9700 (N_9700,N_5549,N_5582);
nor U9701 (N_9701,N_5544,N_5910);
and U9702 (N_9702,N_6764,N_5237);
nor U9703 (N_9703,N_5486,N_5959);
nor U9704 (N_9704,N_5729,N_5704);
or U9705 (N_9705,N_5526,N_5043);
and U9706 (N_9706,N_7079,N_6181);
nor U9707 (N_9707,N_6342,N_7366);
nor U9708 (N_9708,N_5683,N_7055);
or U9709 (N_9709,N_6645,N_7033);
and U9710 (N_9710,N_7215,N_5884);
xor U9711 (N_9711,N_6066,N_6644);
nor U9712 (N_9712,N_5958,N_6269);
nor U9713 (N_9713,N_5385,N_6600);
nand U9714 (N_9714,N_7076,N_5842);
xor U9715 (N_9715,N_6394,N_7368);
or U9716 (N_9716,N_5588,N_6052);
and U9717 (N_9717,N_7038,N_7117);
nand U9718 (N_9718,N_5620,N_5636);
and U9719 (N_9719,N_6777,N_6564);
nand U9720 (N_9720,N_6522,N_6445);
nor U9721 (N_9721,N_5407,N_5725);
and U9722 (N_9722,N_5161,N_6624);
xnor U9723 (N_9723,N_7049,N_7017);
nor U9724 (N_9724,N_7198,N_6231);
nand U9725 (N_9725,N_6723,N_6389);
nor U9726 (N_9726,N_5866,N_5386);
and U9727 (N_9727,N_5035,N_5356);
xor U9728 (N_9728,N_6783,N_5710);
and U9729 (N_9729,N_7326,N_5934);
nand U9730 (N_9730,N_5475,N_5463);
nor U9731 (N_9731,N_7053,N_6170);
nor U9732 (N_9732,N_5043,N_6088);
or U9733 (N_9733,N_5160,N_5023);
and U9734 (N_9734,N_6357,N_6462);
or U9735 (N_9735,N_5935,N_7351);
nand U9736 (N_9736,N_5217,N_6175);
nand U9737 (N_9737,N_6747,N_6959);
or U9738 (N_9738,N_5559,N_5876);
nand U9739 (N_9739,N_6245,N_5930);
and U9740 (N_9740,N_5929,N_5911);
or U9741 (N_9741,N_5771,N_5035);
or U9742 (N_9742,N_5703,N_5282);
nand U9743 (N_9743,N_7257,N_7464);
or U9744 (N_9744,N_7285,N_6798);
nand U9745 (N_9745,N_5164,N_5855);
nand U9746 (N_9746,N_5685,N_7239);
or U9747 (N_9747,N_5021,N_7282);
nand U9748 (N_9748,N_7278,N_6667);
nor U9749 (N_9749,N_5885,N_6913);
nand U9750 (N_9750,N_5488,N_5757);
nor U9751 (N_9751,N_6278,N_7403);
nand U9752 (N_9752,N_6200,N_5747);
xor U9753 (N_9753,N_6402,N_5687);
nand U9754 (N_9754,N_5654,N_5441);
nor U9755 (N_9755,N_6330,N_5519);
xnor U9756 (N_9756,N_6851,N_6793);
and U9757 (N_9757,N_5178,N_6618);
or U9758 (N_9758,N_5143,N_5949);
nor U9759 (N_9759,N_7418,N_7192);
nand U9760 (N_9760,N_6773,N_6167);
nand U9761 (N_9761,N_7169,N_6860);
xor U9762 (N_9762,N_5903,N_6999);
nand U9763 (N_9763,N_5568,N_5287);
nor U9764 (N_9764,N_5320,N_5351);
nand U9765 (N_9765,N_7082,N_7471);
or U9766 (N_9766,N_5597,N_6566);
and U9767 (N_9767,N_5152,N_6599);
nand U9768 (N_9768,N_5910,N_5804);
or U9769 (N_9769,N_7056,N_5495);
xnor U9770 (N_9770,N_5769,N_6075);
nand U9771 (N_9771,N_6934,N_5249);
or U9772 (N_9772,N_6363,N_5332);
xor U9773 (N_9773,N_7403,N_6535);
xnor U9774 (N_9774,N_5743,N_6982);
or U9775 (N_9775,N_7092,N_5056);
or U9776 (N_9776,N_6630,N_6493);
and U9777 (N_9777,N_7426,N_6412);
nor U9778 (N_9778,N_7391,N_7215);
and U9779 (N_9779,N_5839,N_5349);
nand U9780 (N_9780,N_6038,N_5979);
nand U9781 (N_9781,N_7081,N_7456);
nand U9782 (N_9782,N_7473,N_6419);
or U9783 (N_9783,N_5056,N_7205);
and U9784 (N_9784,N_5497,N_5712);
or U9785 (N_9785,N_6282,N_7064);
nor U9786 (N_9786,N_5959,N_5336);
and U9787 (N_9787,N_6670,N_7131);
nand U9788 (N_9788,N_6060,N_5436);
and U9789 (N_9789,N_7050,N_7062);
nand U9790 (N_9790,N_7261,N_5891);
or U9791 (N_9791,N_7389,N_5942);
xor U9792 (N_9792,N_6542,N_5789);
and U9793 (N_9793,N_5750,N_5303);
nand U9794 (N_9794,N_7474,N_5942);
nor U9795 (N_9795,N_6073,N_6373);
nand U9796 (N_9796,N_6053,N_6787);
nand U9797 (N_9797,N_6388,N_6910);
and U9798 (N_9798,N_6376,N_7331);
and U9799 (N_9799,N_6389,N_5374);
nand U9800 (N_9800,N_5107,N_5421);
or U9801 (N_9801,N_5308,N_7065);
nor U9802 (N_9802,N_6414,N_5477);
or U9803 (N_9803,N_5082,N_7277);
nand U9804 (N_9804,N_6877,N_6487);
nor U9805 (N_9805,N_5530,N_5974);
nor U9806 (N_9806,N_6526,N_6772);
nor U9807 (N_9807,N_5941,N_5775);
and U9808 (N_9808,N_7152,N_5991);
nand U9809 (N_9809,N_7242,N_7411);
nor U9810 (N_9810,N_7156,N_7384);
nand U9811 (N_9811,N_5440,N_7214);
or U9812 (N_9812,N_6158,N_6630);
xor U9813 (N_9813,N_5520,N_6360);
nor U9814 (N_9814,N_6690,N_5326);
nand U9815 (N_9815,N_5633,N_7302);
nand U9816 (N_9816,N_7308,N_6107);
and U9817 (N_9817,N_7146,N_6598);
nand U9818 (N_9818,N_6392,N_7382);
nand U9819 (N_9819,N_5261,N_7094);
nor U9820 (N_9820,N_7079,N_6358);
nand U9821 (N_9821,N_6121,N_6700);
nor U9822 (N_9822,N_6724,N_6558);
xor U9823 (N_9823,N_5604,N_5904);
xnor U9824 (N_9824,N_5306,N_6492);
nand U9825 (N_9825,N_5723,N_5951);
or U9826 (N_9826,N_5536,N_7366);
or U9827 (N_9827,N_6579,N_7441);
nand U9828 (N_9828,N_5728,N_6797);
nor U9829 (N_9829,N_7471,N_6716);
nor U9830 (N_9830,N_5185,N_6021);
xnor U9831 (N_9831,N_7155,N_5449);
and U9832 (N_9832,N_6015,N_5518);
nor U9833 (N_9833,N_6222,N_6788);
xor U9834 (N_9834,N_7318,N_5277);
or U9835 (N_9835,N_7214,N_5851);
nor U9836 (N_9836,N_6237,N_5221);
or U9837 (N_9837,N_6582,N_6634);
nand U9838 (N_9838,N_5898,N_6882);
nor U9839 (N_9839,N_6775,N_6273);
nand U9840 (N_9840,N_6435,N_5272);
nand U9841 (N_9841,N_5225,N_5220);
nor U9842 (N_9842,N_5125,N_7110);
nor U9843 (N_9843,N_7162,N_5585);
and U9844 (N_9844,N_5105,N_5685);
xor U9845 (N_9845,N_5983,N_7158);
and U9846 (N_9846,N_5204,N_7247);
nand U9847 (N_9847,N_5767,N_6964);
and U9848 (N_9848,N_6512,N_5334);
or U9849 (N_9849,N_5628,N_5642);
xor U9850 (N_9850,N_6509,N_6845);
xnor U9851 (N_9851,N_7491,N_5812);
and U9852 (N_9852,N_6937,N_5386);
nand U9853 (N_9853,N_7010,N_6446);
and U9854 (N_9854,N_7426,N_5173);
and U9855 (N_9855,N_5366,N_5239);
nor U9856 (N_9856,N_6361,N_5632);
and U9857 (N_9857,N_6085,N_5745);
nand U9858 (N_9858,N_7091,N_5717);
xnor U9859 (N_9859,N_5457,N_6414);
nor U9860 (N_9860,N_6935,N_7238);
nor U9861 (N_9861,N_5424,N_7351);
and U9862 (N_9862,N_6094,N_6208);
nor U9863 (N_9863,N_5758,N_7286);
and U9864 (N_9864,N_6411,N_5296);
nor U9865 (N_9865,N_5934,N_6787);
or U9866 (N_9866,N_6882,N_6233);
and U9867 (N_9867,N_6764,N_6498);
nor U9868 (N_9868,N_6893,N_6934);
or U9869 (N_9869,N_6427,N_7157);
nand U9870 (N_9870,N_7018,N_6938);
and U9871 (N_9871,N_5774,N_6128);
nor U9872 (N_9872,N_6578,N_5722);
nand U9873 (N_9873,N_7072,N_6128);
xor U9874 (N_9874,N_5692,N_6108);
or U9875 (N_9875,N_5557,N_5379);
or U9876 (N_9876,N_7334,N_6974);
nand U9877 (N_9877,N_5985,N_5684);
nor U9878 (N_9878,N_5374,N_5153);
or U9879 (N_9879,N_6054,N_5184);
nor U9880 (N_9880,N_7498,N_6643);
xnor U9881 (N_9881,N_6403,N_5265);
nor U9882 (N_9882,N_7095,N_5919);
or U9883 (N_9883,N_6492,N_5299);
or U9884 (N_9884,N_7446,N_6520);
or U9885 (N_9885,N_7384,N_6460);
and U9886 (N_9886,N_5412,N_7003);
nor U9887 (N_9887,N_6626,N_7005);
nor U9888 (N_9888,N_6747,N_5346);
and U9889 (N_9889,N_7095,N_7177);
and U9890 (N_9890,N_5031,N_6470);
or U9891 (N_9891,N_7298,N_7352);
nand U9892 (N_9892,N_6388,N_7181);
and U9893 (N_9893,N_5754,N_6803);
or U9894 (N_9894,N_6117,N_6672);
and U9895 (N_9895,N_6667,N_6037);
nor U9896 (N_9896,N_5568,N_6088);
or U9897 (N_9897,N_6518,N_5262);
and U9898 (N_9898,N_5071,N_5378);
nand U9899 (N_9899,N_6057,N_7324);
and U9900 (N_9900,N_5063,N_5751);
xor U9901 (N_9901,N_5858,N_5379);
or U9902 (N_9902,N_6778,N_5339);
nand U9903 (N_9903,N_5439,N_5906);
or U9904 (N_9904,N_6571,N_5379);
xnor U9905 (N_9905,N_6962,N_6629);
nand U9906 (N_9906,N_5496,N_5237);
and U9907 (N_9907,N_6177,N_5000);
nor U9908 (N_9908,N_5038,N_5093);
nand U9909 (N_9909,N_5768,N_5890);
nand U9910 (N_9910,N_5001,N_7281);
and U9911 (N_9911,N_5622,N_6693);
and U9912 (N_9912,N_5664,N_5921);
nor U9913 (N_9913,N_5007,N_7397);
and U9914 (N_9914,N_5744,N_5329);
nand U9915 (N_9915,N_6353,N_5962);
or U9916 (N_9916,N_6777,N_6543);
and U9917 (N_9917,N_6729,N_5927);
or U9918 (N_9918,N_7401,N_6165);
xor U9919 (N_9919,N_6500,N_5770);
or U9920 (N_9920,N_5489,N_7323);
nand U9921 (N_9921,N_6744,N_5450);
nand U9922 (N_9922,N_6737,N_6453);
nor U9923 (N_9923,N_6708,N_5129);
or U9924 (N_9924,N_6984,N_5922);
or U9925 (N_9925,N_6122,N_5344);
nand U9926 (N_9926,N_6225,N_6709);
nor U9927 (N_9927,N_5978,N_7257);
or U9928 (N_9928,N_5878,N_6494);
or U9929 (N_9929,N_5355,N_5008);
nand U9930 (N_9930,N_7311,N_5682);
nor U9931 (N_9931,N_5632,N_5449);
nor U9932 (N_9932,N_5830,N_5173);
nand U9933 (N_9933,N_7315,N_5049);
nor U9934 (N_9934,N_7353,N_5890);
or U9935 (N_9935,N_5727,N_7416);
xnor U9936 (N_9936,N_5081,N_7161);
or U9937 (N_9937,N_7450,N_7166);
and U9938 (N_9938,N_5557,N_6727);
nor U9939 (N_9939,N_6322,N_6274);
or U9940 (N_9940,N_6727,N_6879);
nand U9941 (N_9941,N_7176,N_6545);
xnor U9942 (N_9942,N_6243,N_7420);
xor U9943 (N_9943,N_6726,N_5789);
nor U9944 (N_9944,N_5875,N_5669);
or U9945 (N_9945,N_6307,N_7402);
or U9946 (N_9946,N_6129,N_5352);
or U9947 (N_9947,N_6914,N_5298);
nor U9948 (N_9948,N_6530,N_6930);
nand U9949 (N_9949,N_5726,N_6395);
nand U9950 (N_9950,N_7138,N_5610);
and U9951 (N_9951,N_6395,N_6852);
nand U9952 (N_9952,N_7128,N_6358);
nand U9953 (N_9953,N_5257,N_5895);
nand U9954 (N_9954,N_5752,N_6877);
nand U9955 (N_9955,N_6660,N_5819);
and U9956 (N_9956,N_6889,N_6465);
nor U9957 (N_9957,N_5479,N_7021);
nand U9958 (N_9958,N_5583,N_5494);
xor U9959 (N_9959,N_5452,N_7191);
nand U9960 (N_9960,N_6962,N_5134);
nand U9961 (N_9961,N_6260,N_5293);
or U9962 (N_9962,N_5157,N_7370);
or U9963 (N_9963,N_5545,N_6737);
nor U9964 (N_9964,N_7398,N_6844);
and U9965 (N_9965,N_5370,N_5324);
or U9966 (N_9966,N_5728,N_5804);
and U9967 (N_9967,N_5068,N_5642);
or U9968 (N_9968,N_5939,N_6313);
nand U9969 (N_9969,N_7079,N_7066);
nor U9970 (N_9970,N_5357,N_5216);
nor U9971 (N_9971,N_5250,N_5156);
and U9972 (N_9972,N_5765,N_6710);
nor U9973 (N_9973,N_5993,N_5626);
xor U9974 (N_9974,N_7395,N_5535);
xor U9975 (N_9975,N_6181,N_6796);
xor U9976 (N_9976,N_6641,N_6675);
or U9977 (N_9977,N_6291,N_7415);
nor U9978 (N_9978,N_7157,N_6236);
or U9979 (N_9979,N_7158,N_5776);
nand U9980 (N_9980,N_6266,N_5814);
or U9981 (N_9981,N_6553,N_6943);
nor U9982 (N_9982,N_5360,N_5969);
nand U9983 (N_9983,N_5772,N_7309);
and U9984 (N_9984,N_5667,N_6657);
or U9985 (N_9985,N_5405,N_5321);
nor U9986 (N_9986,N_6321,N_5288);
nand U9987 (N_9987,N_6115,N_5323);
nor U9988 (N_9988,N_6318,N_5036);
or U9989 (N_9989,N_5004,N_5982);
nand U9990 (N_9990,N_5354,N_6251);
or U9991 (N_9991,N_7460,N_7272);
nand U9992 (N_9992,N_6463,N_5604);
nand U9993 (N_9993,N_5412,N_6671);
nand U9994 (N_9994,N_5166,N_6896);
xor U9995 (N_9995,N_5476,N_5931);
nor U9996 (N_9996,N_7029,N_5736);
and U9997 (N_9997,N_7242,N_5513);
nor U9998 (N_9998,N_5436,N_7061);
nand U9999 (N_9999,N_6786,N_5034);
nand UO_0 (O_0,N_9199,N_9871);
nor UO_1 (O_1,N_8638,N_8347);
or UO_2 (O_2,N_9458,N_8339);
nand UO_3 (O_3,N_8644,N_8536);
and UO_4 (O_4,N_7718,N_8327);
xnor UO_5 (O_5,N_9221,N_8835);
nand UO_6 (O_6,N_8374,N_9299);
nand UO_7 (O_7,N_7649,N_7747);
nand UO_8 (O_8,N_8175,N_9705);
and UO_9 (O_9,N_9203,N_8025);
nand UO_10 (O_10,N_7650,N_9253);
and UO_11 (O_11,N_8732,N_7825);
nand UO_12 (O_12,N_8600,N_7990);
nor UO_13 (O_13,N_9611,N_9306);
nor UO_14 (O_14,N_9171,N_9113);
or UO_15 (O_15,N_9680,N_8748);
nor UO_16 (O_16,N_8656,N_7844);
xor UO_17 (O_17,N_7814,N_8406);
nand UO_18 (O_18,N_9892,N_9679);
nor UO_19 (O_19,N_9977,N_8125);
nand UO_20 (O_20,N_7622,N_9303);
nor UO_21 (O_21,N_9077,N_8144);
xor UO_22 (O_22,N_8430,N_9998);
nand UO_23 (O_23,N_8287,N_9751);
or UO_24 (O_24,N_7681,N_9169);
nand UO_25 (O_25,N_9534,N_7989);
nor UO_26 (O_26,N_9548,N_9401);
xnor UO_27 (O_27,N_7769,N_7917);
or UO_28 (O_28,N_8167,N_8359);
or UO_29 (O_29,N_8838,N_8940);
nand UO_30 (O_30,N_9730,N_7898);
and UO_31 (O_31,N_9724,N_8106);
and UO_32 (O_32,N_7738,N_9387);
or UO_33 (O_33,N_8087,N_8276);
nor UO_34 (O_34,N_8621,N_8051);
or UO_35 (O_35,N_9276,N_9902);
or UO_36 (O_36,N_9536,N_9432);
nand UO_37 (O_37,N_8229,N_9281);
or UO_38 (O_38,N_8633,N_8995);
or UO_39 (O_39,N_9675,N_9807);
xnor UO_40 (O_40,N_8481,N_8756);
nor UO_41 (O_41,N_9556,N_9987);
nor UO_42 (O_42,N_8804,N_7693);
nor UO_43 (O_43,N_9076,N_8831);
or UO_44 (O_44,N_9592,N_7907);
nand UO_45 (O_45,N_9094,N_9402);
nor UO_46 (O_46,N_7624,N_9634);
nor UO_47 (O_47,N_7656,N_8341);
nor UO_48 (O_48,N_9971,N_8516);
nor UO_49 (O_49,N_9989,N_9835);
and UO_50 (O_50,N_8529,N_9850);
nand UO_51 (O_51,N_9784,N_9275);
xor UO_52 (O_52,N_7831,N_8710);
and UO_53 (O_53,N_7757,N_9563);
nor UO_54 (O_54,N_9547,N_9758);
and UO_55 (O_55,N_8016,N_9443);
or UO_56 (O_56,N_8560,N_7620);
xnor UO_57 (O_57,N_8140,N_9689);
and UO_58 (O_58,N_9124,N_8260);
nor UO_59 (O_59,N_8288,N_8899);
or UO_60 (O_60,N_9263,N_9464);
nand UO_61 (O_61,N_9215,N_8969);
nor UO_62 (O_62,N_8269,N_9994);
nor UO_63 (O_63,N_9629,N_8424);
and UO_64 (O_64,N_9362,N_8258);
nand UO_65 (O_65,N_8188,N_9656);
nand UO_66 (O_66,N_9115,N_8426);
or UO_67 (O_67,N_9390,N_9182);
and UO_68 (O_68,N_9308,N_8095);
xnor UO_69 (O_69,N_7686,N_9213);
nand UO_70 (O_70,N_9144,N_8415);
nand UO_71 (O_71,N_8189,N_9060);
xnor UO_72 (O_72,N_9039,N_9489);
nor UO_73 (O_73,N_9995,N_8538);
or UO_74 (O_74,N_8350,N_8416);
and UO_75 (O_75,N_9301,N_8636);
nand UO_76 (O_76,N_8041,N_7748);
and UO_77 (O_77,N_8963,N_7500);
and UO_78 (O_78,N_9565,N_8300);
nand UO_79 (O_79,N_9941,N_9559);
and UO_80 (O_80,N_8413,N_9176);
or UO_81 (O_81,N_8528,N_9571);
nor UO_82 (O_82,N_9343,N_8403);
or UO_83 (O_83,N_7753,N_9778);
or UO_84 (O_84,N_8314,N_9475);
or UO_85 (O_85,N_7735,N_7873);
nor UO_86 (O_86,N_9555,N_7941);
and UO_87 (O_87,N_7840,N_9787);
and UO_88 (O_88,N_8020,N_9785);
and UO_89 (O_89,N_9319,N_7521);
nand UO_90 (O_90,N_8544,N_8987);
or UO_91 (O_91,N_9716,N_9293);
or UO_92 (O_92,N_9922,N_9980);
or UO_93 (O_93,N_8859,N_7630);
nor UO_94 (O_94,N_9649,N_9480);
nand UO_95 (O_95,N_9921,N_7934);
nor UO_96 (O_96,N_8550,N_7618);
nand UO_97 (O_97,N_9156,N_9430);
and UO_98 (O_98,N_9037,N_8663);
and UO_99 (O_99,N_8027,N_8923);
or UO_100 (O_100,N_9292,N_7691);
nor UO_101 (O_101,N_9631,N_9635);
nand UO_102 (O_102,N_9976,N_9471);
or UO_103 (O_103,N_9827,N_9873);
nand UO_104 (O_104,N_8060,N_8321);
nor UO_105 (O_105,N_7755,N_8142);
nor UO_106 (O_106,N_9075,N_9822);
nor UO_107 (O_107,N_9975,N_7616);
nand UO_108 (O_108,N_8852,N_8553);
or UO_109 (O_109,N_8834,N_8580);
nor UO_110 (O_110,N_8427,N_8344);
nor UO_111 (O_111,N_7996,N_8612);
or UO_112 (O_112,N_9054,N_8883);
and UO_113 (O_113,N_9677,N_7629);
nor UO_114 (O_114,N_8767,N_7929);
or UO_115 (O_115,N_8932,N_7577);
or UO_116 (O_116,N_8019,N_8608);
or UO_117 (O_117,N_9441,N_9371);
or UO_118 (O_118,N_7565,N_8185);
and UO_119 (O_119,N_9044,N_8240);
or UO_120 (O_120,N_9775,N_9396);
nor UO_121 (O_121,N_9021,N_9715);
nand UO_122 (O_122,N_9567,N_7696);
or UO_123 (O_123,N_8851,N_9377);
nor UO_124 (O_124,N_8113,N_8057);
and UO_125 (O_125,N_7692,N_8825);
or UO_126 (O_126,N_8989,N_9662);
and UO_127 (O_127,N_7986,N_7672);
and UO_128 (O_128,N_7984,N_9569);
nand UO_129 (O_129,N_9200,N_9719);
nand UO_130 (O_130,N_9046,N_9435);
and UO_131 (O_131,N_9013,N_8094);
xor UO_132 (O_132,N_8527,N_9884);
nor UO_133 (O_133,N_7612,N_8688);
and UO_134 (O_134,N_9260,N_9118);
and UO_135 (O_135,N_9320,N_8813);
nand UO_136 (O_136,N_7522,N_8784);
or UO_137 (O_137,N_8037,N_7581);
nand UO_138 (O_138,N_9874,N_9544);
and UO_139 (O_139,N_8387,N_8259);
nand UO_140 (O_140,N_9478,N_8872);
or UO_141 (O_141,N_9376,N_9222);
xnor UO_142 (O_142,N_8959,N_9947);
nand UO_143 (O_143,N_7886,N_8283);
nand UO_144 (O_144,N_9476,N_7988);
or UO_145 (O_145,N_8824,N_8043);
nor UO_146 (O_146,N_8653,N_9063);
xnor UO_147 (O_147,N_9878,N_8422);
or UO_148 (O_148,N_7611,N_8482);
nand UO_149 (O_149,N_8614,N_8237);
or UO_150 (O_150,N_8026,N_7955);
nor UO_151 (O_151,N_7883,N_9379);
or UO_152 (O_152,N_8072,N_9473);
and UO_153 (O_153,N_9419,N_7527);
nand UO_154 (O_154,N_9523,N_8483);
nor UO_155 (O_155,N_8626,N_8996);
and UO_156 (O_156,N_9513,N_9288);
nor UO_157 (O_157,N_8924,N_8707);
nand UO_158 (O_158,N_9731,N_8061);
nor UO_159 (O_159,N_9707,N_8058);
nand UO_160 (O_160,N_9918,N_9713);
nor UO_161 (O_161,N_9728,N_9484);
or UO_162 (O_162,N_9851,N_9620);
and UO_163 (O_163,N_9907,N_7517);
xnor UO_164 (O_164,N_8388,N_9696);
nor UO_165 (O_165,N_9290,N_9128);
nand UO_166 (O_166,N_7701,N_9370);
nor UO_167 (O_167,N_7991,N_8428);
nand UO_168 (O_168,N_8267,N_8233);
and UO_169 (O_169,N_7561,N_8050);
nand UO_170 (O_170,N_8377,N_8470);
and UO_171 (O_171,N_9655,N_9912);
or UO_172 (O_172,N_8809,N_9336);
or UO_173 (O_173,N_8593,N_8082);
and UO_174 (O_174,N_7827,N_8193);
or UO_175 (O_175,N_9641,N_7774);
or UO_176 (O_176,N_9624,N_8751);
or UO_177 (O_177,N_9619,N_8418);
or UO_178 (O_178,N_8992,N_7793);
xor UO_179 (O_179,N_8857,N_9261);
and UO_180 (O_180,N_7592,N_9463);
or UO_181 (O_181,N_8137,N_7635);
nand UO_182 (O_182,N_7657,N_9196);
or UO_183 (O_183,N_9442,N_8204);
and UO_184 (O_184,N_8463,N_9088);
or UO_185 (O_185,N_9810,N_8116);
nor UO_186 (O_186,N_8079,N_9467);
xor UO_187 (O_187,N_9726,N_9310);
and UO_188 (O_188,N_9337,N_9152);
nand UO_189 (O_189,N_8561,N_7567);
and UO_190 (O_190,N_9278,N_9274);
nand UO_191 (O_191,N_9951,N_9923);
and UO_192 (O_192,N_8774,N_9839);
or UO_193 (O_193,N_7981,N_9168);
nand UO_194 (O_194,N_9776,N_8657);
nor UO_195 (O_195,N_8122,N_9955);
nor UO_196 (O_196,N_9174,N_9823);
nand UO_197 (O_197,N_7980,N_9436);
xor UO_198 (O_198,N_9940,N_7968);
and UO_199 (O_199,N_8719,N_8531);
xnor UO_200 (O_200,N_7557,N_9640);
xor UO_201 (O_201,N_8209,N_9027);
or UO_202 (O_202,N_9363,N_7528);
nand UO_203 (O_203,N_8955,N_8076);
and UO_204 (O_204,N_7932,N_7790);
nor UO_205 (O_205,N_9539,N_8713);
nand UO_206 (O_206,N_9127,N_8762);
and UO_207 (O_207,N_9305,N_9796);
nand UO_208 (O_208,N_8107,N_8024);
nand UO_209 (O_209,N_9906,N_8964);
nor UO_210 (O_210,N_8780,N_9950);
or UO_211 (O_211,N_8850,N_9350);
and UO_212 (O_212,N_8207,N_7962);
and UO_213 (O_213,N_8983,N_8284);
nand UO_214 (O_214,N_9036,N_7974);
nor UO_215 (O_215,N_8524,N_9177);
nand UO_216 (O_216,N_8123,N_8680);
and UO_217 (O_217,N_7737,N_7868);
nand UO_218 (O_218,N_7711,N_7538);
and UO_219 (O_219,N_9326,N_8431);
xnor UO_220 (O_220,N_7752,N_9015);
nand UO_221 (O_221,N_8837,N_8136);
xnor UO_222 (O_222,N_7939,N_7781);
xnor UO_223 (O_223,N_8908,N_8453);
or UO_224 (O_224,N_9595,N_7815);
and UO_225 (O_225,N_8429,N_7780);
and UO_226 (O_226,N_7874,N_8046);
xor UO_227 (O_227,N_8298,N_9518);
xor UO_228 (O_228,N_8476,N_8309);
nand UO_229 (O_229,N_9136,N_9045);
xnor UO_230 (O_230,N_9840,N_8942);
and UO_231 (O_231,N_8716,N_9602);
nor UO_232 (O_232,N_8689,N_8412);
nor UO_233 (O_233,N_9485,N_8960);
nor UO_234 (O_234,N_8913,N_8897);
or UO_235 (O_235,N_7826,N_9591);
and UO_236 (O_236,N_9404,N_7707);
and UO_237 (O_237,N_7806,N_8948);
or UO_238 (O_238,N_8532,N_8936);
and UO_239 (O_239,N_9636,N_8986);
nor UO_240 (O_240,N_8793,N_7694);
and UO_241 (O_241,N_8383,N_7789);
nand UO_242 (O_242,N_9639,N_8584);
nor UO_243 (O_243,N_8435,N_8334);
nand UO_244 (O_244,N_7913,N_9816);
and UO_245 (O_245,N_7877,N_8715);
nand UO_246 (O_246,N_9845,N_7788);
and UO_247 (O_247,N_8717,N_7663);
nand UO_248 (O_248,N_7654,N_9462);
nor UO_249 (O_249,N_9869,N_9729);
and UO_250 (O_250,N_8890,N_7709);
nand UO_251 (O_251,N_7713,N_7976);
or UO_252 (O_252,N_7746,N_9181);
and UO_253 (O_253,N_9072,N_8293);
nor UO_254 (O_254,N_9521,N_8650);
nand UO_255 (O_255,N_8602,N_7838);
or UO_256 (O_256,N_9806,N_8231);
xor UO_257 (O_257,N_7626,N_8227);
nor UO_258 (O_258,N_8590,N_7901);
and UO_259 (O_259,N_7505,N_8145);
nand UO_260 (O_260,N_8870,N_8569);
or UO_261 (O_261,N_7535,N_9525);
nor UO_262 (O_262,N_9068,N_9145);
nand UO_263 (O_263,N_8084,N_9056);
nand UO_264 (O_264,N_8256,N_9945);
nor UO_265 (O_265,N_9495,N_7640);
and UO_266 (O_266,N_9858,N_9542);
and UO_267 (O_267,N_9526,N_9062);
nor UO_268 (O_268,N_8563,N_8765);
and UO_269 (O_269,N_9109,N_9270);
or UO_270 (O_270,N_9460,N_8363);
nor UO_271 (O_271,N_7760,N_9561);
xor UO_272 (O_272,N_8740,N_7576);
and UO_273 (O_273,N_8928,N_7608);
xor UO_274 (O_274,N_7904,N_9665);
and UO_275 (O_275,N_7975,N_9782);
xor UO_276 (O_276,N_8417,N_9819);
and UO_277 (O_277,N_8727,N_8109);
xor UO_278 (O_278,N_7961,N_8495);
nand UO_279 (O_279,N_9095,N_7889);
nand UO_280 (O_280,N_9865,N_8191);
nand UO_281 (O_281,N_9549,N_9700);
nor UO_282 (O_282,N_9527,N_9825);
or UO_283 (O_283,N_7884,N_9083);
nor UO_284 (O_284,N_8232,N_9560);
nor UO_285 (O_285,N_9609,N_9920);
nand UO_286 (O_286,N_9209,N_8083);
and UO_287 (O_287,N_9447,N_9361);
nor UO_288 (O_288,N_8184,N_8845);
nand UO_289 (O_289,N_7524,N_7578);
nand UO_290 (O_290,N_9138,N_9875);
or UO_291 (O_291,N_8434,N_9391);
nor UO_292 (O_292,N_8789,N_8708);
nor UO_293 (O_293,N_7983,N_8876);
and UO_294 (O_294,N_9709,N_9339);
nand UO_295 (O_295,N_9965,N_8931);
or UO_296 (O_296,N_7764,N_7822);
or UO_297 (O_297,N_9366,N_9407);
nand UO_298 (O_298,N_9237,N_9111);
or UO_299 (O_299,N_9890,N_7928);
nand UO_300 (O_300,N_9736,N_8244);
or UO_301 (O_301,N_9711,N_8196);
or UO_302 (O_302,N_9167,N_9398);
or UO_303 (O_303,N_9828,N_9386);
nor UO_304 (O_304,N_9505,N_7732);
nor UO_305 (O_305,N_7918,N_8030);
nand UO_306 (O_306,N_9277,N_9872);
nor UO_307 (O_307,N_9584,N_9103);
nor UO_308 (O_308,N_9264,N_7563);
and UO_309 (O_309,N_9180,N_9622);
nand UO_310 (O_310,N_7811,N_9269);
nand UO_311 (O_311,N_7900,N_8353);
or UO_312 (O_312,N_8841,N_7710);
and UO_313 (O_313,N_8093,N_8343);
and UO_314 (O_314,N_7926,N_9255);
xor UO_315 (O_315,N_9889,N_8370);
and UO_316 (O_316,N_9623,N_7896);
nor UO_317 (O_317,N_7646,N_7700);
xor UO_318 (O_318,N_9793,N_8056);
nor UO_319 (O_319,N_8183,N_8330);
and UO_320 (O_320,N_8889,N_7698);
or UO_321 (O_321,N_7890,N_7888);
or UO_322 (O_322,N_8368,N_9916);
nor UO_323 (O_323,N_9105,N_9844);
xor UO_324 (O_324,N_8658,N_7756);
nand UO_325 (O_325,N_9486,N_8090);
and UO_326 (O_326,N_9986,N_9030);
or UO_327 (O_327,N_8178,N_9240);
nor UO_328 (O_328,N_9154,N_8295);
or UO_329 (O_329,N_9210,N_8195);
xor UO_330 (O_330,N_9695,N_8139);
or UO_331 (O_331,N_8880,N_9212);
nand UO_332 (O_332,N_8573,N_8760);
xnor UO_333 (O_333,N_8672,N_9374);
xor UO_334 (O_334,N_9389,N_8698);
and UO_335 (O_335,N_9204,N_9250);
or UO_336 (O_336,N_8518,N_9394);
xnor UO_337 (O_337,N_7800,N_8069);
and UO_338 (O_338,N_8764,N_7946);
xnor UO_339 (O_339,N_8381,N_7666);
nor UO_340 (O_340,N_9805,N_9637);
or UO_341 (O_341,N_8176,N_7942);
nor UO_342 (O_342,N_9983,N_9863);
nand UO_343 (O_343,N_9740,N_9187);
and UO_344 (O_344,N_9188,N_8648);
nand UO_345 (O_345,N_8552,N_7785);
and UO_346 (O_346,N_8423,N_8979);
or UO_347 (O_347,N_9382,N_9870);
xnor UO_348 (O_348,N_9335,N_8787);
nor UO_349 (O_349,N_9576,N_7740);
nor UO_350 (O_350,N_9541,N_8998);
xnor UO_351 (O_351,N_8571,N_8456);
or UO_352 (O_352,N_8460,N_8375);
nand UO_353 (O_353,N_9972,N_7816);
nor UO_354 (O_354,N_8669,N_7723);
or UO_355 (O_355,N_8512,N_7967);
nand UO_356 (O_356,N_7726,N_7697);
nand UO_357 (O_357,N_7717,N_8018);
or UO_358 (O_358,N_8182,N_9756);
nor UO_359 (O_359,N_8772,N_9691);
and UO_360 (O_360,N_9812,N_8930);
or UO_361 (O_361,N_9029,N_8034);
or UO_362 (O_362,N_8861,N_8891);
nor UO_363 (O_363,N_8263,N_8678);
or UO_364 (O_364,N_9010,N_9424);
nand UO_365 (O_365,N_9184,N_7745);
and UO_366 (O_366,N_9384,N_9403);
nand UO_367 (O_367,N_9455,N_9586);
or UO_368 (O_368,N_8585,N_9321);
nor UO_369 (O_369,N_7728,N_9507);
nand UO_370 (O_370,N_7559,N_7915);
nand UO_371 (O_371,N_7973,N_7786);
or UO_372 (O_372,N_8049,N_9026);
or UO_373 (O_373,N_8143,N_9625);
and UO_374 (O_374,N_9895,N_8533);
nor UO_375 (O_375,N_9879,N_9059);
or UO_376 (O_376,N_9522,N_9780);
xor UO_377 (O_377,N_9461,N_9747);
nor UO_378 (O_378,N_9824,N_8797);
or UO_379 (O_379,N_8589,N_9820);
or UO_380 (O_380,N_8958,N_8007);
and UO_381 (O_381,N_9032,N_9412);
nand UO_382 (O_382,N_9799,N_9001);
and UO_383 (O_383,N_7882,N_7787);
xor UO_384 (O_384,N_8879,N_9659);
nor UO_385 (O_385,N_8318,N_7817);
nand UO_386 (O_386,N_7706,N_7548);
nor UO_387 (O_387,N_7534,N_8933);
nand UO_388 (O_388,N_9089,N_7631);
nor UO_389 (O_389,N_8031,N_7903);
nor UO_390 (O_390,N_8846,N_9048);
or UO_391 (O_391,N_9750,N_9833);
nor UO_392 (O_392,N_7949,N_8410);
nand UO_393 (O_393,N_8882,N_7652);
and UO_394 (O_394,N_9143,N_8442);
and UO_395 (O_395,N_9451,N_9717);
and UO_396 (O_396,N_9666,N_8272);
xnor UO_397 (O_397,N_7674,N_9420);
and UO_398 (O_398,N_8699,N_9647);
or UO_399 (O_399,N_8855,N_9065);
and UO_400 (O_400,N_9092,N_9147);
nand UO_401 (O_401,N_8530,N_8904);
or UO_402 (O_402,N_8515,N_7940);
xor UO_403 (O_403,N_7503,N_7599);
nand UO_404 (O_404,N_7546,N_9317);
nor UO_405 (O_405,N_9942,N_9004);
nor UO_406 (O_406,N_8886,N_7783);
nor UO_407 (O_407,N_9202,N_9332);
and UO_408 (O_408,N_7562,N_9668);
or UO_409 (O_409,N_7648,N_9843);
nor UO_410 (O_410,N_8355,N_7808);
nor UO_411 (O_411,N_9597,N_7615);
nand UO_412 (O_412,N_9632,N_8570);
nor UO_413 (O_413,N_8332,N_8624);
and UO_414 (O_414,N_9759,N_9114);
nand UO_415 (O_415,N_8130,N_9364);
nand UO_416 (O_416,N_7916,N_9300);
nor UO_417 (O_417,N_8337,N_8395);
nor UO_418 (O_418,N_9198,N_8972);
nand UO_419 (O_419,N_8099,N_9742);
nand UO_420 (O_420,N_8221,N_8469);
and UO_421 (O_421,N_7948,N_8391);
or UO_422 (O_422,N_8687,N_9352);
xnor UO_423 (O_423,N_8639,N_9342);
or UO_424 (O_424,N_8581,N_8742);
and UO_425 (O_425,N_7944,N_8308);
nand UO_426 (O_426,N_8778,N_9749);
or UO_427 (O_427,N_9490,N_8346);
nand UO_428 (O_428,N_7910,N_7938);
xnor UO_429 (O_429,N_9967,N_8135);
xnor UO_430 (O_430,N_8492,N_8398);
and UO_431 (O_431,N_8792,N_9422);
nor UO_432 (O_432,N_8695,N_7589);
xnor UO_433 (O_433,N_8265,N_9378);
nand UO_434 (O_434,N_9448,N_8534);
and UO_435 (O_435,N_7545,N_7775);
nand UO_436 (O_436,N_9993,N_7970);
nand UO_437 (O_437,N_9605,N_7659);
and UO_438 (O_438,N_8691,N_9672);
nand UO_439 (O_439,N_8147,N_9493);
or UO_440 (O_440,N_9826,N_8039);
and UO_441 (O_441,N_7858,N_8329);
and UO_442 (O_442,N_8239,N_7823);
or UO_443 (O_443,N_9081,N_8701);
and UO_444 (O_444,N_7529,N_7751);
nor UO_445 (O_445,N_7643,N_9368);
or UO_446 (O_446,N_8961,N_8489);
nor UO_447 (O_447,N_7598,N_8378);
nand UO_448 (O_448,N_9107,N_8951);
or UO_449 (O_449,N_9973,N_8974);
and UO_450 (O_450,N_8888,N_8322);
nor UO_451 (O_451,N_9648,N_8503);
nand UO_452 (O_452,N_9406,N_9904);
and UO_453 (O_453,N_7813,N_9100);
or UO_454 (O_454,N_7835,N_7594);
nor UO_455 (O_455,N_7647,N_7687);
nor UO_456 (O_456,N_9599,N_7930);
or UO_457 (O_457,N_7602,N_9530);
nor UO_458 (O_458,N_9612,N_8738);
or UO_459 (O_459,N_9483,N_9638);
and UO_460 (O_460,N_8967,N_7951);
and UO_461 (O_461,N_7833,N_8731);
nand UO_462 (O_462,N_7829,N_8040);
nand UO_463 (O_463,N_8721,N_7588);
nand UO_464 (O_464,N_8806,N_8213);
nand UO_465 (O_465,N_8499,N_8336);
and UO_466 (O_466,N_8214,N_9126);
nand UO_467 (O_467,N_9311,N_9185);
or UO_468 (O_468,N_9208,N_8242);
or UO_469 (O_469,N_9223,N_8686);
nor UO_470 (O_470,N_9797,N_8781);
or UO_471 (O_471,N_8664,N_7798);
nor UO_472 (O_472,N_8900,N_8666);
nor UO_473 (O_473,N_9016,N_8487);
or UO_474 (O_474,N_7575,N_9298);
and UO_475 (O_475,N_8860,N_9504);
nor UO_476 (O_476,N_9969,N_9757);
nand UO_477 (O_477,N_7614,N_9466);
and UO_478 (O_478,N_8826,N_8907);
nand UO_479 (O_479,N_8878,N_8316);
xnor UO_480 (O_480,N_8511,N_9957);
nand UO_481 (O_481,N_8615,N_9159);
and UO_482 (O_482,N_9033,N_8980);
or UO_483 (O_483,N_9047,N_8477);
and UO_484 (O_484,N_9738,N_9959);
nor UO_485 (O_485,N_8535,N_9009);
xor UO_486 (O_486,N_7931,N_8827);
xnor UO_487 (O_487,N_7560,N_9146);
nor UO_488 (O_488,N_7762,N_9482);
or UO_489 (O_489,N_9762,N_8582);
xnor UO_490 (O_490,N_8874,N_8541);
nor UO_491 (O_491,N_9020,N_9273);
nor UO_492 (O_492,N_8126,N_7872);
nor UO_493 (O_493,N_8558,N_9894);
and UO_494 (O_494,N_9537,N_9211);
nor UO_495 (O_495,N_8935,N_8394);
and UO_496 (O_496,N_8342,N_9110);
nor UO_497 (O_497,N_7761,N_8683);
nand UO_498 (O_498,N_7739,N_8360);
and UO_499 (O_499,N_9294,N_8086);
xor UO_500 (O_500,N_7714,N_9562);
or UO_501 (O_501,N_8038,N_9494);
nand UO_502 (O_502,N_9671,N_7702);
and UO_503 (O_503,N_9553,N_7543);
xnor UO_504 (O_504,N_9268,N_8508);
nand UO_505 (O_505,N_7556,N_8836);
or UO_506 (O_506,N_8357,N_7644);
and UO_507 (O_507,N_8579,N_9550);
and UO_508 (O_508,N_7573,N_8548);
nand UO_509 (O_509,N_7625,N_8068);
and UO_510 (O_510,N_8916,N_7971);
nor UO_511 (O_511,N_8591,N_7849);
and UO_512 (O_512,N_7770,N_9928);
nand UO_513 (O_513,N_9903,N_8163);
or UO_514 (O_514,N_8975,N_7879);
and UO_515 (O_515,N_9628,N_7636);
and UO_516 (O_516,N_8438,N_8537);
nand UO_517 (O_517,N_9644,N_9664);
nand UO_518 (O_518,N_9139,N_7987);
or UO_519 (O_519,N_9405,N_8519);
and UO_520 (O_520,N_7891,N_9934);
xnor UO_521 (O_521,N_9856,N_8015);
xor UO_522 (O_522,N_9247,N_8407);
or UO_523 (O_523,N_8920,N_8790);
nor UO_524 (O_524,N_9613,N_8386);
nor UO_525 (O_525,N_8199,N_8266);
xnor UO_526 (O_526,N_8501,N_7920);
and UO_527 (O_527,N_8801,N_9120);
nand UO_528 (O_528,N_7856,N_9733);
nor UO_529 (O_529,N_7839,N_8441);
and UO_530 (O_530,N_8364,N_9262);
nand UO_531 (O_531,N_7551,N_8505);
and UO_532 (O_532,N_7773,N_9252);
nand UO_533 (O_533,N_7742,N_8770);
or UO_534 (O_534,N_9685,N_8884);
nor UO_535 (O_535,N_8758,N_8496);
and UO_536 (O_536,N_9218,N_9554);
nor UO_537 (O_537,N_9283,N_8919);
or UO_538 (O_538,N_8264,N_8310);
nor UO_539 (O_539,N_9968,N_9429);
and UO_540 (O_540,N_9328,N_8660);
nor UO_541 (O_541,N_8001,N_7885);
and UO_542 (O_542,N_8864,N_8236);
and UO_543 (O_543,N_8984,N_7606);
xor UO_544 (O_544,N_8023,N_7985);
nor UO_545 (O_545,N_7689,N_8367);
and UO_546 (O_546,N_9795,N_8757);
nand UO_547 (O_547,N_7862,N_8248);
nand UO_548 (O_548,N_9621,N_8566);
or UO_549 (O_549,N_8934,N_9164);
or UO_550 (O_550,N_9446,N_7569);
nand UO_551 (O_551,N_8700,N_9191);
nand UO_552 (O_552,N_8158,N_7679);
and UO_553 (O_553,N_9327,N_7905);
nor UO_554 (O_554,N_9487,N_8003);
xor UO_555 (O_555,N_8539,N_8670);
and UO_556 (O_556,N_7617,N_8223);
or UO_557 (O_557,N_8808,N_9318);
and UO_558 (O_558,N_9763,N_8230);
and UO_559 (O_559,N_9979,N_8583);
nand UO_560 (O_560,N_7669,N_9516);
nand UO_561 (O_561,N_9108,N_8523);
nand UO_562 (O_562,N_7945,N_8149);
nand UO_563 (O_563,N_9469,N_7960);
nor UO_564 (O_564,N_9985,N_9594);
nor UO_565 (O_565,N_9492,N_9285);
and UO_566 (O_566,N_8224,N_7957);
or UO_567 (O_567,N_9383,N_9031);
and UO_568 (O_568,N_9834,N_7724);
nand UO_569 (O_569,N_9090,N_8022);
or UO_570 (O_570,N_8047,N_8782);
or UO_571 (O_571,N_7857,N_9282);
or UO_572 (O_572,N_9614,N_8371);
nand UO_573 (O_573,N_8743,N_9690);
nand UO_574 (O_574,N_9074,N_7555);
nor UO_575 (O_575,N_7914,N_8866);
nand UO_576 (O_576,N_8104,N_8361);
and UO_577 (O_577,N_9924,N_9773);
and UO_578 (O_578,N_9099,N_7749);
nor UO_579 (O_579,N_7662,N_9227);
nor UO_580 (O_580,N_9197,N_8954);
nand UO_581 (O_581,N_9194,N_9997);
xnor UO_582 (O_582,N_9682,N_7867);
nand UO_583 (O_583,N_9104,N_8502);
xnor UO_584 (O_584,N_8171,N_9011);
xor UO_585 (O_585,N_8956,N_9307);
and UO_586 (O_586,N_8720,N_7853);
xor UO_587 (O_587,N_8945,N_9434);
xnor UO_588 (O_588,N_7716,N_7979);
nand UO_589 (O_589,N_7512,N_9939);
and UO_590 (O_590,N_9256,N_8798);
or UO_591 (O_591,N_9474,N_8249);
nor UO_592 (O_592,N_8162,N_9966);
nor UO_593 (O_593,N_8647,N_7660);
and UO_594 (O_594,N_9150,N_9192);
xor UO_595 (O_595,N_9041,N_9910);
and UO_596 (O_596,N_8396,N_9669);
and UO_597 (O_597,N_9633,N_8245);
or UO_598 (O_598,N_9748,N_9761);
or UO_599 (O_599,N_9220,N_8013);
nand UO_600 (O_600,N_9216,N_8217);
and UO_601 (O_601,N_8795,N_9754);
or UO_602 (O_602,N_8966,N_8218);
and UO_603 (O_603,N_8906,N_8235);
nor UO_604 (O_604,N_8603,N_8121);
and UO_605 (O_605,N_8468,N_8830);
nand UO_606 (O_606,N_8807,N_9119);
or UO_607 (O_607,N_9358,N_9477);
or UO_608 (O_608,N_9322,N_8320);
xor UO_609 (O_609,N_7776,N_8105);
or UO_610 (O_610,N_9233,N_8210);
nor UO_611 (O_611,N_9809,N_9877);
and UO_612 (O_612,N_8475,N_8902);
nand UO_613 (O_613,N_9417,N_7922);
and UO_614 (O_614,N_8863,N_7923);
and UO_615 (O_615,N_7995,N_8262);
nor UO_616 (O_616,N_8118,N_9651);
nand UO_617 (O_617,N_8746,N_8498);
nor UO_618 (O_618,N_9859,N_8829);
nand UO_619 (O_619,N_8208,N_9848);
nand UO_620 (O_620,N_9258,N_7766);
or UO_621 (O_621,N_8311,N_9304);
and UO_622 (O_622,N_8029,N_8278);
nand UO_623 (O_623,N_8681,N_8390);
nor UO_624 (O_624,N_9244,N_7730);
or UO_625 (O_625,N_9688,N_8280);
nor UO_626 (O_626,N_9236,N_9978);
nand UO_627 (O_627,N_9926,N_9603);
and UO_628 (O_628,N_8839,N_8750);
or UO_629 (O_629,N_8674,N_8180);
nor UO_630 (O_630,N_8823,N_7664);
and UO_631 (O_631,N_8255,N_7828);
nand UO_632 (O_632,N_8847,N_8042);
nor UO_633 (O_633,N_8509,N_9911);
or UO_634 (O_634,N_8127,N_9932);
nor UO_635 (O_635,N_7863,N_8252);
or UO_636 (O_636,N_9195,N_9178);
and UO_637 (O_637,N_8315,N_9450);
nand UO_638 (O_638,N_8169,N_9345);
nand UO_639 (O_639,N_8325,N_7586);
nand UO_640 (O_640,N_9515,N_7919);
nand UO_641 (O_641,N_9852,N_8822);
nand UO_642 (O_642,N_8455,N_7670);
or UO_643 (O_643,N_8997,N_8291);
nand UO_644 (O_644,N_9743,N_9496);
and UO_645 (O_645,N_9896,N_9771);
nand UO_646 (O_646,N_8576,N_9012);
xnor UO_647 (O_647,N_8922,N_8004);
nand UO_648 (O_648,N_9954,N_9755);
or UO_649 (O_649,N_9900,N_9087);
and UO_650 (O_650,N_9049,N_8285);
nor UO_651 (O_651,N_9886,N_9369);
or UO_652 (O_652,N_7784,N_8243);
xor UO_653 (O_653,N_8212,N_7777);
nand UO_654 (O_654,N_8759,N_9421);
nand UO_655 (O_655,N_9831,N_8755);
nor UO_656 (O_656,N_9347,N_8497);
or UO_657 (O_657,N_8734,N_7703);
or UO_658 (O_658,N_9963,N_8059);
nor UO_659 (O_659,N_8062,N_9249);
nand UO_660 (O_660,N_8439,N_7720);
or UO_661 (O_661,N_8414,N_9946);
nor UO_662 (O_662,N_9053,N_8815);
nor UO_663 (O_663,N_8206,N_9604);
nor UO_664 (O_664,N_9241,N_8655);
or UO_665 (O_665,N_8854,N_8522);
nor UO_666 (O_666,N_9779,N_7846);
or UO_667 (O_667,N_7731,N_8604);
nor UO_668 (O_668,N_9214,N_7880);
or UO_669 (O_669,N_8055,N_8587);
nor UO_670 (O_670,N_9316,N_8376);
or UO_671 (O_671,N_9535,N_9280);
or UO_672 (O_672,N_8521,N_9909);
nor UO_673 (O_673,N_8373,N_9097);
xor UO_674 (O_674,N_9991,N_7515);
or UO_675 (O_675,N_8491,N_9064);
and UO_676 (O_676,N_8131,N_9257);
and UO_677 (O_677,N_9642,N_9042);
xor UO_678 (O_678,N_7583,N_9815);
and UO_679 (O_679,N_8510,N_8723);
or UO_680 (O_680,N_9287,N_9881);
nand UO_681 (O_681,N_9837,N_8129);
nand UO_682 (O_682,N_8304,N_9035);
nand UO_683 (O_683,N_7804,N_8800);
nand UO_684 (O_684,N_8197,N_9598);
nor UO_685 (O_685,N_8791,N_9428);
nand UO_686 (O_686,N_8722,N_8554);
nor UO_687 (O_687,N_7993,N_7591);
and UO_688 (O_688,N_9162,N_8616);
or UO_689 (O_689,N_9007,N_9433);
and UO_690 (O_690,N_9445,N_8673);
nor UO_691 (O_691,N_7570,N_7516);
nand UO_692 (O_692,N_7712,N_7754);
nand UO_693 (O_693,N_7997,N_8464);
xor UO_694 (O_694,N_9086,N_7763);
nor UO_695 (O_695,N_7768,N_9673);
nor UO_696 (O_696,N_9245,N_8944);
or UO_697 (O_697,N_9944,N_8133);
and UO_698 (O_698,N_8526,N_7552);
and UO_699 (O_699,N_8092,N_9789);
or UO_700 (O_700,N_9579,N_8011);
xnor UO_701 (O_701,N_8517,N_8065);
nor UO_702 (O_702,N_9400,N_9459);
nor UO_703 (O_703,N_8070,N_9992);
nand UO_704 (O_704,N_8110,N_7758);
nand UO_705 (O_705,N_8651,N_7959);
and UO_706 (O_706,N_7937,N_7619);
and UO_707 (O_707,N_9974,N_8014);
nand UO_708 (O_708,N_7851,N_9375);
or UO_709 (O_709,N_8564,N_8817);
and UO_710 (O_710,N_7733,N_9416);
or UO_711 (O_711,N_7767,N_9066);
nor UO_712 (O_712,N_8459,N_8598);
and UO_713 (O_713,N_9772,N_9157);
xor UO_714 (O_714,N_8393,N_9657);
or UO_715 (O_715,N_8340,N_7677);
and UO_716 (O_716,N_8556,N_9617);
nor UO_717 (O_717,N_9893,N_7927);
and UO_718 (O_718,N_8111,N_9626);
and UO_719 (O_719,N_8588,N_9808);
nor UO_720 (O_720,N_8372,N_7820);
and UO_721 (O_721,N_7604,N_8643);
or UO_722 (O_722,N_8578,N_8205);
nor UO_723 (O_723,N_9082,N_8811);
and UO_724 (O_724,N_8779,N_9585);
nand UO_725 (O_725,N_8190,N_8705);
nor UO_726 (O_726,N_9545,N_8679);
nor UO_727 (O_727,N_9018,N_8805);
nand UO_728 (O_728,N_7554,N_8382);
nor UO_729 (O_729,N_9324,N_9117);
or UO_730 (O_730,N_7613,N_7909);
nand UO_731 (O_731,N_7607,N_8445);
nand UO_732 (O_732,N_9166,N_7541);
xor UO_733 (O_733,N_9452,N_7964);
or UO_734 (O_734,N_8257,N_8619);
nand UO_735 (O_735,N_8659,N_7935);
nor UO_736 (O_736,N_7912,N_8909);
nand UO_737 (O_737,N_9880,N_9753);
and UO_738 (O_738,N_8021,N_9123);
xor UO_739 (O_739,N_9601,N_9000);
xnor UO_740 (O_740,N_9340,N_9096);
or UO_741 (O_741,N_9866,N_8962);
nor UO_742 (O_742,N_8677,N_9265);
nor UO_743 (O_743,N_8054,N_9832);
nor UO_744 (O_744,N_8551,N_9286);
xnor UO_745 (O_745,N_9140,N_9670);
xor UO_746 (O_746,N_7779,N_8702);
or UO_747 (O_747,N_8247,N_9025);
nand UO_748 (O_748,N_7704,N_9497);
and UO_749 (O_749,N_9829,N_9575);
nand UO_750 (O_750,N_8988,N_8165);
and UO_751 (O_751,N_9266,N_9692);
nand UO_752 (O_752,N_8254,N_7845);
nand UO_753 (O_753,N_9439,N_7574);
or UO_754 (O_754,N_7895,N_8098);
or UO_755 (O_755,N_8773,N_8623);
and UO_756 (O_756,N_8220,N_9137);
nand UO_757 (O_757,N_8451,N_8494);
and UO_758 (O_758,N_9465,N_8842);
or UO_759 (O_759,N_9410,N_8010);
or UO_760 (O_760,N_9392,N_8348);
nand UO_761 (O_761,N_8493,N_7605);
and UO_762 (O_762,N_8148,N_8351);
nor UO_763 (O_763,N_9645,N_7842);
and UO_764 (O_764,N_9267,N_9372);
nor UO_765 (O_765,N_8991,N_7671);
and UO_766 (O_766,N_9234,N_9365);
nor UO_767 (O_767,N_9660,N_7854);
xnor UO_768 (O_768,N_9499,N_9817);
nand UO_769 (O_769,N_9116,N_8138);
or UO_770 (O_770,N_9349,N_9411);
or UO_771 (O_771,N_9179,N_9699);
and UO_772 (O_772,N_9519,N_8222);
or UO_773 (O_773,N_9271,N_8216);
nand UO_774 (O_774,N_8446,N_8035);
or UO_775 (O_775,N_8976,N_7550);
or UO_776 (O_776,N_8887,N_8981);
nand UO_777 (O_777,N_9408,N_9457);
and UO_778 (O_778,N_9122,N_9876);
nand UO_779 (O_779,N_9898,N_8858);
and UO_780 (O_780,N_8379,N_8443);
or UO_781 (O_781,N_7852,N_9057);
or UO_782 (O_782,N_9891,N_8690);
nand UO_783 (O_783,N_9228,N_9792);
or UO_784 (O_784,N_8549,N_8421);
or UO_785 (O_785,N_8654,N_9291);
or UO_786 (O_786,N_9938,N_8622);
and UO_787 (O_787,N_8575,N_8985);
nor UO_788 (O_788,N_8174,N_8472);
nand UO_789 (O_789,N_8437,N_8610);
or UO_790 (O_790,N_8867,N_8063);
nor UO_791 (O_791,N_8354,N_8474);
nor UO_792 (O_792,N_8200,N_8338);
and UO_793 (O_793,N_8323,N_8281);
and UO_794 (O_794,N_8728,N_8630);
nand UO_795 (O_795,N_9802,N_9551);
or UO_796 (O_796,N_8775,N_9073);
nor UO_797 (O_797,N_7860,N_8949);
nand UO_798 (O_798,N_9232,N_8625);
nand UO_799 (O_799,N_9683,N_9901);
and UO_800 (O_800,N_8073,N_8568);
xnor UO_801 (O_801,N_8749,N_8642);
nand UO_802 (O_802,N_9259,N_8771);
nor UO_803 (O_803,N_7683,N_9606);
and UO_804 (O_804,N_8953,N_9847);
nor UO_805 (O_805,N_9235,N_7678);
xor UO_806 (O_806,N_9229,N_8736);
or UO_807 (O_807,N_8349,N_9905);
nor UO_808 (O_808,N_7899,N_8017);
or UO_809 (O_809,N_9777,N_7892);
or UO_810 (O_810,N_9552,N_7834);
and UO_811 (O_811,N_9658,N_8120);
or UO_812 (O_812,N_9051,N_9913);
nor UO_813 (O_813,N_9193,N_8557);
and UO_814 (O_814,N_8794,N_8405);
or UO_815 (O_815,N_7861,N_9468);
or UO_816 (O_816,N_8724,N_8268);
and UO_817 (O_817,N_9888,N_8853);
or UO_818 (O_818,N_9131,N_8168);
xor UO_819 (O_819,N_7797,N_8119);
and UO_820 (O_820,N_9862,N_7906);
nand UO_821 (O_821,N_8618,N_9919);
nand UO_822 (O_822,N_8317,N_7859);
and UO_823 (O_823,N_9760,N_7553);
and UO_824 (O_824,N_8436,N_9050);
xor UO_825 (O_825,N_7539,N_8668);
nand UO_826 (O_826,N_9315,N_8812);
nand UO_827 (O_827,N_7721,N_9811);
xnor UO_828 (O_828,N_8006,N_9506);
and UO_829 (O_829,N_9360,N_8461);
nand UO_830 (O_830,N_9356,N_7540);
nor UO_831 (O_831,N_8306,N_8810);
or UO_832 (O_832,N_8307,N_8753);
and UO_833 (O_833,N_9678,N_9101);
nor UO_834 (O_834,N_8319,N_8671);
or UO_835 (O_835,N_8628,N_9440);
nand UO_836 (O_836,N_8326,N_8172);
xor UO_837 (O_837,N_9153,N_9744);
nor UO_838 (O_838,N_8312,N_8115);
nand UO_839 (O_839,N_9653,N_9708);
or UO_840 (O_840,N_9453,N_8440);
xnor UO_841 (O_841,N_9238,N_7795);
nor UO_842 (O_842,N_8484,N_9503);
or UO_843 (O_843,N_8943,N_9205);
nand UO_844 (O_844,N_9170,N_7544);
and UO_845 (O_845,N_9783,N_9854);
or UO_846 (O_846,N_8915,N_7685);
and UO_847 (O_847,N_9964,N_9135);
or UO_848 (O_848,N_7627,N_8929);
or UO_849 (O_849,N_8730,N_9423);
nor UO_850 (O_850,N_9002,N_9106);
xor UO_851 (O_851,N_9226,N_9289);
and UO_852 (O_852,N_8211,N_8203);
and UO_853 (O_853,N_9588,N_9727);
nor UO_854 (O_854,N_8849,N_9501);
and UO_855 (O_855,N_9488,N_9830);
xnor UO_856 (O_856,N_9470,N_9359);
or UO_857 (O_857,N_8586,N_8362);
nor UO_858 (O_858,N_9803,N_8665);
nand UO_859 (O_859,N_9142,N_8296);
nand UO_860 (O_860,N_9034,N_7809);
xor UO_861 (O_861,N_8128,N_9409);
nor UO_862 (O_862,N_7936,N_9189);
nor UO_863 (O_863,N_7727,N_7792);
or UO_864 (O_864,N_9573,N_9348);
and UO_865 (O_865,N_8875,N_8620);
xor UO_866 (O_866,N_9160,N_8711);
and UO_867 (O_867,N_8652,N_8450);
and UO_868 (O_868,N_8186,N_7722);
xor UO_869 (O_869,N_8617,N_8637);
nor UO_870 (O_870,N_8033,N_8629);
nand UO_871 (O_871,N_8607,N_9132);
nor UO_872 (O_872,N_7847,N_9712);
xnor UO_873 (O_873,N_9512,N_7667);
nor UO_874 (O_874,N_7805,N_9312);
or UO_875 (O_875,N_9915,N_7610);
xor UO_876 (O_876,N_8766,N_7514);
xor UO_877 (O_877,N_8080,N_7632);
or UO_878 (O_878,N_9314,N_9155);
and UO_879 (O_879,N_8384,N_9885);
nand UO_880 (O_880,N_9067,N_9618);
and UO_881 (O_881,N_8994,N_9914);
nand UO_882 (O_882,N_9528,N_9112);
or UO_883 (O_883,N_8977,N_8114);
nand UO_884 (O_884,N_9251,N_8444);
or UO_885 (O_885,N_9331,N_8389);
nand UO_886 (O_886,N_7897,N_9882);
nand UO_887 (O_887,N_9206,N_9663);
or UO_888 (O_888,N_7566,N_8100);
or UO_889 (O_889,N_7876,N_7582);
nor UO_890 (O_890,N_7950,N_7782);
nor UO_891 (O_891,N_9338,N_7966);
nand UO_892 (O_892,N_8071,N_8500);
and UO_893 (O_893,N_7511,N_8356);
nand UO_894 (O_894,N_8177,N_8411);
and UO_895 (O_895,N_7925,N_8366);
nor UO_896 (O_896,N_8228,N_9710);
nand UO_897 (O_897,N_9616,N_7921);
or UO_898 (O_898,N_8170,N_9498);
xnor UO_899 (O_899,N_8202,N_7661);
nor UO_900 (O_900,N_9581,N_8292);
or UO_901 (O_901,N_8744,N_8036);
nand UO_902 (O_902,N_9596,N_8002);
or UO_903 (O_903,N_7507,N_9078);
nor UO_904 (O_904,N_9838,N_9577);
or UO_905 (O_905,N_9351,N_7866);
nand UO_906 (O_906,N_8289,N_8290);
nor UO_907 (O_907,N_9302,N_9373);
nor UO_908 (O_908,N_7999,N_8462);
nand UO_909 (O_909,N_9133,N_8448);
and UO_910 (O_910,N_9960,N_7841);
or UO_911 (O_911,N_9861,N_7609);
and UO_912 (O_912,N_9846,N_8820);
nand UO_913 (O_913,N_8385,N_8101);
nand UO_914 (O_914,N_7832,N_8761);
or UO_915 (O_915,N_9454,N_8091);
nand UO_916 (O_916,N_8286,N_8005);
and UO_917 (O_917,N_8881,N_9990);
nor UO_918 (O_918,N_9529,N_9043);
xor UO_919 (O_919,N_8078,N_9652);
xor UO_920 (O_920,N_9098,N_8692);
nand UO_921 (O_921,N_9608,N_8044);
or UO_922 (O_922,N_7519,N_9770);
xor UO_923 (O_923,N_9055,N_8856);
xnor UO_924 (O_924,N_8970,N_9438);
nor UO_925 (O_925,N_8053,N_8543);
and UO_926 (O_926,N_8641,N_7771);
or UO_927 (O_927,N_8877,N_9627);
or UO_928 (O_928,N_8146,N_9857);
or UO_929 (O_929,N_9610,N_8848);
nand UO_930 (O_930,N_8525,N_9546);
and UO_931 (O_931,N_8488,N_9186);
nand UO_932 (O_932,N_9781,N_9566);
xor UO_933 (O_933,N_8597,N_8274);
or UO_934 (O_934,N_7994,N_9239);
and UO_935 (O_935,N_8194,N_8250);
nor UO_936 (O_936,N_9836,N_7525);
and UO_937 (O_937,N_7579,N_9706);
and UO_938 (O_938,N_8754,N_9533);
nand UO_939 (O_939,N_9491,N_8238);
or UO_940 (O_940,N_7595,N_9344);
and UO_941 (O_941,N_8667,N_7673);
xnor UO_942 (O_942,N_9508,N_8132);
or UO_943 (O_943,N_8741,N_8134);
nor UO_944 (O_944,N_9798,N_9019);
nor UO_945 (O_945,N_9936,N_8905);
nor UO_946 (O_946,N_8627,N_8234);
nor UO_947 (O_947,N_7587,N_8696);
nor UO_948 (O_948,N_9456,N_8074);
nor UO_949 (O_949,N_9325,N_8946);
and UO_950 (O_950,N_8895,N_9243);
and UO_951 (O_951,N_9721,N_8726);
xor UO_952 (O_952,N_9860,N_9141);
or UO_953 (O_953,N_7680,N_9958);
xnor UO_954 (O_954,N_9667,N_8776);
and UO_955 (O_955,N_9583,N_8952);
and UO_956 (O_956,N_9006,N_9791);
nand UO_957 (O_957,N_8045,N_9735);
or UO_958 (O_958,N_7803,N_8862);
or UO_959 (O_959,N_9355,N_9684);
and UO_960 (O_960,N_8685,N_9589);
or UO_961 (O_961,N_8479,N_8662);
nor UO_962 (O_962,N_9295,N_8303);
nor UO_963 (O_963,N_7655,N_7953);
nor UO_964 (O_964,N_7998,N_8661);
and UO_965 (O_965,N_7887,N_8251);
or UO_966 (O_966,N_7992,N_9557);
or UO_967 (O_967,N_7597,N_9774);
and UO_968 (O_968,N_8215,N_8112);
nor UO_969 (O_969,N_9514,N_9800);
nand UO_970 (O_970,N_8279,N_8141);
or UO_971 (O_971,N_9130,N_9868);
xor UO_972 (O_972,N_8124,N_9723);
or UO_973 (O_973,N_9148,N_9272);
or UO_974 (O_974,N_8704,N_8542);
nand UO_975 (O_975,N_8117,N_9058);
and UO_976 (O_976,N_9134,N_7639);
nor UO_977 (O_977,N_8865,N_8225);
nor UO_978 (O_978,N_7601,N_9532);
nor UO_979 (O_979,N_8369,N_7908);
or UO_980 (O_980,N_8028,N_8009);
or UO_981 (O_981,N_9943,N_8990);
nand UO_982 (O_982,N_8433,N_9764);
xnor UO_983 (O_983,N_9079,N_9855);
xnor UO_984 (O_984,N_8480,N_7523);
nand UO_985 (O_985,N_7637,N_7969);
nand UO_986 (O_986,N_9163,N_9161);
nand UO_987 (O_987,N_9615,N_8712);
nand UO_988 (O_988,N_9323,N_9714);
nand UO_989 (O_989,N_8957,N_9786);
nand UO_990 (O_990,N_9397,N_9149);
or UO_991 (O_991,N_7821,N_8783);
nand UO_992 (O_992,N_7810,N_9853);
nor UO_993 (O_993,N_7881,N_8187);
and UO_994 (O_994,N_8763,N_9935);
nor UO_995 (O_995,N_9813,N_9121);
nor UO_996 (O_996,N_9254,N_8646);
xor UO_997 (O_997,N_8595,N_7812);
nand UO_998 (O_998,N_7641,N_7621);
or UO_999 (O_999,N_9085,N_9341);
nor UO_1000 (O_1000,N_8613,N_8684);
nand UO_1001 (O_1001,N_8299,N_8465);
or UO_1002 (O_1002,N_8324,N_9022);
or UO_1003 (O_1003,N_7963,N_8894);
nand UO_1004 (O_1004,N_8871,N_8399);
and UO_1005 (O_1005,N_8788,N_9381);
or UO_1006 (O_1006,N_9158,N_8640);
xnor UO_1007 (O_1007,N_8816,N_9380);
nand UO_1008 (O_1008,N_9357,N_8828);
nand UO_1009 (O_1009,N_8803,N_9734);
xor UO_1010 (O_1010,N_8156,N_9788);
xnor UO_1011 (O_1011,N_8328,N_8982);
nand UO_1012 (O_1012,N_8645,N_9981);
and UO_1013 (O_1013,N_9172,N_8490);
nand UO_1014 (O_1014,N_8706,N_9570);
nor UO_1015 (O_1015,N_8592,N_8676);
nand UO_1016 (O_1016,N_8555,N_8868);
xnor UO_1017 (O_1017,N_7943,N_9481);
nand UO_1018 (O_1018,N_9962,N_9580);
nor UO_1019 (O_1019,N_7510,N_8198);
or UO_1020 (O_1020,N_7526,N_9279);
and UO_1021 (O_1021,N_8103,N_8425);
nand UO_1022 (O_1022,N_9704,N_7824);
nor UO_1023 (O_1023,N_9230,N_8380);
nor UO_1024 (O_1024,N_9607,N_8777);
nand UO_1025 (O_1025,N_7531,N_9284);
nor UO_1026 (O_1026,N_9502,N_9297);
xor UO_1027 (O_1027,N_9765,N_9674);
and UO_1028 (O_1028,N_9982,N_9313);
and UO_1029 (O_1029,N_7537,N_9999);
and UO_1030 (O_1030,N_9080,N_8458);
and UO_1031 (O_1031,N_8634,N_8155);
nand UO_1032 (O_1032,N_8547,N_7958);
nand UO_1033 (O_1033,N_8747,N_7513);
and UO_1034 (O_1034,N_7850,N_9654);
nand UO_1035 (O_1035,N_9931,N_9224);
and UO_1036 (O_1036,N_9500,N_7642);
and UO_1037 (O_1037,N_9346,N_7796);
and UO_1038 (O_1038,N_7600,N_8400);
nand UO_1039 (O_1039,N_8925,N_8594);
nor UO_1040 (O_1040,N_9040,N_8514);
nor UO_1041 (O_1041,N_7837,N_7772);
or UO_1042 (O_1042,N_8901,N_7759);
nand UO_1043 (O_1043,N_9646,N_9248);
or UO_1044 (O_1044,N_9996,N_7634);
and UO_1045 (O_1045,N_7509,N_7668);
and UO_1046 (O_1046,N_9069,N_9008);
nor UO_1047 (O_1047,N_8066,N_9768);
nor UO_1048 (O_1048,N_8993,N_9175);
xnor UO_1049 (O_1049,N_8226,N_7952);
and UO_1050 (O_1050,N_8918,N_8546);
or UO_1051 (O_1051,N_8601,N_7902);
and UO_1052 (O_1052,N_8253,N_7801);
nand UO_1053 (O_1053,N_8910,N_8164);
or UO_1054 (O_1054,N_7651,N_9418);
nand UO_1055 (O_1055,N_9091,N_8457);
nor UO_1056 (O_1056,N_8270,N_9038);
or UO_1057 (O_1057,N_7628,N_9296);
nor UO_1058 (O_1058,N_7665,N_8821);
and UO_1059 (O_1059,N_7933,N_8714);
nand UO_1060 (O_1060,N_8008,N_7506);
and UO_1061 (O_1061,N_9961,N_7658);
and UO_1062 (O_1062,N_9899,N_8965);
or UO_1063 (O_1063,N_9794,N_7836);
or UO_1064 (O_1064,N_9650,N_8157);
nor UO_1065 (O_1065,N_8282,N_8108);
nor UO_1066 (O_1066,N_7734,N_9183);
or UO_1067 (O_1067,N_7520,N_8052);
nor UO_1068 (O_1068,N_9425,N_9543);
xor UO_1069 (O_1069,N_8697,N_9017);
and UO_1070 (O_1070,N_7911,N_7584);
or UO_1071 (O_1071,N_8507,N_7855);
nor UO_1072 (O_1072,N_9084,N_8452);
and UO_1073 (O_1073,N_7675,N_9582);
nand UO_1074 (O_1074,N_8911,N_9426);
or UO_1075 (O_1075,N_7549,N_7954);
nor UO_1076 (O_1076,N_8471,N_8397);
nor UO_1077 (O_1077,N_9190,N_9849);
and UO_1078 (O_1078,N_8840,N_7501);
or UO_1079 (O_1079,N_7871,N_8892);
nor UO_1080 (O_1080,N_8611,N_8152);
nand UO_1081 (O_1081,N_8067,N_7715);
or UO_1082 (O_1082,N_9988,N_9061);
nand UO_1083 (O_1083,N_9821,N_8814);
and UO_1084 (O_1084,N_7708,N_8159);
nor UO_1085 (O_1085,N_9722,N_7799);
nand UO_1086 (O_1086,N_8735,N_9437);
nor UO_1087 (O_1087,N_9509,N_9952);
nand UO_1088 (O_1088,N_8478,N_8818);
nor UO_1089 (O_1089,N_7807,N_9745);
nand UO_1090 (O_1090,N_8649,N_7699);
or UO_1091 (O_1091,N_8192,N_9818);
nand UO_1092 (O_1092,N_7865,N_9698);
nand UO_1093 (O_1093,N_7750,N_9219);
nor UO_1094 (O_1094,N_9814,N_7638);
and UO_1095 (O_1095,N_9329,N_8277);
xor UO_1096 (O_1096,N_8926,N_9395);
nand UO_1097 (O_1097,N_9702,N_8408);
nand UO_1098 (O_1098,N_8032,N_8596);
or UO_1099 (O_1099,N_7778,N_8166);
nand UO_1100 (O_1100,N_9643,N_7869);
xor UO_1101 (O_1101,N_7688,N_7965);
or UO_1102 (O_1102,N_8419,N_9701);
and UO_1103 (O_1103,N_9071,N_9479);
or UO_1104 (O_1104,N_7819,N_9024);
xnor UO_1105 (O_1105,N_8486,N_7947);
nand UO_1106 (O_1106,N_8599,N_8605);
and UO_1107 (O_1107,N_9887,N_8333);
and UO_1108 (O_1108,N_7504,N_9102);
and UO_1109 (O_1109,N_8978,N_8102);
nand UO_1110 (O_1110,N_8769,N_7530);
nor UO_1111 (O_1111,N_8064,N_7603);
nand UO_1112 (O_1112,N_8914,N_9415);
or UO_1113 (O_1113,N_8675,N_9427);
or UO_1114 (O_1114,N_9574,N_8179);
xnor UO_1115 (O_1115,N_8331,N_9630);
nor UO_1116 (O_1116,N_8562,N_9908);
and UO_1117 (O_1117,N_9927,N_9207);
nand UO_1118 (O_1118,N_8409,N_8000);
nand UO_1119 (O_1119,N_7843,N_8950);
xor UO_1120 (O_1120,N_9769,N_9725);
nor UO_1121 (O_1121,N_9005,N_9413);
and UO_1122 (O_1122,N_8606,N_8869);
xor UO_1123 (O_1123,N_8077,N_7743);
or UO_1124 (O_1124,N_9568,N_8160);
or UO_1125 (O_1125,N_8504,N_7645);
xnor UO_1126 (O_1126,N_9246,N_7744);
or UO_1127 (O_1127,N_8939,N_7894);
and UO_1128 (O_1128,N_8294,N_9385);
xnor UO_1129 (O_1129,N_8420,N_8703);
or UO_1130 (O_1130,N_9737,N_7956);
and UO_1131 (O_1131,N_8999,N_8694);
or UO_1132 (O_1132,N_9367,N_8937);
nand UO_1133 (O_1133,N_7508,N_8896);
and UO_1134 (O_1134,N_9687,N_7572);
nor UO_1135 (O_1135,N_7818,N_8567);
nand UO_1136 (O_1136,N_9801,N_7736);
or UO_1137 (O_1137,N_8201,N_8506);
xnor UO_1138 (O_1138,N_9676,N_9697);
and UO_1139 (O_1139,N_7765,N_9804);
nor UO_1140 (O_1140,N_8181,N_8301);
or UO_1141 (O_1141,N_8718,N_9173);
nor UO_1142 (O_1142,N_9984,N_8335);
nand UO_1143 (O_1143,N_8305,N_8173);
or UO_1144 (O_1144,N_9531,N_8485);
nand UO_1145 (O_1145,N_7571,N_8075);
and UO_1146 (O_1146,N_8844,N_8565);
nor UO_1147 (O_1147,N_8635,N_7695);
or UO_1148 (O_1148,N_7623,N_9970);
nor UO_1149 (O_1149,N_9766,N_7558);
or UO_1150 (O_1150,N_9917,N_9151);
nor UO_1151 (O_1151,N_7518,N_7633);
and UO_1152 (O_1152,N_8219,N_9225);
nor UO_1153 (O_1153,N_9558,N_9949);
nor UO_1154 (O_1154,N_8559,N_8682);
and UO_1155 (O_1155,N_9354,N_8785);
nand UO_1156 (O_1156,N_9028,N_9572);
nand UO_1157 (O_1157,N_8153,N_9661);
and UO_1158 (O_1158,N_7580,N_7564);
nand UO_1159 (O_1159,N_8799,N_8941);
or UO_1160 (O_1160,N_8725,N_8729);
and UO_1161 (O_1161,N_9864,N_9752);
nand UO_1162 (O_1162,N_8392,N_8921);
xor UO_1163 (O_1163,N_8927,N_8971);
nor UO_1164 (O_1164,N_7590,N_8454);
nor UO_1165 (O_1165,N_8520,N_8609);
or UO_1166 (O_1166,N_7705,N_9593);
or UO_1167 (O_1167,N_9925,N_8819);
or UO_1168 (O_1168,N_8912,N_8693);
or UO_1169 (O_1169,N_8012,N_9686);
and UO_1170 (O_1170,N_9517,N_7972);
xnor UO_1171 (O_1171,N_8161,N_8358);
and UO_1172 (O_1172,N_9070,N_8973);
nor UO_1173 (O_1173,N_9587,N_9948);
and UO_1174 (O_1174,N_7532,N_8473);
nand UO_1175 (O_1175,N_7542,N_8404);
nor UO_1176 (O_1176,N_8154,N_8739);
xor UO_1177 (O_1177,N_9444,N_8745);
nor UO_1178 (O_1178,N_9023,N_8843);
nor UO_1179 (O_1179,N_8631,N_9449);
nand UO_1180 (O_1180,N_9231,N_9841);
xnor UO_1181 (O_1181,N_7568,N_7729);
or UO_1182 (O_1182,N_9052,N_9353);
xor UO_1183 (O_1183,N_9520,N_7653);
and UO_1184 (O_1184,N_9014,N_8893);
nor UO_1185 (O_1185,N_9790,N_8081);
nand UO_1186 (O_1186,N_9883,N_8402);
xnor UO_1187 (O_1187,N_8345,N_7830);
nand UO_1188 (O_1188,N_9399,N_7924);
nor UO_1189 (O_1189,N_7502,N_7791);
and UO_1190 (O_1190,N_9333,N_8577);
and UO_1191 (O_1191,N_8947,N_9600);
and UO_1192 (O_1192,N_8466,N_9511);
nor UO_1193 (O_1193,N_8151,N_9524);
nor UO_1194 (O_1194,N_8540,N_8903);
nand UO_1195 (O_1195,N_8832,N_7684);
and UO_1196 (O_1196,N_8885,N_9217);
and UO_1197 (O_1197,N_8261,N_7794);
or UO_1198 (O_1198,N_8275,N_9242);
nor UO_1199 (O_1199,N_8241,N_7893);
xor UO_1200 (O_1200,N_9767,N_8709);
and UO_1201 (O_1201,N_8365,N_9510);
and UO_1202 (O_1202,N_9003,N_9956);
xnor UO_1203 (O_1203,N_8401,N_9741);
and UO_1204 (O_1204,N_9414,N_9201);
nor UO_1205 (O_1205,N_9953,N_7802);
and UO_1206 (O_1206,N_9718,N_8467);
or UO_1207 (O_1207,N_7536,N_8273);
nor UO_1208 (O_1208,N_7864,N_8833);
nand UO_1209 (O_1209,N_7741,N_9933);
and UO_1210 (O_1210,N_9739,N_8089);
xor UO_1211 (O_1211,N_9393,N_8271);
or UO_1212 (O_1212,N_9388,N_7547);
or UO_1213 (O_1213,N_7978,N_8246);
or UO_1214 (O_1214,N_9129,N_8150);
nor UO_1215 (O_1215,N_8632,N_9937);
nand UO_1216 (O_1216,N_8449,N_9746);
xor UO_1217 (O_1217,N_9125,N_7690);
nor UO_1218 (O_1218,N_9538,N_8088);
nand UO_1219 (O_1219,N_8302,N_8097);
and UO_1220 (O_1220,N_7848,N_9732);
nor UO_1221 (O_1221,N_9472,N_9564);
nand UO_1222 (O_1222,N_8313,N_7870);
nand UO_1223 (O_1223,N_8752,N_7533);
nor UO_1224 (O_1224,N_8733,N_8352);
xor UO_1225 (O_1225,N_7682,N_7596);
or UO_1226 (O_1226,N_8545,N_9431);
nand UO_1227 (O_1227,N_8917,N_8085);
and UO_1228 (O_1228,N_8297,N_9578);
nand UO_1229 (O_1229,N_9093,N_8898);
nand UO_1230 (O_1230,N_7878,N_8768);
nand UO_1231 (O_1231,N_8572,N_7676);
nand UO_1232 (O_1232,N_7875,N_8968);
nor UO_1233 (O_1233,N_7593,N_9681);
and UO_1234 (O_1234,N_7977,N_9334);
nand UO_1235 (O_1235,N_8796,N_9309);
nor UO_1236 (O_1236,N_8737,N_9165);
and UO_1237 (O_1237,N_9720,N_9703);
nor UO_1238 (O_1238,N_8873,N_7725);
and UO_1239 (O_1239,N_8096,N_8938);
and UO_1240 (O_1240,N_9929,N_9930);
and UO_1241 (O_1241,N_7982,N_9867);
nor UO_1242 (O_1242,N_9540,N_8048);
and UO_1243 (O_1243,N_9693,N_8513);
or UO_1244 (O_1244,N_7719,N_9842);
nand UO_1245 (O_1245,N_9694,N_8574);
or UO_1246 (O_1246,N_8432,N_9897);
and UO_1247 (O_1247,N_8447,N_8786);
nand UO_1248 (O_1248,N_8802,N_9590);
nor UO_1249 (O_1249,N_9330,N_7585);
xnor UO_1250 (O_1250,N_9649,N_7882);
and UO_1251 (O_1251,N_9583,N_8855);
or UO_1252 (O_1252,N_8539,N_7564);
nand UO_1253 (O_1253,N_8465,N_8178);
nand UO_1254 (O_1254,N_9904,N_8426);
or UO_1255 (O_1255,N_7692,N_8982);
xor UO_1256 (O_1256,N_7505,N_8865);
xor UO_1257 (O_1257,N_9001,N_7968);
nand UO_1258 (O_1258,N_9363,N_8104);
or UO_1259 (O_1259,N_9447,N_9388);
and UO_1260 (O_1260,N_8281,N_9962);
and UO_1261 (O_1261,N_8314,N_8687);
nand UO_1262 (O_1262,N_8709,N_9290);
xnor UO_1263 (O_1263,N_9336,N_9944);
and UO_1264 (O_1264,N_9549,N_9150);
nand UO_1265 (O_1265,N_8211,N_8282);
xor UO_1266 (O_1266,N_8972,N_7770);
or UO_1267 (O_1267,N_8792,N_8471);
nor UO_1268 (O_1268,N_9118,N_7697);
and UO_1269 (O_1269,N_9257,N_8731);
or UO_1270 (O_1270,N_9888,N_8828);
nand UO_1271 (O_1271,N_7898,N_8390);
nor UO_1272 (O_1272,N_9321,N_8084);
nand UO_1273 (O_1273,N_7560,N_8261);
or UO_1274 (O_1274,N_7776,N_7999);
nor UO_1275 (O_1275,N_8790,N_8903);
nand UO_1276 (O_1276,N_7843,N_8982);
nand UO_1277 (O_1277,N_9776,N_9507);
or UO_1278 (O_1278,N_8389,N_9701);
or UO_1279 (O_1279,N_7832,N_8329);
nand UO_1280 (O_1280,N_8972,N_7864);
nand UO_1281 (O_1281,N_8610,N_9955);
and UO_1282 (O_1282,N_8751,N_9467);
or UO_1283 (O_1283,N_9543,N_9748);
nor UO_1284 (O_1284,N_7751,N_7880);
nand UO_1285 (O_1285,N_7846,N_8854);
and UO_1286 (O_1286,N_9881,N_9087);
nand UO_1287 (O_1287,N_7773,N_7833);
xor UO_1288 (O_1288,N_8302,N_8178);
nand UO_1289 (O_1289,N_9116,N_8561);
and UO_1290 (O_1290,N_9862,N_8329);
and UO_1291 (O_1291,N_8990,N_8733);
or UO_1292 (O_1292,N_7878,N_9510);
or UO_1293 (O_1293,N_9576,N_8171);
and UO_1294 (O_1294,N_9334,N_8075);
nand UO_1295 (O_1295,N_9992,N_8554);
nor UO_1296 (O_1296,N_9506,N_8429);
and UO_1297 (O_1297,N_8085,N_7940);
or UO_1298 (O_1298,N_9642,N_8600);
and UO_1299 (O_1299,N_8169,N_8391);
and UO_1300 (O_1300,N_8621,N_8461);
nor UO_1301 (O_1301,N_8597,N_7711);
nor UO_1302 (O_1302,N_8715,N_8933);
nor UO_1303 (O_1303,N_8855,N_9556);
nor UO_1304 (O_1304,N_8689,N_9244);
nand UO_1305 (O_1305,N_9848,N_9891);
xnor UO_1306 (O_1306,N_9276,N_9163);
xnor UO_1307 (O_1307,N_8221,N_9873);
nand UO_1308 (O_1308,N_8123,N_9777);
nor UO_1309 (O_1309,N_9641,N_7761);
xor UO_1310 (O_1310,N_7829,N_7609);
and UO_1311 (O_1311,N_9575,N_8511);
xnor UO_1312 (O_1312,N_9514,N_7574);
or UO_1313 (O_1313,N_8918,N_8397);
nand UO_1314 (O_1314,N_9972,N_8348);
or UO_1315 (O_1315,N_8210,N_8916);
nor UO_1316 (O_1316,N_9018,N_9223);
or UO_1317 (O_1317,N_9650,N_9329);
nand UO_1318 (O_1318,N_8263,N_9338);
nor UO_1319 (O_1319,N_7526,N_9899);
nand UO_1320 (O_1320,N_8944,N_9244);
nor UO_1321 (O_1321,N_8521,N_7661);
and UO_1322 (O_1322,N_8907,N_9489);
nor UO_1323 (O_1323,N_9073,N_9117);
nor UO_1324 (O_1324,N_8016,N_8564);
nor UO_1325 (O_1325,N_9199,N_8886);
nor UO_1326 (O_1326,N_8614,N_9251);
or UO_1327 (O_1327,N_7922,N_9537);
and UO_1328 (O_1328,N_8298,N_7626);
or UO_1329 (O_1329,N_8408,N_7957);
or UO_1330 (O_1330,N_9711,N_8730);
nand UO_1331 (O_1331,N_9621,N_8630);
or UO_1332 (O_1332,N_9294,N_9664);
and UO_1333 (O_1333,N_9411,N_8927);
and UO_1334 (O_1334,N_7651,N_8563);
and UO_1335 (O_1335,N_7626,N_7909);
xor UO_1336 (O_1336,N_8907,N_7731);
nor UO_1337 (O_1337,N_9006,N_8143);
nand UO_1338 (O_1338,N_9107,N_9170);
xor UO_1339 (O_1339,N_8485,N_9325);
nor UO_1340 (O_1340,N_8715,N_9441);
nor UO_1341 (O_1341,N_9084,N_9267);
or UO_1342 (O_1342,N_8224,N_9027);
and UO_1343 (O_1343,N_8728,N_8373);
or UO_1344 (O_1344,N_8181,N_8220);
or UO_1345 (O_1345,N_9188,N_8883);
or UO_1346 (O_1346,N_9734,N_9163);
nor UO_1347 (O_1347,N_9722,N_9904);
nand UO_1348 (O_1348,N_8918,N_8514);
or UO_1349 (O_1349,N_8848,N_9155);
and UO_1350 (O_1350,N_9026,N_7735);
and UO_1351 (O_1351,N_9044,N_9685);
nor UO_1352 (O_1352,N_7833,N_8194);
and UO_1353 (O_1353,N_7746,N_9982);
or UO_1354 (O_1354,N_9207,N_9680);
nor UO_1355 (O_1355,N_8535,N_8629);
or UO_1356 (O_1356,N_7780,N_9757);
nand UO_1357 (O_1357,N_9034,N_8396);
xor UO_1358 (O_1358,N_7818,N_9517);
or UO_1359 (O_1359,N_8022,N_7704);
nor UO_1360 (O_1360,N_8114,N_8972);
or UO_1361 (O_1361,N_7585,N_8989);
and UO_1362 (O_1362,N_9366,N_7642);
xnor UO_1363 (O_1363,N_7748,N_8421);
nand UO_1364 (O_1364,N_9687,N_9958);
and UO_1365 (O_1365,N_7545,N_8505);
nand UO_1366 (O_1366,N_9731,N_9188);
nand UO_1367 (O_1367,N_9877,N_7751);
or UO_1368 (O_1368,N_7629,N_7931);
or UO_1369 (O_1369,N_8384,N_7697);
or UO_1370 (O_1370,N_7739,N_9787);
nor UO_1371 (O_1371,N_8380,N_8314);
and UO_1372 (O_1372,N_8541,N_9605);
and UO_1373 (O_1373,N_8497,N_9109);
or UO_1374 (O_1374,N_8989,N_8706);
nand UO_1375 (O_1375,N_8946,N_9709);
nand UO_1376 (O_1376,N_8635,N_7526);
or UO_1377 (O_1377,N_9413,N_9812);
nor UO_1378 (O_1378,N_9206,N_9957);
or UO_1379 (O_1379,N_9339,N_7992);
and UO_1380 (O_1380,N_9402,N_9844);
xor UO_1381 (O_1381,N_8052,N_8865);
nor UO_1382 (O_1382,N_7606,N_9169);
and UO_1383 (O_1383,N_8630,N_8952);
nand UO_1384 (O_1384,N_9583,N_9933);
nor UO_1385 (O_1385,N_9673,N_9376);
or UO_1386 (O_1386,N_8839,N_9110);
or UO_1387 (O_1387,N_9162,N_9650);
and UO_1388 (O_1388,N_8425,N_9511);
or UO_1389 (O_1389,N_8839,N_7543);
and UO_1390 (O_1390,N_7849,N_7613);
nor UO_1391 (O_1391,N_9128,N_8082);
nor UO_1392 (O_1392,N_9433,N_8640);
nand UO_1393 (O_1393,N_8278,N_9767);
or UO_1394 (O_1394,N_8406,N_8578);
nand UO_1395 (O_1395,N_7975,N_9862);
or UO_1396 (O_1396,N_7830,N_8848);
nor UO_1397 (O_1397,N_7972,N_9529);
and UO_1398 (O_1398,N_7833,N_9507);
and UO_1399 (O_1399,N_8211,N_8877);
nor UO_1400 (O_1400,N_7832,N_7754);
nand UO_1401 (O_1401,N_7562,N_9369);
nor UO_1402 (O_1402,N_9233,N_7785);
and UO_1403 (O_1403,N_8302,N_8520);
nor UO_1404 (O_1404,N_9477,N_9551);
nor UO_1405 (O_1405,N_9207,N_8127);
or UO_1406 (O_1406,N_9717,N_9200);
or UO_1407 (O_1407,N_9433,N_7733);
and UO_1408 (O_1408,N_9404,N_9748);
and UO_1409 (O_1409,N_8667,N_9022);
nor UO_1410 (O_1410,N_9147,N_8141);
or UO_1411 (O_1411,N_8660,N_9836);
or UO_1412 (O_1412,N_8291,N_9207);
xnor UO_1413 (O_1413,N_8058,N_9204);
nor UO_1414 (O_1414,N_9536,N_8046);
nor UO_1415 (O_1415,N_8357,N_9206);
xor UO_1416 (O_1416,N_7522,N_8370);
nand UO_1417 (O_1417,N_8128,N_8307);
and UO_1418 (O_1418,N_7578,N_9832);
nand UO_1419 (O_1419,N_9904,N_9198);
nor UO_1420 (O_1420,N_7718,N_9414);
and UO_1421 (O_1421,N_8341,N_8453);
or UO_1422 (O_1422,N_9929,N_9529);
nor UO_1423 (O_1423,N_7836,N_9495);
and UO_1424 (O_1424,N_8145,N_9896);
nor UO_1425 (O_1425,N_8745,N_9373);
and UO_1426 (O_1426,N_9346,N_9979);
nand UO_1427 (O_1427,N_7593,N_8402);
or UO_1428 (O_1428,N_7583,N_7508);
or UO_1429 (O_1429,N_8769,N_8136);
nor UO_1430 (O_1430,N_8574,N_7637);
or UO_1431 (O_1431,N_9232,N_8648);
or UO_1432 (O_1432,N_8656,N_8075);
nor UO_1433 (O_1433,N_7633,N_8936);
nand UO_1434 (O_1434,N_9651,N_8525);
or UO_1435 (O_1435,N_8798,N_8127);
nand UO_1436 (O_1436,N_8942,N_8059);
nand UO_1437 (O_1437,N_8090,N_8756);
nor UO_1438 (O_1438,N_9468,N_7812);
nand UO_1439 (O_1439,N_8119,N_9035);
and UO_1440 (O_1440,N_7943,N_7697);
nand UO_1441 (O_1441,N_7629,N_9544);
or UO_1442 (O_1442,N_8196,N_8934);
and UO_1443 (O_1443,N_7522,N_9414);
and UO_1444 (O_1444,N_9615,N_8462);
or UO_1445 (O_1445,N_7783,N_7898);
nor UO_1446 (O_1446,N_9683,N_8184);
or UO_1447 (O_1447,N_8234,N_8921);
nand UO_1448 (O_1448,N_9609,N_9103);
and UO_1449 (O_1449,N_8338,N_9112);
xnor UO_1450 (O_1450,N_9963,N_7732);
nor UO_1451 (O_1451,N_9206,N_7744);
and UO_1452 (O_1452,N_9937,N_8691);
nor UO_1453 (O_1453,N_9593,N_8349);
and UO_1454 (O_1454,N_8975,N_8217);
nor UO_1455 (O_1455,N_8894,N_7750);
xnor UO_1456 (O_1456,N_8421,N_9234);
and UO_1457 (O_1457,N_9938,N_9106);
nand UO_1458 (O_1458,N_7875,N_8722);
or UO_1459 (O_1459,N_7892,N_9267);
and UO_1460 (O_1460,N_9862,N_8273);
nor UO_1461 (O_1461,N_9006,N_7885);
and UO_1462 (O_1462,N_7517,N_8875);
nand UO_1463 (O_1463,N_9771,N_9477);
nand UO_1464 (O_1464,N_8143,N_9955);
nor UO_1465 (O_1465,N_8218,N_9273);
and UO_1466 (O_1466,N_9497,N_8122);
or UO_1467 (O_1467,N_8272,N_8344);
and UO_1468 (O_1468,N_8931,N_8402);
and UO_1469 (O_1469,N_9325,N_9984);
nand UO_1470 (O_1470,N_9694,N_8580);
nand UO_1471 (O_1471,N_9653,N_8138);
and UO_1472 (O_1472,N_9528,N_7787);
or UO_1473 (O_1473,N_9080,N_8093);
and UO_1474 (O_1474,N_7907,N_9524);
or UO_1475 (O_1475,N_8797,N_7601);
nor UO_1476 (O_1476,N_9702,N_8892);
or UO_1477 (O_1477,N_9144,N_7996);
or UO_1478 (O_1478,N_8827,N_8422);
nor UO_1479 (O_1479,N_9995,N_7827);
nand UO_1480 (O_1480,N_9862,N_8600);
xor UO_1481 (O_1481,N_8101,N_7830);
or UO_1482 (O_1482,N_9077,N_7587);
nor UO_1483 (O_1483,N_8114,N_9079);
or UO_1484 (O_1484,N_8727,N_9084);
or UO_1485 (O_1485,N_9837,N_8312);
and UO_1486 (O_1486,N_7695,N_9550);
nor UO_1487 (O_1487,N_7744,N_9309);
nand UO_1488 (O_1488,N_9737,N_9902);
nand UO_1489 (O_1489,N_8118,N_9762);
and UO_1490 (O_1490,N_9371,N_9570);
and UO_1491 (O_1491,N_9458,N_9022);
nor UO_1492 (O_1492,N_8745,N_8084);
nand UO_1493 (O_1493,N_7898,N_9379);
and UO_1494 (O_1494,N_9357,N_9149);
nor UO_1495 (O_1495,N_9360,N_9017);
or UO_1496 (O_1496,N_8085,N_7881);
or UO_1497 (O_1497,N_8288,N_9091);
nand UO_1498 (O_1498,N_7801,N_7913);
or UO_1499 (O_1499,N_9889,N_8367);
endmodule