module basic_2500_25000_3000_25_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_1668,In_1412);
and U1 (N_1,In_94,In_623);
nand U2 (N_2,In_1643,In_655);
nand U3 (N_3,In_1437,In_1228);
xor U4 (N_4,In_1788,In_1832);
and U5 (N_5,In_1589,In_410);
and U6 (N_6,In_1120,In_398);
nor U7 (N_7,In_934,In_1719);
xor U8 (N_8,In_172,In_2262);
and U9 (N_9,In_241,In_558);
nand U10 (N_10,In_367,In_220);
nand U11 (N_11,In_1445,In_1128);
or U12 (N_12,In_1200,In_546);
nor U13 (N_13,In_1564,In_2103);
nor U14 (N_14,In_628,In_753);
or U15 (N_15,In_920,In_1350);
and U16 (N_16,In_661,In_861);
and U17 (N_17,In_421,In_474);
nor U18 (N_18,In_1787,In_1593);
nand U19 (N_19,In_1214,In_2159);
or U20 (N_20,In_1042,In_432);
xor U21 (N_21,In_1783,In_944);
xor U22 (N_22,In_1226,In_219);
or U23 (N_23,In_98,In_2038);
or U24 (N_24,In_201,In_174);
xnor U25 (N_25,In_563,In_1);
nor U26 (N_26,In_2396,In_1117);
xnor U27 (N_27,In_2242,In_1076);
or U28 (N_28,In_783,In_381);
nand U29 (N_29,In_2042,In_1360);
nand U30 (N_30,In_2344,In_1508);
and U31 (N_31,In_1623,In_109);
nand U32 (N_32,In_1322,In_1365);
xor U33 (N_33,In_956,In_2354);
xnor U34 (N_34,In_2138,In_642);
or U35 (N_35,In_1880,In_591);
nor U36 (N_36,In_2264,In_518);
nor U37 (N_37,In_871,In_1709);
xnor U38 (N_38,In_851,In_2449);
and U39 (N_39,In_1974,In_771);
nor U40 (N_40,In_1418,In_1062);
nor U41 (N_41,In_133,In_1960);
nor U42 (N_42,In_1395,In_415);
nand U43 (N_43,In_1969,In_1924);
and U44 (N_44,In_567,In_1786);
xor U45 (N_45,In_2431,In_1530);
or U46 (N_46,In_1679,In_1081);
and U47 (N_47,In_217,In_1646);
and U48 (N_48,In_1420,In_15);
or U49 (N_49,In_2030,In_490);
nand U50 (N_50,In_941,In_53);
or U51 (N_51,In_1683,In_165);
or U52 (N_52,In_849,In_1381);
xnor U53 (N_53,In_1998,In_1136);
and U54 (N_54,In_1636,In_2274);
xor U55 (N_55,In_1941,In_2395);
xor U56 (N_56,In_509,In_1665);
or U57 (N_57,In_646,In_428);
nor U58 (N_58,In_2417,In_2153);
nor U59 (N_59,In_63,In_643);
and U60 (N_60,In_2209,In_859);
or U61 (N_61,In_2423,In_1949);
xnor U62 (N_62,In_297,In_1246);
and U63 (N_63,In_1003,In_1052);
nand U64 (N_64,In_1304,In_1056);
nor U65 (N_65,In_78,In_1111);
nand U66 (N_66,In_1142,In_190);
and U67 (N_67,In_669,In_2056);
and U68 (N_68,In_2244,In_1410);
or U69 (N_69,In_1194,In_817);
xnor U70 (N_70,In_1116,In_931);
nand U71 (N_71,In_812,In_2425);
or U72 (N_72,In_1385,In_2194);
or U73 (N_73,In_734,In_850);
and U74 (N_74,In_1925,In_1827);
and U75 (N_75,In_1202,In_831);
or U76 (N_76,In_348,In_2422);
and U77 (N_77,In_89,In_2129);
nand U78 (N_78,In_1225,In_728);
and U79 (N_79,In_589,In_491);
or U80 (N_80,In_1298,In_166);
and U81 (N_81,In_1104,In_1990);
nor U82 (N_82,In_2191,In_1959);
nor U83 (N_83,In_1460,In_2022);
or U84 (N_84,In_488,In_664);
or U85 (N_85,In_2066,In_1160);
xor U86 (N_86,In_2321,In_1448);
or U87 (N_87,In_586,In_67);
nor U88 (N_88,In_1963,In_275);
and U89 (N_89,In_696,In_2310);
xnor U90 (N_90,In_1201,In_289);
or U91 (N_91,In_1491,In_306);
xnor U92 (N_92,In_1218,In_672);
nor U93 (N_93,In_878,In_933);
xnor U94 (N_94,In_1957,In_1835);
and U95 (N_95,In_2443,In_131);
xor U96 (N_96,In_1414,In_1720);
nor U97 (N_97,In_2370,In_1625);
or U98 (N_98,In_2095,In_1951);
nand U99 (N_99,In_832,In_435);
or U100 (N_100,In_1635,In_1544);
nor U101 (N_101,In_2466,In_952);
or U102 (N_102,In_1287,In_2491);
or U103 (N_103,In_1729,In_2199);
nor U104 (N_104,In_1687,In_1399);
and U105 (N_105,In_240,In_577);
and U106 (N_106,In_1540,In_2086);
nor U107 (N_107,In_20,In_2338);
nand U108 (N_108,In_310,In_132);
xnor U109 (N_109,In_1041,In_1098);
and U110 (N_110,In_1917,In_498);
nor U111 (N_111,In_691,In_632);
nand U112 (N_112,In_2172,In_1284);
nor U113 (N_113,In_1782,In_2205);
xor U114 (N_114,In_901,In_128);
or U115 (N_115,In_2015,In_343);
nor U116 (N_116,In_1517,In_1475);
and U117 (N_117,In_1693,In_856);
xnor U118 (N_118,In_980,In_1197);
and U119 (N_119,In_1309,In_1223);
and U120 (N_120,In_1691,In_1581);
or U121 (N_121,In_2365,In_2142);
nand U122 (N_122,In_2432,In_1740);
xor U123 (N_123,In_2118,In_1600);
and U124 (N_124,In_2345,In_1572);
nand U125 (N_125,In_722,In_1697);
or U126 (N_126,In_358,In_688);
and U127 (N_127,In_627,In_705);
nor U128 (N_128,In_1770,In_1807);
nor U129 (N_129,In_370,In_62);
and U130 (N_130,In_227,In_2125);
or U131 (N_131,In_329,In_246);
nor U132 (N_132,In_638,In_56);
and U133 (N_133,In_982,In_2412);
and U134 (N_134,In_870,In_465);
or U135 (N_135,In_855,In_2011);
nand U136 (N_136,In_829,In_976);
nor U137 (N_137,In_888,In_1473);
nor U138 (N_138,In_516,In_2104);
or U139 (N_139,In_1670,In_1886);
nand U140 (N_140,In_780,In_1532);
nor U141 (N_141,In_104,In_2411);
or U142 (N_142,In_1597,In_1036);
and U143 (N_143,In_894,In_947);
and U144 (N_144,In_1983,In_804);
nor U145 (N_145,In_887,In_1895);
or U146 (N_146,In_729,In_1909);
and U147 (N_147,In_186,In_30);
nand U148 (N_148,In_234,In_1565);
and U149 (N_149,In_2471,In_1518);
nand U150 (N_150,In_653,In_704);
nand U151 (N_151,In_1192,In_2083);
or U152 (N_152,In_196,In_2130);
nand U153 (N_153,In_147,In_1483);
and U154 (N_154,In_1413,In_1723);
nand U155 (N_155,In_922,In_203);
or U156 (N_156,In_2091,In_71);
nor U157 (N_157,In_2171,In_1255);
nor U158 (N_158,In_755,In_1373);
and U159 (N_159,In_948,In_46);
xor U160 (N_160,In_1332,In_2415);
and U161 (N_161,In_200,In_2406);
and U162 (N_162,In_2419,In_77);
and U163 (N_163,In_808,In_288);
or U164 (N_164,In_1376,In_212);
or U165 (N_165,In_2223,In_1942);
nand U166 (N_166,In_1520,In_1308);
xnor U167 (N_167,In_2385,In_60);
xnor U168 (N_168,In_2486,In_1922);
nor U169 (N_169,In_1617,In_2071);
xnor U170 (N_170,In_479,In_1962);
or U171 (N_171,In_559,In_304);
nand U172 (N_172,In_1888,In_1912);
xnor U173 (N_173,In_1848,In_608);
nand U174 (N_174,In_924,In_1768);
and U175 (N_175,In_1979,In_1588);
and U176 (N_176,In_1569,In_445);
nor U177 (N_177,In_2427,In_885);
and U178 (N_178,In_2455,In_1575);
and U179 (N_179,In_2361,In_493);
nand U180 (N_180,In_501,In_857);
nor U181 (N_181,In_1776,In_2026);
or U182 (N_182,In_2436,In_576);
and U183 (N_183,In_1059,In_156);
nand U184 (N_184,In_716,In_2416);
nor U185 (N_185,In_9,In_469);
or U186 (N_186,In_295,In_754);
nor U187 (N_187,In_1372,In_1889);
nor U188 (N_188,In_587,In_905);
nor U189 (N_189,In_2219,In_112);
and U190 (N_190,In_207,In_703);
or U191 (N_191,In_2243,In_1987);
or U192 (N_192,In_507,In_300);
xnor U193 (N_193,In_351,In_860);
nand U194 (N_194,In_1171,In_631);
or U195 (N_195,In_1604,In_176);
and U196 (N_196,In_1151,In_1290);
or U197 (N_197,In_64,In_1640);
or U198 (N_198,In_1358,In_1337);
nand U199 (N_199,In_1451,In_1738);
or U200 (N_200,In_1083,In_611);
nor U201 (N_201,In_896,In_2369);
nor U202 (N_202,In_1986,In_929);
or U203 (N_203,In_777,In_2231);
nor U204 (N_204,In_2263,In_650);
and U205 (N_205,In_677,In_1557);
or U206 (N_206,In_1237,In_387);
or U207 (N_207,In_1292,In_2300);
or U208 (N_208,In_249,In_1583);
nand U209 (N_209,In_1995,In_13);
nor U210 (N_210,In_1245,In_2034);
nand U211 (N_211,In_1073,In_583);
nand U212 (N_212,In_1749,In_195);
nand U213 (N_213,In_1044,In_1150);
nand U214 (N_214,In_597,In_1512);
nor U215 (N_215,In_588,In_1933);
nor U216 (N_216,In_545,In_450);
or U217 (N_217,In_2311,In_265);
xor U218 (N_218,In_1844,In_1647);
nor U219 (N_219,In_2144,In_1882);
or U220 (N_220,In_2201,In_290);
and U221 (N_221,In_331,In_1836);
xor U222 (N_222,In_1248,In_1898);
nor U223 (N_223,In_1725,In_2331);
nor U224 (N_224,In_1015,In_1459);
xor U225 (N_225,In_1400,In_940);
and U226 (N_226,In_1904,In_1490);
and U227 (N_227,In_1868,In_205);
or U228 (N_228,In_1032,In_120);
nor U229 (N_229,In_764,In_153);
nor U230 (N_230,In_2124,In_2247);
and U231 (N_231,In_87,In_1954);
nor U232 (N_232,In_333,In_2102);
nand U233 (N_233,In_2452,In_845);
nor U234 (N_234,In_1130,In_273);
nand U235 (N_235,In_515,In_2096);
nor U236 (N_236,In_2313,In_1185);
nor U237 (N_237,In_1541,In_2053);
or U238 (N_238,In_1436,In_715);
nand U239 (N_239,In_1580,In_1072);
nand U240 (N_240,In_167,In_407);
nand U241 (N_241,In_1352,In_414);
nor U242 (N_242,In_2013,In_1096);
nand U243 (N_243,In_278,In_2043);
or U244 (N_244,In_1118,In_1531);
xnor U245 (N_245,In_995,In_1433);
or U246 (N_246,In_1270,In_1441);
or U247 (N_247,In_247,In_2012);
xor U248 (N_248,In_1762,In_2101);
and U249 (N_249,In_698,In_1856);
nand U250 (N_250,In_2327,In_745);
xor U251 (N_251,In_1823,In_1037);
xnor U252 (N_252,In_315,In_1966);
nand U253 (N_253,In_622,In_969);
or U254 (N_254,In_2460,In_437);
and U255 (N_255,In_1462,In_732);
and U256 (N_256,In_594,In_1129);
nand U257 (N_257,In_34,In_937);
and U258 (N_258,In_1897,In_429);
xor U259 (N_259,In_1053,In_1145);
xnor U260 (N_260,In_2177,In_897);
or U261 (N_261,In_2348,In_1892);
xor U262 (N_262,In_2413,In_1285);
nor U263 (N_263,In_266,In_1064);
nand U264 (N_264,In_1268,In_1217);
nand U265 (N_265,In_1453,In_1428);
xor U266 (N_266,In_868,In_2484);
nand U267 (N_267,In_1434,In_2170);
or U268 (N_268,In_2081,In_335);
nand U269 (N_269,In_309,In_1272);
nand U270 (N_270,In_447,In_682);
and U271 (N_271,In_746,In_1411);
xnor U272 (N_272,In_1988,In_1497);
nand U273 (N_273,In_1642,In_575);
or U274 (N_274,In_2240,In_1535);
and U275 (N_275,In_2445,In_842);
and U276 (N_276,In_1791,In_1113);
nor U277 (N_277,In_547,In_399);
nor U278 (N_278,In_1103,In_1521);
xnor U279 (N_279,In_1847,In_770);
and U280 (N_280,In_264,In_1769);
and U281 (N_281,In_532,In_1896);
and U282 (N_282,In_1065,In_1254);
nand U283 (N_283,In_1560,In_25);
and U284 (N_284,In_1672,In_2438);
and U285 (N_285,In_1085,In_464);
nor U286 (N_286,In_621,In_139);
nor U287 (N_287,In_449,In_544);
xnor U288 (N_288,In_117,In_340);
nand U289 (N_289,In_797,In_419);
or U290 (N_290,In_97,In_727);
or U291 (N_291,In_1915,In_1877);
or U292 (N_292,In_1108,In_1269);
nand U293 (N_293,In_2324,In_2021);
nand U294 (N_294,In_2155,In_36);
and U295 (N_295,In_1401,In_2383);
or U296 (N_296,In_1476,In_1316);
and U297 (N_297,In_2165,In_2279);
nand U298 (N_298,In_1384,In_882);
nand U299 (N_299,In_1774,In_913);
nand U300 (N_300,In_2010,In_2271);
xnor U301 (N_301,In_1216,In_11);
nand U302 (N_302,In_1916,In_1396);
nand U303 (N_303,In_1137,In_1258);
or U304 (N_304,In_1669,In_1903);
xor U305 (N_305,In_645,In_2210);
or U306 (N_306,In_1566,In_1651);
or U307 (N_307,In_2334,In_83);
xor U308 (N_308,In_2253,In_27);
and U309 (N_309,In_1510,In_1624);
nor U310 (N_310,In_1009,In_2224);
and U311 (N_311,In_2006,In_1492);
xor U312 (N_312,In_765,In_2490);
nor U313 (N_313,In_1961,In_2428);
or U314 (N_314,In_433,In_695);
and U315 (N_315,In_44,In_1523);
and U316 (N_316,In_596,In_1071);
nand U317 (N_317,In_1461,In_803);
xnor U318 (N_318,In_2041,In_1209);
nand U319 (N_319,In_1929,In_1339);
nand U320 (N_320,In_513,In_957);
nor U321 (N_321,In_373,In_1524);
xnor U322 (N_322,In_828,In_1055);
or U323 (N_323,In_2064,In_562);
or U324 (N_324,In_1592,In_303);
xnor U325 (N_325,In_1406,In_379);
or U326 (N_326,In_873,In_1013);
xor U327 (N_327,In_534,In_6);
xnor U328 (N_328,In_1707,In_806);
or U329 (N_329,In_1487,In_1554);
or U330 (N_330,In_2399,In_35);
nand U331 (N_331,In_223,In_2250);
nand U332 (N_332,In_1845,In_946);
and U333 (N_333,In_2197,In_554);
and U334 (N_334,In_1069,In_942);
xor U335 (N_335,In_1944,In_1887);
nor U336 (N_336,In_1378,In_1321);
nand U337 (N_337,In_1463,In_462);
xor U338 (N_338,In_1499,In_101);
nand U339 (N_339,In_720,In_1267);
nand U340 (N_340,In_814,In_2323);
xor U341 (N_341,In_1416,In_709);
nand U342 (N_342,In_2433,In_2414);
or U343 (N_343,In_1975,In_487);
xnor U344 (N_344,In_1379,In_481);
nor U345 (N_345,In_743,In_2418);
xnor U346 (N_346,In_2270,In_424);
xnor U347 (N_347,In_609,In_130);
nor U348 (N_348,In_2157,In_1328);
or U349 (N_349,In_1383,In_2009);
and U350 (N_350,In_907,In_1860);
nand U351 (N_351,In_2248,In_2430);
and U352 (N_352,In_1931,In_1952);
and U353 (N_353,In_209,In_647);
xnor U354 (N_354,In_1934,In_233);
nand U355 (N_355,In_854,In_1872);
or U356 (N_356,In_1455,In_1932);
or U357 (N_357,In_1188,In_838);
nor U358 (N_358,In_1553,In_2000);
nor U359 (N_359,In_4,In_2297);
xnor U360 (N_360,In_2145,In_1031);
nor U361 (N_361,In_1293,In_1910);
nor U362 (N_362,In_1821,In_1191);
or U363 (N_363,In_1386,In_59);
nor U364 (N_364,In_1029,In_1333);
or U365 (N_365,In_65,In_1107);
nand U366 (N_366,In_124,In_438);
nand U367 (N_367,In_1501,In_837);
nand U368 (N_368,In_1800,In_986);
nand U369 (N_369,In_1692,In_2261);
nor U370 (N_370,In_1870,In_29);
or U371 (N_371,In_595,In_569);
or U372 (N_372,In_345,In_269);
or U373 (N_373,In_2057,In_900);
and U374 (N_374,In_2288,In_76);
nand U375 (N_375,In_2320,In_673);
nor U376 (N_376,In_1472,In_1310);
nand U377 (N_377,In_2169,In_1948);
xnor U378 (N_378,In_1450,In_1971);
nor U379 (N_379,In_802,In_665);
and U380 (N_380,In_228,In_108);
and U381 (N_381,In_2454,In_1550);
xnor U382 (N_382,In_1256,In_2273);
xor U383 (N_383,In_640,In_2457);
xor U384 (N_384,In_325,In_150);
xnor U385 (N_385,In_2174,In_2403);
nor U386 (N_386,In_1795,In_1526);
xor U387 (N_387,In_37,In_2234);
nand U388 (N_388,In_1014,In_2150);
xor U389 (N_389,In_1730,In_644);
or U390 (N_390,In_2152,In_283);
xor U391 (N_391,In_1777,In_1573);
nand U392 (N_392,In_884,In_500);
nand U393 (N_393,In_1048,In_107);
nand U394 (N_394,In_1824,In_2285);
nor U395 (N_395,In_235,In_408);
xnor U396 (N_396,In_1489,In_1274);
nand U397 (N_397,In_1712,In_2148);
and U398 (N_398,In_467,In_184);
nand U399 (N_399,In_1250,In_908);
nor U400 (N_400,In_395,In_1846);
nor U401 (N_401,In_185,In_1818);
or U402 (N_402,In_2464,In_144);
nand U403 (N_403,In_1232,In_1803);
or U404 (N_404,In_92,In_881);
nand U405 (N_405,In_899,In_2368);
and U406 (N_406,In_2280,In_489);
and U407 (N_407,In_211,In_675);
or U408 (N_408,In_332,In_2099);
nor U409 (N_409,In_1973,In_1109);
xor U410 (N_410,In_975,In_1480);
nor U411 (N_411,In_510,In_1203);
or U412 (N_412,In_1590,In_1345);
nor U413 (N_413,In_396,In_1562);
nand U414 (N_414,In_148,In_2206);
and U415 (N_415,In_2477,In_1503);
nand U416 (N_416,In_1168,In_23);
nand U417 (N_417,In_91,In_69);
xnor U418 (N_418,In_1721,In_281);
and U419 (N_419,In_2308,In_787);
nor U420 (N_420,In_412,In_2480);
nand U421 (N_421,In_225,In_1112);
and U422 (N_422,In_1249,In_400);
nand U423 (N_423,In_1146,In_1869);
xor U424 (N_424,In_1632,In_2315);
nor U425 (N_425,In_1763,In_1305);
or U426 (N_426,In_1748,In_2173);
and U427 (N_427,In_470,In_157);
nand U428 (N_428,In_21,In_1364);
nand U429 (N_429,In_2003,In_221);
or U430 (N_430,In_173,In_95);
nand U431 (N_431,In_305,In_872);
nor U432 (N_432,In_738,In_85);
and U433 (N_433,In_2487,In_773);
nor U434 (N_434,In_1900,In_1716);
and U435 (N_435,In_1766,In_2070);
nand U436 (N_436,In_431,In_2033);
xor U437 (N_437,In_1866,In_1143);
xor U438 (N_438,In_686,In_1732);
and U439 (N_439,In_1638,In_257);
and U440 (N_440,In_1867,In_127);
and U441 (N_441,In_1528,In_578);
nand U442 (N_442,In_1828,In_1756);
xnor U443 (N_443,In_853,In_2048);
nor U444 (N_444,In_762,In_2218);
nand U445 (N_445,In_2235,In_2494);
nand U446 (N_446,In_981,In_1978);
xnor U447 (N_447,In_1035,In_1746);
and U448 (N_448,In_237,In_336);
nand U449 (N_449,In_1708,In_286);
xnor U450 (N_450,In_1607,In_895);
xor U451 (N_451,In_2291,In_2222);
and U452 (N_452,In_279,In_183);
and U453 (N_453,In_839,In_1348);
nand U454 (N_454,In_2115,In_276);
nor U455 (N_455,In_1063,In_187);
nor U456 (N_456,In_1273,In_1891);
xnor U457 (N_457,In_1853,In_1584);
nand U458 (N_458,In_1264,In_2127);
nand U459 (N_459,In_484,In_1319);
or U460 (N_460,In_604,In_1106);
nor U461 (N_461,In_1481,In_2141);
or U462 (N_462,In_1834,In_1814);
or U463 (N_463,In_1465,In_391);
nand U464 (N_464,In_927,In_1753);
nor U465 (N_465,In_618,In_2497);
or U466 (N_466,In_1792,In_1087);
nor U467 (N_467,In_1519,In_1021);
nand U468 (N_468,In_1813,In_2389);
nand U469 (N_469,In_2175,In_725);
and U470 (N_470,In_911,In_1923);
or U471 (N_471,In_2002,In_2450);
and U472 (N_472,In_180,In_2077);
xnor U473 (N_473,In_1177,In_122);
nor U474 (N_474,In_199,In_811);
or U475 (N_475,In_2133,In_1403);
nor U476 (N_476,In_1389,In_1649);
nand U477 (N_477,In_1755,In_270);
nor U478 (N_478,In_230,In_1559);
xnor U479 (N_479,In_502,In_2364);
nor U480 (N_480,In_494,In_1279);
and U481 (N_481,In_371,In_1294);
nor U482 (N_482,In_566,In_2305);
and U483 (N_483,In_998,In_721);
nand U484 (N_484,In_1387,In_1714);
nand U485 (N_485,In_313,In_1661);
or U486 (N_486,In_48,In_945);
nand U487 (N_487,In_49,In_1057);
nand U488 (N_488,In_1242,In_971);
nor U489 (N_489,In_840,In_1047);
nor U490 (N_490,In_1921,In_82);
nand U491 (N_491,In_1812,In_1645);
xnor U492 (N_492,In_1736,In_12);
xnor U493 (N_493,In_2031,In_1750);
or U494 (N_494,In_816,In_1300);
xnor U495 (N_495,In_2496,In_1193);
nor U496 (N_496,In_321,In_1556);
xor U497 (N_497,In_2162,In_105);
and U498 (N_498,In_2483,In_830);
nand U499 (N_499,In_1017,In_620);
or U500 (N_500,In_496,In_1336);
xor U501 (N_501,In_1608,In_2265);
and U502 (N_502,In_1361,In_74);
nor U503 (N_503,In_1525,In_2404);
nand U504 (N_504,In_452,In_161);
nand U505 (N_505,In_949,In_1049);
nor U506 (N_506,In_1144,In_143);
and U507 (N_507,In_2019,In_2435);
or U508 (N_508,In_193,In_339);
and U509 (N_509,In_2448,In_416);
or U510 (N_510,In_352,In_1377);
and U511 (N_511,In_903,In_2168);
nand U512 (N_512,In_1656,In_1579);
and U513 (N_513,In_271,In_96);
xnor U514 (N_514,In_767,In_1773);
xnor U515 (N_515,In_1878,In_224);
or U516 (N_516,In_1815,In_1680);
nand U517 (N_517,In_324,In_877);
nand U518 (N_518,In_404,In_409);
xnor U519 (N_519,In_2245,In_690);
xnor U520 (N_520,In_1654,In_2356);
nor U521 (N_521,In_1393,In_992);
nor U522 (N_522,In_2330,In_292);
nor U523 (N_523,In_2278,In_1727);
xor U524 (N_524,In_925,In_564);
and U525 (N_525,In_1631,In_598);
and U526 (N_526,In_384,In_2137);
and U527 (N_527,In_1885,In_1811);
nor U528 (N_528,In_605,In_1363);
nand U529 (N_529,In_280,In_1327);
or U530 (N_530,In_926,In_287);
and U531 (N_531,In_2398,In_236);
nor U532 (N_532,In_1101,In_2467);
and U533 (N_533,In_251,In_1210);
or U534 (N_534,In_1198,In_141);
xnor U535 (N_535,In_1516,In_1621);
nand U536 (N_536,In_1905,In_858);
and U537 (N_537,In_1007,In_2342);
nor U538 (N_538,In_813,In_1539);
xnor U539 (N_539,In_1088,In_100);
xor U540 (N_540,In_1630,In_1368);
xnor U541 (N_541,In_2360,In_584);
or U542 (N_542,In_1045,In_751);
and U543 (N_543,In_1612,In_1685);
and U544 (N_544,In_204,In_1391);
nor U545 (N_545,In_1908,In_1174);
xor U546 (N_546,In_1432,In_2329);
nor U547 (N_547,In_1470,In_2207);
xnor U548 (N_548,In_2451,In_1890);
nand U549 (N_549,In_572,In_916);
or U550 (N_550,In_2268,In_1981);
and U551 (N_551,In_1243,In_1667);
or U552 (N_552,In_47,In_38);
and U553 (N_553,In_1555,In_413);
and U554 (N_554,In_2200,In_1090);
or U555 (N_555,In_2446,In_1809);
xnor U556 (N_556,In_2366,In_723);
and U557 (N_557,In_334,In_1928);
and U558 (N_558,In_763,In_439);
nor U559 (N_559,In_2047,In_1307);
nor U560 (N_560,In_2203,In_1231);
and U561 (N_561,In_2226,In_1181);
or U562 (N_562,In_1840,In_260);
nor U563 (N_563,In_2108,In_923);
xnor U564 (N_564,In_114,In_397);
xor U565 (N_565,In_1690,In_548);
and U566 (N_566,In_750,In_1325);
nor U567 (N_567,In_1484,In_1102);
and U568 (N_568,In_2326,In_1970);
xor U569 (N_569,In_1224,In_909);
nand U570 (N_570,In_798,In_2249);
nand U571 (N_571,In_820,In_2190);
and U572 (N_572,In_886,In_113);
or U573 (N_573,In_1675,In_1849);
nand U574 (N_574,In_1999,In_2139);
nor U575 (N_575,In_1236,In_641);
xnor U576 (N_576,In_1089,In_936);
or U577 (N_577,In_2028,In_2470);
nor U578 (N_578,In_1976,In_1852);
xor U579 (N_579,In_1542,In_585);
nor U580 (N_580,In_1700,In_158);
xor U581 (N_581,In_549,In_506);
or U582 (N_582,In_1039,In_90);
xor U583 (N_583,In_2362,In_1686);
and U584 (N_584,In_84,In_668);
nand U585 (N_585,In_955,In_985);
xnor U586 (N_586,In_1251,In_592);
and U587 (N_587,In_1247,In_2420);
nor U588 (N_588,In_1495,In_1012);
or U589 (N_589,In_662,In_766);
and U590 (N_590,In_1182,In_1545);
nor U591 (N_591,In_600,In_2286);
xor U592 (N_592,In_730,In_529);
and U593 (N_593,In_505,In_1810);
nor U594 (N_594,In_556,In_1278);
and U595 (N_595,In_1312,In_1605);
and U596 (N_596,In_2375,In_2405);
nand U597 (N_597,In_31,In_1728);
or U598 (N_598,In_1030,In_2371);
nand U599 (N_599,In_364,In_1235);
xor U600 (N_600,In_436,In_2498);
or U601 (N_601,In_1502,In_1577);
or U602 (N_602,In_1627,In_140);
or U603 (N_603,In_1315,In_2119);
nor U604 (N_604,In_2459,In_2339);
nor U605 (N_605,In_954,In_1789);
nor U606 (N_606,In_2024,In_568);
xor U607 (N_607,In_1169,In_681);
nand U608 (N_608,In_1741,In_2123);
or U609 (N_609,In_993,In_1515);
nand U610 (N_610,In_2098,In_477);
nand U611 (N_611,In_736,In_197);
nor U612 (N_612,In_2289,In_267);
nor U613 (N_613,In_192,In_2252);
xor U614 (N_614,In_473,In_684);
or U615 (N_615,In_2025,In_208);
xor U616 (N_616,In_66,In_2075);
or U617 (N_617,In_1477,In_875);
xor U618 (N_618,In_1747,In_2352);
nand U619 (N_619,In_1159,In_134);
and U620 (N_620,In_2181,In_2134);
xor U621 (N_621,In_483,In_2049);
and U622 (N_622,In_111,In_1291);
or U623 (N_623,In_1563,In_869);
nand U624 (N_624,In_1493,In_966);
or U625 (N_625,In_1861,In_2036);
or U626 (N_626,In_552,In_699);
nor U627 (N_627,In_454,In_1659);
nand U628 (N_628,In_846,In_1710);
or U629 (N_629,In_1939,In_1415);
and U630 (N_630,In_1426,In_2195);
and U631 (N_631,In_243,In_1135);
and U632 (N_632,In_102,In_1040);
and U633 (N_633,In_2179,In_1980);
and U634 (N_634,In_1701,In_1761);
nand U635 (N_635,In_282,In_2088);
nor U636 (N_636,In_962,In_1435);
and U637 (N_637,In_218,In_2151);
nor U638 (N_638,In_659,In_177);
xnor U639 (N_639,In_914,In_1155);
nor U640 (N_640,In_327,In_360);
and U641 (N_641,In_2355,In_1369);
nand U642 (N_642,In_2341,In_2202);
nor U643 (N_643,In_1099,In_1598);
nand U644 (N_644,In_188,In_590);
nor U645 (N_645,In_1176,In_2306);
xnor U646 (N_646,In_458,In_459);
and U647 (N_647,In_1864,In_215);
nor U648 (N_648,In_963,In_2332);
or U649 (N_649,In_1211,In_1694);
or U650 (N_650,In_625,In_1644);
or U651 (N_651,In_514,In_2465);
nor U652 (N_652,In_540,In_1717);
and U653 (N_653,In_361,In_326);
and U654 (N_654,In_1514,In_442);
nand U655 (N_655,In_1994,In_8);
and U656 (N_656,In_1972,In_1879);
nand U657 (N_657,In_318,In_2382);
or U658 (N_658,In_1190,In_1873);
nand U659 (N_659,In_1002,In_1019);
and U660 (N_660,In_1863,In_1529);
nand U661 (N_661,In_2424,In_2221);
or U662 (N_662,In_119,In_635);
xnor U663 (N_663,In_2211,In_1397);
nor U664 (N_664,In_1874,In_323);
xnor U665 (N_665,In_366,In_649);
nor U666 (N_666,In_1619,In_1507);
and U667 (N_667,In_1189,In_1075);
nor U668 (N_668,In_1105,In_737);
or U669 (N_669,In_801,In_32);
xnor U670 (N_670,In_1092,In_1652);
or U671 (N_671,In_1456,In_742);
or U672 (N_672,In_1153,In_2479);
nor U673 (N_673,In_1443,In_639);
nor U674 (N_674,In_714,In_616);
xnor U675 (N_675,In_40,In_574);
and U676 (N_676,In_543,In_427);
xnor U677 (N_677,In_2493,In_960);
or U678 (N_678,In_191,In_1025);
nand U679 (N_679,In_689,In_2400);
xor U680 (N_680,In_633,In_1341);
or U681 (N_681,In_284,In_2397);
nor U682 (N_682,In_1474,In_1838);
or U683 (N_683,In_636,In_1229);
nor U684 (N_684,In_1655,In_2312);
nand U685 (N_685,In_1253,In_2447);
nor U686 (N_686,In_961,In_129);
and U687 (N_687,In_1018,In_1114);
nor U688 (N_688,In_1454,In_1367);
and U689 (N_689,In_262,In_707);
nor U690 (N_690,In_2391,In_248);
xor U691 (N_691,In_1587,In_1469);
xor U692 (N_692,In_2001,In_958);
or U693 (N_693,In_1920,In_1318);
nor U694 (N_694,In_508,In_19);
xor U695 (N_695,In_1662,In_1985);
nand U696 (N_696,In_2357,In_1054);
nand U697 (N_697,In_1425,In_1760);
and U698 (N_698,In_874,In_2116);
xor U699 (N_699,In_1446,In_1252);
and U700 (N_700,In_1482,In_1134);
nand U701 (N_701,In_2410,In_2259);
xor U702 (N_702,In_667,In_2161);
and U703 (N_703,In_1390,In_2363);
nor U704 (N_704,In_530,In_580);
xor U705 (N_705,In_710,In_2187);
and U706 (N_706,In_2230,In_202);
nor U707 (N_707,In_2421,In_815);
or U708 (N_708,In_657,In_748);
nor U709 (N_709,In_666,In_866);
and U710 (N_710,In_2333,In_2186);
or U711 (N_711,In_2160,In_1943);
nor U712 (N_712,In_52,In_155);
xnor U713 (N_713,In_615,In_2090);
nand U714 (N_714,In_1533,In_466);
xor U715 (N_715,In_468,In_2040);
nand U716 (N_716,In_1498,In_311);
and U717 (N_717,In_337,In_1100);
xnor U718 (N_718,In_426,In_1043);
and U719 (N_719,In_357,In_440);
xor U720 (N_720,In_2260,In_73);
or U721 (N_721,In_1074,In_1334);
or U722 (N_722,In_834,In_355);
and U723 (N_723,In_1257,In_1919);
and U724 (N_724,In_943,In_781);
and U725 (N_725,In_1286,In_761);
xnor U726 (N_726,In_2372,In_671);
xor U727 (N_727,In_1739,In_448);
xor U728 (N_728,In_891,In_1280);
nand U729 (N_729,In_239,In_1808);
nor U730 (N_730,In_1726,In_1207);
xnor U731 (N_731,In_1141,In_1068);
nor U732 (N_732,In_2227,In_2407);
nand U733 (N_733,In_1221,In_2309);
or U734 (N_734,In_1552,In_482);
nand U735 (N_735,In_307,In_1682);
nor U736 (N_736,In_61,In_137);
and U737 (N_737,In_821,In_1175);
nand U738 (N_738,In_1338,In_1067);
nor U739 (N_739,In_75,In_1613);
nand U740 (N_740,In_2147,In_555);
nand U741 (N_741,In_2109,In_2065);
nand U742 (N_742,In_906,In_1011);
and U743 (N_743,In_890,In_836);
and U744 (N_744,In_1953,In_1204);
or U745 (N_745,In_451,In_1620);
nor U746 (N_746,In_1023,In_359);
or U747 (N_747,In_1375,In_938);
xor U748 (N_748,In_571,In_1634);
xnor U749 (N_749,In_1775,In_1650);
xor U750 (N_750,In_1158,In_471);
nor U751 (N_751,In_2017,In_2343);
nand U752 (N_752,In_2282,In_378);
nand U753 (N_753,In_1262,In_1051);
nor U754 (N_754,In_1442,In_1947);
and U755 (N_755,In_1301,In_541);
nor U756 (N_756,In_179,In_250);
or U757 (N_757,In_136,In_42);
nand U758 (N_758,In_1875,In_1161);
or U759 (N_759,In_1431,In_619);
or U760 (N_760,In_1140,In_54);
nor U761 (N_761,In_2204,In_446);
and U762 (N_762,In_2167,In_1121);
or U763 (N_763,In_2193,In_2336);
or U764 (N_764,In_2198,In_997);
and U765 (N_765,In_2214,In_919);
xor U766 (N_766,In_1438,In_1778);
nand U767 (N_767,In_2097,In_1568);
nor U768 (N_768,In_827,In_1241);
and U769 (N_769,In_405,In_16);
nand U770 (N_770,In_210,In_759);
nand U771 (N_771,In_2072,In_1609);
nand U772 (N_772,In_1734,In_277);
nand U773 (N_773,In_2275,In_2236);
or U774 (N_774,In_1500,In_375);
or U775 (N_775,In_1883,In_123);
nor U776 (N_776,In_1179,In_1127);
nor U777 (N_777,In_328,In_706);
xnor U778 (N_778,In_1213,In_2296);
xor U779 (N_779,In_256,In_2257);
and U780 (N_780,In_904,In_1326);
or U781 (N_781,In_1317,In_2188);
nand U782 (N_782,In_1936,In_1781);
nand U783 (N_783,In_996,In_1639);
and U784 (N_784,In_792,In_1711);
nand U785 (N_785,In_1230,In_718);
and U786 (N_786,In_932,In_1534);
and U787 (N_787,In_1956,In_1546);
nor U788 (N_788,In_1907,In_2163);
xor U789 (N_789,In_2093,In_685);
or U790 (N_790,In_991,In_2007);
and U791 (N_791,In_1790,In_1820);
nor U792 (N_792,In_362,In_2322);
or U793 (N_793,In_2381,In_1754);
nor U794 (N_794,In_2277,In_726);
or U795 (N_795,In_776,In_1148);
or U796 (N_796,In_1419,In_1842);
and U797 (N_797,In_1826,In_517);
or U798 (N_798,In_1950,In_1733);
xnor U799 (N_799,In_987,In_253);
xor U800 (N_800,In_697,In_2290);
or U801 (N_801,In_1149,In_1302);
and U802 (N_802,In_1859,In_2062);
and U803 (N_803,In_1715,In_1926);
and U804 (N_804,In_538,In_610);
xnor U805 (N_805,In_2225,In_1082);
and U806 (N_806,In_711,In_1833);
and U807 (N_807,In_2076,In_2359);
xnor U808 (N_808,In_2426,In_867);
nor U809 (N_809,In_1060,In_2131);
xor U810 (N_810,In_1091,In_2392);
nor U811 (N_811,In_1282,In_1743);
nand U812 (N_812,In_1240,In_794);
and U813 (N_813,In_930,In_1511);
and U814 (N_814,In_2215,In_708);
xnor U815 (N_815,In_807,In_651);
xnor U816 (N_816,In_2349,In_2039);
nand U817 (N_817,In_2067,In_1421);
or U818 (N_818,In_800,In_1289);
xor U819 (N_819,In_1095,In_1394);
and U820 (N_820,In_999,In_388);
nor U821 (N_821,In_1359,In_1785);
nor U822 (N_822,In_1362,In_658);
nor U823 (N_823,In_1666,In_542);
xnor U824 (N_824,In_356,In_1722);
nand U825 (N_825,In_2080,In_2287);
xnor U826 (N_826,In_1865,In_1696);
nand U827 (N_827,In_163,In_229);
nor U828 (N_828,In_28,In_1388);
or U829 (N_829,In_1938,In_1591);
nor U830 (N_830,In_80,In_2461);
nand U831 (N_831,In_14,In_1699);
or U832 (N_832,In_1735,In_2380);
nor U833 (N_833,In_1937,In_1260);
and U834 (N_834,In_826,In_110);
or U835 (N_835,In_268,In_1172);
nor U836 (N_836,In_2233,In_2112);
xnor U837 (N_837,In_293,In_1671);
and U838 (N_838,In_2373,In_1802);
nand U839 (N_839,In_430,In_977);
nand U840 (N_840,In_1215,In_1930);
nor U841 (N_841,In_457,In_380);
nand U842 (N_842,In_1001,In_26);
nand U843 (N_843,In_2272,In_1382);
xor U844 (N_844,In_1486,In_1817);
or U845 (N_845,In_2472,In_5);
nor U846 (N_846,In_476,In_1303);
xnor U847 (N_847,In_2482,In_735);
xor U848 (N_848,In_1353,In_1967);
nor U849 (N_849,In_2182,In_2473);
or U850 (N_850,In_793,In_973);
nor U851 (N_851,In_1825,In_533);
xor U852 (N_852,In_1407,In_2353);
nand U853 (N_853,In_912,In_1004);
nor U854 (N_854,In_453,In_24);
or U855 (N_855,In_417,In_121);
nor U856 (N_856,In_2390,In_1402);
nor U857 (N_857,In_2337,In_2079);
xor U858 (N_858,In_425,In_1163);
xor U859 (N_859,In_350,In_825);
nor U860 (N_860,In_274,In_2055);
and U861 (N_861,In_2085,In_2241);
nand U862 (N_862,In_1801,In_2178);
and U863 (N_863,In_1028,In_1681);
xnor U864 (N_864,In_2469,In_2393);
xnor U865 (N_865,In_2238,In_1126);
or U866 (N_866,In_1447,In_1906);
nand U867 (N_867,In_390,In_299);
nor U868 (N_868,In_1660,In_2054);
or U869 (N_869,In_2301,In_1703);
nand U870 (N_870,In_1784,In_1993);
and U871 (N_871,In_383,In_2325);
and U872 (N_872,In_1599,In_790);
nand U873 (N_873,In_2340,In_263);
nand U874 (N_874,In_142,In_168);
nand U875 (N_875,In_2051,In_603);
or U876 (N_876,In_1506,In_255);
or U877 (N_877,In_2050,In_1663);
xor U878 (N_878,In_1199,In_687);
and U879 (N_879,In_1259,In_1457);
xnor U880 (N_880,In_1494,In_346);
xnor U881 (N_881,In_1737,In_1538);
or U882 (N_882,In_700,In_2318);
nand U883 (N_883,In_630,In_1548);
nand U884 (N_884,In_39,In_637);
or U885 (N_885,In_2213,In_864);
nor U886 (N_886,In_1006,In_520);
and U887 (N_887,In_893,In_385);
nor U888 (N_888,In_2154,In_918);
nor U889 (N_889,In_1799,In_1992);
or U890 (N_890,In_1170,In_2166);
nor U891 (N_891,In_1423,In_1850);
xor U892 (N_892,In_70,In_485);
nand U893 (N_893,In_1464,In_18);
xnor U894 (N_894,In_1238,In_774);
or U895 (N_895,In_1355,In_1977);
nand U896 (N_896,In_779,In_1724);
nor U897 (N_897,In_1467,In_935);
nand U898 (N_898,In_1094,In_441);
nand U899 (N_899,In_145,In_497);
nand U900 (N_900,In_146,In_756);
nand U901 (N_901,In_2442,In_2164);
xor U902 (N_902,In_1798,In_1558);
xnor U903 (N_903,In_733,In_760);
nor U904 (N_904,In_1626,In_1344);
or U905 (N_905,In_1794,In_1115);
and U906 (N_906,In_1078,In_694);
and U907 (N_907,In_1805,In_118);
or U908 (N_908,In_1261,In_2058);
xor U909 (N_909,In_1603,In_1767);
or U910 (N_910,In_550,In_522);
nor U911 (N_911,In_382,In_1549);
or U912 (N_912,In_1079,In_1744);
and U913 (N_913,In_1323,In_531);
and U914 (N_914,In_613,In_1819);
xor U915 (N_915,In_2078,In_512);
nand U916 (N_916,In_539,In_1222);
xor U917 (N_917,In_2185,In_1208);
nor U918 (N_918,In_2351,In_213);
and U919 (N_919,In_2023,In_1618);
nor U920 (N_920,In_1806,In_504);
or U921 (N_921,In_1296,In_1881);
or U922 (N_922,In_2126,In_1110);
or U923 (N_923,In_1458,In_1610);
xor U924 (N_924,In_678,In_570);
or U925 (N_925,In_724,In_1965);
or U926 (N_926,In_434,In_1946);
or U927 (N_927,In_1265,In_2304);
xor U928 (N_928,In_1125,In_2136);
nand U929 (N_929,In_1187,In_2437);
xnor U930 (N_930,In_1408,In_819);
nand U931 (N_931,In_2319,In_1984);
and U932 (N_932,In_1123,In_1488);
nand U933 (N_933,In_988,In_1537);
xnor U934 (N_934,In_2120,In_169);
nand U935 (N_935,In_579,In_2228);
or U936 (N_936,In_2440,In_159);
xnor U937 (N_937,In_525,In_1658);
and U938 (N_938,In_2140,In_1772);
xor U939 (N_939,In_1409,In_1313);
xor U940 (N_940,In_2018,In_1331);
nand U941 (N_941,In_1281,In_2303);
and U942 (N_942,In_154,In_862);
xor U943 (N_943,In_369,In_1084);
nor U944 (N_944,In_648,In_1184);
nand U945 (N_945,In_372,In_1422);
or U946 (N_946,In_254,In_1271);
nor U947 (N_947,In_1295,In_1165);
nor U948 (N_948,In_1147,In_2488);
or U949 (N_949,In_2295,In_879);
xnor U950 (N_950,In_1771,In_2307);
or U951 (N_951,In_444,In_232);
nand U952 (N_952,In_461,In_1234);
or U953 (N_953,In_2183,In_670);
and U954 (N_954,In_1706,In_285);
nand U955 (N_955,In_799,In_1346);
nand U956 (N_956,In_2298,In_2499);
xor U957 (N_957,In_2386,In_1616);
xor U958 (N_958,In_363,In_2132);
nand U959 (N_959,In_1299,In_1374);
xor U960 (N_960,In_2374,In_1831);
or U961 (N_961,In_1239,In_674);
nor U962 (N_962,In_43,In_72);
or U963 (N_963,In_847,In_2143);
and U964 (N_964,In_2485,In_1876);
or U965 (N_965,In_456,In_1997);
xnor U966 (N_966,In_2434,In_928);
xnor U967 (N_967,In_2087,In_1440);
nor U968 (N_968,In_970,In_892);
xor U969 (N_969,In_1894,In_784);
nand U970 (N_970,In_526,In_2212);
nor U971 (N_971,In_423,In_1927);
and U972 (N_972,In_959,In_1366);
xnor U973 (N_973,In_679,In_951);
xnor U974 (N_974,In_606,In_1154);
nor U975 (N_975,In_2299,In_2158);
or U976 (N_976,In_1162,In_394);
nand U977 (N_977,In_1046,In_1902);
nor U978 (N_978,In_2314,In_1357);
nand U979 (N_979,In_1637,In_1050);
xnor U980 (N_980,In_1676,In_1543);
or U981 (N_981,In_1370,In_805);
nand U982 (N_982,In_314,In_1614);
and U983 (N_983,In_660,In_824);
xnor U984 (N_984,In_258,In_1664);
nand U985 (N_985,In_55,In_557);
nor U986 (N_986,In_599,In_392);
nor U987 (N_987,In_1759,In_1522);
nand U988 (N_988,In_683,In_2114);
or U989 (N_989,In_2481,In_376);
and U990 (N_990,In_162,In_1945);
or U991 (N_991,In_810,In_1452);
nand U992 (N_992,In_1752,In_1070);
or U993 (N_993,In_2032,In_1320);
nand U994 (N_994,In_1427,In_1167);
xor U995 (N_995,In_261,In_1356);
or U996 (N_996,In_967,In_2347);
xnor U997 (N_997,In_1139,In_2100);
or U998 (N_998,In_1404,In_1780);
or U999 (N_999,In_1695,In_511);
and U1000 (N_1000,N_723,N_238);
nand U1001 (N_1001,N_272,N_746);
or U1002 (N_1002,N_806,N_972);
nand U1003 (N_1003,N_741,In_1380);
and U1004 (N_1004,In_553,N_792);
xnor U1005 (N_1005,In_2495,In_486);
or U1006 (N_1006,N_784,N_451);
nand U1007 (N_1007,In_2478,N_671);
nor U1008 (N_1008,N_79,N_404);
xnor U1009 (N_1009,In_374,In_1485);
nand U1010 (N_1010,N_729,N_832);
and U1011 (N_1011,N_433,N_656);
nand U1012 (N_1012,N_481,N_26);
or U1013 (N_1013,N_688,N_253);
xor U1014 (N_1014,In_654,N_10);
xnor U1015 (N_1015,N_733,N_651);
nor U1016 (N_1016,N_391,In_106);
xor U1017 (N_1017,In_2328,N_944);
nor U1018 (N_1018,N_181,N_726);
nor U1019 (N_1019,In_252,In_189);
or U1020 (N_1020,N_340,In_164);
and U1021 (N_1021,N_672,N_948);
nand U1022 (N_1022,N_380,In_171);
nand U1023 (N_1023,In_865,N_157);
nor U1024 (N_1024,N_587,N_809);
and U1025 (N_1025,N_366,In_2468);
xnor U1026 (N_1026,In_1138,N_660);
nand U1027 (N_1027,N_631,N_943);
nand U1028 (N_1028,N_782,N_215);
and U1029 (N_1029,N_425,N_102);
or U1030 (N_1030,N_153,N_146);
nand U1031 (N_1031,N_740,N_622);
nand U1032 (N_1032,In_2444,In_58);
nand U1033 (N_1033,In_2176,N_21);
and U1034 (N_1034,N_402,N_713);
and U1035 (N_1035,N_158,N_178);
xnor U1036 (N_1036,N_675,In_115);
or U1037 (N_1037,N_844,N_930);
and U1038 (N_1038,In_782,N_632);
and U1039 (N_1039,In_1329,N_820);
or U1040 (N_1040,N_498,In_524);
nor U1041 (N_1041,In_880,In_365);
or U1042 (N_1042,In_2476,N_896);
xnor U1043 (N_1043,N_544,N_296);
nand U1044 (N_1044,N_104,N_160);
or U1045 (N_1045,In_2251,In_841);
nand U1046 (N_1046,In_740,N_35);
or U1047 (N_1047,In_206,N_327);
xnor U1048 (N_1048,In_2377,N_322);
or U1049 (N_1049,In_2239,N_356);
and U1050 (N_1050,In_1586,N_696);
nor U1051 (N_1051,N_423,In_1899);
xnor U1052 (N_1052,N_411,N_773);
xor U1053 (N_1053,N_502,In_2105);
and U1054 (N_1054,N_505,N_543);
nand U1055 (N_1055,In_2237,N_879);
or U1056 (N_1056,N_791,In_1347);
or U1057 (N_1057,N_432,N_250);
xor U1058 (N_1058,In_1536,N_332);
and U1059 (N_1059,N_856,N_550);
nand U1060 (N_1060,N_644,In_103);
xor U1061 (N_1061,In_833,In_1314);
nor U1062 (N_1062,N_911,In_2216);
nor U1063 (N_1063,N_576,N_197);
nand U1064 (N_1064,N_396,N_574);
or U1065 (N_1065,In_1796,In_2246);
nand U1066 (N_1066,N_647,N_292);
and U1067 (N_1067,In_1570,N_570);
nand U1068 (N_1068,N_428,In_1779);
or U1069 (N_1069,In_181,In_712);
xor U1070 (N_1070,In_2269,N_617);
and U1071 (N_1071,In_1195,In_1991);
or U1072 (N_1072,N_539,N_129);
nand U1073 (N_1073,In_739,N_825);
and U1074 (N_1074,In_126,N_285);
nor U1075 (N_1075,In_1757,In_316);
nor U1076 (N_1076,N_232,In_1764);
nor U1077 (N_1077,N_616,N_567);
and U1078 (N_1078,N_722,In_294);
nor U1079 (N_1079,N_184,In_10);
or U1080 (N_1080,N_41,N_368);
or U1081 (N_1081,N_922,In_1016);
xnor U1082 (N_1082,N_989,N_932);
or U1083 (N_1083,N_66,N_552);
nand U1084 (N_1084,In_1417,N_348);
nand U1085 (N_1085,In_2441,N_143);
nand U1086 (N_1086,N_707,In_2073);
and U1087 (N_1087,N_492,N_698);
nor U1088 (N_1088,N_601,N_863);
nor U1089 (N_1089,N_152,N_970);
or U1090 (N_1090,N_881,N_662);
or U1091 (N_1091,In_2005,N_486);
nor U1092 (N_1092,In_1061,In_656);
xnor U1093 (N_1093,In_2367,N_287);
xor U1094 (N_1094,In_302,In_1567);
xnor U1095 (N_1095,N_277,In_528);
nor U1096 (N_1096,N_360,N_256);
nand U1097 (N_1097,N_284,N_86);
and U1098 (N_1098,N_816,In_17);
or U1099 (N_1099,In_170,N_845);
and U1100 (N_1100,N_923,N_390);
or U1101 (N_1101,N_935,N_27);
nor U1102 (N_1102,N_997,N_37);
and U1103 (N_1103,In_222,In_2429);
nor U1104 (N_1104,N_446,In_1173);
nand U1105 (N_1105,In_1330,In_1000);
and U1106 (N_1106,N_293,In_1673);
xnor U1107 (N_1107,N_745,N_47);
nor U1108 (N_1108,In_178,In_1276);
nand U1109 (N_1109,N_497,In_1297);
and U1110 (N_1110,N_780,N_11);
nand U1111 (N_1111,N_835,In_2196);
and U1112 (N_1112,In_889,N_925);
and U1113 (N_1113,N_615,In_116);
and U1114 (N_1114,In_2046,N_951);
xnor U1115 (N_1115,In_238,N_589);
xnor U1116 (N_1116,N_799,In_301);
nand U1117 (N_1117,N_53,N_788);
and U1118 (N_1118,N_610,N_639);
and U1119 (N_1119,N_134,In_1547);
and U1120 (N_1120,N_68,N_509);
or U1121 (N_1121,N_165,N_595);
and U1122 (N_1122,N_224,N_394);
or U1123 (N_1123,N_633,N_657);
and U1124 (N_1124,In_818,In_2409);
nor U1125 (N_1125,In_2111,N_233);
xor U1126 (N_1126,In_1561,In_1077);
nand U1127 (N_1127,N_493,N_841);
nand U1128 (N_1128,N_702,In_1122);
nor U1129 (N_1129,N_538,N_359);
nand U1130 (N_1130,N_251,In_1080);
and U1131 (N_1131,In_1816,N_483);
or U1132 (N_1132,In_978,In_1527);
and U1133 (N_1133,N_371,N_525);
and U1134 (N_1134,N_674,In_1582);
nand U1135 (N_1135,In_1595,N_420);
nand U1136 (N_1136,N_96,In_368);
nor U1137 (N_1137,N_161,In_1178);
nor U1138 (N_1138,N_887,N_114);
xor U1139 (N_1139,N_936,In_2110);
nand U1140 (N_1140,N_122,In_1745);
and U1141 (N_1141,In_1479,N_97);
and U1142 (N_1142,N_870,N_728);
and U1143 (N_1143,In_1093,N_926);
nor U1144 (N_1144,In_125,N_758);
xor U1145 (N_1145,In_2192,N_455);
xor U1146 (N_1146,N_223,N_938);
and U1147 (N_1147,N_80,N_400);
nand U1148 (N_1148,N_915,In_1156);
and U1149 (N_1149,In_717,In_2384);
nand U1150 (N_1150,N_584,In_1196);
nand U1151 (N_1151,N_704,In_475);
nor U1152 (N_1152,N_372,N_210);
nand U1153 (N_1153,N_630,In_1585);
or U1154 (N_1154,N_376,N_629);
nand U1155 (N_1155,N_826,In_1444);
or U1156 (N_1156,N_81,N_257);
nor U1157 (N_1157,N_973,N_515);
and U1158 (N_1158,N_450,N_456);
nor U1159 (N_1159,N_494,N_761);
nand U1160 (N_1160,In_1186,N_770);
and U1161 (N_1161,In_994,In_389);
nand U1162 (N_1162,In_1398,In_149);
and U1163 (N_1163,N_818,N_326);
or U1164 (N_1164,N_939,In_1206);
and U1165 (N_1165,N_408,In_182);
nand U1166 (N_1166,In_593,N_488);
xor U1167 (N_1167,N_513,N_140);
or U1168 (N_1168,N_439,N_979);
and U1169 (N_1169,In_2350,In_1277);
xor U1170 (N_1170,N_171,N_619);
or U1171 (N_1171,In_2281,N_363);
xnor U1172 (N_1172,In_386,In_138);
xnor U1173 (N_1173,In_795,N_849);
or U1174 (N_1174,N_899,N_987);
nand U1175 (N_1175,In_796,In_676);
nor U1176 (N_1176,N_294,N_377);
and U1177 (N_1177,In_1066,N_185);
xnor U1178 (N_1178,N_649,N_801);
nor U1179 (N_1179,In_411,In_1504);
xor U1180 (N_1180,N_149,In_1124);
nand U1181 (N_1181,N_523,In_2020);
and U1182 (N_1182,N_785,N_325);
nor U1183 (N_1183,N_247,N_201);
and U1184 (N_1184,N_789,N_116);
xor U1185 (N_1185,N_154,N_229);
xnor U1186 (N_1186,In_565,N_136);
nor U1187 (N_1187,N_222,N_519);
xor U1188 (N_1188,In_523,In_492);
and U1189 (N_1189,N_869,In_2122);
xnor U1190 (N_1190,N_274,In_965);
nor U1191 (N_1191,In_1955,N_207);
xor U1192 (N_1192,In_2008,In_1311);
xnor U1193 (N_1193,N_435,N_169);
xnor U1194 (N_1194,In_535,N_243);
or U1195 (N_1195,N_125,N_33);
xnor U1196 (N_1196,N_388,In_778);
and U1197 (N_1197,N_182,In_2456);
or U1198 (N_1198,N_686,N_307);
and U1199 (N_1199,In_1958,N_941);
nand U1200 (N_1200,N_349,N_280);
and U1201 (N_1201,N_661,N_517);
nand U1202 (N_1202,N_967,In_2027);
nor U1203 (N_1203,N_51,N_861);
or U1204 (N_1204,N_974,In_536);
xnor U1205 (N_1205,N_858,N_600);
xnor U1206 (N_1206,N_638,N_771);
and U1207 (N_1207,N_405,N_429);
nand U1208 (N_1208,In_2184,In_1430);
nor U1209 (N_1209,N_984,N_495);
xor U1210 (N_1210,In_1871,N_817);
and U1211 (N_1211,In_2258,N_769);
nor U1212 (N_1212,N_751,N_426);
or U1213 (N_1213,N_996,In_1505);
or U1214 (N_1214,In_617,N_605);
and U1215 (N_1215,N_95,N_252);
nor U1216 (N_1216,N_555,In_1862);
xor U1217 (N_1217,N_399,N_353);
xnor U1218 (N_1218,N_673,N_444);
xnor U1219 (N_1219,In_272,N_15);
and U1220 (N_1220,N_957,N_314);
nor U1221 (N_1221,N_995,N_38);
and U1222 (N_1222,N_442,N_655);
nand U1223 (N_1223,In_45,N_553);
xnor U1224 (N_1224,N_437,In_519);
xnor U1225 (N_1225,In_1758,N_109);
nand U1226 (N_1226,N_897,N_760);
nand U1227 (N_1227,N_940,N_298);
nand U1228 (N_1228,In_1935,N_705);
xor U1229 (N_1229,In_393,N_46);
xnor U1230 (N_1230,N_738,In_403);
xor U1231 (N_1231,In_1354,In_57);
nand U1232 (N_1232,In_822,In_455);
and U1233 (N_1233,In_152,N_60);
and U1234 (N_1234,N_981,N_663);
and U1235 (N_1235,N_963,In_1342);
xor U1236 (N_1236,N_375,N_504);
and U1237 (N_1237,In_652,N_381);
nand U1238 (N_1238,N_275,N_39);
and U1239 (N_1239,N_626,In_702);
nand U1240 (N_1240,N_88,In_1244);
nand U1241 (N_1241,N_802,N_591);
or U1242 (N_1242,N_346,N_755);
or U1243 (N_1243,N_568,In_2358);
nor U1244 (N_1244,In_1705,N_781);
xor U1245 (N_1245,N_373,N_540);
nor U1246 (N_1246,N_397,N_150);
xnor U1247 (N_1247,N_711,N_886);
nor U1248 (N_1248,In_1212,N_918);
and U1249 (N_1249,N_378,In_320);
nand U1250 (N_1250,N_588,In_1275);
nand U1251 (N_1251,N_531,N_482);
xor U1252 (N_1252,N_883,N_333);
xor U1253 (N_1253,N_775,In_319);
xor U1254 (N_1254,N_2,N_586);
nand U1255 (N_1255,N_447,In_1183);
or U1256 (N_1256,N_934,N_205);
nand U1257 (N_1257,N_72,N_441);
xor U1258 (N_1258,N_246,N_106);
or U1259 (N_1259,N_13,In_495);
or U1260 (N_1260,N_94,N_828);
nor U1261 (N_1261,N_34,In_2489);
and U1262 (N_1262,N_703,N_288);
or U1263 (N_1263,In_2317,In_422);
nand U1264 (N_1264,N_283,N_436);
and U1265 (N_1265,N_848,N_131);
nor U1266 (N_1266,N_575,N_716);
or U1267 (N_1267,N_484,In_402);
xor U1268 (N_1268,In_1765,N_542);
or U1269 (N_1269,N_19,In_2255);
nor U1270 (N_1270,N_6,N_225);
xnor U1271 (N_1271,In_843,N_947);
nor U1272 (N_1272,N_850,N_392);
nor U1273 (N_1273,N_565,N_652);
and U1274 (N_1274,N_459,N_566);
and U1275 (N_1275,N_29,N_458);
or U1276 (N_1276,N_236,In_1964);
xor U1277 (N_1277,In_2189,In_2276);
xor U1278 (N_1278,N_964,N_212);
nor U1279 (N_1279,In_1205,N_58);
nor U1280 (N_1280,N_884,N_216);
or U1281 (N_1281,In_2156,N_401);
xnor U1282 (N_1282,In_876,N_263);
nor U1283 (N_1283,N_862,N_524);
xnor U1284 (N_1284,N_101,N_689);
nand U1285 (N_1285,In_582,N_260);
or U1286 (N_1286,In_1233,N_190);
or U1287 (N_1287,N_49,N_648);
nor U1288 (N_1288,N_815,In_2);
and U1289 (N_1289,N_119,In_1854);
nand U1290 (N_1290,N_724,N_365);
xor U1291 (N_1291,In_537,N_4);
nand U1292 (N_1292,In_1851,N_231);
nand U1293 (N_1293,N_434,N_621);
nand U1294 (N_1294,N_339,In_499);
nor U1295 (N_1295,In_68,N_100);
xnor U1296 (N_1296,N_228,N_514);
nor U1297 (N_1297,In_990,In_741);
nand U1298 (N_1298,N_627,In_1843);
xor U1299 (N_1299,N_659,In_1034);
and U1300 (N_1300,N_699,N_961);
xnor U1301 (N_1301,N_593,N_457);
nor U1302 (N_1302,N_511,N_344);
or U1303 (N_1303,In_347,N_779);
and U1304 (N_1304,N_70,N_440);
nand U1305 (N_1305,In_41,In_1674);
nand U1306 (N_1306,In_198,N_170);
xnor U1307 (N_1307,In_1026,N_308);
or U1308 (N_1308,N_20,N_628);
and U1309 (N_1309,N_547,N_491);
nor U1310 (N_1310,In_338,N_103);
nor U1311 (N_1311,N_798,N_842);
xnor U1312 (N_1312,N_237,In_731);
nor U1313 (N_1313,N_537,In_1008);
nor U1314 (N_1314,N_521,In_1858);
or U1315 (N_1315,N_868,N_692);
and U1316 (N_1316,N_904,In_1713);
nor U1317 (N_1317,In_758,N_144);
nand U1318 (N_1318,In_1157,In_984);
and U1319 (N_1319,N_234,N_120);
or U1320 (N_1320,N_355,N_3);
and U1321 (N_1321,N_919,N_199);
or U1322 (N_1322,In_1914,In_1688);
or U1323 (N_1323,N_151,N_126);
xor U1324 (N_1324,N_966,N_187);
nand U1325 (N_1325,N_445,N_893);
xnor U1326 (N_1326,In_1024,In_1602);
nor U1327 (N_1327,N_874,N_16);
or U1328 (N_1328,In_983,N_410);
or U1329 (N_1329,N_334,N_343);
or U1330 (N_1330,N_814,N_727);
or U1331 (N_1331,N_917,N_73);
nand U1332 (N_1332,N_267,N_752);
and U1333 (N_1333,N_955,In_1731);
and U1334 (N_1334,In_614,N_976);
or U1335 (N_1335,N_937,N_315);
nand U1336 (N_1336,N_138,N_369);
or U1337 (N_1337,N_324,In_786);
nand U1338 (N_1338,N_522,N_685);
nand U1339 (N_1339,N_44,N_737);
or U1340 (N_1340,In_2462,N_331);
and U1341 (N_1341,In_835,N_526);
nor U1342 (N_1342,N_290,N_577);
and U1343 (N_1343,N_192,In_353);
and U1344 (N_1344,N_916,N_510);
nand U1345 (N_1345,N_12,In_33);
nor U1346 (N_1346,N_200,In_2063);
or U1347 (N_1347,N_110,In_626);
nor U1348 (N_1348,N_330,In_2229);
or U1349 (N_1349,N_508,N_777);
xor U1350 (N_1350,N_579,N_969);
nor U1351 (N_1351,In_972,N_419);
and U1352 (N_1352,In_2394,N_905);
or U1353 (N_1353,N_452,N_730);
nor U1354 (N_1354,N_262,N_894);
and U1355 (N_1355,N_921,N_877);
and U1356 (N_1356,N_407,N_808);
or U1357 (N_1357,N_599,N_65);
and U1358 (N_1358,In_2037,In_950);
nor U1359 (N_1359,In_1911,N_393);
and U1360 (N_1360,N_487,N_634);
xnor U1361 (N_1361,In_602,N_9);
or U1362 (N_1362,N_762,N_352);
nand U1363 (N_1363,In_1513,In_915);
and U1364 (N_1364,N_248,N_564);
xor U1365 (N_1365,N_846,In_2107);
nand U1366 (N_1366,N_906,In_1913);
or U1367 (N_1367,In_809,N_83);
xnor U1368 (N_1368,N_875,N_978);
nor U1369 (N_1369,N_183,N_56);
nor U1370 (N_1370,In_1689,N_281);
and U1371 (N_1371,N_30,N_317);
or U1372 (N_1372,In_2379,N_168);
nand U1373 (N_1373,N_807,In_1968);
nand U1374 (N_1374,N_971,N_313);
xnor U1375 (N_1375,N_335,In_989);
xor U1376 (N_1376,In_2388,N_147);
and U1377 (N_1377,N_694,In_2463);
and U1378 (N_1378,N_383,N_173);
or U1379 (N_1379,N_350,N_121);
nand U1380 (N_1380,In_791,N_195);
or U1381 (N_1381,N_471,N_186);
nand U1382 (N_1382,N_571,In_1606);
xor U1383 (N_1383,In_317,N_795);
or U1384 (N_1384,N_929,N_611);
or U1385 (N_1385,N_443,In_607);
nand U1386 (N_1386,In_752,In_1371);
or U1387 (N_1387,N_982,N_8);
or U1388 (N_1388,N_603,In_1989);
and U1389 (N_1389,In_1429,N_562);
nand U1390 (N_1390,N_912,N_778);
or U1391 (N_1391,N_871,N_988);
and U1392 (N_1392,N_466,N_913);
and U1393 (N_1393,N_189,N_836);
nand U1394 (N_1394,N_202,N_908);
or U1395 (N_1395,In_242,N_286);
nor U1396 (N_1396,In_341,N_145);
nand U1397 (N_1397,In_1324,In_898);
and U1398 (N_1398,N_624,N_362);
nand U1399 (N_1399,N_227,N_266);
nor U1400 (N_1400,In_2060,N_596);
xnor U1401 (N_1401,N_889,In_788);
or U1402 (N_1402,N_255,N_361);
nand U1403 (N_1403,In_551,N_54);
xor U1404 (N_1404,N_677,N_418);
or U1405 (N_1405,N_880,In_406);
nand U1406 (N_1406,N_759,In_2082);
nand U1407 (N_1407,N_635,N_99);
nand U1408 (N_1408,N_142,N_316);
nor U1409 (N_1409,N_91,In_1857);
and U1410 (N_1410,N_975,N_833);
or U1411 (N_1411,N_774,N_693);
nor U1412 (N_1412,N_289,In_1266);
and U1413 (N_1413,N_386,N_357);
and U1414 (N_1414,In_910,N_787);
nor U1415 (N_1415,In_1335,N_750);
xnor U1416 (N_1416,N_36,N_318);
or U1417 (N_1417,N_474,N_460);
xnor U1418 (N_1418,N_319,N_614);
or U1419 (N_1419,N_827,N_958);
nor U1420 (N_1420,In_2106,N_715);
or U1421 (N_1421,In_1596,N_415);
nand U1422 (N_1422,N_953,N_276);
and U1423 (N_1423,N_665,N_690);
xor U1424 (N_1424,N_753,N_900);
and U1425 (N_1425,In_1751,In_296);
and U1426 (N_1426,In_245,In_1306);
and U1427 (N_1427,In_1822,N_107);
xnor U1428 (N_1428,N_123,In_560);
nor U1429 (N_1429,N_48,In_3);
or U1430 (N_1430,N_530,In_1611);
xnor U1431 (N_1431,N_668,N_811);
nor U1432 (N_1432,In_2316,N_563);
nand U1433 (N_1433,N_977,N_839);
xor U1434 (N_1434,N_669,In_573);
and U1435 (N_1435,N_909,N_336);
nor U1436 (N_1436,N_559,In_2346);
xor U1437 (N_1437,N_329,N_613);
and U1438 (N_1438,N_960,In_79);
xor U1439 (N_1439,In_1020,N_503);
xnor U1440 (N_1440,N_764,N_890);
and U1441 (N_1441,N_876,N_618);
and U1442 (N_1442,N_414,In_1164);
and U1443 (N_1443,N_162,In_0);
or U1444 (N_1444,In_2113,N_956);
and U1445 (N_1445,In_693,N_535);
nor U1446 (N_1446,N_569,In_979);
xnor U1447 (N_1447,N_763,In_2092);
and U1448 (N_1448,In_624,In_2474);
or U1449 (N_1449,N_516,N_990);
xor U1450 (N_1450,N_541,In_1340);
nand U1451 (N_1451,N_264,In_634);
and U1452 (N_1452,In_757,N_467);
nor U1453 (N_1453,N_637,In_2439);
or U1454 (N_1454,N_873,N_78);
nor U1455 (N_1455,In_2378,In_1392);
xnor U1456 (N_1456,N_735,N_676);
nor U1457 (N_1457,N_812,In_775);
xor U1458 (N_1458,N_824,N_680);
or U1459 (N_1459,In_1551,In_1227);
xnor U1460 (N_1460,N_370,In_1468);
xnor U1461 (N_1461,N_301,In_2061);
or U1462 (N_1462,N_427,N_985);
nand U1463 (N_1463,N_681,N_235);
nand U1464 (N_1464,In_1471,In_1424);
and U1465 (N_1465,In_785,N_670);
and U1466 (N_1466,In_1918,N_320);
xnor U1467 (N_1467,In_1349,N_278);
nor U1468 (N_1468,N_424,N_980);
nand U1469 (N_1469,In_1180,In_2128);
xnor U1470 (N_1470,N_664,In_478);
or U1471 (N_1471,In_2475,N_241);
nor U1472 (N_1472,N_949,N_891);
nand U1473 (N_1473,N_608,N_218);
xnor U1474 (N_1474,N_834,N_597);
nand U1475 (N_1475,N_708,N_417);
or U1476 (N_1476,In_1288,N_485);
nand U1477 (N_1477,N_448,N_691);
or U1478 (N_1478,In_953,N_888);
nor U1479 (N_1479,In_968,In_1343);
xor U1480 (N_1480,In_2117,N_480);
or U1481 (N_1481,In_175,N_767);
and U1482 (N_1482,In_1677,In_2292);
nor U1483 (N_1483,N_45,N_477);
nor U1484 (N_1484,In_291,N_590);
or U1485 (N_1485,N_882,N_895);
and U1486 (N_1486,N_920,In_1648);
or U1487 (N_1487,In_692,N_928);
or U1488 (N_1488,In_1132,N_472);
nand U1489 (N_1489,N_903,N_830);
nand U1490 (N_1490,N_602,In_2217);
or U1491 (N_1491,N_61,In_1010);
nand U1492 (N_1492,In_1166,N_217);
nand U1493 (N_1493,N_612,N_829);
nor U1494 (N_1494,N_69,In_50);
or U1495 (N_1495,In_1576,N_822);
xnor U1496 (N_1496,N_87,N_306);
nand U1497 (N_1497,N_821,N_860);
nor U1498 (N_1498,N_546,N_855);
or U1499 (N_1499,In_22,N_725);
or U1500 (N_1500,N_84,N_25);
and U1501 (N_1501,N_959,N_328);
xor U1502 (N_1502,N_991,N_645);
nand U1503 (N_1503,N_545,In_863);
nand U1504 (N_1504,N_902,N_204);
nor U1505 (N_1505,N_295,N_804);
nand U1506 (N_1506,N_558,N_878);
xor U1507 (N_1507,In_503,In_1615);
and U1508 (N_1508,N_994,N_654);
nor U1509 (N_1509,In_244,N_141);
or U1510 (N_1510,N_226,In_1633);
or U1511 (N_1511,N_666,N_413);
xnor U1512 (N_1512,In_259,N_305);
xnor U1513 (N_1513,N_156,N_983);
nand U1514 (N_1514,N_473,N_403);
or U1515 (N_1515,In_1220,N_259);
nor U1516 (N_1516,N_299,N_323);
or U1517 (N_1517,N_345,N_731);
nand U1518 (N_1518,N_179,N_409);
nor U1519 (N_1519,N_98,N_395);
nand U1520 (N_1520,N_719,N_67);
nor U1521 (N_1521,N_712,N_468);
nand U1522 (N_1522,N_209,N_582);
or U1523 (N_1523,In_1622,In_1940);
and U1524 (N_1524,N_17,In_789);
xnor U1525 (N_1525,N_132,In_844);
nor U1526 (N_1526,N_384,In_2094);
and U1527 (N_1527,In_1742,N_592);
or U1528 (N_1528,In_1594,N_840);
or U1529 (N_1529,N_475,In_322);
nor U1530 (N_1530,N_518,In_1131);
nand U1531 (N_1531,N_85,In_460);
and U1532 (N_1532,N_24,N_128);
and U1533 (N_1533,N_127,N_885);
nor U1534 (N_1534,N_867,N_461);
nand U1535 (N_1535,In_81,N_892);
xor U1536 (N_1536,In_2029,N_130);
nor U1537 (N_1537,In_1893,N_385);
or U1538 (N_1538,N_872,N_536);
and U1539 (N_1539,In_226,In_2293);
xnor U1540 (N_1540,N_810,N_133);
xor U1541 (N_1541,N_520,N_706);
or U1542 (N_1542,In_521,In_51);
nor U1543 (N_1543,N_273,N_609);
and U1544 (N_1544,N_640,In_2408);
nor U1545 (N_1545,N_678,In_308);
nand U1546 (N_1546,In_2453,N_62);
and U1547 (N_1547,N_993,In_902);
xor U1548 (N_1548,N_986,N_166);
xor U1549 (N_1549,In_2149,N_927);
nor U1550 (N_1550,N_714,In_349);
nor U1551 (N_1551,In_1601,N_469);
nand U1552 (N_1552,In_1829,N_744);
nor U1553 (N_1553,In_2089,N_679);
or U1554 (N_1554,N_476,N_551);
xor U1555 (N_1555,In_713,In_701);
nand U1556 (N_1556,In_1793,N_265);
and U1557 (N_1557,N_754,N_527);
xnor U1558 (N_1558,N_998,In_1901);
and U1559 (N_1559,N_412,N_757);
nand U1560 (N_1560,In_1263,N_270);
or U1561 (N_1561,N_374,N_636);
or U1562 (N_1562,In_2121,In_93);
nand U1563 (N_1563,N_506,N_254);
nand U1564 (N_1564,N_642,N_438);
nor U1565 (N_1565,N_244,In_1219);
nand U1566 (N_1566,N_159,In_2401);
and U1567 (N_1567,N_528,N_139);
or U1568 (N_1568,N_239,In_1982);
nand U1569 (N_1569,N_203,In_1097);
xnor U1570 (N_1570,N_721,N_55);
and U1571 (N_1571,N_454,N_108);
nand U1572 (N_1572,In_401,N_695);
nand U1573 (N_1573,In_527,N_717);
and U1574 (N_1574,N_31,In_1629);
nor U1575 (N_1575,N_667,In_2069);
or U1576 (N_1576,In_2376,In_2458);
or U1577 (N_1577,In_2335,N_865);
and U1578 (N_1578,N_623,N_954);
xor U1579 (N_1579,In_214,N_351);
or U1580 (N_1580,N_500,N_115);
or U1581 (N_1581,In_377,N_148);
and U1582 (N_1582,N_556,In_612);
and U1583 (N_1583,N_931,N_797);
or U1584 (N_1584,N_776,N_765);
or U1585 (N_1585,N_71,In_2135);
nand U1586 (N_1586,N_242,N_175);
nor U1587 (N_1587,N_965,N_92);
nor U1588 (N_1588,N_709,N_952);
and U1589 (N_1589,In_1830,N_387);
nor U1590 (N_1590,In_1058,In_1839);
or U1591 (N_1591,In_1684,In_135);
and U1592 (N_1592,N_422,In_2284);
or U1593 (N_1593,N_942,N_529);
nand U1594 (N_1594,N_796,N_561);
nor U1595 (N_1595,N_701,In_344);
xnor U1596 (N_1596,N_489,N_819);
and U1597 (N_1597,N_847,N_910);
or U1598 (N_1598,In_848,N_111);
xnor U1599 (N_1599,In_772,N_193);
nand U1600 (N_1600,N_749,N_220);
xor U1601 (N_1601,In_1653,In_1038);
nand U1602 (N_1602,In_2074,N_950);
and U1603 (N_1603,N_464,N_992);
or U1604 (N_1604,In_1641,N_933);
or U1605 (N_1605,N_534,N_710);
nor U1606 (N_1606,In_2068,N_302);
or U1607 (N_1607,N_300,N_793);
xnor U1608 (N_1608,N_309,N_347);
nand U1609 (N_1609,In_744,N_583);
and U1610 (N_1610,N_683,N_367);
nor U1611 (N_1611,N_163,N_766);
or U1612 (N_1612,In_1657,N_74);
or U1613 (N_1613,N_206,In_1702);
nand U1614 (N_1614,N_620,N_23);
xor U1615 (N_1615,In_480,N_337);
nand U1616 (N_1616,N_853,In_2387);
or U1617 (N_1617,N_478,N_512);
nor U1618 (N_1618,N_261,In_2014);
nor U1619 (N_1619,N_734,In_1628);
xor U1620 (N_1620,In_1283,In_663);
nand U1621 (N_1621,In_2402,N_607);
xnor U1622 (N_1622,N_230,N_720);
xnor U1623 (N_1623,N_430,In_99);
and U1624 (N_1624,N_736,In_463);
or U1625 (N_1625,In_1678,N_898);
nand U1626 (N_1626,N_864,N_40);
nand U1627 (N_1627,In_2302,In_194);
and U1628 (N_1628,N_211,In_917);
nand U1629 (N_1629,N_22,In_420);
xnor U1630 (N_1630,N_18,N_718);
and U1631 (N_1631,N_279,In_581);
nand U1632 (N_1632,In_749,In_1855);
nor U1633 (N_1633,In_747,N_606);
or U1634 (N_1634,In_443,N_338);
nor U1635 (N_1635,In_2045,N_191);
nor U1636 (N_1636,In_1086,N_580);
xor U1637 (N_1637,N_303,N_700);
xor U1638 (N_1638,N_507,In_1837);
nand U1639 (N_1639,In_2044,N_653);
or U1640 (N_1640,N_52,N_594);
and U1641 (N_1641,In_1718,N_838);
xor U1642 (N_1642,In_921,N_63);
xor U1643 (N_1643,N_196,In_2016);
nor U1644 (N_1644,N_641,N_57);
nor U1645 (N_1645,N_194,In_2294);
nand U1646 (N_1646,N_786,N_167);
and U1647 (N_1647,N_463,N_449);
xor U1648 (N_1648,N_968,In_1466);
nand U1649 (N_1649,N_768,N_739);
nand U1650 (N_1650,In_88,In_418);
or U1651 (N_1651,In_2220,N_946);
or U1652 (N_1652,N_282,In_1578);
xnor U1653 (N_1653,In_852,N_82);
or U1654 (N_1654,N_453,N_465);
and U1655 (N_1655,N_548,N_406);
nand U1656 (N_1656,N_682,N_496);
and U1657 (N_1657,N_43,N_851);
xnor U1658 (N_1658,N_0,In_312);
and U1659 (N_1659,N_800,N_379);
and U1660 (N_1660,N_852,N_213);
and U1661 (N_1661,N_962,In_1704);
nand U1662 (N_1662,N_747,N_901);
nand U1663 (N_1663,N_1,N_772);
xnor U1664 (N_1664,In_2283,In_2267);
nand U1665 (N_1665,In_1439,In_2035);
or U1666 (N_1666,In_1804,In_2254);
or U1667 (N_1667,N_93,N_857);
or U1668 (N_1668,N_180,N_310);
or U1669 (N_1669,N_837,N_803);
nor U1670 (N_1670,In_1571,N_77);
nor U1671 (N_1671,N_90,N_554);
or U1672 (N_1672,N_783,N_687);
nor U1673 (N_1673,In_1033,In_1119);
or U1674 (N_1674,N_342,N_431);
xor U1675 (N_1675,N_117,In_1022);
or U1676 (N_1676,In_2084,In_160);
nor U1677 (N_1677,N_557,In_680);
xor U1678 (N_1678,N_291,N_843);
nor U1679 (N_1679,N_249,N_240);
xnor U1680 (N_1680,In_342,In_2208);
nor U1681 (N_1681,N_658,In_2266);
nand U1682 (N_1682,In_1478,In_1449);
xor U1683 (N_1683,N_268,N_742);
xnor U1684 (N_1684,N_5,N_312);
nor U1685 (N_1685,In_719,N_748);
or U1686 (N_1686,In_768,In_1351);
nor U1687 (N_1687,N_462,In_1797);
xor U1688 (N_1688,N_221,N_76);
or U1689 (N_1689,In_86,In_964);
nor U1690 (N_1690,N_533,N_304);
xnor U1691 (N_1691,N_176,In_2256);
nor U1692 (N_1692,N_188,N_113);
nand U1693 (N_1693,In_151,In_769);
nor U1694 (N_1694,N_75,In_601);
nor U1695 (N_1695,N_684,N_164);
or U1696 (N_1696,In_2146,N_732);
nor U1697 (N_1697,In_1405,N_245);
and U1698 (N_1698,N_219,N_364);
nor U1699 (N_1699,In_1133,N_389);
xor U1700 (N_1700,N_174,N_470);
nand U1701 (N_1701,In_1698,N_258);
or U1702 (N_1702,In_472,N_813);
xor U1703 (N_1703,N_271,N_32);
or U1704 (N_1704,N_64,N_499);
or U1705 (N_1705,N_831,N_137);
nand U1706 (N_1706,N_625,N_859);
xor U1707 (N_1707,In_823,N_208);
nor U1708 (N_1708,N_398,N_643);
nand U1709 (N_1709,N_572,In_330);
nand U1710 (N_1710,In_2492,In_2232);
xnor U1711 (N_1711,In_1496,N_581);
xor U1712 (N_1712,In_7,N_214);
or U1713 (N_1713,N_854,N_14);
and U1714 (N_1714,N_756,N_118);
or U1715 (N_1715,N_7,N_650);
nor U1716 (N_1716,N_50,N_907);
nand U1717 (N_1717,N_112,N_945);
or U1718 (N_1718,N_59,N_177);
and U1719 (N_1719,In_561,N_297);
and U1720 (N_1720,In_939,N_560);
or U1721 (N_1721,N_866,In_2180);
and U1722 (N_1722,In_2004,In_1574);
and U1723 (N_1723,In_298,N_311);
or U1724 (N_1724,N_135,N_794);
or U1725 (N_1725,N_42,N_354);
xor U1726 (N_1726,In_1884,N_105);
nand U1727 (N_1727,In_629,N_490);
nand U1728 (N_1728,In_2052,N_573);
and U1729 (N_1729,N_172,N_479);
nand U1730 (N_1730,N_999,In_1996);
and U1731 (N_1731,N_549,In_1152);
or U1732 (N_1732,N_501,In_974);
nor U1733 (N_1733,In_1841,N_805);
xnor U1734 (N_1734,In_2059,N_914);
or U1735 (N_1735,In_1005,N_585);
xnor U1736 (N_1736,N_198,In_231);
nor U1737 (N_1737,In_1027,N_697);
xor U1738 (N_1738,N_269,N_341);
nand U1739 (N_1739,In_354,N_743);
nand U1740 (N_1740,In_883,N_416);
xor U1741 (N_1741,N_124,N_604);
and U1742 (N_1742,N_28,N_155);
nor U1743 (N_1743,In_216,N_321);
nor U1744 (N_1744,N_598,N_358);
and U1745 (N_1745,N_578,N_89);
or U1746 (N_1746,N_646,N_924);
or U1747 (N_1747,N_790,N_382);
xnor U1748 (N_1748,In_1509,N_532);
nor U1749 (N_1749,N_823,N_421);
and U1750 (N_1750,In_1858,In_953);
and U1751 (N_1751,In_614,N_184);
nor U1752 (N_1752,N_518,In_701);
nor U1753 (N_1753,In_374,In_475);
nand U1754 (N_1754,N_489,N_372);
xor U1755 (N_1755,N_952,In_341);
nand U1756 (N_1756,N_707,N_909);
and U1757 (N_1757,N_660,In_216);
nor U1758 (N_1758,N_114,In_1005);
and U1759 (N_1759,In_1297,N_675);
xnor U1760 (N_1760,In_1220,N_117);
nand U1761 (N_1761,N_845,In_1016);
xor U1762 (N_1762,N_524,N_255);
nor U1763 (N_1763,N_920,In_2456);
nand U1764 (N_1764,N_544,N_847);
nor U1765 (N_1765,N_912,N_759);
xor U1766 (N_1766,In_115,N_972);
xor U1767 (N_1767,In_702,N_128);
xor U1768 (N_1768,In_164,N_613);
nand U1769 (N_1769,N_677,In_2456);
xor U1770 (N_1770,N_161,N_127);
nand U1771 (N_1771,N_789,N_376);
nor U1772 (N_1772,N_780,In_712);
xnor U1773 (N_1773,N_801,In_2014);
xor U1774 (N_1774,In_422,N_771);
nand U1775 (N_1775,N_982,N_831);
xnor U1776 (N_1776,N_419,N_520);
nor U1777 (N_1777,N_210,N_39);
and U1778 (N_1778,N_36,N_449);
nand U1779 (N_1779,N_12,N_36);
xnor U1780 (N_1780,N_787,In_164);
nor U1781 (N_1781,N_768,N_408);
or U1782 (N_1782,In_989,In_194);
nor U1783 (N_1783,In_50,In_1283);
xor U1784 (N_1784,In_2082,N_262);
nor U1785 (N_1785,N_879,N_126);
nand U1786 (N_1786,N_746,N_902);
nor U1787 (N_1787,In_478,N_487);
xor U1788 (N_1788,N_728,In_593);
xor U1789 (N_1789,N_589,N_537);
and U1790 (N_1790,N_115,N_455);
nand U1791 (N_1791,N_69,N_758);
nor U1792 (N_1792,In_823,In_634);
xor U1793 (N_1793,N_6,N_473);
nand U1794 (N_1794,N_937,In_316);
and U1795 (N_1795,N_388,In_863);
and U1796 (N_1796,N_351,In_189);
or U1797 (N_1797,In_898,N_547);
xnor U1798 (N_1798,N_268,N_15);
nand U1799 (N_1799,N_964,N_676);
xnor U1800 (N_1800,N_603,In_1843);
or U1801 (N_1801,N_415,N_560);
and U1802 (N_1802,N_984,N_176);
xor U1803 (N_1803,N_943,In_1551);
or U1804 (N_1804,In_2239,In_950);
nand U1805 (N_1805,N_866,In_841);
or U1806 (N_1806,N_77,N_775);
and U1807 (N_1807,N_881,In_2);
and U1808 (N_1808,N_997,In_2092);
nor U1809 (N_1809,N_934,In_2367);
nand U1810 (N_1810,In_1276,N_311);
nor U1811 (N_1811,In_791,N_10);
and U1812 (N_1812,N_151,N_328);
nor U1813 (N_1813,N_78,In_50);
nand U1814 (N_1814,N_829,N_24);
xor U1815 (N_1815,N_765,In_2388);
and U1816 (N_1816,N_548,N_579);
and U1817 (N_1817,N_80,N_155);
nor U1818 (N_1818,N_834,In_1212);
and U1819 (N_1819,N_509,N_672);
xor U1820 (N_1820,In_2107,In_2073);
and U1821 (N_1821,N_826,N_11);
nand U1822 (N_1822,N_633,N_778);
nand U1823 (N_1823,N_263,In_1275);
or U1824 (N_1824,N_971,In_1122);
nand U1825 (N_1825,In_2208,N_351);
nand U1826 (N_1826,N_498,In_607);
or U1827 (N_1827,N_398,N_249);
xnor U1828 (N_1828,In_1751,N_162);
or U1829 (N_1829,N_763,N_479);
nand U1830 (N_1830,N_220,In_106);
xnor U1831 (N_1831,In_536,In_1020);
or U1832 (N_1832,In_330,N_159);
nand U1833 (N_1833,N_833,N_678);
xnor U1834 (N_1834,N_545,N_501);
or U1835 (N_1835,N_838,N_867);
nor U1836 (N_1836,In_455,N_46);
and U1837 (N_1837,In_2367,N_892);
and U1838 (N_1838,N_878,In_238);
xnor U1839 (N_1839,N_930,N_824);
nand U1840 (N_1840,In_758,N_479);
xor U1841 (N_1841,N_180,N_620);
xor U1842 (N_1842,N_713,In_178);
nand U1843 (N_1843,In_2444,N_730);
xor U1844 (N_1844,N_970,N_936);
and U1845 (N_1845,N_978,N_267);
nor U1846 (N_1846,In_1901,N_930);
or U1847 (N_1847,In_231,In_149);
nor U1848 (N_1848,N_165,N_285);
and U1849 (N_1849,N_765,N_668);
or U1850 (N_1850,N_120,N_571);
nand U1851 (N_1851,N_49,N_878);
nand U1852 (N_1852,N_563,N_438);
xor U1853 (N_1853,N_784,In_272);
xor U1854 (N_1854,In_731,N_402);
nor U1855 (N_1855,N_425,In_519);
xor U1856 (N_1856,N_171,N_511);
or U1857 (N_1857,N_212,In_692);
xor U1858 (N_1858,N_215,N_715);
nor U1859 (N_1859,In_472,N_120);
nor U1860 (N_1860,In_1124,N_499);
and U1861 (N_1861,N_271,N_377);
xor U1862 (N_1862,N_449,In_377);
and U1863 (N_1863,In_2035,In_2456);
xnor U1864 (N_1864,In_1567,N_916);
or U1865 (N_1865,N_328,N_564);
or U1866 (N_1866,In_553,N_101);
xnor U1867 (N_1867,In_294,In_115);
nand U1868 (N_1868,N_82,N_869);
and U1869 (N_1869,N_810,N_407);
nor U1870 (N_1870,In_524,N_35);
xnor U1871 (N_1871,N_736,In_1077);
and U1872 (N_1872,In_1816,N_24);
or U1873 (N_1873,In_524,N_449);
and U1874 (N_1874,In_782,N_639);
xnor U1875 (N_1875,N_19,In_1751);
nor U1876 (N_1876,In_2121,In_480);
and U1877 (N_1877,In_354,N_145);
xnor U1878 (N_1878,N_986,N_739);
xnor U1879 (N_1879,N_306,N_508);
xnor U1880 (N_1880,N_757,In_1496);
nor U1881 (N_1881,In_2146,N_135);
or U1882 (N_1882,N_866,In_614);
or U1883 (N_1883,N_46,N_211);
or U1884 (N_1884,N_95,N_965);
nor U1885 (N_1885,In_880,N_896);
and U1886 (N_1886,N_693,In_1468);
xnor U1887 (N_1887,In_1008,N_636);
nor U1888 (N_1888,In_602,N_385);
xor U1889 (N_1889,In_1244,N_655);
or U1890 (N_1890,N_809,In_1935);
nor U1891 (N_1891,N_636,In_1124);
or U1892 (N_1892,N_393,N_272);
and U1893 (N_1893,In_1311,N_116);
or U1894 (N_1894,N_869,N_855);
and U1895 (N_1895,N_275,N_320);
nand U1896 (N_1896,N_719,N_124);
or U1897 (N_1897,In_342,In_22);
and U1898 (N_1898,N_560,N_737);
and U1899 (N_1899,N_495,In_702);
nand U1900 (N_1900,In_1033,In_1022);
nor U1901 (N_1901,N_288,N_149);
and U1902 (N_1902,N_528,In_1705);
nand U1903 (N_1903,In_1674,N_800);
xnor U1904 (N_1904,N_714,In_181);
nor U1905 (N_1905,N_75,N_893);
nor U1906 (N_1906,In_2328,In_2069);
and U1907 (N_1907,N_380,N_953);
or U1908 (N_1908,N_815,N_466);
xnor U1909 (N_1909,N_963,N_859);
nor U1910 (N_1910,N_500,In_2146);
nand U1911 (N_1911,N_627,In_2256);
or U1912 (N_1912,N_198,N_208);
xnor U1913 (N_1913,N_418,N_257);
and U1914 (N_1914,N_330,In_1086);
nand U1915 (N_1915,N_88,N_692);
xor U1916 (N_1916,In_1347,In_1793);
nand U1917 (N_1917,N_832,N_686);
or U1918 (N_1918,In_2196,In_2317);
nand U1919 (N_1919,N_469,N_700);
xnor U1920 (N_1920,N_674,N_249);
or U1921 (N_1921,In_2251,In_1008);
nand U1922 (N_1922,In_88,N_70);
nand U1923 (N_1923,N_833,N_144);
nand U1924 (N_1924,In_2232,N_628);
and U1925 (N_1925,N_879,In_389);
and U1926 (N_1926,N_404,N_61);
or U1927 (N_1927,In_965,N_357);
nor U1928 (N_1928,N_838,N_130);
or U1929 (N_1929,N_275,In_2149);
nor U1930 (N_1930,N_58,In_2246);
nand U1931 (N_1931,N_546,N_49);
nand U1932 (N_1932,In_2068,N_821);
and U1933 (N_1933,N_590,N_592);
nor U1934 (N_1934,N_686,In_2122);
xnor U1935 (N_1935,N_405,In_1340);
nand U1936 (N_1936,N_923,N_550);
nor U1937 (N_1937,N_363,N_341);
or U1938 (N_1938,N_132,N_130);
xnor U1939 (N_1939,N_79,N_324);
xor U1940 (N_1940,In_1131,N_359);
nor U1941 (N_1941,In_194,In_320);
nand U1942 (N_1942,In_744,N_753);
and U1943 (N_1943,N_435,N_587);
nor U1944 (N_1944,In_2106,N_741);
and U1945 (N_1945,N_390,In_2492);
xnor U1946 (N_1946,N_168,N_609);
xnor U1947 (N_1947,In_2346,N_919);
or U1948 (N_1948,N_170,N_37);
nor U1949 (N_1949,In_1349,In_2110);
xnor U1950 (N_1950,N_527,N_731);
nor U1951 (N_1951,N_469,N_956);
or U1952 (N_1952,In_2388,N_733);
xor U1953 (N_1953,N_885,N_505);
and U1954 (N_1954,N_559,N_603);
nand U1955 (N_1955,N_53,In_2052);
or U1956 (N_1956,N_835,N_196);
nor U1957 (N_1957,In_917,N_740);
nor U1958 (N_1958,In_593,N_128);
xor U1959 (N_1959,N_632,In_2068);
and U1960 (N_1960,In_917,In_1731);
nand U1961 (N_1961,N_785,N_937);
nor U1962 (N_1962,N_489,In_2316);
or U1963 (N_1963,N_109,N_657);
and U1964 (N_1964,In_1858,N_218);
nand U1965 (N_1965,N_141,N_874);
or U1966 (N_1966,N_648,N_463);
nor U1967 (N_1967,N_127,N_449);
nor U1968 (N_1968,In_2284,N_525);
xnor U1969 (N_1969,In_50,In_2476);
or U1970 (N_1970,N_48,N_561);
nor U1971 (N_1971,In_2401,In_1745);
nor U1972 (N_1972,N_429,In_1020);
nand U1973 (N_1973,N_377,In_312);
xor U1974 (N_1974,N_718,In_1677);
xnor U1975 (N_1975,N_714,In_2478);
or U1976 (N_1976,N_310,N_803);
nor U1977 (N_1977,N_293,In_602);
or U1978 (N_1978,N_911,N_748);
or U1979 (N_1979,In_463,N_862);
nor U1980 (N_1980,In_1324,N_520);
or U1981 (N_1981,In_1180,N_220);
and U1982 (N_1982,In_983,N_468);
nand U1983 (N_1983,N_229,N_819);
nor U1984 (N_1984,N_576,N_250);
or U1985 (N_1985,N_645,In_519);
nand U1986 (N_1986,N_363,N_506);
xor U1987 (N_1987,N_338,N_205);
nand U1988 (N_1988,N_198,N_217);
or U1989 (N_1989,N_809,In_2350);
and U1990 (N_1990,N_414,In_7);
nor U1991 (N_1991,N_732,N_915);
nand U1992 (N_1992,N_551,N_881);
nand U1993 (N_1993,N_104,N_585);
or U1994 (N_1994,N_772,N_71);
and U1995 (N_1995,N_51,N_837);
or U1996 (N_1996,In_617,N_342);
nand U1997 (N_1997,N_455,N_890);
and U1998 (N_1998,N_740,N_291);
nor U1999 (N_1999,N_603,N_827);
xnor U2000 (N_2000,N_1789,N_1955);
xor U2001 (N_2001,N_1101,N_1905);
nor U2002 (N_2002,N_1743,N_1493);
xor U2003 (N_2003,N_1710,N_1153);
xor U2004 (N_2004,N_1884,N_1533);
nand U2005 (N_2005,N_1257,N_1082);
or U2006 (N_2006,N_1013,N_1632);
or U2007 (N_2007,N_1201,N_1412);
nor U2008 (N_2008,N_1898,N_1599);
and U2009 (N_2009,N_1538,N_1634);
xnor U2010 (N_2010,N_1732,N_1236);
or U2011 (N_2011,N_1446,N_1171);
nand U2012 (N_2012,N_1232,N_1733);
nand U2013 (N_2013,N_1140,N_1172);
or U2014 (N_2014,N_1114,N_1092);
or U2015 (N_2015,N_1550,N_1763);
nand U2016 (N_2016,N_1456,N_1361);
xor U2017 (N_2017,N_1668,N_1139);
or U2018 (N_2018,N_1860,N_1633);
and U2019 (N_2019,N_1751,N_1509);
nand U2020 (N_2020,N_1779,N_1258);
nand U2021 (N_2021,N_1458,N_1304);
or U2022 (N_2022,N_1765,N_1679);
xnor U2023 (N_2023,N_1397,N_1906);
nor U2024 (N_2024,N_1133,N_1930);
and U2025 (N_2025,N_1831,N_1503);
or U2026 (N_2026,N_1323,N_1600);
xnor U2027 (N_2027,N_1769,N_1312);
xor U2028 (N_2028,N_1627,N_1369);
nand U2029 (N_2029,N_1506,N_1249);
or U2030 (N_2030,N_1995,N_1598);
and U2031 (N_2031,N_1650,N_1565);
nor U2032 (N_2032,N_1074,N_1242);
nor U2033 (N_2033,N_1180,N_1534);
nand U2034 (N_2034,N_1519,N_1891);
nand U2035 (N_2035,N_1672,N_1773);
xnor U2036 (N_2036,N_1522,N_1963);
xnor U2037 (N_2037,N_1088,N_1603);
nand U2038 (N_2038,N_1994,N_1929);
xnor U2039 (N_2039,N_1742,N_1871);
or U2040 (N_2040,N_1774,N_1136);
nand U2041 (N_2041,N_1402,N_1681);
nor U2042 (N_2042,N_1965,N_1524);
and U2043 (N_2043,N_1319,N_1273);
and U2044 (N_2044,N_1337,N_1355);
nor U2045 (N_2045,N_1901,N_1941);
and U2046 (N_2046,N_1561,N_1727);
nor U2047 (N_2047,N_1064,N_1240);
xnor U2048 (N_2048,N_1564,N_1025);
nand U2049 (N_2049,N_1676,N_1974);
or U2050 (N_2050,N_1328,N_1935);
nand U2051 (N_2051,N_1462,N_1999);
xor U2052 (N_2052,N_1569,N_1712);
nor U2053 (N_2053,N_1947,N_1996);
nor U2054 (N_2054,N_1078,N_1543);
nor U2055 (N_2055,N_1287,N_1507);
nand U2056 (N_2056,N_1844,N_1539);
nand U2057 (N_2057,N_1017,N_1185);
nand U2058 (N_2058,N_1387,N_1448);
or U2059 (N_2059,N_1515,N_1854);
and U2060 (N_2060,N_1837,N_1120);
and U2061 (N_2061,N_1667,N_1626);
or U2062 (N_2062,N_1188,N_1170);
xor U2063 (N_2063,N_1948,N_1642);
or U2064 (N_2064,N_1640,N_1371);
nand U2065 (N_2065,N_1094,N_1919);
nand U2066 (N_2066,N_1793,N_1848);
or U2067 (N_2067,N_1159,N_1804);
nand U2068 (N_2068,N_1005,N_1708);
xor U2069 (N_2069,N_1581,N_1211);
and U2070 (N_2070,N_1570,N_1969);
xnor U2071 (N_2071,N_1272,N_1436);
and U2072 (N_2072,N_1080,N_1453);
nand U2073 (N_2073,N_1334,N_1066);
or U2074 (N_2074,N_1520,N_1112);
nand U2075 (N_2075,N_1567,N_1239);
or U2076 (N_2076,N_1745,N_1487);
nor U2077 (N_2077,N_1807,N_1032);
nand U2078 (N_2078,N_1942,N_1729);
or U2079 (N_2079,N_1872,N_1091);
and U2080 (N_2080,N_1279,N_1571);
or U2081 (N_2081,N_1812,N_1580);
and U2082 (N_2082,N_1778,N_1476);
or U2083 (N_2083,N_1692,N_1870);
nor U2084 (N_2084,N_1485,N_1018);
nand U2085 (N_2085,N_1490,N_1873);
nand U2086 (N_2086,N_1644,N_1894);
nand U2087 (N_2087,N_1877,N_1531);
nand U2088 (N_2088,N_1728,N_1434);
or U2089 (N_2089,N_1132,N_1103);
nor U2090 (N_2090,N_1788,N_1726);
and U2091 (N_2091,N_1663,N_1081);
or U2092 (N_2092,N_1852,N_1408);
xnor U2093 (N_2093,N_1757,N_1076);
or U2094 (N_2094,N_1843,N_1268);
and U2095 (N_2095,N_1488,N_1959);
and U2096 (N_2096,N_1164,N_1404);
xor U2097 (N_2097,N_1145,N_1719);
and U2098 (N_2098,N_1554,N_1255);
or U2099 (N_2099,N_1622,N_1968);
and U2100 (N_2100,N_1160,N_1563);
xor U2101 (N_2101,N_1973,N_1178);
and U2102 (N_2102,N_1219,N_1698);
nand U2103 (N_2103,N_1875,N_1828);
xor U2104 (N_2104,N_1428,N_1970);
or U2105 (N_2105,N_1115,N_1611);
or U2106 (N_2106,N_1311,N_1984);
xor U2107 (N_2107,N_1466,N_1098);
or U2108 (N_2108,N_1233,N_1855);
or U2109 (N_2109,N_1956,N_1053);
xor U2110 (N_2110,N_1912,N_1004);
or U2111 (N_2111,N_1228,N_1464);
xnor U2112 (N_2112,N_1197,N_1297);
xnor U2113 (N_2113,N_1442,N_1760);
nor U2114 (N_2114,N_1666,N_1479);
nor U2115 (N_2115,N_1780,N_1356);
nand U2116 (N_2116,N_1386,N_1606);
nand U2117 (N_2117,N_1093,N_1484);
and U2118 (N_2118,N_1203,N_1340);
and U2119 (N_2119,N_1890,N_1546);
and U2120 (N_2120,N_1035,N_1011);
or U2121 (N_2121,N_1042,N_1331);
xor U2122 (N_2122,N_1108,N_1235);
xnor U2123 (N_2123,N_1787,N_1986);
nor U2124 (N_2124,N_1753,N_1510);
or U2125 (N_2125,N_1010,N_1186);
nor U2126 (N_2126,N_1913,N_1151);
or U2127 (N_2127,N_1310,N_1975);
xor U2128 (N_2128,N_1750,N_1688);
or U2129 (N_2129,N_1009,N_1578);
nand U2130 (N_2130,N_1477,N_1799);
nor U2131 (N_2131,N_1189,N_1734);
or U2132 (N_2132,N_1585,N_1348);
or U2133 (N_2133,N_1041,N_1922);
nand U2134 (N_2134,N_1266,N_1682);
or U2135 (N_2135,N_1089,N_1154);
and U2136 (N_2136,N_1864,N_1661);
or U2137 (N_2137,N_1654,N_1730);
nand U2138 (N_2138,N_1097,N_1953);
and U2139 (N_2139,N_1724,N_1686);
nor U2140 (N_2140,N_1020,N_1961);
nor U2141 (N_2141,N_1016,N_1949);
xor U2142 (N_2142,N_1617,N_1128);
xnor U2143 (N_2143,N_1339,N_1983);
xnor U2144 (N_2144,N_1892,N_1471);
xor U2145 (N_2145,N_1111,N_1928);
nor U2146 (N_2146,N_1336,N_1940);
nor U2147 (N_2147,N_1687,N_1615);
or U2148 (N_2148,N_1165,N_1338);
and U2149 (N_2149,N_1146,N_1923);
or U2150 (N_2150,N_1879,N_1902);
or U2151 (N_2151,N_1019,N_1579);
xnor U2152 (N_2152,N_1060,N_1288);
nor U2153 (N_2153,N_1226,N_1300);
nor U2154 (N_2154,N_1521,N_1029);
nor U2155 (N_2155,N_1208,N_1869);
nand U2156 (N_2156,N_1370,N_1435);
and U2157 (N_2157,N_1440,N_1196);
nand U2158 (N_2158,N_1985,N_1784);
and U2159 (N_2159,N_1205,N_1911);
and U2160 (N_2160,N_1150,N_1424);
or U2161 (N_2161,N_1480,N_1405);
nand U2162 (N_2162,N_1980,N_1823);
xor U2163 (N_2163,N_1438,N_1392);
and U2164 (N_2164,N_1003,N_1847);
nor U2165 (N_2165,N_1280,N_1702);
or U2166 (N_2166,N_1414,N_1293);
or U2167 (N_2167,N_1330,N_1275);
and U2168 (N_2168,N_1467,N_1641);
nor U2169 (N_2169,N_1212,N_1437);
and U2170 (N_2170,N_1758,N_1937);
nand U2171 (N_2171,N_1991,N_1631);
nor U2172 (N_2172,N_1298,N_1158);
xor U2173 (N_2173,N_1122,N_1006);
nor U2174 (N_2174,N_1499,N_1938);
or U2175 (N_2175,N_1214,N_1075);
xnor U2176 (N_2176,N_1368,N_1327);
nor U2177 (N_2177,N_1262,N_1452);
xnor U2178 (N_2178,N_1142,N_1978);
or U2179 (N_2179,N_1829,N_1358);
nand U2180 (N_2180,N_1116,N_1764);
or U2181 (N_2181,N_1086,N_1678);
nor U2182 (N_2182,N_1785,N_1625);
or U2183 (N_2183,N_1447,N_1776);
and U2184 (N_2184,N_1084,N_1241);
nand U2185 (N_2185,N_1685,N_1762);
or U2186 (N_2186,N_1977,N_1988);
or U2187 (N_2187,N_1796,N_1391);
or U2188 (N_2188,N_1748,N_1992);
nor U2189 (N_2189,N_1276,N_1529);
xor U2190 (N_2190,N_1144,N_1118);
and U2191 (N_2191,N_1989,N_1468);
xor U2192 (N_2192,N_1317,N_1586);
nor U2193 (N_2193,N_1706,N_1691);
or U2194 (N_2194,N_1417,N_1709);
or U2195 (N_2195,N_1878,N_1549);
xnor U2196 (N_2196,N_1489,N_1156);
or U2197 (N_2197,N_1047,N_1362);
and U2198 (N_2198,N_1166,N_1562);
nor U2199 (N_2199,N_1411,N_1289);
and U2200 (N_2200,N_1421,N_1198);
and U2201 (N_2201,N_1836,N_1820);
xor U2202 (N_2202,N_1516,N_1766);
xor U2203 (N_2203,N_1439,N_1958);
xnor U2204 (N_2204,N_1542,N_1474);
and U2205 (N_2205,N_1329,N_1022);
xnor U2206 (N_2206,N_1187,N_1306);
and U2207 (N_2207,N_1926,N_1380);
nand U2208 (N_2208,N_1406,N_1251);
nand U2209 (N_2209,N_1244,N_1577);
nor U2210 (N_2210,N_1997,N_1931);
and U2211 (N_2211,N_1246,N_1110);
or U2212 (N_2212,N_1218,N_1920);
and U2213 (N_2213,N_1810,N_1119);
and U2214 (N_2214,N_1030,N_1693);
xnor U2215 (N_2215,N_1819,N_1070);
xor U2216 (N_2216,N_1419,N_1263);
and U2217 (N_2217,N_1265,N_1375);
or U2218 (N_2218,N_1621,N_1768);
nand U2219 (N_2219,N_1551,N_1826);
nand U2220 (N_2220,N_1000,N_1944);
or U2221 (N_2221,N_1735,N_1602);
nor U2222 (N_2222,N_1537,N_1731);
and U2223 (N_2223,N_1481,N_1595);
nor U2224 (N_2224,N_1250,N_1418);
or U2225 (N_2225,N_1556,N_1707);
xnor U2226 (N_2226,N_1596,N_1376);
nand U2227 (N_2227,N_1701,N_1332);
nand U2228 (N_2228,N_1478,N_1486);
and U2229 (N_2229,N_1495,N_1541);
xnor U2230 (N_2230,N_1222,N_1403);
xor U2231 (N_2231,N_1716,N_1024);
and U2232 (N_2232,N_1143,N_1795);
or U2233 (N_2233,N_1500,N_1713);
xor U2234 (N_2234,N_1281,N_1431);
and U2235 (N_2235,N_1643,N_1518);
or U2236 (N_2236,N_1346,N_1635);
or U2237 (N_2237,N_1248,N_1715);
and U2238 (N_2238,N_1607,N_1646);
xor U2239 (N_2239,N_1059,N_1645);
nor U2240 (N_2240,N_1072,N_1718);
nand U2241 (N_2241,N_1648,N_1231);
xor U2242 (N_2242,N_1857,N_1345);
or U2243 (N_2243,N_1652,N_1192);
or U2244 (N_2244,N_1374,N_1976);
xnor U2245 (N_2245,N_1149,N_1815);
nand U2246 (N_2246,N_1425,N_1107);
xnor U2247 (N_2247,N_1755,N_1697);
and U2248 (N_2248,N_1069,N_1832);
and U2249 (N_2249,N_1962,N_1043);
and U2250 (N_2250,N_1367,N_1651);
nor U2251 (N_2251,N_1597,N_1924);
nor U2252 (N_2252,N_1200,N_1333);
nor U2253 (N_2253,N_1591,N_1703);
nand U2254 (N_2254,N_1925,N_1290);
and U2255 (N_2255,N_1830,N_1838);
nor U2256 (N_2256,N_1987,N_1647);
nand U2257 (N_2257,N_1206,N_1161);
nand U2258 (N_2258,N_1354,N_1135);
nor U2259 (N_2259,N_1443,N_1720);
nand U2260 (N_2260,N_1981,N_1321);
nand U2261 (N_2261,N_1199,N_1463);
nor U2262 (N_2262,N_1343,N_1656);
nand U2263 (N_2263,N_1876,N_1052);
nor U2264 (N_2264,N_1618,N_1612);
xor U2265 (N_2265,N_1155,N_1945);
nor U2266 (N_2266,N_1893,N_1822);
xnor U2267 (N_2267,N_1284,N_1903);
nand U2268 (N_2268,N_1472,N_1415);
nor U2269 (N_2269,N_1866,N_1971);
nor U2270 (N_2270,N_1038,N_1106);
nand U2271 (N_2271,N_1451,N_1058);
or U2272 (N_2272,N_1756,N_1998);
or U2273 (N_2273,N_1460,N_1835);
or U2274 (N_2274,N_1593,N_1324);
xnor U2275 (N_2275,N_1083,N_1552);
xnor U2276 (N_2276,N_1390,N_1040);
nand U2277 (N_2277,N_1470,N_1868);
or U2278 (N_2278,N_1267,N_1002);
nand U2279 (N_2279,N_1744,N_1079);
nor U2280 (N_2280,N_1286,N_1026);
nor U2281 (N_2281,N_1954,N_1982);
or U2282 (N_2282,N_1037,N_1243);
and U2283 (N_2283,N_1572,N_1960);
nor U2284 (N_2284,N_1680,N_1933);
xor U2285 (N_2285,N_1100,N_1366);
and U2286 (N_2286,N_1689,N_1014);
nor U2287 (N_2287,N_1454,N_1547);
and U2288 (N_2288,N_1850,N_1430);
and U2289 (N_2289,N_1175,N_1065);
or U2290 (N_2290,N_1861,N_1806);
xor U2291 (N_2291,N_1385,N_1862);
and U2292 (N_2292,N_1294,N_1675);
nor U2293 (N_2293,N_1056,N_1587);
and U2294 (N_2294,N_1314,N_1502);
and U2295 (N_2295,N_1888,N_1741);
nor U2296 (N_2296,N_1303,N_1409);
nand U2297 (N_2297,N_1781,N_1031);
and U2298 (N_2298,N_1560,N_1341);
nor U2299 (N_2299,N_1530,N_1169);
nand U2300 (N_2300,N_1739,N_1217);
xor U2301 (N_2301,N_1794,N_1821);
nand U2302 (N_2302,N_1313,N_1939);
nor U2303 (N_2303,N_1441,N_1839);
nor U2304 (N_2304,N_1514,N_1604);
or U2305 (N_2305,N_1034,N_1907);
nand U2306 (N_2306,N_1125,N_1445);
or U2307 (N_2307,N_1450,N_1814);
or U2308 (N_2308,N_1594,N_1123);
or U2309 (N_2309,N_1818,N_1696);
or U2310 (N_2310,N_1157,N_1455);
xnor U2311 (N_2311,N_1670,N_1389);
xor U2312 (N_2312,N_1365,N_1853);
nand U2313 (N_2313,N_1129,N_1588);
and U2314 (N_2314,N_1683,N_1316);
xor U2315 (N_2315,N_1229,N_1833);
nor U2316 (N_2316,N_1027,N_1259);
or U2317 (N_2317,N_1152,N_1245);
or U2318 (N_2318,N_1752,N_1895);
and U2319 (N_2319,N_1897,N_1177);
and U2320 (N_2320,N_1138,N_1360);
and U2321 (N_2321,N_1865,N_1071);
or U2322 (N_2322,N_1347,N_1545);
and U2323 (N_2323,N_1230,N_1616);
xnor U2324 (N_2324,N_1797,N_1483);
or U2325 (N_2325,N_1790,N_1061);
and U2326 (N_2326,N_1649,N_1882);
or U2327 (N_2327,N_1432,N_1721);
nand U2328 (N_2328,N_1825,N_1557);
and U2329 (N_2329,N_1301,N_1204);
xor U2330 (N_2330,N_1695,N_1181);
and U2331 (N_2331,N_1957,N_1131);
and U2332 (N_2332,N_1134,N_1372);
and U2333 (N_2333,N_1256,N_1874);
and U2334 (N_2334,N_1881,N_1803);
xnor U2335 (N_2335,N_1711,N_1429);
xnor U2336 (N_2336,N_1817,N_1062);
or U2337 (N_2337,N_1270,N_1399);
xnor U2338 (N_2338,N_1461,N_1496);
or U2339 (N_2339,N_1590,N_1568);
nor U2340 (N_2340,N_1039,N_1377);
or U2341 (N_2341,N_1278,N_1426);
nand U2342 (N_2342,N_1048,N_1224);
nor U2343 (N_2343,N_1917,N_1684);
nor U2344 (N_2344,N_1033,N_1051);
or U2345 (N_2345,N_1809,N_1264);
xor U2346 (N_2346,N_1393,N_1378);
or U2347 (N_2347,N_1636,N_1162);
xnor U2348 (N_2348,N_1527,N_1834);
or U2349 (N_2349,N_1558,N_1416);
nand U2350 (N_2350,N_1722,N_1896);
and U2351 (N_2351,N_1121,N_1523);
and U2352 (N_2352,N_1613,N_1238);
nor U2353 (N_2353,N_1044,N_1225);
xnor U2354 (N_2354,N_1113,N_1574);
nand U2355 (N_2355,N_1609,N_1124);
and U2356 (N_2356,N_1465,N_1964);
and U2357 (N_2357,N_1359,N_1326);
nand U2358 (N_2358,N_1508,N_1269);
or U2359 (N_2359,N_1216,N_1057);
or U2360 (N_2360,N_1993,N_1494);
nor U2361 (N_2361,N_1665,N_1544);
nor U2362 (N_2362,N_1858,N_1786);
nand U2363 (N_2363,N_1179,N_1193);
and U2364 (N_2364,N_1277,N_1282);
nor U2365 (N_2365,N_1754,N_1908);
and U2366 (N_2366,N_1950,N_1395);
or U2367 (N_2367,N_1967,N_1532);
and U2368 (N_2368,N_1400,N_1867);
nand U2369 (N_2369,N_1885,N_1909);
nand U2370 (N_2370,N_1775,N_1252);
nand U2371 (N_2371,N_1528,N_1221);
nand U2372 (N_2372,N_1126,N_1063);
nand U2373 (N_2373,N_1584,N_1457);
and U2374 (N_2374,N_1535,N_1295);
and U2375 (N_2375,N_1916,N_1887);
nor U2376 (N_2376,N_1173,N_1167);
or U2377 (N_2377,N_1087,N_1364);
nand U2378 (N_2378,N_1573,N_1849);
and U2379 (N_2379,N_1202,N_1943);
xor U2380 (N_2380,N_1747,N_1357);
and U2381 (N_2381,N_1717,N_1952);
or U2382 (N_2382,N_1335,N_1704);
and U2383 (N_2383,N_1291,N_1555);
xnor U2384 (N_2384,N_1237,N_1759);
xnor U2385 (N_2385,N_1694,N_1736);
or U2386 (N_2386,N_1677,N_1910);
nand U2387 (N_2387,N_1283,N_1223);
xor U2388 (N_2388,N_1234,N_1036);
nand U2389 (N_2389,N_1285,N_1292);
and U2390 (N_2390,N_1012,N_1767);
nor U2391 (N_2391,N_1883,N_1513);
and U2392 (N_2392,N_1148,N_1183);
and U2393 (N_2393,N_1253,N_1254);
nor U2394 (N_2394,N_1746,N_1946);
nor U2395 (N_2395,N_1210,N_1723);
nor U2396 (N_2396,N_1841,N_1863);
nand U2397 (N_2397,N_1215,N_1344);
or U2398 (N_2398,N_1827,N_1117);
nand U2399 (N_2399,N_1601,N_1049);
or U2400 (N_2400,N_1050,N_1410);
nor U2401 (N_2401,N_1055,N_1511);
and U2402 (N_2402,N_1213,N_1889);
or U2403 (N_2403,N_1401,N_1095);
or U2404 (N_2404,N_1628,N_1605);
nand U2405 (N_2405,N_1227,N_1168);
or U2406 (N_2406,N_1413,N_1318);
nand U2407 (N_2407,N_1761,N_1777);
or U2408 (N_2408,N_1525,N_1536);
or U2409 (N_2409,N_1147,N_1811);
nand U2410 (N_2410,N_1880,N_1576);
and U2411 (N_2411,N_1194,N_1127);
nor U2412 (N_2412,N_1176,N_1067);
xor U2413 (N_2413,N_1859,N_1664);
and U2414 (N_2414,N_1639,N_1109);
nand U2415 (N_2415,N_1271,N_1990);
nor U2416 (N_2416,N_1856,N_1068);
xor U2417 (N_2417,N_1174,N_1592);
and U2418 (N_2418,N_1302,N_1482);
xnor U2419 (N_2419,N_1921,N_1045);
and U2420 (N_2420,N_1501,N_1808);
nor U2421 (N_2421,N_1420,N_1163);
xor U2422 (N_2422,N_1349,N_1629);
and U2423 (N_2423,N_1077,N_1655);
nor U2424 (N_2424,N_1548,N_1914);
nor U2425 (N_2425,N_1444,N_1657);
xnor U2426 (N_2426,N_1904,N_1381);
nor U2427 (N_2427,N_1566,N_1351);
xnor U2428 (N_2428,N_1673,N_1305);
and U2429 (N_2429,N_1073,N_1900);
and U2430 (N_2430,N_1384,N_1363);
xnor U2431 (N_2431,N_1737,N_1315);
and U2432 (N_2432,N_1220,N_1505);
or U2433 (N_2433,N_1422,N_1802);
nor U2434 (N_2434,N_1674,N_1309);
and U2435 (N_2435,N_1260,N_1350);
nor U2436 (N_2436,N_1054,N_1001);
xnor U2437 (N_2437,N_1979,N_1705);
nand U2438 (N_2438,N_1540,N_1342);
nor U2439 (N_2439,N_1700,N_1504);
nand U2440 (N_2440,N_1725,N_1749);
or U2441 (N_2441,N_1619,N_1798);
xnor U2442 (N_2442,N_1783,N_1023);
xor U2443 (N_2443,N_1653,N_1137);
xnor U2444 (N_2444,N_1427,N_1972);
and U2445 (N_2445,N_1559,N_1182);
or U2446 (N_2446,N_1491,N_1379);
nand U2447 (N_2447,N_1459,N_1792);
and U2448 (N_2448,N_1296,N_1610);
nor U2449 (N_2449,N_1851,N_1846);
nor U2450 (N_2450,N_1308,N_1373);
nor U2451 (N_2451,N_1740,N_1699);
and U2452 (N_2452,N_1021,N_1475);
and U2453 (N_2453,N_1388,N_1008);
or U2454 (N_2454,N_1394,N_1469);
or U2455 (N_2455,N_1526,N_1209);
or U2456 (N_2456,N_1191,N_1805);
or U2457 (N_2457,N_1915,N_1398);
nor U2458 (N_2458,N_1782,N_1951);
nand U2459 (N_2459,N_1738,N_1658);
xnor U2460 (N_2460,N_1096,N_1816);
xnor U2461 (N_2461,N_1845,N_1637);
and U2462 (N_2462,N_1353,N_1671);
nand U2463 (N_2463,N_1028,N_1090);
or U2464 (N_2464,N_1007,N_1382);
or U2465 (N_2465,N_1497,N_1583);
and U2466 (N_2466,N_1473,N_1770);
or U2467 (N_2467,N_1492,N_1660);
xor U2468 (N_2468,N_1669,N_1423);
xnor U2469 (N_2469,N_1801,N_1771);
or U2470 (N_2470,N_1383,N_1662);
nand U2471 (N_2471,N_1620,N_1299);
and U2472 (N_2472,N_1842,N_1623);
nand U2473 (N_2473,N_1498,N_1638);
nand U2474 (N_2474,N_1307,N_1932);
xor U2475 (N_2475,N_1046,N_1690);
xor U2476 (N_2476,N_1261,N_1589);
nand U2477 (N_2477,N_1325,N_1015);
or U2478 (N_2478,N_1813,N_1791);
nor U2479 (N_2479,N_1320,N_1918);
nor U2480 (N_2480,N_1274,N_1102);
nor U2481 (N_2481,N_1517,N_1553);
or U2482 (N_2482,N_1207,N_1190);
and U2483 (N_2483,N_1085,N_1407);
nand U2484 (N_2484,N_1608,N_1772);
and U2485 (N_2485,N_1512,N_1886);
xor U2486 (N_2486,N_1396,N_1104);
or U2487 (N_2487,N_1433,N_1130);
xor U2488 (N_2488,N_1449,N_1624);
xnor U2489 (N_2489,N_1247,N_1800);
or U2490 (N_2490,N_1184,N_1659);
and U2491 (N_2491,N_1099,N_1936);
or U2492 (N_2492,N_1899,N_1824);
nor U2493 (N_2493,N_1322,N_1614);
nor U2494 (N_2494,N_1582,N_1141);
or U2495 (N_2495,N_1195,N_1105);
and U2496 (N_2496,N_1840,N_1630);
and U2497 (N_2497,N_1575,N_1714);
nor U2498 (N_2498,N_1966,N_1934);
or U2499 (N_2499,N_1927,N_1352);
or U2500 (N_2500,N_1807,N_1281);
nor U2501 (N_2501,N_1756,N_1289);
and U2502 (N_2502,N_1556,N_1783);
nand U2503 (N_2503,N_1616,N_1247);
nand U2504 (N_2504,N_1181,N_1119);
and U2505 (N_2505,N_1231,N_1163);
and U2506 (N_2506,N_1340,N_1651);
xnor U2507 (N_2507,N_1009,N_1770);
xnor U2508 (N_2508,N_1372,N_1472);
or U2509 (N_2509,N_1422,N_1151);
nand U2510 (N_2510,N_1524,N_1884);
nor U2511 (N_2511,N_1599,N_1577);
and U2512 (N_2512,N_1016,N_1613);
nand U2513 (N_2513,N_1479,N_1505);
nand U2514 (N_2514,N_1419,N_1832);
xor U2515 (N_2515,N_1100,N_1666);
or U2516 (N_2516,N_1768,N_1746);
nand U2517 (N_2517,N_1891,N_1942);
nor U2518 (N_2518,N_1539,N_1204);
nand U2519 (N_2519,N_1718,N_1108);
nand U2520 (N_2520,N_1050,N_1012);
xnor U2521 (N_2521,N_1520,N_1816);
and U2522 (N_2522,N_1715,N_1207);
xor U2523 (N_2523,N_1231,N_1284);
and U2524 (N_2524,N_1525,N_1315);
xnor U2525 (N_2525,N_1430,N_1759);
xnor U2526 (N_2526,N_1627,N_1003);
xor U2527 (N_2527,N_1789,N_1595);
or U2528 (N_2528,N_1158,N_1115);
or U2529 (N_2529,N_1495,N_1880);
xor U2530 (N_2530,N_1119,N_1785);
nor U2531 (N_2531,N_1489,N_1596);
and U2532 (N_2532,N_1570,N_1158);
xnor U2533 (N_2533,N_1093,N_1217);
or U2534 (N_2534,N_1014,N_1144);
or U2535 (N_2535,N_1260,N_1375);
nand U2536 (N_2536,N_1934,N_1550);
xor U2537 (N_2537,N_1817,N_1517);
xor U2538 (N_2538,N_1755,N_1240);
nand U2539 (N_2539,N_1005,N_1049);
xor U2540 (N_2540,N_1152,N_1007);
or U2541 (N_2541,N_1297,N_1156);
nor U2542 (N_2542,N_1991,N_1321);
nand U2543 (N_2543,N_1763,N_1667);
or U2544 (N_2544,N_1999,N_1190);
and U2545 (N_2545,N_1126,N_1904);
xnor U2546 (N_2546,N_1244,N_1067);
nor U2547 (N_2547,N_1130,N_1491);
and U2548 (N_2548,N_1604,N_1823);
or U2549 (N_2549,N_1556,N_1611);
xor U2550 (N_2550,N_1950,N_1017);
nand U2551 (N_2551,N_1890,N_1581);
nand U2552 (N_2552,N_1752,N_1031);
nand U2553 (N_2553,N_1581,N_1207);
nand U2554 (N_2554,N_1814,N_1452);
nor U2555 (N_2555,N_1704,N_1605);
or U2556 (N_2556,N_1473,N_1038);
or U2557 (N_2557,N_1151,N_1214);
nand U2558 (N_2558,N_1584,N_1341);
or U2559 (N_2559,N_1862,N_1572);
nor U2560 (N_2560,N_1749,N_1462);
nand U2561 (N_2561,N_1524,N_1118);
or U2562 (N_2562,N_1957,N_1165);
and U2563 (N_2563,N_1701,N_1504);
nand U2564 (N_2564,N_1061,N_1751);
or U2565 (N_2565,N_1179,N_1321);
xnor U2566 (N_2566,N_1331,N_1524);
or U2567 (N_2567,N_1729,N_1065);
and U2568 (N_2568,N_1458,N_1745);
nor U2569 (N_2569,N_1639,N_1585);
nor U2570 (N_2570,N_1161,N_1520);
nor U2571 (N_2571,N_1829,N_1921);
xor U2572 (N_2572,N_1730,N_1441);
nand U2573 (N_2573,N_1172,N_1783);
xor U2574 (N_2574,N_1225,N_1409);
nand U2575 (N_2575,N_1759,N_1802);
and U2576 (N_2576,N_1134,N_1815);
nand U2577 (N_2577,N_1362,N_1369);
nor U2578 (N_2578,N_1025,N_1870);
or U2579 (N_2579,N_1583,N_1323);
nor U2580 (N_2580,N_1304,N_1615);
and U2581 (N_2581,N_1414,N_1031);
xor U2582 (N_2582,N_1542,N_1118);
nand U2583 (N_2583,N_1832,N_1353);
nand U2584 (N_2584,N_1976,N_1769);
or U2585 (N_2585,N_1998,N_1096);
nor U2586 (N_2586,N_1973,N_1091);
or U2587 (N_2587,N_1478,N_1907);
and U2588 (N_2588,N_1543,N_1084);
and U2589 (N_2589,N_1868,N_1250);
xor U2590 (N_2590,N_1069,N_1856);
nor U2591 (N_2591,N_1768,N_1699);
nor U2592 (N_2592,N_1822,N_1055);
xnor U2593 (N_2593,N_1193,N_1369);
xor U2594 (N_2594,N_1291,N_1673);
nor U2595 (N_2595,N_1349,N_1918);
nor U2596 (N_2596,N_1982,N_1917);
nand U2597 (N_2597,N_1712,N_1065);
nor U2598 (N_2598,N_1601,N_1971);
xnor U2599 (N_2599,N_1767,N_1235);
xnor U2600 (N_2600,N_1291,N_1688);
xnor U2601 (N_2601,N_1011,N_1216);
xor U2602 (N_2602,N_1344,N_1496);
xor U2603 (N_2603,N_1674,N_1863);
xor U2604 (N_2604,N_1255,N_1709);
and U2605 (N_2605,N_1769,N_1217);
nand U2606 (N_2606,N_1900,N_1131);
nand U2607 (N_2607,N_1168,N_1180);
nor U2608 (N_2608,N_1084,N_1802);
xnor U2609 (N_2609,N_1519,N_1059);
nor U2610 (N_2610,N_1326,N_1940);
and U2611 (N_2611,N_1405,N_1460);
nor U2612 (N_2612,N_1233,N_1268);
or U2613 (N_2613,N_1392,N_1266);
and U2614 (N_2614,N_1030,N_1073);
nor U2615 (N_2615,N_1306,N_1041);
nand U2616 (N_2616,N_1392,N_1707);
and U2617 (N_2617,N_1339,N_1190);
nor U2618 (N_2618,N_1611,N_1067);
or U2619 (N_2619,N_1842,N_1840);
xor U2620 (N_2620,N_1578,N_1155);
or U2621 (N_2621,N_1512,N_1836);
nor U2622 (N_2622,N_1962,N_1854);
or U2623 (N_2623,N_1449,N_1789);
xnor U2624 (N_2624,N_1431,N_1954);
nor U2625 (N_2625,N_1319,N_1005);
or U2626 (N_2626,N_1593,N_1077);
nor U2627 (N_2627,N_1980,N_1643);
and U2628 (N_2628,N_1868,N_1881);
nor U2629 (N_2629,N_1260,N_1294);
nand U2630 (N_2630,N_1576,N_1085);
and U2631 (N_2631,N_1263,N_1038);
xnor U2632 (N_2632,N_1132,N_1585);
xor U2633 (N_2633,N_1966,N_1384);
and U2634 (N_2634,N_1174,N_1881);
nor U2635 (N_2635,N_1397,N_1470);
and U2636 (N_2636,N_1505,N_1114);
xnor U2637 (N_2637,N_1598,N_1113);
xor U2638 (N_2638,N_1808,N_1833);
nor U2639 (N_2639,N_1667,N_1219);
nand U2640 (N_2640,N_1868,N_1957);
or U2641 (N_2641,N_1897,N_1153);
xor U2642 (N_2642,N_1588,N_1223);
xnor U2643 (N_2643,N_1809,N_1888);
and U2644 (N_2644,N_1909,N_1488);
nor U2645 (N_2645,N_1129,N_1080);
or U2646 (N_2646,N_1648,N_1062);
and U2647 (N_2647,N_1051,N_1112);
and U2648 (N_2648,N_1778,N_1509);
nor U2649 (N_2649,N_1355,N_1103);
and U2650 (N_2650,N_1559,N_1691);
xor U2651 (N_2651,N_1389,N_1107);
xnor U2652 (N_2652,N_1459,N_1319);
or U2653 (N_2653,N_1083,N_1989);
or U2654 (N_2654,N_1117,N_1497);
nor U2655 (N_2655,N_1688,N_1571);
and U2656 (N_2656,N_1837,N_1180);
or U2657 (N_2657,N_1214,N_1221);
nor U2658 (N_2658,N_1108,N_1309);
nand U2659 (N_2659,N_1824,N_1339);
or U2660 (N_2660,N_1724,N_1394);
and U2661 (N_2661,N_1134,N_1944);
nand U2662 (N_2662,N_1227,N_1273);
nand U2663 (N_2663,N_1023,N_1933);
xor U2664 (N_2664,N_1739,N_1586);
xor U2665 (N_2665,N_1154,N_1425);
xnor U2666 (N_2666,N_1858,N_1557);
nor U2667 (N_2667,N_1754,N_1344);
nand U2668 (N_2668,N_1120,N_1885);
and U2669 (N_2669,N_1869,N_1954);
nor U2670 (N_2670,N_1158,N_1489);
and U2671 (N_2671,N_1947,N_1483);
or U2672 (N_2672,N_1778,N_1278);
and U2673 (N_2673,N_1564,N_1133);
xor U2674 (N_2674,N_1016,N_1569);
nor U2675 (N_2675,N_1625,N_1510);
xor U2676 (N_2676,N_1073,N_1588);
xor U2677 (N_2677,N_1485,N_1772);
nand U2678 (N_2678,N_1407,N_1273);
xor U2679 (N_2679,N_1593,N_1957);
xor U2680 (N_2680,N_1874,N_1468);
nand U2681 (N_2681,N_1960,N_1756);
xnor U2682 (N_2682,N_1103,N_1087);
or U2683 (N_2683,N_1898,N_1570);
or U2684 (N_2684,N_1926,N_1190);
xnor U2685 (N_2685,N_1071,N_1373);
xor U2686 (N_2686,N_1010,N_1498);
nor U2687 (N_2687,N_1793,N_1555);
nand U2688 (N_2688,N_1525,N_1715);
and U2689 (N_2689,N_1740,N_1866);
nor U2690 (N_2690,N_1281,N_1112);
nand U2691 (N_2691,N_1974,N_1323);
nand U2692 (N_2692,N_1777,N_1173);
nor U2693 (N_2693,N_1344,N_1532);
nor U2694 (N_2694,N_1175,N_1320);
or U2695 (N_2695,N_1011,N_1252);
xor U2696 (N_2696,N_1236,N_1301);
xnor U2697 (N_2697,N_1542,N_1639);
and U2698 (N_2698,N_1560,N_1177);
nand U2699 (N_2699,N_1934,N_1209);
and U2700 (N_2700,N_1810,N_1287);
nor U2701 (N_2701,N_1581,N_1675);
or U2702 (N_2702,N_1411,N_1557);
xnor U2703 (N_2703,N_1820,N_1057);
xor U2704 (N_2704,N_1053,N_1112);
nand U2705 (N_2705,N_1448,N_1661);
or U2706 (N_2706,N_1591,N_1881);
or U2707 (N_2707,N_1309,N_1925);
or U2708 (N_2708,N_1366,N_1745);
nand U2709 (N_2709,N_1963,N_1798);
nand U2710 (N_2710,N_1390,N_1448);
nor U2711 (N_2711,N_1236,N_1929);
nor U2712 (N_2712,N_1524,N_1690);
nor U2713 (N_2713,N_1249,N_1275);
or U2714 (N_2714,N_1250,N_1255);
and U2715 (N_2715,N_1463,N_1702);
or U2716 (N_2716,N_1934,N_1302);
or U2717 (N_2717,N_1862,N_1023);
and U2718 (N_2718,N_1338,N_1138);
nor U2719 (N_2719,N_1048,N_1723);
and U2720 (N_2720,N_1824,N_1368);
xor U2721 (N_2721,N_1245,N_1049);
xor U2722 (N_2722,N_1147,N_1116);
nor U2723 (N_2723,N_1639,N_1751);
xor U2724 (N_2724,N_1963,N_1042);
and U2725 (N_2725,N_1487,N_1588);
nand U2726 (N_2726,N_1402,N_1807);
and U2727 (N_2727,N_1541,N_1907);
xor U2728 (N_2728,N_1095,N_1233);
or U2729 (N_2729,N_1894,N_1326);
and U2730 (N_2730,N_1014,N_1791);
and U2731 (N_2731,N_1835,N_1421);
and U2732 (N_2732,N_1622,N_1189);
and U2733 (N_2733,N_1738,N_1917);
and U2734 (N_2734,N_1777,N_1836);
and U2735 (N_2735,N_1431,N_1796);
nand U2736 (N_2736,N_1885,N_1507);
xnor U2737 (N_2737,N_1179,N_1715);
or U2738 (N_2738,N_1859,N_1138);
and U2739 (N_2739,N_1426,N_1881);
nor U2740 (N_2740,N_1985,N_1899);
or U2741 (N_2741,N_1922,N_1326);
and U2742 (N_2742,N_1943,N_1399);
nor U2743 (N_2743,N_1300,N_1778);
xnor U2744 (N_2744,N_1283,N_1804);
nand U2745 (N_2745,N_1537,N_1687);
nor U2746 (N_2746,N_1951,N_1082);
and U2747 (N_2747,N_1992,N_1021);
or U2748 (N_2748,N_1124,N_1133);
xor U2749 (N_2749,N_1322,N_1507);
and U2750 (N_2750,N_1127,N_1761);
nand U2751 (N_2751,N_1081,N_1857);
nand U2752 (N_2752,N_1092,N_1419);
nor U2753 (N_2753,N_1898,N_1016);
xnor U2754 (N_2754,N_1651,N_1551);
and U2755 (N_2755,N_1704,N_1427);
nor U2756 (N_2756,N_1192,N_1895);
xor U2757 (N_2757,N_1470,N_1892);
and U2758 (N_2758,N_1166,N_1528);
nor U2759 (N_2759,N_1869,N_1632);
nor U2760 (N_2760,N_1383,N_1461);
or U2761 (N_2761,N_1047,N_1039);
nand U2762 (N_2762,N_1010,N_1608);
and U2763 (N_2763,N_1819,N_1268);
or U2764 (N_2764,N_1815,N_1657);
and U2765 (N_2765,N_1625,N_1412);
and U2766 (N_2766,N_1941,N_1598);
or U2767 (N_2767,N_1708,N_1175);
and U2768 (N_2768,N_1644,N_1562);
or U2769 (N_2769,N_1439,N_1490);
xor U2770 (N_2770,N_1098,N_1928);
nor U2771 (N_2771,N_1918,N_1073);
nor U2772 (N_2772,N_1080,N_1605);
or U2773 (N_2773,N_1712,N_1317);
nor U2774 (N_2774,N_1050,N_1802);
and U2775 (N_2775,N_1011,N_1117);
xnor U2776 (N_2776,N_1937,N_1331);
nor U2777 (N_2777,N_1248,N_1699);
nor U2778 (N_2778,N_1558,N_1693);
nor U2779 (N_2779,N_1813,N_1804);
nor U2780 (N_2780,N_1589,N_1901);
nor U2781 (N_2781,N_1624,N_1121);
and U2782 (N_2782,N_1892,N_1055);
nor U2783 (N_2783,N_1629,N_1706);
and U2784 (N_2784,N_1818,N_1024);
nand U2785 (N_2785,N_1266,N_1238);
nand U2786 (N_2786,N_1035,N_1472);
and U2787 (N_2787,N_1671,N_1563);
and U2788 (N_2788,N_1067,N_1216);
nor U2789 (N_2789,N_1782,N_1778);
or U2790 (N_2790,N_1266,N_1048);
nand U2791 (N_2791,N_1843,N_1048);
xor U2792 (N_2792,N_1746,N_1139);
nor U2793 (N_2793,N_1251,N_1879);
and U2794 (N_2794,N_1066,N_1526);
nor U2795 (N_2795,N_1296,N_1628);
nand U2796 (N_2796,N_1496,N_1803);
or U2797 (N_2797,N_1327,N_1087);
nor U2798 (N_2798,N_1747,N_1144);
nand U2799 (N_2799,N_1246,N_1728);
or U2800 (N_2800,N_1732,N_1995);
and U2801 (N_2801,N_1891,N_1223);
and U2802 (N_2802,N_1135,N_1167);
and U2803 (N_2803,N_1154,N_1403);
xnor U2804 (N_2804,N_1903,N_1057);
nor U2805 (N_2805,N_1755,N_1824);
nand U2806 (N_2806,N_1005,N_1583);
and U2807 (N_2807,N_1952,N_1704);
nand U2808 (N_2808,N_1207,N_1439);
xnor U2809 (N_2809,N_1855,N_1808);
xor U2810 (N_2810,N_1877,N_1939);
xor U2811 (N_2811,N_1731,N_1381);
and U2812 (N_2812,N_1368,N_1423);
and U2813 (N_2813,N_1461,N_1443);
nor U2814 (N_2814,N_1322,N_1485);
xnor U2815 (N_2815,N_1785,N_1843);
nor U2816 (N_2816,N_1221,N_1370);
and U2817 (N_2817,N_1323,N_1940);
nor U2818 (N_2818,N_1541,N_1396);
nor U2819 (N_2819,N_1242,N_1700);
nand U2820 (N_2820,N_1842,N_1654);
and U2821 (N_2821,N_1361,N_1267);
xnor U2822 (N_2822,N_1946,N_1945);
or U2823 (N_2823,N_1838,N_1686);
nand U2824 (N_2824,N_1086,N_1496);
or U2825 (N_2825,N_1984,N_1155);
or U2826 (N_2826,N_1040,N_1998);
and U2827 (N_2827,N_1601,N_1603);
nor U2828 (N_2828,N_1924,N_1970);
or U2829 (N_2829,N_1910,N_1632);
and U2830 (N_2830,N_1470,N_1929);
and U2831 (N_2831,N_1314,N_1208);
and U2832 (N_2832,N_1043,N_1032);
xnor U2833 (N_2833,N_1475,N_1788);
and U2834 (N_2834,N_1493,N_1272);
nor U2835 (N_2835,N_1367,N_1892);
xnor U2836 (N_2836,N_1326,N_1532);
nor U2837 (N_2837,N_1297,N_1300);
nand U2838 (N_2838,N_1311,N_1044);
nand U2839 (N_2839,N_1766,N_1406);
and U2840 (N_2840,N_1301,N_1660);
nand U2841 (N_2841,N_1653,N_1013);
nand U2842 (N_2842,N_1055,N_1544);
nand U2843 (N_2843,N_1013,N_1756);
nor U2844 (N_2844,N_1116,N_1644);
or U2845 (N_2845,N_1654,N_1003);
xor U2846 (N_2846,N_1369,N_1790);
nand U2847 (N_2847,N_1884,N_1506);
and U2848 (N_2848,N_1230,N_1597);
nor U2849 (N_2849,N_1875,N_1550);
xnor U2850 (N_2850,N_1528,N_1853);
xnor U2851 (N_2851,N_1969,N_1274);
nand U2852 (N_2852,N_1421,N_1756);
xor U2853 (N_2853,N_1430,N_1701);
or U2854 (N_2854,N_1592,N_1531);
xnor U2855 (N_2855,N_1484,N_1804);
or U2856 (N_2856,N_1088,N_1253);
or U2857 (N_2857,N_1014,N_1216);
nand U2858 (N_2858,N_1326,N_1530);
nor U2859 (N_2859,N_1565,N_1530);
or U2860 (N_2860,N_1521,N_1546);
nor U2861 (N_2861,N_1247,N_1589);
and U2862 (N_2862,N_1456,N_1290);
and U2863 (N_2863,N_1383,N_1625);
and U2864 (N_2864,N_1614,N_1427);
or U2865 (N_2865,N_1811,N_1991);
nand U2866 (N_2866,N_1263,N_1567);
and U2867 (N_2867,N_1500,N_1554);
xnor U2868 (N_2868,N_1445,N_1843);
nor U2869 (N_2869,N_1449,N_1178);
and U2870 (N_2870,N_1818,N_1691);
and U2871 (N_2871,N_1707,N_1312);
xnor U2872 (N_2872,N_1251,N_1157);
nand U2873 (N_2873,N_1960,N_1538);
xnor U2874 (N_2874,N_1858,N_1996);
or U2875 (N_2875,N_1480,N_1445);
or U2876 (N_2876,N_1974,N_1129);
nand U2877 (N_2877,N_1793,N_1514);
or U2878 (N_2878,N_1125,N_1403);
or U2879 (N_2879,N_1085,N_1778);
nand U2880 (N_2880,N_1968,N_1547);
and U2881 (N_2881,N_1531,N_1702);
or U2882 (N_2882,N_1664,N_1011);
nor U2883 (N_2883,N_1967,N_1386);
nand U2884 (N_2884,N_1076,N_1539);
nor U2885 (N_2885,N_1612,N_1720);
nor U2886 (N_2886,N_1349,N_1575);
xnor U2887 (N_2887,N_1308,N_1624);
and U2888 (N_2888,N_1807,N_1308);
and U2889 (N_2889,N_1691,N_1633);
nor U2890 (N_2890,N_1378,N_1240);
and U2891 (N_2891,N_1191,N_1382);
or U2892 (N_2892,N_1567,N_1003);
and U2893 (N_2893,N_1265,N_1895);
nor U2894 (N_2894,N_1241,N_1760);
or U2895 (N_2895,N_1638,N_1318);
or U2896 (N_2896,N_1924,N_1091);
nor U2897 (N_2897,N_1925,N_1613);
nand U2898 (N_2898,N_1358,N_1771);
or U2899 (N_2899,N_1967,N_1340);
nor U2900 (N_2900,N_1686,N_1630);
and U2901 (N_2901,N_1958,N_1594);
and U2902 (N_2902,N_1475,N_1312);
and U2903 (N_2903,N_1420,N_1317);
xor U2904 (N_2904,N_1156,N_1488);
or U2905 (N_2905,N_1588,N_1035);
or U2906 (N_2906,N_1734,N_1130);
and U2907 (N_2907,N_1244,N_1853);
xor U2908 (N_2908,N_1986,N_1905);
nor U2909 (N_2909,N_1985,N_1901);
and U2910 (N_2910,N_1427,N_1391);
and U2911 (N_2911,N_1258,N_1617);
or U2912 (N_2912,N_1126,N_1040);
or U2913 (N_2913,N_1488,N_1667);
nand U2914 (N_2914,N_1254,N_1839);
and U2915 (N_2915,N_1958,N_1104);
nand U2916 (N_2916,N_1004,N_1983);
nand U2917 (N_2917,N_1015,N_1452);
nand U2918 (N_2918,N_1436,N_1227);
xor U2919 (N_2919,N_1245,N_1180);
nand U2920 (N_2920,N_1021,N_1486);
xor U2921 (N_2921,N_1267,N_1623);
nand U2922 (N_2922,N_1340,N_1033);
nor U2923 (N_2923,N_1764,N_1035);
xnor U2924 (N_2924,N_1037,N_1091);
nor U2925 (N_2925,N_1466,N_1135);
or U2926 (N_2926,N_1543,N_1472);
and U2927 (N_2927,N_1936,N_1830);
or U2928 (N_2928,N_1256,N_1811);
xnor U2929 (N_2929,N_1773,N_1928);
xnor U2930 (N_2930,N_1298,N_1644);
or U2931 (N_2931,N_1759,N_1102);
and U2932 (N_2932,N_1355,N_1940);
or U2933 (N_2933,N_1569,N_1961);
or U2934 (N_2934,N_1565,N_1204);
or U2935 (N_2935,N_1287,N_1971);
xnor U2936 (N_2936,N_1805,N_1150);
or U2937 (N_2937,N_1334,N_1176);
nand U2938 (N_2938,N_1414,N_1206);
nand U2939 (N_2939,N_1341,N_1441);
or U2940 (N_2940,N_1268,N_1033);
xor U2941 (N_2941,N_1485,N_1169);
or U2942 (N_2942,N_1256,N_1583);
or U2943 (N_2943,N_1171,N_1265);
xor U2944 (N_2944,N_1808,N_1067);
or U2945 (N_2945,N_1355,N_1690);
nor U2946 (N_2946,N_1884,N_1187);
xnor U2947 (N_2947,N_1314,N_1936);
xnor U2948 (N_2948,N_1674,N_1250);
nor U2949 (N_2949,N_1409,N_1573);
or U2950 (N_2950,N_1065,N_1375);
xnor U2951 (N_2951,N_1311,N_1962);
or U2952 (N_2952,N_1437,N_1655);
and U2953 (N_2953,N_1019,N_1009);
or U2954 (N_2954,N_1937,N_1452);
xnor U2955 (N_2955,N_1589,N_1120);
nand U2956 (N_2956,N_1642,N_1086);
xnor U2957 (N_2957,N_1087,N_1284);
and U2958 (N_2958,N_1515,N_1372);
xnor U2959 (N_2959,N_1106,N_1617);
and U2960 (N_2960,N_1783,N_1041);
nand U2961 (N_2961,N_1712,N_1237);
nor U2962 (N_2962,N_1722,N_1822);
or U2963 (N_2963,N_1266,N_1636);
and U2964 (N_2964,N_1485,N_1183);
or U2965 (N_2965,N_1596,N_1206);
or U2966 (N_2966,N_1125,N_1563);
nor U2967 (N_2967,N_1234,N_1376);
nor U2968 (N_2968,N_1114,N_1362);
xnor U2969 (N_2969,N_1197,N_1610);
and U2970 (N_2970,N_1009,N_1464);
nand U2971 (N_2971,N_1488,N_1568);
nor U2972 (N_2972,N_1631,N_1178);
or U2973 (N_2973,N_1169,N_1391);
or U2974 (N_2974,N_1266,N_1734);
nand U2975 (N_2975,N_1100,N_1082);
and U2976 (N_2976,N_1225,N_1682);
nand U2977 (N_2977,N_1015,N_1950);
nand U2978 (N_2978,N_1342,N_1446);
and U2979 (N_2979,N_1853,N_1683);
or U2980 (N_2980,N_1531,N_1549);
xor U2981 (N_2981,N_1169,N_1212);
or U2982 (N_2982,N_1064,N_1951);
nor U2983 (N_2983,N_1293,N_1709);
nand U2984 (N_2984,N_1439,N_1141);
nand U2985 (N_2985,N_1638,N_1307);
nand U2986 (N_2986,N_1833,N_1157);
xor U2987 (N_2987,N_1361,N_1348);
nor U2988 (N_2988,N_1213,N_1442);
xor U2989 (N_2989,N_1278,N_1990);
nand U2990 (N_2990,N_1950,N_1689);
and U2991 (N_2991,N_1117,N_1511);
and U2992 (N_2992,N_1579,N_1753);
or U2993 (N_2993,N_1665,N_1647);
nand U2994 (N_2994,N_1468,N_1019);
xor U2995 (N_2995,N_1866,N_1434);
or U2996 (N_2996,N_1404,N_1954);
nand U2997 (N_2997,N_1249,N_1718);
and U2998 (N_2998,N_1036,N_1476);
nand U2999 (N_2999,N_1982,N_1539);
nand U3000 (N_3000,N_2319,N_2136);
nor U3001 (N_3001,N_2423,N_2882);
nand U3002 (N_3002,N_2913,N_2756);
or U3003 (N_3003,N_2255,N_2888);
or U3004 (N_3004,N_2783,N_2320);
and U3005 (N_3005,N_2724,N_2003);
and U3006 (N_3006,N_2772,N_2037);
xnor U3007 (N_3007,N_2025,N_2899);
and U3008 (N_3008,N_2259,N_2241);
nand U3009 (N_3009,N_2199,N_2696);
nand U3010 (N_3010,N_2642,N_2971);
xor U3011 (N_3011,N_2018,N_2307);
and U3012 (N_3012,N_2252,N_2089);
nor U3013 (N_3013,N_2180,N_2655);
or U3014 (N_3014,N_2308,N_2538);
and U3015 (N_3015,N_2121,N_2457);
nor U3016 (N_3016,N_2851,N_2138);
nor U3017 (N_3017,N_2251,N_2814);
nor U3018 (N_3018,N_2773,N_2948);
xnor U3019 (N_3019,N_2493,N_2631);
nor U3020 (N_3020,N_2049,N_2210);
nor U3021 (N_3021,N_2641,N_2977);
nor U3022 (N_3022,N_2467,N_2455);
nor U3023 (N_3023,N_2329,N_2221);
or U3024 (N_3024,N_2767,N_2539);
nand U3025 (N_3025,N_2123,N_2420);
nand U3026 (N_3026,N_2050,N_2427);
nand U3027 (N_3027,N_2325,N_2609);
nor U3028 (N_3028,N_2793,N_2379);
xor U3029 (N_3029,N_2605,N_2987);
nand U3030 (N_3030,N_2113,N_2440);
and U3031 (N_3031,N_2574,N_2834);
nor U3032 (N_3032,N_2151,N_2410);
nand U3033 (N_3033,N_2600,N_2906);
or U3034 (N_3034,N_2686,N_2964);
nand U3035 (N_3035,N_2230,N_2984);
nor U3036 (N_3036,N_2927,N_2020);
nand U3037 (N_3037,N_2349,N_2026);
xnor U3038 (N_3038,N_2106,N_2816);
nand U3039 (N_3039,N_2873,N_2351);
and U3040 (N_3040,N_2544,N_2664);
nor U3041 (N_3041,N_2378,N_2700);
or U3042 (N_3042,N_2640,N_2802);
nor U3043 (N_3043,N_2891,N_2333);
xnor U3044 (N_3044,N_2261,N_2108);
nand U3045 (N_3045,N_2189,N_2957);
and U3046 (N_3046,N_2334,N_2327);
nand U3047 (N_3047,N_2181,N_2921);
and U3048 (N_3048,N_2549,N_2278);
xnor U3049 (N_3049,N_2552,N_2069);
nand U3050 (N_3050,N_2595,N_2155);
xor U3051 (N_3051,N_2125,N_2200);
nand U3052 (N_3052,N_2736,N_2279);
or U3053 (N_3053,N_2548,N_2706);
nor U3054 (N_3054,N_2999,N_2386);
nand U3055 (N_3055,N_2907,N_2058);
nand U3056 (N_3056,N_2146,N_2864);
or U3057 (N_3057,N_2884,N_2196);
nor U3058 (N_3058,N_2376,N_2061);
or U3059 (N_3059,N_2492,N_2728);
nand U3060 (N_3060,N_2732,N_2713);
nor U3061 (N_3061,N_2438,N_2938);
nand U3062 (N_3062,N_2368,N_2932);
and U3063 (N_3063,N_2212,N_2036);
and U3064 (N_3064,N_2687,N_2436);
nor U3065 (N_3065,N_2924,N_2968);
and U3066 (N_3066,N_2390,N_2601);
nand U3067 (N_3067,N_2893,N_2743);
xnor U3068 (N_3068,N_2391,N_2296);
and U3069 (N_3069,N_2650,N_2480);
nor U3070 (N_3070,N_2116,N_2937);
xnor U3071 (N_3071,N_2998,N_2103);
nand U3072 (N_3072,N_2950,N_2784);
nor U3073 (N_3073,N_2954,N_2017);
nand U3074 (N_3074,N_2709,N_2248);
xnor U3075 (N_3075,N_2623,N_2769);
xor U3076 (N_3076,N_2959,N_2505);
nor U3077 (N_3077,N_2972,N_2651);
or U3078 (N_3078,N_2846,N_2209);
xnor U3079 (N_3079,N_2313,N_2683);
xor U3080 (N_3080,N_2371,N_2303);
or U3081 (N_3081,N_2940,N_2720);
and U3082 (N_3082,N_2403,N_2805);
nand U3083 (N_3083,N_2876,N_2222);
nand U3084 (N_3084,N_2602,N_2463);
nand U3085 (N_3085,N_2073,N_2398);
nor U3086 (N_3086,N_2158,N_2847);
xnor U3087 (N_3087,N_2757,N_2522);
or U3088 (N_3088,N_2031,N_2318);
and U3089 (N_3089,N_2002,N_2949);
and U3090 (N_3090,N_2005,N_2114);
and U3091 (N_3091,N_2345,N_2857);
nor U3092 (N_3092,N_2734,N_2226);
or U3093 (N_3093,N_2202,N_2425);
xnor U3094 (N_3094,N_2942,N_2941);
xnor U3095 (N_3095,N_2040,N_2012);
or U3096 (N_3096,N_2617,N_2304);
nor U3097 (N_3097,N_2082,N_2030);
or U3098 (N_3098,N_2738,N_2813);
and U3099 (N_3099,N_2763,N_2281);
xnor U3100 (N_3100,N_2751,N_2508);
xnor U3101 (N_3101,N_2776,N_2395);
and U3102 (N_3102,N_2903,N_2790);
xnor U3103 (N_3103,N_2016,N_2418);
and U3104 (N_3104,N_2110,N_2055);
and U3105 (N_3105,N_2833,N_2282);
or U3106 (N_3106,N_2288,N_2263);
xor U3107 (N_3107,N_2342,N_2328);
or U3108 (N_3108,N_2855,N_2465);
and U3109 (N_3109,N_2592,N_2515);
xnor U3110 (N_3110,N_2822,N_2231);
xnor U3111 (N_3111,N_2458,N_2407);
xnor U3112 (N_3112,N_2220,N_2022);
nand U3113 (N_3113,N_2748,N_2500);
nand U3114 (N_3114,N_2590,N_2934);
xor U3115 (N_3115,N_2170,N_2764);
nand U3116 (N_3116,N_2550,N_2445);
and U3117 (N_3117,N_2985,N_2203);
nor U3118 (N_3118,N_2678,N_2989);
and U3119 (N_3119,N_2213,N_2393);
nor U3120 (N_3120,N_2287,N_2184);
nand U3121 (N_3121,N_2841,N_2187);
or U3122 (N_3122,N_2039,N_2380);
nor U3123 (N_3123,N_2525,N_2581);
xor U3124 (N_3124,N_2229,N_2662);
and U3125 (N_3125,N_2691,N_2991);
nor U3126 (N_3126,N_2038,N_2446);
xnor U3127 (N_3127,N_2413,N_2659);
or U3128 (N_3128,N_2904,N_2712);
nand U3129 (N_3129,N_2330,N_2292);
nand U3130 (N_3130,N_2853,N_2042);
nor U3131 (N_3131,N_2982,N_2219);
nor U3132 (N_3132,N_2636,N_2658);
and U3133 (N_3133,N_2570,N_2247);
or U3134 (N_3134,N_2321,N_2098);
or U3135 (N_3135,N_2945,N_2337);
and U3136 (N_3136,N_2456,N_2232);
or U3137 (N_3137,N_2406,N_2746);
nor U3138 (N_3138,N_2622,N_2009);
or U3139 (N_3139,N_2533,N_2758);
or U3140 (N_3140,N_2207,N_2536);
xor U3141 (N_3141,N_2235,N_2369);
or U3142 (N_3142,N_2375,N_2530);
nand U3143 (N_3143,N_2929,N_2993);
or U3144 (N_3144,N_2239,N_2867);
nand U3145 (N_3145,N_2863,N_2965);
and U3146 (N_3146,N_2490,N_2461);
xnor U3147 (N_3147,N_2102,N_2159);
or U3148 (N_3148,N_2128,N_2820);
nor U3149 (N_3149,N_2811,N_2010);
or U3150 (N_3150,N_2766,N_2939);
nand U3151 (N_3151,N_2694,N_2374);
nand U3152 (N_3152,N_2542,N_2104);
and U3153 (N_3153,N_2051,N_2546);
or U3154 (N_3154,N_2715,N_2094);
nand U3155 (N_3155,N_2154,N_2566);
nor U3156 (N_3156,N_2412,N_2495);
or U3157 (N_3157,N_2543,N_2537);
and U3158 (N_3158,N_2344,N_2591);
or U3159 (N_3159,N_2208,N_2914);
xor U3160 (N_3160,N_2555,N_2291);
and U3161 (N_3161,N_2778,N_2365);
nor U3162 (N_3162,N_2336,N_2129);
xnor U3163 (N_3163,N_2872,N_2449);
or U3164 (N_3164,N_2933,N_2417);
xor U3165 (N_3165,N_2795,N_2453);
nor U3166 (N_3166,N_2402,N_2635);
xor U3167 (N_3167,N_2264,N_2023);
nor U3168 (N_3168,N_2249,N_2870);
xor U3169 (N_3169,N_2839,N_2830);
and U3170 (N_3170,N_2280,N_2761);
and U3171 (N_3171,N_2975,N_2526);
nor U3172 (N_3172,N_2675,N_2731);
nand U3173 (N_3173,N_2843,N_2062);
and U3174 (N_3174,N_2072,N_2752);
nand U3175 (N_3175,N_2270,N_2698);
xor U3176 (N_3176,N_2798,N_2565);
and U3177 (N_3177,N_2868,N_2771);
nand U3178 (N_3178,N_2314,N_2898);
xnor U3179 (N_3179,N_2111,N_2627);
and U3180 (N_3180,N_2567,N_2100);
xnor U3181 (N_3181,N_2832,N_2521);
or U3182 (N_3182,N_2684,N_2978);
xor U3183 (N_3183,N_2821,N_2699);
xor U3184 (N_3184,N_2124,N_2520);
or U3185 (N_3185,N_2497,N_2141);
nor U3186 (N_3186,N_2916,N_2502);
nor U3187 (N_3187,N_2071,N_2063);
nor U3188 (N_3188,N_2618,N_2849);
and U3189 (N_3189,N_2027,N_2936);
or U3190 (N_3190,N_2667,N_2271);
and U3191 (N_3191,N_2931,N_2826);
and U3192 (N_3192,N_2433,N_2243);
xnor U3193 (N_3193,N_2947,N_2472);
or U3194 (N_3194,N_2416,N_2518);
nor U3195 (N_3195,N_2092,N_2801);
nand U3196 (N_3196,N_2886,N_2324);
xnor U3197 (N_3197,N_2078,N_2167);
nand U3198 (N_3198,N_2045,N_2573);
xnor U3199 (N_3199,N_2781,N_2944);
xnor U3200 (N_3200,N_2885,N_2174);
nor U3201 (N_3201,N_2654,N_2466);
xnor U3202 (N_3202,N_2956,N_2838);
and U3203 (N_3203,N_2859,N_2619);
xnor U3204 (N_3204,N_2507,N_2528);
nor U3205 (N_3205,N_2681,N_2447);
and U3206 (N_3206,N_2861,N_2400);
and U3207 (N_3207,N_2749,N_2354);
nand U3208 (N_3208,N_2594,N_2105);
nor U3209 (N_3209,N_2775,N_2759);
nand U3210 (N_3210,N_2499,N_2952);
nand U3211 (N_3211,N_2172,N_2723);
nor U3212 (N_3212,N_2254,N_2742);
xor U3213 (N_3213,N_2341,N_2663);
or U3214 (N_3214,N_2122,N_2596);
nor U3215 (N_3215,N_2362,N_2044);
or U3216 (N_3216,N_2473,N_2133);
nand U3217 (N_3217,N_2695,N_2346);
or U3218 (N_3218,N_2419,N_2961);
and U3219 (N_3219,N_2477,N_2858);
xor U3220 (N_3220,N_2513,N_2452);
nand U3221 (N_3221,N_2367,N_2083);
xnor U3222 (N_3222,N_2901,N_2117);
xor U3223 (N_3223,N_2874,N_2994);
and U3224 (N_3224,N_2470,N_2032);
and U3225 (N_3225,N_2598,N_2227);
nand U3226 (N_3226,N_2056,N_2580);
or U3227 (N_3227,N_2988,N_2156);
nor U3228 (N_3228,N_2485,N_2647);
xor U3229 (N_3229,N_2177,N_2323);
xor U3230 (N_3230,N_2878,N_2150);
or U3231 (N_3231,N_2065,N_2143);
nand U3232 (N_3232,N_2909,N_2306);
xnor U3233 (N_3233,N_2034,N_2132);
nor U3234 (N_3234,N_2560,N_2482);
and U3235 (N_3235,N_2707,N_2268);
or U3236 (N_3236,N_2540,N_2191);
nand U3237 (N_3237,N_2225,N_2182);
and U3238 (N_3238,N_2340,N_2997);
xor U3239 (N_3239,N_2603,N_2836);
xor U3240 (N_3240,N_2812,N_2604);
or U3241 (N_3241,N_2118,N_2920);
or U3242 (N_3242,N_2708,N_2741);
or U3243 (N_3243,N_2730,N_2648);
nand U3244 (N_3244,N_2780,N_2510);
nand U3245 (N_3245,N_2892,N_2421);
and U3246 (N_3246,N_2719,N_2928);
or U3247 (N_3247,N_2350,N_2671);
and U3248 (N_3248,N_2639,N_2312);
nand U3249 (N_3249,N_2803,N_2943);
or U3250 (N_3250,N_2107,N_2028);
nor U3251 (N_3251,N_2185,N_2572);
nand U3252 (N_3252,N_2842,N_2377);
nand U3253 (N_3253,N_2149,N_2902);
nand U3254 (N_3254,N_2041,N_2523);
and U3255 (N_3255,N_2109,N_2289);
and U3256 (N_3256,N_2139,N_2511);
nor U3257 (N_3257,N_2501,N_2348);
nor U3258 (N_3258,N_2236,N_2064);
xor U3259 (N_3259,N_2087,N_2569);
or U3260 (N_3260,N_2981,N_2652);
or U3261 (N_3261,N_2962,N_2679);
nand U3262 (N_3262,N_2285,N_2689);
nor U3263 (N_3263,N_2381,N_2192);
nand U3264 (N_3264,N_2201,N_2300);
or U3265 (N_3265,N_2875,N_2926);
or U3266 (N_3266,N_2716,N_2534);
or U3267 (N_3267,N_2462,N_2599);
xnor U3268 (N_3268,N_2527,N_2744);
and U3269 (N_3269,N_2915,N_2272);
and U3270 (N_3270,N_2339,N_2649);
nor U3271 (N_3271,N_2228,N_2895);
and U3272 (N_3272,N_2774,N_2211);
and U3273 (N_3273,N_2460,N_2075);
and U3274 (N_3274,N_2283,N_2392);
nor U3275 (N_3275,N_2637,N_2646);
nor U3276 (N_3276,N_2554,N_2361);
nand U3277 (N_3277,N_2946,N_2079);
xor U3278 (N_3278,N_2316,N_2385);
xor U3279 (N_3279,N_2797,N_2399);
nor U3280 (N_3280,N_2722,N_2498);
xnor U3281 (N_3281,N_2808,N_2090);
nor U3282 (N_3282,N_2484,N_2835);
nor U3283 (N_3283,N_2702,N_2444);
or U3284 (N_3284,N_2866,N_2992);
and U3285 (N_3285,N_2953,N_2426);
xor U3286 (N_3286,N_2478,N_2277);
nor U3287 (N_3287,N_2645,N_2575);
xor U3288 (N_3288,N_2673,N_2007);
and U3289 (N_3289,N_2048,N_2725);
and U3290 (N_3290,N_2871,N_2317);
or U3291 (N_3291,N_2195,N_2628);
xnor U3292 (N_3292,N_2331,N_2134);
xor U3293 (N_3293,N_2164,N_2054);
nor U3294 (N_3294,N_2387,N_2559);
nand U3295 (N_3295,N_2397,N_2807);
nand U3296 (N_3296,N_2860,N_2273);
nor U3297 (N_3297,N_2912,N_2353);
xor U3298 (N_3298,N_2973,N_2401);
xnor U3299 (N_3299,N_2237,N_2326);
nor U3300 (N_3300,N_2606,N_2951);
nand U3301 (N_3301,N_2284,N_2597);
xnor U3302 (N_3302,N_2496,N_2454);
xnor U3303 (N_3303,N_2519,N_2524);
or U3304 (N_3304,N_2561,N_2656);
nand U3305 (N_3305,N_2137,N_2424);
nor U3306 (N_3306,N_2338,N_2148);
xor U3307 (N_3307,N_2302,N_2717);
or U3308 (N_3308,N_2762,N_2541);
or U3309 (N_3309,N_2584,N_2266);
or U3310 (N_3310,N_2782,N_2471);
xor U3311 (N_3311,N_2293,N_2918);
nand U3312 (N_3312,N_2356,N_2817);
and U3313 (N_3313,N_2557,N_2481);
or U3314 (N_3314,N_2638,N_2315);
nand U3315 (N_3315,N_2624,N_2532);
xor U3316 (N_3316,N_2373,N_2917);
nor U3317 (N_3317,N_2301,N_2214);
xor U3318 (N_3318,N_2206,N_2176);
nand U3319 (N_3319,N_2244,N_2080);
xnor U3320 (N_3320,N_2753,N_2310);
nand U3321 (N_3321,N_2718,N_2669);
and U3322 (N_3322,N_2256,N_2845);
and U3323 (N_3323,N_2183,N_2024);
and U3324 (N_3324,N_2974,N_2955);
nand U3325 (N_3325,N_2503,N_2585);
and U3326 (N_3326,N_2535,N_2305);
nand U3327 (N_3327,N_2335,N_2428);
xor U3328 (N_3328,N_2869,N_2862);
or U3329 (N_3329,N_2721,N_2754);
nor U3330 (N_3330,N_2171,N_2910);
nand U3331 (N_3331,N_2430,N_2004);
or U3332 (N_3332,N_2364,N_2091);
and U3333 (N_3333,N_2173,N_2163);
nand U3334 (N_3334,N_2611,N_2576);
nor U3335 (N_3335,N_2459,N_2011);
nor U3336 (N_3336,N_2760,N_2966);
nand U3337 (N_3337,N_2976,N_2360);
nor U3338 (N_3338,N_2262,N_2670);
xnor U3339 (N_3339,N_2145,N_2668);
xnor U3340 (N_3340,N_2818,N_2614);
nor U3341 (N_3341,N_2388,N_2265);
xor U3342 (N_3342,N_2483,N_2632);
and U3343 (N_3343,N_2726,N_2823);
or U3344 (N_3344,N_2553,N_2815);
xnor U3345 (N_3345,N_2799,N_2967);
xor U3346 (N_3346,N_2396,N_2516);
and U3347 (N_3347,N_2688,N_2577);
nor U3348 (N_3348,N_2883,N_2286);
nor U3349 (N_3349,N_2383,N_2674);
xor U3350 (N_3350,N_2986,N_2298);
xnor U3351 (N_3351,N_2035,N_2439);
nor U3352 (N_3352,N_2165,N_2188);
nor U3353 (N_3353,N_2630,N_2205);
or U3354 (N_3354,N_2506,N_2408);
nand U3355 (N_3355,N_2889,N_2476);
and U3356 (N_3356,N_2161,N_2352);
nor U3357 (N_3357,N_2238,N_2747);
and U3358 (N_3358,N_2234,N_2442);
or U3359 (N_3359,N_2299,N_2144);
and U3360 (N_3360,N_2370,N_2245);
xor U3361 (N_3361,N_2077,N_2468);
nand U3362 (N_3362,N_2547,N_2015);
nand U3363 (N_3363,N_2809,N_2963);
and U3364 (N_3364,N_2179,N_2001);
nand U3365 (N_3365,N_2274,N_2355);
xnor U3366 (N_3366,N_2127,N_2672);
nand U3367 (N_3367,N_2578,N_2157);
nand U3368 (N_3368,N_2194,N_2160);
or U3369 (N_3369,N_2437,N_2115);
or U3370 (N_3370,N_2070,N_2958);
xnor U3371 (N_3371,N_2119,N_2120);
xnor U3372 (N_3372,N_2588,N_2905);
nor U3373 (N_3373,N_2140,N_2382);
nand U3374 (N_3374,N_2372,N_2198);
and U3375 (N_3375,N_2625,N_2253);
or U3376 (N_3376,N_2765,N_2925);
or U3377 (N_3377,N_2586,N_2366);
xor U3378 (N_3378,N_2930,N_2216);
nor U3379 (N_3379,N_2692,N_2677);
or U3380 (N_3380,N_2384,N_2665);
and U3381 (N_3381,N_2431,N_2739);
xnor U3382 (N_3382,N_2475,N_2634);
or U3383 (N_3383,N_2562,N_2469);
or U3384 (N_3384,N_2311,N_2837);
nor U3385 (N_3385,N_2514,N_2789);
and U3386 (N_3386,N_2794,N_2504);
nand U3387 (N_3387,N_2703,N_2531);
nor U3388 (N_3388,N_2896,N_2297);
or U3389 (N_3389,N_2267,N_2900);
and U3390 (N_3390,N_2777,N_2509);
and U3391 (N_3391,N_2615,N_2359);
xor U3392 (N_3392,N_2911,N_2013);
and U3393 (N_3393,N_2923,N_2043);
nand U3394 (N_3394,N_2996,N_2676);
xnor U3395 (N_3395,N_2394,N_2791);
and U3396 (N_3396,N_2880,N_2705);
xnor U3397 (N_3397,N_2112,N_2215);
xnor U3398 (N_3398,N_2922,N_2620);
xor U3399 (N_3399,N_2414,N_2066);
or U3400 (N_3400,N_2162,N_2682);
xor U3401 (N_3401,N_2970,N_2053);
nand U3402 (N_3402,N_2621,N_2076);
or U3403 (N_3403,N_2792,N_2450);
nand U3404 (N_3404,N_2152,N_2666);
nand U3405 (N_3405,N_2435,N_2242);
and U3406 (N_3406,N_2852,N_2729);
or U3407 (N_3407,N_2644,N_2711);
xnor U3408 (N_3408,N_2464,N_2250);
xnor U3409 (N_3409,N_2033,N_2680);
nand U3410 (N_3410,N_2168,N_2693);
nand U3411 (N_3411,N_2583,N_2479);
nor U3412 (N_3412,N_2019,N_2854);
xor U3413 (N_3413,N_2788,N_2850);
or U3414 (N_3414,N_2517,N_2260);
nor U3415 (N_3415,N_2057,N_2008);
or U3416 (N_3416,N_2643,N_2877);
xor U3417 (N_3417,N_2147,N_2897);
nor U3418 (N_3418,N_2059,N_2246);
or U3419 (N_3419,N_2276,N_2275);
nand U3420 (N_3420,N_2448,N_2879);
xnor U3421 (N_3421,N_2564,N_2607);
xnor U3422 (N_3422,N_2980,N_2856);
nand U3423 (N_3423,N_2785,N_2494);
or U3424 (N_3424,N_2714,N_2204);
nor U3425 (N_3425,N_2142,N_2848);
xor U3426 (N_3426,N_2593,N_2347);
nor U3427 (N_3427,N_2474,N_2701);
and U3428 (N_3428,N_2363,N_2810);
nand U3429 (N_3429,N_2983,N_2101);
nand U3430 (N_3430,N_2060,N_2014);
nor U3431 (N_3431,N_2434,N_2512);
nand U3432 (N_3432,N_2551,N_2081);
xnor U3433 (N_3433,N_2800,N_2825);
xnor U3434 (N_3434,N_2389,N_2491);
xnor U3435 (N_3435,N_2175,N_2224);
nor U3436 (N_3436,N_2322,N_2629);
or U3437 (N_3437,N_2787,N_2052);
or U3438 (N_3438,N_2831,N_2130);
nand U3439 (N_3439,N_2768,N_2332);
nor U3440 (N_3440,N_2021,N_2046);
xnor U3441 (N_3441,N_2919,N_2489);
and U3442 (N_3442,N_2029,N_2294);
and U3443 (N_3443,N_2613,N_2887);
or U3444 (N_3444,N_2840,N_2217);
xor U3445 (N_3445,N_2828,N_2612);
nand U3446 (N_3446,N_2343,N_2558);
nand U3447 (N_3447,N_2153,N_2197);
or U3448 (N_3448,N_2844,N_2582);
xnor U3449 (N_3449,N_2290,N_2908);
or U3450 (N_3450,N_2661,N_2616);
xnor U3451 (N_3451,N_2257,N_2166);
xnor U3452 (N_3452,N_2740,N_2405);
nor U3453 (N_3453,N_2633,N_2404);
nor U3454 (N_3454,N_2589,N_2969);
or U3455 (N_3455,N_2995,N_2240);
and U3456 (N_3456,N_2126,N_2685);
nor U3457 (N_3457,N_2258,N_2084);
nand U3458 (N_3458,N_2186,N_2088);
or U3459 (N_3459,N_2295,N_2824);
or U3460 (N_3460,N_2074,N_2193);
or U3461 (N_3461,N_2710,N_2000);
or U3462 (N_3462,N_2487,N_2608);
nand U3463 (N_3463,N_2804,N_2432);
or U3464 (N_3464,N_2979,N_2935);
and U3465 (N_3465,N_2068,N_2488);
xnor U3466 (N_3466,N_2047,N_2357);
xnor U3467 (N_3467,N_2443,N_2178);
and U3468 (N_3468,N_2415,N_2309);
and U3469 (N_3469,N_2096,N_2086);
nor U3470 (N_3470,N_2131,N_2218);
xor U3471 (N_3471,N_2233,N_2796);
xnor U3472 (N_3472,N_2755,N_2626);
xnor U3473 (N_3473,N_2890,N_2358);
or U3474 (N_3474,N_2737,N_2660);
nor U3475 (N_3475,N_2690,N_2067);
nor U3476 (N_3476,N_2097,N_2881);
nand U3477 (N_3477,N_2411,N_2135);
nor U3478 (N_3478,N_2960,N_2093);
nor U3479 (N_3479,N_2579,N_2819);
nor U3480 (N_3480,N_2529,N_2587);
xnor U3481 (N_3481,N_2806,N_2779);
nand U3482 (N_3482,N_2409,N_2770);
and U3483 (N_3483,N_2750,N_2099);
nor U3484 (N_3484,N_2556,N_2441);
xnor U3485 (N_3485,N_2990,N_2571);
xor U3486 (N_3486,N_2451,N_2727);
or U3487 (N_3487,N_2704,N_2610);
and U3488 (N_3488,N_2735,N_2829);
nand U3489 (N_3489,N_2653,N_2563);
and U3490 (N_3490,N_2422,N_2657);
or U3491 (N_3491,N_2169,N_2095);
nor U3492 (N_3492,N_2486,N_2786);
nand U3493 (N_3493,N_2894,N_2085);
nor U3494 (N_3494,N_2223,N_2190);
or U3495 (N_3495,N_2429,N_2697);
or U3496 (N_3496,N_2269,N_2006);
and U3497 (N_3497,N_2545,N_2733);
nor U3498 (N_3498,N_2568,N_2827);
or U3499 (N_3499,N_2745,N_2865);
nand U3500 (N_3500,N_2436,N_2549);
or U3501 (N_3501,N_2842,N_2429);
xnor U3502 (N_3502,N_2346,N_2149);
and U3503 (N_3503,N_2874,N_2547);
nand U3504 (N_3504,N_2737,N_2911);
and U3505 (N_3505,N_2872,N_2268);
or U3506 (N_3506,N_2861,N_2930);
nand U3507 (N_3507,N_2164,N_2399);
xor U3508 (N_3508,N_2975,N_2905);
and U3509 (N_3509,N_2474,N_2999);
xnor U3510 (N_3510,N_2663,N_2704);
xnor U3511 (N_3511,N_2434,N_2545);
and U3512 (N_3512,N_2071,N_2487);
and U3513 (N_3513,N_2732,N_2149);
nand U3514 (N_3514,N_2187,N_2085);
nor U3515 (N_3515,N_2902,N_2203);
xnor U3516 (N_3516,N_2489,N_2701);
xor U3517 (N_3517,N_2625,N_2544);
nand U3518 (N_3518,N_2870,N_2014);
nor U3519 (N_3519,N_2672,N_2812);
xnor U3520 (N_3520,N_2436,N_2817);
or U3521 (N_3521,N_2295,N_2953);
or U3522 (N_3522,N_2804,N_2338);
nor U3523 (N_3523,N_2178,N_2342);
nand U3524 (N_3524,N_2170,N_2519);
nor U3525 (N_3525,N_2211,N_2314);
nor U3526 (N_3526,N_2433,N_2067);
and U3527 (N_3527,N_2740,N_2367);
xor U3528 (N_3528,N_2720,N_2353);
and U3529 (N_3529,N_2858,N_2276);
nor U3530 (N_3530,N_2859,N_2627);
xnor U3531 (N_3531,N_2844,N_2996);
nor U3532 (N_3532,N_2529,N_2912);
nor U3533 (N_3533,N_2949,N_2503);
and U3534 (N_3534,N_2797,N_2794);
xor U3535 (N_3535,N_2039,N_2637);
nand U3536 (N_3536,N_2554,N_2857);
xnor U3537 (N_3537,N_2285,N_2962);
xor U3538 (N_3538,N_2175,N_2148);
nor U3539 (N_3539,N_2418,N_2865);
nand U3540 (N_3540,N_2684,N_2137);
nand U3541 (N_3541,N_2842,N_2780);
nand U3542 (N_3542,N_2465,N_2033);
and U3543 (N_3543,N_2395,N_2934);
nor U3544 (N_3544,N_2953,N_2738);
nand U3545 (N_3545,N_2759,N_2651);
or U3546 (N_3546,N_2596,N_2111);
nor U3547 (N_3547,N_2289,N_2778);
nor U3548 (N_3548,N_2676,N_2609);
or U3549 (N_3549,N_2779,N_2257);
xor U3550 (N_3550,N_2646,N_2517);
nor U3551 (N_3551,N_2302,N_2364);
nand U3552 (N_3552,N_2792,N_2204);
and U3553 (N_3553,N_2510,N_2280);
nand U3554 (N_3554,N_2060,N_2595);
xor U3555 (N_3555,N_2291,N_2199);
nand U3556 (N_3556,N_2874,N_2773);
or U3557 (N_3557,N_2119,N_2334);
nand U3558 (N_3558,N_2966,N_2016);
nand U3559 (N_3559,N_2473,N_2898);
nand U3560 (N_3560,N_2281,N_2310);
and U3561 (N_3561,N_2144,N_2803);
nand U3562 (N_3562,N_2361,N_2235);
nand U3563 (N_3563,N_2694,N_2964);
nand U3564 (N_3564,N_2469,N_2660);
xor U3565 (N_3565,N_2465,N_2153);
nand U3566 (N_3566,N_2461,N_2431);
and U3567 (N_3567,N_2639,N_2908);
xor U3568 (N_3568,N_2601,N_2854);
xor U3569 (N_3569,N_2821,N_2495);
and U3570 (N_3570,N_2207,N_2328);
xnor U3571 (N_3571,N_2562,N_2831);
or U3572 (N_3572,N_2780,N_2183);
nand U3573 (N_3573,N_2142,N_2189);
or U3574 (N_3574,N_2575,N_2378);
and U3575 (N_3575,N_2830,N_2605);
nor U3576 (N_3576,N_2181,N_2648);
xor U3577 (N_3577,N_2234,N_2122);
xor U3578 (N_3578,N_2802,N_2845);
xor U3579 (N_3579,N_2335,N_2643);
nor U3580 (N_3580,N_2843,N_2135);
nor U3581 (N_3581,N_2173,N_2194);
and U3582 (N_3582,N_2101,N_2619);
xnor U3583 (N_3583,N_2856,N_2277);
xnor U3584 (N_3584,N_2487,N_2325);
and U3585 (N_3585,N_2958,N_2567);
or U3586 (N_3586,N_2363,N_2578);
nor U3587 (N_3587,N_2170,N_2180);
or U3588 (N_3588,N_2104,N_2152);
xnor U3589 (N_3589,N_2912,N_2857);
xor U3590 (N_3590,N_2165,N_2863);
nor U3591 (N_3591,N_2840,N_2854);
nand U3592 (N_3592,N_2332,N_2640);
xnor U3593 (N_3593,N_2734,N_2384);
or U3594 (N_3594,N_2934,N_2822);
and U3595 (N_3595,N_2305,N_2832);
nor U3596 (N_3596,N_2430,N_2686);
xor U3597 (N_3597,N_2816,N_2937);
nor U3598 (N_3598,N_2786,N_2423);
nand U3599 (N_3599,N_2542,N_2599);
xnor U3600 (N_3600,N_2272,N_2800);
and U3601 (N_3601,N_2260,N_2312);
and U3602 (N_3602,N_2439,N_2773);
and U3603 (N_3603,N_2095,N_2774);
nor U3604 (N_3604,N_2163,N_2117);
xnor U3605 (N_3605,N_2102,N_2324);
and U3606 (N_3606,N_2816,N_2100);
or U3607 (N_3607,N_2292,N_2558);
nor U3608 (N_3608,N_2370,N_2604);
or U3609 (N_3609,N_2981,N_2454);
nor U3610 (N_3610,N_2473,N_2681);
nand U3611 (N_3611,N_2055,N_2300);
nand U3612 (N_3612,N_2223,N_2780);
and U3613 (N_3613,N_2366,N_2625);
or U3614 (N_3614,N_2356,N_2328);
and U3615 (N_3615,N_2390,N_2232);
or U3616 (N_3616,N_2536,N_2450);
nor U3617 (N_3617,N_2137,N_2640);
nor U3618 (N_3618,N_2488,N_2976);
or U3619 (N_3619,N_2998,N_2847);
nand U3620 (N_3620,N_2116,N_2017);
nand U3621 (N_3621,N_2838,N_2675);
or U3622 (N_3622,N_2441,N_2580);
or U3623 (N_3623,N_2340,N_2564);
or U3624 (N_3624,N_2712,N_2875);
xnor U3625 (N_3625,N_2206,N_2700);
nor U3626 (N_3626,N_2297,N_2541);
nand U3627 (N_3627,N_2973,N_2084);
and U3628 (N_3628,N_2539,N_2493);
and U3629 (N_3629,N_2304,N_2234);
xor U3630 (N_3630,N_2818,N_2459);
or U3631 (N_3631,N_2852,N_2452);
and U3632 (N_3632,N_2857,N_2803);
and U3633 (N_3633,N_2815,N_2979);
and U3634 (N_3634,N_2542,N_2879);
nor U3635 (N_3635,N_2123,N_2622);
nand U3636 (N_3636,N_2195,N_2641);
xor U3637 (N_3637,N_2335,N_2888);
or U3638 (N_3638,N_2711,N_2575);
nor U3639 (N_3639,N_2948,N_2909);
nand U3640 (N_3640,N_2537,N_2370);
or U3641 (N_3641,N_2864,N_2603);
xor U3642 (N_3642,N_2238,N_2736);
nand U3643 (N_3643,N_2651,N_2149);
or U3644 (N_3644,N_2748,N_2392);
nand U3645 (N_3645,N_2549,N_2078);
nand U3646 (N_3646,N_2095,N_2319);
xnor U3647 (N_3647,N_2609,N_2353);
and U3648 (N_3648,N_2202,N_2831);
nand U3649 (N_3649,N_2038,N_2732);
xnor U3650 (N_3650,N_2111,N_2960);
or U3651 (N_3651,N_2906,N_2883);
nor U3652 (N_3652,N_2210,N_2404);
xor U3653 (N_3653,N_2956,N_2028);
and U3654 (N_3654,N_2576,N_2183);
and U3655 (N_3655,N_2531,N_2825);
nor U3656 (N_3656,N_2025,N_2603);
or U3657 (N_3657,N_2904,N_2009);
nand U3658 (N_3658,N_2742,N_2844);
nand U3659 (N_3659,N_2983,N_2427);
or U3660 (N_3660,N_2561,N_2191);
xor U3661 (N_3661,N_2791,N_2287);
nor U3662 (N_3662,N_2046,N_2978);
nor U3663 (N_3663,N_2103,N_2255);
and U3664 (N_3664,N_2416,N_2987);
nor U3665 (N_3665,N_2537,N_2451);
and U3666 (N_3666,N_2051,N_2239);
or U3667 (N_3667,N_2892,N_2595);
or U3668 (N_3668,N_2942,N_2859);
or U3669 (N_3669,N_2053,N_2847);
xor U3670 (N_3670,N_2034,N_2463);
nor U3671 (N_3671,N_2244,N_2735);
xnor U3672 (N_3672,N_2435,N_2743);
or U3673 (N_3673,N_2916,N_2236);
and U3674 (N_3674,N_2665,N_2580);
and U3675 (N_3675,N_2370,N_2192);
or U3676 (N_3676,N_2363,N_2451);
nand U3677 (N_3677,N_2429,N_2468);
xor U3678 (N_3678,N_2219,N_2683);
and U3679 (N_3679,N_2554,N_2381);
nand U3680 (N_3680,N_2722,N_2902);
and U3681 (N_3681,N_2849,N_2632);
and U3682 (N_3682,N_2242,N_2427);
and U3683 (N_3683,N_2635,N_2128);
and U3684 (N_3684,N_2376,N_2901);
and U3685 (N_3685,N_2397,N_2301);
nor U3686 (N_3686,N_2374,N_2471);
and U3687 (N_3687,N_2145,N_2248);
xnor U3688 (N_3688,N_2126,N_2276);
or U3689 (N_3689,N_2586,N_2482);
nand U3690 (N_3690,N_2654,N_2952);
xor U3691 (N_3691,N_2250,N_2100);
nand U3692 (N_3692,N_2093,N_2974);
nand U3693 (N_3693,N_2316,N_2713);
xor U3694 (N_3694,N_2263,N_2086);
and U3695 (N_3695,N_2777,N_2236);
xor U3696 (N_3696,N_2565,N_2248);
xor U3697 (N_3697,N_2007,N_2261);
or U3698 (N_3698,N_2885,N_2554);
and U3699 (N_3699,N_2787,N_2776);
xor U3700 (N_3700,N_2295,N_2795);
or U3701 (N_3701,N_2382,N_2249);
xor U3702 (N_3702,N_2874,N_2410);
or U3703 (N_3703,N_2449,N_2417);
nor U3704 (N_3704,N_2134,N_2556);
nand U3705 (N_3705,N_2782,N_2282);
xnor U3706 (N_3706,N_2162,N_2898);
nand U3707 (N_3707,N_2185,N_2672);
or U3708 (N_3708,N_2891,N_2836);
and U3709 (N_3709,N_2600,N_2624);
nand U3710 (N_3710,N_2953,N_2247);
or U3711 (N_3711,N_2136,N_2126);
and U3712 (N_3712,N_2088,N_2705);
or U3713 (N_3713,N_2775,N_2255);
and U3714 (N_3714,N_2948,N_2453);
xnor U3715 (N_3715,N_2762,N_2530);
nor U3716 (N_3716,N_2052,N_2184);
xnor U3717 (N_3717,N_2144,N_2180);
nor U3718 (N_3718,N_2528,N_2400);
and U3719 (N_3719,N_2017,N_2695);
xor U3720 (N_3720,N_2334,N_2575);
xnor U3721 (N_3721,N_2535,N_2234);
nor U3722 (N_3722,N_2785,N_2742);
nor U3723 (N_3723,N_2336,N_2890);
and U3724 (N_3724,N_2020,N_2851);
nor U3725 (N_3725,N_2236,N_2218);
or U3726 (N_3726,N_2137,N_2273);
nand U3727 (N_3727,N_2801,N_2363);
or U3728 (N_3728,N_2852,N_2053);
nand U3729 (N_3729,N_2981,N_2070);
or U3730 (N_3730,N_2913,N_2521);
nor U3731 (N_3731,N_2540,N_2491);
nor U3732 (N_3732,N_2972,N_2817);
xor U3733 (N_3733,N_2360,N_2411);
nor U3734 (N_3734,N_2196,N_2847);
nor U3735 (N_3735,N_2551,N_2280);
xnor U3736 (N_3736,N_2251,N_2298);
or U3737 (N_3737,N_2562,N_2607);
or U3738 (N_3738,N_2254,N_2046);
xor U3739 (N_3739,N_2381,N_2497);
xor U3740 (N_3740,N_2209,N_2500);
and U3741 (N_3741,N_2213,N_2426);
xor U3742 (N_3742,N_2397,N_2167);
xor U3743 (N_3743,N_2100,N_2981);
nand U3744 (N_3744,N_2028,N_2637);
nand U3745 (N_3745,N_2434,N_2997);
or U3746 (N_3746,N_2475,N_2062);
xor U3747 (N_3747,N_2796,N_2988);
or U3748 (N_3748,N_2844,N_2292);
nor U3749 (N_3749,N_2086,N_2999);
nand U3750 (N_3750,N_2104,N_2226);
nor U3751 (N_3751,N_2480,N_2019);
nor U3752 (N_3752,N_2246,N_2891);
nor U3753 (N_3753,N_2977,N_2126);
nor U3754 (N_3754,N_2427,N_2574);
and U3755 (N_3755,N_2075,N_2663);
xor U3756 (N_3756,N_2486,N_2959);
xnor U3757 (N_3757,N_2570,N_2404);
and U3758 (N_3758,N_2805,N_2433);
nand U3759 (N_3759,N_2164,N_2439);
xor U3760 (N_3760,N_2141,N_2512);
and U3761 (N_3761,N_2874,N_2080);
xnor U3762 (N_3762,N_2774,N_2890);
and U3763 (N_3763,N_2243,N_2392);
nand U3764 (N_3764,N_2673,N_2488);
xor U3765 (N_3765,N_2745,N_2123);
nand U3766 (N_3766,N_2266,N_2511);
xnor U3767 (N_3767,N_2863,N_2458);
nor U3768 (N_3768,N_2417,N_2297);
and U3769 (N_3769,N_2711,N_2336);
and U3770 (N_3770,N_2246,N_2822);
nand U3771 (N_3771,N_2152,N_2665);
xnor U3772 (N_3772,N_2837,N_2010);
nor U3773 (N_3773,N_2894,N_2333);
nor U3774 (N_3774,N_2054,N_2832);
xor U3775 (N_3775,N_2158,N_2932);
or U3776 (N_3776,N_2272,N_2648);
and U3777 (N_3777,N_2904,N_2225);
nor U3778 (N_3778,N_2385,N_2899);
or U3779 (N_3779,N_2246,N_2256);
nor U3780 (N_3780,N_2348,N_2182);
nor U3781 (N_3781,N_2190,N_2784);
nor U3782 (N_3782,N_2516,N_2648);
nand U3783 (N_3783,N_2507,N_2419);
and U3784 (N_3784,N_2016,N_2337);
and U3785 (N_3785,N_2025,N_2006);
nand U3786 (N_3786,N_2828,N_2560);
nand U3787 (N_3787,N_2272,N_2191);
or U3788 (N_3788,N_2555,N_2200);
and U3789 (N_3789,N_2195,N_2309);
nor U3790 (N_3790,N_2941,N_2594);
xnor U3791 (N_3791,N_2089,N_2638);
xnor U3792 (N_3792,N_2196,N_2198);
xnor U3793 (N_3793,N_2661,N_2830);
and U3794 (N_3794,N_2169,N_2748);
and U3795 (N_3795,N_2558,N_2414);
or U3796 (N_3796,N_2007,N_2128);
xor U3797 (N_3797,N_2978,N_2900);
and U3798 (N_3798,N_2621,N_2974);
nand U3799 (N_3799,N_2338,N_2418);
nor U3800 (N_3800,N_2442,N_2191);
and U3801 (N_3801,N_2105,N_2034);
or U3802 (N_3802,N_2514,N_2553);
nor U3803 (N_3803,N_2408,N_2125);
nor U3804 (N_3804,N_2482,N_2678);
or U3805 (N_3805,N_2909,N_2430);
xor U3806 (N_3806,N_2930,N_2584);
xor U3807 (N_3807,N_2822,N_2540);
xnor U3808 (N_3808,N_2151,N_2114);
nor U3809 (N_3809,N_2515,N_2248);
nand U3810 (N_3810,N_2846,N_2219);
nand U3811 (N_3811,N_2490,N_2622);
or U3812 (N_3812,N_2132,N_2419);
or U3813 (N_3813,N_2614,N_2138);
nor U3814 (N_3814,N_2129,N_2064);
xnor U3815 (N_3815,N_2285,N_2309);
or U3816 (N_3816,N_2204,N_2104);
xnor U3817 (N_3817,N_2991,N_2449);
xor U3818 (N_3818,N_2897,N_2159);
nand U3819 (N_3819,N_2782,N_2777);
and U3820 (N_3820,N_2570,N_2374);
and U3821 (N_3821,N_2200,N_2772);
nand U3822 (N_3822,N_2562,N_2347);
or U3823 (N_3823,N_2912,N_2491);
nand U3824 (N_3824,N_2930,N_2307);
xor U3825 (N_3825,N_2760,N_2820);
xor U3826 (N_3826,N_2069,N_2127);
or U3827 (N_3827,N_2540,N_2381);
xnor U3828 (N_3828,N_2220,N_2683);
nand U3829 (N_3829,N_2949,N_2446);
or U3830 (N_3830,N_2075,N_2893);
and U3831 (N_3831,N_2253,N_2969);
or U3832 (N_3832,N_2083,N_2412);
nor U3833 (N_3833,N_2567,N_2841);
nand U3834 (N_3834,N_2408,N_2415);
xor U3835 (N_3835,N_2294,N_2726);
and U3836 (N_3836,N_2138,N_2608);
nor U3837 (N_3837,N_2676,N_2650);
nand U3838 (N_3838,N_2293,N_2957);
and U3839 (N_3839,N_2604,N_2014);
xnor U3840 (N_3840,N_2901,N_2874);
or U3841 (N_3841,N_2977,N_2195);
nand U3842 (N_3842,N_2072,N_2406);
nand U3843 (N_3843,N_2170,N_2446);
nand U3844 (N_3844,N_2675,N_2049);
or U3845 (N_3845,N_2134,N_2152);
or U3846 (N_3846,N_2678,N_2349);
and U3847 (N_3847,N_2002,N_2459);
or U3848 (N_3848,N_2230,N_2389);
nor U3849 (N_3849,N_2133,N_2477);
and U3850 (N_3850,N_2427,N_2048);
nand U3851 (N_3851,N_2144,N_2311);
xnor U3852 (N_3852,N_2586,N_2079);
and U3853 (N_3853,N_2889,N_2613);
or U3854 (N_3854,N_2706,N_2765);
nand U3855 (N_3855,N_2992,N_2208);
xor U3856 (N_3856,N_2818,N_2776);
and U3857 (N_3857,N_2424,N_2953);
nor U3858 (N_3858,N_2544,N_2735);
and U3859 (N_3859,N_2231,N_2996);
nor U3860 (N_3860,N_2109,N_2421);
nor U3861 (N_3861,N_2679,N_2536);
nand U3862 (N_3862,N_2506,N_2681);
or U3863 (N_3863,N_2899,N_2248);
xnor U3864 (N_3864,N_2100,N_2918);
or U3865 (N_3865,N_2456,N_2870);
and U3866 (N_3866,N_2729,N_2878);
nand U3867 (N_3867,N_2978,N_2734);
nor U3868 (N_3868,N_2738,N_2185);
or U3869 (N_3869,N_2961,N_2716);
nand U3870 (N_3870,N_2180,N_2922);
nand U3871 (N_3871,N_2406,N_2902);
or U3872 (N_3872,N_2897,N_2298);
and U3873 (N_3873,N_2204,N_2923);
xor U3874 (N_3874,N_2350,N_2752);
or U3875 (N_3875,N_2699,N_2764);
xor U3876 (N_3876,N_2645,N_2553);
xnor U3877 (N_3877,N_2660,N_2859);
xor U3878 (N_3878,N_2377,N_2710);
nor U3879 (N_3879,N_2625,N_2047);
or U3880 (N_3880,N_2952,N_2324);
xnor U3881 (N_3881,N_2645,N_2305);
or U3882 (N_3882,N_2012,N_2794);
xor U3883 (N_3883,N_2013,N_2217);
nor U3884 (N_3884,N_2906,N_2603);
and U3885 (N_3885,N_2649,N_2720);
or U3886 (N_3886,N_2691,N_2411);
nand U3887 (N_3887,N_2712,N_2164);
nand U3888 (N_3888,N_2616,N_2969);
xor U3889 (N_3889,N_2727,N_2303);
and U3890 (N_3890,N_2170,N_2595);
and U3891 (N_3891,N_2516,N_2650);
or U3892 (N_3892,N_2906,N_2934);
nand U3893 (N_3893,N_2973,N_2722);
or U3894 (N_3894,N_2006,N_2019);
or U3895 (N_3895,N_2239,N_2611);
or U3896 (N_3896,N_2831,N_2487);
nand U3897 (N_3897,N_2713,N_2562);
xnor U3898 (N_3898,N_2578,N_2262);
and U3899 (N_3899,N_2145,N_2933);
nand U3900 (N_3900,N_2099,N_2088);
or U3901 (N_3901,N_2230,N_2184);
xor U3902 (N_3902,N_2854,N_2441);
or U3903 (N_3903,N_2692,N_2238);
xnor U3904 (N_3904,N_2905,N_2395);
xor U3905 (N_3905,N_2218,N_2576);
nand U3906 (N_3906,N_2900,N_2494);
and U3907 (N_3907,N_2678,N_2589);
nand U3908 (N_3908,N_2781,N_2704);
and U3909 (N_3909,N_2755,N_2351);
or U3910 (N_3910,N_2742,N_2874);
xnor U3911 (N_3911,N_2757,N_2361);
xnor U3912 (N_3912,N_2386,N_2079);
nor U3913 (N_3913,N_2587,N_2721);
or U3914 (N_3914,N_2068,N_2385);
xnor U3915 (N_3915,N_2482,N_2275);
nor U3916 (N_3916,N_2380,N_2640);
xor U3917 (N_3917,N_2508,N_2485);
or U3918 (N_3918,N_2623,N_2509);
nor U3919 (N_3919,N_2063,N_2028);
nor U3920 (N_3920,N_2627,N_2551);
nand U3921 (N_3921,N_2977,N_2382);
nand U3922 (N_3922,N_2565,N_2029);
and U3923 (N_3923,N_2022,N_2471);
and U3924 (N_3924,N_2802,N_2357);
xnor U3925 (N_3925,N_2788,N_2064);
nand U3926 (N_3926,N_2101,N_2757);
and U3927 (N_3927,N_2912,N_2446);
nand U3928 (N_3928,N_2811,N_2282);
nor U3929 (N_3929,N_2595,N_2447);
xor U3930 (N_3930,N_2788,N_2682);
nand U3931 (N_3931,N_2590,N_2765);
xor U3932 (N_3932,N_2835,N_2400);
nand U3933 (N_3933,N_2713,N_2983);
xnor U3934 (N_3934,N_2374,N_2338);
or U3935 (N_3935,N_2308,N_2056);
or U3936 (N_3936,N_2697,N_2104);
nand U3937 (N_3937,N_2961,N_2789);
or U3938 (N_3938,N_2074,N_2241);
nand U3939 (N_3939,N_2713,N_2925);
and U3940 (N_3940,N_2682,N_2327);
nand U3941 (N_3941,N_2089,N_2840);
and U3942 (N_3942,N_2663,N_2771);
and U3943 (N_3943,N_2873,N_2146);
and U3944 (N_3944,N_2367,N_2777);
or U3945 (N_3945,N_2663,N_2629);
xor U3946 (N_3946,N_2898,N_2108);
xnor U3947 (N_3947,N_2051,N_2499);
and U3948 (N_3948,N_2886,N_2401);
nand U3949 (N_3949,N_2450,N_2378);
nor U3950 (N_3950,N_2282,N_2466);
or U3951 (N_3951,N_2767,N_2014);
xnor U3952 (N_3952,N_2560,N_2917);
or U3953 (N_3953,N_2239,N_2707);
nor U3954 (N_3954,N_2935,N_2371);
and U3955 (N_3955,N_2880,N_2991);
nand U3956 (N_3956,N_2211,N_2768);
xnor U3957 (N_3957,N_2451,N_2686);
xor U3958 (N_3958,N_2329,N_2480);
or U3959 (N_3959,N_2946,N_2459);
and U3960 (N_3960,N_2462,N_2987);
xor U3961 (N_3961,N_2030,N_2383);
xnor U3962 (N_3962,N_2561,N_2460);
and U3963 (N_3963,N_2265,N_2295);
and U3964 (N_3964,N_2238,N_2947);
and U3965 (N_3965,N_2570,N_2597);
and U3966 (N_3966,N_2957,N_2392);
nand U3967 (N_3967,N_2073,N_2981);
xnor U3968 (N_3968,N_2619,N_2156);
nor U3969 (N_3969,N_2260,N_2602);
and U3970 (N_3970,N_2381,N_2203);
nor U3971 (N_3971,N_2761,N_2438);
and U3972 (N_3972,N_2351,N_2413);
or U3973 (N_3973,N_2977,N_2292);
and U3974 (N_3974,N_2711,N_2274);
and U3975 (N_3975,N_2684,N_2821);
nand U3976 (N_3976,N_2607,N_2389);
nand U3977 (N_3977,N_2156,N_2984);
and U3978 (N_3978,N_2387,N_2037);
nand U3979 (N_3979,N_2659,N_2573);
nor U3980 (N_3980,N_2996,N_2847);
and U3981 (N_3981,N_2520,N_2207);
and U3982 (N_3982,N_2056,N_2099);
or U3983 (N_3983,N_2585,N_2564);
xor U3984 (N_3984,N_2632,N_2062);
or U3985 (N_3985,N_2628,N_2476);
and U3986 (N_3986,N_2525,N_2793);
nor U3987 (N_3987,N_2718,N_2203);
or U3988 (N_3988,N_2394,N_2049);
nor U3989 (N_3989,N_2450,N_2322);
nand U3990 (N_3990,N_2474,N_2881);
xor U3991 (N_3991,N_2710,N_2720);
nor U3992 (N_3992,N_2603,N_2047);
xor U3993 (N_3993,N_2357,N_2298);
and U3994 (N_3994,N_2191,N_2849);
nand U3995 (N_3995,N_2846,N_2591);
xor U3996 (N_3996,N_2563,N_2855);
or U3997 (N_3997,N_2150,N_2407);
xnor U3998 (N_3998,N_2881,N_2231);
nand U3999 (N_3999,N_2210,N_2689);
nor U4000 (N_4000,N_3673,N_3311);
or U4001 (N_4001,N_3502,N_3517);
xor U4002 (N_4002,N_3855,N_3227);
nand U4003 (N_4003,N_3841,N_3246);
and U4004 (N_4004,N_3678,N_3591);
or U4005 (N_4005,N_3479,N_3388);
nand U4006 (N_4006,N_3395,N_3335);
and U4007 (N_4007,N_3228,N_3033);
and U4008 (N_4008,N_3083,N_3936);
or U4009 (N_4009,N_3533,N_3566);
nand U4010 (N_4010,N_3062,N_3880);
xor U4011 (N_4011,N_3961,N_3409);
and U4012 (N_4012,N_3509,N_3790);
nor U4013 (N_4013,N_3672,N_3028);
xor U4014 (N_4014,N_3941,N_3477);
nand U4015 (N_4015,N_3027,N_3314);
and U4016 (N_4016,N_3039,N_3490);
and U4017 (N_4017,N_3011,N_3698);
and U4018 (N_4018,N_3838,N_3573);
or U4019 (N_4019,N_3156,N_3644);
and U4020 (N_4020,N_3846,N_3580);
xnor U4021 (N_4021,N_3243,N_3373);
nor U4022 (N_4022,N_3784,N_3519);
and U4023 (N_4023,N_3697,N_3840);
xnor U4024 (N_4024,N_3331,N_3076);
nor U4025 (N_4025,N_3912,N_3952);
nor U4026 (N_4026,N_3976,N_3347);
and U4027 (N_4027,N_3878,N_3499);
xnor U4028 (N_4028,N_3748,N_3422);
and U4029 (N_4029,N_3148,N_3398);
xor U4030 (N_4030,N_3590,N_3470);
nand U4031 (N_4031,N_3787,N_3460);
or U4032 (N_4032,N_3351,N_3324);
nand U4033 (N_4033,N_3909,N_3130);
xor U4034 (N_4034,N_3270,N_3825);
and U4035 (N_4035,N_3753,N_3752);
xnor U4036 (N_4036,N_3982,N_3839);
nor U4037 (N_4037,N_3187,N_3997);
xor U4038 (N_4038,N_3273,N_3235);
nor U4039 (N_4039,N_3412,N_3323);
xnor U4040 (N_4040,N_3592,N_3197);
xnor U4041 (N_4041,N_3981,N_3305);
and U4042 (N_4042,N_3109,N_3979);
and U4043 (N_4043,N_3897,N_3377);
nand U4044 (N_4044,N_3929,N_3026);
and U4045 (N_4045,N_3133,N_3240);
xor U4046 (N_4046,N_3047,N_3884);
or U4047 (N_4047,N_3732,N_3201);
nor U4048 (N_4048,N_3986,N_3332);
nor U4049 (N_4049,N_3847,N_3088);
xor U4050 (N_4050,N_3819,N_3193);
nand U4051 (N_4051,N_3290,N_3397);
or U4052 (N_4052,N_3551,N_3129);
nand U4053 (N_4053,N_3171,N_3087);
or U4054 (N_4054,N_3462,N_3914);
xor U4055 (N_4055,N_3413,N_3809);
nor U4056 (N_4056,N_3777,N_3730);
nand U4057 (N_4057,N_3858,N_3346);
or U4058 (N_4058,N_3706,N_3774);
and U4059 (N_4059,N_3209,N_3424);
or U4060 (N_4060,N_3905,N_3713);
nand U4061 (N_4061,N_3518,N_3217);
nor U4062 (N_4062,N_3029,N_3439);
xor U4063 (N_4063,N_3159,N_3435);
nand U4064 (N_4064,N_3091,N_3155);
or U4065 (N_4065,N_3670,N_3110);
nor U4066 (N_4066,N_3703,N_3535);
xnor U4067 (N_4067,N_3264,N_3971);
or U4068 (N_4068,N_3105,N_3946);
or U4069 (N_4069,N_3434,N_3214);
xnor U4070 (N_4070,N_3379,N_3891);
or U4071 (N_4071,N_3765,N_3722);
nor U4072 (N_4072,N_3671,N_3226);
and U4073 (N_4073,N_3627,N_3973);
or U4074 (N_4074,N_3402,N_3131);
nand U4075 (N_4075,N_3805,N_3447);
xor U4076 (N_4076,N_3547,N_3530);
nor U4077 (N_4077,N_3684,N_3860);
nand U4078 (N_4078,N_3983,N_3330);
xnor U4079 (N_4079,N_3716,N_3189);
xor U4080 (N_4080,N_3608,N_3553);
nand U4081 (N_4081,N_3137,N_3861);
nand U4082 (N_4082,N_3183,N_3296);
nand U4083 (N_4083,N_3792,N_3212);
nand U4084 (N_4084,N_3167,N_3987);
xor U4085 (N_4085,N_3911,N_3350);
xnor U4086 (N_4086,N_3272,N_3190);
nand U4087 (N_4087,N_3688,N_3779);
nor U4088 (N_4088,N_3814,N_3248);
xor U4089 (N_4089,N_3475,N_3116);
and U4090 (N_4090,N_3181,N_3123);
and U4091 (N_4091,N_3401,N_3628);
or U4092 (N_4092,N_3606,N_3431);
or U4093 (N_4093,N_3122,N_3542);
or U4094 (N_4094,N_3045,N_3938);
or U4095 (N_4095,N_3104,N_3165);
xnor U4096 (N_4096,N_3180,N_3658);
nor U4097 (N_4097,N_3913,N_3822);
nand U4098 (N_4098,N_3354,N_3005);
nand U4099 (N_4099,N_3618,N_3344);
nor U4100 (N_4100,N_3966,N_3310);
or U4101 (N_4101,N_3830,N_3561);
nor U4102 (N_4102,N_3650,N_3112);
or U4103 (N_4103,N_3136,N_3036);
or U4104 (N_4104,N_3299,N_3154);
xor U4105 (N_4105,N_3124,N_3828);
nor U4106 (N_4106,N_3877,N_3457);
or U4107 (N_4107,N_3666,N_3236);
nand U4108 (N_4108,N_3169,N_3994);
or U4109 (N_4109,N_3019,N_3003);
xnor U4110 (N_4110,N_3195,N_3466);
nor U4111 (N_4111,N_3661,N_3705);
or U4112 (N_4112,N_3051,N_3843);
nand U4113 (N_4113,N_3364,N_3500);
xor U4114 (N_4114,N_3651,N_3559);
nand U4115 (N_4115,N_3662,N_3623);
xor U4116 (N_4116,N_3338,N_3325);
and U4117 (N_4117,N_3511,N_3333);
and U4118 (N_4118,N_3601,N_3725);
or U4119 (N_4119,N_3001,N_3773);
or U4120 (N_4120,N_3506,N_3149);
nand U4121 (N_4121,N_3077,N_3778);
or U4122 (N_4122,N_3943,N_3985);
nor U4123 (N_4123,N_3414,N_3140);
and U4124 (N_4124,N_3150,N_3921);
xnor U4125 (N_4125,N_3892,N_3292);
xnor U4126 (N_4126,N_3630,N_3875);
and U4127 (N_4127,N_3358,N_3262);
and U4128 (N_4128,N_3285,N_3527);
and U4129 (N_4129,N_3539,N_3253);
or U4130 (N_4130,N_3526,N_3883);
or U4131 (N_4131,N_3229,N_3524);
nand U4132 (N_4132,N_3761,N_3611);
xnor U4133 (N_4133,N_3655,N_3505);
or U4134 (N_4134,N_3249,N_3378);
nor U4135 (N_4135,N_3629,N_3933);
or U4136 (N_4136,N_3329,N_3081);
or U4137 (N_4137,N_3867,N_3121);
xor U4138 (N_4138,N_3782,N_3799);
xnor U4139 (N_4139,N_3967,N_3614);
or U4140 (N_4140,N_3563,N_3465);
or U4141 (N_4141,N_3558,N_3836);
nor U4142 (N_4142,N_3175,N_3991);
nand U4143 (N_4143,N_3009,N_3764);
nand U4144 (N_4144,N_3297,N_3536);
and U4145 (N_4145,N_3334,N_3522);
and U4146 (N_4146,N_3489,N_3743);
xnor U4147 (N_4147,N_3996,N_3342);
xor U4148 (N_4148,N_3158,N_3676);
nor U4149 (N_4149,N_3652,N_3544);
nand U4150 (N_4150,N_3701,N_3570);
nor U4151 (N_4151,N_3886,N_3486);
or U4152 (N_4152,N_3138,N_3053);
or U4153 (N_4153,N_3746,N_3284);
nand U4154 (N_4154,N_3793,N_3709);
or U4155 (N_4155,N_3492,N_3244);
xnor U4156 (N_4156,N_3796,N_3487);
and U4157 (N_4157,N_3755,N_3404);
or U4158 (N_4158,N_3926,N_3862);
and U4159 (N_4159,N_3633,N_3071);
nand U4160 (N_4160,N_3857,N_3308);
or U4161 (N_4161,N_3128,N_3501);
nand U4162 (N_4162,N_3920,N_3694);
or U4163 (N_4163,N_3554,N_3776);
nor U4164 (N_4164,N_3034,N_3198);
xor U4165 (N_4165,N_3800,N_3215);
xnor U4166 (N_4166,N_3969,N_3281);
and U4167 (N_4167,N_3010,N_3636);
and U4168 (N_4168,N_3795,N_3202);
nor U4169 (N_4169,N_3049,N_3221);
nor U4170 (N_4170,N_3718,N_3280);
nand U4171 (N_4171,N_3978,N_3361);
nor U4172 (N_4172,N_3758,N_3469);
nand U4173 (N_4173,N_3147,N_3854);
xnor U4174 (N_4174,N_3251,N_3020);
or U4175 (N_4175,N_3459,N_3549);
and U4176 (N_4176,N_3476,N_3096);
xor U4177 (N_4177,N_3609,N_3733);
and U4178 (N_4178,N_3869,N_3894);
and U4179 (N_4179,N_3211,N_3375);
or U4180 (N_4180,N_3493,N_3844);
or U4181 (N_4181,N_3863,N_3394);
nor U4182 (N_4182,N_3495,N_3974);
and U4183 (N_4183,N_3355,N_3620);
and U4184 (N_4184,N_3163,N_3507);
or U4185 (N_4185,N_3277,N_3679);
and U4186 (N_4186,N_3832,N_3889);
nand U4187 (N_4187,N_3184,N_3744);
xor U4188 (N_4188,N_3007,N_3279);
xor U4189 (N_4189,N_3372,N_3739);
or U4190 (N_4190,N_3977,N_3833);
and U4191 (N_4191,N_3515,N_3135);
nand U4192 (N_4192,N_3616,N_3728);
nand U4193 (N_4193,N_3213,N_3427);
nor U4194 (N_4194,N_3516,N_3428);
xor U4195 (N_4195,N_3496,N_3399);
or U4196 (N_4196,N_3808,N_3798);
nor U4197 (N_4197,N_3182,N_3474);
nor U4198 (N_4198,N_3696,N_3637);
xor U4199 (N_4199,N_3812,N_3306);
nor U4200 (N_4200,N_3174,N_3455);
and U4201 (N_4201,N_3579,N_3494);
or U4202 (N_4202,N_3864,N_3056);
nand U4203 (N_4203,N_3360,N_3786);
and U4204 (N_4204,N_3908,N_3995);
and U4205 (N_4205,N_3815,N_3328);
and U4206 (N_4206,N_3960,N_3754);
and U4207 (N_4207,N_3803,N_3031);
and U4208 (N_4208,N_3529,N_3014);
xnor U4209 (N_4209,N_3956,N_3008);
or U4210 (N_4210,N_3757,N_3200);
and U4211 (N_4211,N_3321,N_3856);
and U4212 (N_4212,N_3667,N_3421);
nand U4213 (N_4213,N_3120,N_3613);
and U4214 (N_4214,N_3371,N_3783);
xnor U4215 (N_4215,N_3680,N_3589);
nor U4216 (N_4216,N_3456,N_3035);
nor U4217 (N_4217,N_3153,N_3384);
nor U4218 (N_4218,N_3102,N_3999);
or U4219 (N_4219,N_3572,N_3263);
nand U4220 (N_4220,N_3513,N_3626);
nand U4221 (N_4221,N_3576,N_3924);
nand U4222 (N_4222,N_3937,N_3851);
xor U4223 (N_4223,N_3093,N_3313);
nor U4224 (N_4224,N_3052,N_3600);
and U4225 (N_4225,N_3044,N_3834);
nand U4226 (N_4226,N_3873,N_3898);
nor U4227 (N_4227,N_3239,N_3993);
or U4228 (N_4228,N_3910,N_3257);
or U4229 (N_4229,N_3002,N_3641);
nor U4230 (N_4230,N_3022,N_3018);
and U4231 (N_4231,N_3132,N_3704);
and U4232 (N_4232,N_3635,N_3980);
or U4233 (N_4233,N_3681,N_3692);
and U4234 (N_4234,N_3433,N_3508);
xor U4235 (N_4235,N_3726,N_3144);
nor U4236 (N_4236,N_3082,N_3759);
xnor U4237 (N_4237,N_3359,N_3737);
nand U4238 (N_4238,N_3567,N_3293);
nor U4239 (N_4239,N_3139,N_3170);
and U4240 (N_4240,N_3177,N_3231);
xor U4241 (N_4241,N_3578,N_3069);
and U4242 (N_4242,N_3318,N_3598);
nand U4243 (N_4243,N_3420,N_3942);
xor U4244 (N_4244,N_3634,N_3070);
xnor U4245 (N_4245,N_3497,N_3315);
or U4246 (N_4246,N_3464,N_3972);
xor U4247 (N_4247,N_3975,N_3958);
xnor U4248 (N_4248,N_3023,N_3168);
nor U4249 (N_4249,N_3042,N_3254);
and U4250 (N_4250,N_3788,N_3848);
and U4251 (N_4251,N_3657,N_3396);
nor U4252 (N_4252,N_3368,N_3574);
xnor U4253 (N_4253,N_3024,N_3899);
or U4254 (N_4254,N_3829,N_3407);
or U4255 (N_4255,N_3453,N_3702);
nor U4256 (N_4256,N_3811,N_3593);
nor U4257 (N_4257,N_3890,N_3481);
nand U4258 (N_4258,N_3649,N_3260);
and U4259 (N_4259,N_3970,N_3117);
nor U4260 (N_4260,N_3562,N_3349);
and U4261 (N_4261,N_3690,N_3341);
xnor U4262 (N_4262,N_3068,N_3677);
or U4263 (N_4263,N_3157,N_3689);
nor U4264 (N_4264,N_3963,N_3919);
nor U4265 (N_4265,N_3432,N_3237);
nand U4266 (N_4266,N_3640,N_3686);
or U4267 (N_4267,N_3065,N_3648);
nand U4268 (N_4268,N_3365,N_3055);
or U4269 (N_4269,N_3707,N_3719);
nor U4270 (N_4270,N_3419,N_3988);
and U4271 (N_4271,N_3269,N_3232);
xnor U4272 (N_4272,N_3588,N_3442);
nand U4273 (N_4273,N_3250,N_3738);
xnor U4274 (N_4274,N_3204,N_3415);
xor U4275 (N_4275,N_3727,N_3691);
or U4276 (N_4276,N_3780,N_3656);
nand U4277 (N_4277,N_3115,N_3653);
xor U4278 (N_4278,N_3438,N_3556);
nand U4279 (N_4279,N_3143,N_3763);
nor U4280 (N_4280,N_3537,N_3896);
nor U4281 (N_4281,N_3472,N_3859);
nor U4282 (N_4282,N_3079,N_3741);
nand U4283 (N_4283,N_3760,N_3199);
and U4284 (N_4284,N_3309,N_3944);
and U4285 (N_4285,N_3906,N_3503);
nor U4286 (N_4286,N_3160,N_3196);
xor U4287 (N_4287,N_3430,N_3810);
xor U4288 (N_4288,N_3451,N_3080);
and U4289 (N_4289,N_3876,N_3006);
nor U4290 (N_4290,N_3085,N_3723);
nor U4291 (N_4291,N_3103,N_3370);
nor U4292 (N_4292,N_3827,N_3514);
nand U4293 (N_4293,N_3710,N_3203);
nor U4294 (N_4294,N_3882,N_3048);
or U4295 (N_4295,N_3317,N_3916);
or U4296 (N_4296,N_3928,N_3258);
or U4297 (N_4297,N_3931,N_3186);
nand U4298 (N_4298,N_3669,N_3842);
and U4299 (N_4299,N_3113,N_3577);
nor U4300 (N_4300,N_3098,N_3504);
nor U4301 (N_4301,N_3918,N_3852);
nor U4302 (N_4302,N_3107,N_3478);
nand U4303 (N_4303,N_3473,N_3904);
or U4304 (N_4304,N_3327,N_3715);
nor U4305 (N_4305,N_3756,N_3801);
xnor U4306 (N_4306,N_3724,N_3312);
or U4307 (N_4307,N_3298,N_3021);
and U4308 (N_4308,N_3063,N_3583);
and U4309 (N_4309,N_3708,N_3145);
xor U4310 (N_4310,N_3271,N_3736);
nand U4311 (N_4311,N_3188,N_3223);
nand U4312 (N_4312,N_3295,N_3826);
xnor U4313 (N_4313,N_3408,N_3903);
nand U4314 (N_4314,N_3423,N_3114);
nand U4315 (N_4315,N_3984,N_3654);
or U4316 (N_4316,N_3820,N_3289);
nor U4317 (N_4317,N_3222,N_3804);
xnor U4318 (N_4318,N_3276,N_3286);
or U4319 (N_4319,N_3381,N_3385);
nor U4320 (N_4320,N_3612,N_3353);
nand U4321 (N_4321,N_3871,N_3550);
nand U4322 (N_4322,N_3386,N_3134);
or U4323 (N_4323,N_3278,N_3017);
xnor U4324 (N_4324,N_3721,N_3441);
xor U4325 (N_4325,N_3340,N_3030);
nor U4326 (N_4326,N_3543,N_3769);
nor U4327 (N_4327,N_3604,N_3205);
and U4328 (N_4328,N_3595,N_3745);
or U4329 (N_4329,N_3552,N_3821);
nor U4330 (N_4330,N_3720,N_3078);
and U4331 (N_4331,N_3234,N_3599);
and U4332 (N_4332,N_3638,N_3066);
nor U4333 (N_4333,N_3772,N_3521);
or U4334 (N_4334,N_3224,N_3480);
nor U4335 (N_4335,N_3060,N_3099);
nor U4336 (N_4336,N_3300,N_3872);
xor U4337 (N_4337,N_3336,N_3925);
xor U4338 (N_4338,N_3714,N_3075);
xnor U4339 (N_4339,N_3437,N_3619);
and U4340 (N_4340,N_3092,N_3206);
nor U4341 (N_4341,N_3108,N_3040);
nor U4342 (N_4342,N_3191,N_3711);
nand U4343 (N_4343,N_3268,N_3443);
or U4344 (N_4344,N_3603,N_3885);
xor U4345 (N_4345,N_3225,N_3930);
nor U4346 (N_4346,N_3454,N_3125);
and U4347 (N_4347,N_3747,N_3301);
xor U4348 (N_4348,N_3000,N_3436);
and U4349 (N_4349,N_3957,N_3953);
nand U4350 (N_4350,N_3220,N_3951);
nand U4351 (N_4351,N_3639,N_3740);
nand U4352 (N_4352,N_3194,N_3964);
nor U4353 (N_4353,N_3176,N_3094);
and U4354 (N_4354,N_3596,N_3917);
xnor U4355 (N_4355,N_3564,N_3850);
nor U4356 (N_4356,N_3389,N_3768);
nor U4357 (N_4357,N_3319,N_3357);
nand U4358 (N_4358,N_3127,N_3059);
and U4359 (N_4359,N_3173,N_3675);
xor U4360 (N_4360,N_3569,N_3693);
nand U4361 (N_4361,N_3038,N_3687);
and U4362 (N_4362,N_3448,N_3410);
nand U4363 (N_4363,N_3089,N_3712);
nand U4364 (N_4364,N_3161,N_3207);
nand U4365 (N_4365,N_3868,N_3084);
xnor U4366 (N_4366,N_3785,N_3491);
and U4367 (N_4367,N_3621,N_3597);
and U4368 (N_4368,N_3631,N_3106);
or U4369 (N_4369,N_3735,N_3512);
and U4370 (N_4370,N_3445,N_3870);
nand U4371 (N_4371,N_3267,N_3927);
nand U4372 (N_4372,N_3699,N_3646);
and U4373 (N_4373,N_3731,N_3050);
and U4374 (N_4374,N_3751,N_3775);
and U4375 (N_4375,N_3902,N_3162);
nand U4376 (N_4376,N_3320,N_3179);
or U4377 (N_4377,N_3900,N_3352);
and U4378 (N_4378,N_3146,N_3767);
and U4379 (N_4379,N_3922,N_3949);
or U4380 (N_4380,N_3418,N_3887);
xnor U4381 (N_4381,N_3054,N_3417);
and U4382 (N_4382,N_3945,N_3762);
nor U4383 (N_4383,N_3817,N_3797);
nor U4384 (N_4384,N_3450,N_3452);
nor U4385 (N_4385,N_3742,N_3695);
nor U4386 (N_4386,N_3625,N_3990);
or U4387 (N_4387,N_3645,N_3528);
nand U4388 (N_4388,N_3560,N_3241);
nor U4389 (N_4389,N_3057,N_3178);
and U4390 (N_4390,N_3291,N_3643);
and U4391 (N_4391,N_3393,N_3283);
and U4392 (N_4392,N_3164,N_3895);
or U4393 (N_4393,N_3934,N_3090);
nor U4394 (N_4394,N_3565,N_3510);
nor U4395 (N_4395,N_3400,N_3073);
and U4396 (N_4396,N_3383,N_3274);
and U4397 (N_4397,N_3520,N_3749);
or U4398 (N_4398,N_3345,N_3682);
or U4399 (N_4399,N_3256,N_3532);
xnor U4400 (N_4400,N_3893,N_3586);
nor U4401 (N_4401,N_3865,N_3879);
xor U4402 (N_4402,N_3192,N_3247);
or U4403 (N_4403,N_3288,N_3208);
xor U4404 (N_4404,N_3545,N_3622);
or U4405 (N_4405,N_3700,N_3664);
or U4406 (N_4406,N_3482,N_3575);
and U4407 (N_4407,N_3266,N_3659);
or U4408 (N_4408,N_3366,N_3259);
nor U4409 (N_4409,N_3101,N_3807);
and U4410 (N_4410,N_3152,N_3037);
or U4411 (N_4411,N_3304,N_3369);
or U4412 (N_4412,N_3923,N_3218);
and U4413 (N_4413,N_3376,N_3853);
nor U4414 (N_4414,N_3907,N_3647);
nand U4415 (N_4415,N_3275,N_3940);
nand U4416 (N_4416,N_3791,N_3411);
nor U4417 (N_4417,N_3568,N_3594);
xnor U4418 (N_4418,N_3245,N_3548);
and U4419 (N_4419,N_3185,N_3348);
nor U4420 (N_4420,N_3959,N_3151);
or U4421 (N_4421,N_3816,N_3962);
or U4422 (N_4422,N_3555,N_3584);
nand U4423 (N_4423,N_3074,N_3086);
nor U4424 (N_4424,N_3717,N_3498);
or U4425 (N_4425,N_3605,N_3525);
or U4426 (N_4426,N_3233,N_3467);
nor U4427 (N_4427,N_3343,N_3632);
or U4428 (N_4428,N_3356,N_3965);
or U4429 (N_4429,N_3043,N_3734);
or U4430 (N_4430,N_3013,N_3581);
nor U4431 (N_4431,N_3390,N_3642);
nor U4432 (N_4432,N_3531,N_3770);
or U4433 (N_4433,N_3337,N_3483);
nor U4434 (N_4434,N_3668,N_3238);
and U4435 (N_4435,N_3947,N_3302);
or U4436 (N_4436,N_3025,N_3939);
and U4437 (N_4437,N_3416,N_3072);
nor U4438 (N_4438,N_3463,N_3771);
nor U4439 (N_4439,N_3219,N_3287);
nand U4440 (N_4440,N_3582,N_3488);
nor U4441 (N_4441,N_3665,N_3968);
and U4442 (N_4442,N_3663,N_3046);
or U4443 (N_4443,N_3935,N_3403);
nor U4444 (N_4444,N_3380,N_3387);
nand U4445 (N_4445,N_3172,N_3265);
nor U4446 (N_4446,N_3624,N_3585);
nor U4447 (N_4447,N_3750,N_3367);
and U4448 (N_4448,N_3824,N_3866);
or U4449 (N_4449,N_3901,N_3362);
or U4450 (N_4450,N_3538,N_3316);
or U4451 (N_4451,N_3041,N_3426);
or U4452 (N_4452,N_3032,N_3541);
nor U4453 (N_4453,N_3294,N_3835);
nor U4454 (N_4454,N_3449,N_3789);
and U4455 (N_4455,N_3406,N_3660);
xnor U4456 (N_4456,N_3557,N_3485);
or U4457 (N_4457,N_3405,N_3948);
and U4458 (N_4458,N_3339,N_3461);
or U4459 (N_4459,N_3119,N_3216);
and U4460 (N_4460,N_3881,N_3837);
nor U4461 (N_4461,N_3061,N_3915);
and U4462 (N_4462,N_3794,N_3118);
nor U4463 (N_4463,N_3012,N_3615);
nand U4464 (N_4464,N_3813,N_3992);
xnor U4465 (N_4465,N_3818,N_3429);
nor U4466 (N_4466,N_3602,N_3391);
xnor U4467 (N_4467,N_3307,N_3230);
or U4468 (N_4468,N_3058,N_3440);
and U4469 (N_4469,N_3888,N_3523);
nand U4470 (N_4470,N_3374,N_3874);
and U4471 (N_4471,N_3950,N_3849);
or U4472 (N_4472,N_3571,N_3067);
or U4473 (N_4473,N_3111,N_3004);
or U4474 (N_4474,N_3610,N_3458);
and U4475 (N_4475,N_3781,N_3425);
and U4476 (N_4476,N_3255,N_3955);
or U4477 (N_4477,N_3100,N_3142);
xor U4478 (N_4478,N_3261,N_3015);
xor U4479 (N_4479,N_3242,N_3766);
xnor U4480 (N_4480,N_3683,N_3322);
xnor U4481 (N_4481,N_3444,N_3806);
nand U4482 (N_4482,N_3831,N_3685);
xnor U4483 (N_4483,N_3607,N_3382);
nor U4484 (N_4484,N_3471,N_3468);
nand U4485 (N_4485,N_3823,N_3484);
xnor U4486 (N_4486,N_3845,N_3989);
nand U4487 (N_4487,N_3326,N_3095);
nand U4488 (N_4488,N_3016,N_3097);
xnor U4489 (N_4489,N_3932,N_3729);
or U4490 (N_4490,N_3674,N_3210);
xor U4491 (N_4491,N_3954,N_3252);
nor U4492 (N_4492,N_3998,N_3064);
nor U4493 (N_4493,N_3282,N_3587);
xnor U4494 (N_4494,N_3617,N_3363);
and U4495 (N_4495,N_3392,N_3303);
or U4496 (N_4496,N_3802,N_3141);
nor U4497 (N_4497,N_3126,N_3546);
and U4498 (N_4498,N_3540,N_3534);
nand U4499 (N_4499,N_3446,N_3166);
xor U4500 (N_4500,N_3976,N_3241);
or U4501 (N_4501,N_3453,N_3736);
and U4502 (N_4502,N_3438,N_3036);
and U4503 (N_4503,N_3052,N_3442);
or U4504 (N_4504,N_3838,N_3397);
nor U4505 (N_4505,N_3549,N_3550);
or U4506 (N_4506,N_3787,N_3537);
or U4507 (N_4507,N_3108,N_3945);
nand U4508 (N_4508,N_3497,N_3659);
nor U4509 (N_4509,N_3876,N_3746);
or U4510 (N_4510,N_3113,N_3604);
and U4511 (N_4511,N_3144,N_3376);
nand U4512 (N_4512,N_3954,N_3251);
xor U4513 (N_4513,N_3458,N_3400);
or U4514 (N_4514,N_3664,N_3420);
nor U4515 (N_4515,N_3559,N_3831);
and U4516 (N_4516,N_3259,N_3383);
or U4517 (N_4517,N_3534,N_3931);
or U4518 (N_4518,N_3422,N_3563);
and U4519 (N_4519,N_3465,N_3562);
xnor U4520 (N_4520,N_3798,N_3091);
xor U4521 (N_4521,N_3794,N_3522);
and U4522 (N_4522,N_3156,N_3958);
nor U4523 (N_4523,N_3149,N_3056);
nand U4524 (N_4524,N_3170,N_3630);
xnor U4525 (N_4525,N_3498,N_3764);
nand U4526 (N_4526,N_3379,N_3062);
xor U4527 (N_4527,N_3969,N_3466);
nor U4528 (N_4528,N_3611,N_3013);
or U4529 (N_4529,N_3141,N_3110);
and U4530 (N_4530,N_3170,N_3295);
nand U4531 (N_4531,N_3718,N_3238);
nand U4532 (N_4532,N_3437,N_3515);
nor U4533 (N_4533,N_3602,N_3411);
nand U4534 (N_4534,N_3068,N_3299);
nor U4535 (N_4535,N_3672,N_3690);
and U4536 (N_4536,N_3144,N_3898);
nand U4537 (N_4537,N_3157,N_3494);
and U4538 (N_4538,N_3300,N_3572);
or U4539 (N_4539,N_3246,N_3237);
nor U4540 (N_4540,N_3539,N_3935);
nor U4541 (N_4541,N_3930,N_3588);
nand U4542 (N_4542,N_3903,N_3969);
or U4543 (N_4543,N_3748,N_3676);
nand U4544 (N_4544,N_3581,N_3819);
nand U4545 (N_4545,N_3353,N_3352);
or U4546 (N_4546,N_3589,N_3005);
nor U4547 (N_4547,N_3276,N_3168);
and U4548 (N_4548,N_3157,N_3514);
or U4549 (N_4549,N_3553,N_3718);
or U4550 (N_4550,N_3562,N_3714);
or U4551 (N_4551,N_3014,N_3192);
and U4552 (N_4552,N_3131,N_3996);
and U4553 (N_4553,N_3110,N_3696);
xor U4554 (N_4554,N_3342,N_3206);
xor U4555 (N_4555,N_3360,N_3217);
or U4556 (N_4556,N_3210,N_3715);
or U4557 (N_4557,N_3811,N_3878);
nor U4558 (N_4558,N_3071,N_3852);
or U4559 (N_4559,N_3785,N_3637);
nor U4560 (N_4560,N_3844,N_3692);
xor U4561 (N_4561,N_3011,N_3874);
and U4562 (N_4562,N_3501,N_3190);
xnor U4563 (N_4563,N_3668,N_3781);
nor U4564 (N_4564,N_3557,N_3710);
or U4565 (N_4565,N_3066,N_3844);
nand U4566 (N_4566,N_3175,N_3700);
xor U4567 (N_4567,N_3247,N_3167);
or U4568 (N_4568,N_3958,N_3153);
and U4569 (N_4569,N_3232,N_3624);
or U4570 (N_4570,N_3704,N_3316);
nand U4571 (N_4571,N_3591,N_3077);
and U4572 (N_4572,N_3572,N_3399);
nand U4573 (N_4573,N_3120,N_3737);
or U4574 (N_4574,N_3848,N_3039);
nand U4575 (N_4575,N_3965,N_3958);
nor U4576 (N_4576,N_3767,N_3201);
nand U4577 (N_4577,N_3315,N_3554);
nor U4578 (N_4578,N_3756,N_3325);
nor U4579 (N_4579,N_3226,N_3524);
or U4580 (N_4580,N_3723,N_3826);
or U4581 (N_4581,N_3381,N_3554);
nand U4582 (N_4582,N_3062,N_3437);
nor U4583 (N_4583,N_3785,N_3032);
nor U4584 (N_4584,N_3064,N_3867);
or U4585 (N_4585,N_3274,N_3497);
and U4586 (N_4586,N_3017,N_3423);
and U4587 (N_4587,N_3197,N_3125);
nor U4588 (N_4588,N_3676,N_3254);
xnor U4589 (N_4589,N_3090,N_3730);
nand U4590 (N_4590,N_3591,N_3187);
nor U4591 (N_4591,N_3290,N_3782);
nand U4592 (N_4592,N_3352,N_3566);
nand U4593 (N_4593,N_3184,N_3232);
or U4594 (N_4594,N_3667,N_3535);
xor U4595 (N_4595,N_3687,N_3033);
nand U4596 (N_4596,N_3580,N_3637);
and U4597 (N_4597,N_3892,N_3286);
and U4598 (N_4598,N_3492,N_3692);
nor U4599 (N_4599,N_3120,N_3638);
or U4600 (N_4600,N_3743,N_3970);
or U4601 (N_4601,N_3454,N_3705);
nor U4602 (N_4602,N_3330,N_3867);
nor U4603 (N_4603,N_3424,N_3733);
nor U4604 (N_4604,N_3276,N_3347);
nand U4605 (N_4605,N_3967,N_3628);
and U4606 (N_4606,N_3851,N_3795);
or U4607 (N_4607,N_3475,N_3587);
nand U4608 (N_4608,N_3644,N_3987);
nor U4609 (N_4609,N_3670,N_3891);
nand U4610 (N_4610,N_3699,N_3621);
and U4611 (N_4611,N_3995,N_3145);
and U4612 (N_4612,N_3454,N_3485);
or U4613 (N_4613,N_3433,N_3340);
xnor U4614 (N_4614,N_3216,N_3372);
or U4615 (N_4615,N_3115,N_3991);
and U4616 (N_4616,N_3800,N_3179);
nand U4617 (N_4617,N_3835,N_3620);
and U4618 (N_4618,N_3487,N_3229);
nand U4619 (N_4619,N_3788,N_3899);
xnor U4620 (N_4620,N_3373,N_3490);
nor U4621 (N_4621,N_3463,N_3799);
xnor U4622 (N_4622,N_3512,N_3836);
nor U4623 (N_4623,N_3778,N_3749);
nor U4624 (N_4624,N_3962,N_3865);
xnor U4625 (N_4625,N_3765,N_3753);
nand U4626 (N_4626,N_3036,N_3271);
nand U4627 (N_4627,N_3475,N_3274);
nand U4628 (N_4628,N_3360,N_3296);
xor U4629 (N_4629,N_3182,N_3201);
and U4630 (N_4630,N_3730,N_3486);
or U4631 (N_4631,N_3781,N_3283);
and U4632 (N_4632,N_3398,N_3571);
xnor U4633 (N_4633,N_3820,N_3508);
xor U4634 (N_4634,N_3632,N_3425);
or U4635 (N_4635,N_3714,N_3287);
nor U4636 (N_4636,N_3446,N_3988);
and U4637 (N_4637,N_3393,N_3086);
nor U4638 (N_4638,N_3708,N_3182);
or U4639 (N_4639,N_3031,N_3100);
or U4640 (N_4640,N_3735,N_3899);
nand U4641 (N_4641,N_3342,N_3001);
and U4642 (N_4642,N_3337,N_3017);
nand U4643 (N_4643,N_3564,N_3106);
or U4644 (N_4644,N_3319,N_3293);
and U4645 (N_4645,N_3835,N_3364);
nand U4646 (N_4646,N_3899,N_3676);
nand U4647 (N_4647,N_3659,N_3780);
xor U4648 (N_4648,N_3975,N_3269);
xor U4649 (N_4649,N_3002,N_3240);
nor U4650 (N_4650,N_3024,N_3829);
and U4651 (N_4651,N_3925,N_3907);
or U4652 (N_4652,N_3914,N_3543);
xor U4653 (N_4653,N_3178,N_3012);
nor U4654 (N_4654,N_3724,N_3859);
nand U4655 (N_4655,N_3236,N_3011);
or U4656 (N_4656,N_3306,N_3256);
nand U4657 (N_4657,N_3292,N_3034);
or U4658 (N_4658,N_3808,N_3107);
xor U4659 (N_4659,N_3821,N_3896);
nand U4660 (N_4660,N_3367,N_3653);
or U4661 (N_4661,N_3790,N_3011);
or U4662 (N_4662,N_3989,N_3971);
xor U4663 (N_4663,N_3007,N_3853);
nor U4664 (N_4664,N_3070,N_3392);
nand U4665 (N_4665,N_3208,N_3959);
nand U4666 (N_4666,N_3059,N_3274);
nand U4667 (N_4667,N_3471,N_3023);
and U4668 (N_4668,N_3172,N_3794);
nor U4669 (N_4669,N_3793,N_3002);
nor U4670 (N_4670,N_3370,N_3622);
nand U4671 (N_4671,N_3818,N_3951);
or U4672 (N_4672,N_3509,N_3182);
nand U4673 (N_4673,N_3454,N_3384);
nor U4674 (N_4674,N_3639,N_3628);
and U4675 (N_4675,N_3667,N_3032);
xor U4676 (N_4676,N_3602,N_3729);
xor U4677 (N_4677,N_3815,N_3851);
and U4678 (N_4678,N_3637,N_3826);
or U4679 (N_4679,N_3215,N_3927);
and U4680 (N_4680,N_3249,N_3795);
and U4681 (N_4681,N_3490,N_3375);
or U4682 (N_4682,N_3023,N_3068);
or U4683 (N_4683,N_3904,N_3802);
and U4684 (N_4684,N_3772,N_3245);
nor U4685 (N_4685,N_3657,N_3365);
nor U4686 (N_4686,N_3079,N_3953);
xor U4687 (N_4687,N_3440,N_3966);
and U4688 (N_4688,N_3074,N_3947);
or U4689 (N_4689,N_3770,N_3831);
or U4690 (N_4690,N_3381,N_3546);
or U4691 (N_4691,N_3162,N_3635);
nand U4692 (N_4692,N_3739,N_3909);
nor U4693 (N_4693,N_3549,N_3911);
xnor U4694 (N_4694,N_3845,N_3872);
xnor U4695 (N_4695,N_3924,N_3721);
nand U4696 (N_4696,N_3413,N_3745);
and U4697 (N_4697,N_3117,N_3596);
xnor U4698 (N_4698,N_3951,N_3207);
nor U4699 (N_4699,N_3198,N_3860);
xor U4700 (N_4700,N_3644,N_3268);
xor U4701 (N_4701,N_3877,N_3795);
and U4702 (N_4702,N_3784,N_3889);
and U4703 (N_4703,N_3648,N_3758);
xor U4704 (N_4704,N_3700,N_3995);
and U4705 (N_4705,N_3862,N_3148);
nor U4706 (N_4706,N_3231,N_3770);
nand U4707 (N_4707,N_3132,N_3691);
and U4708 (N_4708,N_3162,N_3673);
nor U4709 (N_4709,N_3895,N_3915);
nor U4710 (N_4710,N_3768,N_3491);
and U4711 (N_4711,N_3612,N_3137);
nand U4712 (N_4712,N_3801,N_3293);
and U4713 (N_4713,N_3279,N_3924);
nand U4714 (N_4714,N_3969,N_3204);
nor U4715 (N_4715,N_3791,N_3668);
xnor U4716 (N_4716,N_3188,N_3654);
nor U4717 (N_4717,N_3488,N_3198);
xor U4718 (N_4718,N_3117,N_3229);
nor U4719 (N_4719,N_3533,N_3703);
nand U4720 (N_4720,N_3228,N_3822);
nor U4721 (N_4721,N_3880,N_3379);
nor U4722 (N_4722,N_3918,N_3073);
nand U4723 (N_4723,N_3730,N_3738);
nand U4724 (N_4724,N_3658,N_3228);
nand U4725 (N_4725,N_3335,N_3972);
xnor U4726 (N_4726,N_3289,N_3020);
and U4727 (N_4727,N_3625,N_3790);
and U4728 (N_4728,N_3006,N_3998);
nor U4729 (N_4729,N_3392,N_3096);
nand U4730 (N_4730,N_3651,N_3612);
or U4731 (N_4731,N_3064,N_3683);
and U4732 (N_4732,N_3401,N_3583);
nand U4733 (N_4733,N_3731,N_3279);
or U4734 (N_4734,N_3997,N_3120);
xnor U4735 (N_4735,N_3825,N_3445);
or U4736 (N_4736,N_3715,N_3437);
and U4737 (N_4737,N_3822,N_3627);
nor U4738 (N_4738,N_3347,N_3799);
or U4739 (N_4739,N_3832,N_3746);
nand U4740 (N_4740,N_3015,N_3867);
or U4741 (N_4741,N_3853,N_3506);
or U4742 (N_4742,N_3375,N_3015);
and U4743 (N_4743,N_3440,N_3833);
xnor U4744 (N_4744,N_3249,N_3329);
or U4745 (N_4745,N_3475,N_3127);
and U4746 (N_4746,N_3232,N_3033);
nand U4747 (N_4747,N_3894,N_3049);
or U4748 (N_4748,N_3252,N_3901);
nor U4749 (N_4749,N_3593,N_3758);
nor U4750 (N_4750,N_3328,N_3134);
xor U4751 (N_4751,N_3463,N_3384);
or U4752 (N_4752,N_3011,N_3083);
and U4753 (N_4753,N_3995,N_3582);
nor U4754 (N_4754,N_3180,N_3805);
nand U4755 (N_4755,N_3069,N_3078);
xor U4756 (N_4756,N_3107,N_3623);
and U4757 (N_4757,N_3883,N_3068);
xor U4758 (N_4758,N_3193,N_3051);
or U4759 (N_4759,N_3831,N_3524);
and U4760 (N_4760,N_3945,N_3683);
or U4761 (N_4761,N_3273,N_3804);
xnor U4762 (N_4762,N_3802,N_3498);
nand U4763 (N_4763,N_3674,N_3138);
and U4764 (N_4764,N_3172,N_3787);
and U4765 (N_4765,N_3216,N_3033);
and U4766 (N_4766,N_3340,N_3905);
or U4767 (N_4767,N_3967,N_3914);
and U4768 (N_4768,N_3741,N_3647);
nor U4769 (N_4769,N_3016,N_3512);
nor U4770 (N_4770,N_3458,N_3197);
xor U4771 (N_4771,N_3525,N_3867);
or U4772 (N_4772,N_3242,N_3849);
and U4773 (N_4773,N_3357,N_3155);
or U4774 (N_4774,N_3314,N_3261);
nand U4775 (N_4775,N_3473,N_3472);
or U4776 (N_4776,N_3903,N_3094);
nand U4777 (N_4777,N_3930,N_3505);
or U4778 (N_4778,N_3261,N_3748);
nor U4779 (N_4779,N_3745,N_3799);
or U4780 (N_4780,N_3708,N_3206);
nand U4781 (N_4781,N_3225,N_3525);
xnor U4782 (N_4782,N_3542,N_3642);
nor U4783 (N_4783,N_3354,N_3785);
and U4784 (N_4784,N_3601,N_3285);
nand U4785 (N_4785,N_3029,N_3382);
and U4786 (N_4786,N_3583,N_3484);
xor U4787 (N_4787,N_3782,N_3615);
or U4788 (N_4788,N_3933,N_3499);
nor U4789 (N_4789,N_3501,N_3464);
nor U4790 (N_4790,N_3399,N_3458);
nor U4791 (N_4791,N_3279,N_3624);
and U4792 (N_4792,N_3844,N_3031);
and U4793 (N_4793,N_3584,N_3387);
and U4794 (N_4794,N_3644,N_3124);
xnor U4795 (N_4795,N_3953,N_3876);
and U4796 (N_4796,N_3811,N_3319);
xnor U4797 (N_4797,N_3817,N_3601);
or U4798 (N_4798,N_3816,N_3789);
and U4799 (N_4799,N_3294,N_3063);
or U4800 (N_4800,N_3820,N_3464);
and U4801 (N_4801,N_3556,N_3467);
nor U4802 (N_4802,N_3519,N_3033);
nor U4803 (N_4803,N_3536,N_3932);
nand U4804 (N_4804,N_3003,N_3451);
nor U4805 (N_4805,N_3310,N_3211);
nor U4806 (N_4806,N_3397,N_3224);
nand U4807 (N_4807,N_3656,N_3112);
or U4808 (N_4808,N_3498,N_3581);
xnor U4809 (N_4809,N_3117,N_3998);
and U4810 (N_4810,N_3783,N_3477);
xor U4811 (N_4811,N_3976,N_3855);
xor U4812 (N_4812,N_3736,N_3719);
nand U4813 (N_4813,N_3838,N_3285);
xor U4814 (N_4814,N_3564,N_3050);
and U4815 (N_4815,N_3409,N_3534);
or U4816 (N_4816,N_3990,N_3530);
nor U4817 (N_4817,N_3002,N_3752);
nand U4818 (N_4818,N_3156,N_3618);
nand U4819 (N_4819,N_3689,N_3739);
and U4820 (N_4820,N_3294,N_3567);
nand U4821 (N_4821,N_3371,N_3767);
xor U4822 (N_4822,N_3996,N_3300);
or U4823 (N_4823,N_3897,N_3281);
and U4824 (N_4824,N_3622,N_3311);
and U4825 (N_4825,N_3313,N_3818);
and U4826 (N_4826,N_3708,N_3386);
or U4827 (N_4827,N_3570,N_3921);
and U4828 (N_4828,N_3526,N_3866);
and U4829 (N_4829,N_3821,N_3089);
or U4830 (N_4830,N_3147,N_3924);
or U4831 (N_4831,N_3338,N_3489);
and U4832 (N_4832,N_3150,N_3384);
or U4833 (N_4833,N_3207,N_3404);
nor U4834 (N_4834,N_3344,N_3693);
nor U4835 (N_4835,N_3548,N_3262);
or U4836 (N_4836,N_3638,N_3474);
or U4837 (N_4837,N_3307,N_3964);
nand U4838 (N_4838,N_3092,N_3997);
or U4839 (N_4839,N_3613,N_3206);
or U4840 (N_4840,N_3559,N_3816);
and U4841 (N_4841,N_3156,N_3369);
and U4842 (N_4842,N_3109,N_3418);
nand U4843 (N_4843,N_3514,N_3991);
or U4844 (N_4844,N_3893,N_3780);
nor U4845 (N_4845,N_3166,N_3833);
and U4846 (N_4846,N_3408,N_3444);
xor U4847 (N_4847,N_3398,N_3791);
and U4848 (N_4848,N_3909,N_3548);
nor U4849 (N_4849,N_3032,N_3706);
nor U4850 (N_4850,N_3401,N_3245);
nor U4851 (N_4851,N_3014,N_3088);
nand U4852 (N_4852,N_3414,N_3758);
nor U4853 (N_4853,N_3851,N_3833);
nor U4854 (N_4854,N_3053,N_3070);
nor U4855 (N_4855,N_3774,N_3855);
and U4856 (N_4856,N_3989,N_3332);
or U4857 (N_4857,N_3216,N_3480);
nand U4858 (N_4858,N_3165,N_3263);
xor U4859 (N_4859,N_3033,N_3379);
xor U4860 (N_4860,N_3972,N_3581);
xor U4861 (N_4861,N_3333,N_3958);
nor U4862 (N_4862,N_3584,N_3078);
or U4863 (N_4863,N_3446,N_3470);
xnor U4864 (N_4864,N_3821,N_3383);
nor U4865 (N_4865,N_3515,N_3395);
and U4866 (N_4866,N_3584,N_3657);
or U4867 (N_4867,N_3711,N_3317);
nor U4868 (N_4868,N_3108,N_3228);
xor U4869 (N_4869,N_3177,N_3100);
nand U4870 (N_4870,N_3547,N_3007);
xor U4871 (N_4871,N_3412,N_3893);
nor U4872 (N_4872,N_3229,N_3064);
nor U4873 (N_4873,N_3160,N_3996);
nand U4874 (N_4874,N_3243,N_3549);
or U4875 (N_4875,N_3323,N_3600);
nor U4876 (N_4876,N_3792,N_3498);
nand U4877 (N_4877,N_3541,N_3146);
and U4878 (N_4878,N_3276,N_3653);
or U4879 (N_4879,N_3967,N_3933);
nand U4880 (N_4880,N_3325,N_3175);
and U4881 (N_4881,N_3542,N_3798);
xor U4882 (N_4882,N_3176,N_3438);
nor U4883 (N_4883,N_3924,N_3906);
xor U4884 (N_4884,N_3983,N_3387);
xor U4885 (N_4885,N_3011,N_3349);
nand U4886 (N_4886,N_3191,N_3354);
xnor U4887 (N_4887,N_3942,N_3256);
and U4888 (N_4888,N_3508,N_3197);
or U4889 (N_4889,N_3004,N_3553);
and U4890 (N_4890,N_3922,N_3102);
nand U4891 (N_4891,N_3571,N_3254);
xor U4892 (N_4892,N_3234,N_3597);
or U4893 (N_4893,N_3578,N_3250);
nand U4894 (N_4894,N_3072,N_3332);
and U4895 (N_4895,N_3917,N_3653);
or U4896 (N_4896,N_3691,N_3337);
or U4897 (N_4897,N_3363,N_3007);
and U4898 (N_4898,N_3600,N_3711);
or U4899 (N_4899,N_3649,N_3572);
and U4900 (N_4900,N_3156,N_3491);
and U4901 (N_4901,N_3465,N_3066);
or U4902 (N_4902,N_3408,N_3083);
and U4903 (N_4903,N_3277,N_3224);
and U4904 (N_4904,N_3118,N_3366);
nand U4905 (N_4905,N_3327,N_3014);
nor U4906 (N_4906,N_3880,N_3280);
nand U4907 (N_4907,N_3905,N_3246);
xor U4908 (N_4908,N_3848,N_3876);
or U4909 (N_4909,N_3610,N_3619);
nand U4910 (N_4910,N_3123,N_3984);
and U4911 (N_4911,N_3660,N_3415);
nand U4912 (N_4912,N_3717,N_3966);
nand U4913 (N_4913,N_3908,N_3292);
nor U4914 (N_4914,N_3201,N_3791);
nand U4915 (N_4915,N_3050,N_3379);
nand U4916 (N_4916,N_3964,N_3908);
nor U4917 (N_4917,N_3844,N_3172);
nor U4918 (N_4918,N_3485,N_3857);
xnor U4919 (N_4919,N_3340,N_3844);
xnor U4920 (N_4920,N_3631,N_3511);
nor U4921 (N_4921,N_3280,N_3620);
or U4922 (N_4922,N_3083,N_3749);
or U4923 (N_4923,N_3333,N_3952);
nor U4924 (N_4924,N_3900,N_3692);
xnor U4925 (N_4925,N_3192,N_3425);
or U4926 (N_4926,N_3495,N_3304);
nor U4927 (N_4927,N_3879,N_3151);
nand U4928 (N_4928,N_3396,N_3259);
xnor U4929 (N_4929,N_3840,N_3263);
or U4930 (N_4930,N_3436,N_3185);
nor U4931 (N_4931,N_3699,N_3934);
or U4932 (N_4932,N_3958,N_3586);
or U4933 (N_4933,N_3676,N_3994);
xor U4934 (N_4934,N_3180,N_3939);
and U4935 (N_4935,N_3420,N_3176);
nand U4936 (N_4936,N_3752,N_3205);
nor U4937 (N_4937,N_3660,N_3847);
xor U4938 (N_4938,N_3465,N_3758);
xnor U4939 (N_4939,N_3702,N_3360);
xnor U4940 (N_4940,N_3582,N_3031);
xor U4941 (N_4941,N_3156,N_3393);
or U4942 (N_4942,N_3756,N_3694);
nor U4943 (N_4943,N_3344,N_3333);
and U4944 (N_4944,N_3250,N_3890);
xnor U4945 (N_4945,N_3455,N_3147);
nand U4946 (N_4946,N_3431,N_3864);
xor U4947 (N_4947,N_3042,N_3516);
or U4948 (N_4948,N_3162,N_3265);
nand U4949 (N_4949,N_3597,N_3965);
or U4950 (N_4950,N_3059,N_3808);
xor U4951 (N_4951,N_3251,N_3513);
nor U4952 (N_4952,N_3467,N_3549);
and U4953 (N_4953,N_3267,N_3931);
or U4954 (N_4954,N_3413,N_3058);
and U4955 (N_4955,N_3411,N_3587);
nor U4956 (N_4956,N_3172,N_3219);
nor U4957 (N_4957,N_3572,N_3161);
nor U4958 (N_4958,N_3741,N_3308);
nor U4959 (N_4959,N_3857,N_3649);
nand U4960 (N_4960,N_3918,N_3794);
nand U4961 (N_4961,N_3847,N_3763);
nor U4962 (N_4962,N_3243,N_3310);
and U4963 (N_4963,N_3212,N_3668);
and U4964 (N_4964,N_3070,N_3726);
nor U4965 (N_4965,N_3990,N_3655);
or U4966 (N_4966,N_3429,N_3122);
nand U4967 (N_4967,N_3934,N_3406);
nand U4968 (N_4968,N_3459,N_3568);
nor U4969 (N_4969,N_3079,N_3048);
nor U4970 (N_4970,N_3357,N_3813);
or U4971 (N_4971,N_3400,N_3380);
and U4972 (N_4972,N_3982,N_3295);
or U4973 (N_4973,N_3146,N_3164);
xnor U4974 (N_4974,N_3403,N_3858);
xnor U4975 (N_4975,N_3917,N_3418);
xnor U4976 (N_4976,N_3531,N_3064);
nor U4977 (N_4977,N_3056,N_3296);
and U4978 (N_4978,N_3428,N_3933);
and U4979 (N_4979,N_3373,N_3658);
nand U4980 (N_4980,N_3535,N_3986);
nand U4981 (N_4981,N_3804,N_3305);
xnor U4982 (N_4982,N_3455,N_3788);
and U4983 (N_4983,N_3559,N_3976);
nand U4984 (N_4984,N_3814,N_3149);
and U4985 (N_4985,N_3776,N_3491);
xor U4986 (N_4986,N_3948,N_3770);
or U4987 (N_4987,N_3599,N_3556);
nand U4988 (N_4988,N_3036,N_3440);
nand U4989 (N_4989,N_3646,N_3477);
nor U4990 (N_4990,N_3269,N_3075);
xnor U4991 (N_4991,N_3150,N_3296);
or U4992 (N_4992,N_3829,N_3537);
or U4993 (N_4993,N_3975,N_3982);
nor U4994 (N_4994,N_3144,N_3822);
or U4995 (N_4995,N_3916,N_3865);
nor U4996 (N_4996,N_3203,N_3372);
and U4997 (N_4997,N_3484,N_3974);
and U4998 (N_4998,N_3471,N_3076);
or U4999 (N_4999,N_3943,N_3345);
or U5000 (N_5000,N_4165,N_4685);
or U5001 (N_5001,N_4188,N_4997);
xnor U5002 (N_5002,N_4496,N_4507);
or U5003 (N_5003,N_4231,N_4099);
nor U5004 (N_5004,N_4925,N_4715);
and U5005 (N_5005,N_4641,N_4594);
and U5006 (N_5006,N_4215,N_4678);
nand U5007 (N_5007,N_4145,N_4491);
or U5008 (N_5008,N_4271,N_4088);
and U5009 (N_5009,N_4010,N_4295);
and U5010 (N_5010,N_4984,N_4541);
or U5011 (N_5011,N_4958,N_4636);
xnor U5012 (N_5012,N_4943,N_4481);
or U5013 (N_5013,N_4763,N_4954);
and U5014 (N_5014,N_4696,N_4385);
xnor U5015 (N_5015,N_4578,N_4094);
nor U5016 (N_5016,N_4966,N_4913);
nand U5017 (N_5017,N_4276,N_4151);
nor U5018 (N_5018,N_4645,N_4826);
or U5019 (N_5019,N_4164,N_4421);
nor U5020 (N_5020,N_4484,N_4005);
nor U5021 (N_5021,N_4803,N_4887);
nor U5022 (N_5022,N_4513,N_4509);
or U5023 (N_5023,N_4390,N_4771);
nor U5024 (N_5024,N_4173,N_4840);
xnor U5025 (N_5025,N_4653,N_4700);
and U5026 (N_5026,N_4764,N_4508);
nor U5027 (N_5027,N_4945,N_4667);
and U5028 (N_5028,N_4948,N_4460);
nor U5029 (N_5029,N_4790,N_4168);
xnor U5030 (N_5030,N_4120,N_4776);
xor U5031 (N_5031,N_4238,N_4643);
nand U5032 (N_5032,N_4569,N_4581);
nand U5033 (N_5033,N_4050,N_4918);
xor U5034 (N_5034,N_4848,N_4301);
and U5035 (N_5035,N_4247,N_4758);
nand U5036 (N_5036,N_4349,N_4822);
or U5037 (N_5037,N_4064,N_4703);
and U5038 (N_5038,N_4206,N_4072);
nand U5039 (N_5039,N_4767,N_4798);
nand U5040 (N_5040,N_4690,N_4038);
or U5041 (N_5041,N_4867,N_4724);
xor U5042 (N_5042,N_4116,N_4939);
nand U5043 (N_5043,N_4419,N_4067);
or U5044 (N_5044,N_4381,N_4191);
nor U5045 (N_5045,N_4051,N_4666);
xor U5046 (N_5046,N_4552,N_4418);
xnor U5047 (N_5047,N_4405,N_4792);
xor U5048 (N_5048,N_4772,N_4664);
or U5049 (N_5049,N_4674,N_4189);
and U5050 (N_5050,N_4902,N_4570);
xnor U5051 (N_5051,N_4382,N_4656);
or U5052 (N_5052,N_4222,N_4018);
nand U5053 (N_5053,N_4937,N_4808);
or U5054 (N_5054,N_4928,N_4519);
nand U5055 (N_5055,N_4981,N_4695);
xor U5056 (N_5056,N_4579,N_4609);
nor U5057 (N_5057,N_4339,N_4037);
nand U5058 (N_5058,N_4806,N_4103);
and U5059 (N_5059,N_4008,N_4976);
xnor U5060 (N_5060,N_4399,N_4490);
nand U5061 (N_5061,N_4911,N_4459);
and U5062 (N_5062,N_4415,N_4108);
and U5063 (N_5063,N_4726,N_4322);
and U5064 (N_5064,N_4982,N_4900);
or U5065 (N_5065,N_4081,N_4585);
nor U5066 (N_5066,N_4035,N_4029);
xnor U5067 (N_5067,N_4425,N_4175);
nand U5068 (N_5068,N_4102,N_4161);
nand U5069 (N_5069,N_4398,N_4407);
or U5070 (N_5070,N_4647,N_4410);
nor U5071 (N_5071,N_4422,N_4435);
and U5072 (N_5072,N_4548,N_4015);
or U5073 (N_5073,N_4528,N_4130);
and U5074 (N_5074,N_4242,N_4259);
nand U5075 (N_5075,N_4924,N_4572);
nor U5076 (N_5076,N_4575,N_4012);
or U5077 (N_5077,N_4992,N_4923);
xnor U5078 (N_5078,N_4794,N_4115);
and U5079 (N_5079,N_4731,N_4040);
and U5080 (N_5080,N_4371,N_4797);
xnor U5081 (N_5081,N_4174,N_4379);
nor U5082 (N_5082,N_4657,N_4553);
nand U5083 (N_5083,N_4394,N_4973);
nor U5084 (N_5084,N_4097,N_4563);
nor U5085 (N_5085,N_4733,N_4235);
nor U5086 (N_5086,N_4527,N_4250);
and U5087 (N_5087,N_4021,N_4256);
or U5088 (N_5088,N_4111,N_4178);
nand U5089 (N_5089,N_4310,N_4049);
and U5090 (N_5090,N_4327,N_4547);
or U5091 (N_5091,N_4367,N_4427);
nand U5092 (N_5092,N_4251,N_4866);
and U5093 (N_5093,N_4843,N_4677);
and U5094 (N_5094,N_4241,N_4908);
or U5095 (N_5095,N_4823,N_4558);
or U5096 (N_5096,N_4034,N_4462);
nand U5097 (N_5097,N_4068,N_4582);
or U5098 (N_5098,N_4863,N_4497);
or U5099 (N_5099,N_4078,N_4028);
nor U5100 (N_5100,N_4941,N_4538);
nand U5101 (N_5101,N_4543,N_4093);
nand U5102 (N_5102,N_4517,N_4603);
nand U5103 (N_5103,N_4030,N_4658);
xor U5104 (N_5104,N_4629,N_4267);
nor U5105 (N_5105,N_4205,N_4487);
xor U5106 (N_5106,N_4857,N_4488);
xor U5107 (N_5107,N_4395,N_4632);
nor U5108 (N_5108,N_4045,N_4545);
nand U5109 (N_5109,N_4475,N_4869);
nor U5110 (N_5110,N_4542,N_4461);
xnor U5111 (N_5111,N_4392,N_4186);
or U5112 (N_5112,N_4016,N_4779);
or U5113 (N_5113,N_4535,N_4146);
nand U5114 (N_5114,N_4725,N_4978);
xnor U5115 (N_5115,N_4634,N_4249);
xnor U5116 (N_5116,N_4680,N_4033);
and U5117 (N_5117,N_4386,N_4555);
nor U5118 (N_5118,N_4739,N_4470);
and U5119 (N_5119,N_4302,N_4159);
or U5120 (N_5120,N_4445,N_4619);
xor U5121 (N_5121,N_4252,N_4142);
and U5122 (N_5122,N_4495,N_4775);
or U5123 (N_5123,N_4163,N_4787);
and U5124 (N_5124,N_4350,N_4639);
and U5125 (N_5125,N_4584,N_4439);
nand U5126 (N_5126,N_4932,N_4181);
nor U5127 (N_5127,N_4782,N_4860);
or U5128 (N_5128,N_4246,N_4140);
nor U5129 (N_5129,N_4988,N_4816);
nor U5130 (N_5130,N_4313,N_4032);
xor U5131 (N_5131,N_4047,N_4883);
xnor U5132 (N_5132,N_4156,N_4865);
and U5133 (N_5133,N_4679,N_4574);
xor U5134 (N_5134,N_4478,N_4952);
and U5135 (N_5135,N_4373,N_4214);
and U5136 (N_5136,N_4384,N_4209);
nand U5137 (N_5137,N_4013,N_4606);
and U5138 (N_5138,N_4514,N_4127);
nand U5139 (N_5139,N_4525,N_4633);
xor U5140 (N_5140,N_4537,N_4710);
nand U5141 (N_5141,N_4309,N_4280);
xor U5142 (N_5142,N_4592,N_4659);
xnor U5143 (N_5143,N_4721,N_4221);
and U5144 (N_5144,N_4176,N_4287);
xnor U5145 (N_5145,N_4101,N_4056);
and U5146 (N_5146,N_4505,N_4261);
and U5147 (N_5147,N_4896,N_4812);
nand U5148 (N_5148,N_4691,N_4232);
or U5149 (N_5149,N_4065,N_4224);
xnor U5150 (N_5150,N_4123,N_4849);
xor U5151 (N_5151,N_4587,N_4198);
nand U5152 (N_5152,N_4638,N_4270);
xnor U5153 (N_5153,N_4536,N_4388);
and U5154 (N_5154,N_4121,N_4380);
and U5155 (N_5155,N_4391,N_4042);
nor U5156 (N_5156,N_4300,N_4964);
xor U5157 (N_5157,N_4279,N_4712);
nand U5158 (N_5158,N_4903,N_4152);
or U5159 (N_5159,N_4599,N_4912);
nand U5160 (N_5160,N_4858,N_4778);
xor U5161 (N_5161,N_4856,N_4566);
and U5162 (N_5162,N_4967,N_4172);
nor U5163 (N_5163,N_4149,N_4830);
and U5164 (N_5164,N_4624,N_4550);
or U5165 (N_5165,N_4502,N_4239);
nand U5166 (N_5166,N_4894,N_4483);
xor U5167 (N_5167,N_4414,N_4342);
and U5168 (N_5168,N_4053,N_4137);
nand U5169 (N_5169,N_4991,N_4735);
xnor U5170 (N_5170,N_4757,N_4087);
xor U5171 (N_5171,N_4885,N_4133);
and U5172 (N_5172,N_4393,N_4676);
nand U5173 (N_5173,N_4568,N_4969);
or U5174 (N_5174,N_4098,N_4752);
nor U5175 (N_5175,N_4534,N_4644);
or U5176 (N_5176,N_4167,N_4909);
nor U5177 (N_5177,N_4262,N_4441);
and U5178 (N_5178,N_4651,N_4933);
nor U5179 (N_5179,N_4452,N_4283);
nor U5180 (N_5180,N_4456,N_4880);
or U5181 (N_5181,N_4026,N_4955);
nor U5182 (N_5182,N_4871,N_4916);
or U5183 (N_5183,N_4075,N_4717);
nor U5184 (N_5184,N_4268,N_4070);
xor U5185 (N_5185,N_4637,N_4227);
or U5186 (N_5186,N_4009,N_4815);
nor U5187 (N_5187,N_4358,N_4448);
nand U5188 (N_5188,N_4260,N_4323);
nor U5189 (N_5189,N_4253,N_4876);
nor U5190 (N_5190,N_4203,N_4213);
and U5191 (N_5191,N_4990,N_4950);
xnor U5192 (N_5192,N_4361,N_4458);
xnor U5193 (N_5193,N_4987,N_4714);
xor U5194 (N_5194,N_4022,N_4118);
nand U5195 (N_5195,N_4832,N_4202);
nand U5196 (N_5196,N_4306,N_4546);
xnor U5197 (N_5197,N_4374,N_4336);
nor U5198 (N_5198,N_4104,N_4357);
xor U5199 (N_5199,N_4804,N_4959);
xor U5200 (N_5200,N_4077,N_4389);
nand U5201 (N_5201,N_4332,N_4036);
xnor U5202 (N_5202,N_4503,N_4963);
xnor U5203 (N_5203,N_4124,N_4652);
or U5204 (N_5204,N_4906,N_4835);
or U5205 (N_5205,N_4947,N_4851);
xor U5206 (N_5206,N_4755,N_4926);
and U5207 (N_5207,N_4316,N_4084);
nand U5208 (N_5208,N_4837,N_4212);
or U5209 (N_5209,N_4489,N_4387);
and U5210 (N_5210,N_4884,N_4041);
nand U5211 (N_5211,N_4248,N_4229);
nor U5212 (N_5212,N_4451,N_4063);
nor U5213 (N_5213,N_4881,N_4827);
and U5214 (N_5214,N_4591,N_4288);
nor U5215 (N_5215,N_4711,N_4431);
and U5216 (N_5216,N_4877,N_4512);
and U5217 (N_5217,N_4972,N_4303);
nor U5218 (N_5218,N_4946,N_4898);
or U5219 (N_5219,N_4317,N_4833);
xor U5220 (N_5220,N_4225,N_4376);
or U5221 (N_5221,N_4277,N_4836);
xor U5222 (N_5222,N_4184,N_4061);
and U5223 (N_5223,N_4291,N_4626);
nand U5224 (N_5224,N_4750,N_4531);
or U5225 (N_5225,N_4264,N_4975);
or U5226 (N_5226,N_4980,N_4683);
xor U5227 (N_5227,N_4905,N_4853);
nand U5228 (N_5228,N_4868,N_4554);
nor U5229 (N_5229,N_4500,N_4620);
and U5230 (N_5230,N_4708,N_4675);
xnor U5231 (N_5231,N_4193,N_4071);
nand U5232 (N_5232,N_4893,N_4048);
nand U5233 (N_5233,N_4293,N_4718);
nand U5234 (N_5234,N_4299,N_4355);
or U5235 (N_5235,N_4919,N_4760);
nand U5236 (N_5236,N_4890,N_4577);
or U5237 (N_5237,N_4597,N_4083);
nand U5238 (N_5238,N_4069,N_4974);
or U5239 (N_5239,N_4351,N_4155);
nand U5240 (N_5240,N_4621,N_4789);
nor U5241 (N_5241,N_4737,N_4131);
or U5242 (N_5242,N_4492,N_4873);
nor U5243 (N_5243,N_4162,N_4608);
nor U5244 (N_5244,N_4786,N_4119);
and U5245 (N_5245,N_4002,N_4234);
nand U5246 (N_5246,N_4716,N_4818);
and U5247 (N_5247,N_4437,N_4821);
xnor U5248 (N_5248,N_4366,N_4499);
and U5249 (N_5249,N_4192,N_4031);
or U5250 (N_5250,N_4586,N_4687);
nor U5251 (N_5251,N_4995,N_4682);
xor U5252 (N_5252,N_4180,N_4204);
nor U5253 (N_5253,N_4243,N_4265);
or U5254 (N_5254,N_4962,N_4039);
and U5255 (N_5255,N_4024,N_4829);
or U5256 (N_5256,N_4774,N_4017);
xor U5257 (N_5257,N_4160,N_4862);
xor U5258 (N_5258,N_4109,N_4681);
xnor U5259 (N_5259,N_4631,N_4436);
nand U5260 (N_5260,N_4328,N_4530);
xnor U5261 (N_5261,N_4296,N_4562);
nand U5262 (N_5262,N_4169,N_4540);
nand U5263 (N_5263,N_4614,N_4136);
nor U5264 (N_5264,N_4612,N_4258);
nand U5265 (N_5265,N_4748,N_4095);
nor U5266 (N_5266,N_4917,N_4401);
and U5267 (N_5267,N_4082,N_4648);
nor U5268 (N_5268,N_4370,N_4326);
nor U5269 (N_5269,N_4197,N_4971);
or U5270 (N_5270,N_4257,N_4308);
nor U5271 (N_5271,N_4770,N_4549);
nor U5272 (N_5272,N_4780,N_4785);
and U5273 (N_5273,N_4669,N_4471);
nand U5274 (N_5274,N_4240,N_4922);
nor U5275 (N_5275,N_4960,N_4741);
xor U5276 (N_5276,N_4333,N_4122);
and U5277 (N_5277,N_4986,N_4573);
xnor U5278 (N_5278,N_4810,N_4403);
nand U5279 (N_5279,N_4730,N_4433);
and U5280 (N_5280,N_4272,N_4430);
nor U5281 (N_5281,N_4230,N_4914);
xor U5282 (N_5282,N_4699,N_4426);
nand U5283 (N_5283,N_4236,N_4315);
xor U5284 (N_5284,N_4511,N_4520);
nor U5285 (N_5285,N_4889,N_4524);
or U5286 (N_5286,N_4551,N_4820);
or U5287 (N_5287,N_4529,N_4211);
xnor U5288 (N_5288,N_4020,N_4940);
xnor U5289 (N_5289,N_4622,N_4266);
and U5290 (N_5290,N_4761,N_4319);
or U5291 (N_5291,N_4968,N_4245);
or U5292 (N_5292,N_4625,N_4556);
and U5293 (N_5293,N_4544,N_4200);
nand U5294 (N_5294,N_4058,N_4989);
nor U5295 (N_5295,N_4589,N_4754);
nor U5296 (N_5296,N_4874,N_4707);
or U5297 (N_5297,N_4294,N_4698);
and U5298 (N_5298,N_4521,N_4477);
and U5299 (N_5299,N_4465,N_4353);
xor U5300 (N_5300,N_4055,N_4286);
and U5301 (N_5301,N_4934,N_4408);
nand U5302 (N_5302,N_4751,N_4595);
or U5303 (N_5303,N_4814,N_4290);
and U5304 (N_5304,N_4931,N_4692);
or U5305 (N_5305,N_4765,N_4125);
and U5306 (N_5306,N_4143,N_4208);
and U5307 (N_5307,N_4417,N_4004);
and U5308 (N_5308,N_4066,N_4879);
and U5309 (N_5309,N_4216,N_4665);
or U5310 (N_5310,N_4498,N_4560);
and U5311 (N_5311,N_4985,N_4640);
and U5312 (N_5312,N_4977,N_4583);
xor U5313 (N_5313,N_4443,N_4942);
and U5314 (N_5314,N_4642,N_4994);
and U5315 (N_5315,N_4628,N_4539);
and U5316 (N_5316,N_4515,N_4444);
nor U5317 (N_5317,N_4742,N_4311);
nor U5318 (N_5318,N_4559,N_4590);
or U5319 (N_5319,N_4738,N_4702);
and U5320 (N_5320,N_4107,N_4689);
or U5321 (N_5321,N_4359,N_4429);
or U5322 (N_5322,N_4557,N_4784);
nand U5323 (N_5323,N_4057,N_4196);
nand U5324 (N_5324,N_4870,N_4468);
and U5325 (N_5325,N_4709,N_4649);
nand U5326 (N_5326,N_4144,N_4105);
nor U5327 (N_5327,N_4364,N_4510);
and U5328 (N_5328,N_4930,N_4727);
or U5329 (N_5329,N_4791,N_4844);
or U5330 (N_5330,N_4610,N_4096);
nor U5331 (N_5331,N_4961,N_4504);
and U5332 (N_5332,N_4979,N_4949);
xor U5333 (N_5333,N_4464,N_4073);
nand U5334 (N_5334,N_4434,N_4891);
nand U5335 (N_5335,N_4892,N_4713);
nand U5336 (N_5336,N_4719,N_4183);
xor U5337 (N_5337,N_4668,N_4522);
xor U5338 (N_5338,N_4601,N_4532);
and U5339 (N_5339,N_4404,N_4607);
or U5340 (N_5340,N_4759,N_4375);
or U5341 (N_5341,N_4076,N_4796);
or U5342 (N_5342,N_4729,N_4630);
nand U5343 (N_5343,N_4195,N_4686);
nor U5344 (N_5344,N_4207,N_4957);
xnor U5345 (N_5345,N_4915,N_4795);
nand U5346 (N_5346,N_4348,N_4377);
nand U5347 (N_5347,N_4278,N_4054);
and U5348 (N_5348,N_4611,N_4341);
nand U5349 (N_5349,N_4330,N_4747);
nand U5350 (N_5350,N_4263,N_4019);
nor U5351 (N_5351,N_4190,N_4298);
or U5352 (N_5352,N_4720,N_4372);
nor U5353 (N_5353,N_4838,N_4485);
xnor U5354 (N_5354,N_4218,N_4324);
and U5355 (N_5355,N_4001,N_4732);
and U5356 (N_5356,N_4199,N_4882);
xor U5357 (N_5357,N_4354,N_4693);
xor U5358 (N_5358,N_4673,N_4201);
xor U5359 (N_5359,N_4809,N_4847);
and U5360 (N_5360,N_4623,N_4396);
nand U5361 (N_5361,N_4074,N_4297);
nand U5362 (N_5362,N_4356,N_4846);
nand U5363 (N_5363,N_4139,N_4480);
nor U5364 (N_5364,N_4670,N_4023);
nor U5365 (N_5365,N_4533,N_4340);
and U5366 (N_5366,N_4839,N_4613);
nand U5367 (N_5367,N_4043,N_4412);
xor U5368 (N_5368,N_4025,N_4153);
xnor U5369 (N_5369,N_4362,N_4331);
nor U5370 (N_5370,N_4226,N_4811);
nand U5371 (N_5371,N_4929,N_4397);
or U5372 (N_5372,N_4334,N_4185);
and U5373 (N_5373,N_4831,N_4805);
nand U5374 (N_5374,N_4453,N_4723);
and U5375 (N_5375,N_4344,N_4825);
or U5376 (N_5376,N_4325,N_4244);
xor U5377 (N_5377,N_4841,N_4605);
and U5378 (N_5378,N_4888,N_4457);
xor U5379 (N_5379,N_4166,N_4440);
xor U5380 (N_5380,N_4079,N_4416);
nor U5381 (N_5381,N_4895,N_4598);
nand U5382 (N_5382,N_4921,N_4329);
nand U5383 (N_5383,N_4428,N_4935);
or U5384 (N_5384,N_4878,N_4147);
and U5385 (N_5385,N_4970,N_4616);
nand U5386 (N_5386,N_4704,N_4233);
nand U5387 (N_5387,N_4722,N_4661);
xor U5388 (N_5388,N_4187,N_4134);
nor U5389 (N_5389,N_4085,N_4129);
nor U5390 (N_5390,N_4864,N_4688);
and U5391 (N_5391,N_4734,N_4663);
xnor U5392 (N_5392,N_4756,N_4567);
and U5393 (N_5393,N_4466,N_4766);
or U5394 (N_5394,N_4106,N_4217);
and U5395 (N_5395,N_4854,N_4335);
nor U5396 (N_5396,N_4936,N_4337);
xnor U5397 (N_5397,N_4694,N_4210);
nor U5398 (N_5398,N_4768,N_4273);
nor U5399 (N_5399,N_4455,N_4824);
nand U5400 (N_5400,N_4314,N_4788);
or U5401 (N_5401,N_4007,N_4564);
xor U5402 (N_5402,N_4062,N_4449);
nand U5403 (N_5403,N_4424,N_4128);
nor U5404 (N_5404,N_4951,N_4845);
or U5405 (N_5405,N_4493,N_4275);
or U5406 (N_5406,N_4132,N_4801);
nand U5407 (N_5407,N_4646,N_4292);
nand U5408 (N_5408,N_4117,N_4479);
or U5409 (N_5409,N_4363,N_4223);
nor U5410 (N_5410,N_4897,N_4154);
and U5411 (N_5411,N_4571,N_4565);
nor U5412 (N_5412,N_4467,N_4100);
or U5413 (N_5413,N_4938,N_4454);
or U5414 (N_5414,N_4219,N_4904);
and U5415 (N_5415,N_4378,N_4650);
nor U5416 (N_5416,N_4170,N_4138);
xnor U5417 (N_5417,N_4516,N_4899);
nand U5418 (N_5418,N_4060,N_4802);
nor U5419 (N_5419,N_4182,N_4736);
or U5420 (N_5420,N_4000,N_4604);
and U5421 (N_5421,N_4706,N_4910);
nand U5422 (N_5422,N_4561,N_4052);
or U5423 (N_5423,N_4743,N_4369);
or U5424 (N_5424,N_4998,N_4494);
xor U5425 (N_5425,N_4114,N_4027);
and U5426 (N_5426,N_4834,N_4438);
xnor U5427 (N_5427,N_4112,N_4011);
or U5428 (N_5428,N_4697,N_4655);
nand U5429 (N_5429,N_4749,N_4255);
nand U5430 (N_5430,N_4501,N_4705);
and U5431 (N_5431,N_4783,N_4852);
nor U5432 (N_5432,N_4753,N_4365);
xor U5433 (N_5433,N_4842,N_4284);
nor U5434 (N_5434,N_4126,N_4158);
and U5435 (N_5435,N_4850,N_4318);
xor U5436 (N_5436,N_4442,N_4091);
nand U5437 (N_5437,N_4450,N_4006);
or U5438 (N_5438,N_4281,N_4684);
or U5439 (N_5439,N_4828,N_4635);
nor U5440 (N_5440,N_4777,N_4411);
nand U5441 (N_5441,N_4983,N_4282);
nor U5442 (N_5442,N_4523,N_4228);
xor U5443 (N_5443,N_4602,N_4345);
xor U5444 (N_5444,N_4409,N_4432);
nor U5445 (N_5445,N_4800,N_4177);
nor U5446 (N_5446,N_4321,N_4875);
and U5447 (N_5447,N_4044,N_4907);
and U5448 (N_5448,N_4194,N_4157);
and U5449 (N_5449,N_4701,N_4672);
xor U5450 (N_5450,N_4807,N_4953);
xnor U5451 (N_5451,N_4307,N_4745);
nand U5452 (N_5452,N_4237,N_4446);
xor U5453 (N_5453,N_4615,N_4769);
xor U5454 (N_5454,N_4617,N_4855);
and U5455 (N_5455,N_4762,N_4993);
and U5456 (N_5456,N_4289,N_4944);
xor U5457 (N_5457,N_4799,N_4148);
nor U5458 (N_5458,N_4588,N_4113);
or U5459 (N_5459,N_4526,N_4171);
nand U5460 (N_5460,N_4744,N_4861);
and U5461 (N_5461,N_4886,N_4872);
nor U5462 (N_5462,N_4476,N_4420);
or U5463 (N_5463,N_4817,N_4090);
nor U5464 (N_5464,N_4343,N_4996);
xnor U5465 (N_5465,N_4596,N_4660);
xor U5466 (N_5466,N_4593,N_4773);
nor U5467 (N_5467,N_4474,N_4920);
and U5468 (N_5468,N_4086,N_4482);
or U5469 (N_5469,N_4089,N_4014);
xor U5470 (N_5470,N_4901,N_4305);
nand U5471 (N_5471,N_4654,N_4220);
xnor U5472 (N_5472,N_4618,N_4740);
nand U5473 (N_5473,N_4627,N_4472);
xor U5474 (N_5474,N_4580,N_4368);
or U5475 (N_5475,N_4927,N_4999);
and U5476 (N_5476,N_4965,N_4347);
xnor U5477 (N_5477,N_4141,N_4463);
and U5478 (N_5478,N_4304,N_4092);
or U5479 (N_5479,N_4150,N_4793);
and U5480 (N_5480,N_4352,N_4179);
nor U5481 (N_5481,N_4269,N_4671);
nand U5482 (N_5482,N_4285,N_4080);
nand U5483 (N_5483,N_4320,N_4346);
nor U5484 (N_5484,N_4059,N_4003);
nor U5485 (N_5485,N_4813,N_4110);
and U5486 (N_5486,N_4338,N_4413);
or U5487 (N_5487,N_4662,N_4274);
or U5488 (N_5488,N_4473,N_4859);
nand U5489 (N_5489,N_4469,N_4360);
and U5490 (N_5490,N_4518,N_4600);
xnor U5491 (N_5491,N_4819,N_4254);
and U5492 (N_5492,N_4383,N_4312);
or U5493 (N_5493,N_4046,N_4486);
and U5494 (N_5494,N_4447,N_4576);
xor U5495 (N_5495,N_4406,N_4402);
nand U5496 (N_5496,N_4506,N_4746);
xor U5497 (N_5497,N_4728,N_4781);
nand U5498 (N_5498,N_4956,N_4135);
nand U5499 (N_5499,N_4400,N_4423);
or U5500 (N_5500,N_4527,N_4580);
and U5501 (N_5501,N_4153,N_4678);
nand U5502 (N_5502,N_4707,N_4733);
xnor U5503 (N_5503,N_4420,N_4705);
xnor U5504 (N_5504,N_4145,N_4345);
nor U5505 (N_5505,N_4467,N_4407);
or U5506 (N_5506,N_4597,N_4577);
nand U5507 (N_5507,N_4120,N_4858);
and U5508 (N_5508,N_4119,N_4744);
nand U5509 (N_5509,N_4599,N_4161);
and U5510 (N_5510,N_4633,N_4552);
nand U5511 (N_5511,N_4767,N_4116);
and U5512 (N_5512,N_4192,N_4224);
nor U5513 (N_5513,N_4153,N_4050);
nor U5514 (N_5514,N_4261,N_4210);
nor U5515 (N_5515,N_4803,N_4628);
and U5516 (N_5516,N_4675,N_4736);
nand U5517 (N_5517,N_4033,N_4930);
or U5518 (N_5518,N_4930,N_4711);
nor U5519 (N_5519,N_4291,N_4016);
xor U5520 (N_5520,N_4479,N_4208);
nor U5521 (N_5521,N_4733,N_4892);
nor U5522 (N_5522,N_4402,N_4271);
or U5523 (N_5523,N_4692,N_4734);
nand U5524 (N_5524,N_4976,N_4628);
nor U5525 (N_5525,N_4574,N_4666);
or U5526 (N_5526,N_4923,N_4472);
or U5527 (N_5527,N_4788,N_4537);
nand U5528 (N_5528,N_4007,N_4846);
or U5529 (N_5529,N_4078,N_4280);
nand U5530 (N_5530,N_4846,N_4720);
nand U5531 (N_5531,N_4523,N_4703);
nor U5532 (N_5532,N_4753,N_4300);
xnor U5533 (N_5533,N_4052,N_4275);
nand U5534 (N_5534,N_4986,N_4305);
nand U5535 (N_5535,N_4334,N_4295);
nand U5536 (N_5536,N_4268,N_4492);
nor U5537 (N_5537,N_4749,N_4248);
xnor U5538 (N_5538,N_4495,N_4940);
and U5539 (N_5539,N_4518,N_4482);
xor U5540 (N_5540,N_4443,N_4811);
xor U5541 (N_5541,N_4753,N_4170);
nand U5542 (N_5542,N_4844,N_4287);
nor U5543 (N_5543,N_4591,N_4458);
nor U5544 (N_5544,N_4527,N_4160);
nand U5545 (N_5545,N_4145,N_4835);
nand U5546 (N_5546,N_4534,N_4688);
xnor U5547 (N_5547,N_4730,N_4209);
nor U5548 (N_5548,N_4681,N_4560);
and U5549 (N_5549,N_4754,N_4762);
xor U5550 (N_5550,N_4656,N_4128);
and U5551 (N_5551,N_4316,N_4264);
nor U5552 (N_5552,N_4771,N_4809);
nand U5553 (N_5553,N_4610,N_4938);
xnor U5554 (N_5554,N_4148,N_4635);
nor U5555 (N_5555,N_4473,N_4890);
nor U5556 (N_5556,N_4691,N_4548);
xnor U5557 (N_5557,N_4340,N_4113);
xor U5558 (N_5558,N_4184,N_4264);
nand U5559 (N_5559,N_4187,N_4570);
and U5560 (N_5560,N_4446,N_4637);
or U5561 (N_5561,N_4485,N_4391);
or U5562 (N_5562,N_4290,N_4261);
nand U5563 (N_5563,N_4374,N_4100);
nor U5564 (N_5564,N_4471,N_4495);
nand U5565 (N_5565,N_4748,N_4463);
and U5566 (N_5566,N_4302,N_4280);
nand U5567 (N_5567,N_4489,N_4055);
and U5568 (N_5568,N_4518,N_4575);
nor U5569 (N_5569,N_4761,N_4759);
xnor U5570 (N_5570,N_4351,N_4147);
nand U5571 (N_5571,N_4412,N_4696);
xnor U5572 (N_5572,N_4497,N_4468);
nor U5573 (N_5573,N_4501,N_4844);
or U5574 (N_5574,N_4459,N_4602);
xor U5575 (N_5575,N_4989,N_4565);
and U5576 (N_5576,N_4800,N_4978);
nor U5577 (N_5577,N_4060,N_4864);
xnor U5578 (N_5578,N_4544,N_4188);
or U5579 (N_5579,N_4230,N_4674);
xnor U5580 (N_5580,N_4816,N_4020);
nor U5581 (N_5581,N_4726,N_4381);
or U5582 (N_5582,N_4725,N_4399);
or U5583 (N_5583,N_4508,N_4840);
and U5584 (N_5584,N_4263,N_4129);
xnor U5585 (N_5585,N_4385,N_4001);
and U5586 (N_5586,N_4620,N_4793);
nand U5587 (N_5587,N_4224,N_4477);
xor U5588 (N_5588,N_4770,N_4662);
xnor U5589 (N_5589,N_4283,N_4537);
and U5590 (N_5590,N_4835,N_4261);
and U5591 (N_5591,N_4407,N_4843);
and U5592 (N_5592,N_4816,N_4701);
nor U5593 (N_5593,N_4803,N_4524);
xor U5594 (N_5594,N_4336,N_4684);
or U5595 (N_5595,N_4983,N_4962);
nor U5596 (N_5596,N_4103,N_4042);
or U5597 (N_5597,N_4308,N_4446);
nand U5598 (N_5598,N_4814,N_4477);
nor U5599 (N_5599,N_4730,N_4892);
nor U5600 (N_5600,N_4766,N_4674);
nor U5601 (N_5601,N_4210,N_4368);
xor U5602 (N_5602,N_4915,N_4639);
or U5603 (N_5603,N_4297,N_4162);
nand U5604 (N_5604,N_4121,N_4045);
nand U5605 (N_5605,N_4636,N_4458);
xor U5606 (N_5606,N_4464,N_4181);
nand U5607 (N_5607,N_4822,N_4847);
nand U5608 (N_5608,N_4579,N_4129);
or U5609 (N_5609,N_4268,N_4520);
nor U5610 (N_5610,N_4226,N_4003);
nor U5611 (N_5611,N_4287,N_4668);
nor U5612 (N_5612,N_4800,N_4780);
or U5613 (N_5613,N_4241,N_4422);
nor U5614 (N_5614,N_4194,N_4215);
nor U5615 (N_5615,N_4957,N_4744);
nor U5616 (N_5616,N_4107,N_4940);
nand U5617 (N_5617,N_4327,N_4068);
nand U5618 (N_5618,N_4811,N_4145);
nand U5619 (N_5619,N_4463,N_4867);
or U5620 (N_5620,N_4412,N_4238);
or U5621 (N_5621,N_4101,N_4876);
or U5622 (N_5622,N_4283,N_4688);
nor U5623 (N_5623,N_4727,N_4810);
or U5624 (N_5624,N_4900,N_4387);
nor U5625 (N_5625,N_4121,N_4177);
or U5626 (N_5626,N_4528,N_4909);
and U5627 (N_5627,N_4369,N_4459);
or U5628 (N_5628,N_4288,N_4628);
and U5629 (N_5629,N_4559,N_4278);
or U5630 (N_5630,N_4978,N_4103);
and U5631 (N_5631,N_4630,N_4733);
or U5632 (N_5632,N_4494,N_4546);
nor U5633 (N_5633,N_4943,N_4760);
nor U5634 (N_5634,N_4222,N_4859);
nand U5635 (N_5635,N_4745,N_4108);
and U5636 (N_5636,N_4072,N_4127);
nor U5637 (N_5637,N_4091,N_4073);
nor U5638 (N_5638,N_4142,N_4106);
or U5639 (N_5639,N_4152,N_4257);
and U5640 (N_5640,N_4739,N_4826);
and U5641 (N_5641,N_4074,N_4274);
or U5642 (N_5642,N_4397,N_4651);
or U5643 (N_5643,N_4105,N_4441);
xor U5644 (N_5644,N_4602,N_4618);
and U5645 (N_5645,N_4989,N_4103);
or U5646 (N_5646,N_4907,N_4683);
or U5647 (N_5647,N_4798,N_4005);
nor U5648 (N_5648,N_4586,N_4164);
nand U5649 (N_5649,N_4839,N_4243);
or U5650 (N_5650,N_4046,N_4849);
xor U5651 (N_5651,N_4431,N_4969);
nand U5652 (N_5652,N_4866,N_4513);
nor U5653 (N_5653,N_4390,N_4009);
nor U5654 (N_5654,N_4626,N_4878);
nor U5655 (N_5655,N_4177,N_4384);
and U5656 (N_5656,N_4321,N_4157);
nor U5657 (N_5657,N_4268,N_4255);
and U5658 (N_5658,N_4879,N_4109);
nor U5659 (N_5659,N_4706,N_4211);
or U5660 (N_5660,N_4524,N_4689);
nand U5661 (N_5661,N_4996,N_4158);
nor U5662 (N_5662,N_4970,N_4749);
and U5663 (N_5663,N_4971,N_4190);
or U5664 (N_5664,N_4211,N_4025);
xnor U5665 (N_5665,N_4961,N_4845);
nor U5666 (N_5666,N_4156,N_4253);
and U5667 (N_5667,N_4890,N_4503);
xnor U5668 (N_5668,N_4999,N_4090);
nand U5669 (N_5669,N_4544,N_4779);
xor U5670 (N_5670,N_4907,N_4716);
nand U5671 (N_5671,N_4093,N_4684);
or U5672 (N_5672,N_4618,N_4563);
xor U5673 (N_5673,N_4312,N_4765);
or U5674 (N_5674,N_4528,N_4413);
or U5675 (N_5675,N_4255,N_4320);
and U5676 (N_5676,N_4986,N_4577);
or U5677 (N_5677,N_4611,N_4972);
and U5678 (N_5678,N_4774,N_4877);
nor U5679 (N_5679,N_4753,N_4808);
nand U5680 (N_5680,N_4340,N_4606);
xor U5681 (N_5681,N_4611,N_4404);
nand U5682 (N_5682,N_4000,N_4417);
nor U5683 (N_5683,N_4891,N_4946);
or U5684 (N_5684,N_4917,N_4997);
and U5685 (N_5685,N_4227,N_4246);
nor U5686 (N_5686,N_4386,N_4301);
or U5687 (N_5687,N_4777,N_4221);
xnor U5688 (N_5688,N_4987,N_4190);
or U5689 (N_5689,N_4903,N_4808);
and U5690 (N_5690,N_4772,N_4381);
and U5691 (N_5691,N_4115,N_4862);
xor U5692 (N_5692,N_4517,N_4109);
nand U5693 (N_5693,N_4014,N_4815);
nor U5694 (N_5694,N_4559,N_4732);
xor U5695 (N_5695,N_4399,N_4599);
or U5696 (N_5696,N_4977,N_4185);
and U5697 (N_5697,N_4935,N_4838);
or U5698 (N_5698,N_4117,N_4470);
xor U5699 (N_5699,N_4728,N_4151);
xor U5700 (N_5700,N_4339,N_4523);
nand U5701 (N_5701,N_4244,N_4820);
or U5702 (N_5702,N_4961,N_4214);
and U5703 (N_5703,N_4314,N_4592);
nand U5704 (N_5704,N_4563,N_4419);
and U5705 (N_5705,N_4248,N_4404);
nand U5706 (N_5706,N_4405,N_4603);
nor U5707 (N_5707,N_4497,N_4452);
and U5708 (N_5708,N_4534,N_4248);
nand U5709 (N_5709,N_4458,N_4622);
nor U5710 (N_5710,N_4447,N_4085);
xor U5711 (N_5711,N_4868,N_4701);
nor U5712 (N_5712,N_4775,N_4038);
nor U5713 (N_5713,N_4047,N_4080);
and U5714 (N_5714,N_4378,N_4047);
nand U5715 (N_5715,N_4128,N_4905);
or U5716 (N_5716,N_4959,N_4941);
nand U5717 (N_5717,N_4170,N_4858);
and U5718 (N_5718,N_4192,N_4713);
or U5719 (N_5719,N_4125,N_4880);
or U5720 (N_5720,N_4871,N_4307);
nand U5721 (N_5721,N_4894,N_4917);
nand U5722 (N_5722,N_4364,N_4012);
nor U5723 (N_5723,N_4598,N_4216);
nand U5724 (N_5724,N_4151,N_4233);
nor U5725 (N_5725,N_4562,N_4704);
nand U5726 (N_5726,N_4832,N_4633);
nand U5727 (N_5727,N_4350,N_4758);
or U5728 (N_5728,N_4351,N_4774);
or U5729 (N_5729,N_4332,N_4722);
and U5730 (N_5730,N_4234,N_4570);
or U5731 (N_5731,N_4563,N_4437);
xor U5732 (N_5732,N_4609,N_4441);
nor U5733 (N_5733,N_4094,N_4361);
xnor U5734 (N_5734,N_4273,N_4791);
or U5735 (N_5735,N_4014,N_4672);
or U5736 (N_5736,N_4555,N_4406);
and U5737 (N_5737,N_4580,N_4831);
nand U5738 (N_5738,N_4457,N_4772);
or U5739 (N_5739,N_4693,N_4653);
nor U5740 (N_5740,N_4937,N_4583);
xor U5741 (N_5741,N_4431,N_4317);
xor U5742 (N_5742,N_4567,N_4354);
xor U5743 (N_5743,N_4238,N_4386);
or U5744 (N_5744,N_4953,N_4577);
xnor U5745 (N_5745,N_4493,N_4203);
nand U5746 (N_5746,N_4980,N_4772);
nand U5747 (N_5747,N_4421,N_4842);
nand U5748 (N_5748,N_4457,N_4721);
or U5749 (N_5749,N_4955,N_4495);
nor U5750 (N_5750,N_4109,N_4714);
nand U5751 (N_5751,N_4572,N_4857);
nor U5752 (N_5752,N_4237,N_4007);
or U5753 (N_5753,N_4454,N_4263);
xor U5754 (N_5754,N_4816,N_4441);
nand U5755 (N_5755,N_4886,N_4929);
and U5756 (N_5756,N_4265,N_4919);
xor U5757 (N_5757,N_4635,N_4652);
and U5758 (N_5758,N_4245,N_4849);
nor U5759 (N_5759,N_4471,N_4026);
and U5760 (N_5760,N_4920,N_4293);
nor U5761 (N_5761,N_4778,N_4139);
nor U5762 (N_5762,N_4598,N_4870);
or U5763 (N_5763,N_4506,N_4689);
or U5764 (N_5764,N_4065,N_4714);
xnor U5765 (N_5765,N_4698,N_4624);
nor U5766 (N_5766,N_4457,N_4087);
xnor U5767 (N_5767,N_4730,N_4422);
or U5768 (N_5768,N_4729,N_4740);
nand U5769 (N_5769,N_4871,N_4189);
or U5770 (N_5770,N_4674,N_4139);
or U5771 (N_5771,N_4848,N_4440);
xor U5772 (N_5772,N_4749,N_4516);
nor U5773 (N_5773,N_4822,N_4699);
xor U5774 (N_5774,N_4836,N_4373);
or U5775 (N_5775,N_4422,N_4988);
and U5776 (N_5776,N_4061,N_4867);
nand U5777 (N_5777,N_4491,N_4009);
nand U5778 (N_5778,N_4013,N_4263);
or U5779 (N_5779,N_4687,N_4477);
xor U5780 (N_5780,N_4167,N_4155);
xor U5781 (N_5781,N_4883,N_4222);
nand U5782 (N_5782,N_4951,N_4196);
nor U5783 (N_5783,N_4356,N_4226);
or U5784 (N_5784,N_4385,N_4027);
nand U5785 (N_5785,N_4169,N_4166);
xnor U5786 (N_5786,N_4924,N_4218);
xor U5787 (N_5787,N_4483,N_4775);
and U5788 (N_5788,N_4514,N_4989);
or U5789 (N_5789,N_4798,N_4808);
and U5790 (N_5790,N_4716,N_4821);
and U5791 (N_5791,N_4613,N_4056);
xor U5792 (N_5792,N_4809,N_4823);
and U5793 (N_5793,N_4217,N_4952);
xor U5794 (N_5794,N_4826,N_4024);
and U5795 (N_5795,N_4001,N_4410);
nor U5796 (N_5796,N_4060,N_4433);
and U5797 (N_5797,N_4985,N_4432);
xor U5798 (N_5798,N_4025,N_4689);
and U5799 (N_5799,N_4631,N_4408);
or U5800 (N_5800,N_4014,N_4713);
nand U5801 (N_5801,N_4396,N_4683);
or U5802 (N_5802,N_4783,N_4990);
nand U5803 (N_5803,N_4804,N_4100);
nand U5804 (N_5804,N_4266,N_4410);
and U5805 (N_5805,N_4784,N_4418);
and U5806 (N_5806,N_4602,N_4530);
and U5807 (N_5807,N_4470,N_4336);
xor U5808 (N_5808,N_4810,N_4610);
or U5809 (N_5809,N_4366,N_4061);
and U5810 (N_5810,N_4783,N_4184);
nand U5811 (N_5811,N_4905,N_4612);
nand U5812 (N_5812,N_4366,N_4380);
xor U5813 (N_5813,N_4175,N_4225);
nor U5814 (N_5814,N_4949,N_4568);
and U5815 (N_5815,N_4301,N_4548);
and U5816 (N_5816,N_4855,N_4245);
xor U5817 (N_5817,N_4571,N_4337);
or U5818 (N_5818,N_4645,N_4979);
nand U5819 (N_5819,N_4195,N_4782);
or U5820 (N_5820,N_4089,N_4842);
nand U5821 (N_5821,N_4256,N_4470);
nand U5822 (N_5822,N_4385,N_4937);
or U5823 (N_5823,N_4856,N_4539);
nor U5824 (N_5824,N_4946,N_4597);
and U5825 (N_5825,N_4616,N_4385);
or U5826 (N_5826,N_4939,N_4703);
nor U5827 (N_5827,N_4710,N_4431);
nor U5828 (N_5828,N_4760,N_4882);
xor U5829 (N_5829,N_4685,N_4825);
nor U5830 (N_5830,N_4544,N_4612);
nand U5831 (N_5831,N_4313,N_4823);
and U5832 (N_5832,N_4003,N_4106);
or U5833 (N_5833,N_4357,N_4966);
and U5834 (N_5834,N_4656,N_4099);
and U5835 (N_5835,N_4177,N_4579);
xor U5836 (N_5836,N_4630,N_4778);
nor U5837 (N_5837,N_4633,N_4726);
or U5838 (N_5838,N_4000,N_4258);
and U5839 (N_5839,N_4486,N_4364);
or U5840 (N_5840,N_4535,N_4151);
nor U5841 (N_5841,N_4970,N_4820);
and U5842 (N_5842,N_4648,N_4876);
nand U5843 (N_5843,N_4372,N_4229);
and U5844 (N_5844,N_4301,N_4947);
and U5845 (N_5845,N_4803,N_4551);
xnor U5846 (N_5846,N_4663,N_4388);
nand U5847 (N_5847,N_4599,N_4059);
nand U5848 (N_5848,N_4087,N_4531);
xnor U5849 (N_5849,N_4552,N_4289);
nor U5850 (N_5850,N_4331,N_4206);
or U5851 (N_5851,N_4360,N_4219);
nand U5852 (N_5852,N_4433,N_4609);
nand U5853 (N_5853,N_4648,N_4804);
nor U5854 (N_5854,N_4184,N_4864);
and U5855 (N_5855,N_4499,N_4681);
or U5856 (N_5856,N_4844,N_4947);
nand U5857 (N_5857,N_4816,N_4044);
nand U5858 (N_5858,N_4605,N_4826);
or U5859 (N_5859,N_4997,N_4169);
xnor U5860 (N_5860,N_4142,N_4251);
xor U5861 (N_5861,N_4427,N_4950);
or U5862 (N_5862,N_4654,N_4403);
xnor U5863 (N_5863,N_4947,N_4768);
xnor U5864 (N_5864,N_4800,N_4968);
nand U5865 (N_5865,N_4314,N_4014);
nand U5866 (N_5866,N_4378,N_4019);
xor U5867 (N_5867,N_4594,N_4264);
nand U5868 (N_5868,N_4822,N_4307);
or U5869 (N_5869,N_4168,N_4315);
nand U5870 (N_5870,N_4158,N_4043);
and U5871 (N_5871,N_4457,N_4391);
or U5872 (N_5872,N_4777,N_4186);
nand U5873 (N_5873,N_4539,N_4780);
and U5874 (N_5874,N_4847,N_4482);
xor U5875 (N_5875,N_4913,N_4222);
xor U5876 (N_5876,N_4479,N_4569);
or U5877 (N_5877,N_4892,N_4066);
nor U5878 (N_5878,N_4293,N_4037);
nand U5879 (N_5879,N_4223,N_4513);
xor U5880 (N_5880,N_4548,N_4589);
or U5881 (N_5881,N_4557,N_4361);
or U5882 (N_5882,N_4071,N_4291);
xnor U5883 (N_5883,N_4579,N_4973);
nor U5884 (N_5884,N_4524,N_4044);
and U5885 (N_5885,N_4571,N_4199);
nor U5886 (N_5886,N_4252,N_4269);
nand U5887 (N_5887,N_4290,N_4706);
nand U5888 (N_5888,N_4357,N_4088);
nor U5889 (N_5889,N_4537,N_4080);
nand U5890 (N_5890,N_4400,N_4330);
nor U5891 (N_5891,N_4235,N_4419);
or U5892 (N_5892,N_4386,N_4547);
nand U5893 (N_5893,N_4097,N_4988);
nor U5894 (N_5894,N_4821,N_4958);
nand U5895 (N_5895,N_4011,N_4254);
or U5896 (N_5896,N_4332,N_4019);
and U5897 (N_5897,N_4817,N_4637);
or U5898 (N_5898,N_4257,N_4302);
and U5899 (N_5899,N_4071,N_4237);
nor U5900 (N_5900,N_4644,N_4648);
nor U5901 (N_5901,N_4439,N_4498);
and U5902 (N_5902,N_4339,N_4317);
and U5903 (N_5903,N_4162,N_4058);
nor U5904 (N_5904,N_4949,N_4533);
nand U5905 (N_5905,N_4639,N_4776);
nor U5906 (N_5906,N_4765,N_4295);
xnor U5907 (N_5907,N_4393,N_4995);
or U5908 (N_5908,N_4084,N_4394);
xnor U5909 (N_5909,N_4822,N_4667);
nor U5910 (N_5910,N_4342,N_4766);
nor U5911 (N_5911,N_4334,N_4651);
and U5912 (N_5912,N_4054,N_4414);
nand U5913 (N_5913,N_4863,N_4407);
or U5914 (N_5914,N_4159,N_4600);
nand U5915 (N_5915,N_4853,N_4858);
nand U5916 (N_5916,N_4965,N_4874);
or U5917 (N_5917,N_4720,N_4148);
xnor U5918 (N_5918,N_4328,N_4894);
xnor U5919 (N_5919,N_4227,N_4568);
or U5920 (N_5920,N_4170,N_4714);
nand U5921 (N_5921,N_4356,N_4680);
or U5922 (N_5922,N_4123,N_4081);
nor U5923 (N_5923,N_4760,N_4874);
or U5924 (N_5924,N_4890,N_4458);
and U5925 (N_5925,N_4805,N_4301);
nand U5926 (N_5926,N_4483,N_4832);
or U5927 (N_5927,N_4005,N_4914);
xor U5928 (N_5928,N_4064,N_4303);
or U5929 (N_5929,N_4443,N_4104);
nand U5930 (N_5930,N_4515,N_4926);
and U5931 (N_5931,N_4660,N_4531);
nand U5932 (N_5932,N_4563,N_4013);
nor U5933 (N_5933,N_4589,N_4005);
nor U5934 (N_5934,N_4673,N_4314);
nand U5935 (N_5935,N_4537,N_4117);
and U5936 (N_5936,N_4328,N_4532);
xnor U5937 (N_5937,N_4828,N_4830);
and U5938 (N_5938,N_4831,N_4937);
or U5939 (N_5939,N_4779,N_4231);
nand U5940 (N_5940,N_4949,N_4154);
nor U5941 (N_5941,N_4839,N_4345);
xor U5942 (N_5942,N_4905,N_4243);
nand U5943 (N_5943,N_4928,N_4797);
or U5944 (N_5944,N_4895,N_4805);
and U5945 (N_5945,N_4071,N_4088);
and U5946 (N_5946,N_4008,N_4316);
nand U5947 (N_5947,N_4680,N_4496);
or U5948 (N_5948,N_4276,N_4372);
nor U5949 (N_5949,N_4785,N_4122);
and U5950 (N_5950,N_4222,N_4852);
and U5951 (N_5951,N_4650,N_4563);
xor U5952 (N_5952,N_4604,N_4290);
or U5953 (N_5953,N_4781,N_4802);
nand U5954 (N_5954,N_4805,N_4358);
nor U5955 (N_5955,N_4164,N_4340);
or U5956 (N_5956,N_4514,N_4798);
or U5957 (N_5957,N_4671,N_4615);
nor U5958 (N_5958,N_4181,N_4305);
xnor U5959 (N_5959,N_4742,N_4825);
or U5960 (N_5960,N_4320,N_4738);
or U5961 (N_5961,N_4976,N_4267);
or U5962 (N_5962,N_4324,N_4222);
and U5963 (N_5963,N_4259,N_4227);
and U5964 (N_5964,N_4043,N_4927);
or U5965 (N_5965,N_4102,N_4185);
or U5966 (N_5966,N_4118,N_4704);
nand U5967 (N_5967,N_4903,N_4436);
nor U5968 (N_5968,N_4371,N_4134);
nor U5969 (N_5969,N_4731,N_4124);
nand U5970 (N_5970,N_4876,N_4606);
nor U5971 (N_5971,N_4712,N_4317);
xnor U5972 (N_5972,N_4411,N_4907);
or U5973 (N_5973,N_4534,N_4620);
nand U5974 (N_5974,N_4994,N_4001);
xnor U5975 (N_5975,N_4397,N_4674);
and U5976 (N_5976,N_4310,N_4762);
and U5977 (N_5977,N_4174,N_4659);
nor U5978 (N_5978,N_4941,N_4009);
nand U5979 (N_5979,N_4347,N_4684);
and U5980 (N_5980,N_4186,N_4927);
nor U5981 (N_5981,N_4808,N_4036);
and U5982 (N_5982,N_4179,N_4581);
and U5983 (N_5983,N_4543,N_4315);
xnor U5984 (N_5984,N_4634,N_4286);
or U5985 (N_5985,N_4480,N_4220);
xnor U5986 (N_5986,N_4479,N_4886);
xor U5987 (N_5987,N_4532,N_4646);
xor U5988 (N_5988,N_4146,N_4556);
and U5989 (N_5989,N_4776,N_4259);
and U5990 (N_5990,N_4818,N_4131);
nor U5991 (N_5991,N_4328,N_4247);
and U5992 (N_5992,N_4244,N_4713);
nand U5993 (N_5993,N_4329,N_4384);
or U5994 (N_5994,N_4441,N_4147);
xor U5995 (N_5995,N_4920,N_4368);
and U5996 (N_5996,N_4716,N_4623);
xor U5997 (N_5997,N_4580,N_4923);
xnor U5998 (N_5998,N_4001,N_4155);
or U5999 (N_5999,N_4002,N_4009);
nor U6000 (N_6000,N_5428,N_5232);
xor U6001 (N_6001,N_5560,N_5688);
nor U6002 (N_6002,N_5581,N_5627);
and U6003 (N_6003,N_5454,N_5360);
xor U6004 (N_6004,N_5378,N_5589);
nor U6005 (N_6005,N_5515,N_5122);
nor U6006 (N_6006,N_5608,N_5738);
nand U6007 (N_6007,N_5583,N_5200);
or U6008 (N_6008,N_5114,N_5807);
or U6009 (N_6009,N_5546,N_5486);
and U6010 (N_6010,N_5708,N_5240);
or U6011 (N_6011,N_5293,N_5464);
nand U6012 (N_6012,N_5385,N_5528);
nand U6013 (N_6013,N_5874,N_5032);
or U6014 (N_6014,N_5451,N_5535);
and U6015 (N_6015,N_5315,N_5380);
nor U6016 (N_6016,N_5747,N_5055);
or U6017 (N_6017,N_5012,N_5426);
or U6018 (N_6018,N_5376,N_5552);
nand U6019 (N_6019,N_5933,N_5333);
nand U6020 (N_6020,N_5472,N_5176);
nor U6021 (N_6021,N_5058,N_5229);
or U6022 (N_6022,N_5618,N_5906);
xnor U6023 (N_6023,N_5812,N_5703);
and U6024 (N_6024,N_5720,N_5357);
xor U6025 (N_6025,N_5201,N_5828);
nand U6026 (N_6026,N_5503,N_5001);
xor U6027 (N_6027,N_5516,N_5913);
nand U6028 (N_6028,N_5872,N_5407);
nor U6029 (N_6029,N_5649,N_5716);
and U6030 (N_6030,N_5067,N_5917);
or U6031 (N_6031,N_5047,N_5825);
and U6032 (N_6032,N_5714,N_5994);
xor U6033 (N_6033,N_5956,N_5158);
nor U6034 (N_6034,N_5118,N_5071);
xnor U6035 (N_6035,N_5383,N_5525);
nor U6036 (N_6036,N_5753,N_5263);
nor U6037 (N_6037,N_5004,N_5553);
or U6038 (N_6038,N_5039,N_5886);
xor U6039 (N_6039,N_5624,N_5659);
and U6040 (N_6040,N_5375,N_5892);
nor U6041 (N_6041,N_5041,N_5655);
nand U6042 (N_6042,N_5588,N_5558);
xor U6043 (N_6043,N_5261,N_5466);
and U6044 (N_6044,N_5936,N_5203);
nand U6045 (N_6045,N_5749,N_5813);
nand U6046 (N_6046,N_5676,N_5362);
nand U6047 (N_6047,N_5251,N_5117);
xor U6048 (N_6048,N_5142,N_5615);
nor U6049 (N_6049,N_5636,N_5606);
nor U6050 (N_6050,N_5363,N_5254);
nand U6051 (N_6051,N_5386,N_5252);
xor U6052 (N_6052,N_5264,N_5346);
and U6053 (N_6053,N_5578,N_5431);
and U6054 (N_6054,N_5074,N_5123);
nor U6055 (N_6055,N_5998,N_5083);
or U6056 (N_6056,N_5406,N_5740);
nand U6057 (N_6057,N_5392,N_5051);
nand U6058 (N_6058,N_5188,N_5015);
or U6059 (N_6059,N_5631,N_5482);
or U6060 (N_6060,N_5831,N_5793);
xor U6061 (N_6061,N_5954,N_5895);
xor U6062 (N_6062,N_5002,N_5093);
or U6063 (N_6063,N_5729,N_5511);
and U6064 (N_6064,N_5648,N_5213);
or U6065 (N_6065,N_5163,N_5672);
xor U6066 (N_6066,N_5955,N_5628);
xor U6067 (N_6067,N_5202,N_5418);
nor U6068 (N_6068,N_5169,N_5830);
nand U6069 (N_6069,N_5199,N_5322);
nor U6070 (N_6070,N_5258,N_5410);
or U6071 (N_6071,N_5524,N_5253);
or U6072 (N_6072,N_5030,N_5999);
and U6073 (N_6073,N_5846,N_5037);
xor U6074 (N_6074,N_5223,N_5265);
nand U6075 (N_6075,N_5343,N_5149);
xor U6076 (N_6076,N_5331,N_5371);
nand U6077 (N_6077,N_5962,N_5177);
or U6078 (N_6078,N_5046,N_5996);
nor U6079 (N_6079,N_5125,N_5057);
or U6080 (N_6080,N_5810,N_5971);
nor U6081 (N_6081,N_5834,N_5541);
nand U6082 (N_6082,N_5043,N_5904);
and U6083 (N_6083,N_5619,N_5782);
xnor U6084 (N_6084,N_5860,N_5567);
nand U6085 (N_6085,N_5653,N_5011);
and U6086 (N_6086,N_5498,N_5922);
or U6087 (N_6087,N_5036,N_5774);
xnor U6088 (N_6088,N_5306,N_5197);
and U6089 (N_6089,N_5267,N_5246);
nor U6090 (N_6090,N_5959,N_5457);
or U6091 (N_6091,N_5884,N_5526);
or U6092 (N_6092,N_5434,N_5739);
nand U6093 (N_6093,N_5328,N_5193);
nor U6094 (N_6094,N_5190,N_5304);
xnor U6095 (N_6095,N_5509,N_5372);
and U6096 (N_6096,N_5300,N_5437);
nor U6097 (N_6097,N_5354,N_5334);
nor U6098 (N_6098,N_5900,N_5512);
or U6099 (N_6099,N_5910,N_5762);
nor U6100 (N_6100,N_5502,N_5271);
and U6101 (N_6101,N_5920,N_5964);
or U6102 (N_6102,N_5186,N_5480);
and U6103 (N_6103,N_5856,N_5645);
and U6104 (N_6104,N_5517,N_5598);
nor U6105 (N_6105,N_5275,N_5325);
and U6106 (N_6106,N_5592,N_5908);
nor U6107 (N_6107,N_5818,N_5440);
xnor U6108 (N_6108,N_5417,N_5128);
xor U6109 (N_6109,N_5469,N_5280);
nand U6110 (N_6110,N_5997,N_5847);
nor U6111 (N_6111,N_5775,N_5070);
xor U6112 (N_6112,N_5722,N_5062);
xor U6113 (N_6113,N_5858,N_5685);
xnor U6114 (N_6114,N_5496,N_5035);
nand U6115 (N_6115,N_5465,N_5941);
and U6116 (N_6116,N_5759,N_5096);
and U6117 (N_6117,N_5850,N_5413);
nor U6118 (N_6118,N_5102,N_5862);
nor U6119 (N_6119,N_5899,N_5794);
or U6120 (N_6120,N_5311,N_5210);
and U6121 (N_6121,N_5673,N_5634);
or U6122 (N_6122,N_5602,N_5967);
xnor U6123 (N_6123,N_5785,N_5724);
nand U6124 (N_6124,N_5605,N_5888);
and U6125 (N_6125,N_5629,N_5756);
and U6126 (N_6126,N_5717,N_5501);
xnor U6127 (N_6127,N_5402,N_5013);
xor U6128 (N_6128,N_5789,N_5798);
and U6129 (N_6129,N_5819,N_5119);
nand U6130 (N_6130,N_5586,N_5727);
xnor U6131 (N_6131,N_5788,N_5064);
and U6132 (N_6132,N_5319,N_5268);
and U6133 (N_6133,N_5702,N_5781);
or U6134 (N_6134,N_5162,N_5108);
nand U6135 (N_6135,N_5172,N_5554);
and U6136 (N_6136,N_5518,N_5934);
nand U6137 (N_6137,N_5390,N_5768);
nand U6138 (N_6138,N_5905,N_5249);
nor U6139 (N_6139,N_5278,N_5243);
or U6140 (N_6140,N_5338,N_5427);
nor U6141 (N_6141,N_5990,N_5814);
nand U6142 (N_6142,N_5355,N_5857);
nor U6143 (N_6143,N_5393,N_5625);
xnor U6144 (N_6144,N_5519,N_5561);
nor U6145 (N_6145,N_5520,N_5167);
or U6146 (N_6146,N_5483,N_5088);
and U6147 (N_6147,N_5504,N_5993);
nor U6148 (N_6148,N_5989,N_5690);
or U6149 (N_6149,N_5231,N_5575);
nor U6150 (N_6150,N_5237,N_5136);
nor U6151 (N_6151,N_5532,N_5744);
xor U6152 (N_6152,N_5965,N_5914);
nand U6153 (N_6153,N_5130,N_5924);
or U6154 (N_6154,N_5205,N_5408);
xnor U6155 (N_6155,N_5196,N_5140);
and U6156 (N_6156,N_5715,N_5038);
xor U6157 (N_6157,N_5220,N_5907);
nand U6158 (N_6158,N_5034,N_5766);
nand U6159 (N_6159,N_5481,N_5446);
xnor U6160 (N_6160,N_5299,N_5986);
or U6161 (N_6161,N_5443,N_5335);
or U6162 (N_6162,N_5048,N_5143);
and U6163 (N_6163,N_5550,N_5239);
xnor U6164 (N_6164,N_5556,N_5151);
nor U6165 (N_6165,N_5174,N_5534);
nand U6166 (N_6166,N_5820,N_5613);
or U6167 (N_6167,N_5484,N_5356);
nor U6168 (N_6168,N_5091,N_5405);
nor U6169 (N_6169,N_5221,N_5514);
xor U6170 (N_6170,N_5467,N_5684);
and U6171 (N_6171,N_5422,N_5180);
or U6172 (N_6172,N_5421,N_5795);
or U6173 (N_6173,N_5923,N_5379);
or U6174 (N_6174,N_5607,N_5885);
and U6175 (N_6175,N_5911,N_5262);
xor U6176 (N_6176,N_5488,N_5233);
nor U6177 (N_6177,N_5758,N_5080);
and U6178 (N_6178,N_5751,N_5358);
and U6179 (N_6179,N_5241,N_5182);
nand U6180 (N_6180,N_5981,N_5170);
and U6181 (N_6181,N_5450,N_5564);
xor U6182 (N_6182,N_5786,N_5737);
nand U6183 (N_6183,N_5745,N_5569);
or U6184 (N_6184,N_5801,N_5284);
nor U6185 (N_6185,N_5638,N_5822);
nand U6186 (N_6186,N_5460,N_5441);
and U6187 (N_6187,N_5864,N_5103);
and U6188 (N_6188,N_5215,N_5754);
nand U6189 (N_6189,N_5972,N_5696);
nor U6190 (N_6190,N_5445,N_5797);
nand U6191 (N_6191,N_5208,N_5870);
nand U6192 (N_6192,N_5365,N_5282);
nand U6193 (N_6193,N_5225,N_5497);
or U6194 (N_6194,N_5211,N_5007);
and U6195 (N_6195,N_5733,N_5838);
xnor U6196 (N_6196,N_5340,N_5770);
xor U6197 (N_6197,N_5670,N_5308);
xor U6198 (N_6198,N_5218,N_5719);
nor U6199 (N_6199,N_5320,N_5018);
or U6200 (N_6200,N_5978,N_5166);
nor U6201 (N_6201,N_5661,N_5713);
nor U6202 (N_6202,N_5783,N_5059);
and U6203 (N_6203,N_5337,N_5614);
and U6204 (N_6204,N_5593,N_5976);
or U6205 (N_6205,N_5458,N_5764);
xnor U6206 (N_6206,N_5219,N_5823);
and U6207 (N_6207,N_5269,N_5478);
and U6208 (N_6208,N_5341,N_5042);
or U6209 (N_6209,N_5662,N_5621);
xnor U6210 (N_6210,N_5635,N_5784);
and U6211 (N_6211,N_5543,N_5353);
or U6212 (N_6212,N_5226,N_5429);
or U6213 (N_6213,N_5682,N_5024);
and U6214 (N_6214,N_5141,N_5292);
nor U6215 (N_6215,N_5887,N_5022);
xnor U6216 (N_6216,N_5677,N_5777);
xor U6217 (N_6217,N_5164,N_5124);
and U6218 (N_6218,N_5949,N_5531);
xnor U6219 (N_6219,N_5580,N_5711);
or U6220 (N_6220,N_5082,N_5671);
xnor U6221 (N_6221,N_5943,N_5826);
nor U6222 (N_6222,N_5214,N_5792);
nand U6223 (N_6223,N_5309,N_5617);
or U6224 (N_6224,N_5277,N_5804);
nor U6225 (N_6225,N_5098,N_5120);
nand U6226 (N_6226,N_5640,N_5367);
and U6227 (N_6227,N_5686,N_5843);
xor U6228 (N_6228,N_5487,N_5494);
xnor U6229 (N_6229,N_5126,N_5929);
and U6230 (N_6230,N_5297,N_5448);
nor U6231 (N_6231,N_5799,N_5880);
nand U6232 (N_6232,N_5266,N_5779);
xor U6233 (N_6233,N_5366,N_5152);
nand U6234 (N_6234,N_5005,N_5324);
xor U6235 (N_6235,N_5153,N_5155);
and U6236 (N_6236,N_5701,N_5397);
or U6237 (N_6237,N_5411,N_5479);
nor U6238 (N_6238,N_5599,N_5522);
and U6239 (N_6239,N_5937,N_5891);
nor U6240 (N_6240,N_5350,N_5395);
nand U6241 (N_6241,N_5837,N_5732);
or U6242 (N_6242,N_5216,N_5085);
xnor U6243 (N_6243,N_5289,N_5938);
nand U6244 (N_6244,N_5841,N_5321);
nand U6245 (N_6245,N_5660,N_5548);
and U6246 (N_6246,N_5709,N_5290);
nand U6247 (N_6247,N_5099,N_5272);
or U6248 (N_6248,N_5361,N_5204);
and U6249 (N_6249,N_5415,N_5148);
or U6250 (N_6250,N_5185,N_5650);
and U6251 (N_6251,N_5966,N_5869);
or U6252 (N_6252,N_5332,N_5139);
and U6253 (N_6253,N_5946,N_5352);
or U6254 (N_6254,N_5305,N_5313);
nand U6255 (N_6255,N_5896,N_5926);
nor U6256 (N_6256,N_5398,N_5761);
or U6257 (N_6257,N_5054,N_5995);
xnor U6258 (N_6258,N_5156,N_5591);
nor U6259 (N_6259,N_5302,N_5664);
xor U6260 (N_6260,N_5069,N_5028);
or U6261 (N_6261,N_5898,N_5270);
or U6262 (N_6262,N_5742,N_5595);
nand U6263 (N_6263,N_5571,N_5287);
xor U6264 (N_6264,N_5961,N_5228);
nand U6265 (N_6265,N_5245,N_5476);
or U6266 (N_6266,N_5016,N_5138);
or U6267 (N_6267,N_5493,N_5442);
and U6268 (N_6268,N_5259,N_5565);
or U6269 (N_6269,N_5439,N_5087);
nand U6270 (N_6270,N_5980,N_5681);
or U6271 (N_6271,N_5930,N_5707);
or U6272 (N_6272,N_5572,N_5175);
nand U6273 (N_6273,N_5377,N_5928);
nor U6274 (N_6274,N_5373,N_5563);
xnor U6275 (N_6275,N_5712,N_5470);
or U6276 (N_6276,N_5090,N_5957);
or U6277 (N_6277,N_5609,N_5985);
nor U6278 (N_6278,N_5063,N_5835);
xnor U6279 (N_6279,N_5115,N_5414);
nor U6280 (N_6280,N_5436,N_5652);
nor U6281 (N_6281,N_5697,N_5050);
and U6282 (N_6282,N_5146,N_5555);
or U6283 (N_6283,N_5008,N_5817);
xnor U6284 (N_6284,N_5121,N_5209);
xnor U6285 (N_6285,N_5693,N_5207);
xor U6286 (N_6286,N_5014,N_5939);
nor U6287 (N_6287,N_5601,N_5963);
or U6288 (N_6288,N_5610,N_5023);
nor U6289 (N_6289,N_5633,N_5691);
nor U6290 (N_6290,N_5079,N_5665);
nand U6291 (N_6291,N_5988,N_5903);
nor U6292 (N_6292,N_5604,N_5927);
and U6293 (N_6293,N_5491,N_5894);
xnor U6294 (N_6294,N_5296,N_5699);
and U6295 (N_6295,N_5212,N_5286);
xor U6296 (N_6296,N_5310,N_5726);
and U6297 (N_6297,N_5678,N_5529);
and U6298 (N_6298,N_5168,N_5728);
and U6299 (N_6299,N_5611,N_5330);
or U6300 (N_6300,N_5829,N_5116);
nand U6301 (N_6301,N_5979,N_5616);
xor U6302 (N_6302,N_5984,N_5045);
nor U6303 (N_6303,N_5298,N_5157);
nand U6304 (N_6304,N_5384,N_5452);
xor U6305 (N_6305,N_5875,N_5184);
xnor U6306 (N_6306,N_5791,N_5897);
nor U6307 (N_6307,N_5165,N_5106);
xor U6308 (N_6308,N_5500,N_5113);
nand U6309 (N_6309,N_5597,N_5944);
nand U6310 (N_6310,N_5776,N_5412);
xor U6311 (N_6311,N_5396,N_5867);
nand U6312 (N_6312,N_5871,N_5735);
nor U6313 (N_6313,N_5435,N_5545);
nand U6314 (N_6314,N_5626,N_5760);
nor U6315 (N_6315,N_5559,N_5003);
and U6316 (N_6316,N_5477,N_5100);
or U6317 (N_6317,N_5364,N_5033);
or U6318 (N_6318,N_5710,N_5388);
nor U6319 (N_6319,N_5741,N_5370);
or U6320 (N_6320,N_5950,N_5235);
nand U6321 (N_6321,N_5808,N_5861);
nand U6322 (N_6322,N_5419,N_5183);
nand U6323 (N_6323,N_5510,N_5468);
nor U6324 (N_6324,N_5010,N_5755);
and U6325 (N_6325,N_5463,N_5983);
xor U6326 (N_6326,N_5179,N_5765);
or U6327 (N_6327,N_5582,N_5919);
nor U6328 (N_6328,N_5456,N_5029);
xor U6329 (N_6329,N_5746,N_5973);
and U6330 (N_6330,N_5803,N_5181);
nor U6331 (N_6331,N_5095,N_5447);
nor U6332 (N_6332,N_5952,N_5072);
nor U6333 (N_6333,N_5077,N_5101);
nand U6334 (N_6334,N_5506,N_5842);
and U6335 (N_6335,N_5658,N_5730);
xnor U6336 (N_6336,N_5021,N_5656);
or U6337 (N_6337,N_5533,N_5195);
nor U6338 (N_6338,N_5620,N_5889);
xor U6339 (N_6339,N_5075,N_5839);
nand U6340 (N_6340,N_5382,N_5049);
or U6341 (N_6341,N_5323,N_5314);
and U6342 (N_6342,N_5991,N_5694);
or U6343 (N_6343,N_5796,N_5958);
nor U6344 (N_6344,N_5863,N_5111);
nor U6345 (N_6345,N_5668,N_5866);
and U6346 (N_6346,N_5094,N_5692);
or U6347 (N_6347,N_5723,N_5250);
and U6348 (N_6348,N_5394,N_5086);
or U6349 (N_6349,N_5137,N_5743);
and U6350 (N_6350,N_5663,N_5081);
nand U6351 (N_6351,N_5171,N_5260);
xor U6352 (N_6352,N_5513,N_5206);
xor U6353 (N_6353,N_5790,N_5721);
xor U6354 (N_6354,N_5731,N_5368);
nand U6355 (N_6355,N_5844,N_5288);
nor U6356 (N_6356,N_5025,N_5222);
xor U6357 (N_6357,N_5683,N_5912);
and U6358 (N_6358,N_5767,N_5006);
nor U6359 (N_6359,N_5351,N_5772);
or U6360 (N_6360,N_5178,N_5893);
xor U6361 (N_6361,N_5150,N_5925);
nand U6362 (N_6362,N_5129,N_5521);
xor U6363 (N_6363,N_5424,N_5757);
xnor U6364 (N_6364,N_5455,N_5705);
nand U6365 (N_6365,N_5053,N_5301);
xnor U6366 (N_6366,N_5940,N_5399);
xnor U6367 (N_6367,N_5189,N_5107);
or U6368 (N_6368,N_5078,N_5734);
nand U6369 (N_6369,N_5587,N_5173);
nand U6370 (N_6370,N_5851,N_5044);
xor U6371 (N_6371,N_5666,N_5566);
xor U6372 (N_6372,N_5865,N_5000);
xnor U6373 (N_6373,N_5017,N_5073);
or U6374 (N_6374,N_5780,N_5942);
nor U6375 (N_6375,N_5811,N_5092);
nor U6376 (N_6376,N_5603,N_5538);
nor U6377 (N_6377,N_5987,N_5704);
xnor U6378 (N_6378,N_5453,N_5632);
or U6379 (N_6379,N_5342,N_5307);
xor U6380 (N_6380,N_5135,N_5027);
and U6381 (N_6381,N_5570,N_5285);
nand U6382 (N_6382,N_5953,N_5247);
xor U6383 (N_6383,N_5089,N_5833);
nand U6384 (N_6384,N_5159,N_5527);
and U6385 (N_6385,N_5105,N_5462);
nor U6386 (N_6386,N_5316,N_5579);
nor U6387 (N_6387,N_5574,N_5549);
xnor U6388 (N_6388,N_5110,N_5474);
and U6389 (N_6389,N_5590,N_5495);
nand U6390 (N_6390,N_5982,N_5339);
xnor U6391 (N_6391,N_5577,N_5909);
and U6392 (N_6392,N_5420,N_5242);
and U6393 (N_6393,N_5291,N_5187);
nand U6394 (N_6394,N_5236,N_5404);
and U6395 (N_6395,N_5192,N_5132);
nor U6396 (N_6396,N_5918,N_5669);
nor U6397 (N_6397,N_5061,N_5974);
nand U6398 (N_6398,N_5680,N_5066);
or U6399 (N_6399,N_5687,N_5257);
or U6400 (N_6400,N_5718,N_5131);
xnor U6401 (N_6401,N_5433,N_5492);
xor U6402 (N_6402,N_5945,N_5104);
xor U6403 (N_6403,N_5256,N_5901);
nand U6404 (N_6404,N_5444,N_5540);
and U6405 (N_6405,N_5438,N_5161);
or U6406 (N_6406,N_5679,N_5327);
nor U6407 (N_6407,N_5584,N_5145);
nand U6408 (N_6408,N_5312,N_5430);
or U6409 (N_6409,N_5623,N_5471);
and U6410 (N_6410,N_5459,N_5542);
nor U6411 (N_6411,N_5281,N_5879);
nor U6412 (N_6412,N_5651,N_5381);
xor U6413 (N_6413,N_5273,N_5854);
xor U6414 (N_6414,N_5675,N_5736);
and U6415 (N_6415,N_5931,N_5748);
or U6416 (N_6416,N_5191,N_5855);
and U6417 (N_6417,N_5134,N_5112);
xnor U6418 (N_6418,N_5065,N_5508);
nand U6419 (N_6419,N_5935,N_5530);
nor U6420 (N_6420,N_5127,N_5667);
nand U6421 (N_6421,N_5133,N_5283);
xnor U6422 (N_6422,N_5674,N_5840);
and U6423 (N_6423,N_5778,N_5816);
nor U6424 (N_6424,N_5802,N_5809);
or U6425 (N_6425,N_5750,N_5947);
or U6426 (N_6426,N_5097,N_5646);
xor U6427 (N_6427,N_5449,N_5992);
or U6428 (N_6428,N_5932,N_5853);
nor U6429 (N_6429,N_5596,N_5374);
xor U6430 (N_6430,N_5279,N_5916);
nor U6431 (N_6431,N_5622,N_5369);
nand U6432 (N_6432,N_5409,N_5975);
or U6433 (N_6433,N_5969,N_5868);
or U6434 (N_6434,N_5544,N_5084);
or U6435 (N_6435,N_5425,N_5160);
or U6436 (N_6436,N_5432,N_5876);
nand U6437 (N_6437,N_5295,N_5695);
nand U6438 (N_6438,N_5769,N_5639);
nand U6439 (N_6439,N_5594,N_5849);
xor U6440 (N_6440,N_5523,N_5568);
and U6441 (N_6441,N_5832,N_5318);
nand U6442 (N_6442,N_5052,N_5423);
nand U6443 (N_6443,N_5562,N_5499);
and U6444 (N_6444,N_5040,N_5238);
or U6445 (N_6445,N_5227,N_5347);
and U6446 (N_6446,N_5031,N_5951);
xor U6447 (N_6447,N_5706,N_5657);
xnor U6448 (N_6448,N_5507,N_5144);
or U6449 (N_6449,N_5576,N_5147);
or U6450 (N_6450,N_5771,N_5647);
nor U6451 (N_6451,N_5020,N_5836);
or U6452 (N_6452,N_5019,N_5060);
or U6453 (N_6453,N_5303,N_5198);
nand U6454 (N_6454,N_5882,N_5348);
or U6455 (N_6455,N_5154,N_5400);
or U6456 (N_6456,N_5921,N_5547);
nand U6457 (N_6457,N_5960,N_5401);
xnor U6458 (N_6458,N_5873,N_5349);
or U6459 (N_6459,N_5878,N_5763);
and U6460 (N_6460,N_5573,N_5336);
nand U6461 (N_6461,N_5881,N_5902);
xnor U6462 (N_6462,N_5224,N_5700);
or U6463 (N_6463,N_5805,N_5644);
nor U6464 (N_6464,N_5970,N_5637);
and U6465 (N_6465,N_5217,N_5948);
and U6466 (N_6466,N_5600,N_5643);
nor U6467 (N_6467,N_5326,N_5248);
and U6468 (N_6468,N_5654,N_5473);
xor U6469 (N_6469,N_5536,N_5505);
nor U6470 (N_6470,N_5806,N_5585);
and U6471 (N_6471,N_5852,N_5815);
and U6472 (N_6472,N_5244,N_5725);
and U6473 (N_6473,N_5109,N_5859);
xor U6474 (N_6474,N_5009,N_5274);
xor U6475 (N_6475,N_5557,N_5890);
and U6476 (N_6476,N_5800,N_5752);
nand U6477 (N_6477,N_5345,N_5977);
xnor U6478 (N_6478,N_5689,N_5824);
or U6479 (N_6479,N_5475,N_5915);
xor U6480 (N_6480,N_5359,N_5294);
xor U6481 (N_6481,N_5848,N_5630);
or U6482 (N_6482,N_5234,N_5551);
nor U6483 (N_6483,N_5317,N_5537);
xor U6484 (N_6484,N_5056,N_5773);
nand U6485 (N_6485,N_5276,N_5230);
and U6486 (N_6486,N_5642,N_5845);
or U6487 (N_6487,N_5329,N_5461);
and U6488 (N_6488,N_5068,N_5255);
xnor U6489 (N_6489,N_5821,N_5827);
nand U6490 (N_6490,N_5641,N_5539);
nand U6491 (N_6491,N_5485,N_5883);
xor U6492 (N_6492,N_5194,N_5389);
or U6493 (N_6493,N_5416,N_5387);
nand U6494 (N_6494,N_5026,N_5612);
or U6495 (N_6495,N_5490,N_5968);
nor U6496 (N_6496,N_5344,N_5489);
nor U6497 (N_6497,N_5391,N_5076);
and U6498 (N_6498,N_5698,N_5403);
xor U6499 (N_6499,N_5877,N_5787);
xnor U6500 (N_6500,N_5560,N_5674);
nor U6501 (N_6501,N_5017,N_5964);
nor U6502 (N_6502,N_5722,N_5294);
nand U6503 (N_6503,N_5256,N_5250);
nand U6504 (N_6504,N_5040,N_5656);
or U6505 (N_6505,N_5619,N_5647);
or U6506 (N_6506,N_5555,N_5215);
or U6507 (N_6507,N_5835,N_5200);
nand U6508 (N_6508,N_5552,N_5315);
nand U6509 (N_6509,N_5196,N_5824);
or U6510 (N_6510,N_5497,N_5582);
and U6511 (N_6511,N_5023,N_5002);
or U6512 (N_6512,N_5002,N_5064);
or U6513 (N_6513,N_5737,N_5557);
xnor U6514 (N_6514,N_5752,N_5279);
and U6515 (N_6515,N_5979,N_5981);
nor U6516 (N_6516,N_5980,N_5809);
or U6517 (N_6517,N_5625,N_5554);
nor U6518 (N_6518,N_5269,N_5859);
or U6519 (N_6519,N_5530,N_5402);
or U6520 (N_6520,N_5140,N_5929);
nor U6521 (N_6521,N_5207,N_5792);
nand U6522 (N_6522,N_5638,N_5746);
nand U6523 (N_6523,N_5303,N_5027);
or U6524 (N_6524,N_5116,N_5005);
nand U6525 (N_6525,N_5811,N_5925);
xnor U6526 (N_6526,N_5367,N_5058);
nor U6527 (N_6527,N_5073,N_5636);
nor U6528 (N_6528,N_5376,N_5528);
and U6529 (N_6529,N_5355,N_5471);
and U6530 (N_6530,N_5824,N_5505);
nand U6531 (N_6531,N_5479,N_5781);
and U6532 (N_6532,N_5043,N_5651);
xor U6533 (N_6533,N_5076,N_5490);
or U6534 (N_6534,N_5069,N_5124);
nand U6535 (N_6535,N_5030,N_5368);
and U6536 (N_6536,N_5266,N_5848);
nand U6537 (N_6537,N_5031,N_5489);
xor U6538 (N_6538,N_5806,N_5334);
nand U6539 (N_6539,N_5866,N_5392);
nor U6540 (N_6540,N_5062,N_5534);
nand U6541 (N_6541,N_5950,N_5020);
and U6542 (N_6542,N_5672,N_5063);
or U6543 (N_6543,N_5322,N_5926);
nor U6544 (N_6544,N_5144,N_5642);
nand U6545 (N_6545,N_5000,N_5753);
xnor U6546 (N_6546,N_5960,N_5728);
xor U6547 (N_6547,N_5559,N_5361);
and U6548 (N_6548,N_5812,N_5449);
or U6549 (N_6549,N_5941,N_5110);
and U6550 (N_6550,N_5611,N_5115);
xor U6551 (N_6551,N_5377,N_5823);
nand U6552 (N_6552,N_5506,N_5623);
nor U6553 (N_6553,N_5754,N_5216);
and U6554 (N_6554,N_5745,N_5365);
or U6555 (N_6555,N_5413,N_5772);
nor U6556 (N_6556,N_5701,N_5611);
nand U6557 (N_6557,N_5886,N_5653);
xnor U6558 (N_6558,N_5029,N_5620);
xnor U6559 (N_6559,N_5140,N_5953);
xor U6560 (N_6560,N_5329,N_5415);
or U6561 (N_6561,N_5330,N_5635);
nor U6562 (N_6562,N_5394,N_5577);
xnor U6563 (N_6563,N_5148,N_5341);
nor U6564 (N_6564,N_5698,N_5336);
nand U6565 (N_6565,N_5232,N_5539);
nand U6566 (N_6566,N_5067,N_5840);
nor U6567 (N_6567,N_5319,N_5233);
or U6568 (N_6568,N_5934,N_5521);
or U6569 (N_6569,N_5489,N_5403);
nor U6570 (N_6570,N_5346,N_5471);
or U6571 (N_6571,N_5880,N_5691);
xor U6572 (N_6572,N_5145,N_5627);
nand U6573 (N_6573,N_5803,N_5401);
nand U6574 (N_6574,N_5042,N_5063);
xnor U6575 (N_6575,N_5143,N_5352);
and U6576 (N_6576,N_5237,N_5696);
nor U6577 (N_6577,N_5593,N_5797);
nor U6578 (N_6578,N_5088,N_5591);
nor U6579 (N_6579,N_5051,N_5769);
nand U6580 (N_6580,N_5156,N_5281);
xor U6581 (N_6581,N_5015,N_5689);
nand U6582 (N_6582,N_5802,N_5856);
or U6583 (N_6583,N_5304,N_5760);
and U6584 (N_6584,N_5048,N_5865);
nor U6585 (N_6585,N_5360,N_5779);
xor U6586 (N_6586,N_5079,N_5993);
or U6587 (N_6587,N_5674,N_5871);
nor U6588 (N_6588,N_5492,N_5597);
xor U6589 (N_6589,N_5088,N_5662);
and U6590 (N_6590,N_5984,N_5884);
nand U6591 (N_6591,N_5764,N_5367);
or U6592 (N_6592,N_5740,N_5090);
nand U6593 (N_6593,N_5915,N_5070);
nand U6594 (N_6594,N_5507,N_5940);
or U6595 (N_6595,N_5764,N_5285);
or U6596 (N_6596,N_5850,N_5664);
nor U6597 (N_6597,N_5818,N_5223);
or U6598 (N_6598,N_5575,N_5248);
nand U6599 (N_6599,N_5286,N_5691);
and U6600 (N_6600,N_5838,N_5195);
and U6601 (N_6601,N_5566,N_5849);
and U6602 (N_6602,N_5981,N_5413);
nor U6603 (N_6603,N_5452,N_5290);
or U6604 (N_6604,N_5220,N_5795);
and U6605 (N_6605,N_5333,N_5517);
nand U6606 (N_6606,N_5846,N_5712);
nor U6607 (N_6607,N_5294,N_5175);
xor U6608 (N_6608,N_5969,N_5307);
and U6609 (N_6609,N_5101,N_5485);
and U6610 (N_6610,N_5611,N_5634);
xor U6611 (N_6611,N_5722,N_5657);
and U6612 (N_6612,N_5111,N_5761);
xor U6613 (N_6613,N_5252,N_5300);
or U6614 (N_6614,N_5844,N_5164);
and U6615 (N_6615,N_5602,N_5448);
nor U6616 (N_6616,N_5932,N_5732);
and U6617 (N_6617,N_5458,N_5047);
xor U6618 (N_6618,N_5352,N_5669);
nand U6619 (N_6619,N_5701,N_5087);
and U6620 (N_6620,N_5866,N_5286);
xor U6621 (N_6621,N_5756,N_5031);
xor U6622 (N_6622,N_5107,N_5946);
and U6623 (N_6623,N_5838,N_5250);
and U6624 (N_6624,N_5254,N_5336);
xor U6625 (N_6625,N_5573,N_5494);
nand U6626 (N_6626,N_5115,N_5788);
and U6627 (N_6627,N_5152,N_5083);
xnor U6628 (N_6628,N_5037,N_5707);
nand U6629 (N_6629,N_5090,N_5966);
or U6630 (N_6630,N_5810,N_5747);
nor U6631 (N_6631,N_5337,N_5765);
xnor U6632 (N_6632,N_5475,N_5195);
nand U6633 (N_6633,N_5919,N_5556);
xnor U6634 (N_6634,N_5665,N_5084);
nor U6635 (N_6635,N_5434,N_5354);
or U6636 (N_6636,N_5454,N_5233);
xnor U6637 (N_6637,N_5619,N_5337);
nand U6638 (N_6638,N_5135,N_5639);
xor U6639 (N_6639,N_5469,N_5529);
or U6640 (N_6640,N_5869,N_5890);
and U6641 (N_6641,N_5699,N_5673);
or U6642 (N_6642,N_5079,N_5512);
nand U6643 (N_6643,N_5718,N_5478);
or U6644 (N_6644,N_5806,N_5992);
nor U6645 (N_6645,N_5226,N_5716);
or U6646 (N_6646,N_5666,N_5991);
or U6647 (N_6647,N_5405,N_5315);
xnor U6648 (N_6648,N_5023,N_5878);
or U6649 (N_6649,N_5863,N_5779);
xnor U6650 (N_6650,N_5709,N_5783);
and U6651 (N_6651,N_5193,N_5092);
or U6652 (N_6652,N_5294,N_5688);
xor U6653 (N_6653,N_5331,N_5250);
xnor U6654 (N_6654,N_5971,N_5848);
nand U6655 (N_6655,N_5785,N_5562);
nor U6656 (N_6656,N_5539,N_5433);
nand U6657 (N_6657,N_5701,N_5665);
or U6658 (N_6658,N_5829,N_5114);
xnor U6659 (N_6659,N_5892,N_5237);
or U6660 (N_6660,N_5820,N_5125);
and U6661 (N_6661,N_5176,N_5955);
xnor U6662 (N_6662,N_5896,N_5756);
nand U6663 (N_6663,N_5273,N_5267);
nand U6664 (N_6664,N_5195,N_5849);
nor U6665 (N_6665,N_5896,N_5300);
nor U6666 (N_6666,N_5766,N_5984);
nand U6667 (N_6667,N_5840,N_5286);
and U6668 (N_6668,N_5860,N_5246);
and U6669 (N_6669,N_5764,N_5242);
or U6670 (N_6670,N_5865,N_5733);
xor U6671 (N_6671,N_5837,N_5281);
nand U6672 (N_6672,N_5299,N_5117);
or U6673 (N_6673,N_5854,N_5359);
and U6674 (N_6674,N_5855,N_5791);
or U6675 (N_6675,N_5312,N_5969);
xnor U6676 (N_6676,N_5105,N_5092);
or U6677 (N_6677,N_5028,N_5360);
nor U6678 (N_6678,N_5640,N_5486);
or U6679 (N_6679,N_5615,N_5696);
or U6680 (N_6680,N_5274,N_5609);
or U6681 (N_6681,N_5848,N_5932);
and U6682 (N_6682,N_5114,N_5856);
and U6683 (N_6683,N_5925,N_5012);
and U6684 (N_6684,N_5529,N_5102);
and U6685 (N_6685,N_5975,N_5733);
nor U6686 (N_6686,N_5472,N_5241);
nor U6687 (N_6687,N_5475,N_5192);
nand U6688 (N_6688,N_5996,N_5057);
nor U6689 (N_6689,N_5369,N_5092);
nor U6690 (N_6690,N_5834,N_5857);
xor U6691 (N_6691,N_5956,N_5614);
and U6692 (N_6692,N_5503,N_5204);
and U6693 (N_6693,N_5150,N_5147);
nand U6694 (N_6694,N_5178,N_5434);
xnor U6695 (N_6695,N_5073,N_5965);
or U6696 (N_6696,N_5274,N_5865);
nor U6697 (N_6697,N_5306,N_5523);
and U6698 (N_6698,N_5177,N_5042);
or U6699 (N_6699,N_5145,N_5089);
nand U6700 (N_6700,N_5468,N_5677);
xor U6701 (N_6701,N_5053,N_5898);
or U6702 (N_6702,N_5772,N_5085);
nand U6703 (N_6703,N_5106,N_5595);
xor U6704 (N_6704,N_5978,N_5325);
xnor U6705 (N_6705,N_5396,N_5226);
or U6706 (N_6706,N_5235,N_5150);
or U6707 (N_6707,N_5411,N_5346);
nor U6708 (N_6708,N_5202,N_5408);
xor U6709 (N_6709,N_5153,N_5132);
or U6710 (N_6710,N_5182,N_5685);
nand U6711 (N_6711,N_5146,N_5075);
nor U6712 (N_6712,N_5126,N_5589);
or U6713 (N_6713,N_5120,N_5528);
or U6714 (N_6714,N_5488,N_5885);
nand U6715 (N_6715,N_5106,N_5785);
xor U6716 (N_6716,N_5373,N_5463);
nor U6717 (N_6717,N_5462,N_5148);
xnor U6718 (N_6718,N_5656,N_5414);
nand U6719 (N_6719,N_5976,N_5795);
nand U6720 (N_6720,N_5063,N_5040);
nor U6721 (N_6721,N_5697,N_5465);
nand U6722 (N_6722,N_5883,N_5025);
and U6723 (N_6723,N_5039,N_5399);
and U6724 (N_6724,N_5992,N_5302);
nor U6725 (N_6725,N_5747,N_5076);
xor U6726 (N_6726,N_5180,N_5508);
and U6727 (N_6727,N_5790,N_5409);
xor U6728 (N_6728,N_5058,N_5835);
xnor U6729 (N_6729,N_5433,N_5079);
nor U6730 (N_6730,N_5077,N_5090);
and U6731 (N_6731,N_5687,N_5073);
nor U6732 (N_6732,N_5333,N_5832);
and U6733 (N_6733,N_5361,N_5827);
nor U6734 (N_6734,N_5876,N_5600);
nand U6735 (N_6735,N_5489,N_5418);
nor U6736 (N_6736,N_5008,N_5621);
nand U6737 (N_6737,N_5815,N_5775);
nor U6738 (N_6738,N_5453,N_5196);
and U6739 (N_6739,N_5840,N_5191);
or U6740 (N_6740,N_5490,N_5508);
or U6741 (N_6741,N_5106,N_5030);
nor U6742 (N_6742,N_5634,N_5459);
nand U6743 (N_6743,N_5564,N_5336);
and U6744 (N_6744,N_5390,N_5249);
or U6745 (N_6745,N_5294,N_5822);
and U6746 (N_6746,N_5675,N_5785);
or U6747 (N_6747,N_5727,N_5359);
nor U6748 (N_6748,N_5843,N_5879);
xor U6749 (N_6749,N_5467,N_5213);
nor U6750 (N_6750,N_5184,N_5451);
xor U6751 (N_6751,N_5823,N_5616);
xnor U6752 (N_6752,N_5338,N_5986);
and U6753 (N_6753,N_5377,N_5288);
nor U6754 (N_6754,N_5585,N_5622);
xnor U6755 (N_6755,N_5011,N_5164);
and U6756 (N_6756,N_5637,N_5085);
or U6757 (N_6757,N_5296,N_5416);
nand U6758 (N_6758,N_5246,N_5711);
nor U6759 (N_6759,N_5467,N_5784);
or U6760 (N_6760,N_5603,N_5556);
nand U6761 (N_6761,N_5840,N_5425);
nor U6762 (N_6762,N_5913,N_5180);
nand U6763 (N_6763,N_5808,N_5788);
nor U6764 (N_6764,N_5529,N_5360);
or U6765 (N_6765,N_5023,N_5201);
nor U6766 (N_6766,N_5338,N_5243);
or U6767 (N_6767,N_5362,N_5554);
and U6768 (N_6768,N_5069,N_5346);
nand U6769 (N_6769,N_5594,N_5342);
nor U6770 (N_6770,N_5240,N_5842);
and U6771 (N_6771,N_5186,N_5682);
nor U6772 (N_6772,N_5402,N_5918);
nand U6773 (N_6773,N_5700,N_5219);
or U6774 (N_6774,N_5215,N_5779);
and U6775 (N_6775,N_5718,N_5217);
nor U6776 (N_6776,N_5730,N_5693);
or U6777 (N_6777,N_5914,N_5715);
or U6778 (N_6778,N_5907,N_5786);
xor U6779 (N_6779,N_5426,N_5203);
nor U6780 (N_6780,N_5727,N_5666);
or U6781 (N_6781,N_5720,N_5860);
or U6782 (N_6782,N_5177,N_5099);
nor U6783 (N_6783,N_5534,N_5245);
nand U6784 (N_6784,N_5044,N_5394);
nor U6785 (N_6785,N_5551,N_5613);
xnor U6786 (N_6786,N_5104,N_5541);
nand U6787 (N_6787,N_5481,N_5327);
and U6788 (N_6788,N_5765,N_5902);
nor U6789 (N_6789,N_5508,N_5987);
xor U6790 (N_6790,N_5704,N_5168);
nor U6791 (N_6791,N_5916,N_5828);
and U6792 (N_6792,N_5406,N_5220);
nand U6793 (N_6793,N_5263,N_5626);
and U6794 (N_6794,N_5109,N_5666);
nand U6795 (N_6795,N_5254,N_5231);
xor U6796 (N_6796,N_5646,N_5645);
xor U6797 (N_6797,N_5949,N_5153);
and U6798 (N_6798,N_5755,N_5273);
or U6799 (N_6799,N_5035,N_5998);
nand U6800 (N_6800,N_5432,N_5805);
nand U6801 (N_6801,N_5488,N_5507);
nor U6802 (N_6802,N_5445,N_5216);
xor U6803 (N_6803,N_5416,N_5286);
and U6804 (N_6804,N_5460,N_5562);
or U6805 (N_6805,N_5073,N_5362);
xnor U6806 (N_6806,N_5450,N_5309);
nand U6807 (N_6807,N_5381,N_5628);
xor U6808 (N_6808,N_5297,N_5367);
nor U6809 (N_6809,N_5700,N_5209);
nand U6810 (N_6810,N_5153,N_5126);
xor U6811 (N_6811,N_5068,N_5805);
nand U6812 (N_6812,N_5497,N_5946);
nand U6813 (N_6813,N_5382,N_5070);
or U6814 (N_6814,N_5212,N_5160);
or U6815 (N_6815,N_5551,N_5279);
or U6816 (N_6816,N_5214,N_5635);
nor U6817 (N_6817,N_5593,N_5694);
xor U6818 (N_6818,N_5203,N_5910);
nand U6819 (N_6819,N_5315,N_5154);
nor U6820 (N_6820,N_5833,N_5304);
nand U6821 (N_6821,N_5011,N_5598);
xnor U6822 (N_6822,N_5655,N_5868);
nor U6823 (N_6823,N_5144,N_5333);
and U6824 (N_6824,N_5639,N_5047);
nor U6825 (N_6825,N_5817,N_5182);
nor U6826 (N_6826,N_5788,N_5512);
or U6827 (N_6827,N_5579,N_5857);
nor U6828 (N_6828,N_5045,N_5811);
and U6829 (N_6829,N_5155,N_5829);
nand U6830 (N_6830,N_5809,N_5469);
xor U6831 (N_6831,N_5240,N_5387);
xnor U6832 (N_6832,N_5763,N_5692);
nand U6833 (N_6833,N_5591,N_5483);
nand U6834 (N_6834,N_5761,N_5158);
nor U6835 (N_6835,N_5736,N_5147);
xnor U6836 (N_6836,N_5368,N_5369);
nand U6837 (N_6837,N_5968,N_5280);
and U6838 (N_6838,N_5760,N_5619);
xor U6839 (N_6839,N_5087,N_5446);
nor U6840 (N_6840,N_5650,N_5543);
nand U6841 (N_6841,N_5072,N_5992);
and U6842 (N_6842,N_5859,N_5107);
nand U6843 (N_6843,N_5615,N_5116);
and U6844 (N_6844,N_5187,N_5981);
xor U6845 (N_6845,N_5419,N_5059);
or U6846 (N_6846,N_5608,N_5669);
nand U6847 (N_6847,N_5146,N_5223);
or U6848 (N_6848,N_5419,N_5436);
or U6849 (N_6849,N_5863,N_5353);
or U6850 (N_6850,N_5139,N_5752);
xor U6851 (N_6851,N_5799,N_5159);
nand U6852 (N_6852,N_5206,N_5154);
xnor U6853 (N_6853,N_5894,N_5256);
and U6854 (N_6854,N_5665,N_5129);
or U6855 (N_6855,N_5069,N_5886);
xnor U6856 (N_6856,N_5090,N_5487);
or U6857 (N_6857,N_5814,N_5088);
nor U6858 (N_6858,N_5320,N_5398);
or U6859 (N_6859,N_5778,N_5615);
nor U6860 (N_6860,N_5821,N_5516);
xnor U6861 (N_6861,N_5441,N_5510);
nand U6862 (N_6862,N_5791,N_5403);
and U6863 (N_6863,N_5081,N_5508);
or U6864 (N_6864,N_5447,N_5053);
or U6865 (N_6865,N_5846,N_5771);
xnor U6866 (N_6866,N_5568,N_5500);
or U6867 (N_6867,N_5576,N_5788);
xnor U6868 (N_6868,N_5991,N_5773);
and U6869 (N_6869,N_5372,N_5221);
and U6870 (N_6870,N_5963,N_5270);
xnor U6871 (N_6871,N_5274,N_5022);
nor U6872 (N_6872,N_5275,N_5538);
xnor U6873 (N_6873,N_5197,N_5987);
or U6874 (N_6874,N_5503,N_5892);
xnor U6875 (N_6875,N_5815,N_5716);
nand U6876 (N_6876,N_5340,N_5342);
and U6877 (N_6877,N_5535,N_5301);
nor U6878 (N_6878,N_5490,N_5823);
and U6879 (N_6879,N_5833,N_5412);
nor U6880 (N_6880,N_5252,N_5686);
nand U6881 (N_6881,N_5167,N_5569);
and U6882 (N_6882,N_5885,N_5092);
nor U6883 (N_6883,N_5833,N_5151);
or U6884 (N_6884,N_5532,N_5549);
nand U6885 (N_6885,N_5517,N_5910);
xor U6886 (N_6886,N_5669,N_5900);
nor U6887 (N_6887,N_5942,N_5521);
and U6888 (N_6888,N_5927,N_5424);
and U6889 (N_6889,N_5395,N_5895);
and U6890 (N_6890,N_5164,N_5159);
and U6891 (N_6891,N_5170,N_5008);
xnor U6892 (N_6892,N_5071,N_5947);
or U6893 (N_6893,N_5648,N_5610);
nor U6894 (N_6894,N_5596,N_5739);
xor U6895 (N_6895,N_5231,N_5302);
or U6896 (N_6896,N_5721,N_5191);
and U6897 (N_6897,N_5647,N_5864);
and U6898 (N_6898,N_5725,N_5428);
nand U6899 (N_6899,N_5895,N_5530);
nand U6900 (N_6900,N_5145,N_5905);
nand U6901 (N_6901,N_5235,N_5945);
nand U6902 (N_6902,N_5015,N_5038);
xnor U6903 (N_6903,N_5530,N_5790);
and U6904 (N_6904,N_5813,N_5553);
nor U6905 (N_6905,N_5013,N_5146);
nand U6906 (N_6906,N_5432,N_5724);
xnor U6907 (N_6907,N_5225,N_5019);
xnor U6908 (N_6908,N_5613,N_5513);
nor U6909 (N_6909,N_5188,N_5161);
and U6910 (N_6910,N_5178,N_5020);
nor U6911 (N_6911,N_5818,N_5045);
nor U6912 (N_6912,N_5893,N_5192);
nand U6913 (N_6913,N_5963,N_5877);
nand U6914 (N_6914,N_5802,N_5947);
nor U6915 (N_6915,N_5680,N_5848);
nor U6916 (N_6916,N_5106,N_5643);
nor U6917 (N_6917,N_5085,N_5796);
nand U6918 (N_6918,N_5782,N_5445);
or U6919 (N_6919,N_5916,N_5556);
and U6920 (N_6920,N_5315,N_5426);
nand U6921 (N_6921,N_5055,N_5709);
xor U6922 (N_6922,N_5985,N_5475);
xor U6923 (N_6923,N_5608,N_5407);
xnor U6924 (N_6924,N_5576,N_5627);
nor U6925 (N_6925,N_5621,N_5542);
xor U6926 (N_6926,N_5055,N_5396);
and U6927 (N_6927,N_5826,N_5020);
nand U6928 (N_6928,N_5116,N_5172);
and U6929 (N_6929,N_5799,N_5850);
nand U6930 (N_6930,N_5416,N_5484);
or U6931 (N_6931,N_5213,N_5426);
nand U6932 (N_6932,N_5387,N_5381);
nor U6933 (N_6933,N_5763,N_5526);
and U6934 (N_6934,N_5029,N_5065);
or U6935 (N_6935,N_5255,N_5308);
nand U6936 (N_6936,N_5076,N_5155);
and U6937 (N_6937,N_5676,N_5765);
or U6938 (N_6938,N_5831,N_5707);
xnor U6939 (N_6939,N_5294,N_5828);
nor U6940 (N_6940,N_5303,N_5135);
nand U6941 (N_6941,N_5790,N_5285);
nor U6942 (N_6942,N_5057,N_5564);
nand U6943 (N_6943,N_5856,N_5846);
or U6944 (N_6944,N_5268,N_5187);
nor U6945 (N_6945,N_5963,N_5237);
nor U6946 (N_6946,N_5313,N_5151);
and U6947 (N_6947,N_5079,N_5460);
nor U6948 (N_6948,N_5209,N_5041);
nand U6949 (N_6949,N_5473,N_5607);
nor U6950 (N_6950,N_5458,N_5103);
xor U6951 (N_6951,N_5698,N_5840);
nand U6952 (N_6952,N_5846,N_5893);
nand U6953 (N_6953,N_5689,N_5821);
nand U6954 (N_6954,N_5568,N_5130);
nand U6955 (N_6955,N_5628,N_5073);
nor U6956 (N_6956,N_5071,N_5172);
or U6957 (N_6957,N_5332,N_5411);
and U6958 (N_6958,N_5646,N_5415);
nor U6959 (N_6959,N_5023,N_5910);
nand U6960 (N_6960,N_5197,N_5867);
nand U6961 (N_6961,N_5878,N_5929);
and U6962 (N_6962,N_5537,N_5651);
and U6963 (N_6963,N_5062,N_5304);
nor U6964 (N_6964,N_5510,N_5149);
or U6965 (N_6965,N_5214,N_5333);
nor U6966 (N_6966,N_5518,N_5026);
or U6967 (N_6967,N_5057,N_5438);
nand U6968 (N_6968,N_5066,N_5418);
or U6969 (N_6969,N_5859,N_5230);
nand U6970 (N_6970,N_5717,N_5132);
or U6971 (N_6971,N_5170,N_5117);
nand U6972 (N_6972,N_5997,N_5691);
nand U6973 (N_6973,N_5133,N_5563);
nand U6974 (N_6974,N_5396,N_5143);
and U6975 (N_6975,N_5651,N_5993);
or U6976 (N_6976,N_5711,N_5167);
nor U6977 (N_6977,N_5806,N_5558);
nand U6978 (N_6978,N_5736,N_5221);
or U6979 (N_6979,N_5781,N_5189);
nor U6980 (N_6980,N_5918,N_5747);
nor U6981 (N_6981,N_5744,N_5546);
nand U6982 (N_6982,N_5119,N_5218);
nand U6983 (N_6983,N_5803,N_5984);
and U6984 (N_6984,N_5104,N_5177);
or U6985 (N_6985,N_5911,N_5789);
or U6986 (N_6986,N_5736,N_5117);
or U6987 (N_6987,N_5331,N_5209);
xor U6988 (N_6988,N_5974,N_5776);
or U6989 (N_6989,N_5561,N_5102);
and U6990 (N_6990,N_5309,N_5711);
nand U6991 (N_6991,N_5312,N_5226);
or U6992 (N_6992,N_5581,N_5725);
xnor U6993 (N_6993,N_5812,N_5278);
nand U6994 (N_6994,N_5942,N_5492);
xor U6995 (N_6995,N_5844,N_5991);
or U6996 (N_6996,N_5792,N_5806);
nand U6997 (N_6997,N_5126,N_5402);
and U6998 (N_6998,N_5855,N_5227);
and U6999 (N_6999,N_5488,N_5892);
or U7000 (N_7000,N_6908,N_6965);
or U7001 (N_7001,N_6317,N_6637);
xnor U7002 (N_7002,N_6935,N_6680);
and U7003 (N_7003,N_6944,N_6755);
or U7004 (N_7004,N_6600,N_6806);
and U7005 (N_7005,N_6252,N_6159);
or U7006 (N_7006,N_6256,N_6595);
and U7007 (N_7007,N_6464,N_6423);
or U7008 (N_7008,N_6791,N_6892);
nand U7009 (N_7009,N_6591,N_6724);
nand U7010 (N_7010,N_6112,N_6067);
or U7011 (N_7011,N_6707,N_6047);
and U7012 (N_7012,N_6108,N_6874);
and U7013 (N_7013,N_6174,N_6436);
or U7014 (N_7014,N_6150,N_6635);
nor U7015 (N_7015,N_6456,N_6249);
nor U7016 (N_7016,N_6016,N_6924);
nand U7017 (N_7017,N_6206,N_6381);
and U7018 (N_7018,N_6620,N_6147);
nor U7019 (N_7019,N_6702,N_6109);
and U7020 (N_7020,N_6862,N_6066);
nor U7021 (N_7021,N_6043,N_6575);
nand U7022 (N_7022,N_6838,N_6449);
and U7023 (N_7023,N_6093,N_6795);
nand U7024 (N_7024,N_6408,N_6647);
and U7025 (N_7025,N_6484,N_6192);
nand U7026 (N_7026,N_6071,N_6049);
xnor U7027 (N_7027,N_6075,N_6401);
and U7028 (N_7028,N_6937,N_6783);
nand U7029 (N_7029,N_6120,N_6297);
xnor U7030 (N_7030,N_6288,N_6846);
and U7031 (N_7031,N_6726,N_6732);
and U7032 (N_7032,N_6887,N_6185);
xor U7033 (N_7033,N_6366,N_6094);
nand U7034 (N_7034,N_6718,N_6845);
or U7035 (N_7035,N_6352,N_6660);
and U7036 (N_7036,N_6590,N_6648);
and U7037 (N_7037,N_6546,N_6662);
nand U7038 (N_7038,N_6440,N_6764);
or U7039 (N_7039,N_6385,N_6750);
nand U7040 (N_7040,N_6902,N_6947);
nand U7041 (N_7041,N_6765,N_6044);
or U7042 (N_7042,N_6645,N_6952);
nor U7043 (N_7043,N_6746,N_6835);
nand U7044 (N_7044,N_6447,N_6751);
or U7045 (N_7045,N_6657,N_6936);
nor U7046 (N_7046,N_6189,N_6499);
and U7047 (N_7047,N_6998,N_6850);
or U7048 (N_7048,N_6302,N_6968);
xnor U7049 (N_7049,N_6267,N_6020);
nand U7050 (N_7050,N_6674,N_6097);
xnor U7051 (N_7051,N_6646,N_6177);
nand U7052 (N_7052,N_6954,N_6217);
nand U7053 (N_7053,N_6226,N_6325);
or U7054 (N_7054,N_6743,N_6781);
nor U7055 (N_7055,N_6530,N_6091);
xnor U7056 (N_7056,N_6276,N_6540);
nand U7057 (N_7057,N_6753,N_6913);
nor U7058 (N_7058,N_6733,N_6344);
xnor U7059 (N_7059,N_6475,N_6809);
xor U7060 (N_7060,N_6455,N_6052);
nand U7061 (N_7061,N_6428,N_6294);
nor U7062 (N_7062,N_6742,N_6322);
or U7063 (N_7063,N_6496,N_6019);
or U7064 (N_7064,N_6115,N_6639);
or U7065 (N_7065,N_6670,N_6446);
or U7066 (N_7066,N_6383,N_6962);
nand U7067 (N_7067,N_6190,N_6992);
and U7068 (N_7068,N_6898,N_6196);
and U7069 (N_7069,N_6041,N_6508);
nor U7070 (N_7070,N_6506,N_6321);
xnor U7071 (N_7071,N_6134,N_6896);
nand U7072 (N_7072,N_6543,N_6841);
xnor U7073 (N_7073,N_6000,N_6013);
or U7074 (N_7074,N_6882,N_6730);
or U7075 (N_7075,N_6495,N_6258);
or U7076 (N_7076,N_6933,N_6232);
xor U7077 (N_7077,N_6945,N_6878);
or U7078 (N_7078,N_6659,N_6153);
nor U7079 (N_7079,N_6415,N_6972);
nand U7080 (N_7080,N_6342,N_6981);
nor U7081 (N_7081,N_6144,N_6246);
nand U7082 (N_7082,N_6711,N_6914);
and U7083 (N_7083,N_6717,N_6710);
and U7084 (N_7084,N_6400,N_6176);
xor U7085 (N_7085,N_6950,N_6823);
nor U7086 (N_7086,N_6092,N_6168);
nand U7087 (N_7087,N_6550,N_6099);
nor U7088 (N_7088,N_6796,N_6934);
nor U7089 (N_7089,N_6787,N_6187);
or U7090 (N_7090,N_6327,N_6493);
and U7091 (N_7091,N_6445,N_6334);
nand U7092 (N_7092,N_6319,N_6920);
nand U7093 (N_7093,N_6769,N_6122);
nand U7094 (N_7094,N_6009,N_6866);
xor U7095 (N_7095,N_6669,N_6369);
or U7096 (N_7096,N_6471,N_6556);
and U7097 (N_7097,N_6214,N_6259);
xor U7098 (N_7098,N_6608,N_6429);
xor U7099 (N_7099,N_6613,N_6046);
xnor U7100 (N_7100,N_6404,N_6227);
and U7101 (N_7101,N_6465,N_6593);
nand U7102 (N_7102,N_6215,N_6301);
xnor U7103 (N_7103,N_6008,N_6739);
nand U7104 (N_7104,N_6967,N_6272);
nand U7105 (N_7105,N_6048,N_6572);
xnor U7106 (N_7106,N_6129,N_6700);
and U7107 (N_7107,N_6209,N_6736);
nand U7108 (N_7108,N_6064,N_6966);
nor U7109 (N_7109,N_6494,N_6164);
nand U7110 (N_7110,N_6566,N_6855);
or U7111 (N_7111,N_6194,N_6228);
xnor U7112 (N_7112,N_6712,N_6157);
xnor U7113 (N_7113,N_6513,N_6116);
nor U7114 (N_7114,N_6254,N_6814);
xnor U7115 (N_7115,N_6413,N_6457);
nand U7116 (N_7116,N_6666,N_6949);
nand U7117 (N_7117,N_6314,N_6958);
nor U7118 (N_7118,N_6792,N_6812);
and U7119 (N_7119,N_6713,N_6738);
and U7120 (N_7120,N_6087,N_6433);
nor U7121 (N_7121,N_6481,N_6123);
or U7122 (N_7122,N_6316,N_6070);
or U7123 (N_7123,N_6017,N_6309);
nor U7124 (N_7124,N_6126,N_6402);
xor U7125 (N_7125,N_6247,N_6368);
or U7126 (N_7126,N_6721,N_6725);
nand U7127 (N_7127,N_6901,N_6875);
and U7128 (N_7128,N_6022,N_6643);
nor U7129 (N_7129,N_6354,N_6173);
xor U7130 (N_7130,N_6837,N_6586);
or U7131 (N_7131,N_6458,N_6472);
nor U7132 (N_7132,N_6679,N_6610);
and U7133 (N_7133,N_6904,N_6351);
or U7134 (N_7134,N_6957,N_6592);
and U7135 (N_7135,N_6754,N_6040);
or U7136 (N_7136,N_6876,N_6060);
or U7137 (N_7137,N_6827,N_6925);
nor U7138 (N_7138,N_6890,N_6438);
or U7139 (N_7139,N_6452,N_6531);
xor U7140 (N_7140,N_6237,N_6558);
and U7141 (N_7141,N_6379,N_6089);
nand U7142 (N_7142,N_6698,N_6574);
nand U7143 (N_7143,N_6629,N_6163);
and U7144 (N_7144,N_6104,N_6262);
nand U7145 (N_7145,N_6539,N_6030);
and U7146 (N_7146,N_6058,N_6828);
nor U7147 (N_7147,N_6996,N_6544);
and U7148 (N_7148,N_6160,N_6004);
nor U7149 (N_7149,N_6807,N_6218);
or U7150 (N_7150,N_6326,N_6435);
or U7151 (N_7151,N_6195,N_6220);
and U7152 (N_7152,N_6273,N_6365);
or U7153 (N_7153,N_6772,N_6025);
nor U7154 (N_7154,N_6729,N_6392);
nor U7155 (N_7155,N_6308,N_6984);
and U7156 (N_7156,N_6375,N_6072);
xor U7157 (N_7157,N_6037,N_6377);
or U7158 (N_7158,N_6561,N_6614);
xor U7159 (N_7159,N_6480,N_6239);
nor U7160 (N_7160,N_6527,N_6830);
nand U7161 (N_7161,N_6555,N_6167);
or U7162 (N_7162,N_6100,N_6356);
xnor U7163 (N_7163,N_6861,N_6175);
nand U7164 (N_7164,N_6650,N_6976);
nand U7165 (N_7165,N_6582,N_6589);
xnor U7166 (N_7166,N_6774,N_6995);
or U7167 (N_7167,N_6503,N_6641);
and U7168 (N_7168,N_6251,N_6961);
xnor U7169 (N_7169,N_6763,N_6983);
or U7170 (N_7170,N_6205,N_6955);
nor U7171 (N_7171,N_6820,N_6619);
and U7172 (N_7172,N_6021,N_6844);
nor U7173 (N_7173,N_6031,N_6490);
nor U7174 (N_7174,N_6672,N_6014);
xnor U7175 (N_7175,N_6790,N_6709);
or U7176 (N_7176,N_6974,N_6923);
xnor U7177 (N_7177,N_6241,N_6811);
nor U7178 (N_7178,N_6797,N_6510);
or U7179 (N_7179,N_6001,N_6242);
or U7180 (N_7180,N_6303,N_6181);
nand U7181 (N_7181,N_6997,N_6825);
nor U7182 (N_7182,N_6675,N_6015);
nor U7183 (N_7183,N_6912,N_6624);
nand U7184 (N_7184,N_6893,N_6604);
and U7185 (N_7185,N_6534,N_6114);
xor U7186 (N_7186,N_6842,N_6979);
nor U7187 (N_7187,N_6565,N_6621);
xor U7188 (N_7188,N_6424,N_6005);
and U7189 (N_7189,N_6758,N_6722);
or U7190 (N_7190,N_6441,N_6526);
or U7191 (N_7191,N_6581,N_6879);
or U7192 (N_7192,N_6171,N_6061);
nand U7193 (N_7193,N_6461,N_6155);
or U7194 (N_7194,N_6599,N_6389);
nor U7195 (N_7195,N_6360,N_6833);
and U7196 (N_7196,N_6138,N_6193);
nor U7197 (N_7197,N_6113,N_6601);
xor U7198 (N_7198,N_6329,N_6474);
nor U7199 (N_7199,N_6971,N_6466);
nand U7200 (N_7200,N_6263,N_6250);
nand U7201 (N_7201,N_6393,N_6364);
nor U7202 (N_7202,N_6607,N_6065);
and U7203 (N_7203,N_6468,N_6524);
xor U7204 (N_7204,N_6261,N_6623);
nor U7205 (N_7205,N_6024,N_6376);
and U7206 (N_7206,N_6012,N_6859);
xnor U7207 (N_7207,N_6305,N_6767);
nand U7208 (N_7208,N_6172,N_6491);
nand U7209 (N_7209,N_6895,N_6940);
xor U7210 (N_7210,N_6824,N_6361);
xnor U7211 (N_7211,N_6692,N_6202);
nor U7212 (N_7212,N_6110,N_6340);
and U7213 (N_7213,N_6422,N_6459);
nand U7214 (N_7214,N_6057,N_6941);
xor U7215 (N_7215,N_6023,N_6689);
and U7216 (N_7216,N_6785,N_6333);
nand U7217 (N_7217,N_6870,N_6911);
or U7218 (N_7218,N_6201,N_6084);
nor U7219 (N_7219,N_6849,N_6028);
or U7220 (N_7220,N_6124,N_6985);
or U7221 (N_7221,N_6492,N_6860);
or U7222 (N_7222,N_6213,N_6264);
nand U7223 (N_7223,N_6567,N_6951);
nand U7224 (N_7224,N_6118,N_6625);
or U7225 (N_7225,N_6691,N_6542);
and U7226 (N_7226,N_6602,N_6324);
nor U7227 (N_7227,N_6018,N_6290);
nand U7228 (N_7228,N_6617,N_6969);
or U7229 (N_7229,N_6872,N_6665);
nor U7230 (N_7230,N_6839,N_6397);
or U7231 (N_7231,N_6255,N_6180);
nor U7232 (N_7232,N_6603,N_6834);
xor U7233 (N_7233,N_6654,N_6311);
xnor U7234 (N_7234,N_6162,N_6088);
nand U7235 (N_7235,N_6585,N_6002);
and U7236 (N_7236,N_6338,N_6685);
and U7237 (N_7237,N_6386,N_6131);
nor U7238 (N_7238,N_6773,N_6989);
nor U7239 (N_7239,N_6432,N_6973);
or U7240 (N_7240,N_6128,N_6328);
and U7241 (N_7241,N_6341,N_6136);
xor U7242 (N_7242,N_6502,N_6483);
or U7243 (N_7243,N_6384,N_6339);
or U7244 (N_7244,N_6442,N_6234);
xor U7245 (N_7245,N_6676,N_6050);
and U7246 (N_7246,N_6551,N_6299);
or U7247 (N_7247,N_6596,N_6740);
xnor U7248 (N_7248,N_6805,N_6749);
or U7249 (N_7249,N_6421,N_6082);
nor U7250 (N_7250,N_6414,N_6125);
nor U7251 (N_7251,N_6628,N_6038);
and U7252 (N_7252,N_6557,N_6467);
and U7253 (N_7253,N_6832,N_6248);
nand U7254 (N_7254,N_6735,N_6518);
nand U7255 (N_7255,N_6517,N_6371);
or U7256 (N_7256,N_6885,N_6668);
xnor U7257 (N_7257,N_6430,N_6525);
nor U7258 (N_7258,N_6938,N_6287);
xnor U7259 (N_7259,N_6053,N_6265);
nand U7260 (N_7260,N_6417,N_6096);
xnor U7261 (N_7261,N_6528,N_6269);
or U7262 (N_7262,N_6652,N_6387);
and U7263 (N_7263,N_6813,N_6587);
and U7264 (N_7264,N_6487,N_6877);
xnor U7265 (N_7265,N_6549,N_6188);
nand U7266 (N_7266,N_6293,N_6501);
and U7267 (N_7267,N_6410,N_6395);
nand U7268 (N_7268,N_6516,N_6426);
xor U7269 (N_7269,N_6956,N_6627);
and U7270 (N_7270,N_6815,N_6800);
nor U7271 (N_7271,N_6407,N_6137);
nor U7272 (N_7272,N_6651,N_6683);
or U7273 (N_7273,N_6026,N_6987);
or U7274 (N_7274,N_6488,N_6761);
nor U7275 (N_7275,N_6768,N_6045);
and U7276 (N_7276,N_6822,N_6148);
nor U7277 (N_7277,N_6318,N_6076);
nor U7278 (N_7278,N_6391,N_6611);
nand U7279 (N_7279,N_6946,N_6856);
and U7280 (N_7280,N_6681,N_6538);
nor U7281 (N_7281,N_6444,N_6152);
xnor U7282 (N_7282,N_6451,N_6708);
or U7283 (N_7283,N_6682,N_6078);
or U7284 (N_7284,N_6982,N_6106);
xor U7285 (N_7285,N_6253,N_6900);
xor U7286 (N_7286,N_6584,N_6184);
nand U7287 (N_7287,N_6673,N_6035);
and U7288 (N_7288,N_6541,N_6664);
xor U7289 (N_7289,N_6922,N_6081);
and U7290 (N_7290,N_6706,N_6817);
and U7291 (N_7291,N_6266,N_6649);
nand U7292 (N_7292,N_6868,N_6888);
xor U7293 (N_7293,N_6759,N_6918);
and U7294 (N_7294,N_6169,N_6597);
and U7295 (N_7295,N_6776,N_6240);
nor U7296 (N_7296,N_6003,N_6310);
and U7297 (N_7297,N_6609,N_6348);
nand U7298 (N_7298,N_6042,N_6409);
or U7299 (N_7299,N_6644,N_6335);
and U7300 (N_7300,N_6212,N_6286);
or U7301 (N_7301,N_6068,N_6362);
nand U7302 (N_7302,N_6548,N_6851);
or U7303 (N_7303,N_6396,N_6616);
xnor U7304 (N_7304,N_6762,N_6357);
nor U7305 (N_7305,N_6705,N_6151);
or U7306 (N_7306,N_6964,N_6270);
nand U7307 (N_7307,N_6080,N_6208);
xnor U7308 (N_7308,N_6915,N_6994);
or U7309 (N_7309,N_6006,N_6268);
and U7310 (N_7310,N_6370,N_6752);
and U7311 (N_7311,N_6577,N_6568);
nand U7312 (N_7312,N_6304,N_6704);
and U7313 (N_7313,N_6942,N_6988);
xnor U7314 (N_7314,N_6478,N_6281);
nand U7315 (N_7315,N_6010,N_6307);
xnor U7316 (N_7316,N_6063,N_6418);
and U7317 (N_7317,N_6186,N_6497);
nor U7318 (N_7318,N_6355,N_6182);
or U7319 (N_7319,N_6142,N_6831);
xnor U7320 (N_7320,N_6963,N_6880);
xor U7321 (N_7321,N_6374,N_6747);
xnor U7322 (N_7322,N_6867,N_6032);
nor U7323 (N_7323,N_6990,N_6529);
xnor U7324 (N_7324,N_6786,N_6883);
nor U7325 (N_7325,N_6696,N_6521);
nor U7326 (N_7326,N_6460,N_6658);
nand U7327 (N_7327,N_6522,N_6836);
and U7328 (N_7328,N_6622,N_6229);
and U7329 (N_7329,N_6479,N_6580);
nand U7330 (N_7330,N_6107,N_6978);
nand U7331 (N_7331,N_6378,N_6233);
xor U7332 (N_7332,N_6086,N_6916);
or U7333 (N_7333,N_6715,N_6779);
xnor U7334 (N_7334,N_6312,N_6511);
nand U7335 (N_7335,N_6298,N_6406);
xnor U7336 (N_7336,N_6257,N_6211);
nor U7337 (N_7337,N_6881,N_6179);
nor U7338 (N_7338,N_6403,N_6055);
nand U7339 (N_7339,N_6011,N_6007);
or U7340 (N_7340,N_6507,N_6728);
or U7341 (N_7341,N_6291,N_6380);
nor U7342 (N_7342,N_6808,N_6139);
or U7343 (N_7343,N_6230,N_6083);
or U7344 (N_7344,N_6336,N_6745);
xor U7345 (N_7345,N_6631,N_6578);
xnor U7346 (N_7346,N_6295,N_6198);
nor U7347 (N_7347,N_6903,N_6149);
nor U7348 (N_7348,N_6993,N_6894);
or U7349 (N_7349,N_6489,N_6509);
and U7350 (N_7350,N_6802,N_6358);
xor U7351 (N_7351,N_6416,N_6606);
xor U7352 (N_7352,N_6183,N_6929);
and U7353 (N_7353,N_6277,N_6448);
and U7354 (N_7354,N_6090,N_6798);
and U7355 (N_7355,N_6353,N_6111);
xor U7356 (N_7356,N_6615,N_6437);
xor U7357 (N_7357,N_6686,N_6821);
or U7358 (N_7358,N_6141,N_6425);
nand U7359 (N_7359,N_6170,N_6210);
nand U7360 (N_7360,N_6583,N_6694);
nand U7361 (N_7361,N_6737,N_6547);
nor U7362 (N_7362,N_6146,N_6970);
and U7363 (N_7363,N_6482,N_6642);
nand U7364 (N_7364,N_6036,N_6275);
or U7365 (N_7365,N_6485,N_6103);
or U7366 (N_7366,N_6419,N_6236);
xor U7367 (N_7367,N_6778,N_6165);
nand U7368 (N_7368,N_6079,N_6858);
and U7369 (N_7369,N_6863,N_6626);
nor U7370 (N_7370,N_6843,N_6382);
xnor U7371 (N_7371,N_6315,N_6770);
or U7372 (N_7372,N_6537,N_6282);
or U7373 (N_7373,N_6411,N_6907);
and U7374 (N_7374,N_6390,N_6562);
xnor U7375 (N_7375,N_6656,N_6102);
nor U7376 (N_7376,N_6598,N_6098);
xor U7377 (N_7377,N_6279,N_6869);
or U7378 (N_7378,N_6033,N_6127);
xor U7379 (N_7379,N_6801,N_6051);
nor U7380 (N_7380,N_6323,N_6532);
or U7381 (N_7381,N_6101,N_6731);
or U7382 (N_7382,N_6074,N_6693);
nor U7383 (N_7383,N_6612,N_6405);
nor U7384 (N_7384,N_6221,N_6135);
xnor U7385 (N_7385,N_6453,N_6771);
and U7386 (N_7386,N_6454,N_6799);
xnor U7387 (N_7387,N_6630,N_6161);
and U7388 (N_7388,N_6166,N_6156);
nor U7389 (N_7389,N_6520,N_6523);
nor U7390 (N_7390,N_6931,N_6140);
nand U7391 (N_7391,N_6278,N_6703);
or U7392 (N_7392,N_6238,N_6948);
or U7393 (N_7393,N_6677,N_6741);
xor U7394 (N_7394,N_6756,N_6243);
nand U7395 (N_7395,N_6848,N_6977);
nor U7396 (N_7396,N_6618,N_6347);
nand U7397 (N_7397,N_6399,N_6563);
xor U7398 (N_7398,N_6498,N_6039);
nor U7399 (N_7399,N_6191,N_6274);
xor U7400 (N_7400,N_6930,N_6363);
xnor U7401 (N_7401,N_6204,N_6200);
and U7402 (N_7402,N_6062,N_6300);
and U7403 (N_7403,N_6671,N_6701);
nand U7404 (N_7404,N_6853,N_6143);
nor U7405 (N_7405,N_6943,N_6780);
nand U7406 (N_7406,N_6225,N_6980);
xnor U7407 (N_7407,N_6678,N_6054);
nand U7408 (N_7408,N_6926,N_6512);
xor U7409 (N_7409,N_6343,N_6871);
or U7410 (N_7410,N_6450,N_6789);
or U7411 (N_7411,N_6533,N_6991);
and U7412 (N_7412,N_6223,N_6222);
and U7413 (N_7413,N_6245,N_6349);
nor U7414 (N_7414,N_6463,N_6847);
and U7415 (N_7415,N_6119,N_6899);
or U7416 (N_7416,N_6398,N_6766);
nand U7417 (N_7417,N_6133,N_6029);
or U7418 (N_7418,N_6697,N_6292);
nor U7419 (N_7419,N_6178,N_6760);
nand U7420 (N_7420,N_6373,N_6331);
xnor U7421 (N_7421,N_6552,N_6588);
xnor U7422 (N_7422,N_6158,N_6999);
nand U7423 (N_7423,N_6219,N_6431);
xnor U7424 (N_7424,N_6788,N_6632);
nor U7425 (N_7425,N_6897,N_6727);
nor U7426 (N_7426,N_6313,N_6959);
or U7427 (N_7427,N_6695,N_6564);
nand U7428 (N_7428,N_6891,N_6285);
nor U7429 (N_7429,N_6594,N_6854);
and U7430 (N_7430,N_6203,N_6289);
xor U7431 (N_7431,N_6804,N_6576);
nor U7432 (N_7432,N_6284,N_6427);
and U7433 (N_7433,N_6154,N_6554);
xor U7434 (N_7434,N_6921,N_6818);
nand U7435 (N_7435,N_6653,N_6332);
nor U7436 (N_7436,N_6816,N_6077);
or U7437 (N_7437,N_6462,N_6553);
and U7438 (N_7438,N_6909,N_6346);
nor U7439 (N_7439,N_6939,N_6634);
nor U7440 (N_7440,N_6231,N_6829);
or U7441 (N_7441,N_6199,N_6235);
and U7442 (N_7442,N_6056,N_6121);
xor U7443 (N_7443,N_6296,N_6699);
nand U7444 (N_7444,N_6476,N_6953);
and U7445 (N_7445,N_6640,N_6687);
xnor U7446 (N_7446,N_6784,N_6350);
nor U7447 (N_7447,N_6864,N_6757);
or U7448 (N_7448,N_6690,N_6477);
xnor U7449 (N_7449,N_6744,N_6873);
nand U7450 (N_7450,N_6059,N_6782);
and U7451 (N_7451,N_6857,N_6069);
xnor U7452 (N_7452,N_6545,N_6280);
or U7453 (N_7453,N_6986,N_6519);
xor U7454 (N_7454,N_6720,N_6330);
and U7455 (N_7455,N_6271,N_6810);
xor U7456 (N_7456,N_6095,N_6105);
nand U7457 (N_7457,N_6573,N_6579);
and U7458 (N_7458,N_6714,N_6748);
nand U7459 (N_7459,N_6536,N_6337);
xor U7460 (N_7460,N_6073,N_6917);
xnor U7461 (N_7461,N_6840,N_6283);
xnor U7462 (N_7462,N_6723,N_6306);
nor U7463 (N_7463,N_6367,N_6775);
or U7464 (N_7464,N_6505,N_6826);
and U7465 (N_7465,N_6412,N_6473);
or U7466 (N_7466,N_6372,N_6569);
and U7467 (N_7467,N_6469,N_6655);
nand U7468 (N_7468,N_6320,N_6927);
and U7469 (N_7469,N_6865,N_6638);
nand U7470 (N_7470,N_6734,N_6719);
xor U7471 (N_7471,N_6515,N_6928);
or U7472 (N_7472,N_6684,N_6688);
or U7473 (N_7473,N_6439,N_6117);
nor U7474 (N_7474,N_6906,N_6884);
or U7475 (N_7475,N_6420,N_6636);
xor U7476 (N_7476,N_6932,N_6975);
xnor U7477 (N_7477,N_6504,N_6661);
and U7478 (N_7478,N_6605,N_6027);
nand U7479 (N_7479,N_6819,N_6889);
nand U7480 (N_7480,N_6197,N_6434);
or U7481 (N_7481,N_6571,N_6560);
nand U7482 (N_7482,N_6905,N_6244);
xnor U7483 (N_7483,N_6886,N_6663);
xor U7484 (N_7484,N_6345,N_6145);
nor U7485 (N_7485,N_6514,N_6443);
nor U7486 (N_7486,N_6132,N_6486);
nor U7487 (N_7487,N_6803,N_6130);
xnor U7488 (N_7488,N_6960,N_6535);
nor U7489 (N_7489,N_6793,N_6919);
nor U7490 (N_7490,N_6777,N_6224);
or U7491 (N_7491,N_6207,N_6910);
xor U7492 (N_7492,N_6794,N_6034);
nor U7493 (N_7493,N_6852,N_6388);
nand U7494 (N_7494,N_6716,N_6470);
nand U7495 (N_7495,N_6260,N_6559);
nand U7496 (N_7496,N_6394,N_6570);
nor U7497 (N_7497,N_6500,N_6216);
or U7498 (N_7498,N_6359,N_6085);
and U7499 (N_7499,N_6667,N_6633);
xor U7500 (N_7500,N_6846,N_6211);
xor U7501 (N_7501,N_6626,N_6008);
and U7502 (N_7502,N_6833,N_6565);
nor U7503 (N_7503,N_6857,N_6292);
or U7504 (N_7504,N_6996,N_6470);
nand U7505 (N_7505,N_6027,N_6937);
and U7506 (N_7506,N_6102,N_6535);
nor U7507 (N_7507,N_6801,N_6709);
xnor U7508 (N_7508,N_6705,N_6082);
and U7509 (N_7509,N_6993,N_6032);
and U7510 (N_7510,N_6492,N_6554);
nor U7511 (N_7511,N_6188,N_6710);
nor U7512 (N_7512,N_6681,N_6388);
and U7513 (N_7513,N_6704,N_6601);
xnor U7514 (N_7514,N_6949,N_6784);
and U7515 (N_7515,N_6535,N_6460);
or U7516 (N_7516,N_6082,N_6486);
nor U7517 (N_7517,N_6478,N_6606);
xnor U7518 (N_7518,N_6498,N_6690);
or U7519 (N_7519,N_6797,N_6811);
or U7520 (N_7520,N_6399,N_6356);
nor U7521 (N_7521,N_6666,N_6672);
xnor U7522 (N_7522,N_6156,N_6990);
or U7523 (N_7523,N_6850,N_6698);
and U7524 (N_7524,N_6262,N_6683);
nand U7525 (N_7525,N_6608,N_6915);
nor U7526 (N_7526,N_6782,N_6112);
and U7527 (N_7527,N_6895,N_6027);
xor U7528 (N_7528,N_6531,N_6550);
nor U7529 (N_7529,N_6593,N_6332);
or U7530 (N_7530,N_6142,N_6409);
and U7531 (N_7531,N_6709,N_6287);
nand U7532 (N_7532,N_6736,N_6883);
and U7533 (N_7533,N_6768,N_6596);
and U7534 (N_7534,N_6176,N_6079);
xor U7535 (N_7535,N_6862,N_6696);
or U7536 (N_7536,N_6741,N_6913);
or U7537 (N_7537,N_6723,N_6667);
or U7538 (N_7538,N_6897,N_6431);
nand U7539 (N_7539,N_6174,N_6431);
or U7540 (N_7540,N_6962,N_6236);
or U7541 (N_7541,N_6818,N_6851);
xnor U7542 (N_7542,N_6347,N_6432);
xnor U7543 (N_7543,N_6228,N_6659);
nor U7544 (N_7544,N_6378,N_6363);
xnor U7545 (N_7545,N_6597,N_6271);
and U7546 (N_7546,N_6598,N_6246);
nand U7547 (N_7547,N_6135,N_6042);
or U7548 (N_7548,N_6124,N_6341);
and U7549 (N_7549,N_6825,N_6883);
nand U7550 (N_7550,N_6390,N_6327);
and U7551 (N_7551,N_6191,N_6350);
nand U7552 (N_7552,N_6951,N_6063);
nand U7553 (N_7553,N_6811,N_6291);
nor U7554 (N_7554,N_6370,N_6960);
nor U7555 (N_7555,N_6671,N_6975);
and U7556 (N_7556,N_6147,N_6252);
and U7557 (N_7557,N_6680,N_6457);
nor U7558 (N_7558,N_6482,N_6038);
or U7559 (N_7559,N_6423,N_6035);
or U7560 (N_7560,N_6954,N_6562);
nand U7561 (N_7561,N_6334,N_6966);
or U7562 (N_7562,N_6248,N_6596);
nand U7563 (N_7563,N_6278,N_6247);
nand U7564 (N_7564,N_6253,N_6606);
and U7565 (N_7565,N_6576,N_6812);
and U7566 (N_7566,N_6601,N_6772);
and U7567 (N_7567,N_6786,N_6957);
nor U7568 (N_7568,N_6346,N_6402);
xnor U7569 (N_7569,N_6512,N_6190);
or U7570 (N_7570,N_6672,N_6728);
or U7571 (N_7571,N_6053,N_6459);
nand U7572 (N_7572,N_6889,N_6614);
xor U7573 (N_7573,N_6433,N_6673);
nand U7574 (N_7574,N_6244,N_6397);
nand U7575 (N_7575,N_6533,N_6157);
or U7576 (N_7576,N_6915,N_6056);
or U7577 (N_7577,N_6272,N_6644);
xnor U7578 (N_7578,N_6521,N_6519);
xnor U7579 (N_7579,N_6178,N_6662);
xor U7580 (N_7580,N_6006,N_6502);
xor U7581 (N_7581,N_6394,N_6715);
xor U7582 (N_7582,N_6530,N_6097);
or U7583 (N_7583,N_6277,N_6538);
xor U7584 (N_7584,N_6023,N_6814);
nand U7585 (N_7585,N_6406,N_6321);
or U7586 (N_7586,N_6780,N_6940);
or U7587 (N_7587,N_6591,N_6205);
xor U7588 (N_7588,N_6603,N_6479);
and U7589 (N_7589,N_6576,N_6993);
nor U7590 (N_7590,N_6365,N_6411);
or U7591 (N_7591,N_6393,N_6184);
xnor U7592 (N_7592,N_6532,N_6203);
xnor U7593 (N_7593,N_6449,N_6466);
and U7594 (N_7594,N_6394,N_6240);
or U7595 (N_7595,N_6773,N_6040);
nor U7596 (N_7596,N_6957,N_6425);
or U7597 (N_7597,N_6683,N_6797);
xor U7598 (N_7598,N_6375,N_6917);
and U7599 (N_7599,N_6389,N_6948);
nor U7600 (N_7600,N_6281,N_6307);
and U7601 (N_7601,N_6481,N_6135);
or U7602 (N_7602,N_6358,N_6673);
and U7603 (N_7603,N_6374,N_6067);
or U7604 (N_7604,N_6968,N_6595);
nand U7605 (N_7605,N_6613,N_6757);
nor U7606 (N_7606,N_6925,N_6338);
nand U7607 (N_7607,N_6178,N_6613);
and U7608 (N_7608,N_6820,N_6891);
and U7609 (N_7609,N_6673,N_6203);
nand U7610 (N_7610,N_6896,N_6741);
and U7611 (N_7611,N_6166,N_6785);
and U7612 (N_7612,N_6360,N_6051);
xnor U7613 (N_7613,N_6956,N_6080);
nand U7614 (N_7614,N_6079,N_6259);
nor U7615 (N_7615,N_6580,N_6213);
nand U7616 (N_7616,N_6479,N_6597);
or U7617 (N_7617,N_6049,N_6131);
nand U7618 (N_7618,N_6443,N_6813);
xor U7619 (N_7619,N_6727,N_6820);
or U7620 (N_7620,N_6984,N_6641);
nand U7621 (N_7621,N_6080,N_6638);
or U7622 (N_7622,N_6960,N_6176);
or U7623 (N_7623,N_6437,N_6050);
or U7624 (N_7624,N_6448,N_6168);
or U7625 (N_7625,N_6271,N_6700);
and U7626 (N_7626,N_6077,N_6444);
nand U7627 (N_7627,N_6026,N_6661);
xnor U7628 (N_7628,N_6271,N_6526);
and U7629 (N_7629,N_6912,N_6550);
xor U7630 (N_7630,N_6214,N_6588);
or U7631 (N_7631,N_6035,N_6531);
xnor U7632 (N_7632,N_6149,N_6042);
or U7633 (N_7633,N_6670,N_6486);
and U7634 (N_7634,N_6131,N_6938);
xor U7635 (N_7635,N_6421,N_6515);
xor U7636 (N_7636,N_6071,N_6630);
nor U7637 (N_7637,N_6340,N_6182);
and U7638 (N_7638,N_6784,N_6036);
xor U7639 (N_7639,N_6635,N_6138);
xnor U7640 (N_7640,N_6158,N_6599);
and U7641 (N_7641,N_6524,N_6020);
xnor U7642 (N_7642,N_6246,N_6113);
nand U7643 (N_7643,N_6252,N_6062);
nand U7644 (N_7644,N_6542,N_6308);
nand U7645 (N_7645,N_6164,N_6790);
xnor U7646 (N_7646,N_6699,N_6243);
or U7647 (N_7647,N_6527,N_6295);
nor U7648 (N_7648,N_6257,N_6520);
nand U7649 (N_7649,N_6091,N_6183);
or U7650 (N_7650,N_6218,N_6258);
nand U7651 (N_7651,N_6358,N_6994);
and U7652 (N_7652,N_6724,N_6295);
or U7653 (N_7653,N_6892,N_6089);
or U7654 (N_7654,N_6350,N_6049);
nand U7655 (N_7655,N_6303,N_6403);
nor U7656 (N_7656,N_6647,N_6483);
nand U7657 (N_7657,N_6528,N_6828);
or U7658 (N_7658,N_6798,N_6794);
or U7659 (N_7659,N_6100,N_6639);
and U7660 (N_7660,N_6273,N_6004);
and U7661 (N_7661,N_6089,N_6743);
and U7662 (N_7662,N_6335,N_6486);
xnor U7663 (N_7663,N_6271,N_6407);
and U7664 (N_7664,N_6828,N_6889);
nor U7665 (N_7665,N_6921,N_6329);
nor U7666 (N_7666,N_6356,N_6050);
nand U7667 (N_7667,N_6899,N_6966);
nand U7668 (N_7668,N_6901,N_6982);
and U7669 (N_7669,N_6955,N_6261);
and U7670 (N_7670,N_6273,N_6039);
or U7671 (N_7671,N_6644,N_6192);
and U7672 (N_7672,N_6394,N_6657);
nor U7673 (N_7673,N_6152,N_6615);
or U7674 (N_7674,N_6134,N_6345);
xnor U7675 (N_7675,N_6998,N_6585);
xnor U7676 (N_7676,N_6754,N_6400);
or U7677 (N_7677,N_6570,N_6026);
and U7678 (N_7678,N_6913,N_6025);
or U7679 (N_7679,N_6266,N_6839);
or U7680 (N_7680,N_6186,N_6238);
xnor U7681 (N_7681,N_6379,N_6462);
nor U7682 (N_7682,N_6168,N_6075);
nand U7683 (N_7683,N_6547,N_6666);
and U7684 (N_7684,N_6957,N_6949);
and U7685 (N_7685,N_6531,N_6072);
xor U7686 (N_7686,N_6202,N_6760);
xnor U7687 (N_7687,N_6073,N_6494);
or U7688 (N_7688,N_6068,N_6323);
nor U7689 (N_7689,N_6004,N_6889);
nor U7690 (N_7690,N_6578,N_6943);
and U7691 (N_7691,N_6990,N_6784);
nor U7692 (N_7692,N_6126,N_6950);
nor U7693 (N_7693,N_6781,N_6922);
xnor U7694 (N_7694,N_6314,N_6650);
nor U7695 (N_7695,N_6433,N_6856);
nor U7696 (N_7696,N_6621,N_6551);
and U7697 (N_7697,N_6773,N_6618);
nand U7698 (N_7698,N_6616,N_6938);
nor U7699 (N_7699,N_6627,N_6072);
xnor U7700 (N_7700,N_6288,N_6457);
or U7701 (N_7701,N_6187,N_6751);
or U7702 (N_7702,N_6305,N_6089);
nor U7703 (N_7703,N_6969,N_6826);
nand U7704 (N_7704,N_6073,N_6800);
and U7705 (N_7705,N_6005,N_6563);
or U7706 (N_7706,N_6315,N_6724);
xnor U7707 (N_7707,N_6858,N_6697);
xor U7708 (N_7708,N_6247,N_6907);
nor U7709 (N_7709,N_6264,N_6707);
and U7710 (N_7710,N_6358,N_6874);
nor U7711 (N_7711,N_6219,N_6142);
xor U7712 (N_7712,N_6951,N_6905);
or U7713 (N_7713,N_6394,N_6000);
and U7714 (N_7714,N_6979,N_6943);
or U7715 (N_7715,N_6505,N_6352);
nand U7716 (N_7716,N_6501,N_6614);
and U7717 (N_7717,N_6525,N_6535);
nand U7718 (N_7718,N_6408,N_6130);
or U7719 (N_7719,N_6532,N_6592);
and U7720 (N_7720,N_6101,N_6215);
and U7721 (N_7721,N_6660,N_6710);
nor U7722 (N_7722,N_6130,N_6531);
nand U7723 (N_7723,N_6724,N_6515);
or U7724 (N_7724,N_6757,N_6802);
or U7725 (N_7725,N_6609,N_6472);
or U7726 (N_7726,N_6118,N_6287);
and U7727 (N_7727,N_6872,N_6630);
nor U7728 (N_7728,N_6512,N_6739);
xor U7729 (N_7729,N_6251,N_6416);
xnor U7730 (N_7730,N_6344,N_6387);
nor U7731 (N_7731,N_6855,N_6514);
xor U7732 (N_7732,N_6286,N_6373);
nor U7733 (N_7733,N_6147,N_6979);
xnor U7734 (N_7734,N_6946,N_6709);
xnor U7735 (N_7735,N_6071,N_6349);
nand U7736 (N_7736,N_6914,N_6439);
xnor U7737 (N_7737,N_6881,N_6731);
and U7738 (N_7738,N_6841,N_6415);
xnor U7739 (N_7739,N_6482,N_6586);
nand U7740 (N_7740,N_6008,N_6559);
nor U7741 (N_7741,N_6847,N_6491);
nor U7742 (N_7742,N_6476,N_6226);
and U7743 (N_7743,N_6405,N_6061);
xnor U7744 (N_7744,N_6010,N_6909);
and U7745 (N_7745,N_6574,N_6610);
and U7746 (N_7746,N_6353,N_6768);
nor U7747 (N_7747,N_6617,N_6324);
nor U7748 (N_7748,N_6914,N_6555);
and U7749 (N_7749,N_6634,N_6152);
xnor U7750 (N_7750,N_6371,N_6019);
nor U7751 (N_7751,N_6327,N_6015);
or U7752 (N_7752,N_6276,N_6397);
nand U7753 (N_7753,N_6720,N_6202);
nand U7754 (N_7754,N_6975,N_6412);
nand U7755 (N_7755,N_6577,N_6937);
xnor U7756 (N_7756,N_6857,N_6991);
xnor U7757 (N_7757,N_6622,N_6819);
or U7758 (N_7758,N_6911,N_6754);
nor U7759 (N_7759,N_6294,N_6574);
nand U7760 (N_7760,N_6246,N_6090);
nor U7761 (N_7761,N_6198,N_6255);
or U7762 (N_7762,N_6776,N_6345);
nand U7763 (N_7763,N_6309,N_6559);
xnor U7764 (N_7764,N_6650,N_6748);
and U7765 (N_7765,N_6664,N_6870);
xor U7766 (N_7766,N_6049,N_6640);
xor U7767 (N_7767,N_6632,N_6873);
and U7768 (N_7768,N_6222,N_6799);
nand U7769 (N_7769,N_6217,N_6518);
nand U7770 (N_7770,N_6350,N_6707);
or U7771 (N_7771,N_6982,N_6184);
and U7772 (N_7772,N_6159,N_6738);
or U7773 (N_7773,N_6209,N_6111);
xnor U7774 (N_7774,N_6409,N_6597);
nor U7775 (N_7775,N_6653,N_6021);
xnor U7776 (N_7776,N_6597,N_6963);
nor U7777 (N_7777,N_6815,N_6166);
nand U7778 (N_7778,N_6006,N_6409);
xor U7779 (N_7779,N_6614,N_6685);
or U7780 (N_7780,N_6014,N_6087);
xnor U7781 (N_7781,N_6412,N_6646);
and U7782 (N_7782,N_6567,N_6142);
nor U7783 (N_7783,N_6809,N_6060);
xor U7784 (N_7784,N_6856,N_6930);
or U7785 (N_7785,N_6084,N_6380);
nand U7786 (N_7786,N_6916,N_6486);
or U7787 (N_7787,N_6234,N_6619);
xor U7788 (N_7788,N_6278,N_6335);
nor U7789 (N_7789,N_6999,N_6216);
and U7790 (N_7790,N_6535,N_6123);
and U7791 (N_7791,N_6996,N_6318);
and U7792 (N_7792,N_6764,N_6748);
xor U7793 (N_7793,N_6369,N_6692);
or U7794 (N_7794,N_6507,N_6188);
xor U7795 (N_7795,N_6580,N_6913);
nor U7796 (N_7796,N_6895,N_6063);
and U7797 (N_7797,N_6534,N_6059);
nor U7798 (N_7798,N_6758,N_6689);
and U7799 (N_7799,N_6809,N_6821);
and U7800 (N_7800,N_6096,N_6973);
xnor U7801 (N_7801,N_6043,N_6523);
or U7802 (N_7802,N_6763,N_6284);
or U7803 (N_7803,N_6771,N_6948);
or U7804 (N_7804,N_6731,N_6629);
and U7805 (N_7805,N_6802,N_6109);
and U7806 (N_7806,N_6066,N_6192);
xnor U7807 (N_7807,N_6979,N_6701);
nand U7808 (N_7808,N_6648,N_6996);
or U7809 (N_7809,N_6152,N_6274);
and U7810 (N_7810,N_6729,N_6737);
and U7811 (N_7811,N_6516,N_6560);
nand U7812 (N_7812,N_6474,N_6069);
or U7813 (N_7813,N_6467,N_6451);
and U7814 (N_7814,N_6501,N_6994);
nor U7815 (N_7815,N_6717,N_6530);
and U7816 (N_7816,N_6865,N_6600);
xor U7817 (N_7817,N_6509,N_6940);
and U7818 (N_7818,N_6737,N_6902);
nand U7819 (N_7819,N_6951,N_6128);
xor U7820 (N_7820,N_6103,N_6953);
or U7821 (N_7821,N_6640,N_6951);
xnor U7822 (N_7822,N_6089,N_6851);
nor U7823 (N_7823,N_6862,N_6551);
or U7824 (N_7824,N_6659,N_6433);
or U7825 (N_7825,N_6618,N_6731);
or U7826 (N_7826,N_6624,N_6514);
nor U7827 (N_7827,N_6400,N_6024);
and U7828 (N_7828,N_6502,N_6653);
nand U7829 (N_7829,N_6381,N_6698);
and U7830 (N_7830,N_6022,N_6755);
xor U7831 (N_7831,N_6860,N_6776);
or U7832 (N_7832,N_6920,N_6113);
nor U7833 (N_7833,N_6248,N_6685);
nor U7834 (N_7834,N_6684,N_6069);
nor U7835 (N_7835,N_6209,N_6518);
or U7836 (N_7836,N_6165,N_6556);
nor U7837 (N_7837,N_6400,N_6167);
nor U7838 (N_7838,N_6631,N_6061);
nor U7839 (N_7839,N_6200,N_6629);
or U7840 (N_7840,N_6303,N_6711);
and U7841 (N_7841,N_6759,N_6989);
or U7842 (N_7842,N_6999,N_6571);
xor U7843 (N_7843,N_6212,N_6827);
nor U7844 (N_7844,N_6973,N_6957);
or U7845 (N_7845,N_6746,N_6453);
xor U7846 (N_7846,N_6380,N_6447);
nor U7847 (N_7847,N_6603,N_6634);
nor U7848 (N_7848,N_6523,N_6300);
xnor U7849 (N_7849,N_6775,N_6328);
and U7850 (N_7850,N_6062,N_6533);
or U7851 (N_7851,N_6249,N_6278);
and U7852 (N_7852,N_6315,N_6031);
nor U7853 (N_7853,N_6888,N_6231);
nand U7854 (N_7854,N_6725,N_6181);
nand U7855 (N_7855,N_6023,N_6534);
or U7856 (N_7856,N_6346,N_6808);
xnor U7857 (N_7857,N_6081,N_6874);
and U7858 (N_7858,N_6072,N_6398);
or U7859 (N_7859,N_6631,N_6770);
xnor U7860 (N_7860,N_6898,N_6583);
and U7861 (N_7861,N_6228,N_6930);
nand U7862 (N_7862,N_6360,N_6036);
or U7863 (N_7863,N_6945,N_6094);
and U7864 (N_7864,N_6086,N_6632);
nor U7865 (N_7865,N_6415,N_6278);
or U7866 (N_7866,N_6725,N_6465);
nor U7867 (N_7867,N_6376,N_6791);
xor U7868 (N_7868,N_6076,N_6978);
nand U7869 (N_7869,N_6638,N_6337);
nor U7870 (N_7870,N_6003,N_6382);
and U7871 (N_7871,N_6297,N_6614);
nand U7872 (N_7872,N_6678,N_6785);
and U7873 (N_7873,N_6163,N_6313);
xnor U7874 (N_7874,N_6562,N_6850);
nand U7875 (N_7875,N_6833,N_6015);
and U7876 (N_7876,N_6208,N_6030);
nor U7877 (N_7877,N_6337,N_6127);
xor U7878 (N_7878,N_6926,N_6986);
and U7879 (N_7879,N_6026,N_6922);
or U7880 (N_7880,N_6398,N_6338);
or U7881 (N_7881,N_6123,N_6088);
or U7882 (N_7882,N_6691,N_6828);
or U7883 (N_7883,N_6379,N_6442);
nand U7884 (N_7884,N_6199,N_6069);
or U7885 (N_7885,N_6260,N_6966);
or U7886 (N_7886,N_6559,N_6702);
nor U7887 (N_7887,N_6465,N_6240);
nor U7888 (N_7888,N_6681,N_6702);
and U7889 (N_7889,N_6720,N_6988);
xor U7890 (N_7890,N_6602,N_6256);
nand U7891 (N_7891,N_6912,N_6473);
or U7892 (N_7892,N_6672,N_6915);
xnor U7893 (N_7893,N_6000,N_6946);
xnor U7894 (N_7894,N_6575,N_6583);
nor U7895 (N_7895,N_6368,N_6878);
and U7896 (N_7896,N_6928,N_6694);
xnor U7897 (N_7897,N_6650,N_6038);
and U7898 (N_7898,N_6213,N_6375);
nor U7899 (N_7899,N_6980,N_6056);
or U7900 (N_7900,N_6519,N_6563);
xnor U7901 (N_7901,N_6149,N_6091);
nand U7902 (N_7902,N_6571,N_6077);
nor U7903 (N_7903,N_6950,N_6652);
and U7904 (N_7904,N_6034,N_6611);
and U7905 (N_7905,N_6950,N_6128);
or U7906 (N_7906,N_6324,N_6325);
xnor U7907 (N_7907,N_6948,N_6038);
or U7908 (N_7908,N_6128,N_6003);
and U7909 (N_7909,N_6651,N_6208);
nand U7910 (N_7910,N_6414,N_6348);
or U7911 (N_7911,N_6187,N_6341);
or U7912 (N_7912,N_6851,N_6662);
xnor U7913 (N_7913,N_6507,N_6584);
or U7914 (N_7914,N_6435,N_6212);
xnor U7915 (N_7915,N_6242,N_6352);
and U7916 (N_7916,N_6367,N_6851);
or U7917 (N_7917,N_6188,N_6907);
or U7918 (N_7918,N_6792,N_6565);
nand U7919 (N_7919,N_6221,N_6907);
and U7920 (N_7920,N_6811,N_6729);
nor U7921 (N_7921,N_6942,N_6886);
nand U7922 (N_7922,N_6370,N_6484);
xnor U7923 (N_7923,N_6697,N_6756);
nand U7924 (N_7924,N_6391,N_6464);
and U7925 (N_7925,N_6378,N_6997);
and U7926 (N_7926,N_6025,N_6542);
and U7927 (N_7927,N_6024,N_6394);
nor U7928 (N_7928,N_6155,N_6205);
nand U7929 (N_7929,N_6592,N_6523);
and U7930 (N_7930,N_6593,N_6679);
nor U7931 (N_7931,N_6824,N_6133);
nor U7932 (N_7932,N_6140,N_6587);
or U7933 (N_7933,N_6654,N_6724);
nand U7934 (N_7934,N_6629,N_6374);
or U7935 (N_7935,N_6935,N_6209);
or U7936 (N_7936,N_6541,N_6699);
nand U7937 (N_7937,N_6488,N_6441);
xnor U7938 (N_7938,N_6435,N_6730);
or U7939 (N_7939,N_6591,N_6453);
and U7940 (N_7940,N_6397,N_6285);
and U7941 (N_7941,N_6374,N_6063);
xor U7942 (N_7942,N_6500,N_6657);
nor U7943 (N_7943,N_6726,N_6699);
nand U7944 (N_7944,N_6944,N_6045);
xor U7945 (N_7945,N_6891,N_6877);
xnor U7946 (N_7946,N_6667,N_6457);
nand U7947 (N_7947,N_6218,N_6802);
nand U7948 (N_7948,N_6652,N_6962);
or U7949 (N_7949,N_6343,N_6143);
nand U7950 (N_7950,N_6138,N_6376);
xor U7951 (N_7951,N_6291,N_6077);
nor U7952 (N_7952,N_6027,N_6701);
xnor U7953 (N_7953,N_6517,N_6650);
xor U7954 (N_7954,N_6466,N_6186);
nand U7955 (N_7955,N_6150,N_6311);
xor U7956 (N_7956,N_6874,N_6699);
and U7957 (N_7957,N_6113,N_6748);
or U7958 (N_7958,N_6913,N_6868);
nand U7959 (N_7959,N_6101,N_6684);
or U7960 (N_7960,N_6063,N_6085);
or U7961 (N_7961,N_6299,N_6998);
and U7962 (N_7962,N_6323,N_6128);
xnor U7963 (N_7963,N_6707,N_6060);
and U7964 (N_7964,N_6383,N_6565);
and U7965 (N_7965,N_6017,N_6047);
nor U7966 (N_7966,N_6898,N_6689);
and U7967 (N_7967,N_6186,N_6387);
nor U7968 (N_7968,N_6266,N_6938);
and U7969 (N_7969,N_6226,N_6644);
nor U7970 (N_7970,N_6795,N_6761);
nand U7971 (N_7971,N_6937,N_6078);
nand U7972 (N_7972,N_6698,N_6635);
xnor U7973 (N_7973,N_6776,N_6326);
nand U7974 (N_7974,N_6928,N_6358);
nor U7975 (N_7975,N_6910,N_6342);
xor U7976 (N_7976,N_6181,N_6593);
nor U7977 (N_7977,N_6464,N_6761);
nand U7978 (N_7978,N_6828,N_6927);
xnor U7979 (N_7979,N_6876,N_6482);
nand U7980 (N_7980,N_6306,N_6272);
xor U7981 (N_7981,N_6030,N_6784);
xor U7982 (N_7982,N_6968,N_6548);
and U7983 (N_7983,N_6294,N_6882);
nor U7984 (N_7984,N_6770,N_6739);
nand U7985 (N_7985,N_6974,N_6250);
xor U7986 (N_7986,N_6774,N_6990);
nor U7987 (N_7987,N_6261,N_6863);
nor U7988 (N_7988,N_6377,N_6448);
or U7989 (N_7989,N_6280,N_6417);
xnor U7990 (N_7990,N_6165,N_6835);
nand U7991 (N_7991,N_6180,N_6060);
nor U7992 (N_7992,N_6781,N_6703);
nand U7993 (N_7993,N_6344,N_6777);
nor U7994 (N_7994,N_6167,N_6724);
or U7995 (N_7995,N_6917,N_6272);
xor U7996 (N_7996,N_6127,N_6757);
or U7997 (N_7997,N_6596,N_6435);
and U7998 (N_7998,N_6053,N_6449);
nor U7999 (N_7999,N_6499,N_6611);
or U8000 (N_8000,N_7772,N_7137);
and U8001 (N_8001,N_7273,N_7672);
xor U8002 (N_8002,N_7382,N_7854);
nand U8003 (N_8003,N_7206,N_7057);
and U8004 (N_8004,N_7601,N_7512);
or U8005 (N_8005,N_7465,N_7887);
xor U8006 (N_8006,N_7931,N_7626);
nor U8007 (N_8007,N_7677,N_7515);
nand U8008 (N_8008,N_7207,N_7650);
or U8009 (N_8009,N_7370,N_7778);
xnor U8010 (N_8010,N_7424,N_7656);
and U8011 (N_8011,N_7686,N_7071);
nor U8012 (N_8012,N_7551,N_7398);
nor U8013 (N_8013,N_7932,N_7103);
nand U8014 (N_8014,N_7605,N_7482);
nand U8015 (N_8015,N_7969,N_7183);
or U8016 (N_8016,N_7599,N_7736);
xor U8017 (N_8017,N_7441,N_7507);
nor U8018 (N_8018,N_7224,N_7361);
nor U8019 (N_8019,N_7709,N_7245);
nand U8020 (N_8020,N_7602,N_7479);
xor U8021 (N_8021,N_7421,N_7776);
and U8022 (N_8022,N_7393,N_7270);
xor U8023 (N_8023,N_7338,N_7905);
or U8024 (N_8024,N_7452,N_7204);
nand U8025 (N_8025,N_7590,N_7352);
nand U8026 (N_8026,N_7826,N_7483);
or U8027 (N_8027,N_7464,N_7819);
and U8028 (N_8028,N_7453,N_7023);
nand U8029 (N_8029,N_7331,N_7033);
or U8030 (N_8030,N_7450,N_7915);
nor U8031 (N_8031,N_7566,N_7713);
and U8032 (N_8032,N_7746,N_7520);
nor U8033 (N_8033,N_7274,N_7378);
nand U8034 (N_8034,N_7291,N_7049);
and U8035 (N_8035,N_7865,N_7187);
nand U8036 (N_8036,N_7024,N_7981);
nor U8037 (N_8037,N_7165,N_7847);
nor U8038 (N_8038,N_7784,N_7570);
or U8039 (N_8039,N_7839,N_7807);
xnor U8040 (N_8040,N_7523,N_7619);
or U8041 (N_8041,N_7930,N_7917);
nor U8042 (N_8042,N_7946,N_7792);
and U8043 (N_8043,N_7173,N_7959);
or U8044 (N_8044,N_7690,N_7624);
nor U8045 (N_8045,N_7330,N_7783);
nand U8046 (N_8046,N_7800,N_7853);
nand U8047 (N_8047,N_7010,N_7284);
and U8048 (N_8048,N_7265,N_7864);
nor U8049 (N_8049,N_7387,N_7194);
and U8050 (N_8050,N_7868,N_7996);
nor U8051 (N_8051,N_7022,N_7164);
and U8052 (N_8052,N_7610,N_7445);
or U8053 (N_8053,N_7489,N_7580);
nor U8054 (N_8054,N_7423,N_7689);
or U8055 (N_8055,N_7789,N_7416);
or U8056 (N_8056,N_7428,N_7615);
nand U8057 (N_8057,N_7474,N_7434);
nor U8058 (N_8058,N_7034,N_7252);
nand U8059 (N_8059,N_7712,N_7621);
nor U8060 (N_8060,N_7112,N_7798);
nand U8061 (N_8061,N_7942,N_7253);
and U8062 (N_8062,N_7758,N_7732);
xnor U8063 (N_8063,N_7442,N_7038);
nor U8064 (N_8064,N_7018,N_7162);
xnor U8065 (N_8065,N_7659,N_7111);
or U8066 (N_8066,N_7501,N_7041);
or U8067 (N_8067,N_7129,N_7353);
xnor U8068 (N_8068,N_7589,N_7584);
nand U8069 (N_8069,N_7449,N_7524);
and U8070 (N_8070,N_7205,N_7062);
xnor U8071 (N_8071,N_7841,N_7168);
or U8072 (N_8072,N_7664,N_7364);
nand U8073 (N_8073,N_7567,N_7803);
xnor U8074 (N_8074,N_7851,N_7506);
nor U8075 (N_8075,N_7997,N_7029);
xor U8076 (N_8076,N_7240,N_7325);
and U8077 (N_8077,N_7134,N_7215);
nor U8078 (N_8078,N_7903,N_7059);
nand U8079 (N_8079,N_7249,N_7140);
nor U8080 (N_8080,N_7322,N_7283);
nand U8081 (N_8081,N_7052,N_7994);
nand U8082 (N_8082,N_7461,N_7375);
xnor U8083 (N_8083,N_7978,N_7993);
nand U8084 (N_8084,N_7899,N_7420);
or U8085 (N_8085,N_7949,N_7559);
or U8086 (N_8086,N_7318,N_7568);
nor U8087 (N_8087,N_7725,N_7092);
nand U8088 (N_8088,N_7830,N_7500);
xnor U8089 (N_8089,N_7646,N_7124);
and U8090 (N_8090,N_7358,N_7473);
or U8091 (N_8091,N_7926,N_7925);
and U8092 (N_8092,N_7212,N_7292);
xnor U8093 (N_8093,N_7480,N_7678);
and U8094 (N_8094,N_7333,N_7365);
xnor U8095 (N_8095,N_7403,N_7629);
or U8096 (N_8096,N_7790,N_7005);
nand U8097 (N_8097,N_7904,N_7153);
xnor U8098 (N_8098,N_7756,N_7475);
and U8099 (N_8099,N_7869,N_7402);
nor U8100 (N_8100,N_7995,N_7574);
nor U8101 (N_8101,N_7963,N_7635);
xnor U8102 (N_8102,N_7486,N_7829);
nand U8103 (N_8103,N_7235,N_7303);
or U8104 (N_8104,N_7127,N_7576);
nor U8105 (N_8105,N_7004,N_7104);
xor U8106 (N_8106,N_7857,N_7940);
and U8107 (N_8107,N_7669,N_7765);
nand U8108 (N_8108,N_7799,N_7553);
xnor U8109 (N_8109,N_7290,N_7060);
and U8110 (N_8110,N_7924,N_7189);
or U8111 (N_8111,N_7132,N_7457);
nor U8112 (N_8112,N_7115,N_7612);
nand U8113 (N_8113,N_7053,N_7150);
nor U8114 (N_8114,N_7907,N_7349);
xor U8115 (N_8115,N_7269,N_7101);
xnor U8116 (N_8116,N_7594,N_7710);
nand U8117 (N_8117,N_7469,N_7888);
and U8118 (N_8118,N_7722,N_7301);
nor U8119 (N_8119,N_7233,N_7462);
and U8120 (N_8120,N_7302,N_7455);
and U8121 (N_8121,N_7572,N_7562);
or U8122 (N_8122,N_7747,N_7064);
nand U8123 (N_8123,N_7945,N_7724);
or U8124 (N_8124,N_7431,N_7607);
nand U8125 (N_8125,N_7496,N_7446);
and U8126 (N_8126,N_7791,N_7716);
or U8127 (N_8127,N_7817,N_7222);
and U8128 (N_8128,N_7195,N_7844);
xnor U8129 (N_8129,N_7545,N_7967);
nand U8130 (N_8130,N_7935,N_7078);
nor U8131 (N_8131,N_7176,N_7311);
xor U8132 (N_8132,N_7682,N_7648);
and U8133 (N_8133,N_7999,N_7759);
nand U8134 (N_8134,N_7138,N_7761);
or U8135 (N_8135,N_7694,N_7381);
nor U8136 (N_8136,N_7914,N_7396);
nand U8137 (N_8137,N_7200,N_7987);
or U8138 (N_8138,N_7019,N_7780);
or U8139 (N_8139,N_7435,N_7961);
xor U8140 (N_8140,N_7699,N_7984);
and U8141 (N_8141,N_7404,N_7182);
nor U8142 (N_8142,N_7076,N_7988);
nor U8143 (N_8143,N_7871,N_7861);
nor U8144 (N_8144,N_7426,N_7372);
nor U8145 (N_8145,N_7406,N_7796);
nand U8146 (N_8146,N_7502,N_7117);
nor U8147 (N_8147,N_7571,N_7050);
or U8148 (N_8148,N_7055,N_7389);
or U8149 (N_8149,N_7866,N_7802);
nand U8150 (N_8150,N_7476,N_7118);
nor U8151 (N_8151,N_7676,N_7897);
or U8152 (N_8152,N_7108,N_7578);
xor U8153 (N_8153,N_7095,N_7685);
nor U8154 (N_8154,N_7696,N_7898);
xor U8155 (N_8155,N_7105,N_7636);
and U8156 (N_8156,N_7341,N_7237);
and U8157 (N_8157,N_7856,N_7691);
nor U8158 (N_8158,N_7146,N_7246);
xnor U8159 (N_8159,N_7219,N_7002);
nand U8160 (N_8160,N_7849,N_7394);
and U8161 (N_8161,N_7742,N_7367);
xor U8162 (N_8162,N_7573,N_7561);
xor U8163 (N_8163,N_7745,N_7279);
nand U8164 (N_8164,N_7822,N_7390);
and U8165 (N_8165,N_7068,N_7654);
nand U8166 (N_8166,N_7100,N_7250);
xnor U8167 (N_8167,N_7516,N_7016);
nor U8168 (N_8168,N_7409,N_7543);
nor U8169 (N_8169,N_7448,N_7779);
or U8170 (N_8170,N_7889,N_7070);
nand U8171 (N_8171,N_7876,N_7360);
nor U8172 (N_8172,N_7976,N_7848);
nor U8173 (N_8173,N_7007,N_7386);
and U8174 (N_8174,N_7335,N_7217);
xor U8175 (N_8175,N_7110,N_7313);
xnor U8176 (N_8176,N_7706,N_7180);
and U8177 (N_8177,N_7158,N_7762);
nor U8178 (N_8178,N_7884,N_7384);
nand U8179 (N_8179,N_7310,N_7090);
nand U8180 (N_8180,N_7198,N_7950);
or U8181 (N_8181,N_7102,N_7718);
or U8182 (N_8182,N_7651,N_7665);
nor U8183 (N_8183,N_7555,N_7009);
and U8184 (N_8184,N_7161,N_7348);
xnor U8185 (N_8185,N_7846,N_7466);
xor U8186 (N_8186,N_7517,N_7199);
nand U8187 (N_8187,N_7838,N_7125);
xor U8188 (N_8188,N_7873,N_7340);
and U8189 (N_8189,N_7518,N_7460);
and U8190 (N_8190,N_7521,N_7508);
and U8191 (N_8191,N_7788,N_7363);
xor U8192 (N_8192,N_7282,N_7632);
and U8193 (N_8193,N_7494,N_7616);
and U8194 (N_8194,N_7259,N_7047);
nor U8195 (N_8195,N_7356,N_7837);
nor U8196 (N_8196,N_7355,N_7777);
and U8197 (N_8197,N_7063,N_7326);
nand U8198 (N_8198,N_7089,N_7731);
nand U8199 (N_8199,N_7463,N_7391);
xnor U8200 (N_8200,N_7001,N_7281);
nand U8201 (N_8201,N_7201,N_7723);
nor U8202 (N_8202,N_7587,N_7708);
nand U8203 (N_8203,N_7763,N_7858);
nand U8204 (N_8204,N_7417,N_7261);
and U8205 (N_8205,N_7226,N_7294);
xnor U8206 (N_8206,N_7098,N_7174);
or U8207 (N_8207,N_7548,N_7514);
nor U8208 (N_8208,N_7843,N_7692);
xnor U8209 (N_8209,N_7618,N_7305);
and U8210 (N_8210,N_7850,N_7671);
xor U8211 (N_8211,N_7597,N_7879);
nand U8212 (N_8212,N_7135,N_7151);
and U8213 (N_8213,N_7885,N_7894);
and U8214 (N_8214,N_7828,N_7181);
nand U8215 (N_8215,N_7529,N_7919);
and U8216 (N_8216,N_7234,N_7878);
and U8217 (N_8217,N_7972,N_7027);
xnor U8218 (N_8218,N_7003,N_7046);
nor U8219 (N_8219,N_7640,N_7860);
or U8220 (N_8220,N_7097,N_7093);
and U8221 (N_8221,N_7037,N_7149);
xnor U8222 (N_8222,N_7160,N_7120);
nor U8223 (N_8223,N_7971,N_7412);
xnor U8224 (N_8224,N_7192,N_7008);
nand U8225 (N_8225,N_7304,N_7923);
nor U8226 (N_8226,N_7141,N_7220);
nor U8227 (N_8227,N_7955,N_7197);
xor U8228 (N_8228,N_7921,N_7603);
nor U8229 (N_8229,N_7721,N_7411);
and U8230 (N_8230,N_7155,N_7244);
or U8231 (N_8231,N_7373,N_7436);
xor U8232 (N_8232,N_7069,N_7755);
and U8233 (N_8233,N_7522,N_7541);
nand U8234 (N_8234,N_7067,N_7072);
or U8235 (N_8235,N_7422,N_7749);
and U8236 (N_8236,N_7503,N_7196);
nand U8237 (N_8237,N_7152,N_7272);
nor U8238 (N_8238,N_7751,N_7526);
and U8239 (N_8239,N_7805,N_7683);
xnor U8240 (N_8240,N_7558,N_7729);
nand U8241 (N_8241,N_7613,N_7020);
nand U8242 (N_8242,N_7432,N_7719);
or U8243 (N_8243,N_7179,N_7345);
nor U8244 (N_8244,N_7951,N_7734);
xor U8245 (N_8245,N_7286,N_7171);
and U8246 (N_8246,N_7744,N_7238);
or U8247 (N_8247,N_7513,N_7015);
nand U8248 (N_8248,N_7447,N_7701);
nor U8249 (N_8249,N_7357,N_7549);
or U8250 (N_8250,N_7628,N_7498);
or U8251 (N_8251,N_7680,N_7495);
or U8252 (N_8252,N_7661,N_7831);
nor U8253 (N_8253,N_7278,N_7738);
nor U8254 (N_8254,N_7663,N_7277);
and U8255 (N_8255,N_7908,N_7577);
nand U8256 (N_8256,N_7099,N_7223);
nand U8257 (N_8257,N_7214,N_7209);
nand U8258 (N_8258,N_7752,N_7730);
nor U8259 (N_8259,N_7938,N_7630);
xor U8260 (N_8260,N_7585,N_7407);
and U8261 (N_8261,N_7782,N_7642);
nand U8262 (N_8262,N_7280,N_7859);
nand U8263 (N_8263,N_7845,N_7643);
xor U8264 (N_8264,N_7821,N_7021);
nor U8265 (N_8265,N_7119,N_7232);
or U8266 (N_8266,N_7287,N_7637);
nor U8267 (N_8267,N_7490,N_7026);
or U8268 (N_8268,N_7241,N_7816);
nand U8269 (N_8269,N_7877,N_7986);
nor U8270 (N_8270,N_7852,N_7258);
nor U8271 (N_8271,N_7968,N_7257);
and U8272 (N_8272,N_7957,N_7874);
nor U8273 (N_8273,N_7880,N_7644);
nor U8274 (N_8274,N_7296,N_7264);
nand U8275 (N_8275,N_7983,N_7397);
nor U8276 (N_8276,N_7172,N_7666);
and U8277 (N_8277,N_7592,N_7148);
or U8278 (N_8278,N_7693,N_7528);
nor U8279 (N_8279,N_7084,N_7324);
nand U8280 (N_8280,N_7467,N_7727);
nand U8281 (N_8281,N_7346,N_7900);
or U8282 (N_8282,N_7660,N_7825);
xor U8283 (N_8283,N_7344,N_7263);
nor U8284 (N_8284,N_7649,N_7956);
xnor U8285 (N_8285,N_7992,N_7748);
nor U8286 (N_8286,N_7320,N_7557);
nor U8287 (N_8287,N_7886,N_7048);
nor U8288 (N_8288,N_7824,N_7948);
and U8289 (N_8289,N_7014,N_7647);
or U8290 (N_8290,N_7668,N_7918);
nand U8291 (N_8291,N_7532,N_7371);
nand U8292 (N_8292,N_7260,N_7025);
and U8293 (N_8293,N_7415,N_7684);
xnor U8294 (N_8294,N_7906,N_7964);
xor U8295 (N_8295,N_7741,N_7218);
nand U8296 (N_8296,N_7519,N_7347);
or U8297 (N_8297,N_7399,N_7083);
and U8298 (N_8298,N_7631,N_7753);
or U8299 (N_8299,N_7211,N_7444);
and U8300 (N_8300,N_7116,N_7653);
and U8301 (N_8301,N_7883,N_7109);
nor U8302 (N_8302,N_7377,N_7901);
nand U8303 (N_8303,N_7031,N_7236);
nor U8304 (N_8304,N_7096,N_7812);
xor U8305 (N_8305,N_7842,N_7035);
or U8306 (N_8306,N_7609,N_7509);
nand U8307 (N_8307,N_7113,N_7953);
nand U8308 (N_8308,N_7634,N_7814);
and U8309 (N_8309,N_7596,N_7032);
and U8310 (N_8310,N_7936,N_7221);
xor U8311 (N_8311,N_7892,N_7922);
or U8312 (N_8312,N_7891,N_7641);
nand U8313 (N_8313,N_7459,N_7400);
nand U8314 (N_8314,N_7662,N_7937);
or U8315 (N_8315,N_7652,N_7875);
nor U8316 (N_8316,N_7617,N_7472);
nand U8317 (N_8317,N_7768,N_7639);
nand U8318 (N_8318,N_7339,N_7623);
and U8319 (N_8319,N_7427,N_7510);
nand U8320 (N_8320,N_7638,N_7739);
xnor U8321 (N_8321,N_7960,N_7088);
nand U8322 (N_8322,N_7156,N_7947);
or U8323 (N_8323,N_7965,N_7657);
or U8324 (N_8324,N_7836,N_7916);
nor U8325 (N_8325,N_7369,N_7268);
xnor U8326 (N_8326,N_7985,N_7210);
nand U8327 (N_8327,N_7655,N_7362);
and U8328 (N_8328,N_7308,N_7579);
xnor U8329 (N_8329,N_7039,N_7456);
xor U8330 (N_8330,N_7000,N_7797);
xnor U8331 (N_8331,N_7419,N_7633);
xor U8332 (N_8332,N_7620,N_7306);
and U8333 (N_8333,N_7276,N_7136);
nor U8334 (N_8334,N_7085,N_7248);
nor U8335 (N_8335,N_7343,N_7328);
and U8336 (N_8336,N_7982,N_7504);
nand U8337 (N_8337,N_7833,N_7611);
nor U8338 (N_8338,N_7801,N_7401);
nand U8339 (N_8339,N_7006,N_7227);
xnor U8340 (N_8340,N_7608,N_7977);
nor U8341 (N_8341,N_7929,N_7547);
nand U8342 (N_8342,N_7531,N_7332);
and U8343 (N_8343,N_7715,N_7271);
nand U8344 (N_8344,N_7429,N_7795);
nand U8345 (N_8345,N_7533,N_7595);
xor U8346 (N_8346,N_7144,N_7870);
and U8347 (N_8347,N_7028,N_7970);
nor U8348 (N_8348,N_7809,N_7159);
nor U8349 (N_8349,N_7735,N_7228);
nor U8350 (N_8350,N_7359,N_7073);
or U8351 (N_8351,N_7262,N_7893);
nand U8352 (N_8352,N_7213,N_7430);
or U8353 (N_8353,N_7823,N_7082);
and U8354 (N_8354,N_7044,N_7334);
and U8355 (N_8355,N_7913,N_7530);
and U8356 (N_8356,N_7058,N_7771);
xor U8357 (N_8357,N_7535,N_7536);
nand U8358 (N_8358,N_7484,N_7872);
xnor U8359 (N_8359,N_7586,N_7203);
or U8360 (N_8360,N_7319,N_7061);
nor U8361 (N_8361,N_7505,N_7133);
nand U8362 (N_8362,N_7928,N_7040);
nor U8363 (N_8363,N_7990,N_7114);
or U8364 (N_8364,N_7697,N_7491);
and U8365 (N_8365,N_7775,N_7733);
or U8366 (N_8366,N_7711,N_7065);
or U8367 (N_8367,N_7374,N_7720);
nor U8368 (N_8368,N_7556,N_7525);
nand U8369 (N_8369,N_7499,N_7695);
nand U8370 (N_8370,N_7354,N_7740);
nor U8371 (N_8371,N_7862,N_7679);
and U8372 (N_8372,N_7760,N_7750);
and U8373 (N_8373,N_7493,N_7583);
nand U8374 (N_8374,N_7564,N_7974);
xor U8375 (N_8375,N_7167,N_7321);
nor U8376 (N_8376,N_7289,N_7770);
nor U8377 (N_8377,N_7835,N_7413);
xor U8378 (N_8378,N_7471,N_7042);
nor U8379 (N_8379,N_7470,N_7317);
or U8380 (N_8380,N_7086,N_7147);
or U8381 (N_8381,N_7497,N_7175);
nand U8382 (N_8382,N_7440,N_7477);
and U8383 (N_8383,N_7075,N_7944);
or U8384 (N_8384,N_7606,N_7939);
nand U8385 (N_8385,N_7658,N_7418);
nor U8386 (N_8386,N_7810,N_7645);
xor U8387 (N_8387,N_7670,N_7043);
nor U8388 (N_8388,N_7293,N_7454);
and U8389 (N_8389,N_7106,N_7840);
nand U8390 (N_8390,N_7737,N_7208);
nand U8391 (N_8391,N_7902,N_7910);
and U8392 (N_8392,N_7781,N_7309);
xnor U8393 (N_8393,N_7764,N_7056);
nor U8394 (N_8394,N_7488,N_7582);
and U8395 (N_8395,N_7934,N_7342);
xnor U8396 (N_8396,N_7973,N_7184);
or U8397 (N_8397,N_7154,N_7933);
and U8398 (N_8398,N_7080,N_7832);
xnor U8399 (N_8399,N_7980,N_7077);
xnor U8400 (N_8400,N_7593,N_7468);
xnor U8401 (N_8401,N_7376,N_7170);
or U8402 (N_8402,N_7912,N_7481);
xor U8403 (N_8403,N_7337,N_7704);
nand U8404 (N_8404,N_7705,N_7327);
nand U8405 (N_8405,N_7368,N_7811);
or U8406 (N_8406,N_7813,N_7591);
nand U8407 (N_8407,N_7011,N_7054);
or U8408 (N_8408,N_7251,N_7550);
nand U8409 (N_8409,N_7909,N_7408);
or U8410 (N_8410,N_7143,N_7216);
or U8411 (N_8411,N_7266,N_7794);
or U8412 (N_8412,N_7229,N_7688);
nand U8413 (N_8413,N_7145,N_7079);
xor U8414 (N_8414,N_7051,N_7177);
nand U8415 (N_8415,N_7863,N_7329);
xor U8416 (N_8416,N_7437,N_7989);
nand U8417 (N_8417,N_7242,N_7674);
nor U8418 (N_8418,N_7804,N_7726);
xor U8419 (N_8419,N_7350,N_7681);
nand U8420 (N_8420,N_7169,N_7379);
or U8421 (N_8421,N_7130,N_7163);
xor U8422 (N_8422,N_7754,N_7703);
or U8423 (N_8423,N_7012,N_7625);
xor U8424 (N_8424,N_7121,N_7546);
nand U8425 (N_8425,N_7538,N_7458);
nand U8426 (N_8426,N_7757,N_7438);
xor U8427 (N_8427,N_7698,N_7091);
nand U8428 (N_8428,N_7896,N_7614);
xor U8429 (N_8429,N_7895,N_7074);
or U8430 (N_8430,N_7107,N_7087);
or U8431 (N_8431,N_7433,N_7588);
or U8432 (N_8432,N_7239,N_7941);
nor U8433 (N_8433,N_7787,N_7539);
or U8434 (N_8434,N_7139,N_7920);
or U8435 (N_8435,N_7815,N_7998);
or U8436 (N_8436,N_7122,N_7806);
nor U8437 (N_8437,N_7300,N_7178);
nand U8438 (N_8438,N_7312,N_7492);
nand U8439 (N_8439,N_7793,N_7622);
xnor U8440 (N_8440,N_7185,N_7439);
and U8441 (N_8441,N_7707,N_7288);
or U8442 (N_8442,N_7927,N_7380);
nand U8443 (N_8443,N_7366,N_7414);
and U8444 (N_8444,N_7243,N_7425);
xor U8445 (N_8445,N_7254,N_7563);
nor U8446 (N_8446,N_7785,N_7094);
xor U8447 (N_8447,N_7979,N_7275);
xor U8448 (N_8448,N_7820,N_7231);
nand U8449 (N_8449,N_7581,N_7126);
nand U8450 (N_8450,N_7193,N_7767);
xnor U8451 (N_8451,N_7066,N_7769);
nor U8452 (N_8452,N_7827,N_7166);
nand U8453 (N_8453,N_7527,N_7534);
or U8454 (N_8454,N_7188,N_7540);
and U8455 (N_8455,N_7045,N_7190);
and U8456 (N_8456,N_7336,N_7255);
xor U8457 (N_8457,N_7728,N_7307);
nor U8458 (N_8458,N_7267,N_7766);
nand U8459 (N_8459,N_7351,N_7552);
xor U8460 (N_8460,N_7991,N_7673);
and U8461 (N_8461,N_7383,N_7627);
and U8462 (N_8462,N_7443,N_7943);
xnor U8463 (N_8463,N_7881,N_7714);
nor U8464 (N_8464,N_7247,N_7537);
nor U8465 (N_8465,N_7882,N_7225);
and U8466 (N_8466,N_7890,N_7478);
xnor U8467 (N_8467,N_7818,N_7451);
or U8468 (N_8468,N_7485,N_7128);
or U8469 (N_8469,N_7966,N_7230);
nor U8470 (N_8470,N_7131,N_7297);
nand U8471 (N_8471,N_7186,N_7554);
or U8472 (N_8472,N_7142,N_7773);
and U8473 (N_8473,N_7560,N_7385);
and U8474 (N_8474,N_7388,N_7954);
or U8475 (N_8475,N_7123,N_7030);
nor U8476 (N_8476,N_7808,N_7600);
xnor U8477 (N_8477,N_7743,N_7395);
or U8478 (N_8478,N_7544,N_7687);
or U8479 (N_8479,N_7157,N_7604);
nor U8480 (N_8480,N_7295,N_7392);
nand U8481 (N_8481,N_7867,N_7036);
nor U8482 (N_8482,N_7316,N_7202);
xnor U8483 (N_8483,N_7565,N_7834);
nand U8484 (N_8484,N_7081,N_7958);
nand U8485 (N_8485,N_7314,N_7542);
nor U8486 (N_8486,N_7511,N_7256);
and U8487 (N_8487,N_7285,N_7962);
xor U8488 (N_8488,N_7569,N_7405);
nand U8489 (N_8489,N_7911,N_7410);
and U8490 (N_8490,N_7667,N_7774);
and U8491 (N_8491,N_7952,N_7702);
nor U8492 (N_8492,N_7013,N_7975);
or U8493 (N_8493,N_7700,N_7598);
nor U8494 (N_8494,N_7786,N_7315);
nand U8495 (N_8495,N_7855,N_7575);
nand U8496 (N_8496,N_7191,N_7323);
or U8497 (N_8497,N_7017,N_7717);
xnor U8498 (N_8498,N_7298,N_7675);
nor U8499 (N_8499,N_7487,N_7299);
xnor U8500 (N_8500,N_7915,N_7340);
xnor U8501 (N_8501,N_7833,N_7381);
nand U8502 (N_8502,N_7162,N_7793);
and U8503 (N_8503,N_7151,N_7217);
and U8504 (N_8504,N_7643,N_7970);
xnor U8505 (N_8505,N_7297,N_7387);
nand U8506 (N_8506,N_7922,N_7912);
xnor U8507 (N_8507,N_7145,N_7373);
and U8508 (N_8508,N_7958,N_7720);
and U8509 (N_8509,N_7027,N_7909);
or U8510 (N_8510,N_7963,N_7456);
nor U8511 (N_8511,N_7243,N_7031);
or U8512 (N_8512,N_7139,N_7472);
xor U8513 (N_8513,N_7625,N_7923);
or U8514 (N_8514,N_7652,N_7337);
and U8515 (N_8515,N_7304,N_7682);
xnor U8516 (N_8516,N_7765,N_7350);
nor U8517 (N_8517,N_7332,N_7088);
xor U8518 (N_8518,N_7040,N_7785);
nor U8519 (N_8519,N_7767,N_7712);
or U8520 (N_8520,N_7406,N_7185);
nand U8521 (N_8521,N_7083,N_7298);
nor U8522 (N_8522,N_7747,N_7732);
nor U8523 (N_8523,N_7114,N_7173);
or U8524 (N_8524,N_7330,N_7807);
and U8525 (N_8525,N_7854,N_7681);
nor U8526 (N_8526,N_7903,N_7951);
and U8527 (N_8527,N_7218,N_7674);
xnor U8528 (N_8528,N_7352,N_7133);
nor U8529 (N_8529,N_7095,N_7062);
or U8530 (N_8530,N_7581,N_7878);
xnor U8531 (N_8531,N_7279,N_7338);
or U8532 (N_8532,N_7511,N_7519);
nand U8533 (N_8533,N_7924,N_7384);
or U8534 (N_8534,N_7619,N_7062);
nand U8535 (N_8535,N_7146,N_7268);
nor U8536 (N_8536,N_7182,N_7602);
xnor U8537 (N_8537,N_7626,N_7365);
and U8538 (N_8538,N_7026,N_7740);
nand U8539 (N_8539,N_7858,N_7453);
or U8540 (N_8540,N_7790,N_7984);
xor U8541 (N_8541,N_7916,N_7984);
nor U8542 (N_8542,N_7978,N_7999);
or U8543 (N_8543,N_7132,N_7879);
xor U8544 (N_8544,N_7523,N_7212);
or U8545 (N_8545,N_7902,N_7716);
nor U8546 (N_8546,N_7720,N_7647);
nand U8547 (N_8547,N_7839,N_7104);
xor U8548 (N_8548,N_7127,N_7708);
and U8549 (N_8549,N_7870,N_7893);
nand U8550 (N_8550,N_7449,N_7022);
nor U8551 (N_8551,N_7674,N_7089);
or U8552 (N_8552,N_7560,N_7821);
and U8553 (N_8553,N_7219,N_7966);
or U8554 (N_8554,N_7610,N_7717);
or U8555 (N_8555,N_7290,N_7778);
nand U8556 (N_8556,N_7878,N_7789);
xnor U8557 (N_8557,N_7290,N_7706);
nand U8558 (N_8558,N_7986,N_7520);
or U8559 (N_8559,N_7906,N_7040);
or U8560 (N_8560,N_7054,N_7659);
nor U8561 (N_8561,N_7666,N_7445);
nor U8562 (N_8562,N_7594,N_7055);
or U8563 (N_8563,N_7313,N_7868);
and U8564 (N_8564,N_7080,N_7652);
nand U8565 (N_8565,N_7584,N_7059);
xnor U8566 (N_8566,N_7756,N_7229);
xor U8567 (N_8567,N_7924,N_7574);
or U8568 (N_8568,N_7498,N_7757);
or U8569 (N_8569,N_7356,N_7196);
or U8570 (N_8570,N_7727,N_7959);
nand U8571 (N_8571,N_7778,N_7921);
and U8572 (N_8572,N_7026,N_7576);
nand U8573 (N_8573,N_7847,N_7719);
nor U8574 (N_8574,N_7177,N_7354);
and U8575 (N_8575,N_7582,N_7983);
and U8576 (N_8576,N_7711,N_7861);
and U8577 (N_8577,N_7849,N_7357);
and U8578 (N_8578,N_7524,N_7274);
or U8579 (N_8579,N_7823,N_7926);
nor U8580 (N_8580,N_7927,N_7740);
and U8581 (N_8581,N_7958,N_7203);
and U8582 (N_8582,N_7591,N_7638);
and U8583 (N_8583,N_7645,N_7082);
xnor U8584 (N_8584,N_7127,N_7417);
or U8585 (N_8585,N_7213,N_7565);
nand U8586 (N_8586,N_7870,N_7068);
and U8587 (N_8587,N_7994,N_7831);
or U8588 (N_8588,N_7284,N_7281);
or U8589 (N_8589,N_7214,N_7887);
xnor U8590 (N_8590,N_7973,N_7840);
xnor U8591 (N_8591,N_7551,N_7730);
nor U8592 (N_8592,N_7961,N_7654);
xor U8593 (N_8593,N_7070,N_7596);
nor U8594 (N_8594,N_7949,N_7478);
or U8595 (N_8595,N_7580,N_7053);
nor U8596 (N_8596,N_7080,N_7442);
nor U8597 (N_8597,N_7553,N_7427);
xnor U8598 (N_8598,N_7345,N_7667);
nor U8599 (N_8599,N_7739,N_7807);
nor U8600 (N_8600,N_7454,N_7027);
nor U8601 (N_8601,N_7266,N_7432);
and U8602 (N_8602,N_7923,N_7221);
nor U8603 (N_8603,N_7187,N_7059);
or U8604 (N_8604,N_7333,N_7151);
or U8605 (N_8605,N_7004,N_7550);
and U8606 (N_8606,N_7820,N_7393);
nor U8607 (N_8607,N_7461,N_7493);
nor U8608 (N_8608,N_7504,N_7860);
nor U8609 (N_8609,N_7461,N_7474);
nand U8610 (N_8610,N_7434,N_7730);
and U8611 (N_8611,N_7373,N_7322);
xnor U8612 (N_8612,N_7418,N_7808);
nand U8613 (N_8613,N_7233,N_7493);
or U8614 (N_8614,N_7801,N_7978);
nand U8615 (N_8615,N_7365,N_7160);
xor U8616 (N_8616,N_7085,N_7961);
xor U8617 (N_8617,N_7651,N_7628);
or U8618 (N_8618,N_7009,N_7151);
nor U8619 (N_8619,N_7143,N_7274);
xnor U8620 (N_8620,N_7615,N_7495);
nand U8621 (N_8621,N_7580,N_7207);
and U8622 (N_8622,N_7872,N_7144);
nand U8623 (N_8623,N_7048,N_7872);
or U8624 (N_8624,N_7917,N_7945);
nand U8625 (N_8625,N_7098,N_7093);
nand U8626 (N_8626,N_7951,N_7060);
nand U8627 (N_8627,N_7516,N_7332);
nand U8628 (N_8628,N_7807,N_7536);
nor U8629 (N_8629,N_7129,N_7748);
nor U8630 (N_8630,N_7759,N_7325);
or U8631 (N_8631,N_7506,N_7788);
or U8632 (N_8632,N_7192,N_7871);
or U8633 (N_8633,N_7802,N_7988);
or U8634 (N_8634,N_7090,N_7088);
nor U8635 (N_8635,N_7873,N_7658);
xnor U8636 (N_8636,N_7177,N_7414);
and U8637 (N_8637,N_7775,N_7176);
nand U8638 (N_8638,N_7168,N_7928);
xor U8639 (N_8639,N_7251,N_7898);
and U8640 (N_8640,N_7313,N_7471);
xor U8641 (N_8641,N_7242,N_7723);
or U8642 (N_8642,N_7262,N_7812);
nor U8643 (N_8643,N_7771,N_7487);
and U8644 (N_8644,N_7608,N_7957);
and U8645 (N_8645,N_7110,N_7559);
nand U8646 (N_8646,N_7228,N_7630);
nor U8647 (N_8647,N_7606,N_7911);
and U8648 (N_8648,N_7094,N_7560);
nand U8649 (N_8649,N_7322,N_7247);
xnor U8650 (N_8650,N_7749,N_7019);
nor U8651 (N_8651,N_7464,N_7286);
or U8652 (N_8652,N_7426,N_7310);
nand U8653 (N_8653,N_7173,N_7069);
xnor U8654 (N_8654,N_7177,N_7009);
nand U8655 (N_8655,N_7320,N_7504);
nand U8656 (N_8656,N_7514,N_7496);
xnor U8657 (N_8657,N_7308,N_7950);
nor U8658 (N_8658,N_7680,N_7724);
and U8659 (N_8659,N_7856,N_7813);
xor U8660 (N_8660,N_7656,N_7898);
nand U8661 (N_8661,N_7462,N_7090);
nand U8662 (N_8662,N_7192,N_7778);
xnor U8663 (N_8663,N_7814,N_7537);
and U8664 (N_8664,N_7674,N_7661);
and U8665 (N_8665,N_7940,N_7768);
xor U8666 (N_8666,N_7870,N_7282);
and U8667 (N_8667,N_7723,N_7848);
and U8668 (N_8668,N_7415,N_7141);
and U8669 (N_8669,N_7525,N_7567);
and U8670 (N_8670,N_7481,N_7348);
nand U8671 (N_8671,N_7192,N_7506);
and U8672 (N_8672,N_7726,N_7742);
nand U8673 (N_8673,N_7012,N_7020);
and U8674 (N_8674,N_7114,N_7762);
xnor U8675 (N_8675,N_7113,N_7848);
or U8676 (N_8676,N_7932,N_7637);
and U8677 (N_8677,N_7142,N_7284);
or U8678 (N_8678,N_7613,N_7716);
or U8679 (N_8679,N_7694,N_7217);
and U8680 (N_8680,N_7423,N_7406);
and U8681 (N_8681,N_7695,N_7831);
or U8682 (N_8682,N_7271,N_7566);
xor U8683 (N_8683,N_7047,N_7599);
nor U8684 (N_8684,N_7969,N_7297);
or U8685 (N_8685,N_7676,N_7390);
or U8686 (N_8686,N_7420,N_7482);
nand U8687 (N_8687,N_7369,N_7556);
or U8688 (N_8688,N_7203,N_7160);
nand U8689 (N_8689,N_7616,N_7522);
or U8690 (N_8690,N_7662,N_7257);
and U8691 (N_8691,N_7890,N_7555);
nor U8692 (N_8692,N_7730,N_7634);
nand U8693 (N_8693,N_7216,N_7933);
nor U8694 (N_8694,N_7715,N_7513);
and U8695 (N_8695,N_7385,N_7952);
xnor U8696 (N_8696,N_7717,N_7827);
or U8697 (N_8697,N_7651,N_7068);
xor U8698 (N_8698,N_7131,N_7055);
nand U8699 (N_8699,N_7775,N_7491);
and U8700 (N_8700,N_7482,N_7048);
and U8701 (N_8701,N_7250,N_7041);
and U8702 (N_8702,N_7051,N_7372);
nand U8703 (N_8703,N_7670,N_7062);
or U8704 (N_8704,N_7714,N_7595);
nand U8705 (N_8705,N_7690,N_7576);
or U8706 (N_8706,N_7515,N_7475);
xor U8707 (N_8707,N_7232,N_7032);
nor U8708 (N_8708,N_7620,N_7212);
xnor U8709 (N_8709,N_7773,N_7974);
or U8710 (N_8710,N_7885,N_7020);
xor U8711 (N_8711,N_7841,N_7221);
nor U8712 (N_8712,N_7267,N_7409);
xnor U8713 (N_8713,N_7052,N_7456);
xor U8714 (N_8714,N_7667,N_7724);
nor U8715 (N_8715,N_7531,N_7649);
or U8716 (N_8716,N_7448,N_7144);
and U8717 (N_8717,N_7992,N_7506);
or U8718 (N_8718,N_7274,N_7750);
xnor U8719 (N_8719,N_7960,N_7776);
nand U8720 (N_8720,N_7590,N_7599);
or U8721 (N_8721,N_7640,N_7002);
or U8722 (N_8722,N_7294,N_7302);
or U8723 (N_8723,N_7454,N_7066);
nor U8724 (N_8724,N_7175,N_7719);
and U8725 (N_8725,N_7511,N_7925);
and U8726 (N_8726,N_7436,N_7812);
xnor U8727 (N_8727,N_7754,N_7208);
nand U8728 (N_8728,N_7207,N_7232);
nand U8729 (N_8729,N_7961,N_7956);
and U8730 (N_8730,N_7627,N_7877);
or U8731 (N_8731,N_7856,N_7406);
nand U8732 (N_8732,N_7352,N_7060);
and U8733 (N_8733,N_7753,N_7374);
nand U8734 (N_8734,N_7660,N_7266);
and U8735 (N_8735,N_7710,N_7411);
or U8736 (N_8736,N_7076,N_7594);
nor U8737 (N_8737,N_7768,N_7424);
or U8738 (N_8738,N_7631,N_7181);
nand U8739 (N_8739,N_7663,N_7972);
or U8740 (N_8740,N_7586,N_7879);
xnor U8741 (N_8741,N_7270,N_7925);
xnor U8742 (N_8742,N_7178,N_7299);
nor U8743 (N_8743,N_7793,N_7450);
xor U8744 (N_8744,N_7837,N_7788);
nor U8745 (N_8745,N_7354,N_7256);
or U8746 (N_8746,N_7669,N_7333);
nand U8747 (N_8747,N_7945,N_7498);
nand U8748 (N_8748,N_7756,N_7450);
xnor U8749 (N_8749,N_7282,N_7917);
and U8750 (N_8750,N_7063,N_7248);
nand U8751 (N_8751,N_7835,N_7293);
or U8752 (N_8752,N_7905,N_7690);
nand U8753 (N_8753,N_7178,N_7250);
nand U8754 (N_8754,N_7278,N_7284);
xor U8755 (N_8755,N_7382,N_7541);
nor U8756 (N_8756,N_7219,N_7621);
or U8757 (N_8757,N_7030,N_7961);
xnor U8758 (N_8758,N_7370,N_7756);
or U8759 (N_8759,N_7906,N_7807);
and U8760 (N_8760,N_7753,N_7301);
or U8761 (N_8761,N_7198,N_7258);
xnor U8762 (N_8762,N_7710,N_7089);
nor U8763 (N_8763,N_7956,N_7177);
or U8764 (N_8764,N_7119,N_7152);
or U8765 (N_8765,N_7748,N_7223);
or U8766 (N_8766,N_7021,N_7928);
nand U8767 (N_8767,N_7279,N_7722);
xnor U8768 (N_8768,N_7778,N_7927);
nand U8769 (N_8769,N_7372,N_7299);
and U8770 (N_8770,N_7995,N_7733);
or U8771 (N_8771,N_7289,N_7590);
nand U8772 (N_8772,N_7059,N_7569);
nand U8773 (N_8773,N_7165,N_7976);
nand U8774 (N_8774,N_7939,N_7830);
nor U8775 (N_8775,N_7773,N_7934);
xnor U8776 (N_8776,N_7544,N_7617);
xor U8777 (N_8777,N_7280,N_7889);
xor U8778 (N_8778,N_7799,N_7673);
and U8779 (N_8779,N_7726,N_7007);
and U8780 (N_8780,N_7658,N_7426);
or U8781 (N_8781,N_7322,N_7756);
nand U8782 (N_8782,N_7946,N_7386);
and U8783 (N_8783,N_7364,N_7767);
or U8784 (N_8784,N_7144,N_7656);
and U8785 (N_8785,N_7237,N_7830);
xor U8786 (N_8786,N_7983,N_7355);
nand U8787 (N_8787,N_7613,N_7072);
xnor U8788 (N_8788,N_7824,N_7746);
xnor U8789 (N_8789,N_7052,N_7076);
and U8790 (N_8790,N_7801,N_7544);
and U8791 (N_8791,N_7618,N_7677);
and U8792 (N_8792,N_7095,N_7048);
xor U8793 (N_8793,N_7328,N_7909);
xor U8794 (N_8794,N_7387,N_7420);
or U8795 (N_8795,N_7163,N_7948);
nand U8796 (N_8796,N_7028,N_7125);
or U8797 (N_8797,N_7334,N_7285);
xor U8798 (N_8798,N_7337,N_7353);
nor U8799 (N_8799,N_7500,N_7955);
and U8800 (N_8800,N_7989,N_7169);
nor U8801 (N_8801,N_7663,N_7080);
xnor U8802 (N_8802,N_7511,N_7923);
xnor U8803 (N_8803,N_7587,N_7219);
nand U8804 (N_8804,N_7560,N_7344);
and U8805 (N_8805,N_7093,N_7364);
nor U8806 (N_8806,N_7660,N_7726);
nand U8807 (N_8807,N_7418,N_7097);
or U8808 (N_8808,N_7679,N_7155);
xnor U8809 (N_8809,N_7779,N_7288);
or U8810 (N_8810,N_7063,N_7486);
and U8811 (N_8811,N_7494,N_7283);
xor U8812 (N_8812,N_7318,N_7727);
or U8813 (N_8813,N_7476,N_7529);
nand U8814 (N_8814,N_7773,N_7972);
nand U8815 (N_8815,N_7926,N_7698);
xnor U8816 (N_8816,N_7927,N_7787);
or U8817 (N_8817,N_7185,N_7566);
nor U8818 (N_8818,N_7849,N_7666);
nand U8819 (N_8819,N_7467,N_7435);
nor U8820 (N_8820,N_7800,N_7351);
xnor U8821 (N_8821,N_7999,N_7112);
or U8822 (N_8822,N_7842,N_7033);
nand U8823 (N_8823,N_7139,N_7068);
and U8824 (N_8824,N_7089,N_7220);
nand U8825 (N_8825,N_7151,N_7681);
and U8826 (N_8826,N_7012,N_7441);
nand U8827 (N_8827,N_7208,N_7767);
and U8828 (N_8828,N_7257,N_7486);
and U8829 (N_8829,N_7809,N_7666);
nand U8830 (N_8830,N_7048,N_7360);
xor U8831 (N_8831,N_7560,N_7846);
xnor U8832 (N_8832,N_7058,N_7417);
nor U8833 (N_8833,N_7467,N_7562);
or U8834 (N_8834,N_7734,N_7725);
nand U8835 (N_8835,N_7688,N_7570);
or U8836 (N_8836,N_7543,N_7667);
xor U8837 (N_8837,N_7067,N_7342);
nand U8838 (N_8838,N_7733,N_7213);
nand U8839 (N_8839,N_7634,N_7933);
nor U8840 (N_8840,N_7762,N_7054);
or U8841 (N_8841,N_7571,N_7540);
or U8842 (N_8842,N_7535,N_7217);
xor U8843 (N_8843,N_7316,N_7733);
nand U8844 (N_8844,N_7846,N_7774);
nor U8845 (N_8845,N_7751,N_7548);
and U8846 (N_8846,N_7621,N_7940);
and U8847 (N_8847,N_7164,N_7631);
or U8848 (N_8848,N_7006,N_7312);
nor U8849 (N_8849,N_7976,N_7303);
nor U8850 (N_8850,N_7618,N_7460);
xor U8851 (N_8851,N_7123,N_7153);
or U8852 (N_8852,N_7119,N_7227);
nor U8853 (N_8853,N_7755,N_7062);
xor U8854 (N_8854,N_7571,N_7963);
xnor U8855 (N_8855,N_7313,N_7153);
and U8856 (N_8856,N_7053,N_7436);
or U8857 (N_8857,N_7370,N_7007);
nand U8858 (N_8858,N_7786,N_7987);
nand U8859 (N_8859,N_7385,N_7653);
xnor U8860 (N_8860,N_7013,N_7183);
or U8861 (N_8861,N_7628,N_7204);
nand U8862 (N_8862,N_7894,N_7555);
nand U8863 (N_8863,N_7706,N_7494);
or U8864 (N_8864,N_7885,N_7679);
nand U8865 (N_8865,N_7466,N_7917);
and U8866 (N_8866,N_7139,N_7440);
nand U8867 (N_8867,N_7926,N_7100);
and U8868 (N_8868,N_7566,N_7054);
nand U8869 (N_8869,N_7655,N_7100);
xor U8870 (N_8870,N_7723,N_7650);
nand U8871 (N_8871,N_7538,N_7758);
xor U8872 (N_8872,N_7475,N_7238);
nand U8873 (N_8873,N_7276,N_7508);
nand U8874 (N_8874,N_7840,N_7363);
or U8875 (N_8875,N_7227,N_7536);
nand U8876 (N_8876,N_7596,N_7288);
and U8877 (N_8877,N_7748,N_7556);
nor U8878 (N_8878,N_7699,N_7731);
nand U8879 (N_8879,N_7835,N_7977);
or U8880 (N_8880,N_7519,N_7571);
xnor U8881 (N_8881,N_7462,N_7896);
xnor U8882 (N_8882,N_7855,N_7082);
and U8883 (N_8883,N_7794,N_7377);
and U8884 (N_8884,N_7388,N_7427);
and U8885 (N_8885,N_7201,N_7079);
nor U8886 (N_8886,N_7344,N_7298);
xnor U8887 (N_8887,N_7568,N_7168);
nor U8888 (N_8888,N_7214,N_7393);
and U8889 (N_8889,N_7151,N_7436);
nand U8890 (N_8890,N_7938,N_7900);
or U8891 (N_8891,N_7193,N_7364);
nand U8892 (N_8892,N_7489,N_7332);
or U8893 (N_8893,N_7496,N_7958);
and U8894 (N_8894,N_7695,N_7188);
and U8895 (N_8895,N_7960,N_7303);
and U8896 (N_8896,N_7113,N_7746);
and U8897 (N_8897,N_7597,N_7183);
and U8898 (N_8898,N_7542,N_7538);
or U8899 (N_8899,N_7171,N_7653);
xor U8900 (N_8900,N_7346,N_7582);
or U8901 (N_8901,N_7618,N_7431);
nor U8902 (N_8902,N_7762,N_7540);
nand U8903 (N_8903,N_7265,N_7710);
and U8904 (N_8904,N_7444,N_7108);
nand U8905 (N_8905,N_7844,N_7699);
or U8906 (N_8906,N_7389,N_7388);
nor U8907 (N_8907,N_7375,N_7448);
or U8908 (N_8908,N_7388,N_7707);
and U8909 (N_8909,N_7844,N_7219);
nand U8910 (N_8910,N_7160,N_7780);
or U8911 (N_8911,N_7767,N_7839);
nor U8912 (N_8912,N_7014,N_7816);
nand U8913 (N_8913,N_7615,N_7475);
or U8914 (N_8914,N_7240,N_7749);
nor U8915 (N_8915,N_7981,N_7197);
and U8916 (N_8916,N_7451,N_7166);
and U8917 (N_8917,N_7693,N_7479);
nand U8918 (N_8918,N_7179,N_7278);
xnor U8919 (N_8919,N_7797,N_7298);
and U8920 (N_8920,N_7584,N_7722);
nor U8921 (N_8921,N_7979,N_7842);
nand U8922 (N_8922,N_7334,N_7172);
or U8923 (N_8923,N_7865,N_7653);
xor U8924 (N_8924,N_7011,N_7432);
xor U8925 (N_8925,N_7022,N_7165);
nand U8926 (N_8926,N_7420,N_7087);
or U8927 (N_8927,N_7834,N_7025);
xnor U8928 (N_8928,N_7914,N_7981);
nor U8929 (N_8929,N_7184,N_7315);
nor U8930 (N_8930,N_7072,N_7042);
nor U8931 (N_8931,N_7204,N_7772);
xnor U8932 (N_8932,N_7034,N_7653);
nand U8933 (N_8933,N_7374,N_7451);
xor U8934 (N_8934,N_7044,N_7894);
nand U8935 (N_8935,N_7495,N_7195);
nor U8936 (N_8936,N_7059,N_7750);
nor U8937 (N_8937,N_7620,N_7143);
and U8938 (N_8938,N_7124,N_7836);
nand U8939 (N_8939,N_7175,N_7492);
nand U8940 (N_8940,N_7653,N_7792);
nor U8941 (N_8941,N_7150,N_7286);
xnor U8942 (N_8942,N_7950,N_7732);
or U8943 (N_8943,N_7566,N_7897);
and U8944 (N_8944,N_7636,N_7408);
or U8945 (N_8945,N_7382,N_7354);
or U8946 (N_8946,N_7880,N_7184);
xnor U8947 (N_8947,N_7272,N_7392);
xnor U8948 (N_8948,N_7247,N_7870);
nand U8949 (N_8949,N_7854,N_7067);
nor U8950 (N_8950,N_7463,N_7136);
and U8951 (N_8951,N_7932,N_7481);
and U8952 (N_8952,N_7766,N_7329);
nor U8953 (N_8953,N_7247,N_7963);
xnor U8954 (N_8954,N_7964,N_7117);
and U8955 (N_8955,N_7974,N_7414);
nand U8956 (N_8956,N_7547,N_7648);
nor U8957 (N_8957,N_7533,N_7612);
xor U8958 (N_8958,N_7051,N_7655);
nor U8959 (N_8959,N_7701,N_7747);
nand U8960 (N_8960,N_7772,N_7380);
or U8961 (N_8961,N_7716,N_7922);
nor U8962 (N_8962,N_7552,N_7609);
nor U8963 (N_8963,N_7076,N_7001);
or U8964 (N_8964,N_7447,N_7135);
nand U8965 (N_8965,N_7503,N_7895);
xor U8966 (N_8966,N_7526,N_7094);
nand U8967 (N_8967,N_7200,N_7395);
and U8968 (N_8968,N_7333,N_7043);
xor U8969 (N_8969,N_7733,N_7078);
xnor U8970 (N_8970,N_7897,N_7556);
xor U8971 (N_8971,N_7697,N_7892);
or U8972 (N_8972,N_7754,N_7089);
or U8973 (N_8973,N_7832,N_7468);
nand U8974 (N_8974,N_7968,N_7947);
xor U8975 (N_8975,N_7603,N_7062);
nand U8976 (N_8976,N_7366,N_7531);
xor U8977 (N_8977,N_7723,N_7814);
xnor U8978 (N_8978,N_7725,N_7672);
nand U8979 (N_8979,N_7513,N_7157);
nand U8980 (N_8980,N_7469,N_7645);
and U8981 (N_8981,N_7293,N_7561);
xnor U8982 (N_8982,N_7005,N_7696);
nor U8983 (N_8983,N_7692,N_7137);
nand U8984 (N_8984,N_7103,N_7556);
or U8985 (N_8985,N_7339,N_7827);
nand U8986 (N_8986,N_7023,N_7474);
nand U8987 (N_8987,N_7035,N_7200);
nand U8988 (N_8988,N_7896,N_7936);
or U8989 (N_8989,N_7037,N_7873);
nor U8990 (N_8990,N_7374,N_7491);
xor U8991 (N_8991,N_7564,N_7309);
or U8992 (N_8992,N_7441,N_7121);
and U8993 (N_8993,N_7418,N_7520);
and U8994 (N_8994,N_7394,N_7936);
or U8995 (N_8995,N_7336,N_7649);
nand U8996 (N_8996,N_7849,N_7663);
and U8997 (N_8997,N_7002,N_7609);
nand U8998 (N_8998,N_7842,N_7050);
nand U8999 (N_8999,N_7065,N_7892);
and U9000 (N_9000,N_8502,N_8142);
nor U9001 (N_9001,N_8500,N_8710);
nand U9002 (N_9002,N_8685,N_8618);
and U9003 (N_9003,N_8783,N_8503);
or U9004 (N_9004,N_8115,N_8845);
nand U9005 (N_9005,N_8980,N_8914);
nand U9006 (N_9006,N_8918,N_8517);
xor U9007 (N_9007,N_8775,N_8300);
and U9008 (N_9008,N_8823,N_8647);
nand U9009 (N_9009,N_8921,N_8522);
and U9010 (N_9010,N_8005,N_8784);
nand U9011 (N_9011,N_8679,N_8063);
nor U9012 (N_9012,N_8424,N_8272);
xor U9013 (N_9013,N_8144,N_8334);
and U9014 (N_9014,N_8123,N_8733);
and U9015 (N_9015,N_8003,N_8730);
nor U9016 (N_9016,N_8567,N_8542);
nand U9017 (N_9017,N_8943,N_8904);
and U9018 (N_9018,N_8229,N_8853);
nor U9019 (N_9019,N_8555,N_8960);
and U9020 (N_9020,N_8094,N_8535);
nor U9021 (N_9021,N_8954,N_8852);
nor U9022 (N_9022,N_8291,N_8377);
xor U9023 (N_9023,N_8372,N_8885);
or U9024 (N_9024,N_8975,N_8600);
nor U9025 (N_9025,N_8330,N_8350);
and U9026 (N_9026,N_8514,N_8586);
nand U9027 (N_9027,N_8982,N_8268);
nand U9028 (N_9028,N_8041,N_8989);
and U9029 (N_9029,N_8327,N_8070);
and U9030 (N_9030,N_8037,N_8961);
nand U9031 (N_9031,N_8749,N_8688);
nand U9032 (N_9032,N_8270,N_8298);
and U9033 (N_9033,N_8831,N_8024);
and U9034 (N_9034,N_8745,N_8842);
xor U9035 (N_9035,N_8707,N_8058);
or U9036 (N_9036,N_8414,N_8684);
and U9037 (N_9037,N_8103,N_8338);
or U9038 (N_9038,N_8344,N_8172);
xor U9039 (N_9039,N_8076,N_8322);
and U9040 (N_9040,N_8520,N_8341);
nor U9041 (N_9041,N_8256,N_8169);
nor U9042 (N_9042,N_8219,N_8443);
and U9043 (N_9043,N_8218,N_8597);
and U9044 (N_9044,N_8881,N_8049);
nor U9045 (N_9045,N_8576,N_8035);
nor U9046 (N_9046,N_8366,N_8480);
xor U9047 (N_9047,N_8355,N_8027);
xnor U9048 (N_9048,N_8947,N_8721);
nor U9049 (N_9049,N_8483,N_8561);
nand U9050 (N_9050,N_8451,N_8620);
and U9051 (N_9051,N_8922,N_8209);
or U9052 (N_9052,N_8747,N_8609);
xor U9053 (N_9053,N_8902,N_8036);
or U9054 (N_9054,N_8441,N_8112);
xnor U9055 (N_9055,N_8716,N_8352);
and U9056 (N_9056,N_8602,N_8171);
xnor U9057 (N_9057,N_8762,N_8486);
nand U9058 (N_9058,N_8471,N_8430);
and U9059 (N_9059,N_8438,N_8621);
nor U9060 (N_9060,N_8120,N_8109);
and U9061 (N_9061,N_8636,N_8856);
xor U9062 (N_9062,N_8162,N_8860);
and U9063 (N_9063,N_8955,N_8497);
and U9064 (N_9064,N_8368,N_8985);
or U9065 (N_9065,N_8155,N_8981);
or U9066 (N_9066,N_8164,N_8454);
nor U9067 (N_9067,N_8997,N_8869);
nor U9068 (N_9068,N_8400,N_8077);
nand U9069 (N_9069,N_8066,N_8953);
or U9070 (N_9070,N_8217,N_8059);
or U9071 (N_9071,N_8401,N_8106);
or U9072 (N_9072,N_8202,N_8292);
xnor U9073 (N_9073,N_8548,N_8131);
and U9074 (N_9074,N_8667,N_8890);
nor U9075 (N_9075,N_8245,N_8701);
xor U9076 (N_9076,N_8868,N_8148);
and U9077 (N_9077,N_8487,N_8072);
and U9078 (N_9078,N_8055,N_8593);
nand U9079 (N_9079,N_8014,N_8818);
nand U9080 (N_9080,N_8858,N_8630);
and U9081 (N_9081,N_8578,N_8524);
xnor U9082 (N_9082,N_8010,N_8391);
or U9083 (N_9083,N_8864,N_8269);
nand U9084 (N_9084,N_8507,N_8098);
or U9085 (N_9085,N_8089,N_8894);
nor U9086 (N_9086,N_8175,N_8791);
and U9087 (N_9087,N_8968,N_8797);
nor U9088 (N_9088,N_8848,N_8316);
nand U9089 (N_9089,N_8302,N_8867);
and U9090 (N_9090,N_8819,N_8840);
and U9091 (N_9091,N_8495,N_8937);
and U9092 (N_9092,N_8773,N_8444);
xor U9093 (N_9093,N_8697,N_8187);
nand U9094 (N_9094,N_8192,N_8671);
xnor U9095 (N_9095,N_8595,N_8396);
or U9096 (N_9096,N_8389,N_8884);
xnor U9097 (N_9097,N_8594,N_8157);
nand U9098 (N_9098,N_8457,N_8122);
and U9099 (N_9099,N_8891,N_8538);
nor U9100 (N_9100,N_8184,N_8442);
and U9101 (N_9101,N_8932,N_8725);
or U9102 (N_9102,N_8200,N_8404);
and U9103 (N_9103,N_8962,N_8562);
or U9104 (N_9104,N_8080,N_8518);
xnor U9105 (N_9105,N_8043,N_8477);
xnor U9106 (N_9106,N_8988,N_8761);
nand U9107 (N_9107,N_8001,N_8614);
nor U9108 (N_9108,N_8494,N_8794);
nand U9109 (N_9109,N_8363,N_8608);
nor U9110 (N_9110,N_8052,N_8336);
nand U9111 (N_9111,N_8167,N_8537);
xnor U9112 (N_9112,N_8478,N_8303);
nor U9113 (N_9113,N_8248,N_8166);
nand U9114 (N_9114,N_8912,N_8908);
nor U9115 (N_9115,N_8545,N_8754);
or U9116 (N_9116,N_8455,N_8698);
nand U9117 (N_9117,N_8023,N_8850);
or U9118 (N_9118,N_8820,N_8504);
and U9119 (N_9119,N_8149,N_8326);
or U9120 (N_9120,N_8727,N_8657);
nor U9121 (N_9121,N_8787,N_8228);
nor U9122 (N_9122,N_8785,N_8592);
xor U9123 (N_9123,N_8097,N_8910);
and U9124 (N_9124,N_8750,N_8459);
and U9125 (N_9125,N_8689,N_8277);
xor U9126 (N_9126,N_8481,N_8473);
nor U9127 (N_9127,N_8623,N_8990);
and U9128 (N_9128,N_8876,N_8861);
nor U9129 (N_9129,N_8060,N_8544);
xnor U9130 (N_9130,N_8051,N_8660);
and U9131 (N_9131,N_8723,N_8738);
nor U9132 (N_9132,N_8111,N_8411);
or U9133 (N_9133,N_8057,N_8339);
or U9134 (N_9134,N_8516,N_8911);
or U9135 (N_9135,N_8901,N_8752);
or U9136 (N_9136,N_8371,N_8583);
xnor U9137 (N_9137,N_8464,N_8511);
xor U9138 (N_9138,N_8095,N_8267);
nor U9139 (N_9139,N_8129,N_8484);
and U9140 (N_9140,N_8233,N_8474);
nor U9141 (N_9141,N_8694,N_8488);
nor U9142 (N_9142,N_8616,N_8116);
nor U9143 (N_9143,N_8604,N_8615);
nor U9144 (N_9144,N_8826,N_8413);
or U9145 (N_9145,N_8976,N_8665);
and U9146 (N_9146,N_8903,N_8333);
nor U9147 (N_9147,N_8417,N_8812);
nand U9148 (N_9148,N_8439,N_8559);
or U9149 (N_9149,N_8917,N_8046);
nor U9150 (N_9150,N_8288,N_8729);
nor U9151 (N_9151,N_8654,N_8798);
nand U9152 (N_9152,N_8436,N_8458);
xnor U9153 (N_9153,N_8191,N_8728);
xor U9154 (N_9154,N_8993,N_8580);
xnor U9155 (N_9155,N_8427,N_8532);
xor U9156 (N_9156,N_8216,N_8713);
nand U9157 (N_9157,N_8346,N_8809);
nor U9158 (N_9158,N_8755,N_8412);
nor U9159 (N_9159,N_8469,N_8977);
nor U9160 (N_9160,N_8470,N_8779);
nor U9161 (N_9161,N_8979,N_8627);
nand U9162 (N_9162,N_8475,N_8744);
nor U9163 (N_9163,N_8748,N_8824);
and U9164 (N_9164,N_8632,N_8138);
nand U9165 (N_9165,N_8663,N_8032);
xor U9166 (N_9166,N_8179,N_8570);
nor U9167 (N_9167,N_8306,N_8662);
or U9168 (N_9168,N_8073,N_8093);
nor U9169 (N_9169,N_8311,N_8974);
nor U9170 (N_9170,N_8033,N_8053);
nand U9171 (N_9171,N_8530,N_8380);
xnor U9172 (N_9172,N_8558,N_8044);
xor U9173 (N_9173,N_8998,N_8930);
and U9174 (N_9174,N_8619,N_8612);
nand U9175 (N_9175,N_8923,N_8531);
or U9176 (N_9176,N_8203,N_8603);
or U9177 (N_9177,N_8577,N_8739);
xnor U9178 (N_9178,N_8509,N_8950);
nand U9179 (N_9179,N_8714,N_8581);
or U9180 (N_9180,N_8587,N_8638);
or U9181 (N_9181,N_8347,N_8141);
nand U9182 (N_9182,N_8362,N_8007);
or U9183 (N_9183,N_8758,N_8238);
and U9184 (N_9184,N_8395,N_8100);
and U9185 (N_9185,N_8512,N_8045);
nand U9186 (N_9186,N_8243,N_8241);
xor U9187 (N_9187,N_8666,N_8952);
nor U9188 (N_9188,N_8276,N_8656);
and U9189 (N_9189,N_8074,N_8168);
nand U9190 (N_9190,N_8190,N_8337);
and U9191 (N_9191,N_8026,N_8235);
or U9192 (N_9192,N_8147,N_8956);
nor U9193 (N_9193,N_8879,N_8403);
and U9194 (N_9194,N_8220,N_8145);
and U9195 (N_9195,N_8692,N_8492);
or U9196 (N_9196,N_8317,N_8221);
xnor U9197 (N_9197,N_8645,N_8434);
nor U9198 (N_9198,N_8971,N_8022);
and U9199 (N_9199,N_8970,N_8485);
xnor U9200 (N_9200,N_8348,N_8181);
xnor U9201 (N_9201,N_8318,N_8153);
xnor U9202 (N_9202,N_8081,N_8892);
nor U9203 (N_9203,N_8260,N_8004);
nor U9204 (N_9204,N_8320,N_8789);
nand U9205 (N_9205,N_8539,N_8087);
or U9206 (N_9206,N_8199,N_8703);
nand U9207 (N_9207,N_8139,N_8626);
or U9208 (N_9208,N_8564,N_8527);
nand U9209 (N_9209,N_8415,N_8385);
xor U9210 (N_9210,N_8641,N_8084);
nand U9211 (N_9211,N_8437,N_8513);
nor U9212 (N_9212,N_8176,N_8965);
nand U9213 (N_9213,N_8499,N_8813);
nand U9214 (N_9214,N_8222,N_8855);
nor U9215 (N_9215,N_8900,N_8646);
or U9216 (N_9216,N_8801,N_8865);
nor U9217 (N_9217,N_8331,N_8482);
or U9218 (N_9218,N_8031,N_8622);
nand U9219 (N_9219,N_8648,N_8040);
or U9220 (N_9220,N_8143,N_8661);
and U9221 (N_9221,N_8939,N_8599);
and U9222 (N_9222,N_8397,N_8874);
and U9223 (N_9223,N_8390,N_8572);
xnor U9224 (N_9224,N_8030,N_8983);
and U9225 (N_9225,N_8768,N_8405);
nand U9226 (N_9226,N_8329,N_8054);
or U9227 (N_9227,N_8285,N_8793);
xnor U9228 (N_9228,N_8828,N_8704);
or U9229 (N_9229,N_8510,N_8025);
or U9230 (N_9230,N_8948,N_8899);
or U9231 (N_9231,N_8357,N_8283);
or U9232 (N_9232,N_8695,N_8432);
and U9233 (N_9233,N_8696,N_8601);
and U9234 (N_9234,N_8996,N_8655);
and U9235 (N_9235,N_8829,N_8584);
nor U9236 (N_9236,N_8286,N_8772);
and U9237 (N_9237,N_8259,N_8686);
and U9238 (N_9238,N_8673,N_8136);
nor U9239 (N_9239,N_8712,N_8195);
nor U9240 (N_9240,N_8223,N_8582);
xor U9241 (N_9241,N_8928,N_8064);
xor U9242 (N_9242,N_8546,N_8197);
xnor U9243 (N_9243,N_8585,N_8050);
or U9244 (N_9244,N_8849,N_8994);
xor U9245 (N_9245,N_8523,N_8871);
xnor U9246 (N_9246,N_8308,N_8140);
xnor U9247 (N_9247,N_8447,N_8491);
xnor U9248 (N_9248,N_8261,N_8958);
nand U9249 (N_9249,N_8731,N_8722);
or U9250 (N_9250,N_8463,N_8128);
nand U9251 (N_9251,N_8501,N_8183);
and U9252 (N_9252,N_8916,N_8895);
nor U9253 (N_9253,N_8158,N_8254);
nand U9254 (N_9254,N_8406,N_8806);
and U9255 (N_9255,N_8194,N_8508);
nor U9256 (N_9256,N_8549,N_8999);
xor U9257 (N_9257,N_8575,N_8383);
or U9258 (N_9258,N_8253,N_8332);
or U9259 (N_9259,N_8717,N_8560);
or U9260 (N_9260,N_8225,N_8935);
xnor U9261 (N_9261,N_8893,N_8882);
xnor U9262 (N_9262,N_8307,N_8110);
nor U9263 (N_9263,N_8515,N_8675);
nand U9264 (N_9264,N_8816,N_8554);
nand U9265 (N_9265,N_8863,N_8418);
and U9266 (N_9266,N_8013,N_8808);
nand U9267 (N_9267,N_8872,N_8929);
xnor U9268 (N_9268,N_8264,N_8295);
and U9269 (N_9269,N_8117,N_8720);
and U9270 (N_9270,N_8551,N_8769);
and U9271 (N_9271,N_8681,N_8841);
xor U9272 (N_9272,N_8668,N_8015);
or U9273 (N_9273,N_8170,N_8843);
and U9274 (N_9274,N_8847,N_8294);
or U9275 (N_9275,N_8541,N_8342);
xor U9276 (N_9276,N_8068,N_8062);
nand U9277 (N_9277,N_8314,N_8114);
and U9278 (N_9278,N_8653,N_8009);
nor U9279 (N_9279,N_8433,N_8156);
or U9280 (N_9280,N_8016,N_8319);
nand U9281 (N_9281,N_8237,N_8297);
nor U9282 (N_9282,N_8821,N_8741);
nor U9283 (N_9283,N_8658,N_8506);
and U9284 (N_9284,N_8101,N_8519);
nor U9285 (N_9285,N_8328,N_8568);
nand U9286 (N_9286,N_8090,N_8118);
nor U9287 (N_9287,N_8827,N_8940);
and U9288 (N_9288,N_8177,N_8732);
and U9289 (N_9289,N_8425,N_8931);
nor U9290 (N_9290,N_8198,N_8765);
xnor U9291 (N_9291,N_8649,N_8764);
nor U9292 (N_9292,N_8651,N_8724);
and U9293 (N_9293,N_8693,N_8378);
or U9294 (N_9294,N_8907,N_8699);
or U9295 (N_9295,N_8065,N_8282);
nor U9296 (N_9296,N_8132,N_8774);
nor U9297 (N_9297,N_8251,N_8607);
nand U9298 (N_9298,N_8373,N_8146);
nor U9299 (N_9299,N_8605,N_8674);
nor U9300 (N_9300,N_8002,N_8244);
nor U9301 (N_9301,N_8263,N_8866);
xor U9302 (N_9302,N_8836,N_8777);
nand U9303 (N_9303,N_8669,N_8886);
and U9304 (N_9304,N_8275,N_8945);
and U9305 (N_9305,N_8811,N_8625);
xnor U9306 (N_9306,N_8107,N_8782);
nand U9307 (N_9307,N_8310,N_8422);
xor U9308 (N_9308,N_8078,N_8165);
xnor U9309 (N_9309,N_8759,N_8796);
or U9310 (N_9310,N_8624,N_8213);
nand U9311 (N_9311,N_8029,N_8854);
nand U9312 (N_9312,N_8325,N_8652);
nand U9313 (N_9313,N_8825,N_8008);
and U9314 (N_9314,N_8448,N_8056);
nand U9315 (N_9315,N_8231,N_8351);
nor U9316 (N_9316,N_8239,N_8643);
nand U9317 (N_9317,N_8419,N_8924);
nor U9318 (N_9318,N_8212,N_8019);
and U9319 (N_9319,N_8185,N_8814);
and U9320 (N_9320,N_8152,N_8092);
nand U9321 (N_9321,N_8951,N_8851);
nor U9322 (N_9322,N_8410,N_8018);
or U9323 (N_9323,N_8211,N_8529);
or U9324 (N_9324,N_8573,N_8906);
nor U9325 (N_9325,N_8472,N_8792);
nor U9326 (N_9326,N_8151,N_8613);
and U9327 (N_9327,N_8967,N_8178);
or U9328 (N_9328,N_8534,N_8161);
nand U9329 (N_9329,N_8296,N_8767);
or U9330 (N_9330,N_8973,N_8683);
nand U9331 (N_9331,N_8556,N_8271);
nand U9332 (N_9332,N_8189,N_8431);
xnor U9333 (N_9333,N_8521,N_8963);
or U9334 (N_9334,N_8274,N_8986);
xor U9335 (N_9335,N_8186,N_8370);
or U9336 (N_9336,N_8536,N_8552);
nand U9337 (N_9337,N_8069,N_8420);
xnor U9338 (N_9338,N_8995,N_8540);
nor U9339 (N_9339,N_8315,N_8246);
xnor U9340 (N_9340,N_8354,N_8880);
nand U9341 (N_9341,N_8440,N_8832);
nor U9342 (N_9342,N_8833,N_8279);
or U9343 (N_9343,N_8349,N_8941);
nand U9344 (N_9344,N_8343,N_8265);
nor U9345 (N_9345,N_8105,N_8174);
or U9346 (N_9346,N_8588,N_8252);
xnor U9347 (N_9347,N_8163,N_8687);
nand U9348 (N_9348,N_8456,N_8611);
and U9349 (N_9349,N_8207,N_8644);
nor U9350 (N_9350,N_8565,N_8173);
nand U9351 (N_9351,N_8817,N_8896);
xor U9352 (N_9352,N_8596,N_8388);
nor U9353 (N_9353,N_8991,N_8079);
xor U9354 (N_9354,N_8925,N_8445);
nand U9355 (N_9355,N_8345,N_8670);
or U9356 (N_9356,N_8676,N_8071);
nand U9357 (N_9357,N_8706,N_8610);
xor U9358 (N_9358,N_8690,N_8489);
nand U9359 (N_9359,N_8547,N_8134);
nor U9360 (N_9360,N_8305,N_8096);
and U9361 (N_9361,N_8795,N_8757);
and U9362 (N_9362,N_8498,N_8708);
nor U9363 (N_9363,N_8234,N_8365);
and U9364 (N_9364,N_8086,N_8778);
nor U9365 (N_9365,N_8208,N_8805);
xor U9366 (N_9366,N_8642,N_8591);
nor U9367 (N_9367,N_8038,N_8946);
or U9368 (N_9368,N_8273,N_8802);
nor U9369 (N_9369,N_8386,N_8409);
or U9370 (N_9370,N_8313,N_8740);
nor U9371 (N_9371,N_8119,N_8230);
or U9372 (N_9372,N_8374,N_8737);
xnor U9373 (N_9373,N_8505,N_8700);
and U9374 (N_9374,N_8124,N_8889);
and U9375 (N_9375,N_8934,N_8938);
or U9376 (N_9376,N_8048,N_8672);
nor U9377 (N_9377,N_8214,N_8525);
and U9378 (N_9378,N_8429,N_8160);
nand U9379 (N_9379,N_8449,N_8631);
nand U9380 (N_9380,N_8113,N_8857);
nor U9381 (N_9381,N_8299,N_8844);
and U9382 (N_9382,N_8392,N_8137);
nor U9383 (N_9383,N_8878,N_8028);
or U9384 (N_9384,N_8240,N_8490);
or U9385 (N_9385,N_8376,N_8799);
nand U9386 (N_9386,N_8574,N_8726);
xnor U9387 (N_9387,N_8742,N_8659);
nand U9388 (N_9388,N_8936,N_8121);
nand U9389 (N_9389,N_8598,N_8082);
xor U9390 (N_9390,N_8944,N_8450);
and U9391 (N_9391,N_8734,N_8807);
or U9392 (N_9392,N_8159,N_8476);
and U9393 (N_9393,N_8188,N_8426);
xor U9394 (N_9394,N_8247,N_8803);
xor U9395 (N_9395,N_8800,N_8705);
nor U9396 (N_9396,N_8870,N_8375);
or U9397 (N_9397,N_8091,N_8839);
or U9398 (N_9398,N_8290,N_8280);
xor U9399 (N_9399,N_8369,N_8108);
or U9400 (N_9400,N_8266,N_8353);
and U9401 (N_9401,N_8579,N_8000);
and U9402 (N_9402,N_8606,N_8017);
nand U9403 (N_9403,N_8719,N_8193);
or U9404 (N_9404,N_8398,N_8702);
and U9405 (N_9405,N_8637,N_8862);
and U9406 (N_9406,N_8972,N_8533);
and U9407 (N_9407,N_8526,N_8321);
nor U9408 (N_9408,N_8127,N_8763);
nor U9409 (N_9409,N_8629,N_8205);
or U9410 (N_9410,N_8987,N_8650);
xnor U9411 (N_9411,N_8751,N_8743);
or U9412 (N_9412,N_8557,N_8047);
nand U9413 (N_9413,N_8566,N_8920);
nand U9414 (N_9414,N_8543,N_8846);
nand U9415 (N_9415,N_8790,N_8678);
nand U9416 (N_9416,N_8428,N_8293);
and U9417 (N_9417,N_8387,N_8201);
nand U9418 (N_9418,N_8736,N_8709);
and U9419 (N_9419,N_8639,N_8359);
nand U9420 (N_9420,N_8224,N_8766);
or U9421 (N_9421,N_8617,N_8249);
nand U9422 (N_9422,N_8949,N_8788);
and U9423 (N_9423,N_8897,N_8150);
xnor U9424 (N_9424,N_8830,N_8933);
nand U9425 (N_9425,N_8232,N_8493);
and U9426 (N_9426,N_8834,N_8407);
nand U9427 (N_9427,N_8553,N_8822);
xnor U9428 (N_9428,N_8416,N_8550);
or U9429 (N_9429,N_8964,N_8978);
and U9430 (N_9430,N_8452,N_8992);
nor U9431 (N_9431,N_8284,N_8888);
and U9432 (N_9432,N_8746,N_8682);
nor U9433 (N_9433,N_8691,N_8154);
nor U9434 (N_9434,N_8927,N_8135);
xnor U9435 (N_9435,N_8460,N_8324);
nor U9436 (N_9436,N_8356,N_8875);
and U9437 (N_9437,N_8210,N_8061);
and U9438 (N_9438,N_8771,N_8301);
nor U9439 (N_9439,N_8196,N_8304);
nor U9440 (N_9440,N_8984,N_8628);
xnor U9441 (N_9441,N_8715,N_8909);
and U9442 (N_9442,N_8468,N_8360);
or U9443 (N_9443,N_8640,N_8182);
nand U9444 (N_9444,N_8012,N_8133);
xnor U9445 (N_9445,N_8287,N_8104);
nor U9446 (N_9446,N_8571,N_8421);
xnor U9447 (N_9447,N_8255,N_8204);
or U9448 (N_9448,N_8810,N_8563);
xnor U9449 (N_9449,N_8770,N_8312);
and U9450 (N_9450,N_8453,N_8278);
or U9451 (N_9451,N_8289,N_8381);
and U9452 (N_9452,N_8226,N_8394);
xnor U9453 (N_9453,N_8959,N_8838);
xnor U9454 (N_9454,N_8467,N_8569);
or U9455 (N_9455,N_8664,N_8753);
xnor U9456 (N_9456,N_8680,N_8042);
nand U9457 (N_9457,N_8837,N_8085);
nand U9458 (N_9458,N_8815,N_8262);
xnor U9459 (N_9459,N_8130,N_8718);
and U9460 (N_9460,N_8358,N_8479);
nand U9461 (N_9461,N_8067,N_8781);
nor U9462 (N_9462,N_8126,N_8633);
nor U9463 (N_9463,N_8257,N_8034);
nor U9464 (N_9464,N_8180,N_8887);
nand U9465 (N_9465,N_8883,N_8835);
xor U9466 (N_9466,N_8011,N_8335);
nand U9467 (N_9467,N_8361,N_8461);
nor U9468 (N_9468,N_8125,N_8913);
xor U9469 (N_9469,N_8898,N_8340);
nand U9470 (N_9470,N_8075,N_8496);
and U9471 (N_9471,N_8590,N_8957);
or U9472 (N_9472,N_8102,N_8227);
and U9473 (N_9473,N_8915,N_8408);
nand U9474 (N_9474,N_8384,N_8088);
nor U9475 (N_9475,N_8760,N_8969);
and U9476 (N_9476,N_8756,N_8465);
or U9477 (N_9477,N_8528,N_8466);
nand U9478 (N_9478,N_8905,N_8942);
xor U9479 (N_9479,N_8735,N_8323);
xnor U9480 (N_9480,N_8423,N_8926);
or U9481 (N_9481,N_8250,N_8367);
xor U9482 (N_9482,N_8039,N_8786);
nand U9483 (N_9483,N_8635,N_8393);
xor U9484 (N_9484,N_8873,N_8776);
and U9485 (N_9485,N_8309,N_8634);
xor U9486 (N_9486,N_8006,N_8364);
and U9487 (N_9487,N_8206,N_8215);
or U9488 (N_9488,N_8020,N_8236);
or U9489 (N_9489,N_8780,N_8462);
xnor U9490 (N_9490,N_8242,N_8435);
nand U9491 (N_9491,N_8379,N_8402);
or U9492 (N_9492,N_8589,N_8399);
or U9493 (N_9493,N_8877,N_8711);
nor U9494 (N_9494,N_8804,N_8859);
nand U9495 (N_9495,N_8281,N_8919);
and U9496 (N_9496,N_8966,N_8083);
nor U9497 (N_9497,N_8382,N_8258);
or U9498 (N_9498,N_8677,N_8446);
or U9499 (N_9499,N_8099,N_8021);
and U9500 (N_9500,N_8743,N_8336);
xor U9501 (N_9501,N_8787,N_8896);
xnor U9502 (N_9502,N_8069,N_8296);
or U9503 (N_9503,N_8273,N_8785);
nand U9504 (N_9504,N_8457,N_8357);
nand U9505 (N_9505,N_8047,N_8753);
or U9506 (N_9506,N_8076,N_8777);
nand U9507 (N_9507,N_8292,N_8555);
xnor U9508 (N_9508,N_8634,N_8933);
nor U9509 (N_9509,N_8016,N_8413);
nor U9510 (N_9510,N_8535,N_8150);
xor U9511 (N_9511,N_8052,N_8158);
nand U9512 (N_9512,N_8520,N_8155);
or U9513 (N_9513,N_8327,N_8639);
nor U9514 (N_9514,N_8990,N_8800);
and U9515 (N_9515,N_8796,N_8534);
xnor U9516 (N_9516,N_8551,N_8199);
or U9517 (N_9517,N_8860,N_8801);
nand U9518 (N_9518,N_8083,N_8756);
nor U9519 (N_9519,N_8302,N_8752);
nand U9520 (N_9520,N_8896,N_8135);
xnor U9521 (N_9521,N_8929,N_8909);
or U9522 (N_9522,N_8171,N_8257);
or U9523 (N_9523,N_8338,N_8823);
and U9524 (N_9524,N_8046,N_8503);
nor U9525 (N_9525,N_8847,N_8576);
nor U9526 (N_9526,N_8157,N_8845);
nand U9527 (N_9527,N_8067,N_8233);
or U9528 (N_9528,N_8741,N_8268);
xor U9529 (N_9529,N_8696,N_8450);
and U9530 (N_9530,N_8980,N_8083);
nor U9531 (N_9531,N_8921,N_8722);
xor U9532 (N_9532,N_8172,N_8168);
and U9533 (N_9533,N_8963,N_8129);
and U9534 (N_9534,N_8876,N_8934);
nand U9535 (N_9535,N_8711,N_8952);
xor U9536 (N_9536,N_8644,N_8729);
nand U9537 (N_9537,N_8580,N_8284);
nand U9538 (N_9538,N_8348,N_8788);
nor U9539 (N_9539,N_8324,N_8071);
xnor U9540 (N_9540,N_8960,N_8050);
and U9541 (N_9541,N_8490,N_8013);
and U9542 (N_9542,N_8715,N_8460);
xor U9543 (N_9543,N_8934,N_8299);
xnor U9544 (N_9544,N_8824,N_8999);
nor U9545 (N_9545,N_8541,N_8369);
nor U9546 (N_9546,N_8075,N_8741);
xnor U9547 (N_9547,N_8204,N_8450);
xor U9548 (N_9548,N_8606,N_8321);
nor U9549 (N_9549,N_8707,N_8664);
or U9550 (N_9550,N_8155,N_8091);
xnor U9551 (N_9551,N_8476,N_8905);
or U9552 (N_9552,N_8356,N_8325);
or U9553 (N_9553,N_8893,N_8062);
or U9554 (N_9554,N_8619,N_8478);
nand U9555 (N_9555,N_8238,N_8125);
or U9556 (N_9556,N_8537,N_8097);
xor U9557 (N_9557,N_8123,N_8638);
nor U9558 (N_9558,N_8010,N_8564);
nand U9559 (N_9559,N_8616,N_8337);
nand U9560 (N_9560,N_8114,N_8434);
xor U9561 (N_9561,N_8755,N_8986);
or U9562 (N_9562,N_8136,N_8938);
and U9563 (N_9563,N_8113,N_8288);
nand U9564 (N_9564,N_8280,N_8571);
nor U9565 (N_9565,N_8945,N_8552);
xor U9566 (N_9566,N_8648,N_8380);
nand U9567 (N_9567,N_8929,N_8082);
nor U9568 (N_9568,N_8138,N_8042);
xnor U9569 (N_9569,N_8776,N_8703);
nor U9570 (N_9570,N_8781,N_8601);
nor U9571 (N_9571,N_8968,N_8475);
and U9572 (N_9572,N_8401,N_8510);
xnor U9573 (N_9573,N_8856,N_8942);
and U9574 (N_9574,N_8229,N_8238);
or U9575 (N_9575,N_8517,N_8147);
nor U9576 (N_9576,N_8432,N_8328);
and U9577 (N_9577,N_8698,N_8141);
nand U9578 (N_9578,N_8750,N_8308);
xnor U9579 (N_9579,N_8644,N_8092);
and U9580 (N_9580,N_8999,N_8203);
or U9581 (N_9581,N_8627,N_8407);
nor U9582 (N_9582,N_8381,N_8614);
nor U9583 (N_9583,N_8528,N_8899);
xnor U9584 (N_9584,N_8799,N_8593);
and U9585 (N_9585,N_8674,N_8550);
or U9586 (N_9586,N_8787,N_8018);
xnor U9587 (N_9587,N_8717,N_8917);
nand U9588 (N_9588,N_8802,N_8397);
nor U9589 (N_9589,N_8979,N_8953);
xnor U9590 (N_9590,N_8519,N_8409);
or U9591 (N_9591,N_8637,N_8370);
nand U9592 (N_9592,N_8573,N_8461);
nand U9593 (N_9593,N_8860,N_8298);
nor U9594 (N_9594,N_8568,N_8882);
nor U9595 (N_9595,N_8271,N_8275);
nand U9596 (N_9596,N_8781,N_8510);
or U9597 (N_9597,N_8296,N_8254);
and U9598 (N_9598,N_8825,N_8355);
or U9599 (N_9599,N_8451,N_8702);
and U9600 (N_9600,N_8616,N_8630);
nand U9601 (N_9601,N_8418,N_8286);
nand U9602 (N_9602,N_8716,N_8150);
or U9603 (N_9603,N_8900,N_8162);
nor U9604 (N_9604,N_8416,N_8712);
or U9605 (N_9605,N_8746,N_8396);
nand U9606 (N_9606,N_8180,N_8423);
nor U9607 (N_9607,N_8166,N_8874);
or U9608 (N_9608,N_8862,N_8010);
nor U9609 (N_9609,N_8785,N_8219);
nand U9610 (N_9610,N_8798,N_8663);
xnor U9611 (N_9611,N_8815,N_8400);
nand U9612 (N_9612,N_8698,N_8652);
and U9613 (N_9613,N_8689,N_8832);
or U9614 (N_9614,N_8470,N_8129);
and U9615 (N_9615,N_8304,N_8451);
nor U9616 (N_9616,N_8975,N_8163);
or U9617 (N_9617,N_8094,N_8343);
or U9618 (N_9618,N_8001,N_8704);
and U9619 (N_9619,N_8844,N_8201);
xnor U9620 (N_9620,N_8839,N_8740);
and U9621 (N_9621,N_8728,N_8130);
nor U9622 (N_9622,N_8132,N_8293);
and U9623 (N_9623,N_8374,N_8238);
nand U9624 (N_9624,N_8039,N_8222);
nand U9625 (N_9625,N_8839,N_8975);
or U9626 (N_9626,N_8971,N_8452);
xnor U9627 (N_9627,N_8854,N_8008);
nand U9628 (N_9628,N_8865,N_8692);
nand U9629 (N_9629,N_8198,N_8078);
nand U9630 (N_9630,N_8630,N_8503);
nor U9631 (N_9631,N_8626,N_8664);
nor U9632 (N_9632,N_8629,N_8291);
and U9633 (N_9633,N_8097,N_8336);
nand U9634 (N_9634,N_8008,N_8193);
xor U9635 (N_9635,N_8391,N_8971);
or U9636 (N_9636,N_8290,N_8981);
or U9637 (N_9637,N_8356,N_8121);
or U9638 (N_9638,N_8812,N_8023);
nor U9639 (N_9639,N_8517,N_8685);
xor U9640 (N_9640,N_8864,N_8324);
nor U9641 (N_9641,N_8722,N_8056);
or U9642 (N_9642,N_8806,N_8095);
xnor U9643 (N_9643,N_8963,N_8006);
and U9644 (N_9644,N_8656,N_8315);
nor U9645 (N_9645,N_8971,N_8577);
xnor U9646 (N_9646,N_8818,N_8839);
nor U9647 (N_9647,N_8955,N_8883);
xor U9648 (N_9648,N_8009,N_8462);
xor U9649 (N_9649,N_8405,N_8936);
or U9650 (N_9650,N_8799,N_8583);
and U9651 (N_9651,N_8823,N_8739);
or U9652 (N_9652,N_8047,N_8829);
or U9653 (N_9653,N_8064,N_8728);
xnor U9654 (N_9654,N_8889,N_8780);
and U9655 (N_9655,N_8598,N_8261);
nor U9656 (N_9656,N_8774,N_8777);
and U9657 (N_9657,N_8048,N_8541);
or U9658 (N_9658,N_8736,N_8876);
nand U9659 (N_9659,N_8553,N_8241);
nand U9660 (N_9660,N_8318,N_8957);
or U9661 (N_9661,N_8419,N_8621);
xor U9662 (N_9662,N_8754,N_8215);
and U9663 (N_9663,N_8669,N_8246);
and U9664 (N_9664,N_8084,N_8804);
nor U9665 (N_9665,N_8680,N_8475);
or U9666 (N_9666,N_8773,N_8906);
nand U9667 (N_9667,N_8348,N_8066);
xor U9668 (N_9668,N_8298,N_8304);
nand U9669 (N_9669,N_8943,N_8103);
xnor U9670 (N_9670,N_8044,N_8370);
nand U9671 (N_9671,N_8897,N_8660);
or U9672 (N_9672,N_8682,N_8060);
nor U9673 (N_9673,N_8795,N_8303);
nand U9674 (N_9674,N_8953,N_8994);
nor U9675 (N_9675,N_8587,N_8420);
xor U9676 (N_9676,N_8703,N_8541);
or U9677 (N_9677,N_8246,N_8249);
and U9678 (N_9678,N_8696,N_8966);
nand U9679 (N_9679,N_8509,N_8927);
nor U9680 (N_9680,N_8165,N_8943);
nor U9681 (N_9681,N_8643,N_8629);
nor U9682 (N_9682,N_8260,N_8429);
nor U9683 (N_9683,N_8066,N_8045);
nor U9684 (N_9684,N_8357,N_8785);
nor U9685 (N_9685,N_8059,N_8132);
and U9686 (N_9686,N_8087,N_8998);
or U9687 (N_9687,N_8390,N_8639);
or U9688 (N_9688,N_8501,N_8733);
or U9689 (N_9689,N_8854,N_8130);
nor U9690 (N_9690,N_8440,N_8875);
nor U9691 (N_9691,N_8040,N_8524);
xnor U9692 (N_9692,N_8020,N_8692);
and U9693 (N_9693,N_8514,N_8884);
xnor U9694 (N_9694,N_8051,N_8306);
nor U9695 (N_9695,N_8552,N_8112);
or U9696 (N_9696,N_8420,N_8044);
nor U9697 (N_9697,N_8717,N_8061);
or U9698 (N_9698,N_8005,N_8632);
or U9699 (N_9699,N_8156,N_8826);
nor U9700 (N_9700,N_8987,N_8106);
or U9701 (N_9701,N_8429,N_8013);
nor U9702 (N_9702,N_8665,N_8456);
nand U9703 (N_9703,N_8017,N_8762);
nand U9704 (N_9704,N_8976,N_8260);
nor U9705 (N_9705,N_8750,N_8500);
xnor U9706 (N_9706,N_8557,N_8739);
nand U9707 (N_9707,N_8183,N_8546);
or U9708 (N_9708,N_8474,N_8276);
nor U9709 (N_9709,N_8023,N_8598);
and U9710 (N_9710,N_8411,N_8558);
or U9711 (N_9711,N_8581,N_8586);
and U9712 (N_9712,N_8767,N_8329);
nand U9713 (N_9713,N_8290,N_8251);
nand U9714 (N_9714,N_8013,N_8940);
and U9715 (N_9715,N_8008,N_8200);
nand U9716 (N_9716,N_8650,N_8064);
or U9717 (N_9717,N_8971,N_8207);
nand U9718 (N_9718,N_8783,N_8300);
nand U9719 (N_9719,N_8721,N_8246);
nand U9720 (N_9720,N_8482,N_8739);
xor U9721 (N_9721,N_8779,N_8925);
nor U9722 (N_9722,N_8087,N_8272);
xnor U9723 (N_9723,N_8437,N_8746);
nand U9724 (N_9724,N_8536,N_8628);
or U9725 (N_9725,N_8971,N_8609);
nor U9726 (N_9726,N_8774,N_8061);
xor U9727 (N_9727,N_8728,N_8471);
xnor U9728 (N_9728,N_8037,N_8363);
xnor U9729 (N_9729,N_8959,N_8002);
and U9730 (N_9730,N_8812,N_8154);
nand U9731 (N_9731,N_8169,N_8987);
or U9732 (N_9732,N_8764,N_8816);
nand U9733 (N_9733,N_8475,N_8805);
nand U9734 (N_9734,N_8044,N_8708);
or U9735 (N_9735,N_8725,N_8078);
and U9736 (N_9736,N_8547,N_8757);
and U9737 (N_9737,N_8765,N_8732);
xnor U9738 (N_9738,N_8602,N_8565);
xnor U9739 (N_9739,N_8476,N_8478);
nand U9740 (N_9740,N_8204,N_8310);
or U9741 (N_9741,N_8710,N_8349);
and U9742 (N_9742,N_8785,N_8866);
nand U9743 (N_9743,N_8542,N_8748);
nor U9744 (N_9744,N_8970,N_8774);
nor U9745 (N_9745,N_8330,N_8709);
xnor U9746 (N_9746,N_8601,N_8545);
nor U9747 (N_9747,N_8142,N_8783);
and U9748 (N_9748,N_8081,N_8339);
nor U9749 (N_9749,N_8615,N_8000);
and U9750 (N_9750,N_8538,N_8403);
xor U9751 (N_9751,N_8311,N_8567);
or U9752 (N_9752,N_8136,N_8880);
or U9753 (N_9753,N_8984,N_8178);
xnor U9754 (N_9754,N_8771,N_8273);
nand U9755 (N_9755,N_8299,N_8498);
and U9756 (N_9756,N_8788,N_8770);
nor U9757 (N_9757,N_8683,N_8128);
nor U9758 (N_9758,N_8542,N_8976);
nand U9759 (N_9759,N_8117,N_8702);
xor U9760 (N_9760,N_8101,N_8181);
xor U9761 (N_9761,N_8267,N_8835);
nor U9762 (N_9762,N_8508,N_8167);
xnor U9763 (N_9763,N_8949,N_8526);
nor U9764 (N_9764,N_8160,N_8224);
xor U9765 (N_9765,N_8077,N_8226);
and U9766 (N_9766,N_8994,N_8917);
xor U9767 (N_9767,N_8586,N_8143);
or U9768 (N_9768,N_8445,N_8259);
nor U9769 (N_9769,N_8143,N_8021);
xnor U9770 (N_9770,N_8254,N_8258);
nor U9771 (N_9771,N_8070,N_8697);
nor U9772 (N_9772,N_8386,N_8924);
or U9773 (N_9773,N_8178,N_8553);
nor U9774 (N_9774,N_8225,N_8951);
nor U9775 (N_9775,N_8855,N_8324);
nand U9776 (N_9776,N_8981,N_8578);
and U9777 (N_9777,N_8792,N_8418);
nand U9778 (N_9778,N_8822,N_8500);
and U9779 (N_9779,N_8943,N_8157);
and U9780 (N_9780,N_8632,N_8246);
or U9781 (N_9781,N_8255,N_8874);
xnor U9782 (N_9782,N_8043,N_8096);
xnor U9783 (N_9783,N_8185,N_8533);
xnor U9784 (N_9784,N_8436,N_8856);
or U9785 (N_9785,N_8337,N_8452);
xor U9786 (N_9786,N_8363,N_8137);
and U9787 (N_9787,N_8721,N_8203);
nand U9788 (N_9788,N_8335,N_8960);
nand U9789 (N_9789,N_8407,N_8320);
xor U9790 (N_9790,N_8641,N_8816);
and U9791 (N_9791,N_8500,N_8122);
or U9792 (N_9792,N_8990,N_8807);
and U9793 (N_9793,N_8651,N_8164);
or U9794 (N_9794,N_8953,N_8036);
nor U9795 (N_9795,N_8918,N_8212);
nor U9796 (N_9796,N_8358,N_8881);
or U9797 (N_9797,N_8413,N_8446);
or U9798 (N_9798,N_8971,N_8731);
and U9799 (N_9799,N_8764,N_8280);
or U9800 (N_9800,N_8232,N_8636);
nand U9801 (N_9801,N_8992,N_8519);
nor U9802 (N_9802,N_8149,N_8264);
nor U9803 (N_9803,N_8210,N_8234);
or U9804 (N_9804,N_8600,N_8079);
and U9805 (N_9805,N_8469,N_8694);
nor U9806 (N_9806,N_8829,N_8027);
nand U9807 (N_9807,N_8618,N_8730);
and U9808 (N_9808,N_8861,N_8097);
or U9809 (N_9809,N_8619,N_8262);
or U9810 (N_9810,N_8860,N_8452);
nand U9811 (N_9811,N_8166,N_8255);
and U9812 (N_9812,N_8827,N_8514);
or U9813 (N_9813,N_8110,N_8631);
xor U9814 (N_9814,N_8768,N_8703);
xnor U9815 (N_9815,N_8155,N_8454);
xnor U9816 (N_9816,N_8575,N_8179);
nand U9817 (N_9817,N_8514,N_8832);
nor U9818 (N_9818,N_8917,N_8209);
nor U9819 (N_9819,N_8694,N_8413);
nand U9820 (N_9820,N_8606,N_8884);
and U9821 (N_9821,N_8038,N_8011);
xor U9822 (N_9822,N_8215,N_8040);
nand U9823 (N_9823,N_8346,N_8400);
xor U9824 (N_9824,N_8481,N_8766);
and U9825 (N_9825,N_8806,N_8791);
or U9826 (N_9826,N_8305,N_8159);
nand U9827 (N_9827,N_8911,N_8024);
nand U9828 (N_9828,N_8387,N_8285);
and U9829 (N_9829,N_8508,N_8621);
nor U9830 (N_9830,N_8260,N_8890);
or U9831 (N_9831,N_8269,N_8877);
and U9832 (N_9832,N_8812,N_8466);
xnor U9833 (N_9833,N_8041,N_8635);
or U9834 (N_9834,N_8441,N_8702);
xnor U9835 (N_9835,N_8348,N_8972);
or U9836 (N_9836,N_8674,N_8917);
xor U9837 (N_9837,N_8821,N_8964);
nor U9838 (N_9838,N_8759,N_8139);
xnor U9839 (N_9839,N_8716,N_8996);
or U9840 (N_9840,N_8100,N_8399);
or U9841 (N_9841,N_8207,N_8472);
nor U9842 (N_9842,N_8204,N_8456);
and U9843 (N_9843,N_8603,N_8149);
nand U9844 (N_9844,N_8373,N_8564);
or U9845 (N_9845,N_8044,N_8382);
xor U9846 (N_9846,N_8675,N_8311);
nand U9847 (N_9847,N_8737,N_8848);
or U9848 (N_9848,N_8257,N_8670);
nand U9849 (N_9849,N_8137,N_8160);
nand U9850 (N_9850,N_8904,N_8689);
xnor U9851 (N_9851,N_8388,N_8639);
and U9852 (N_9852,N_8684,N_8193);
nor U9853 (N_9853,N_8905,N_8090);
nand U9854 (N_9854,N_8687,N_8189);
xor U9855 (N_9855,N_8940,N_8419);
xnor U9856 (N_9856,N_8603,N_8369);
and U9857 (N_9857,N_8684,N_8053);
and U9858 (N_9858,N_8957,N_8912);
and U9859 (N_9859,N_8714,N_8777);
nand U9860 (N_9860,N_8287,N_8203);
nor U9861 (N_9861,N_8065,N_8279);
nand U9862 (N_9862,N_8954,N_8787);
nand U9863 (N_9863,N_8311,N_8469);
nor U9864 (N_9864,N_8643,N_8947);
nand U9865 (N_9865,N_8539,N_8321);
xor U9866 (N_9866,N_8209,N_8101);
nand U9867 (N_9867,N_8525,N_8902);
and U9868 (N_9868,N_8380,N_8025);
and U9869 (N_9869,N_8284,N_8626);
and U9870 (N_9870,N_8968,N_8895);
xor U9871 (N_9871,N_8637,N_8884);
nor U9872 (N_9872,N_8677,N_8265);
nand U9873 (N_9873,N_8820,N_8364);
nand U9874 (N_9874,N_8712,N_8846);
or U9875 (N_9875,N_8569,N_8597);
nor U9876 (N_9876,N_8798,N_8761);
nor U9877 (N_9877,N_8354,N_8082);
xnor U9878 (N_9878,N_8558,N_8419);
or U9879 (N_9879,N_8347,N_8800);
and U9880 (N_9880,N_8148,N_8736);
and U9881 (N_9881,N_8978,N_8309);
nand U9882 (N_9882,N_8249,N_8607);
and U9883 (N_9883,N_8946,N_8204);
xnor U9884 (N_9884,N_8508,N_8722);
xnor U9885 (N_9885,N_8551,N_8779);
nor U9886 (N_9886,N_8836,N_8688);
nand U9887 (N_9887,N_8527,N_8232);
nor U9888 (N_9888,N_8376,N_8102);
nor U9889 (N_9889,N_8719,N_8953);
nor U9890 (N_9890,N_8538,N_8586);
and U9891 (N_9891,N_8417,N_8256);
or U9892 (N_9892,N_8056,N_8813);
and U9893 (N_9893,N_8021,N_8384);
nor U9894 (N_9894,N_8801,N_8398);
and U9895 (N_9895,N_8693,N_8168);
nor U9896 (N_9896,N_8326,N_8860);
nand U9897 (N_9897,N_8835,N_8226);
and U9898 (N_9898,N_8394,N_8635);
or U9899 (N_9899,N_8437,N_8743);
xor U9900 (N_9900,N_8961,N_8494);
xor U9901 (N_9901,N_8390,N_8658);
or U9902 (N_9902,N_8951,N_8825);
or U9903 (N_9903,N_8211,N_8214);
and U9904 (N_9904,N_8218,N_8649);
nor U9905 (N_9905,N_8062,N_8404);
xor U9906 (N_9906,N_8143,N_8418);
nor U9907 (N_9907,N_8103,N_8802);
or U9908 (N_9908,N_8857,N_8670);
nand U9909 (N_9909,N_8967,N_8959);
or U9910 (N_9910,N_8054,N_8582);
nand U9911 (N_9911,N_8649,N_8283);
or U9912 (N_9912,N_8444,N_8763);
or U9913 (N_9913,N_8132,N_8885);
or U9914 (N_9914,N_8189,N_8294);
and U9915 (N_9915,N_8577,N_8718);
nand U9916 (N_9916,N_8951,N_8661);
and U9917 (N_9917,N_8993,N_8532);
or U9918 (N_9918,N_8800,N_8213);
nand U9919 (N_9919,N_8747,N_8011);
xor U9920 (N_9920,N_8077,N_8799);
or U9921 (N_9921,N_8757,N_8329);
and U9922 (N_9922,N_8501,N_8827);
nor U9923 (N_9923,N_8546,N_8430);
xor U9924 (N_9924,N_8580,N_8231);
or U9925 (N_9925,N_8232,N_8443);
and U9926 (N_9926,N_8159,N_8917);
and U9927 (N_9927,N_8819,N_8418);
or U9928 (N_9928,N_8703,N_8143);
nand U9929 (N_9929,N_8507,N_8324);
or U9930 (N_9930,N_8386,N_8621);
or U9931 (N_9931,N_8483,N_8643);
nand U9932 (N_9932,N_8233,N_8222);
or U9933 (N_9933,N_8961,N_8527);
nor U9934 (N_9934,N_8024,N_8189);
xor U9935 (N_9935,N_8013,N_8037);
nand U9936 (N_9936,N_8935,N_8768);
nor U9937 (N_9937,N_8313,N_8735);
nand U9938 (N_9938,N_8942,N_8921);
and U9939 (N_9939,N_8884,N_8974);
nor U9940 (N_9940,N_8931,N_8147);
and U9941 (N_9941,N_8407,N_8046);
or U9942 (N_9942,N_8209,N_8093);
or U9943 (N_9943,N_8329,N_8476);
nor U9944 (N_9944,N_8589,N_8438);
and U9945 (N_9945,N_8706,N_8444);
nand U9946 (N_9946,N_8326,N_8952);
nor U9947 (N_9947,N_8066,N_8892);
or U9948 (N_9948,N_8089,N_8378);
nor U9949 (N_9949,N_8951,N_8658);
or U9950 (N_9950,N_8461,N_8675);
nor U9951 (N_9951,N_8131,N_8679);
nor U9952 (N_9952,N_8295,N_8340);
nor U9953 (N_9953,N_8264,N_8860);
or U9954 (N_9954,N_8698,N_8281);
and U9955 (N_9955,N_8608,N_8939);
nand U9956 (N_9956,N_8002,N_8780);
and U9957 (N_9957,N_8233,N_8025);
and U9958 (N_9958,N_8971,N_8034);
xor U9959 (N_9959,N_8573,N_8050);
nor U9960 (N_9960,N_8623,N_8490);
nor U9961 (N_9961,N_8797,N_8069);
nor U9962 (N_9962,N_8804,N_8831);
xor U9963 (N_9963,N_8175,N_8672);
or U9964 (N_9964,N_8082,N_8117);
nand U9965 (N_9965,N_8488,N_8881);
xnor U9966 (N_9966,N_8514,N_8959);
nand U9967 (N_9967,N_8056,N_8175);
xnor U9968 (N_9968,N_8758,N_8952);
or U9969 (N_9969,N_8992,N_8294);
or U9970 (N_9970,N_8885,N_8741);
nand U9971 (N_9971,N_8700,N_8796);
and U9972 (N_9972,N_8576,N_8991);
xor U9973 (N_9973,N_8543,N_8628);
nand U9974 (N_9974,N_8356,N_8221);
nand U9975 (N_9975,N_8185,N_8540);
nand U9976 (N_9976,N_8063,N_8100);
nand U9977 (N_9977,N_8669,N_8506);
nand U9978 (N_9978,N_8682,N_8236);
nand U9979 (N_9979,N_8468,N_8973);
xnor U9980 (N_9980,N_8471,N_8651);
or U9981 (N_9981,N_8271,N_8282);
or U9982 (N_9982,N_8045,N_8371);
xor U9983 (N_9983,N_8612,N_8394);
or U9984 (N_9984,N_8074,N_8643);
xor U9985 (N_9985,N_8159,N_8021);
nor U9986 (N_9986,N_8961,N_8966);
xor U9987 (N_9987,N_8413,N_8188);
nand U9988 (N_9988,N_8145,N_8535);
and U9989 (N_9989,N_8865,N_8930);
nor U9990 (N_9990,N_8757,N_8803);
nor U9991 (N_9991,N_8091,N_8396);
nor U9992 (N_9992,N_8080,N_8863);
and U9993 (N_9993,N_8473,N_8593);
xor U9994 (N_9994,N_8210,N_8535);
or U9995 (N_9995,N_8755,N_8290);
nand U9996 (N_9996,N_8452,N_8101);
or U9997 (N_9997,N_8325,N_8323);
nor U9998 (N_9998,N_8016,N_8764);
nor U9999 (N_9999,N_8858,N_8004);
nand U10000 (N_10000,N_9519,N_9370);
nand U10001 (N_10001,N_9546,N_9912);
nand U10002 (N_10002,N_9385,N_9134);
nor U10003 (N_10003,N_9412,N_9976);
xor U10004 (N_10004,N_9434,N_9752);
or U10005 (N_10005,N_9941,N_9391);
nor U10006 (N_10006,N_9492,N_9486);
nor U10007 (N_10007,N_9766,N_9446);
and U10008 (N_10008,N_9871,N_9664);
nand U10009 (N_10009,N_9631,N_9720);
nand U10010 (N_10010,N_9414,N_9275);
and U10011 (N_10011,N_9255,N_9508);
nor U10012 (N_10012,N_9171,N_9571);
nand U10013 (N_10013,N_9149,N_9049);
nand U10014 (N_10014,N_9212,N_9153);
nor U10015 (N_10015,N_9621,N_9036);
and U10016 (N_10016,N_9292,N_9359);
nand U10017 (N_10017,N_9205,N_9884);
nand U10018 (N_10018,N_9395,N_9987);
xnor U10019 (N_10019,N_9407,N_9903);
nand U10020 (N_10020,N_9161,N_9151);
xor U10021 (N_10021,N_9783,N_9267);
nand U10022 (N_10022,N_9327,N_9040);
xor U10023 (N_10023,N_9892,N_9390);
xor U10024 (N_10024,N_9394,N_9488);
nor U10025 (N_10025,N_9633,N_9236);
and U10026 (N_10026,N_9551,N_9587);
or U10027 (N_10027,N_9744,N_9944);
xnor U10028 (N_10028,N_9289,N_9464);
or U10029 (N_10029,N_9355,N_9991);
or U10030 (N_10030,N_9132,N_9405);
and U10031 (N_10031,N_9600,N_9223);
xor U10032 (N_10032,N_9676,N_9023);
xnor U10033 (N_10033,N_9691,N_9636);
nor U10034 (N_10034,N_9445,N_9726);
and U10035 (N_10035,N_9938,N_9896);
or U10036 (N_10036,N_9058,N_9417);
or U10037 (N_10037,N_9831,N_9811);
nor U10038 (N_10038,N_9969,N_9942);
nand U10039 (N_10039,N_9680,N_9328);
and U10040 (N_10040,N_9876,N_9031);
nor U10041 (N_10041,N_9276,N_9886);
xor U10042 (N_10042,N_9737,N_9072);
nand U10043 (N_10043,N_9061,N_9329);
nand U10044 (N_10044,N_9823,N_9834);
nor U10045 (N_10045,N_9846,N_9813);
or U10046 (N_10046,N_9281,N_9282);
or U10047 (N_10047,N_9785,N_9772);
xor U10048 (N_10048,N_9866,N_9437);
xnor U10049 (N_10049,N_9634,N_9793);
nor U10050 (N_10050,N_9403,N_9577);
nor U10051 (N_10051,N_9699,N_9343);
and U10052 (N_10052,N_9173,N_9420);
or U10053 (N_10053,N_9812,N_9165);
nand U10054 (N_10054,N_9597,N_9917);
nor U10055 (N_10055,N_9448,N_9792);
and U10056 (N_10056,N_9684,N_9042);
or U10057 (N_10057,N_9156,N_9190);
or U10058 (N_10058,N_9207,N_9254);
nand U10059 (N_10059,N_9076,N_9294);
nand U10060 (N_10060,N_9511,N_9353);
nand U10061 (N_10061,N_9191,N_9443);
and U10062 (N_10062,N_9291,N_9230);
nor U10063 (N_10063,N_9169,N_9999);
and U10064 (N_10064,N_9761,N_9046);
xnor U10065 (N_10065,N_9543,N_9295);
nor U10066 (N_10066,N_9925,N_9142);
and U10067 (N_10067,N_9091,N_9389);
and U10068 (N_10068,N_9654,N_9650);
nand U10069 (N_10069,N_9854,N_9330);
xnor U10070 (N_10070,N_9096,N_9378);
or U10071 (N_10071,N_9313,N_9233);
and U10072 (N_10072,N_9954,N_9452);
or U10073 (N_10073,N_9364,N_9759);
nand U10074 (N_10074,N_9973,N_9369);
xnor U10075 (N_10075,N_9283,N_9714);
or U10076 (N_10076,N_9002,N_9931);
nor U10077 (N_10077,N_9086,N_9438);
xnor U10078 (N_10078,N_9174,N_9424);
or U10079 (N_10079,N_9777,N_9729);
and U10080 (N_10080,N_9979,N_9570);
or U10081 (N_10081,N_9232,N_9559);
xnor U10082 (N_10082,N_9179,N_9534);
or U10083 (N_10083,N_9731,N_9129);
xnor U10084 (N_10084,N_9008,N_9164);
nor U10085 (N_10085,N_9929,N_9399);
and U10086 (N_10086,N_9657,N_9767);
nand U10087 (N_10087,N_9272,N_9997);
or U10088 (N_10088,N_9019,N_9351);
xor U10089 (N_10089,N_9485,N_9264);
nand U10090 (N_10090,N_9248,N_9145);
and U10091 (N_10091,N_9249,N_9853);
nand U10092 (N_10092,N_9373,N_9566);
or U10093 (N_10093,N_9167,N_9933);
or U10094 (N_10094,N_9195,N_9835);
xor U10095 (N_10095,N_9743,N_9182);
nand U10096 (N_10096,N_9322,N_9116);
or U10097 (N_10097,N_9060,N_9126);
xor U10098 (N_10098,N_9995,N_9560);
nand U10099 (N_10099,N_9569,N_9415);
xor U10100 (N_10100,N_9017,N_9382);
and U10101 (N_10101,N_9316,N_9937);
xnor U10102 (N_10102,N_9050,N_9352);
or U10103 (N_10103,N_9041,N_9270);
and U10104 (N_10104,N_9655,N_9806);
xor U10105 (N_10105,N_9034,N_9895);
and U10106 (N_10106,N_9055,N_9462);
xnor U10107 (N_10107,N_9719,N_9975);
or U10108 (N_10108,N_9807,N_9221);
nor U10109 (N_10109,N_9818,N_9540);
nand U10110 (N_10110,N_9503,N_9105);
nand U10111 (N_10111,N_9111,N_9589);
nand U10112 (N_10112,N_9288,N_9647);
xnor U10113 (N_10113,N_9102,N_9709);
xor U10114 (N_10114,N_9614,N_9319);
or U10115 (N_10115,N_9079,N_9428);
or U10116 (N_10116,N_9694,N_9038);
nand U10117 (N_10117,N_9757,N_9645);
nand U10118 (N_10118,N_9368,N_9764);
nor U10119 (N_10119,N_9906,N_9943);
xnor U10120 (N_10120,N_9640,N_9756);
nor U10121 (N_10121,N_9769,N_9280);
and U10122 (N_10122,N_9686,N_9860);
or U10123 (N_10123,N_9609,N_9260);
or U10124 (N_10124,N_9572,N_9136);
nand U10125 (N_10125,N_9518,N_9606);
nand U10126 (N_10126,N_9541,N_9580);
and U10127 (N_10127,N_9423,N_9955);
xor U10128 (N_10128,N_9456,N_9748);
or U10129 (N_10129,N_9939,N_9401);
and U10130 (N_10130,N_9215,N_9977);
or U10131 (N_10131,N_9104,N_9905);
and U10132 (N_10132,N_9659,N_9039);
and U10133 (N_10133,N_9796,N_9159);
nand U10134 (N_10134,N_9004,N_9185);
nor U10135 (N_10135,N_9745,N_9338);
nand U10136 (N_10136,N_9155,N_9642);
and U10137 (N_10137,N_9583,N_9466);
and U10138 (N_10138,N_9139,N_9304);
nand U10139 (N_10139,N_9599,N_9458);
nand U10140 (N_10140,N_9472,N_9346);
nand U10141 (N_10141,N_9930,N_9422);
nand U10142 (N_10142,N_9525,N_9051);
nor U10143 (N_10143,N_9515,N_9376);
or U10144 (N_10144,N_9154,N_9475);
nor U10145 (N_10145,N_9990,N_9344);
or U10146 (N_10146,N_9323,N_9651);
nand U10147 (N_10147,N_9901,N_9106);
nand U10148 (N_10148,N_9241,N_9962);
nand U10149 (N_10149,N_9562,N_9803);
nor U10150 (N_10150,N_9468,N_9162);
nand U10151 (N_10151,N_9902,N_9801);
xor U10152 (N_10152,N_9301,N_9514);
nand U10153 (N_10153,N_9122,N_9698);
nand U10154 (N_10154,N_9791,N_9003);
or U10155 (N_10155,N_9608,N_9829);
or U10156 (N_10156,N_9591,N_9052);
xnor U10157 (N_10157,N_9605,N_9561);
xor U10158 (N_10158,N_9278,N_9348);
and U10159 (N_10159,N_9321,N_9484);
nor U10160 (N_10160,N_9697,N_9604);
or U10161 (N_10161,N_9774,N_9137);
nand U10162 (N_10162,N_9817,N_9271);
nand U10163 (N_10163,N_9457,N_9258);
or U10164 (N_10164,N_9374,N_9918);
and U10165 (N_10165,N_9203,N_9266);
nand U10166 (N_10166,N_9998,N_9277);
nand U10167 (N_10167,N_9384,N_9845);
nand U10168 (N_10168,N_9682,N_9952);
xnor U10169 (N_10169,N_9240,N_9579);
xor U10170 (N_10170,N_9163,N_9495);
nand U10171 (N_10171,N_9856,N_9778);
nand U10172 (N_10172,N_9160,N_9520);
xnor U10173 (N_10173,N_9320,N_9483);
xor U10174 (N_10174,N_9516,N_9878);
nor U10175 (N_10175,N_9213,N_9660);
nor U10176 (N_10176,N_9749,N_9784);
nand U10177 (N_10177,N_9469,N_9910);
or U10178 (N_10178,N_9765,N_9035);
or U10179 (N_10179,N_9947,N_9114);
nor U10180 (N_10180,N_9971,N_9287);
and U10181 (N_10181,N_9927,N_9147);
nor U10182 (N_10182,N_9696,N_9113);
or U10183 (N_10183,N_9493,N_9148);
nor U10184 (N_10184,N_9658,N_9265);
nor U10185 (N_10185,N_9557,N_9433);
or U10186 (N_10186,N_9689,N_9435);
nor U10187 (N_10187,N_9109,N_9668);
xnor U10188 (N_10188,N_9082,N_9187);
xor U10189 (N_10189,N_9128,N_9197);
nor U10190 (N_10190,N_9538,N_9563);
or U10191 (N_10191,N_9622,N_9883);
nor U10192 (N_10192,N_9934,N_9206);
nor U10193 (N_10193,N_9909,N_9358);
or U10194 (N_10194,N_9723,N_9945);
xnor U10195 (N_10195,N_9711,N_9891);
nor U10196 (N_10196,N_9146,N_9547);
xor U10197 (N_10197,N_9357,N_9302);
nand U10198 (N_10198,N_9926,N_9612);
nand U10199 (N_10199,N_9773,N_9099);
nand U10200 (N_10200,N_9669,N_9646);
xor U10201 (N_10201,N_9225,N_9625);
nand U10202 (N_10202,N_9112,N_9607);
nand U10203 (N_10203,N_9509,N_9377);
xor U10204 (N_10204,N_9262,N_9450);
or U10205 (N_10205,N_9297,N_9960);
or U10206 (N_10206,N_9127,N_9703);
and U10207 (N_10207,N_9582,N_9229);
nand U10208 (N_10208,N_9666,N_9740);
or U10209 (N_10209,N_9951,N_9875);
nand U10210 (N_10210,N_9734,N_9712);
xnor U10211 (N_10211,N_9054,N_9011);
nor U10212 (N_10212,N_9889,N_9471);
nor U10213 (N_10213,N_9470,N_9819);
xor U10214 (N_10214,N_9717,N_9261);
and U10215 (N_10215,N_9879,N_9226);
and U10216 (N_10216,N_9841,N_9406);
nor U10217 (N_10217,N_9652,N_9474);
xnor U10218 (N_10218,N_9674,N_9381);
xor U10219 (N_10219,N_9629,N_9386);
and U10220 (N_10220,N_9180,N_9150);
xor U10221 (N_10221,N_9594,N_9873);
nor U10222 (N_10222,N_9950,N_9269);
nor U10223 (N_10223,N_9416,N_9242);
nor U10224 (N_10224,N_9994,N_9175);
or U10225 (N_10225,N_9314,N_9168);
xnor U10226 (N_10226,N_9108,N_9836);
and U10227 (N_10227,N_9528,N_9400);
and U10228 (N_10228,N_9710,N_9649);
and U10229 (N_10229,N_9263,N_9115);
xnor U10230 (N_10230,N_9898,N_9476);
or U10231 (N_10231,N_9821,N_9965);
xor U10232 (N_10232,N_9914,N_9980);
nor U10233 (N_10233,N_9888,N_9648);
nand U10234 (N_10234,N_9628,N_9855);
nor U10235 (N_10235,N_9983,N_9393);
xor U10236 (N_10236,N_9166,N_9881);
nand U10237 (N_10237,N_9170,N_9978);
nand U10238 (N_10238,N_9363,N_9332);
and U10239 (N_10239,N_9549,N_9588);
nand U10240 (N_10240,N_9858,N_9118);
nand U10241 (N_10241,N_9045,N_9360);
and U10242 (N_10242,N_9670,N_9787);
xor U10243 (N_10243,N_9194,N_9837);
and U10244 (N_10244,N_9238,N_9981);
or U10245 (N_10245,N_9885,N_9454);
and U10246 (N_10246,N_9693,N_9497);
nor U10247 (N_10247,N_9279,N_9832);
or U10248 (N_10248,N_9618,N_9956);
or U10249 (N_10249,N_9317,N_9140);
nand U10250 (N_10250,N_9234,N_9963);
or U10251 (N_10251,N_9713,N_9820);
nor U10252 (N_10252,N_9771,N_9071);
nor U10253 (N_10253,N_9298,N_9685);
nor U10254 (N_10254,N_9808,N_9781);
nor U10255 (N_10255,N_9144,N_9198);
or U10256 (N_10256,N_9005,N_9256);
xnor U10257 (N_10257,N_9123,N_9957);
and U10258 (N_10258,N_9754,N_9887);
nor U10259 (N_10259,N_9677,N_9101);
and U10260 (N_10260,N_9616,N_9037);
nor U10261 (N_10261,N_9988,N_9565);
or U10262 (N_10262,N_9923,N_9958);
xor U10263 (N_10263,N_9522,N_9724);
or U10264 (N_10264,N_9989,N_9309);
xnor U10265 (N_10265,N_9015,N_9066);
or U10266 (N_10266,N_9593,N_9851);
or U10267 (N_10267,N_9441,N_9542);
xor U10268 (N_10268,N_9334,N_9315);
nand U10269 (N_10269,N_9318,N_9993);
nand U10270 (N_10270,N_9843,N_9200);
xnor U10271 (N_10271,N_9214,N_9619);
xnor U10272 (N_10272,N_9461,N_9815);
nand U10273 (N_10273,N_9576,N_9790);
nor U10274 (N_10274,N_9966,N_9453);
and U10275 (N_10275,N_9868,N_9010);
and U10276 (N_10276,N_9780,N_9967);
nor U10277 (N_10277,N_9581,N_9117);
nor U10278 (N_10278,N_9573,N_9554);
nor U10279 (N_10279,N_9638,N_9959);
nor U10280 (N_10280,N_9172,N_9656);
nand U10281 (N_10281,N_9133,N_9718);
or U10282 (N_10282,N_9311,N_9333);
nand U10283 (N_10283,N_9575,N_9303);
or U10284 (N_10284,N_9012,N_9009);
and U10285 (N_10285,N_9158,N_9928);
nor U10286 (N_10286,N_9284,N_9574);
nand U10287 (N_10287,N_9919,N_9916);
nor U10288 (N_10288,N_9533,N_9776);
or U10289 (N_10289,N_9864,N_9907);
or U10290 (N_10290,N_9671,N_9615);
and U10291 (N_10291,N_9915,N_9564);
or U10292 (N_10292,N_9984,N_9218);
or U10293 (N_10293,N_9513,N_9220);
xor U10294 (N_10294,N_9427,N_9308);
xor U10295 (N_10295,N_9874,N_9637);
or U10296 (N_10296,N_9953,N_9728);
nand U10297 (N_10297,N_9350,N_9857);
or U10298 (N_10298,N_9530,N_9065);
nor U10299 (N_10299,N_9539,N_9770);
xor U10300 (N_10300,N_9088,N_9822);
xor U10301 (N_10301,N_9335,N_9077);
or U10302 (N_10302,N_9325,N_9429);
nor U10303 (N_10303,N_9030,N_9788);
xnor U10304 (N_10304,N_9025,N_9722);
nor U10305 (N_10305,N_9924,N_9816);
xor U10306 (N_10306,N_9499,N_9644);
xnor U10307 (N_10307,N_9482,N_9001);
nor U10308 (N_10308,N_9585,N_9404);
or U10309 (N_10309,N_9548,N_9440);
xnor U10310 (N_10310,N_9306,N_9794);
nand U10311 (N_10311,N_9863,N_9613);
nor U10312 (N_10312,N_9568,N_9535);
and U10313 (N_10313,N_9839,N_9592);
nand U10314 (N_10314,N_9544,N_9882);
xor U10315 (N_10315,N_9069,N_9296);
and U10316 (N_10316,N_9380,N_9290);
nand U10317 (N_10317,N_9014,N_9442);
and U10318 (N_10318,N_9013,N_9070);
and U10319 (N_10319,N_9135,N_9188);
and U10320 (N_10320,N_9838,N_9419);
nor U10321 (N_10321,N_9336,N_9704);
and U10322 (N_10322,N_9932,N_9246);
nor U10323 (N_10323,N_9068,N_9131);
or U10324 (N_10324,N_9601,N_9502);
nand U10325 (N_10325,N_9473,N_9125);
nand U10326 (N_10326,N_9326,N_9746);
or U10327 (N_10327,N_9869,N_9421);
and U10328 (N_10328,N_9250,N_9211);
and U10329 (N_10329,N_9331,N_9477);
and U10330 (N_10330,N_9349,N_9016);
or U10331 (N_10331,N_9750,N_9586);
and U10332 (N_10332,N_9970,N_9510);
and U10333 (N_10333,N_9911,N_9087);
and U10334 (N_10334,N_9620,N_9402);
or U10335 (N_10335,N_9899,N_9506);
nand U10336 (N_10336,N_9392,N_9480);
nor U10337 (N_10337,N_9500,N_9595);
nand U10338 (N_10338,N_9231,N_9733);
nor U10339 (N_10339,N_9192,N_9894);
nand U10340 (N_10340,N_9021,N_9293);
nand U10341 (N_10341,N_9189,N_9397);
xor U10342 (N_10342,N_9603,N_9063);
or U10343 (N_10343,N_9985,N_9244);
xnor U10344 (N_10344,N_9208,N_9690);
and U10345 (N_10345,N_9598,N_9681);
nand U10346 (N_10346,N_9227,N_9196);
or U10347 (N_10347,N_9948,N_9365);
xor U10348 (N_10348,N_9183,N_9623);
and U10349 (N_10349,N_9814,N_9083);
and U10350 (N_10350,N_9436,N_9545);
or U10351 (N_10351,N_9387,N_9018);
nand U10352 (N_10352,N_9610,N_9100);
nor U10353 (N_10353,N_9523,N_9312);
or U10354 (N_10354,N_9219,N_9596);
nand U10355 (N_10355,N_9340,N_9177);
nand U10356 (N_10356,N_9643,N_9398);
nand U10357 (N_10357,N_9425,N_9531);
nor U10358 (N_10358,N_9641,N_9665);
nand U10359 (N_10359,N_9235,N_9467);
nor U10360 (N_10360,N_9449,N_9840);
or U10361 (N_10361,N_9299,N_9496);
nor U10362 (N_10362,N_9632,N_9043);
xnor U10363 (N_10363,N_9768,N_9537);
xnor U10364 (N_10364,N_9624,N_9692);
nand U10365 (N_10365,N_9904,N_9463);
or U10366 (N_10366,N_9141,N_9590);
and U10367 (N_10367,N_9532,N_9849);
xor U10368 (N_10368,N_9237,N_9057);
xnor U10369 (N_10369,N_9064,N_9826);
nor U10370 (N_10370,N_9120,N_9553);
or U10371 (N_10371,N_9431,N_9124);
nor U10372 (N_10372,N_9371,N_9810);
xnor U10373 (N_10373,N_9372,N_9430);
xor U10374 (N_10374,N_9922,N_9865);
or U10375 (N_10375,N_9257,N_9341);
or U10376 (N_10376,N_9735,N_9202);
xor U10377 (N_10377,N_9968,N_9210);
xnor U10378 (N_10378,N_9081,N_9053);
nor U10379 (N_10379,N_9307,N_9550);
nor U10380 (N_10380,N_9578,N_9090);
nand U10381 (N_10381,N_9702,N_9732);
or U10382 (N_10382,N_9310,N_9700);
or U10383 (N_10383,N_9982,N_9251);
nand U10384 (N_10384,N_9204,N_9092);
and U10385 (N_10385,N_9324,N_9805);
nand U10386 (N_10386,N_9526,N_9584);
or U10387 (N_10387,N_9908,N_9465);
nor U10388 (N_10388,N_9558,N_9048);
and U10389 (N_10389,N_9130,N_9833);
xnor U10390 (N_10390,N_9751,N_9367);
nand U10391 (N_10391,N_9736,N_9490);
nor U10392 (N_10392,N_9517,N_9489);
nor U10393 (N_10393,N_9409,N_9940);
nand U10394 (N_10394,N_9521,N_9800);
or U10395 (N_10395,N_9339,N_9755);
nand U10396 (N_10396,N_9848,N_9913);
and U10397 (N_10397,N_9738,N_9852);
nor U10398 (N_10398,N_9224,N_9239);
and U10399 (N_10399,N_9494,N_9611);
xnor U10400 (N_10400,N_9662,N_9809);
xor U10401 (N_10401,N_9782,N_9529);
nand U10402 (N_10402,N_9078,N_9418);
and U10403 (N_10403,N_9027,N_9789);
nor U10404 (N_10404,N_9062,N_9354);
or U10405 (N_10405,N_9683,N_9824);
nor U10406 (N_10406,N_9741,N_9715);
nand U10407 (N_10407,N_9653,N_9627);
or U10408 (N_10408,N_9026,N_9753);
nor U10409 (N_10409,N_9524,N_9413);
nand U10410 (N_10410,N_9721,N_9602);
nor U10411 (N_10411,N_9974,N_9716);
nand U10412 (N_10412,N_9253,N_9786);
and U10413 (N_10413,N_9763,N_9695);
nand U10414 (N_10414,N_9033,N_9775);
and U10415 (N_10415,N_9567,N_9047);
xnor U10416 (N_10416,N_9507,N_9897);
nor U10417 (N_10417,N_9199,N_9356);
xor U10418 (N_10418,N_9121,N_9687);
and U10419 (N_10419,N_9217,N_9996);
or U10420 (N_10420,N_9411,N_9617);
nor U10421 (N_10421,N_9094,N_9758);
and U10422 (N_10422,N_9186,N_9626);
nor U10423 (N_10423,N_9872,N_9459);
nand U10424 (N_10424,N_9245,N_9193);
and U10425 (N_10425,N_9862,N_9708);
and U10426 (N_10426,N_9804,N_9056);
and U10427 (N_10427,N_9478,N_9707);
and U10428 (N_10428,N_9501,N_9032);
nor U10429 (N_10429,N_9799,N_9706);
nor U10430 (N_10430,N_9089,N_9487);
or U10431 (N_10431,N_9867,N_9844);
nand U10432 (N_10432,N_9388,N_9408);
nor U10433 (N_10433,N_9444,N_9020);
nand U10434 (N_10434,N_9481,N_9337);
nor U10435 (N_10435,N_9935,N_9029);
xor U10436 (N_10436,N_9268,N_9157);
nor U10437 (N_10437,N_9828,N_9228);
nand U10438 (N_10438,N_9222,N_9080);
and U10439 (N_10439,N_9964,N_9342);
nor U10440 (N_10440,N_9439,N_9143);
or U10441 (N_10441,N_9663,N_9247);
nand U10442 (N_10442,N_9345,N_9512);
nand U10443 (N_10443,N_9725,N_9961);
xor U10444 (N_10444,N_9073,N_9527);
or U10445 (N_10445,N_9000,N_9110);
nor U10446 (N_10446,N_9460,N_9176);
or U10447 (N_10447,N_9181,N_9085);
nor U10448 (N_10448,N_9098,N_9305);
nand U10449 (N_10449,N_9184,N_9095);
or U10450 (N_10450,N_9447,N_9243);
and U10451 (N_10451,N_9747,N_9742);
nand U10452 (N_10452,N_9286,N_9022);
xnor U10453 (N_10453,N_9498,N_9890);
nor U10454 (N_10454,N_9798,N_9007);
or U10455 (N_10455,N_9877,N_9209);
and U10456 (N_10456,N_9795,N_9138);
nor U10457 (N_10457,N_9097,N_9847);
nand U10458 (N_10458,N_9152,N_9936);
or U10459 (N_10459,N_9920,N_9093);
nor U10460 (N_10460,N_9859,N_9727);
xor U10461 (N_10461,N_9536,N_9075);
or U10462 (N_10462,N_9504,N_9259);
and U10463 (N_10463,N_9491,N_9949);
xnor U10464 (N_10464,N_9024,N_9556);
nor U10465 (N_10465,N_9635,N_9679);
nor U10466 (N_10466,N_9739,N_9273);
xor U10467 (N_10467,N_9830,N_9059);
or U10468 (N_10468,N_9675,N_9252);
nor U10469 (N_10469,N_9396,N_9178);
and U10470 (N_10470,N_9383,N_9119);
nand U10471 (N_10471,N_9688,N_9366);
nor U10472 (N_10472,N_9630,N_9673);
nor U10473 (N_10473,N_9842,N_9361);
nand U10474 (N_10474,N_9067,N_9300);
xnor U10475 (N_10475,N_9705,N_9701);
nand U10476 (N_10476,N_9797,N_9451);
xor U10477 (N_10477,N_9921,N_9827);
or U10478 (N_10478,N_9555,N_9992);
nor U10479 (N_10479,N_9285,N_9103);
nand U10480 (N_10480,N_9107,N_9084);
and U10481 (N_10481,N_9986,N_9893);
and U10482 (N_10482,N_9410,N_9861);
nor U10483 (N_10483,N_9362,N_9044);
nand U10484 (N_10484,N_9972,N_9505);
or U10485 (N_10485,N_9274,N_9760);
xnor U10486 (N_10486,N_9552,N_9870);
xor U10487 (N_10487,N_9672,N_9216);
xnor U10488 (N_10488,N_9479,N_9661);
nor U10489 (N_10489,N_9347,N_9379);
xor U10490 (N_10490,N_9426,N_9762);
nor U10491 (N_10491,N_9779,N_9802);
or U10492 (N_10492,N_9455,N_9825);
nand U10493 (N_10493,N_9432,N_9850);
and U10494 (N_10494,N_9730,N_9201);
nor U10495 (N_10495,N_9639,N_9667);
nand U10496 (N_10496,N_9880,N_9900);
and U10497 (N_10497,N_9028,N_9006);
and U10498 (N_10498,N_9946,N_9678);
nor U10499 (N_10499,N_9375,N_9074);
or U10500 (N_10500,N_9832,N_9545);
or U10501 (N_10501,N_9880,N_9110);
and U10502 (N_10502,N_9397,N_9399);
or U10503 (N_10503,N_9540,N_9703);
nand U10504 (N_10504,N_9533,N_9027);
and U10505 (N_10505,N_9023,N_9015);
xor U10506 (N_10506,N_9926,N_9874);
nand U10507 (N_10507,N_9640,N_9254);
or U10508 (N_10508,N_9969,N_9124);
and U10509 (N_10509,N_9192,N_9546);
nor U10510 (N_10510,N_9944,N_9674);
nand U10511 (N_10511,N_9144,N_9960);
nand U10512 (N_10512,N_9297,N_9655);
nand U10513 (N_10513,N_9865,N_9913);
and U10514 (N_10514,N_9996,N_9136);
nor U10515 (N_10515,N_9391,N_9624);
and U10516 (N_10516,N_9275,N_9560);
nand U10517 (N_10517,N_9555,N_9646);
or U10518 (N_10518,N_9308,N_9084);
nor U10519 (N_10519,N_9009,N_9899);
nand U10520 (N_10520,N_9938,N_9086);
and U10521 (N_10521,N_9854,N_9228);
xnor U10522 (N_10522,N_9983,N_9004);
or U10523 (N_10523,N_9999,N_9671);
nand U10524 (N_10524,N_9894,N_9431);
and U10525 (N_10525,N_9576,N_9809);
nor U10526 (N_10526,N_9527,N_9509);
or U10527 (N_10527,N_9746,N_9361);
nor U10528 (N_10528,N_9124,N_9003);
nor U10529 (N_10529,N_9763,N_9717);
xnor U10530 (N_10530,N_9938,N_9562);
xnor U10531 (N_10531,N_9066,N_9248);
nor U10532 (N_10532,N_9208,N_9592);
nor U10533 (N_10533,N_9145,N_9909);
nor U10534 (N_10534,N_9229,N_9774);
xnor U10535 (N_10535,N_9395,N_9929);
and U10536 (N_10536,N_9507,N_9111);
xnor U10537 (N_10537,N_9579,N_9856);
nor U10538 (N_10538,N_9198,N_9639);
or U10539 (N_10539,N_9360,N_9349);
xor U10540 (N_10540,N_9237,N_9337);
and U10541 (N_10541,N_9183,N_9487);
nand U10542 (N_10542,N_9119,N_9156);
nor U10543 (N_10543,N_9728,N_9963);
nor U10544 (N_10544,N_9240,N_9130);
xnor U10545 (N_10545,N_9326,N_9179);
xnor U10546 (N_10546,N_9943,N_9481);
xor U10547 (N_10547,N_9532,N_9570);
nand U10548 (N_10548,N_9784,N_9633);
nand U10549 (N_10549,N_9063,N_9928);
and U10550 (N_10550,N_9203,N_9999);
or U10551 (N_10551,N_9990,N_9982);
and U10552 (N_10552,N_9934,N_9002);
or U10553 (N_10553,N_9442,N_9369);
and U10554 (N_10554,N_9154,N_9749);
nor U10555 (N_10555,N_9041,N_9816);
xor U10556 (N_10556,N_9589,N_9107);
nand U10557 (N_10557,N_9964,N_9330);
nor U10558 (N_10558,N_9752,N_9980);
xnor U10559 (N_10559,N_9112,N_9405);
and U10560 (N_10560,N_9824,N_9177);
nor U10561 (N_10561,N_9114,N_9866);
nor U10562 (N_10562,N_9587,N_9915);
nor U10563 (N_10563,N_9466,N_9550);
and U10564 (N_10564,N_9469,N_9253);
xnor U10565 (N_10565,N_9618,N_9204);
or U10566 (N_10566,N_9045,N_9028);
xnor U10567 (N_10567,N_9571,N_9075);
or U10568 (N_10568,N_9504,N_9568);
and U10569 (N_10569,N_9737,N_9210);
nor U10570 (N_10570,N_9437,N_9704);
nand U10571 (N_10571,N_9627,N_9724);
or U10572 (N_10572,N_9079,N_9549);
nand U10573 (N_10573,N_9656,N_9600);
and U10574 (N_10574,N_9320,N_9321);
and U10575 (N_10575,N_9464,N_9795);
nand U10576 (N_10576,N_9795,N_9829);
nand U10577 (N_10577,N_9717,N_9256);
nor U10578 (N_10578,N_9589,N_9847);
and U10579 (N_10579,N_9288,N_9354);
xor U10580 (N_10580,N_9400,N_9331);
nor U10581 (N_10581,N_9139,N_9906);
nor U10582 (N_10582,N_9390,N_9299);
and U10583 (N_10583,N_9309,N_9842);
nand U10584 (N_10584,N_9975,N_9597);
nand U10585 (N_10585,N_9097,N_9457);
nor U10586 (N_10586,N_9069,N_9174);
or U10587 (N_10587,N_9501,N_9260);
nand U10588 (N_10588,N_9048,N_9900);
or U10589 (N_10589,N_9098,N_9913);
xnor U10590 (N_10590,N_9754,N_9836);
nand U10591 (N_10591,N_9429,N_9905);
xor U10592 (N_10592,N_9022,N_9782);
and U10593 (N_10593,N_9676,N_9756);
nor U10594 (N_10594,N_9571,N_9682);
or U10595 (N_10595,N_9979,N_9646);
nor U10596 (N_10596,N_9477,N_9628);
and U10597 (N_10597,N_9460,N_9026);
or U10598 (N_10598,N_9400,N_9724);
xnor U10599 (N_10599,N_9579,N_9930);
or U10600 (N_10600,N_9803,N_9983);
xor U10601 (N_10601,N_9469,N_9996);
or U10602 (N_10602,N_9822,N_9559);
and U10603 (N_10603,N_9816,N_9013);
xnor U10604 (N_10604,N_9535,N_9502);
xnor U10605 (N_10605,N_9821,N_9738);
xnor U10606 (N_10606,N_9369,N_9020);
or U10607 (N_10607,N_9536,N_9024);
nor U10608 (N_10608,N_9807,N_9207);
and U10609 (N_10609,N_9814,N_9878);
xnor U10610 (N_10610,N_9447,N_9008);
xor U10611 (N_10611,N_9447,N_9302);
xnor U10612 (N_10612,N_9535,N_9348);
or U10613 (N_10613,N_9215,N_9634);
xnor U10614 (N_10614,N_9873,N_9581);
nand U10615 (N_10615,N_9908,N_9357);
nand U10616 (N_10616,N_9298,N_9927);
and U10617 (N_10617,N_9725,N_9822);
or U10618 (N_10618,N_9242,N_9867);
xor U10619 (N_10619,N_9701,N_9459);
nand U10620 (N_10620,N_9646,N_9942);
nor U10621 (N_10621,N_9144,N_9028);
xnor U10622 (N_10622,N_9081,N_9899);
nand U10623 (N_10623,N_9573,N_9021);
xor U10624 (N_10624,N_9951,N_9326);
and U10625 (N_10625,N_9674,N_9788);
or U10626 (N_10626,N_9379,N_9109);
nor U10627 (N_10627,N_9784,N_9630);
xor U10628 (N_10628,N_9010,N_9184);
nand U10629 (N_10629,N_9801,N_9443);
or U10630 (N_10630,N_9231,N_9104);
or U10631 (N_10631,N_9676,N_9975);
xor U10632 (N_10632,N_9497,N_9155);
and U10633 (N_10633,N_9451,N_9344);
or U10634 (N_10634,N_9734,N_9344);
nand U10635 (N_10635,N_9448,N_9395);
nor U10636 (N_10636,N_9378,N_9268);
and U10637 (N_10637,N_9727,N_9175);
xnor U10638 (N_10638,N_9595,N_9215);
and U10639 (N_10639,N_9549,N_9869);
or U10640 (N_10640,N_9449,N_9916);
nor U10641 (N_10641,N_9200,N_9422);
nand U10642 (N_10642,N_9893,N_9099);
nor U10643 (N_10643,N_9200,N_9829);
or U10644 (N_10644,N_9140,N_9527);
nand U10645 (N_10645,N_9485,N_9973);
nand U10646 (N_10646,N_9804,N_9081);
nor U10647 (N_10647,N_9019,N_9229);
nand U10648 (N_10648,N_9025,N_9288);
xnor U10649 (N_10649,N_9156,N_9613);
xnor U10650 (N_10650,N_9592,N_9845);
xor U10651 (N_10651,N_9441,N_9167);
or U10652 (N_10652,N_9407,N_9928);
nand U10653 (N_10653,N_9875,N_9267);
nand U10654 (N_10654,N_9058,N_9365);
xnor U10655 (N_10655,N_9176,N_9834);
xnor U10656 (N_10656,N_9463,N_9079);
nand U10657 (N_10657,N_9725,N_9373);
nand U10658 (N_10658,N_9978,N_9078);
and U10659 (N_10659,N_9815,N_9571);
or U10660 (N_10660,N_9662,N_9195);
xor U10661 (N_10661,N_9453,N_9390);
nor U10662 (N_10662,N_9161,N_9950);
or U10663 (N_10663,N_9885,N_9516);
and U10664 (N_10664,N_9088,N_9599);
nor U10665 (N_10665,N_9881,N_9087);
or U10666 (N_10666,N_9573,N_9132);
and U10667 (N_10667,N_9298,N_9011);
and U10668 (N_10668,N_9879,N_9535);
nor U10669 (N_10669,N_9124,N_9049);
nor U10670 (N_10670,N_9028,N_9277);
xnor U10671 (N_10671,N_9721,N_9909);
or U10672 (N_10672,N_9719,N_9613);
nor U10673 (N_10673,N_9202,N_9104);
or U10674 (N_10674,N_9089,N_9825);
and U10675 (N_10675,N_9603,N_9522);
xnor U10676 (N_10676,N_9101,N_9863);
nor U10677 (N_10677,N_9018,N_9492);
and U10678 (N_10678,N_9622,N_9462);
nand U10679 (N_10679,N_9114,N_9241);
or U10680 (N_10680,N_9154,N_9477);
or U10681 (N_10681,N_9304,N_9106);
or U10682 (N_10682,N_9728,N_9814);
nor U10683 (N_10683,N_9351,N_9005);
xnor U10684 (N_10684,N_9212,N_9765);
nand U10685 (N_10685,N_9827,N_9333);
or U10686 (N_10686,N_9720,N_9747);
and U10687 (N_10687,N_9345,N_9858);
nor U10688 (N_10688,N_9561,N_9942);
and U10689 (N_10689,N_9454,N_9841);
xnor U10690 (N_10690,N_9284,N_9214);
or U10691 (N_10691,N_9544,N_9586);
and U10692 (N_10692,N_9672,N_9995);
and U10693 (N_10693,N_9096,N_9638);
or U10694 (N_10694,N_9977,N_9832);
nand U10695 (N_10695,N_9910,N_9009);
xor U10696 (N_10696,N_9694,N_9482);
or U10697 (N_10697,N_9763,N_9314);
xnor U10698 (N_10698,N_9811,N_9901);
and U10699 (N_10699,N_9990,N_9143);
nand U10700 (N_10700,N_9331,N_9498);
nor U10701 (N_10701,N_9291,N_9728);
nand U10702 (N_10702,N_9715,N_9284);
nand U10703 (N_10703,N_9536,N_9246);
nor U10704 (N_10704,N_9458,N_9917);
or U10705 (N_10705,N_9876,N_9174);
nand U10706 (N_10706,N_9910,N_9862);
nor U10707 (N_10707,N_9067,N_9623);
or U10708 (N_10708,N_9708,N_9616);
or U10709 (N_10709,N_9088,N_9470);
and U10710 (N_10710,N_9602,N_9807);
nor U10711 (N_10711,N_9081,N_9207);
nand U10712 (N_10712,N_9446,N_9577);
nand U10713 (N_10713,N_9771,N_9157);
and U10714 (N_10714,N_9170,N_9520);
nor U10715 (N_10715,N_9432,N_9830);
and U10716 (N_10716,N_9590,N_9610);
or U10717 (N_10717,N_9127,N_9440);
xnor U10718 (N_10718,N_9515,N_9554);
nand U10719 (N_10719,N_9484,N_9170);
or U10720 (N_10720,N_9703,N_9386);
or U10721 (N_10721,N_9186,N_9505);
xnor U10722 (N_10722,N_9565,N_9451);
or U10723 (N_10723,N_9224,N_9256);
or U10724 (N_10724,N_9806,N_9101);
nor U10725 (N_10725,N_9661,N_9378);
and U10726 (N_10726,N_9689,N_9063);
or U10727 (N_10727,N_9886,N_9131);
nor U10728 (N_10728,N_9428,N_9012);
xor U10729 (N_10729,N_9802,N_9730);
xor U10730 (N_10730,N_9940,N_9454);
or U10731 (N_10731,N_9211,N_9780);
and U10732 (N_10732,N_9828,N_9773);
and U10733 (N_10733,N_9918,N_9706);
and U10734 (N_10734,N_9630,N_9383);
nand U10735 (N_10735,N_9109,N_9454);
or U10736 (N_10736,N_9444,N_9281);
or U10737 (N_10737,N_9013,N_9927);
nor U10738 (N_10738,N_9772,N_9032);
xor U10739 (N_10739,N_9074,N_9303);
nand U10740 (N_10740,N_9235,N_9179);
xnor U10741 (N_10741,N_9189,N_9911);
and U10742 (N_10742,N_9433,N_9540);
nor U10743 (N_10743,N_9197,N_9993);
nand U10744 (N_10744,N_9268,N_9049);
xor U10745 (N_10745,N_9411,N_9915);
and U10746 (N_10746,N_9245,N_9274);
and U10747 (N_10747,N_9075,N_9421);
xnor U10748 (N_10748,N_9231,N_9517);
and U10749 (N_10749,N_9412,N_9950);
nor U10750 (N_10750,N_9658,N_9216);
and U10751 (N_10751,N_9489,N_9032);
or U10752 (N_10752,N_9678,N_9874);
nand U10753 (N_10753,N_9317,N_9319);
nand U10754 (N_10754,N_9178,N_9383);
nor U10755 (N_10755,N_9343,N_9072);
nand U10756 (N_10756,N_9240,N_9633);
or U10757 (N_10757,N_9226,N_9178);
nor U10758 (N_10758,N_9269,N_9744);
xnor U10759 (N_10759,N_9916,N_9525);
and U10760 (N_10760,N_9247,N_9408);
nand U10761 (N_10761,N_9806,N_9430);
or U10762 (N_10762,N_9381,N_9789);
xor U10763 (N_10763,N_9895,N_9490);
nand U10764 (N_10764,N_9112,N_9808);
nand U10765 (N_10765,N_9051,N_9408);
and U10766 (N_10766,N_9721,N_9293);
nor U10767 (N_10767,N_9025,N_9342);
nand U10768 (N_10768,N_9266,N_9201);
nand U10769 (N_10769,N_9711,N_9894);
nor U10770 (N_10770,N_9375,N_9854);
or U10771 (N_10771,N_9130,N_9371);
xnor U10772 (N_10772,N_9549,N_9119);
and U10773 (N_10773,N_9273,N_9132);
nand U10774 (N_10774,N_9128,N_9656);
and U10775 (N_10775,N_9016,N_9303);
xor U10776 (N_10776,N_9890,N_9174);
or U10777 (N_10777,N_9522,N_9358);
and U10778 (N_10778,N_9534,N_9985);
xor U10779 (N_10779,N_9522,N_9444);
nand U10780 (N_10780,N_9176,N_9264);
or U10781 (N_10781,N_9792,N_9605);
xnor U10782 (N_10782,N_9550,N_9749);
nand U10783 (N_10783,N_9952,N_9441);
nand U10784 (N_10784,N_9862,N_9153);
or U10785 (N_10785,N_9956,N_9015);
or U10786 (N_10786,N_9890,N_9685);
nand U10787 (N_10787,N_9106,N_9479);
nor U10788 (N_10788,N_9953,N_9497);
nand U10789 (N_10789,N_9109,N_9460);
and U10790 (N_10790,N_9095,N_9065);
nor U10791 (N_10791,N_9596,N_9177);
and U10792 (N_10792,N_9486,N_9324);
and U10793 (N_10793,N_9365,N_9817);
or U10794 (N_10794,N_9510,N_9119);
nor U10795 (N_10795,N_9320,N_9078);
xor U10796 (N_10796,N_9770,N_9959);
nand U10797 (N_10797,N_9889,N_9017);
xor U10798 (N_10798,N_9745,N_9054);
nand U10799 (N_10799,N_9709,N_9300);
nor U10800 (N_10800,N_9029,N_9998);
nor U10801 (N_10801,N_9739,N_9618);
nor U10802 (N_10802,N_9542,N_9475);
xor U10803 (N_10803,N_9208,N_9377);
nand U10804 (N_10804,N_9369,N_9365);
or U10805 (N_10805,N_9274,N_9921);
xnor U10806 (N_10806,N_9164,N_9099);
or U10807 (N_10807,N_9879,N_9899);
nand U10808 (N_10808,N_9149,N_9108);
nand U10809 (N_10809,N_9531,N_9022);
nor U10810 (N_10810,N_9263,N_9699);
nor U10811 (N_10811,N_9810,N_9577);
nor U10812 (N_10812,N_9991,N_9261);
nand U10813 (N_10813,N_9326,N_9776);
or U10814 (N_10814,N_9505,N_9841);
nand U10815 (N_10815,N_9586,N_9588);
nand U10816 (N_10816,N_9962,N_9323);
xnor U10817 (N_10817,N_9089,N_9095);
nand U10818 (N_10818,N_9927,N_9879);
nand U10819 (N_10819,N_9589,N_9184);
xnor U10820 (N_10820,N_9792,N_9878);
xor U10821 (N_10821,N_9068,N_9716);
xnor U10822 (N_10822,N_9122,N_9672);
and U10823 (N_10823,N_9567,N_9093);
or U10824 (N_10824,N_9728,N_9245);
and U10825 (N_10825,N_9938,N_9638);
and U10826 (N_10826,N_9989,N_9176);
nand U10827 (N_10827,N_9049,N_9626);
xor U10828 (N_10828,N_9903,N_9249);
or U10829 (N_10829,N_9855,N_9925);
and U10830 (N_10830,N_9128,N_9637);
xor U10831 (N_10831,N_9481,N_9389);
and U10832 (N_10832,N_9551,N_9182);
and U10833 (N_10833,N_9760,N_9523);
nor U10834 (N_10834,N_9712,N_9488);
nand U10835 (N_10835,N_9219,N_9971);
xor U10836 (N_10836,N_9705,N_9564);
or U10837 (N_10837,N_9990,N_9512);
xor U10838 (N_10838,N_9735,N_9685);
nand U10839 (N_10839,N_9625,N_9156);
nand U10840 (N_10840,N_9945,N_9573);
nor U10841 (N_10841,N_9105,N_9816);
xnor U10842 (N_10842,N_9243,N_9803);
nor U10843 (N_10843,N_9831,N_9289);
or U10844 (N_10844,N_9299,N_9900);
nand U10845 (N_10845,N_9481,N_9367);
nor U10846 (N_10846,N_9231,N_9497);
and U10847 (N_10847,N_9863,N_9573);
xnor U10848 (N_10848,N_9877,N_9534);
or U10849 (N_10849,N_9465,N_9540);
nand U10850 (N_10850,N_9398,N_9602);
and U10851 (N_10851,N_9569,N_9493);
and U10852 (N_10852,N_9302,N_9003);
xor U10853 (N_10853,N_9654,N_9027);
and U10854 (N_10854,N_9712,N_9031);
or U10855 (N_10855,N_9188,N_9615);
nor U10856 (N_10856,N_9795,N_9583);
and U10857 (N_10857,N_9497,N_9954);
nand U10858 (N_10858,N_9673,N_9603);
nor U10859 (N_10859,N_9344,N_9126);
nor U10860 (N_10860,N_9393,N_9601);
and U10861 (N_10861,N_9051,N_9131);
or U10862 (N_10862,N_9387,N_9416);
xnor U10863 (N_10863,N_9070,N_9006);
nand U10864 (N_10864,N_9019,N_9798);
xnor U10865 (N_10865,N_9906,N_9735);
nor U10866 (N_10866,N_9317,N_9274);
xnor U10867 (N_10867,N_9687,N_9619);
nand U10868 (N_10868,N_9869,N_9457);
and U10869 (N_10869,N_9506,N_9684);
and U10870 (N_10870,N_9298,N_9649);
xor U10871 (N_10871,N_9219,N_9080);
or U10872 (N_10872,N_9153,N_9311);
or U10873 (N_10873,N_9337,N_9702);
xor U10874 (N_10874,N_9489,N_9594);
nor U10875 (N_10875,N_9721,N_9396);
xnor U10876 (N_10876,N_9881,N_9136);
nor U10877 (N_10877,N_9011,N_9426);
nand U10878 (N_10878,N_9453,N_9571);
nand U10879 (N_10879,N_9715,N_9744);
nand U10880 (N_10880,N_9649,N_9055);
nor U10881 (N_10881,N_9552,N_9616);
or U10882 (N_10882,N_9036,N_9037);
nand U10883 (N_10883,N_9382,N_9739);
xnor U10884 (N_10884,N_9164,N_9690);
and U10885 (N_10885,N_9829,N_9455);
or U10886 (N_10886,N_9097,N_9057);
or U10887 (N_10887,N_9925,N_9429);
and U10888 (N_10888,N_9382,N_9858);
and U10889 (N_10889,N_9280,N_9272);
or U10890 (N_10890,N_9490,N_9574);
or U10891 (N_10891,N_9437,N_9903);
and U10892 (N_10892,N_9797,N_9475);
or U10893 (N_10893,N_9471,N_9409);
nand U10894 (N_10894,N_9407,N_9639);
xor U10895 (N_10895,N_9514,N_9862);
or U10896 (N_10896,N_9364,N_9216);
and U10897 (N_10897,N_9483,N_9395);
xnor U10898 (N_10898,N_9582,N_9023);
nand U10899 (N_10899,N_9225,N_9881);
nand U10900 (N_10900,N_9359,N_9062);
xnor U10901 (N_10901,N_9974,N_9769);
nand U10902 (N_10902,N_9269,N_9997);
nor U10903 (N_10903,N_9317,N_9080);
nand U10904 (N_10904,N_9231,N_9537);
nor U10905 (N_10905,N_9720,N_9567);
or U10906 (N_10906,N_9325,N_9511);
nor U10907 (N_10907,N_9912,N_9594);
xor U10908 (N_10908,N_9024,N_9181);
nand U10909 (N_10909,N_9022,N_9822);
nor U10910 (N_10910,N_9484,N_9860);
nor U10911 (N_10911,N_9631,N_9173);
nand U10912 (N_10912,N_9917,N_9289);
nand U10913 (N_10913,N_9571,N_9631);
nor U10914 (N_10914,N_9072,N_9470);
nand U10915 (N_10915,N_9726,N_9639);
and U10916 (N_10916,N_9788,N_9866);
xor U10917 (N_10917,N_9617,N_9941);
nand U10918 (N_10918,N_9405,N_9745);
xor U10919 (N_10919,N_9088,N_9909);
or U10920 (N_10920,N_9260,N_9259);
or U10921 (N_10921,N_9988,N_9197);
and U10922 (N_10922,N_9422,N_9919);
and U10923 (N_10923,N_9764,N_9734);
or U10924 (N_10924,N_9882,N_9409);
and U10925 (N_10925,N_9892,N_9061);
or U10926 (N_10926,N_9702,N_9954);
and U10927 (N_10927,N_9066,N_9582);
xnor U10928 (N_10928,N_9250,N_9013);
or U10929 (N_10929,N_9883,N_9193);
nand U10930 (N_10930,N_9922,N_9061);
nand U10931 (N_10931,N_9756,N_9960);
and U10932 (N_10932,N_9110,N_9702);
or U10933 (N_10933,N_9536,N_9677);
nor U10934 (N_10934,N_9686,N_9407);
and U10935 (N_10935,N_9555,N_9816);
and U10936 (N_10936,N_9103,N_9316);
or U10937 (N_10937,N_9305,N_9803);
nand U10938 (N_10938,N_9138,N_9013);
and U10939 (N_10939,N_9389,N_9900);
xor U10940 (N_10940,N_9303,N_9268);
nand U10941 (N_10941,N_9765,N_9968);
and U10942 (N_10942,N_9554,N_9172);
nand U10943 (N_10943,N_9679,N_9222);
nand U10944 (N_10944,N_9929,N_9818);
xor U10945 (N_10945,N_9149,N_9720);
xnor U10946 (N_10946,N_9010,N_9325);
xor U10947 (N_10947,N_9313,N_9330);
nor U10948 (N_10948,N_9877,N_9533);
and U10949 (N_10949,N_9657,N_9465);
nand U10950 (N_10950,N_9144,N_9957);
or U10951 (N_10951,N_9670,N_9825);
or U10952 (N_10952,N_9030,N_9403);
and U10953 (N_10953,N_9647,N_9134);
nand U10954 (N_10954,N_9688,N_9829);
and U10955 (N_10955,N_9192,N_9828);
nor U10956 (N_10956,N_9990,N_9069);
nor U10957 (N_10957,N_9461,N_9639);
xnor U10958 (N_10958,N_9057,N_9968);
xor U10959 (N_10959,N_9330,N_9974);
or U10960 (N_10960,N_9174,N_9948);
xnor U10961 (N_10961,N_9321,N_9842);
xnor U10962 (N_10962,N_9215,N_9945);
and U10963 (N_10963,N_9527,N_9810);
or U10964 (N_10964,N_9224,N_9007);
and U10965 (N_10965,N_9466,N_9591);
nor U10966 (N_10966,N_9695,N_9026);
xor U10967 (N_10967,N_9196,N_9747);
and U10968 (N_10968,N_9854,N_9223);
nor U10969 (N_10969,N_9859,N_9252);
nor U10970 (N_10970,N_9213,N_9269);
and U10971 (N_10971,N_9979,N_9021);
or U10972 (N_10972,N_9063,N_9115);
and U10973 (N_10973,N_9002,N_9745);
or U10974 (N_10974,N_9828,N_9247);
nor U10975 (N_10975,N_9210,N_9627);
nand U10976 (N_10976,N_9756,N_9324);
nand U10977 (N_10977,N_9635,N_9659);
nor U10978 (N_10978,N_9373,N_9346);
and U10979 (N_10979,N_9735,N_9336);
nand U10980 (N_10980,N_9002,N_9257);
and U10981 (N_10981,N_9830,N_9472);
or U10982 (N_10982,N_9236,N_9724);
nand U10983 (N_10983,N_9051,N_9537);
nor U10984 (N_10984,N_9516,N_9268);
or U10985 (N_10985,N_9396,N_9193);
and U10986 (N_10986,N_9862,N_9138);
or U10987 (N_10987,N_9130,N_9615);
or U10988 (N_10988,N_9079,N_9778);
or U10989 (N_10989,N_9856,N_9674);
xor U10990 (N_10990,N_9474,N_9006);
nand U10991 (N_10991,N_9945,N_9801);
nor U10992 (N_10992,N_9498,N_9366);
nor U10993 (N_10993,N_9967,N_9892);
or U10994 (N_10994,N_9686,N_9865);
nor U10995 (N_10995,N_9060,N_9218);
and U10996 (N_10996,N_9876,N_9153);
or U10997 (N_10997,N_9115,N_9488);
and U10998 (N_10998,N_9513,N_9222);
xor U10999 (N_10999,N_9723,N_9824);
nor U11000 (N_11000,N_10614,N_10995);
nor U11001 (N_11001,N_10713,N_10832);
or U11002 (N_11002,N_10356,N_10010);
or U11003 (N_11003,N_10666,N_10409);
or U11004 (N_11004,N_10205,N_10689);
xor U11005 (N_11005,N_10911,N_10078);
or U11006 (N_11006,N_10853,N_10969);
and U11007 (N_11007,N_10525,N_10470);
or U11008 (N_11008,N_10512,N_10464);
and U11009 (N_11009,N_10918,N_10753);
nor U11010 (N_11010,N_10871,N_10496);
nor U11011 (N_11011,N_10137,N_10655);
nor U11012 (N_11012,N_10772,N_10179);
nand U11013 (N_11013,N_10703,N_10377);
and U11014 (N_11014,N_10695,N_10516);
nor U11015 (N_11015,N_10349,N_10505);
or U11016 (N_11016,N_10828,N_10773);
and U11017 (N_11017,N_10293,N_10158);
and U11018 (N_11018,N_10716,N_10542);
nand U11019 (N_11019,N_10860,N_10774);
or U11020 (N_11020,N_10439,N_10107);
or U11021 (N_11021,N_10881,N_10507);
nor U11022 (N_11022,N_10261,N_10462);
xor U11023 (N_11023,N_10769,N_10906);
xor U11024 (N_11024,N_10836,N_10761);
nor U11025 (N_11025,N_10143,N_10213);
and U11026 (N_11026,N_10958,N_10531);
nand U11027 (N_11027,N_10019,N_10636);
nand U11028 (N_11028,N_10175,N_10087);
nand U11029 (N_11029,N_10754,N_10206);
and U11030 (N_11030,N_10745,N_10109);
nand U11031 (N_11031,N_10279,N_10351);
nand U11032 (N_11032,N_10931,N_10541);
and U11033 (N_11033,N_10567,N_10764);
nand U11034 (N_11034,N_10849,N_10125);
nor U11035 (N_11035,N_10028,N_10993);
xnor U11036 (N_11036,N_10629,N_10050);
nand U11037 (N_11037,N_10469,N_10942);
or U11038 (N_11038,N_10110,N_10641);
and U11039 (N_11039,N_10341,N_10168);
xnor U11040 (N_11040,N_10862,N_10480);
nor U11041 (N_11041,N_10956,N_10581);
or U11042 (N_11042,N_10685,N_10526);
nand U11043 (N_11043,N_10103,N_10159);
xnor U11044 (N_11044,N_10845,N_10659);
xor U11045 (N_11045,N_10642,N_10442);
nand U11046 (N_11046,N_10215,N_10527);
and U11047 (N_11047,N_10289,N_10556);
and U11048 (N_11048,N_10971,N_10840);
xnor U11049 (N_11049,N_10669,N_10009);
nor U11050 (N_11050,N_10933,N_10684);
nor U11051 (N_11051,N_10692,N_10352);
and U11052 (N_11052,N_10679,N_10064);
nand U11053 (N_11053,N_10976,N_10375);
nor U11054 (N_11054,N_10301,N_10374);
nor U11055 (N_11055,N_10468,N_10463);
or U11056 (N_11056,N_10667,N_10590);
nor U11057 (N_11057,N_10072,N_10891);
and U11058 (N_11058,N_10285,N_10668);
nor U11059 (N_11059,N_10079,N_10458);
xor U11060 (N_11060,N_10309,N_10705);
or U11061 (N_11061,N_10337,N_10591);
and U11062 (N_11062,N_10571,N_10012);
or U11063 (N_11063,N_10287,N_10700);
nand U11064 (N_11064,N_10876,N_10198);
and U11065 (N_11065,N_10886,N_10015);
or U11066 (N_11066,N_10691,N_10304);
xnor U11067 (N_11067,N_10018,N_10965);
and U11068 (N_11068,N_10718,N_10077);
and U11069 (N_11069,N_10503,N_10132);
xnor U11070 (N_11070,N_10837,N_10059);
xor U11071 (N_11071,N_10658,N_10214);
and U11072 (N_11072,N_10466,N_10224);
or U11073 (N_11073,N_10418,N_10791);
nor U11074 (N_11074,N_10176,N_10486);
and U11075 (N_11075,N_10093,N_10719);
nand U11076 (N_11076,N_10264,N_10178);
and U11077 (N_11077,N_10998,N_10366);
and U11078 (N_11078,N_10278,N_10405);
or U11079 (N_11079,N_10621,N_10454);
or U11080 (N_11080,N_10733,N_10857);
or U11081 (N_11081,N_10120,N_10286);
nor U11082 (N_11082,N_10736,N_10492);
nor U11083 (N_11083,N_10238,N_10795);
nor U11084 (N_11084,N_10847,N_10574);
nand U11085 (N_11085,N_10217,N_10709);
or U11086 (N_11086,N_10748,N_10811);
and U11087 (N_11087,N_10834,N_10276);
nor U11088 (N_11088,N_10649,N_10343);
nand U11089 (N_11089,N_10829,N_10057);
and U11090 (N_11090,N_10407,N_10323);
or U11091 (N_11091,N_10076,N_10555);
xor U11092 (N_11092,N_10450,N_10779);
or U11093 (N_11093,N_10485,N_10426);
nand U11094 (N_11094,N_10780,N_10623);
xnor U11095 (N_11095,N_10319,N_10167);
and U11096 (N_11096,N_10966,N_10024);
or U11097 (N_11097,N_10537,N_10031);
or U11098 (N_11098,N_10524,N_10620);
nand U11099 (N_11099,N_10706,N_10484);
nor U11100 (N_11100,N_10036,N_10661);
nor U11101 (N_11101,N_10164,N_10711);
nand U11102 (N_11102,N_10386,N_10633);
or U11103 (N_11103,N_10533,N_10271);
nand U11104 (N_11104,N_10095,N_10677);
nor U11105 (N_11105,N_10983,N_10570);
xor U11106 (N_11106,N_10927,N_10855);
nor U11107 (N_11107,N_10563,N_10550);
nor U11108 (N_11108,N_10201,N_10473);
xnor U11109 (N_11109,N_10979,N_10844);
nor U11110 (N_11110,N_10743,N_10495);
nor U11111 (N_11111,N_10548,N_10021);
or U11112 (N_11112,N_10543,N_10529);
nand U11113 (N_11113,N_10895,N_10506);
nor U11114 (N_11114,N_10456,N_10449);
and U11115 (N_11115,N_10731,N_10790);
or U11116 (N_11116,N_10850,N_10569);
and U11117 (N_11117,N_10777,N_10187);
nand U11118 (N_11118,N_10608,N_10568);
nand U11119 (N_11119,N_10562,N_10263);
nand U11120 (N_11120,N_10963,N_10062);
nor U11121 (N_11121,N_10978,N_10482);
nand U11122 (N_11122,N_10382,N_10363);
nor U11123 (N_11123,N_10693,N_10421);
or U11124 (N_11124,N_10902,N_10274);
nor U11125 (N_11125,N_10387,N_10866);
xor U11126 (N_11126,N_10166,N_10887);
nand U11127 (N_11127,N_10557,N_10964);
or U11128 (N_11128,N_10822,N_10594);
nor U11129 (N_11129,N_10115,N_10868);
and U11130 (N_11130,N_10023,N_10919);
xor U11131 (N_11131,N_10243,N_10910);
xor U11132 (N_11132,N_10502,N_10626);
nand U11133 (N_11133,N_10814,N_10508);
nand U11134 (N_11134,N_10219,N_10465);
nand U11135 (N_11135,N_10129,N_10535);
nand U11136 (N_11136,N_10598,N_10712);
nand U11137 (N_11137,N_10913,N_10231);
nor U11138 (N_11138,N_10500,N_10230);
xnor U11139 (N_11139,N_10003,N_10900);
nand U11140 (N_11140,N_10235,N_10767);
and U11141 (N_11141,N_10404,N_10270);
and U11142 (N_11142,N_10317,N_10262);
nor U11143 (N_11143,N_10987,N_10930);
and U11144 (N_11144,N_10967,N_10281);
xnor U11145 (N_11145,N_10472,N_10924);
nor U11146 (N_11146,N_10101,N_10068);
nand U11147 (N_11147,N_10904,N_10841);
and U11148 (N_11148,N_10671,N_10242);
nand U11149 (N_11149,N_10846,N_10367);
xnor U11150 (N_11150,N_10029,N_10856);
nor U11151 (N_11151,N_10413,N_10872);
or U11152 (N_11152,N_10605,N_10237);
or U11153 (N_11153,N_10096,N_10457);
or U11154 (N_11154,N_10826,N_10750);
or U11155 (N_11155,N_10152,N_10153);
or U11156 (N_11156,N_10354,N_10157);
nand U11157 (N_11157,N_10091,N_10277);
and U11158 (N_11158,N_10172,N_10347);
nor U11159 (N_11159,N_10060,N_10739);
and U11160 (N_11160,N_10597,N_10460);
nor U11161 (N_11161,N_10427,N_10092);
nor U11162 (N_11162,N_10290,N_10752);
xnor U11163 (N_11163,N_10756,N_10702);
nor U11164 (N_11164,N_10252,N_10578);
nor U11165 (N_11165,N_10114,N_10735);
xnor U11166 (N_11166,N_10990,N_10625);
nand U11167 (N_11167,N_10135,N_10573);
and U11168 (N_11168,N_10448,N_10624);
nand U11169 (N_11169,N_10121,N_10402);
xor U11170 (N_11170,N_10088,N_10809);
or U11171 (N_11171,N_10478,N_10334);
xnor U11172 (N_11172,N_10851,N_10991);
and U11173 (N_11173,N_10196,N_10288);
nand U11174 (N_11174,N_10561,N_10226);
xnor U11175 (N_11175,N_10306,N_10424);
or U11176 (N_11176,N_10229,N_10035);
and U11177 (N_11177,N_10720,N_10221);
xnor U11178 (N_11178,N_10223,N_10962);
nand U11179 (N_11179,N_10732,N_10295);
xnor U11180 (N_11180,N_10047,N_10162);
nor U11181 (N_11181,N_10957,N_10051);
or U11182 (N_11182,N_10313,N_10054);
nand U11183 (N_11183,N_10303,N_10657);
nor U11184 (N_11184,N_10130,N_10199);
nand U11185 (N_11185,N_10080,N_10396);
xnor U11186 (N_11186,N_10170,N_10372);
or U11187 (N_11187,N_10789,N_10459);
and U11188 (N_11188,N_10183,N_10371);
and U11189 (N_11189,N_10156,N_10678);
and U11190 (N_11190,N_10233,N_10848);
xor U11191 (N_11191,N_10610,N_10083);
xor U11192 (N_11192,N_10858,N_10937);
xnor U11193 (N_11193,N_10332,N_10250);
xor U11194 (N_11194,N_10227,N_10007);
nand U11195 (N_11195,N_10483,N_10020);
nor U11196 (N_11196,N_10558,N_10879);
or U11197 (N_11197,N_10428,N_10805);
nor U11198 (N_11198,N_10914,N_10786);
nor U11199 (N_11199,N_10086,N_10934);
nor U11200 (N_11200,N_10744,N_10113);
and U11201 (N_11201,N_10340,N_10635);
or U11202 (N_11202,N_10042,N_10785);
nor U11203 (N_11203,N_10241,N_10002);
or U11204 (N_11204,N_10683,N_10835);
or U11205 (N_11205,N_10333,N_10833);
nor U11206 (N_11206,N_10792,N_10838);
nand U11207 (N_11207,N_10968,N_10244);
and U11208 (N_11208,N_10075,N_10266);
and U11209 (N_11209,N_10410,N_10001);
xnor U11210 (N_11210,N_10422,N_10896);
or U11211 (N_11211,N_10149,N_10280);
or U11212 (N_11212,N_10599,N_10842);
or U11213 (N_11213,N_10335,N_10787);
nand U11214 (N_11214,N_10939,N_10467);
and U11215 (N_11215,N_10884,N_10203);
or U11216 (N_11216,N_10399,N_10551);
nand U11217 (N_11217,N_10725,N_10673);
nor U11218 (N_11218,N_10816,N_10751);
xor U11219 (N_11219,N_10348,N_10056);
nand U11220 (N_11220,N_10312,N_10344);
or U11221 (N_11221,N_10165,N_10515);
nor U11222 (N_11222,N_10318,N_10188);
or U11223 (N_11223,N_10701,N_10944);
and U11224 (N_11224,N_10194,N_10359);
nand U11225 (N_11225,N_10697,N_10553);
nand U11226 (N_11226,N_10328,N_10097);
xor U11227 (N_11227,N_10812,N_10742);
xor U11228 (N_11228,N_10532,N_10863);
or U11229 (N_11229,N_10126,N_10727);
nor U11230 (N_11230,N_10654,N_10622);
and U11231 (N_11231,N_10245,N_10576);
and U11232 (N_11232,N_10030,N_10053);
xnor U11233 (N_11233,N_10069,N_10602);
nand U11234 (N_11234,N_10817,N_10256);
and U11235 (N_11235,N_10825,N_10609);
nand U11236 (N_11236,N_10821,N_10297);
and U11237 (N_11237,N_10981,N_10559);
nor U11238 (N_11238,N_10451,N_10081);
nor U11239 (N_11239,N_10033,N_10431);
and U11240 (N_11240,N_10248,N_10730);
xor U11241 (N_11241,N_10315,N_10320);
xor U11242 (N_11242,N_10336,N_10412);
and U11243 (N_11243,N_10184,N_10195);
nor U11244 (N_11244,N_10191,N_10022);
or U11245 (N_11245,N_10425,N_10329);
xor U11246 (N_11246,N_10370,N_10173);
nand U11247 (N_11247,N_10564,N_10908);
nand U11248 (N_11248,N_10331,N_10634);
nor U11249 (N_11249,N_10122,N_10310);
nor U11250 (N_11250,N_10615,N_10381);
nor U11251 (N_11251,N_10249,N_10586);
or U11252 (N_11252,N_10082,N_10181);
nand U11253 (N_11253,N_10111,N_10807);
or U11254 (N_11254,N_10267,N_10269);
nor U11255 (N_11255,N_10151,N_10606);
or U11256 (N_11256,N_10453,N_10708);
or U11257 (N_11257,N_10831,N_10094);
nor U11258 (N_11258,N_10136,N_10923);
nor U11259 (N_11259,N_10182,N_10444);
nor U11260 (N_11260,N_10216,N_10493);
nand U11261 (N_11261,N_10044,N_10870);
nor U11262 (N_11262,N_10688,N_10681);
or U11263 (N_11263,N_10759,N_10034);
nand U11264 (N_11264,N_10728,N_10547);
and U11265 (N_11265,N_10992,N_10133);
nor U11266 (N_11266,N_10150,N_10255);
nand U11267 (N_11267,N_10384,N_10400);
and U11268 (N_11268,N_10146,N_10342);
nor U11269 (N_11269,N_10544,N_10651);
nand U11270 (N_11270,N_10726,N_10960);
nand U11271 (N_11271,N_10740,N_10741);
xnor U11272 (N_11272,N_10888,N_10218);
or U11273 (N_11273,N_10653,N_10202);
or U11274 (N_11274,N_10210,N_10128);
xnor U11275 (N_11275,N_10899,N_10545);
and U11276 (N_11276,N_10803,N_10510);
nor U11277 (N_11277,N_10160,N_10662);
nand U11278 (N_11278,N_10443,N_10994);
and U11279 (N_11279,N_10938,N_10067);
or U11280 (N_11280,N_10327,N_10192);
xor U11281 (N_11281,N_10810,N_10762);
nor U11282 (N_11282,N_10717,N_10768);
or U11283 (N_11283,N_10494,N_10275);
xnor U11284 (N_11284,N_10040,N_10890);
or U11285 (N_11285,N_10305,N_10360);
and U11286 (N_11286,N_10511,N_10584);
and U11287 (N_11287,N_10039,N_10799);
or U11288 (N_11288,N_10758,N_10099);
nor U11289 (N_11289,N_10648,N_10061);
nand U11290 (N_11290,N_10065,N_10643);
and U11291 (N_11291,N_10043,N_10925);
or U11292 (N_11292,N_10936,N_10124);
nand U11293 (N_11293,N_10147,N_10922);
and U11294 (N_11294,N_10268,N_10011);
and U11295 (N_11295,N_10501,N_10308);
nand U11296 (N_11296,N_10801,N_10721);
nor U11297 (N_11297,N_10746,N_10528);
nand U11298 (N_11298,N_10358,N_10475);
and U11299 (N_11299,N_10596,N_10788);
nor U11300 (N_11300,N_10572,N_10246);
and U11301 (N_11301,N_10307,N_10680);
nor U11302 (N_11302,N_10907,N_10155);
and U11303 (N_11303,N_10038,N_10148);
or U11304 (N_11304,N_10445,N_10696);
xnor U11305 (N_11305,N_10778,N_10257);
xnor U11306 (N_11306,N_10253,N_10105);
nand U11307 (N_11307,N_10260,N_10970);
nor U11308 (N_11308,N_10420,N_10647);
nand U11309 (N_11309,N_10102,N_10793);
nor U11310 (N_11310,N_10291,N_10108);
xnor U11311 (N_11311,N_10436,N_10066);
xor U11312 (N_11312,N_10715,N_10771);
and U11313 (N_11313,N_10350,N_10380);
nand U11314 (N_11314,N_10593,N_10820);
nor U11315 (N_11315,N_10220,N_10950);
xnor U11316 (N_11316,N_10376,N_10729);
nand U11317 (N_11317,N_10112,N_10985);
and U11318 (N_11318,N_10770,N_10819);
and U11319 (N_11319,N_10587,N_10583);
xor U11320 (N_11320,N_10883,N_10935);
nand U11321 (N_11321,N_10865,N_10560);
and U11322 (N_11322,N_10014,N_10430);
or U11323 (N_11323,N_10522,N_10714);
nor U11324 (N_11324,N_10325,N_10055);
or U11325 (N_11325,N_10316,N_10197);
nor U11326 (N_11326,N_10640,N_10698);
nor U11327 (N_11327,N_10611,N_10588);
and U11328 (N_11328,N_10447,N_10905);
xnor U11329 (N_11329,N_10379,N_10322);
or U11330 (N_11330,N_10123,N_10540);
xnor U11331 (N_11331,N_10999,N_10225);
and U11332 (N_11332,N_10074,N_10476);
and U11333 (N_11333,N_10901,N_10504);
or U11334 (N_11334,N_10784,N_10131);
and U11335 (N_11335,N_10982,N_10554);
or U11336 (N_11336,N_10321,N_10637);
nor U11337 (N_11337,N_10403,N_10200);
nor U11338 (N_11338,N_10892,N_10948);
nor U11339 (N_11339,N_10813,N_10283);
and U11340 (N_11340,N_10854,N_10498);
or U11341 (N_11341,N_10154,N_10265);
nand U11342 (N_11342,N_10984,N_10026);
nor U11343 (N_11343,N_10357,N_10045);
xor U11344 (N_11344,N_10766,N_10006);
and U11345 (N_11345,N_10630,N_10479);
nand U11346 (N_11346,N_10808,N_10674);
nand U11347 (N_11347,N_10952,N_10394);
nor U11348 (N_11348,N_10383,N_10875);
and U11349 (N_11349,N_10204,N_10259);
or U11350 (N_11350,N_10481,N_10882);
xnor U11351 (N_11351,N_10520,N_10595);
or U11352 (N_11352,N_10046,N_10839);
or U11353 (N_11353,N_10228,N_10037);
xor U11354 (N_11354,N_10915,N_10361);
and U11355 (N_11355,N_10723,N_10738);
or U11356 (N_11356,N_10916,N_10355);
xnor U11357 (N_11357,N_10440,N_10941);
nand U11358 (N_11358,N_10894,N_10408);
and U11359 (N_11359,N_10251,N_10100);
nand U11360 (N_11360,N_10818,N_10209);
and U11361 (N_11361,N_10663,N_10660);
nand U11362 (N_11362,N_10830,N_10294);
xor U11363 (N_11363,N_10763,N_10687);
and U11364 (N_11364,N_10893,N_10806);
or U11365 (N_11365,N_10239,N_10536);
nand U11366 (N_11366,N_10646,N_10185);
xnor U11367 (N_11367,N_10177,N_10138);
nor U11368 (N_11368,N_10628,N_10490);
nand U11369 (N_11369,N_10063,N_10645);
nor U11370 (N_11370,N_10676,N_10867);
nor U11371 (N_11371,N_10211,N_10298);
or U11372 (N_11372,N_10208,N_10926);
nor U11373 (N_11373,N_10955,N_10519);
xor U11374 (N_11374,N_10488,N_10546);
nor U11375 (N_11375,N_10311,N_10058);
or U11376 (N_11376,N_10917,N_10292);
nand U11377 (N_11377,N_10940,N_10980);
nor U11378 (N_11378,N_10282,N_10945);
or U11379 (N_11379,N_10406,N_10682);
or U11380 (N_11380,N_10362,N_10212);
nor U11381 (N_11381,N_10411,N_10704);
or U11382 (N_11382,N_10592,N_10174);
nand U11383 (N_11383,N_10049,N_10299);
nor U11384 (N_11384,N_10207,N_10710);
xnor U11385 (N_11385,N_10119,N_10782);
and U11386 (N_11386,N_10776,N_10664);
or U11387 (N_11387,N_10423,N_10656);
xnor U11388 (N_11388,N_10675,N_10169);
xnor U11389 (N_11389,N_10639,N_10765);
and U11390 (N_11390,N_10734,N_10071);
and U11391 (N_11391,N_10338,N_10798);
and U11392 (N_11392,N_10190,N_10052);
xnor U11393 (N_11393,N_10432,N_10946);
nor U11394 (N_11394,N_10880,N_10446);
xor U11395 (N_11395,N_10189,N_10254);
and U11396 (N_11396,N_10089,N_10098);
xor U11397 (N_11397,N_10013,N_10385);
nand U11398 (N_11398,N_10565,N_10041);
nor U11399 (N_11399,N_10441,N_10521);
and U11400 (N_11400,N_10368,N_10815);
nor U11401 (N_11401,N_10008,N_10247);
and U11402 (N_11402,N_10804,N_10017);
nor U11403 (N_11403,N_10977,N_10437);
or U11404 (N_11404,N_10824,N_10603);
and U11405 (N_11405,N_10296,N_10461);
xor U11406 (N_11406,N_10414,N_10222);
nand U11407 (N_11407,N_10487,N_10989);
xnor U11408 (N_11408,N_10234,N_10997);
nor U11409 (N_11409,N_10929,N_10416);
or U11410 (N_11410,N_10909,N_10800);
and U11411 (N_11411,N_10747,N_10090);
nand U11412 (N_11412,N_10885,N_10949);
nor U11413 (N_11413,N_10434,N_10391);
or U11414 (N_11414,N_10757,N_10415);
nand U11415 (N_11415,N_10903,N_10118);
nand U11416 (N_11416,N_10530,N_10988);
nand U11417 (N_11417,N_10474,N_10632);
nor U11418 (N_11418,N_10106,N_10390);
xnor U11419 (N_11419,N_10797,N_10694);
and U11420 (N_11420,N_10986,N_10722);
nand U11421 (N_11421,N_10140,N_10085);
xor U11422 (N_11422,N_10134,N_10393);
nand U11423 (N_11423,N_10193,N_10491);
nor U11424 (N_11424,N_10300,N_10070);
or U11425 (N_11425,N_10144,N_10873);
or U11426 (N_11426,N_10517,N_10513);
and U11427 (N_11427,N_10670,N_10145);
xnor U11428 (N_11428,N_10345,N_10921);
and U11429 (N_11429,N_10781,N_10796);
and U11430 (N_11430,N_10617,N_10273);
nor U11431 (N_11431,N_10961,N_10000);
or U11432 (N_11432,N_10638,N_10928);
xor U11433 (N_11433,N_10724,N_10353);
and U11434 (N_11434,N_10104,N_10972);
and U11435 (N_11435,N_10048,N_10373);
nand U11436 (N_11436,N_10852,N_10877);
or U11437 (N_11437,N_10912,N_10398);
and U11438 (N_11438,N_10604,N_10388);
xnor U11439 (N_11439,N_10878,N_10497);
and U11440 (N_11440,N_10330,N_10612);
or U11441 (N_11441,N_10644,N_10141);
and U11442 (N_11442,N_10802,N_10760);
or U11443 (N_11443,N_10389,N_10509);
nand U11444 (N_11444,N_10631,N_10613);
xnor U11445 (N_11445,N_10665,N_10514);
and U11446 (N_11446,N_10539,N_10650);
or U11447 (N_11447,N_10580,N_10794);
or U11448 (N_11448,N_10452,N_10954);
and U11449 (N_11449,N_10116,N_10016);
or U11450 (N_11450,N_10627,N_10272);
xnor U11451 (N_11451,N_10823,N_10139);
nand U11452 (N_11452,N_10672,N_10616);
or U11453 (N_11453,N_10284,N_10142);
and U11454 (N_11454,N_10025,N_10392);
or U11455 (N_11455,N_10240,N_10186);
nand U11456 (N_11456,N_10365,N_10898);
or U11457 (N_11457,N_10232,N_10117);
xor U11458 (N_11458,N_10607,N_10619);
xor U11459 (N_11459,N_10004,N_10314);
or U11460 (N_11460,N_10600,N_10589);
and U11461 (N_11461,N_10401,N_10161);
xnor U11462 (N_11462,N_10489,N_10084);
nand U11463 (N_11463,N_10073,N_10861);
and U11464 (N_11464,N_10326,N_10523);
nor U11465 (N_11465,N_10419,N_10843);
or U11466 (N_11466,N_10378,N_10951);
nor U11467 (N_11467,N_10324,N_10601);
or U11468 (N_11468,N_10455,N_10932);
nand U11469 (N_11469,N_10897,N_10920);
xor U11470 (N_11470,N_10534,N_10417);
xor U11471 (N_11471,N_10737,N_10582);
nor U11472 (N_11472,N_10827,N_10236);
or U11473 (N_11473,N_10869,N_10996);
or U11474 (N_11474,N_10127,N_10364);
and U11475 (N_11475,N_10585,N_10577);
or U11476 (N_11476,N_10435,N_10749);
nor U11477 (N_11477,N_10395,N_10579);
and U11478 (N_11478,N_10755,N_10538);
or U11479 (N_11479,N_10397,N_10707);
and U11480 (N_11480,N_10864,N_10171);
xnor U11481 (N_11481,N_10471,N_10369);
xor U11482 (N_11482,N_10686,N_10438);
nor U11483 (N_11483,N_10552,N_10339);
nor U11484 (N_11484,N_10953,N_10346);
and U11485 (N_11485,N_10775,N_10302);
nand U11486 (N_11486,N_10566,N_10258);
and U11487 (N_11487,N_10859,N_10433);
nor U11488 (N_11488,N_10699,N_10975);
nand U11489 (N_11489,N_10163,N_10652);
nor U11490 (N_11490,N_10575,N_10477);
nor U11491 (N_11491,N_10943,N_10180);
xor U11492 (N_11492,N_10690,N_10499);
or U11493 (N_11493,N_10947,N_10549);
nand U11494 (N_11494,N_10973,N_10027);
nand U11495 (N_11495,N_10005,N_10518);
nor U11496 (N_11496,N_10783,N_10974);
xnor U11497 (N_11497,N_10429,N_10032);
or U11498 (N_11498,N_10618,N_10959);
or U11499 (N_11499,N_10874,N_10889);
nand U11500 (N_11500,N_10254,N_10181);
xnor U11501 (N_11501,N_10289,N_10400);
and U11502 (N_11502,N_10493,N_10348);
nand U11503 (N_11503,N_10537,N_10745);
and U11504 (N_11504,N_10508,N_10874);
and U11505 (N_11505,N_10538,N_10980);
xnor U11506 (N_11506,N_10675,N_10610);
xnor U11507 (N_11507,N_10739,N_10261);
or U11508 (N_11508,N_10115,N_10905);
xnor U11509 (N_11509,N_10360,N_10308);
and U11510 (N_11510,N_10392,N_10433);
or U11511 (N_11511,N_10041,N_10857);
nand U11512 (N_11512,N_10368,N_10602);
or U11513 (N_11513,N_10623,N_10496);
and U11514 (N_11514,N_10422,N_10836);
nor U11515 (N_11515,N_10583,N_10038);
xor U11516 (N_11516,N_10639,N_10477);
or U11517 (N_11517,N_10121,N_10714);
or U11518 (N_11518,N_10028,N_10775);
nor U11519 (N_11519,N_10657,N_10269);
xnor U11520 (N_11520,N_10931,N_10301);
or U11521 (N_11521,N_10764,N_10609);
xor U11522 (N_11522,N_10719,N_10694);
or U11523 (N_11523,N_10115,N_10892);
nand U11524 (N_11524,N_10106,N_10837);
nor U11525 (N_11525,N_10320,N_10681);
and U11526 (N_11526,N_10607,N_10151);
or U11527 (N_11527,N_10256,N_10842);
and U11528 (N_11528,N_10423,N_10413);
nand U11529 (N_11529,N_10777,N_10824);
nor U11530 (N_11530,N_10124,N_10604);
or U11531 (N_11531,N_10706,N_10908);
nor U11532 (N_11532,N_10392,N_10500);
nor U11533 (N_11533,N_10133,N_10548);
and U11534 (N_11534,N_10712,N_10115);
nor U11535 (N_11535,N_10698,N_10277);
or U11536 (N_11536,N_10753,N_10660);
or U11537 (N_11537,N_10178,N_10675);
nor U11538 (N_11538,N_10615,N_10963);
or U11539 (N_11539,N_10214,N_10947);
or U11540 (N_11540,N_10482,N_10233);
nand U11541 (N_11541,N_10867,N_10959);
xnor U11542 (N_11542,N_10718,N_10595);
nand U11543 (N_11543,N_10286,N_10428);
and U11544 (N_11544,N_10264,N_10920);
xor U11545 (N_11545,N_10606,N_10352);
nand U11546 (N_11546,N_10604,N_10947);
and U11547 (N_11547,N_10935,N_10326);
xnor U11548 (N_11548,N_10640,N_10696);
and U11549 (N_11549,N_10768,N_10854);
nand U11550 (N_11550,N_10568,N_10343);
xnor U11551 (N_11551,N_10389,N_10139);
nor U11552 (N_11552,N_10443,N_10831);
nand U11553 (N_11553,N_10134,N_10762);
nor U11554 (N_11554,N_10738,N_10991);
xnor U11555 (N_11555,N_10632,N_10679);
and U11556 (N_11556,N_10709,N_10772);
nor U11557 (N_11557,N_10071,N_10669);
nand U11558 (N_11558,N_10598,N_10213);
or U11559 (N_11559,N_10065,N_10634);
nor U11560 (N_11560,N_10238,N_10561);
nand U11561 (N_11561,N_10149,N_10628);
nand U11562 (N_11562,N_10632,N_10551);
nand U11563 (N_11563,N_10445,N_10535);
nand U11564 (N_11564,N_10952,N_10970);
and U11565 (N_11565,N_10178,N_10373);
nor U11566 (N_11566,N_10556,N_10546);
and U11567 (N_11567,N_10309,N_10373);
nor U11568 (N_11568,N_10777,N_10753);
nand U11569 (N_11569,N_10354,N_10178);
nand U11570 (N_11570,N_10294,N_10716);
nor U11571 (N_11571,N_10957,N_10234);
xnor U11572 (N_11572,N_10986,N_10014);
or U11573 (N_11573,N_10813,N_10293);
nand U11574 (N_11574,N_10288,N_10007);
nand U11575 (N_11575,N_10538,N_10853);
nand U11576 (N_11576,N_10792,N_10625);
nor U11577 (N_11577,N_10003,N_10139);
and U11578 (N_11578,N_10510,N_10220);
xnor U11579 (N_11579,N_10471,N_10727);
xnor U11580 (N_11580,N_10990,N_10654);
nor U11581 (N_11581,N_10576,N_10003);
xor U11582 (N_11582,N_10645,N_10752);
nor U11583 (N_11583,N_10246,N_10360);
xnor U11584 (N_11584,N_10191,N_10428);
xnor U11585 (N_11585,N_10705,N_10962);
nor U11586 (N_11586,N_10246,N_10150);
xnor U11587 (N_11587,N_10013,N_10931);
nor U11588 (N_11588,N_10898,N_10391);
and U11589 (N_11589,N_10546,N_10441);
xnor U11590 (N_11590,N_10591,N_10071);
and U11591 (N_11591,N_10420,N_10202);
or U11592 (N_11592,N_10436,N_10782);
xnor U11593 (N_11593,N_10908,N_10531);
nor U11594 (N_11594,N_10136,N_10788);
and U11595 (N_11595,N_10135,N_10517);
nand U11596 (N_11596,N_10317,N_10085);
xnor U11597 (N_11597,N_10508,N_10749);
or U11598 (N_11598,N_10731,N_10600);
xnor U11599 (N_11599,N_10487,N_10094);
nand U11600 (N_11600,N_10343,N_10840);
or U11601 (N_11601,N_10477,N_10104);
or U11602 (N_11602,N_10604,N_10760);
nand U11603 (N_11603,N_10087,N_10822);
and U11604 (N_11604,N_10382,N_10787);
nand U11605 (N_11605,N_10313,N_10770);
nor U11606 (N_11606,N_10099,N_10797);
xor U11607 (N_11607,N_10678,N_10848);
nand U11608 (N_11608,N_10260,N_10112);
or U11609 (N_11609,N_10104,N_10795);
nor U11610 (N_11610,N_10615,N_10789);
nand U11611 (N_11611,N_10554,N_10253);
and U11612 (N_11612,N_10082,N_10617);
or U11613 (N_11613,N_10770,N_10617);
or U11614 (N_11614,N_10821,N_10920);
nor U11615 (N_11615,N_10188,N_10789);
nand U11616 (N_11616,N_10721,N_10678);
or U11617 (N_11617,N_10838,N_10962);
and U11618 (N_11618,N_10544,N_10258);
and U11619 (N_11619,N_10394,N_10701);
or U11620 (N_11620,N_10975,N_10686);
or U11621 (N_11621,N_10464,N_10720);
and U11622 (N_11622,N_10029,N_10829);
xor U11623 (N_11623,N_10295,N_10930);
or U11624 (N_11624,N_10692,N_10903);
nand U11625 (N_11625,N_10702,N_10855);
and U11626 (N_11626,N_10079,N_10848);
nor U11627 (N_11627,N_10907,N_10773);
nor U11628 (N_11628,N_10733,N_10740);
xor U11629 (N_11629,N_10150,N_10771);
and U11630 (N_11630,N_10539,N_10146);
xnor U11631 (N_11631,N_10547,N_10063);
and U11632 (N_11632,N_10669,N_10708);
and U11633 (N_11633,N_10497,N_10345);
xor U11634 (N_11634,N_10965,N_10785);
or U11635 (N_11635,N_10295,N_10508);
or U11636 (N_11636,N_10731,N_10210);
or U11637 (N_11637,N_10685,N_10702);
nor U11638 (N_11638,N_10109,N_10012);
or U11639 (N_11639,N_10558,N_10665);
and U11640 (N_11640,N_10856,N_10134);
and U11641 (N_11641,N_10164,N_10658);
or U11642 (N_11642,N_10942,N_10968);
xnor U11643 (N_11643,N_10581,N_10343);
nand U11644 (N_11644,N_10007,N_10089);
or U11645 (N_11645,N_10012,N_10412);
nor U11646 (N_11646,N_10384,N_10279);
or U11647 (N_11647,N_10066,N_10431);
and U11648 (N_11648,N_10113,N_10536);
and U11649 (N_11649,N_10218,N_10428);
xnor U11650 (N_11650,N_10718,N_10945);
nand U11651 (N_11651,N_10976,N_10650);
nor U11652 (N_11652,N_10894,N_10883);
nor U11653 (N_11653,N_10620,N_10835);
and U11654 (N_11654,N_10480,N_10531);
and U11655 (N_11655,N_10302,N_10074);
xor U11656 (N_11656,N_10366,N_10857);
nand U11657 (N_11657,N_10497,N_10762);
xor U11658 (N_11658,N_10354,N_10046);
nand U11659 (N_11659,N_10472,N_10385);
and U11660 (N_11660,N_10081,N_10621);
or U11661 (N_11661,N_10652,N_10183);
or U11662 (N_11662,N_10468,N_10077);
nor U11663 (N_11663,N_10538,N_10659);
xnor U11664 (N_11664,N_10378,N_10927);
nor U11665 (N_11665,N_10457,N_10322);
xnor U11666 (N_11666,N_10635,N_10892);
nor U11667 (N_11667,N_10852,N_10054);
nand U11668 (N_11668,N_10843,N_10319);
nor U11669 (N_11669,N_10971,N_10140);
xor U11670 (N_11670,N_10992,N_10263);
or U11671 (N_11671,N_10680,N_10486);
nor U11672 (N_11672,N_10958,N_10250);
or U11673 (N_11673,N_10596,N_10712);
nor U11674 (N_11674,N_10805,N_10785);
or U11675 (N_11675,N_10292,N_10064);
or U11676 (N_11676,N_10711,N_10395);
xnor U11677 (N_11677,N_10634,N_10535);
nand U11678 (N_11678,N_10797,N_10247);
or U11679 (N_11679,N_10645,N_10113);
and U11680 (N_11680,N_10920,N_10204);
and U11681 (N_11681,N_10392,N_10087);
and U11682 (N_11682,N_10239,N_10289);
or U11683 (N_11683,N_10471,N_10498);
or U11684 (N_11684,N_10144,N_10071);
xnor U11685 (N_11685,N_10680,N_10007);
nor U11686 (N_11686,N_10878,N_10603);
or U11687 (N_11687,N_10643,N_10296);
and U11688 (N_11688,N_10095,N_10438);
or U11689 (N_11689,N_10378,N_10463);
xor U11690 (N_11690,N_10199,N_10480);
nor U11691 (N_11691,N_10848,N_10376);
and U11692 (N_11692,N_10586,N_10137);
xnor U11693 (N_11693,N_10483,N_10532);
xnor U11694 (N_11694,N_10824,N_10347);
nor U11695 (N_11695,N_10284,N_10299);
nor U11696 (N_11696,N_10491,N_10452);
nor U11697 (N_11697,N_10849,N_10729);
and U11698 (N_11698,N_10796,N_10318);
nand U11699 (N_11699,N_10603,N_10394);
nand U11700 (N_11700,N_10816,N_10662);
nor U11701 (N_11701,N_10821,N_10887);
and U11702 (N_11702,N_10944,N_10685);
or U11703 (N_11703,N_10203,N_10679);
and U11704 (N_11704,N_10099,N_10694);
nor U11705 (N_11705,N_10465,N_10849);
nor U11706 (N_11706,N_10147,N_10706);
nor U11707 (N_11707,N_10728,N_10706);
nand U11708 (N_11708,N_10331,N_10124);
xor U11709 (N_11709,N_10565,N_10190);
or U11710 (N_11710,N_10823,N_10685);
or U11711 (N_11711,N_10125,N_10994);
nand U11712 (N_11712,N_10265,N_10076);
or U11713 (N_11713,N_10128,N_10891);
nor U11714 (N_11714,N_10794,N_10828);
xor U11715 (N_11715,N_10977,N_10905);
nand U11716 (N_11716,N_10566,N_10170);
xor U11717 (N_11717,N_10018,N_10601);
xor U11718 (N_11718,N_10706,N_10847);
nor U11719 (N_11719,N_10368,N_10323);
xor U11720 (N_11720,N_10435,N_10057);
and U11721 (N_11721,N_10146,N_10814);
nand U11722 (N_11722,N_10190,N_10821);
xor U11723 (N_11723,N_10930,N_10206);
nor U11724 (N_11724,N_10065,N_10649);
xnor U11725 (N_11725,N_10261,N_10243);
xor U11726 (N_11726,N_10319,N_10611);
xor U11727 (N_11727,N_10174,N_10100);
nor U11728 (N_11728,N_10767,N_10774);
nand U11729 (N_11729,N_10239,N_10697);
xnor U11730 (N_11730,N_10073,N_10756);
or U11731 (N_11731,N_10053,N_10235);
nand U11732 (N_11732,N_10572,N_10839);
or U11733 (N_11733,N_10461,N_10030);
and U11734 (N_11734,N_10875,N_10089);
nor U11735 (N_11735,N_10283,N_10754);
or U11736 (N_11736,N_10117,N_10643);
nor U11737 (N_11737,N_10176,N_10955);
nor U11738 (N_11738,N_10907,N_10671);
nor U11739 (N_11739,N_10954,N_10383);
nand U11740 (N_11740,N_10163,N_10790);
or U11741 (N_11741,N_10678,N_10291);
or U11742 (N_11742,N_10243,N_10336);
xnor U11743 (N_11743,N_10477,N_10346);
xor U11744 (N_11744,N_10670,N_10136);
nor U11745 (N_11745,N_10126,N_10286);
nor U11746 (N_11746,N_10584,N_10096);
or U11747 (N_11747,N_10038,N_10899);
nor U11748 (N_11748,N_10178,N_10097);
nand U11749 (N_11749,N_10956,N_10303);
nor U11750 (N_11750,N_10786,N_10533);
nor U11751 (N_11751,N_10195,N_10861);
or U11752 (N_11752,N_10856,N_10670);
and U11753 (N_11753,N_10017,N_10243);
and U11754 (N_11754,N_10214,N_10221);
xor U11755 (N_11755,N_10360,N_10008);
nand U11756 (N_11756,N_10713,N_10139);
nor U11757 (N_11757,N_10359,N_10890);
or U11758 (N_11758,N_10452,N_10244);
nor U11759 (N_11759,N_10940,N_10978);
and U11760 (N_11760,N_10792,N_10805);
nor U11761 (N_11761,N_10025,N_10317);
xnor U11762 (N_11762,N_10326,N_10985);
and U11763 (N_11763,N_10293,N_10233);
xnor U11764 (N_11764,N_10213,N_10978);
nand U11765 (N_11765,N_10496,N_10967);
xor U11766 (N_11766,N_10407,N_10223);
or U11767 (N_11767,N_10642,N_10531);
or U11768 (N_11768,N_10798,N_10142);
nor U11769 (N_11769,N_10055,N_10052);
nand U11770 (N_11770,N_10666,N_10483);
xor U11771 (N_11771,N_10179,N_10917);
and U11772 (N_11772,N_10707,N_10444);
xor U11773 (N_11773,N_10470,N_10701);
or U11774 (N_11774,N_10345,N_10162);
xnor U11775 (N_11775,N_10015,N_10248);
or U11776 (N_11776,N_10812,N_10204);
and U11777 (N_11777,N_10983,N_10034);
xor U11778 (N_11778,N_10344,N_10499);
xor U11779 (N_11779,N_10632,N_10126);
nor U11780 (N_11780,N_10784,N_10884);
nor U11781 (N_11781,N_10980,N_10795);
and U11782 (N_11782,N_10027,N_10956);
and U11783 (N_11783,N_10131,N_10471);
nand U11784 (N_11784,N_10936,N_10966);
nor U11785 (N_11785,N_10290,N_10376);
or U11786 (N_11786,N_10762,N_10515);
nor U11787 (N_11787,N_10661,N_10395);
and U11788 (N_11788,N_10897,N_10800);
nor U11789 (N_11789,N_10867,N_10645);
or U11790 (N_11790,N_10792,N_10810);
or U11791 (N_11791,N_10153,N_10371);
nand U11792 (N_11792,N_10354,N_10098);
or U11793 (N_11793,N_10089,N_10378);
nand U11794 (N_11794,N_10663,N_10689);
nor U11795 (N_11795,N_10863,N_10722);
xnor U11796 (N_11796,N_10848,N_10440);
nand U11797 (N_11797,N_10656,N_10116);
nor U11798 (N_11798,N_10156,N_10559);
nand U11799 (N_11799,N_10849,N_10601);
nor U11800 (N_11800,N_10641,N_10098);
nand U11801 (N_11801,N_10772,N_10874);
nor U11802 (N_11802,N_10417,N_10192);
xnor U11803 (N_11803,N_10959,N_10197);
or U11804 (N_11804,N_10993,N_10475);
or U11805 (N_11805,N_10788,N_10907);
or U11806 (N_11806,N_10094,N_10279);
or U11807 (N_11807,N_10931,N_10529);
nand U11808 (N_11808,N_10355,N_10545);
nand U11809 (N_11809,N_10676,N_10846);
xor U11810 (N_11810,N_10263,N_10909);
nand U11811 (N_11811,N_10043,N_10286);
nor U11812 (N_11812,N_10746,N_10830);
and U11813 (N_11813,N_10637,N_10849);
nor U11814 (N_11814,N_10563,N_10411);
or U11815 (N_11815,N_10753,N_10924);
nand U11816 (N_11816,N_10466,N_10307);
or U11817 (N_11817,N_10397,N_10812);
or U11818 (N_11818,N_10705,N_10156);
xor U11819 (N_11819,N_10583,N_10030);
nand U11820 (N_11820,N_10397,N_10733);
and U11821 (N_11821,N_10885,N_10882);
and U11822 (N_11822,N_10855,N_10799);
or U11823 (N_11823,N_10060,N_10256);
nor U11824 (N_11824,N_10637,N_10946);
or U11825 (N_11825,N_10228,N_10124);
xor U11826 (N_11826,N_10118,N_10233);
nor U11827 (N_11827,N_10055,N_10654);
nor U11828 (N_11828,N_10214,N_10297);
and U11829 (N_11829,N_10419,N_10180);
or U11830 (N_11830,N_10930,N_10612);
and U11831 (N_11831,N_10811,N_10157);
nor U11832 (N_11832,N_10331,N_10957);
nand U11833 (N_11833,N_10064,N_10701);
or U11834 (N_11834,N_10478,N_10047);
and U11835 (N_11835,N_10559,N_10292);
nor U11836 (N_11836,N_10053,N_10341);
nand U11837 (N_11837,N_10939,N_10807);
or U11838 (N_11838,N_10862,N_10939);
nor U11839 (N_11839,N_10723,N_10012);
nor U11840 (N_11840,N_10718,N_10399);
nor U11841 (N_11841,N_10732,N_10085);
nand U11842 (N_11842,N_10061,N_10331);
xnor U11843 (N_11843,N_10155,N_10738);
nand U11844 (N_11844,N_10389,N_10021);
xnor U11845 (N_11845,N_10096,N_10195);
nor U11846 (N_11846,N_10675,N_10700);
and U11847 (N_11847,N_10852,N_10407);
and U11848 (N_11848,N_10079,N_10794);
nand U11849 (N_11849,N_10112,N_10101);
and U11850 (N_11850,N_10901,N_10071);
or U11851 (N_11851,N_10778,N_10373);
nor U11852 (N_11852,N_10825,N_10376);
or U11853 (N_11853,N_10212,N_10625);
nor U11854 (N_11854,N_10143,N_10551);
or U11855 (N_11855,N_10223,N_10021);
xnor U11856 (N_11856,N_10918,N_10929);
and U11857 (N_11857,N_10569,N_10126);
nor U11858 (N_11858,N_10099,N_10764);
nand U11859 (N_11859,N_10808,N_10480);
or U11860 (N_11860,N_10767,N_10983);
or U11861 (N_11861,N_10612,N_10680);
or U11862 (N_11862,N_10579,N_10439);
xnor U11863 (N_11863,N_10671,N_10178);
and U11864 (N_11864,N_10779,N_10362);
and U11865 (N_11865,N_10799,N_10730);
and U11866 (N_11866,N_10253,N_10297);
xor U11867 (N_11867,N_10279,N_10779);
nor U11868 (N_11868,N_10067,N_10016);
nor U11869 (N_11869,N_10217,N_10251);
nand U11870 (N_11870,N_10231,N_10651);
and U11871 (N_11871,N_10753,N_10052);
nor U11872 (N_11872,N_10995,N_10643);
and U11873 (N_11873,N_10491,N_10922);
and U11874 (N_11874,N_10880,N_10125);
or U11875 (N_11875,N_10130,N_10712);
xor U11876 (N_11876,N_10675,N_10649);
nand U11877 (N_11877,N_10025,N_10535);
nor U11878 (N_11878,N_10632,N_10703);
or U11879 (N_11879,N_10497,N_10305);
nand U11880 (N_11880,N_10694,N_10218);
or U11881 (N_11881,N_10511,N_10732);
nor U11882 (N_11882,N_10290,N_10282);
nand U11883 (N_11883,N_10648,N_10493);
nand U11884 (N_11884,N_10446,N_10470);
and U11885 (N_11885,N_10063,N_10453);
or U11886 (N_11886,N_10060,N_10246);
nand U11887 (N_11887,N_10046,N_10802);
nand U11888 (N_11888,N_10974,N_10865);
and U11889 (N_11889,N_10847,N_10668);
and U11890 (N_11890,N_10376,N_10648);
nand U11891 (N_11891,N_10241,N_10960);
or U11892 (N_11892,N_10630,N_10792);
or U11893 (N_11893,N_10548,N_10408);
nand U11894 (N_11894,N_10679,N_10176);
or U11895 (N_11895,N_10513,N_10538);
and U11896 (N_11896,N_10746,N_10367);
and U11897 (N_11897,N_10429,N_10113);
and U11898 (N_11898,N_10284,N_10657);
nor U11899 (N_11899,N_10331,N_10793);
xnor U11900 (N_11900,N_10562,N_10679);
or U11901 (N_11901,N_10170,N_10214);
nor U11902 (N_11902,N_10477,N_10951);
nor U11903 (N_11903,N_10893,N_10915);
nor U11904 (N_11904,N_10693,N_10548);
xor U11905 (N_11905,N_10141,N_10433);
and U11906 (N_11906,N_10945,N_10103);
nor U11907 (N_11907,N_10716,N_10389);
nand U11908 (N_11908,N_10876,N_10456);
nand U11909 (N_11909,N_10484,N_10006);
and U11910 (N_11910,N_10476,N_10960);
xnor U11911 (N_11911,N_10044,N_10731);
and U11912 (N_11912,N_10135,N_10952);
xor U11913 (N_11913,N_10923,N_10253);
or U11914 (N_11914,N_10282,N_10159);
xor U11915 (N_11915,N_10294,N_10845);
nor U11916 (N_11916,N_10042,N_10658);
xnor U11917 (N_11917,N_10192,N_10434);
or U11918 (N_11918,N_10766,N_10310);
nand U11919 (N_11919,N_10362,N_10449);
nand U11920 (N_11920,N_10500,N_10671);
nand U11921 (N_11921,N_10012,N_10065);
nand U11922 (N_11922,N_10388,N_10698);
and U11923 (N_11923,N_10507,N_10306);
nor U11924 (N_11924,N_10856,N_10957);
nor U11925 (N_11925,N_10362,N_10452);
xnor U11926 (N_11926,N_10343,N_10097);
nand U11927 (N_11927,N_10172,N_10616);
and U11928 (N_11928,N_10136,N_10894);
xnor U11929 (N_11929,N_10929,N_10937);
xnor U11930 (N_11930,N_10732,N_10621);
and U11931 (N_11931,N_10945,N_10639);
and U11932 (N_11932,N_10171,N_10109);
and U11933 (N_11933,N_10070,N_10395);
nor U11934 (N_11934,N_10122,N_10561);
and U11935 (N_11935,N_10941,N_10150);
or U11936 (N_11936,N_10056,N_10590);
or U11937 (N_11937,N_10585,N_10098);
nand U11938 (N_11938,N_10017,N_10103);
xor U11939 (N_11939,N_10674,N_10928);
or U11940 (N_11940,N_10524,N_10302);
or U11941 (N_11941,N_10766,N_10624);
and U11942 (N_11942,N_10722,N_10430);
xor U11943 (N_11943,N_10630,N_10582);
and U11944 (N_11944,N_10709,N_10386);
and U11945 (N_11945,N_10098,N_10627);
nand U11946 (N_11946,N_10738,N_10751);
xor U11947 (N_11947,N_10333,N_10369);
and U11948 (N_11948,N_10000,N_10278);
xor U11949 (N_11949,N_10757,N_10237);
or U11950 (N_11950,N_10336,N_10947);
nor U11951 (N_11951,N_10894,N_10496);
nor U11952 (N_11952,N_10190,N_10727);
xnor U11953 (N_11953,N_10969,N_10542);
nand U11954 (N_11954,N_10697,N_10054);
or U11955 (N_11955,N_10420,N_10877);
nand U11956 (N_11956,N_10331,N_10753);
or U11957 (N_11957,N_10667,N_10937);
xor U11958 (N_11958,N_10617,N_10853);
and U11959 (N_11959,N_10083,N_10741);
or U11960 (N_11960,N_10563,N_10511);
nand U11961 (N_11961,N_10476,N_10764);
and U11962 (N_11962,N_10507,N_10621);
nand U11963 (N_11963,N_10697,N_10355);
nor U11964 (N_11964,N_10431,N_10313);
nand U11965 (N_11965,N_10410,N_10106);
and U11966 (N_11966,N_10313,N_10921);
nand U11967 (N_11967,N_10047,N_10248);
xnor U11968 (N_11968,N_10062,N_10453);
or U11969 (N_11969,N_10010,N_10892);
or U11970 (N_11970,N_10900,N_10157);
nand U11971 (N_11971,N_10115,N_10113);
and U11972 (N_11972,N_10999,N_10316);
nor U11973 (N_11973,N_10184,N_10339);
nor U11974 (N_11974,N_10569,N_10696);
and U11975 (N_11975,N_10885,N_10371);
nor U11976 (N_11976,N_10280,N_10143);
and U11977 (N_11977,N_10223,N_10344);
and U11978 (N_11978,N_10968,N_10016);
or U11979 (N_11979,N_10167,N_10522);
nand U11980 (N_11980,N_10683,N_10288);
nand U11981 (N_11981,N_10635,N_10188);
nor U11982 (N_11982,N_10920,N_10659);
or U11983 (N_11983,N_10752,N_10419);
xnor U11984 (N_11984,N_10394,N_10481);
nor U11985 (N_11985,N_10890,N_10041);
xnor U11986 (N_11986,N_10554,N_10056);
xnor U11987 (N_11987,N_10029,N_10212);
and U11988 (N_11988,N_10311,N_10762);
or U11989 (N_11989,N_10703,N_10884);
xor U11990 (N_11990,N_10283,N_10120);
nor U11991 (N_11991,N_10669,N_10491);
xor U11992 (N_11992,N_10729,N_10113);
xnor U11993 (N_11993,N_10892,N_10206);
nand U11994 (N_11994,N_10145,N_10418);
nand U11995 (N_11995,N_10020,N_10662);
or U11996 (N_11996,N_10358,N_10253);
xor U11997 (N_11997,N_10476,N_10025);
nor U11998 (N_11998,N_10687,N_10168);
xnor U11999 (N_11999,N_10029,N_10412);
and U12000 (N_12000,N_11834,N_11964);
nand U12001 (N_12001,N_11800,N_11136);
or U12002 (N_12002,N_11357,N_11916);
nand U12003 (N_12003,N_11815,N_11752);
or U12004 (N_12004,N_11207,N_11593);
nor U12005 (N_12005,N_11313,N_11228);
or U12006 (N_12006,N_11899,N_11151);
xor U12007 (N_12007,N_11306,N_11883);
xor U12008 (N_12008,N_11147,N_11809);
and U12009 (N_12009,N_11940,N_11219);
or U12010 (N_12010,N_11702,N_11912);
nand U12011 (N_12011,N_11995,N_11783);
and U12012 (N_12012,N_11250,N_11072);
and U12013 (N_12013,N_11638,N_11927);
xnor U12014 (N_12014,N_11477,N_11914);
nand U12015 (N_12015,N_11644,N_11792);
nand U12016 (N_12016,N_11768,N_11600);
nand U12017 (N_12017,N_11101,N_11324);
or U12018 (N_12018,N_11734,N_11462);
nand U12019 (N_12019,N_11440,N_11703);
xnor U12020 (N_12020,N_11669,N_11695);
or U12021 (N_12021,N_11478,N_11741);
xor U12022 (N_12022,N_11632,N_11276);
xor U12023 (N_12023,N_11712,N_11023);
nor U12024 (N_12024,N_11405,N_11329);
xor U12025 (N_12025,N_11791,N_11260);
and U12026 (N_12026,N_11002,N_11090);
nor U12027 (N_12027,N_11731,N_11381);
or U12028 (N_12028,N_11653,N_11689);
or U12029 (N_12029,N_11528,N_11924);
nand U12030 (N_12030,N_11108,N_11256);
nand U12031 (N_12031,N_11929,N_11534);
and U12032 (N_12032,N_11105,N_11781);
nor U12033 (N_12033,N_11616,N_11141);
nor U12034 (N_12034,N_11327,N_11699);
nor U12035 (N_12035,N_11842,N_11866);
nor U12036 (N_12036,N_11513,N_11213);
xor U12037 (N_12037,N_11038,N_11142);
xor U12038 (N_12038,N_11379,N_11015);
or U12039 (N_12039,N_11227,N_11846);
nor U12040 (N_12040,N_11540,N_11861);
and U12041 (N_12041,N_11320,N_11220);
or U12042 (N_12042,N_11655,N_11085);
or U12043 (N_12043,N_11216,N_11976);
and U12044 (N_12044,N_11847,N_11458);
or U12045 (N_12045,N_11547,N_11434);
nand U12046 (N_12046,N_11596,N_11167);
xnor U12047 (N_12047,N_11884,N_11523);
nand U12048 (N_12048,N_11612,N_11541);
nand U12049 (N_12049,N_11749,N_11340);
and U12050 (N_12050,N_11121,N_11131);
xnor U12051 (N_12051,N_11195,N_11806);
xor U12052 (N_12052,N_11971,N_11438);
nor U12053 (N_12053,N_11139,N_11660);
nor U12054 (N_12054,N_11039,N_11410);
nor U12055 (N_12055,N_11646,N_11514);
xor U12056 (N_12056,N_11175,N_11822);
and U12057 (N_12057,N_11897,N_11425);
or U12058 (N_12058,N_11177,N_11988);
nor U12059 (N_12059,N_11074,N_11608);
nand U12060 (N_12060,N_11642,N_11271);
nand U12061 (N_12061,N_11209,N_11331);
xnor U12062 (N_12062,N_11365,N_11698);
and U12063 (N_12063,N_11919,N_11651);
or U12064 (N_12064,N_11443,N_11268);
xor U12065 (N_12065,N_11186,N_11479);
xnor U12066 (N_12066,N_11265,N_11771);
nor U12067 (N_12067,N_11215,N_11587);
or U12068 (N_12068,N_11965,N_11150);
or U12069 (N_12069,N_11701,N_11886);
xnor U12070 (N_12070,N_11686,N_11132);
nor U12071 (N_12071,N_11051,N_11233);
nand U12072 (N_12072,N_11526,N_11722);
or U12073 (N_12073,N_11003,N_11188);
or U12074 (N_12074,N_11625,N_11426);
nand U12075 (N_12075,N_11252,N_11432);
nand U12076 (N_12076,N_11048,N_11640);
xor U12077 (N_12077,N_11521,N_11077);
nor U12078 (N_12078,N_11575,N_11578);
nand U12079 (N_12079,N_11647,N_11400);
nor U12080 (N_12080,N_11774,N_11730);
nand U12081 (N_12081,N_11095,N_11392);
and U12082 (N_12082,N_11495,N_11355);
xnor U12083 (N_12083,N_11394,N_11614);
xnor U12084 (N_12084,N_11423,N_11981);
xnor U12085 (N_12085,N_11527,N_11556);
or U12086 (N_12086,N_11571,N_11404);
or U12087 (N_12087,N_11374,N_11648);
or U12088 (N_12088,N_11214,N_11588);
nor U12089 (N_12089,N_11737,N_11533);
nor U12090 (N_12090,N_11020,N_11166);
or U12091 (N_12091,N_11302,N_11990);
nor U12092 (N_12092,N_11532,N_11145);
nand U12093 (N_12093,N_11247,N_11202);
nand U12094 (N_12094,N_11187,N_11645);
or U12095 (N_12095,N_11603,N_11429);
or U12096 (N_12096,N_11666,N_11558);
nand U12097 (N_12097,N_11871,N_11945);
or U12098 (N_12098,N_11333,N_11129);
nor U12099 (N_12099,N_11909,N_11637);
xnor U12100 (N_12100,N_11467,N_11218);
xnor U12101 (N_12101,N_11933,N_11344);
and U12102 (N_12102,N_11113,N_11179);
xnor U12103 (N_12103,N_11253,N_11386);
nand U12104 (N_12104,N_11862,N_11497);
nor U12105 (N_12105,N_11622,N_11254);
and U12106 (N_12106,N_11041,N_11615);
or U12107 (N_12107,N_11384,N_11713);
and U12108 (N_12108,N_11165,N_11977);
and U12109 (N_12109,N_11626,N_11738);
or U12110 (N_12110,N_11144,N_11787);
nand U12111 (N_12111,N_11110,N_11249);
or U12112 (N_12112,N_11934,N_11821);
nand U12113 (N_12113,N_11500,N_11865);
nand U12114 (N_12114,N_11753,N_11760);
and U12115 (N_12115,N_11062,N_11114);
nand U12116 (N_12116,N_11750,N_11989);
nor U12117 (N_12117,N_11745,N_11631);
and U12118 (N_12118,N_11829,N_11030);
or U12119 (N_12119,N_11830,N_11696);
nor U12120 (N_12120,N_11487,N_11880);
xnor U12121 (N_12121,N_11430,N_11162);
nand U12122 (N_12122,N_11305,N_11549);
nand U12123 (N_12123,N_11224,N_11818);
or U12124 (N_12124,N_11568,N_11287);
nand U12125 (N_12125,N_11820,N_11735);
or U12126 (N_12126,N_11468,N_11805);
nand U12127 (N_12127,N_11721,N_11785);
xor U12128 (N_12128,N_11751,N_11649);
nand U12129 (N_12129,N_11053,N_11456);
xnor U12130 (N_12130,N_11788,N_11087);
nor U12131 (N_12131,N_11494,N_11295);
nand U12132 (N_12132,N_11368,N_11470);
and U12133 (N_12133,N_11481,N_11773);
and U12134 (N_12134,N_11537,N_11480);
nand U12135 (N_12135,N_11986,N_11552);
xor U12136 (N_12136,N_11402,N_11812);
and U12137 (N_12137,N_11396,N_11421);
nor U12138 (N_12138,N_11780,N_11611);
or U12139 (N_12139,N_11706,N_11678);
xor U12140 (N_12140,N_11503,N_11281);
nand U12141 (N_12141,N_11399,N_11086);
xnor U12142 (N_12142,N_11684,N_11566);
nand U12143 (N_12143,N_11951,N_11453);
and U12144 (N_12144,N_11855,N_11754);
xnor U12145 (N_12145,N_11153,N_11089);
nand U12146 (N_12146,N_11512,N_11868);
or U12147 (N_12147,N_11967,N_11229);
and U12148 (N_12148,N_11825,N_11044);
nor U12149 (N_12149,N_11992,N_11941);
nand U12150 (N_12150,N_11289,N_11057);
nor U12151 (N_12151,N_11583,N_11665);
or U12152 (N_12152,N_11601,N_11431);
nor U12153 (N_12153,N_11518,N_11908);
nor U12154 (N_12154,N_11406,N_11504);
and U12155 (N_12155,N_11314,N_11437);
or U12156 (N_12156,N_11688,N_11881);
and U12157 (N_12157,N_11275,N_11635);
nand U12158 (N_12158,N_11102,N_11624);
and U12159 (N_12159,N_11683,N_11409);
and U12160 (N_12160,N_11729,N_11137);
and U12161 (N_12161,N_11459,N_11192);
and U12162 (N_12162,N_11234,N_11982);
nor U12163 (N_12163,N_11138,N_11762);
xnor U12164 (N_12164,N_11032,N_11975);
xnor U12165 (N_12165,N_11063,N_11013);
nor U12166 (N_12166,N_11336,N_11980);
nand U12167 (N_12167,N_11045,N_11170);
nor U12168 (N_12168,N_11303,N_11391);
or U12169 (N_12169,N_11100,N_11461);
or U12170 (N_12170,N_11873,N_11180);
or U12171 (N_12171,N_11326,N_11067);
nor U12172 (N_12172,N_11439,N_11661);
or U12173 (N_12173,N_11064,N_11682);
or U12174 (N_12174,N_11913,N_11872);
nand U12175 (N_12175,N_11577,N_11312);
nand U12176 (N_12176,N_11841,N_11562);
and U12177 (N_12177,N_11525,N_11375);
xor U12178 (N_12178,N_11485,N_11436);
nor U12179 (N_12179,N_11049,N_11888);
and U12180 (N_12180,N_11026,N_11538);
and U12181 (N_12181,N_11621,N_11910);
xnor U12182 (N_12182,N_11553,N_11206);
nor U12183 (N_12183,N_11304,N_11168);
nand U12184 (N_12184,N_11455,N_11288);
nand U12185 (N_12185,N_11733,N_11770);
xor U12186 (N_12186,N_11687,N_11955);
nor U12187 (N_12187,N_11911,N_11850);
or U12188 (N_12188,N_11483,N_11623);
and U12189 (N_12189,N_11383,N_11418);
xnor U12190 (N_12190,N_11799,N_11226);
or U12191 (N_12191,N_11146,N_11189);
or U12192 (N_12192,N_11205,N_11958);
nor U12193 (N_12193,N_11983,N_11663);
and U12194 (N_12194,N_11726,N_11870);
and U12195 (N_12195,N_11991,N_11435);
or U12196 (N_12196,N_11125,N_11922);
nand U12197 (N_12197,N_11671,N_11832);
and U12198 (N_12198,N_11382,N_11096);
xnor U12199 (N_12199,N_11349,N_11710);
nand U12200 (N_12200,N_11511,N_11182);
nor U12201 (N_12201,N_11860,N_11119);
nor U12202 (N_12202,N_11836,N_11874);
nand U12203 (N_12203,N_11973,N_11807);
and U12204 (N_12204,N_11319,N_11516);
nor U12205 (N_12205,N_11554,N_11474);
nor U12206 (N_12206,N_11446,N_11427);
nor U12207 (N_12207,N_11551,N_11068);
and U12208 (N_12208,N_11307,N_11111);
and U12209 (N_12209,N_11814,N_11962);
nand U12210 (N_12210,N_11273,N_11109);
xnor U12211 (N_12211,N_11609,N_11920);
nor U12212 (N_12212,N_11490,N_11269);
nor U12213 (N_12213,N_11579,N_11697);
and U12214 (N_12214,N_11035,N_11029);
or U12215 (N_12215,N_11448,N_11585);
nor U12216 (N_12216,N_11171,N_11685);
nand U12217 (N_12217,N_11341,N_11159);
and U12218 (N_12218,N_11184,N_11274);
nor U12219 (N_12219,N_11471,N_11546);
nand U12220 (N_12220,N_11676,N_11947);
and U12221 (N_12221,N_11237,N_11444);
nand U12222 (N_12222,N_11183,N_11008);
nor U12223 (N_12223,N_11708,N_11457);
or U12224 (N_12224,N_11084,N_11407);
nand U12225 (N_12225,N_11217,N_11393);
or U12226 (N_12226,N_11460,N_11923);
or U12227 (N_12227,N_11094,N_11321);
xnor U12228 (N_12228,N_11043,N_11364);
xor U12229 (N_12229,N_11024,N_11659);
xnor U12230 (N_12230,N_11864,N_11739);
or U12231 (N_12231,N_11816,N_11309);
or U12232 (N_12232,N_11317,N_11387);
xnor U12233 (N_12233,N_11376,N_11465);
nor U12234 (N_12234,N_11979,N_11694);
nand U12235 (N_12235,N_11529,N_11117);
nand U12236 (N_12236,N_11009,N_11058);
xnor U12237 (N_12237,N_11956,N_11763);
nand U12238 (N_12238,N_11299,N_11291);
or U12239 (N_12239,N_11498,N_11796);
nor U12240 (N_12240,N_11025,N_11362);
and U12241 (N_12241,N_11031,N_11510);
nor U12242 (N_12242,N_11681,N_11801);
xnor U12243 (N_12243,N_11335,N_11397);
or U12244 (N_12244,N_11776,N_11747);
xnor U12245 (N_12245,N_11559,N_11743);
or U12246 (N_12246,N_11416,N_11006);
nor U12247 (N_12247,N_11069,N_11598);
xnor U12248 (N_12248,N_11194,N_11853);
nand U12249 (N_12249,N_11939,N_11415);
nor U12250 (N_12250,N_11719,N_11813);
or U12251 (N_12251,N_11690,N_11264);
nand U12252 (N_12252,N_11744,N_11938);
xor U12253 (N_12253,N_11723,N_11968);
or U12254 (N_12254,N_11450,N_11879);
or U12255 (N_12255,N_11210,N_11449);
xnor U12256 (N_12256,N_11970,N_11567);
nor U12257 (N_12257,N_11769,N_11388);
xnor U12258 (N_12258,N_11896,N_11837);
nor U12259 (N_12259,N_11932,N_11042);
nand U12260 (N_12260,N_11126,N_11928);
xnor U12261 (N_12261,N_11176,N_11088);
xnor U12262 (N_12262,N_11849,N_11946);
nor U12263 (N_12263,N_11065,N_11679);
xor U12264 (N_12264,N_11358,N_11034);
nand U12265 (N_12265,N_11576,N_11059);
xor U12266 (N_12266,N_11482,N_11169);
xnor U12267 (N_12267,N_11412,N_11135);
or U12268 (N_12268,N_11654,N_11246);
xor U12269 (N_12269,N_11680,N_11627);
nand U12270 (N_12270,N_11005,N_11040);
xnor U12271 (N_12271,N_11353,N_11066);
or U12272 (N_12272,N_11520,N_11772);
xor U12273 (N_12273,N_11133,N_11011);
and U12274 (N_12274,N_11906,N_11251);
nand U12275 (N_12275,N_11036,N_11828);
nand U12276 (N_12276,N_11509,N_11028);
or U12277 (N_12277,N_11359,N_11027);
or U12278 (N_12278,N_11966,N_11301);
xor U12279 (N_12279,N_11629,N_11606);
nor U12280 (N_12280,N_11953,N_11325);
nand U12281 (N_12281,N_11047,N_11272);
nand U12282 (N_12282,N_11451,N_11351);
or U12283 (N_12283,N_11263,N_11996);
nor U12284 (N_12284,N_11954,N_11328);
or U12285 (N_12285,N_11727,N_11081);
or U12286 (N_12286,N_11347,N_11193);
nor U12287 (N_12287,N_11584,N_11949);
or U12288 (N_12288,N_11904,N_11848);
nor U12289 (N_12289,N_11728,N_11157);
and U12290 (N_12290,N_11742,N_11935);
xor U12291 (N_12291,N_11185,N_11984);
and U12292 (N_12292,N_11900,N_11890);
nand U12293 (N_12293,N_11613,N_11944);
nand U12294 (N_12294,N_11824,N_11658);
nor U12295 (N_12295,N_11550,N_11574);
nor U12296 (N_12296,N_11242,N_11106);
xor U12297 (N_12297,N_11310,N_11501);
nor U12298 (N_12298,N_11535,N_11506);
or U12299 (N_12299,N_11433,N_11677);
xnor U12300 (N_12300,N_11422,N_11893);
or U12301 (N_12301,N_11280,N_11270);
nand U12302 (N_12302,N_11782,N_11191);
xor U12303 (N_12303,N_11802,N_11997);
or U12304 (N_12304,N_11856,N_11942);
and U12305 (N_12305,N_11572,N_11517);
xor U12306 (N_12306,N_11486,N_11311);
or U12307 (N_12307,N_11746,N_11238);
xor U12308 (N_12308,N_11755,N_11284);
nor U12309 (N_12309,N_11725,N_11985);
xor U12310 (N_12310,N_11158,N_11798);
xnor U12311 (N_12311,N_11972,N_11267);
nand U12312 (N_12312,N_11604,N_11122);
nand U12313 (N_12313,N_11952,N_11628);
xnor U12314 (N_12314,N_11070,N_11403);
xor U12315 (N_12315,N_11582,N_11428);
and U12316 (N_12316,N_11371,N_11083);
and U12317 (N_12317,N_11515,N_11892);
nand U12318 (N_12318,N_11931,N_11107);
nor U12319 (N_12319,N_11163,N_11491);
or U12320 (N_12320,N_11826,N_11017);
or U12321 (N_12321,N_11519,N_11877);
and U12322 (N_12322,N_11561,N_11670);
nor U12323 (N_12323,N_11367,N_11492);
nor U12324 (N_12324,N_11693,N_11573);
nor U12325 (N_12325,N_11235,N_11994);
and U12326 (N_12326,N_11560,N_11858);
or U12327 (N_12327,N_11636,N_11756);
xnor U12328 (N_12328,N_11499,N_11472);
xor U12329 (N_12329,N_11748,N_11208);
nand U12330 (N_12330,N_11948,N_11539);
and U12331 (N_12331,N_11203,N_11610);
or U12332 (N_12332,N_11212,N_11097);
or U12333 (N_12333,N_11732,N_11236);
or U12334 (N_12334,N_11673,N_11118);
xnor U12335 (N_12335,N_11718,N_11643);
xor U12336 (N_12336,N_11545,N_11859);
nand U12337 (N_12337,N_11010,N_11543);
or U12338 (N_12338,N_11290,N_11441);
or U12339 (N_12339,N_11369,N_11366);
and U12340 (N_12340,N_11707,N_11767);
nand U12341 (N_12341,N_11103,N_11876);
nor U12342 (N_12342,N_11389,N_11476);
or U12343 (N_12343,N_11259,N_11898);
nand U12344 (N_12344,N_11810,N_11116);
and U12345 (N_12345,N_11895,N_11508);
nand U12346 (N_12346,N_11078,N_11385);
xor U12347 (N_12347,N_11292,N_11338);
nand U12348 (N_12348,N_11000,N_11257);
xnor U12349 (N_12349,N_11007,N_11595);
xnor U12350 (N_12350,N_11071,N_11091);
xor U12351 (N_12351,N_11797,N_11445);
or U12352 (N_12352,N_11761,N_11123);
or U12353 (N_12353,N_11469,N_11804);
xnor U12354 (N_12354,N_11395,N_11765);
nand U12355 (N_12355,N_11925,N_11817);
nor U12356 (N_12356,N_11466,N_11452);
nor U12357 (N_12357,N_11974,N_11297);
nand U12358 (N_12358,N_11279,N_11827);
and U12359 (N_12359,N_11414,N_11076);
xor U12360 (N_12360,N_11803,N_11104);
nor U12361 (N_12361,N_11322,N_11668);
or U12362 (N_12362,N_11507,N_11843);
nor U12363 (N_12363,N_11882,N_11473);
nand U12364 (N_12364,N_11618,N_11419);
xor U12365 (N_12365,N_11149,N_11667);
xor U12366 (N_12366,N_11789,N_11092);
and U12367 (N_12367,N_11937,N_11867);
or U12368 (N_12368,N_11599,N_11323);
xor U12369 (N_12369,N_11590,N_11244);
or U12370 (N_12370,N_11190,N_11339);
and U12371 (N_12371,N_11037,N_11811);
xor U12372 (N_12372,N_11705,N_11565);
xnor U12373 (N_12373,N_11201,N_11308);
and U12374 (N_12374,N_11390,N_11156);
nor U12375 (N_12375,N_11408,N_11963);
nor U12376 (N_12376,N_11581,N_11050);
xor U12377 (N_12377,N_11283,N_11332);
nor U12378 (N_12378,N_11363,N_11709);
and U12379 (N_12379,N_11046,N_11620);
xor U12380 (N_12380,N_11542,N_11300);
or U12381 (N_12381,N_11160,N_11840);
nor U12382 (N_12382,N_11716,N_11370);
and U12383 (N_12383,N_11266,N_11969);
and U12384 (N_12384,N_11674,N_11764);
and U12385 (N_12385,N_11093,N_11346);
nand U12386 (N_12386,N_11724,N_11901);
nand U12387 (N_12387,N_11650,N_11330);
or U12388 (N_12388,N_11959,N_11348);
and U12389 (N_12389,N_11672,N_11277);
and U12390 (N_12390,N_11352,N_11127);
nand U12391 (N_12391,N_11838,N_11261);
and U12392 (N_12392,N_11484,N_11488);
nand U12393 (N_12393,N_11298,N_11278);
nand U12394 (N_12394,N_11978,N_11987);
nand U12395 (N_12395,N_11001,N_11373);
and U12396 (N_12396,N_11591,N_11350);
or U12397 (N_12397,N_11602,N_11420);
xnor U12398 (N_12398,N_11115,N_11522);
and U12399 (N_12399,N_11055,N_11926);
and U12400 (N_12400,N_11943,N_11961);
nor U12401 (N_12401,N_11079,N_11222);
nand U12402 (N_12402,N_11711,N_11502);
nand U12403 (N_12403,N_11819,N_11221);
nand U12404 (N_12404,N_11907,N_11758);
and U12405 (N_12405,N_11736,N_11835);
xnor U12406 (N_12406,N_11173,N_11960);
xor U12407 (N_12407,N_11240,N_11424);
or U12408 (N_12408,N_11164,N_11021);
or U12409 (N_12409,N_11902,N_11875);
xor U12410 (N_12410,N_11851,N_11592);
nand U12411 (N_12411,N_11905,N_11564);
or U12412 (N_12412,N_11199,N_11152);
xnor U12413 (N_12413,N_11605,N_11634);
nand U12414 (N_12414,N_11061,N_11936);
or U12415 (N_12415,N_11282,N_11148);
nand U12416 (N_12416,N_11225,N_11793);
nor U12417 (N_12417,N_11652,N_11633);
xor U12418 (N_12418,N_11315,N_11891);
xor U12419 (N_12419,N_11915,N_11442);
xnor U12420 (N_12420,N_11285,N_11293);
and U12421 (N_12421,N_11921,N_11903);
nor U12422 (N_12422,N_11957,N_11181);
and U12423 (N_12423,N_11717,N_11174);
or U12424 (N_12424,N_11857,N_11808);
xnor U12425 (N_12425,N_11714,N_11197);
nand U12426 (N_12426,N_11286,N_11918);
or U12427 (N_12427,N_11656,N_11243);
nand U12428 (N_12428,N_11475,N_11950);
nand U12429 (N_12429,N_11248,N_11447);
or U12430 (N_12430,N_11073,N_11354);
nand U12431 (N_12431,N_11361,N_11833);
nand U12432 (N_12432,N_11230,N_11178);
or U12433 (N_12433,N_11563,N_11334);
or U12434 (N_12434,N_11143,N_11245);
and U12435 (N_12435,N_11124,N_11657);
xnor U12436 (N_12436,N_11917,N_11885);
nand U12437 (N_12437,N_11134,N_11154);
or U12438 (N_12438,N_11715,N_11530);
nand U12439 (N_12439,N_11794,N_11316);
and U12440 (N_12440,N_11536,N_11255);
nor U12441 (N_12441,N_11128,N_11993);
and U12442 (N_12442,N_11200,N_11548);
nand U12443 (N_12443,N_11380,N_11417);
xnor U12444 (N_12444,N_11531,N_11544);
or U12445 (N_12445,N_11675,N_11778);
nor U12446 (N_12446,N_11413,N_11691);
or U12447 (N_12447,N_11786,N_11662);
nor U12448 (N_12448,N_11823,N_11496);
nor U12449 (N_12449,N_11524,N_11463);
nor U12450 (N_12450,N_11557,N_11777);
or U12451 (N_12451,N_11075,N_11998);
or U12452 (N_12452,N_11231,N_11296);
or U12453 (N_12453,N_11022,N_11060);
or U12454 (N_12454,N_11505,N_11795);
xnor U12455 (N_12455,N_11570,N_11080);
nor U12456 (N_12456,N_11790,N_11589);
and U12457 (N_12457,N_11869,N_11619);
nand U12458 (N_12458,N_11555,N_11757);
and U12459 (N_12459,N_11337,N_11845);
or U12460 (N_12460,N_11360,N_11014);
and U12461 (N_12461,N_11372,N_11641);
nand U12462 (N_12462,N_11894,N_11839);
xor U12463 (N_12463,N_11889,N_11082);
nor U12464 (N_12464,N_11630,N_11398);
or U12465 (N_12465,N_11239,N_11318);
nor U12466 (N_12466,N_11098,N_11198);
or U12467 (N_12467,N_11878,N_11356);
nand U12468 (N_12468,N_11378,N_11759);
or U12469 (N_12469,N_11343,N_11112);
nor U12470 (N_12470,N_11140,N_11664);
xor U12471 (N_12471,N_11033,N_11999);
and U12472 (N_12472,N_11004,N_11155);
nor U12473 (N_12473,N_11054,N_11377);
nor U12474 (N_12474,N_11852,N_11345);
nor U12475 (N_12475,N_11052,N_11012);
and U12476 (N_12476,N_11740,N_11831);
xor U12477 (N_12477,N_11161,N_11720);
or U12478 (N_12478,N_11493,N_11019);
and U12479 (N_12479,N_11258,N_11241);
xnor U12480 (N_12480,N_11223,N_11464);
xor U12481 (N_12481,N_11172,N_11196);
nand U12482 (N_12482,N_11775,N_11232);
nor U12483 (N_12483,N_11120,N_11597);
nand U12484 (N_12484,N_11692,N_11779);
nor U12485 (N_12485,N_11016,N_11580);
xnor U12486 (N_12486,N_11401,N_11639);
or U12487 (N_12487,N_11863,N_11262);
nand U12488 (N_12488,N_11784,N_11294);
and U12489 (N_12489,N_11607,N_11342);
and U12490 (N_12490,N_11454,N_11211);
nor U12491 (N_12491,N_11569,N_11056);
and U12492 (N_12492,N_11844,N_11887);
nor U12493 (N_12493,N_11018,N_11700);
nor U12494 (N_12494,N_11594,N_11489);
and U12495 (N_12495,N_11099,N_11130);
xor U12496 (N_12496,N_11617,N_11930);
xnor U12497 (N_12497,N_11411,N_11766);
or U12498 (N_12498,N_11704,N_11854);
nand U12499 (N_12499,N_11586,N_11204);
or U12500 (N_12500,N_11827,N_11215);
or U12501 (N_12501,N_11873,N_11865);
or U12502 (N_12502,N_11283,N_11643);
or U12503 (N_12503,N_11444,N_11541);
nor U12504 (N_12504,N_11278,N_11150);
xnor U12505 (N_12505,N_11692,N_11603);
xnor U12506 (N_12506,N_11340,N_11400);
nand U12507 (N_12507,N_11088,N_11648);
xnor U12508 (N_12508,N_11545,N_11617);
nor U12509 (N_12509,N_11737,N_11609);
or U12510 (N_12510,N_11823,N_11777);
and U12511 (N_12511,N_11435,N_11961);
and U12512 (N_12512,N_11273,N_11155);
xor U12513 (N_12513,N_11623,N_11488);
and U12514 (N_12514,N_11251,N_11966);
nand U12515 (N_12515,N_11831,N_11061);
nor U12516 (N_12516,N_11010,N_11630);
nor U12517 (N_12517,N_11265,N_11633);
and U12518 (N_12518,N_11790,N_11883);
nand U12519 (N_12519,N_11324,N_11191);
or U12520 (N_12520,N_11445,N_11229);
xnor U12521 (N_12521,N_11072,N_11340);
nor U12522 (N_12522,N_11601,N_11682);
nor U12523 (N_12523,N_11309,N_11589);
nand U12524 (N_12524,N_11106,N_11666);
xor U12525 (N_12525,N_11688,N_11885);
or U12526 (N_12526,N_11024,N_11369);
or U12527 (N_12527,N_11145,N_11139);
xnor U12528 (N_12528,N_11257,N_11954);
or U12529 (N_12529,N_11886,N_11400);
nor U12530 (N_12530,N_11980,N_11049);
nor U12531 (N_12531,N_11529,N_11866);
and U12532 (N_12532,N_11868,N_11635);
nor U12533 (N_12533,N_11031,N_11147);
nor U12534 (N_12534,N_11067,N_11131);
nor U12535 (N_12535,N_11834,N_11511);
xor U12536 (N_12536,N_11801,N_11379);
nand U12537 (N_12537,N_11103,N_11299);
nor U12538 (N_12538,N_11485,N_11246);
or U12539 (N_12539,N_11777,N_11672);
xnor U12540 (N_12540,N_11866,N_11506);
and U12541 (N_12541,N_11075,N_11770);
xor U12542 (N_12542,N_11565,N_11059);
or U12543 (N_12543,N_11335,N_11048);
and U12544 (N_12544,N_11237,N_11581);
xnor U12545 (N_12545,N_11815,N_11549);
nor U12546 (N_12546,N_11312,N_11968);
or U12547 (N_12547,N_11012,N_11832);
or U12548 (N_12548,N_11789,N_11095);
nand U12549 (N_12549,N_11917,N_11254);
xor U12550 (N_12550,N_11479,N_11545);
nand U12551 (N_12551,N_11597,N_11851);
or U12552 (N_12552,N_11204,N_11555);
or U12553 (N_12553,N_11264,N_11879);
and U12554 (N_12554,N_11254,N_11521);
nand U12555 (N_12555,N_11864,N_11544);
nand U12556 (N_12556,N_11752,N_11697);
or U12557 (N_12557,N_11530,N_11351);
nand U12558 (N_12558,N_11949,N_11324);
nor U12559 (N_12559,N_11317,N_11672);
and U12560 (N_12560,N_11539,N_11565);
nand U12561 (N_12561,N_11911,N_11348);
nand U12562 (N_12562,N_11933,N_11177);
nor U12563 (N_12563,N_11243,N_11598);
nor U12564 (N_12564,N_11614,N_11619);
nor U12565 (N_12565,N_11631,N_11955);
nor U12566 (N_12566,N_11122,N_11245);
and U12567 (N_12567,N_11335,N_11175);
and U12568 (N_12568,N_11255,N_11482);
or U12569 (N_12569,N_11887,N_11306);
nor U12570 (N_12570,N_11467,N_11366);
xor U12571 (N_12571,N_11494,N_11149);
and U12572 (N_12572,N_11342,N_11363);
and U12573 (N_12573,N_11708,N_11539);
nor U12574 (N_12574,N_11338,N_11807);
nor U12575 (N_12575,N_11133,N_11813);
or U12576 (N_12576,N_11557,N_11735);
nor U12577 (N_12577,N_11001,N_11675);
nor U12578 (N_12578,N_11953,N_11902);
and U12579 (N_12579,N_11019,N_11784);
nand U12580 (N_12580,N_11268,N_11703);
and U12581 (N_12581,N_11352,N_11774);
xnor U12582 (N_12582,N_11032,N_11606);
and U12583 (N_12583,N_11161,N_11460);
xnor U12584 (N_12584,N_11927,N_11411);
nor U12585 (N_12585,N_11116,N_11400);
and U12586 (N_12586,N_11581,N_11871);
xnor U12587 (N_12587,N_11854,N_11024);
or U12588 (N_12588,N_11998,N_11232);
xor U12589 (N_12589,N_11689,N_11532);
nand U12590 (N_12590,N_11005,N_11505);
or U12591 (N_12591,N_11637,N_11718);
and U12592 (N_12592,N_11264,N_11582);
nand U12593 (N_12593,N_11223,N_11077);
nor U12594 (N_12594,N_11613,N_11181);
and U12595 (N_12595,N_11705,N_11472);
and U12596 (N_12596,N_11577,N_11010);
nor U12597 (N_12597,N_11606,N_11903);
or U12598 (N_12598,N_11639,N_11245);
nor U12599 (N_12599,N_11327,N_11767);
nand U12600 (N_12600,N_11997,N_11477);
xnor U12601 (N_12601,N_11817,N_11561);
nand U12602 (N_12602,N_11166,N_11373);
nor U12603 (N_12603,N_11318,N_11378);
and U12604 (N_12604,N_11895,N_11146);
and U12605 (N_12605,N_11810,N_11300);
or U12606 (N_12606,N_11305,N_11286);
nand U12607 (N_12607,N_11929,N_11369);
nand U12608 (N_12608,N_11384,N_11725);
nand U12609 (N_12609,N_11862,N_11773);
nand U12610 (N_12610,N_11363,N_11538);
nor U12611 (N_12611,N_11107,N_11430);
nor U12612 (N_12612,N_11346,N_11574);
xnor U12613 (N_12613,N_11588,N_11415);
or U12614 (N_12614,N_11507,N_11982);
or U12615 (N_12615,N_11115,N_11307);
or U12616 (N_12616,N_11986,N_11792);
nand U12617 (N_12617,N_11110,N_11634);
nand U12618 (N_12618,N_11652,N_11766);
nand U12619 (N_12619,N_11532,N_11399);
or U12620 (N_12620,N_11840,N_11850);
xor U12621 (N_12621,N_11861,N_11654);
xor U12622 (N_12622,N_11533,N_11806);
nor U12623 (N_12623,N_11168,N_11966);
xor U12624 (N_12624,N_11091,N_11542);
nand U12625 (N_12625,N_11855,N_11736);
and U12626 (N_12626,N_11261,N_11963);
or U12627 (N_12627,N_11749,N_11972);
and U12628 (N_12628,N_11106,N_11366);
and U12629 (N_12629,N_11830,N_11427);
or U12630 (N_12630,N_11293,N_11506);
nor U12631 (N_12631,N_11104,N_11656);
nor U12632 (N_12632,N_11414,N_11959);
xnor U12633 (N_12633,N_11375,N_11916);
xnor U12634 (N_12634,N_11869,N_11060);
nand U12635 (N_12635,N_11995,N_11799);
nand U12636 (N_12636,N_11195,N_11086);
and U12637 (N_12637,N_11554,N_11584);
xor U12638 (N_12638,N_11601,N_11481);
or U12639 (N_12639,N_11668,N_11897);
or U12640 (N_12640,N_11721,N_11816);
nor U12641 (N_12641,N_11218,N_11786);
or U12642 (N_12642,N_11130,N_11226);
nand U12643 (N_12643,N_11250,N_11393);
and U12644 (N_12644,N_11574,N_11303);
and U12645 (N_12645,N_11704,N_11304);
nor U12646 (N_12646,N_11983,N_11087);
and U12647 (N_12647,N_11690,N_11603);
and U12648 (N_12648,N_11837,N_11757);
or U12649 (N_12649,N_11849,N_11626);
nor U12650 (N_12650,N_11867,N_11627);
nor U12651 (N_12651,N_11935,N_11394);
nor U12652 (N_12652,N_11745,N_11039);
and U12653 (N_12653,N_11346,N_11456);
nand U12654 (N_12654,N_11079,N_11268);
xnor U12655 (N_12655,N_11275,N_11184);
nor U12656 (N_12656,N_11972,N_11751);
nand U12657 (N_12657,N_11540,N_11590);
xor U12658 (N_12658,N_11075,N_11164);
or U12659 (N_12659,N_11941,N_11284);
nor U12660 (N_12660,N_11516,N_11889);
and U12661 (N_12661,N_11925,N_11089);
or U12662 (N_12662,N_11124,N_11563);
nand U12663 (N_12663,N_11282,N_11918);
or U12664 (N_12664,N_11610,N_11055);
and U12665 (N_12665,N_11293,N_11519);
xor U12666 (N_12666,N_11855,N_11829);
and U12667 (N_12667,N_11409,N_11765);
and U12668 (N_12668,N_11074,N_11449);
and U12669 (N_12669,N_11105,N_11186);
nor U12670 (N_12670,N_11405,N_11091);
or U12671 (N_12671,N_11562,N_11853);
or U12672 (N_12672,N_11707,N_11406);
nor U12673 (N_12673,N_11199,N_11460);
and U12674 (N_12674,N_11502,N_11717);
nor U12675 (N_12675,N_11661,N_11009);
xnor U12676 (N_12676,N_11052,N_11367);
xnor U12677 (N_12677,N_11365,N_11177);
or U12678 (N_12678,N_11366,N_11880);
xor U12679 (N_12679,N_11020,N_11790);
xnor U12680 (N_12680,N_11419,N_11157);
or U12681 (N_12681,N_11106,N_11023);
xor U12682 (N_12682,N_11404,N_11550);
and U12683 (N_12683,N_11329,N_11357);
or U12684 (N_12684,N_11807,N_11872);
or U12685 (N_12685,N_11466,N_11214);
xor U12686 (N_12686,N_11922,N_11582);
and U12687 (N_12687,N_11879,N_11906);
and U12688 (N_12688,N_11113,N_11372);
nor U12689 (N_12689,N_11149,N_11095);
and U12690 (N_12690,N_11682,N_11203);
nor U12691 (N_12691,N_11743,N_11689);
and U12692 (N_12692,N_11305,N_11333);
or U12693 (N_12693,N_11048,N_11318);
nand U12694 (N_12694,N_11761,N_11701);
nor U12695 (N_12695,N_11041,N_11707);
nor U12696 (N_12696,N_11699,N_11398);
nand U12697 (N_12697,N_11461,N_11498);
and U12698 (N_12698,N_11215,N_11162);
xnor U12699 (N_12699,N_11985,N_11537);
nand U12700 (N_12700,N_11118,N_11494);
or U12701 (N_12701,N_11691,N_11084);
or U12702 (N_12702,N_11843,N_11531);
or U12703 (N_12703,N_11958,N_11294);
nor U12704 (N_12704,N_11692,N_11381);
xor U12705 (N_12705,N_11458,N_11066);
and U12706 (N_12706,N_11278,N_11438);
nor U12707 (N_12707,N_11317,N_11015);
and U12708 (N_12708,N_11573,N_11795);
xor U12709 (N_12709,N_11059,N_11053);
or U12710 (N_12710,N_11900,N_11822);
or U12711 (N_12711,N_11906,N_11244);
xor U12712 (N_12712,N_11580,N_11975);
or U12713 (N_12713,N_11269,N_11031);
or U12714 (N_12714,N_11661,N_11404);
nor U12715 (N_12715,N_11835,N_11588);
and U12716 (N_12716,N_11587,N_11241);
and U12717 (N_12717,N_11567,N_11862);
nand U12718 (N_12718,N_11479,N_11162);
and U12719 (N_12719,N_11368,N_11178);
nor U12720 (N_12720,N_11339,N_11102);
nor U12721 (N_12721,N_11514,N_11526);
nand U12722 (N_12722,N_11887,N_11174);
and U12723 (N_12723,N_11831,N_11896);
xor U12724 (N_12724,N_11463,N_11115);
nand U12725 (N_12725,N_11983,N_11687);
xnor U12726 (N_12726,N_11005,N_11050);
and U12727 (N_12727,N_11243,N_11621);
or U12728 (N_12728,N_11503,N_11561);
xnor U12729 (N_12729,N_11177,N_11465);
nand U12730 (N_12730,N_11977,N_11580);
nand U12731 (N_12731,N_11891,N_11763);
xor U12732 (N_12732,N_11785,N_11800);
nand U12733 (N_12733,N_11255,N_11917);
and U12734 (N_12734,N_11240,N_11162);
xnor U12735 (N_12735,N_11257,N_11609);
nor U12736 (N_12736,N_11450,N_11688);
or U12737 (N_12737,N_11805,N_11906);
nand U12738 (N_12738,N_11760,N_11869);
nor U12739 (N_12739,N_11527,N_11710);
or U12740 (N_12740,N_11485,N_11526);
nor U12741 (N_12741,N_11325,N_11006);
nand U12742 (N_12742,N_11612,N_11987);
nand U12743 (N_12743,N_11335,N_11194);
nor U12744 (N_12744,N_11817,N_11737);
xnor U12745 (N_12745,N_11480,N_11906);
nand U12746 (N_12746,N_11713,N_11877);
nor U12747 (N_12747,N_11620,N_11972);
nor U12748 (N_12748,N_11852,N_11312);
nand U12749 (N_12749,N_11230,N_11884);
or U12750 (N_12750,N_11786,N_11727);
nand U12751 (N_12751,N_11051,N_11876);
xor U12752 (N_12752,N_11666,N_11685);
xnor U12753 (N_12753,N_11340,N_11126);
xnor U12754 (N_12754,N_11094,N_11080);
nand U12755 (N_12755,N_11432,N_11349);
nor U12756 (N_12756,N_11995,N_11750);
nand U12757 (N_12757,N_11633,N_11170);
and U12758 (N_12758,N_11189,N_11426);
nor U12759 (N_12759,N_11715,N_11783);
nor U12760 (N_12760,N_11261,N_11854);
or U12761 (N_12761,N_11745,N_11672);
nor U12762 (N_12762,N_11888,N_11300);
nand U12763 (N_12763,N_11749,N_11643);
nand U12764 (N_12764,N_11616,N_11796);
xor U12765 (N_12765,N_11657,N_11115);
xnor U12766 (N_12766,N_11360,N_11212);
nand U12767 (N_12767,N_11349,N_11606);
and U12768 (N_12768,N_11705,N_11354);
xor U12769 (N_12769,N_11254,N_11111);
nand U12770 (N_12770,N_11010,N_11410);
xor U12771 (N_12771,N_11670,N_11571);
nand U12772 (N_12772,N_11017,N_11354);
nand U12773 (N_12773,N_11593,N_11800);
xnor U12774 (N_12774,N_11476,N_11481);
xnor U12775 (N_12775,N_11272,N_11117);
and U12776 (N_12776,N_11572,N_11617);
and U12777 (N_12777,N_11866,N_11685);
nand U12778 (N_12778,N_11300,N_11805);
xor U12779 (N_12779,N_11995,N_11618);
nand U12780 (N_12780,N_11594,N_11511);
xnor U12781 (N_12781,N_11060,N_11929);
nand U12782 (N_12782,N_11456,N_11886);
nor U12783 (N_12783,N_11752,N_11830);
xnor U12784 (N_12784,N_11907,N_11950);
nand U12785 (N_12785,N_11910,N_11783);
and U12786 (N_12786,N_11914,N_11126);
nand U12787 (N_12787,N_11314,N_11946);
xnor U12788 (N_12788,N_11788,N_11147);
and U12789 (N_12789,N_11705,N_11282);
and U12790 (N_12790,N_11877,N_11006);
and U12791 (N_12791,N_11719,N_11763);
nor U12792 (N_12792,N_11720,N_11397);
nor U12793 (N_12793,N_11989,N_11361);
and U12794 (N_12794,N_11085,N_11268);
or U12795 (N_12795,N_11574,N_11061);
nor U12796 (N_12796,N_11700,N_11454);
nor U12797 (N_12797,N_11886,N_11518);
or U12798 (N_12798,N_11208,N_11606);
or U12799 (N_12799,N_11421,N_11133);
nand U12800 (N_12800,N_11875,N_11437);
or U12801 (N_12801,N_11613,N_11008);
xnor U12802 (N_12802,N_11931,N_11012);
xnor U12803 (N_12803,N_11372,N_11869);
or U12804 (N_12804,N_11792,N_11674);
and U12805 (N_12805,N_11089,N_11098);
xnor U12806 (N_12806,N_11325,N_11965);
xor U12807 (N_12807,N_11259,N_11593);
xnor U12808 (N_12808,N_11504,N_11580);
xnor U12809 (N_12809,N_11038,N_11114);
nor U12810 (N_12810,N_11321,N_11728);
and U12811 (N_12811,N_11724,N_11788);
nand U12812 (N_12812,N_11894,N_11427);
nand U12813 (N_12813,N_11597,N_11367);
and U12814 (N_12814,N_11093,N_11766);
or U12815 (N_12815,N_11260,N_11750);
nand U12816 (N_12816,N_11090,N_11447);
nand U12817 (N_12817,N_11551,N_11093);
xor U12818 (N_12818,N_11210,N_11518);
nand U12819 (N_12819,N_11090,N_11084);
nand U12820 (N_12820,N_11905,N_11414);
xnor U12821 (N_12821,N_11452,N_11583);
and U12822 (N_12822,N_11065,N_11368);
and U12823 (N_12823,N_11115,N_11147);
and U12824 (N_12824,N_11855,N_11224);
or U12825 (N_12825,N_11512,N_11149);
xor U12826 (N_12826,N_11257,N_11769);
xnor U12827 (N_12827,N_11669,N_11146);
nand U12828 (N_12828,N_11002,N_11533);
nand U12829 (N_12829,N_11253,N_11168);
and U12830 (N_12830,N_11909,N_11639);
xor U12831 (N_12831,N_11899,N_11807);
nand U12832 (N_12832,N_11688,N_11072);
or U12833 (N_12833,N_11054,N_11042);
nand U12834 (N_12834,N_11626,N_11271);
xor U12835 (N_12835,N_11002,N_11994);
xor U12836 (N_12836,N_11396,N_11794);
nor U12837 (N_12837,N_11345,N_11926);
and U12838 (N_12838,N_11378,N_11791);
xnor U12839 (N_12839,N_11212,N_11512);
or U12840 (N_12840,N_11782,N_11748);
or U12841 (N_12841,N_11466,N_11908);
xor U12842 (N_12842,N_11637,N_11805);
nor U12843 (N_12843,N_11695,N_11081);
nand U12844 (N_12844,N_11531,N_11285);
nand U12845 (N_12845,N_11218,N_11899);
or U12846 (N_12846,N_11217,N_11395);
and U12847 (N_12847,N_11389,N_11483);
and U12848 (N_12848,N_11075,N_11559);
nor U12849 (N_12849,N_11395,N_11785);
nor U12850 (N_12850,N_11584,N_11294);
and U12851 (N_12851,N_11753,N_11531);
and U12852 (N_12852,N_11027,N_11155);
nand U12853 (N_12853,N_11053,N_11877);
xor U12854 (N_12854,N_11485,N_11269);
nor U12855 (N_12855,N_11226,N_11188);
xnor U12856 (N_12856,N_11124,N_11185);
and U12857 (N_12857,N_11780,N_11119);
xnor U12858 (N_12858,N_11595,N_11743);
nor U12859 (N_12859,N_11851,N_11385);
and U12860 (N_12860,N_11553,N_11644);
or U12861 (N_12861,N_11906,N_11543);
xnor U12862 (N_12862,N_11789,N_11101);
and U12863 (N_12863,N_11546,N_11879);
nand U12864 (N_12864,N_11470,N_11004);
nor U12865 (N_12865,N_11378,N_11649);
nand U12866 (N_12866,N_11997,N_11130);
or U12867 (N_12867,N_11849,N_11264);
or U12868 (N_12868,N_11863,N_11717);
nand U12869 (N_12869,N_11826,N_11303);
xnor U12870 (N_12870,N_11468,N_11700);
nand U12871 (N_12871,N_11753,N_11077);
or U12872 (N_12872,N_11802,N_11266);
xor U12873 (N_12873,N_11864,N_11769);
nor U12874 (N_12874,N_11822,N_11588);
or U12875 (N_12875,N_11908,N_11912);
nor U12876 (N_12876,N_11610,N_11646);
or U12877 (N_12877,N_11745,N_11875);
and U12878 (N_12878,N_11478,N_11705);
and U12879 (N_12879,N_11576,N_11335);
nand U12880 (N_12880,N_11806,N_11690);
nor U12881 (N_12881,N_11825,N_11666);
nand U12882 (N_12882,N_11817,N_11555);
nand U12883 (N_12883,N_11977,N_11704);
xnor U12884 (N_12884,N_11405,N_11877);
or U12885 (N_12885,N_11939,N_11969);
xor U12886 (N_12886,N_11733,N_11038);
nor U12887 (N_12887,N_11801,N_11210);
nor U12888 (N_12888,N_11132,N_11695);
or U12889 (N_12889,N_11437,N_11035);
or U12890 (N_12890,N_11827,N_11817);
or U12891 (N_12891,N_11923,N_11651);
nor U12892 (N_12892,N_11618,N_11746);
nand U12893 (N_12893,N_11154,N_11351);
nor U12894 (N_12894,N_11439,N_11536);
xnor U12895 (N_12895,N_11757,N_11571);
or U12896 (N_12896,N_11894,N_11102);
nand U12897 (N_12897,N_11740,N_11403);
or U12898 (N_12898,N_11758,N_11464);
nand U12899 (N_12899,N_11122,N_11460);
nor U12900 (N_12900,N_11519,N_11570);
and U12901 (N_12901,N_11989,N_11823);
or U12902 (N_12902,N_11272,N_11192);
or U12903 (N_12903,N_11976,N_11461);
nor U12904 (N_12904,N_11439,N_11625);
xor U12905 (N_12905,N_11024,N_11789);
xor U12906 (N_12906,N_11061,N_11850);
nand U12907 (N_12907,N_11323,N_11897);
or U12908 (N_12908,N_11502,N_11840);
or U12909 (N_12909,N_11689,N_11774);
or U12910 (N_12910,N_11959,N_11764);
nand U12911 (N_12911,N_11997,N_11598);
nor U12912 (N_12912,N_11560,N_11060);
xnor U12913 (N_12913,N_11759,N_11175);
or U12914 (N_12914,N_11968,N_11703);
nor U12915 (N_12915,N_11393,N_11981);
or U12916 (N_12916,N_11256,N_11222);
nand U12917 (N_12917,N_11522,N_11532);
or U12918 (N_12918,N_11711,N_11044);
and U12919 (N_12919,N_11706,N_11200);
xnor U12920 (N_12920,N_11901,N_11334);
nand U12921 (N_12921,N_11458,N_11881);
or U12922 (N_12922,N_11841,N_11893);
nand U12923 (N_12923,N_11858,N_11015);
nor U12924 (N_12924,N_11070,N_11601);
xnor U12925 (N_12925,N_11442,N_11781);
or U12926 (N_12926,N_11479,N_11523);
nand U12927 (N_12927,N_11611,N_11861);
or U12928 (N_12928,N_11484,N_11874);
xnor U12929 (N_12929,N_11634,N_11078);
nand U12930 (N_12930,N_11202,N_11798);
xnor U12931 (N_12931,N_11362,N_11761);
or U12932 (N_12932,N_11005,N_11691);
or U12933 (N_12933,N_11093,N_11716);
or U12934 (N_12934,N_11075,N_11954);
and U12935 (N_12935,N_11277,N_11605);
nand U12936 (N_12936,N_11778,N_11686);
and U12937 (N_12937,N_11983,N_11774);
or U12938 (N_12938,N_11606,N_11814);
and U12939 (N_12939,N_11734,N_11571);
nand U12940 (N_12940,N_11416,N_11861);
nor U12941 (N_12941,N_11003,N_11745);
and U12942 (N_12942,N_11556,N_11534);
and U12943 (N_12943,N_11382,N_11872);
or U12944 (N_12944,N_11657,N_11682);
and U12945 (N_12945,N_11810,N_11545);
or U12946 (N_12946,N_11624,N_11654);
xnor U12947 (N_12947,N_11099,N_11353);
nor U12948 (N_12948,N_11071,N_11992);
or U12949 (N_12949,N_11201,N_11913);
nor U12950 (N_12950,N_11994,N_11225);
nand U12951 (N_12951,N_11174,N_11306);
and U12952 (N_12952,N_11270,N_11829);
nand U12953 (N_12953,N_11463,N_11647);
nand U12954 (N_12954,N_11799,N_11737);
and U12955 (N_12955,N_11409,N_11262);
or U12956 (N_12956,N_11857,N_11678);
nand U12957 (N_12957,N_11944,N_11756);
and U12958 (N_12958,N_11570,N_11363);
nor U12959 (N_12959,N_11495,N_11960);
xor U12960 (N_12960,N_11047,N_11691);
xor U12961 (N_12961,N_11201,N_11119);
or U12962 (N_12962,N_11559,N_11108);
or U12963 (N_12963,N_11341,N_11912);
xnor U12964 (N_12964,N_11450,N_11009);
nor U12965 (N_12965,N_11399,N_11866);
or U12966 (N_12966,N_11112,N_11732);
nand U12967 (N_12967,N_11700,N_11851);
and U12968 (N_12968,N_11125,N_11129);
xor U12969 (N_12969,N_11862,N_11187);
nand U12970 (N_12970,N_11623,N_11293);
or U12971 (N_12971,N_11493,N_11884);
xor U12972 (N_12972,N_11679,N_11978);
nor U12973 (N_12973,N_11252,N_11265);
xor U12974 (N_12974,N_11140,N_11649);
and U12975 (N_12975,N_11291,N_11384);
and U12976 (N_12976,N_11591,N_11991);
xor U12977 (N_12977,N_11799,N_11557);
and U12978 (N_12978,N_11886,N_11138);
xor U12979 (N_12979,N_11714,N_11262);
and U12980 (N_12980,N_11099,N_11336);
or U12981 (N_12981,N_11172,N_11464);
xor U12982 (N_12982,N_11866,N_11145);
or U12983 (N_12983,N_11920,N_11034);
xnor U12984 (N_12984,N_11106,N_11754);
or U12985 (N_12985,N_11835,N_11413);
or U12986 (N_12986,N_11673,N_11056);
xnor U12987 (N_12987,N_11633,N_11151);
nor U12988 (N_12988,N_11824,N_11855);
and U12989 (N_12989,N_11675,N_11337);
and U12990 (N_12990,N_11921,N_11420);
and U12991 (N_12991,N_11304,N_11526);
nand U12992 (N_12992,N_11220,N_11491);
or U12993 (N_12993,N_11835,N_11474);
and U12994 (N_12994,N_11031,N_11059);
and U12995 (N_12995,N_11604,N_11737);
and U12996 (N_12996,N_11329,N_11015);
and U12997 (N_12997,N_11702,N_11352);
nor U12998 (N_12998,N_11042,N_11674);
nor U12999 (N_12999,N_11700,N_11046);
and U13000 (N_13000,N_12353,N_12144);
nand U13001 (N_13001,N_12078,N_12926);
xnor U13002 (N_13002,N_12503,N_12706);
and U13003 (N_13003,N_12857,N_12120);
and U13004 (N_13004,N_12343,N_12692);
xnor U13005 (N_13005,N_12345,N_12365);
and U13006 (N_13006,N_12132,N_12054);
nor U13007 (N_13007,N_12377,N_12707);
nor U13008 (N_13008,N_12143,N_12769);
xnor U13009 (N_13009,N_12510,N_12423);
nor U13010 (N_13010,N_12397,N_12033);
nor U13011 (N_13011,N_12273,N_12942);
and U13012 (N_13012,N_12504,N_12406);
or U13013 (N_13013,N_12096,N_12505);
nand U13014 (N_13014,N_12000,N_12590);
and U13015 (N_13015,N_12981,N_12572);
nand U13016 (N_13016,N_12863,N_12242);
xnor U13017 (N_13017,N_12104,N_12904);
and U13018 (N_13018,N_12410,N_12917);
nor U13019 (N_13019,N_12500,N_12815);
nand U13020 (N_13020,N_12465,N_12937);
xnor U13021 (N_13021,N_12086,N_12574);
nor U13022 (N_13022,N_12998,N_12002);
xor U13023 (N_13023,N_12085,N_12071);
or U13024 (N_13024,N_12667,N_12717);
nor U13025 (N_13025,N_12385,N_12948);
and U13026 (N_13026,N_12653,N_12809);
nor U13027 (N_13027,N_12580,N_12989);
nand U13028 (N_13028,N_12371,N_12197);
or U13029 (N_13029,N_12562,N_12065);
xnor U13030 (N_13030,N_12452,N_12180);
or U13031 (N_13031,N_12460,N_12641);
or U13032 (N_13032,N_12502,N_12128);
or U13033 (N_13033,N_12886,N_12927);
xnor U13034 (N_13034,N_12796,N_12954);
and U13035 (N_13035,N_12324,N_12646);
or U13036 (N_13036,N_12280,N_12755);
and U13037 (N_13037,N_12845,N_12015);
nor U13038 (N_13038,N_12265,N_12721);
and U13039 (N_13039,N_12779,N_12175);
and U13040 (N_13040,N_12561,N_12891);
and U13041 (N_13041,N_12093,N_12799);
nor U13042 (N_13042,N_12805,N_12330);
or U13043 (N_13043,N_12124,N_12684);
or U13044 (N_13044,N_12847,N_12759);
nand U13045 (N_13045,N_12591,N_12516);
and U13046 (N_13046,N_12340,N_12425);
nand U13047 (N_13047,N_12158,N_12295);
and U13048 (N_13048,N_12416,N_12987);
and U13049 (N_13049,N_12888,N_12127);
or U13050 (N_13050,N_12312,N_12678);
or U13051 (N_13051,N_12966,N_12457);
nor U13052 (N_13052,N_12670,N_12328);
xnor U13053 (N_13053,N_12620,N_12800);
and U13054 (N_13054,N_12971,N_12696);
and U13055 (N_13055,N_12936,N_12492);
and U13056 (N_13056,N_12911,N_12428);
nand U13057 (N_13057,N_12107,N_12355);
nand U13058 (N_13058,N_12166,N_12008);
nor U13059 (N_13059,N_12017,N_12157);
or U13060 (N_13060,N_12765,N_12476);
nand U13061 (N_13061,N_12323,N_12013);
xnor U13062 (N_13062,N_12626,N_12952);
and U13063 (N_13063,N_12066,N_12228);
and U13064 (N_13064,N_12632,N_12337);
nand U13065 (N_13065,N_12342,N_12152);
nand U13066 (N_13066,N_12209,N_12551);
nand U13067 (N_13067,N_12032,N_12790);
and U13068 (N_13068,N_12634,N_12348);
and U13069 (N_13069,N_12262,N_12094);
nand U13070 (N_13070,N_12518,N_12718);
or U13071 (N_13071,N_12732,N_12865);
or U13072 (N_13072,N_12907,N_12320);
nor U13073 (N_13073,N_12450,N_12633);
nand U13074 (N_13074,N_12169,N_12165);
and U13075 (N_13075,N_12034,N_12635);
nor U13076 (N_13076,N_12223,N_12967);
nand U13077 (N_13077,N_12434,N_12766);
xor U13078 (N_13078,N_12931,N_12376);
or U13079 (N_13079,N_12184,N_12662);
xnor U13080 (N_13080,N_12637,N_12254);
nand U13081 (N_13081,N_12945,N_12139);
and U13082 (N_13082,N_12623,N_12045);
nor U13083 (N_13083,N_12758,N_12618);
and U13084 (N_13084,N_12752,N_12610);
nor U13085 (N_13085,N_12011,N_12473);
or U13086 (N_13086,N_12768,N_12609);
nand U13087 (N_13087,N_12161,N_12248);
nand U13088 (N_13088,N_12074,N_12554);
or U13089 (N_13089,N_12488,N_12813);
or U13090 (N_13090,N_12775,N_12668);
and U13091 (N_13091,N_12556,N_12229);
nand U13092 (N_13092,N_12527,N_12309);
nand U13093 (N_13093,N_12714,N_12407);
or U13094 (N_13094,N_12982,N_12743);
nor U13095 (N_13095,N_12628,N_12780);
or U13096 (N_13096,N_12621,N_12046);
xor U13097 (N_13097,N_12056,N_12053);
xnor U13098 (N_13098,N_12921,N_12463);
xor U13099 (N_13099,N_12833,N_12199);
or U13100 (N_13100,N_12928,N_12964);
xnor U13101 (N_13101,N_12261,N_12501);
nor U13102 (N_13102,N_12613,N_12403);
xor U13103 (N_13103,N_12177,N_12876);
or U13104 (N_13104,N_12461,N_12807);
or U13105 (N_13105,N_12963,N_12855);
or U13106 (N_13106,N_12910,N_12319);
xnor U13107 (N_13107,N_12399,N_12351);
xor U13108 (N_13108,N_12702,N_12358);
or U13109 (N_13109,N_12676,N_12680);
nor U13110 (N_13110,N_12108,N_12988);
nand U13111 (N_13111,N_12977,N_12185);
and U13112 (N_13112,N_12213,N_12063);
nand U13113 (N_13113,N_12350,N_12880);
nor U13114 (N_13114,N_12025,N_12822);
nor U13115 (N_13115,N_12617,N_12658);
xor U13116 (N_13116,N_12255,N_12899);
or U13117 (N_13117,N_12485,N_12830);
and U13118 (N_13118,N_12630,N_12316);
nor U13119 (N_13119,N_12691,N_12673);
nand U13120 (N_13120,N_12850,N_12567);
xnor U13121 (N_13121,N_12302,N_12204);
and U13122 (N_13122,N_12436,N_12163);
nand U13123 (N_13123,N_12705,N_12872);
nor U13124 (N_13124,N_12479,N_12352);
or U13125 (N_13125,N_12234,N_12136);
xnor U13126 (N_13126,N_12601,N_12624);
xnor U13127 (N_13127,N_12887,N_12266);
xnor U13128 (N_13128,N_12250,N_12918);
nand U13129 (N_13129,N_12782,N_12125);
and U13130 (N_13130,N_12315,N_12398);
or U13131 (N_13131,N_12467,N_12729);
nand U13132 (N_13132,N_12441,N_12150);
nor U13133 (N_13133,N_12097,N_12194);
nand U13134 (N_13134,N_12995,N_12512);
and U13135 (N_13135,N_12602,N_12604);
and U13136 (N_13136,N_12730,N_12260);
and U13137 (N_13137,N_12867,N_12726);
xnor U13138 (N_13138,N_12683,N_12770);
xor U13139 (N_13139,N_12313,N_12837);
nor U13140 (N_13140,N_12497,N_12258);
xnor U13141 (N_13141,N_12949,N_12905);
or U13142 (N_13142,N_12924,N_12072);
or U13143 (N_13143,N_12061,N_12080);
nor U13144 (N_13144,N_12115,N_12146);
and U13145 (N_13145,N_12135,N_12508);
nand U13146 (N_13146,N_12823,N_12232);
and U13147 (N_13147,N_12294,N_12293);
nand U13148 (N_13148,N_12023,N_12838);
nor U13149 (N_13149,N_12844,N_12846);
xor U13150 (N_13150,N_12734,N_12835);
and U13151 (N_13151,N_12070,N_12012);
xnor U13152 (N_13152,N_12119,N_12737);
xnor U13153 (N_13153,N_12007,N_12305);
xor U13154 (N_13154,N_12111,N_12241);
and U13155 (N_13155,N_12019,N_12322);
or U13156 (N_13156,N_12470,N_12841);
or U13157 (N_13157,N_12221,N_12546);
and U13158 (N_13158,N_12238,N_12908);
or U13159 (N_13159,N_12049,N_12958);
xnor U13160 (N_13160,N_12525,N_12672);
xnor U13161 (N_13161,N_12271,N_12171);
or U13162 (N_13162,N_12912,N_12215);
nand U13163 (N_13163,N_12110,N_12363);
and U13164 (N_13164,N_12716,N_12748);
or U13165 (N_13165,N_12349,N_12099);
xnor U13166 (N_13166,N_12311,N_12898);
and U13167 (N_13167,N_12777,N_12036);
nand U13168 (N_13168,N_12244,N_12875);
and U13169 (N_13169,N_12840,N_12188);
or U13170 (N_13170,N_12474,N_12181);
and U13171 (N_13171,N_12515,N_12206);
and U13172 (N_13172,N_12130,N_12060);
and U13173 (N_13173,N_12774,N_12665);
and U13174 (N_13174,N_12993,N_12587);
nand U13175 (N_13175,N_12881,N_12659);
xor U13176 (N_13176,N_12751,N_12715);
or U13177 (N_13177,N_12861,N_12024);
nand U13178 (N_13178,N_12442,N_12892);
and U13179 (N_13179,N_12938,N_12573);
nand U13180 (N_13180,N_12731,N_12786);
nor U13181 (N_13181,N_12622,N_12552);
and U13182 (N_13182,N_12446,N_12092);
and U13183 (N_13183,N_12222,N_12122);
or U13184 (N_13184,N_12784,N_12374);
nand U13185 (N_13185,N_12879,N_12109);
and U13186 (N_13186,N_12321,N_12897);
xnor U13187 (N_13187,N_12415,N_12695);
nor U13188 (N_13188,N_12419,N_12596);
nand U13189 (N_13189,N_12923,N_12230);
nand U13190 (N_13190,N_12816,N_12037);
xor U13191 (N_13191,N_12657,N_12332);
nor U13192 (N_13192,N_12694,N_12405);
and U13193 (N_13193,N_12728,N_12597);
and U13194 (N_13194,N_12693,N_12818);
xor U13195 (N_13195,N_12168,N_12589);
nand U13196 (N_13196,N_12660,N_12583);
nand U13197 (N_13197,N_12429,N_12381);
nand U13198 (N_13198,N_12042,N_12020);
nor U13199 (N_13199,N_12384,N_12089);
and U13200 (N_13200,N_12961,N_12114);
and U13201 (N_13201,N_12953,N_12156);
and U13202 (N_13202,N_12486,N_12129);
and U13203 (N_13203,N_12878,N_12920);
xor U13204 (N_13204,N_12028,N_12549);
xor U13205 (N_13205,N_12532,N_12448);
nor U13206 (N_13206,N_12956,N_12133);
xnor U13207 (N_13207,N_12514,N_12484);
xnor U13208 (N_13208,N_12664,N_12040);
xnor U13209 (N_13209,N_12690,N_12939);
xor U13210 (N_13210,N_12076,N_12101);
and U13211 (N_13211,N_12742,N_12297);
and U13212 (N_13212,N_12877,N_12394);
xor U13213 (N_13213,N_12588,N_12559);
or U13214 (N_13214,N_12675,N_12654);
or U13215 (N_13215,N_12016,N_12048);
and U13216 (N_13216,N_12550,N_12490);
nand U13217 (N_13217,N_12477,N_12946);
nand U13218 (N_13218,N_12383,N_12885);
nor U13219 (N_13219,N_12827,N_12159);
nor U13220 (N_13220,N_12491,N_12439);
or U13221 (N_13221,N_12579,N_12083);
nor U13222 (N_13222,N_12778,N_12018);
nand U13223 (N_13223,N_12824,N_12247);
nor U13224 (N_13224,N_12370,N_12999);
and U13225 (N_13225,N_12493,N_12825);
or U13226 (N_13226,N_12334,N_12974);
nand U13227 (N_13227,N_12489,N_12560);
xor U13228 (N_13228,N_12750,N_12521);
or U13229 (N_13229,N_12747,N_12997);
or U13230 (N_13230,N_12585,N_12256);
or U13231 (N_13231,N_12192,N_12544);
nor U13232 (N_13232,N_12299,N_12014);
and U13233 (N_13233,N_12102,N_12226);
xor U13234 (N_13234,N_12186,N_12272);
and U13235 (N_13235,N_12711,N_12581);
or U13236 (N_13236,N_12317,N_12113);
nor U13237 (N_13237,N_12137,N_12090);
nor U13238 (N_13238,N_12239,N_12703);
xnor U13239 (N_13239,N_12052,N_12699);
nand U13240 (N_13240,N_12389,N_12059);
nand U13241 (N_13241,N_12178,N_12772);
and U13242 (N_13242,N_12227,N_12520);
nor U13243 (N_13243,N_12839,N_12496);
nor U13244 (N_13244,N_12445,N_12906);
nor U13245 (N_13245,N_12739,N_12160);
nand U13246 (N_13246,N_12536,N_12277);
or U13247 (N_13247,N_12432,N_12073);
and U13248 (N_13248,N_12438,N_12400);
nand U13249 (N_13249,N_12220,N_12393);
and U13250 (N_13250,N_12117,N_12252);
or U13251 (N_13251,N_12047,N_12055);
and U13252 (N_13252,N_12978,N_12331);
or U13253 (N_13253,N_12529,N_12116);
and U13254 (N_13254,N_12860,N_12466);
nand U13255 (N_13255,N_12831,N_12785);
and U13256 (N_13256,N_12142,N_12645);
or U13257 (N_13257,N_12724,N_12494);
nand U13258 (N_13258,N_12903,N_12735);
and U13259 (N_13259,N_12788,N_12627);
nand U13260 (N_13260,N_12578,N_12557);
nand U13261 (N_13261,N_12575,N_12754);
nand U13262 (N_13262,N_12563,N_12341);
or U13263 (N_13263,N_12338,N_12611);
nor U13264 (N_13264,N_12141,N_12456);
xnor U13265 (N_13265,N_12329,N_12968);
and U13266 (N_13266,N_12929,N_12854);
xnor U13267 (N_13267,N_12368,N_12021);
xor U13268 (N_13268,N_12592,N_12095);
nor U13269 (N_13269,N_12803,N_12426);
nand U13270 (N_13270,N_12354,N_12362);
nor U13271 (N_13271,N_12858,N_12131);
nor U13272 (N_13272,N_12487,N_12864);
xnor U13273 (N_13273,N_12203,N_12198);
or U13274 (N_13274,N_12994,N_12041);
and U13275 (N_13275,N_12868,N_12638);
and U13276 (N_13276,N_12303,N_12733);
and U13277 (N_13277,N_12246,N_12566);
and U13278 (N_13278,N_12039,N_12663);
or U13279 (N_13279,N_12652,N_12523);
nand U13280 (N_13280,N_12240,N_12914);
xnor U13281 (N_13281,N_12372,N_12539);
and U13282 (N_13282,N_12586,N_12084);
nor U13283 (N_13283,N_12571,N_12069);
or U13284 (N_13284,N_12593,N_12607);
nor U13285 (N_13285,N_12509,N_12424);
nand U13286 (N_13286,N_12314,N_12214);
nor U13287 (N_13287,N_12797,N_12565);
nor U13288 (N_13288,N_12615,N_12972);
nand U13289 (N_13289,N_12577,N_12951);
and U13290 (N_13290,N_12873,N_12375);
nor U13291 (N_13291,N_12026,N_12806);
nor U13292 (N_13292,N_12511,N_12112);
or U13293 (N_13293,N_12746,N_12736);
nand U13294 (N_13294,N_12555,N_12741);
xnor U13295 (N_13295,N_12333,N_12915);
nand U13296 (N_13296,N_12882,N_12225);
nor U13297 (N_13297,N_12005,N_12421);
and U13298 (N_13298,N_12216,N_12401);
nand U13299 (N_13299,N_12412,N_12934);
and U13300 (N_13300,N_12464,N_12991);
nor U13301 (N_13301,N_12106,N_12173);
nor U13302 (N_13302,N_12155,N_12409);
nand U13303 (N_13303,N_12212,N_12792);
nor U13304 (N_13304,N_12541,N_12866);
and U13305 (N_13305,N_12883,N_12264);
or U13306 (N_13306,N_12965,N_12304);
nand U13307 (N_13307,N_12677,N_12245);
nand U13308 (N_13308,N_12568,N_12195);
nand U13309 (N_13309,N_12207,N_12079);
nor U13310 (N_13310,N_12826,N_12361);
or U13311 (N_13311,N_12697,N_12674);
xor U13312 (N_13312,N_12679,N_12817);
and U13313 (N_13313,N_12513,N_12656);
and U13314 (N_13314,N_12408,N_12373);
and U13315 (N_13315,N_12543,N_12640);
nor U13316 (N_13316,N_12001,N_12196);
and U13317 (N_13317,N_12614,N_12764);
xnor U13318 (N_13318,N_12189,N_12360);
and U13319 (N_13319,N_12386,N_12859);
and U13320 (N_13320,N_12829,N_12336);
xnor U13321 (N_13321,N_12075,N_12745);
or U13322 (N_13322,N_12979,N_12138);
and U13323 (N_13323,N_12689,N_12417);
or U13324 (N_13324,N_12451,N_12950);
or U13325 (N_13325,N_12498,N_12856);
nor U13326 (N_13326,N_12832,N_12802);
xnor U13327 (N_13327,N_12279,N_12848);
and U13328 (N_13328,N_12027,N_12183);
nand U13329 (N_13329,N_12267,N_12233);
xnor U13330 (N_13330,N_12996,N_12444);
and U13331 (N_13331,N_12851,N_12576);
and U13332 (N_13332,N_12288,N_12287);
nand U13333 (N_13333,N_12147,N_12725);
nor U13334 (N_13334,N_12202,N_12275);
xor U13335 (N_13335,N_12347,N_12356);
xor U13336 (N_13336,N_12268,N_12955);
nand U13337 (N_13337,N_12308,N_12584);
nand U13338 (N_13338,N_12973,N_12148);
nand U13339 (N_13339,N_12922,N_12170);
nor U13340 (N_13340,N_12776,N_12537);
nor U13341 (N_13341,N_12595,N_12925);
nand U13342 (N_13342,N_12648,N_12631);
nor U13343 (N_13343,N_12594,N_12700);
or U13344 (N_13344,N_12517,N_12547);
and U13345 (N_13345,N_12990,N_12357);
xnor U13346 (N_13346,N_12980,N_12843);
nor U13347 (N_13347,N_12793,N_12378);
nand U13348 (N_13348,N_12335,N_12030);
xor U13349 (N_13349,N_12327,N_12895);
nand U13350 (N_13350,N_12771,N_12688);
and U13351 (N_13351,N_12871,N_12387);
or U13352 (N_13352,N_12528,N_12043);
and U13353 (N_13353,N_12003,N_12454);
or U13354 (N_13354,N_12339,N_12281);
or U13355 (N_13355,N_12187,N_12193);
xnor U13356 (N_13356,N_12612,N_12081);
nor U13357 (N_13357,N_12682,N_12420);
nand U13358 (N_13358,N_12068,N_12453);
xnor U13359 (N_13359,N_12636,N_12263);
nand U13360 (N_13360,N_12392,N_12449);
nor U13361 (N_13361,N_12763,N_12306);
xor U13362 (N_13362,N_12787,N_12808);
and U13363 (N_13363,N_12603,N_12217);
nand U13364 (N_13364,N_12647,N_12270);
nand U13365 (N_13365,N_12091,N_12251);
xnor U13366 (N_13366,N_12440,N_12538);
xnor U13367 (N_13367,N_12179,N_12300);
xor U13368 (N_13368,N_12298,N_12274);
or U13369 (N_13369,N_12810,N_12478);
nand U13370 (N_13370,N_12849,N_12190);
and U13371 (N_13371,N_12499,N_12598);
and U13372 (N_13372,N_12526,N_12224);
and U13373 (N_13373,N_12642,N_12545);
nand U13374 (N_13374,N_12744,N_12902);
and U13375 (N_13375,N_12391,N_12738);
nand U13376 (N_13376,N_12804,N_12757);
nand U13377 (N_13377,N_12103,N_12082);
and U13378 (N_13378,N_12767,N_12390);
or U13379 (N_13379,N_12218,N_12960);
and U13380 (N_13380,N_12639,N_12852);
or U13381 (N_13381,N_12346,N_12459);
and U13382 (N_13382,N_12121,N_12781);
nor U13383 (N_13383,N_12483,N_12427);
nor U13384 (N_13384,N_12167,N_12307);
and U13385 (N_13385,N_12794,N_12282);
and U13386 (N_13386,N_12686,N_12957);
nand U13387 (N_13387,N_12983,N_12798);
nor U13388 (N_13388,N_12862,N_12482);
and U13389 (N_13389,N_12643,N_12976);
or U13390 (N_13390,N_12944,N_12380);
and U13391 (N_13391,N_12708,N_12471);
or U13392 (N_13392,N_12285,N_12710);
and U13393 (N_13393,N_12153,N_12773);
nand U13394 (N_13394,N_12208,N_12118);
nand U13395 (N_13395,N_12932,N_12257);
nor U13396 (N_13396,N_12462,N_12723);
nor U13397 (N_13397,N_12430,N_12940);
nand U13398 (N_13398,N_12388,N_12475);
xnor U13399 (N_13399,N_12722,N_12962);
nor U13400 (N_13400,N_12836,N_12524);
or U13401 (N_13401,N_12100,N_12644);
nor U13402 (N_13402,N_12890,N_12975);
nand U13403 (N_13403,N_12098,N_12051);
nor U13404 (N_13404,N_12900,N_12164);
nand U13405 (N_13405,N_12004,N_12364);
or U13406 (N_13406,N_12749,N_12874);
xor U13407 (N_13407,N_12236,N_12687);
nor U13408 (N_13408,N_12970,N_12869);
xor U13409 (N_13409,N_12801,N_12548);
or U13410 (N_13410,N_12182,N_12359);
or U13411 (N_13411,N_12259,N_12010);
nor U13412 (N_13412,N_12088,N_12468);
xnor U13413 (N_13413,N_12713,N_12819);
or U13414 (N_13414,N_12472,N_12600);
nand U13415 (N_13415,N_12172,N_12941);
xnor U13416 (N_13416,N_12029,N_12211);
or U13417 (N_13417,N_12756,N_12753);
xnor U13418 (N_13418,N_12326,N_12290);
or U13419 (N_13419,N_12443,N_12050);
nand U13420 (N_13420,N_12174,N_12795);
xnor U13421 (N_13421,N_12145,N_12535);
nand U13422 (N_13422,N_12284,N_12413);
nand U13423 (N_13423,N_12210,N_12649);
and U13424 (N_13424,N_12783,N_12134);
nor U13425 (N_13425,N_12828,N_12901);
nand U13426 (N_13426,N_12893,N_12414);
nand U13427 (N_13427,N_12985,N_12812);
nand U13428 (N_13428,N_12035,N_12447);
and U13429 (N_13429,N_12553,N_12530);
xnor U13430 (N_13430,N_12959,N_12276);
nor U13431 (N_13431,N_12651,N_12231);
and U13432 (N_13432,N_12655,N_12986);
nand U13433 (N_13433,N_12616,N_12123);
nand U13434 (N_13434,N_12943,N_12205);
xor U13435 (N_13435,N_12286,N_12433);
xor U13436 (N_13436,N_12191,N_12671);
xor U13437 (N_13437,N_12495,N_12067);
xnor U13438 (N_13438,N_12044,N_12564);
xnor U13439 (N_13439,N_12947,N_12704);
and U13440 (N_13440,N_12269,N_12992);
and U13441 (N_13441,N_12278,N_12542);
xor U13442 (N_13442,N_12369,N_12919);
and U13443 (N_13443,N_12522,N_12606);
nor U13444 (N_13444,N_12009,N_12570);
nor U13445 (N_13445,N_12969,N_12006);
xor U13446 (N_13446,N_12064,N_12396);
and U13447 (N_13447,N_12154,N_12253);
or U13448 (N_13448,N_12712,N_12762);
and U13449 (N_13449,N_12894,N_12814);
or U13450 (N_13450,N_12292,N_12431);
nand U13451 (N_13451,N_12740,N_12719);
xnor U13452 (N_13452,N_12811,N_12435);
and U13453 (N_13453,N_12935,N_12455);
nor U13454 (N_13454,N_12519,N_12650);
or U13455 (N_13455,N_12243,N_12507);
and U13456 (N_13456,N_12219,N_12404);
nor U13457 (N_13457,N_12289,N_12201);
or U13458 (N_13458,N_12418,N_12367);
nand U13459 (N_13459,N_12062,N_12720);
and U13460 (N_13460,N_12625,N_12291);
nand U13461 (N_13461,N_12318,N_12698);
xor U13462 (N_13462,N_12140,N_12126);
and U13463 (N_13463,N_12296,N_12853);
and U13464 (N_13464,N_12534,N_12382);
nand U13465 (N_13465,N_12151,N_12681);
xnor U13466 (N_13466,N_12301,N_12031);
nand U13467 (N_13467,N_12870,N_12411);
nor U13468 (N_13468,N_12889,N_12569);
nor U13469 (N_13469,N_12791,N_12933);
nor U13470 (N_13470,N_12896,N_12629);
or U13471 (N_13471,N_12402,N_12761);
and U13472 (N_13472,N_12176,N_12760);
or U13473 (N_13473,N_12087,N_12379);
nand U13474 (N_13474,N_12310,N_12661);
or U13475 (N_13475,N_12984,N_12058);
and U13476 (N_13476,N_12249,N_12437);
xor U13477 (N_13477,N_12149,N_12237);
or U13478 (N_13478,N_12325,N_12685);
nor U13479 (N_13479,N_12506,N_12105);
or U13480 (N_13480,N_12727,N_12619);
nand U13481 (N_13481,N_12666,N_12842);
or U13482 (N_13482,N_12235,N_12038);
xnor U13483 (N_13483,N_12709,N_12669);
xor U13484 (N_13484,N_12884,N_12200);
nor U13485 (N_13485,N_12469,N_12701);
xor U13486 (N_13486,N_12599,N_12422);
xnor U13487 (N_13487,N_12480,N_12608);
nand U13488 (N_13488,N_12540,N_12481);
or U13489 (N_13489,N_12834,N_12458);
nand U13490 (N_13490,N_12820,N_12913);
nand U13491 (N_13491,N_12531,N_12077);
and U13492 (N_13492,N_12395,N_12366);
or U13493 (N_13493,N_12344,N_12916);
xnor U13494 (N_13494,N_12821,N_12789);
and U13495 (N_13495,N_12533,N_12283);
nor U13496 (N_13496,N_12022,N_12930);
nor U13497 (N_13497,N_12909,N_12057);
xnor U13498 (N_13498,N_12605,N_12582);
xnor U13499 (N_13499,N_12162,N_12558);
and U13500 (N_13500,N_12722,N_12559);
nand U13501 (N_13501,N_12426,N_12933);
xnor U13502 (N_13502,N_12672,N_12928);
and U13503 (N_13503,N_12401,N_12208);
nand U13504 (N_13504,N_12493,N_12697);
nor U13505 (N_13505,N_12033,N_12461);
nor U13506 (N_13506,N_12326,N_12039);
nand U13507 (N_13507,N_12499,N_12049);
and U13508 (N_13508,N_12120,N_12286);
and U13509 (N_13509,N_12341,N_12848);
and U13510 (N_13510,N_12749,N_12177);
or U13511 (N_13511,N_12421,N_12987);
xnor U13512 (N_13512,N_12323,N_12365);
xor U13513 (N_13513,N_12915,N_12448);
nand U13514 (N_13514,N_12500,N_12111);
or U13515 (N_13515,N_12878,N_12195);
nor U13516 (N_13516,N_12303,N_12669);
nor U13517 (N_13517,N_12705,N_12319);
or U13518 (N_13518,N_12737,N_12135);
or U13519 (N_13519,N_12704,N_12414);
and U13520 (N_13520,N_12515,N_12234);
nand U13521 (N_13521,N_12833,N_12665);
nand U13522 (N_13522,N_12195,N_12826);
or U13523 (N_13523,N_12555,N_12804);
nand U13524 (N_13524,N_12261,N_12234);
and U13525 (N_13525,N_12034,N_12888);
nor U13526 (N_13526,N_12580,N_12915);
nor U13527 (N_13527,N_12520,N_12385);
and U13528 (N_13528,N_12628,N_12900);
nor U13529 (N_13529,N_12357,N_12795);
or U13530 (N_13530,N_12606,N_12640);
nor U13531 (N_13531,N_12440,N_12340);
nand U13532 (N_13532,N_12861,N_12723);
nand U13533 (N_13533,N_12058,N_12288);
nor U13534 (N_13534,N_12805,N_12785);
or U13535 (N_13535,N_12356,N_12673);
nor U13536 (N_13536,N_12572,N_12475);
or U13537 (N_13537,N_12473,N_12098);
and U13538 (N_13538,N_12639,N_12410);
xor U13539 (N_13539,N_12491,N_12076);
xnor U13540 (N_13540,N_12256,N_12388);
xnor U13541 (N_13541,N_12827,N_12618);
xor U13542 (N_13542,N_12131,N_12309);
nand U13543 (N_13543,N_12429,N_12849);
and U13544 (N_13544,N_12491,N_12907);
nor U13545 (N_13545,N_12532,N_12484);
xnor U13546 (N_13546,N_12069,N_12683);
nand U13547 (N_13547,N_12441,N_12602);
nor U13548 (N_13548,N_12677,N_12734);
or U13549 (N_13549,N_12767,N_12332);
and U13550 (N_13550,N_12402,N_12663);
or U13551 (N_13551,N_12422,N_12607);
and U13552 (N_13552,N_12455,N_12220);
nor U13553 (N_13553,N_12134,N_12543);
nor U13554 (N_13554,N_12271,N_12498);
or U13555 (N_13555,N_12261,N_12295);
nor U13556 (N_13556,N_12903,N_12365);
or U13557 (N_13557,N_12933,N_12097);
and U13558 (N_13558,N_12705,N_12478);
and U13559 (N_13559,N_12390,N_12305);
or U13560 (N_13560,N_12911,N_12001);
or U13561 (N_13561,N_12764,N_12690);
and U13562 (N_13562,N_12248,N_12323);
nor U13563 (N_13563,N_12571,N_12518);
and U13564 (N_13564,N_12842,N_12991);
xor U13565 (N_13565,N_12304,N_12078);
nand U13566 (N_13566,N_12298,N_12841);
or U13567 (N_13567,N_12272,N_12997);
xnor U13568 (N_13568,N_12873,N_12392);
or U13569 (N_13569,N_12455,N_12721);
xor U13570 (N_13570,N_12885,N_12302);
or U13571 (N_13571,N_12353,N_12593);
and U13572 (N_13572,N_12601,N_12576);
or U13573 (N_13573,N_12009,N_12913);
and U13574 (N_13574,N_12476,N_12597);
nor U13575 (N_13575,N_12939,N_12686);
xor U13576 (N_13576,N_12106,N_12269);
nand U13577 (N_13577,N_12693,N_12945);
and U13578 (N_13578,N_12953,N_12631);
or U13579 (N_13579,N_12611,N_12323);
and U13580 (N_13580,N_12940,N_12957);
xnor U13581 (N_13581,N_12049,N_12824);
xor U13582 (N_13582,N_12005,N_12712);
and U13583 (N_13583,N_12008,N_12033);
nand U13584 (N_13584,N_12967,N_12566);
and U13585 (N_13585,N_12570,N_12006);
and U13586 (N_13586,N_12781,N_12289);
and U13587 (N_13587,N_12326,N_12637);
nand U13588 (N_13588,N_12808,N_12626);
and U13589 (N_13589,N_12182,N_12869);
xnor U13590 (N_13590,N_12991,N_12637);
xnor U13591 (N_13591,N_12673,N_12172);
and U13592 (N_13592,N_12181,N_12631);
nor U13593 (N_13593,N_12841,N_12315);
xor U13594 (N_13594,N_12739,N_12497);
nand U13595 (N_13595,N_12300,N_12924);
nor U13596 (N_13596,N_12370,N_12400);
nor U13597 (N_13597,N_12783,N_12614);
nor U13598 (N_13598,N_12138,N_12422);
and U13599 (N_13599,N_12902,N_12262);
or U13600 (N_13600,N_12647,N_12355);
nand U13601 (N_13601,N_12750,N_12828);
and U13602 (N_13602,N_12919,N_12382);
nor U13603 (N_13603,N_12553,N_12811);
xor U13604 (N_13604,N_12969,N_12120);
or U13605 (N_13605,N_12347,N_12583);
or U13606 (N_13606,N_12190,N_12786);
nor U13607 (N_13607,N_12734,N_12367);
or U13608 (N_13608,N_12817,N_12851);
or U13609 (N_13609,N_12474,N_12707);
nand U13610 (N_13610,N_12801,N_12985);
or U13611 (N_13611,N_12359,N_12977);
xor U13612 (N_13612,N_12159,N_12835);
nor U13613 (N_13613,N_12124,N_12474);
nor U13614 (N_13614,N_12621,N_12848);
or U13615 (N_13615,N_12187,N_12098);
nand U13616 (N_13616,N_12642,N_12352);
nand U13617 (N_13617,N_12504,N_12147);
or U13618 (N_13618,N_12741,N_12054);
and U13619 (N_13619,N_12354,N_12766);
or U13620 (N_13620,N_12139,N_12065);
nor U13621 (N_13621,N_12641,N_12227);
nor U13622 (N_13622,N_12453,N_12827);
and U13623 (N_13623,N_12593,N_12294);
nand U13624 (N_13624,N_12486,N_12809);
nor U13625 (N_13625,N_12405,N_12416);
xnor U13626 (N_13626,N_12590,N_12562);
and U13627 (N_13627,N_12215,N_12087);
xnor U13628 (N_13628,N_12185,N_12252);
nand U13629 (N_13629,N_12896,N_12366);
nand U13630 (N_13630,N_12487,N_12557);
nor U13631 (N_13631,N_12876,N_12792);
xor U13632 (N_13632,N_12488,N_12071);
or U13633 (N_13633,N_12121,N_12735);
or U13634 (N_13634,N_12220,N_12238);
xnor U13635 (N_13635,N_12303,N_12131);
nor U13636 (N_13636,N_12950,N_12980);
nor U13637 (N_13637,N_12528,N_12143);
nand U13638 (N_13638,N_12610,N_12358);
xor U13639 (N_13639,N_12234,N_12266);
nor U13640 (N_13640,N_12468,N_12218);
xnor U13641 (N_13641,N_12166,N_12164);
xnor U13642 (N_13642,N_12046,N_12041);
nor U13643 (N_13643,N_12459,N_12327);
xor U13644 (N_13644,N_12688,N_12492);
nand U13645 (N_13645,N_12303,N_12695);
and U13646 (N_13646,N_12942,N_12327);
xnor U13647 (N_13647,N_12736,N_12560);
or U13648 (N_13648,N_12528,N_12617);
or U13649 (N_13649,N_12270,N_12710);
xor U13650 (N_13650,N_12637,N_12916);
or U13651 (N_13651,N_12679,N_12806);
nor U13652 (N_13652,N_12759,N_12002);
or U13653 (N_13653,N_12742,N_12092);
or U13654 (N_13654,N_12403,N_12180);
nand U13655 (N_13655,N_12559,N_12117);
and U13656 (N_13656,N_12107,N_12273);
nor U13657 (N_13657,N_12243,N_12338);
nor U13658 (N_13658,N_12802,N_12940);
xor U13659 (N_13659,N_12799,N_12175);
and U13660 (N_13660,N_12136,N_12406);
and U13661 (N_13661,N_12267,N_12443);
and U13662 (N_13662,N_12053,N_12554);
or U13663 (N_13663,N_12528,N_12727);
xor U13664 (N_13664,N_12418,N_12505);
xnor U13665 (N_13665,N_12476,N_12073);
nand U13666 (N_13666,N_12466,N_12442);
or U13667 (N_13667,N_12145,N_12518);
nor U13668 (N_13668,N_12171,N_12819);
or U13669 (N_13669,N_12254,N_12736);
or U13670 (N_13670,N_12154,N_12088);
or U13671 (N_13671,N_12696,N_12224);
nand U13672 (N_13672,N_12608,N_12252);
and U13673 (N_13673,N_12011,N_12384);
and U13674 (N_13674,N_12078,N_12794);
nand U13675 (N_13675,N_12122,N_12552);
nand U13676 (N_13676,N_12935,N_12650);
and U13677 (N_13677,N_12940,N_12303);
and U13678 (N_13678,N_12233,N_12973);
nor U13679 (N_13679,N_12098,N_12754);
or U13680 (N_13680,N_12450,N_12056);
nor U13681 (N_13681,N_12513,N_12708);
nor U13682 (N_13682,N_12033,N_12428);
and U13683 (N_13683,N_12196,N_12769);
xnor U13684 (N_13684,N_12329,N_12651);
and U13685 (N_13685,N_12313,N_12496);
nor U13686 (N_13686,N_12643,N_12025);
or U13687 (N_13687,N_12599,N_12795);
nor U13688 (N_13688,N_12756,N_12579);
nand U13689 (N_13689,N_12246,N_12765);
nand U13690 (N_13690,N_12708,N_12447);
nor U13691 (N_13691,N_12246,N_12263);
or U13692 (N_13692,N_12932,N_12332);
or U13693 (N_13693,N_12739,N_12533);
nand U13694 (N_13694,N_12469,N_12566);
nor U13695 (N_13695,N_12921,N_12899);
nor U13696 (N_13696,N_12530,N_12709);
xor U13697 (N_13697,N_12941,N_12195);
and U13698 (N_13698,N_12574,N_12776);
nor U13699 (N_13699,N_12151,N_12218);
nand U13700 (N_13700,N_12230,N_12407);
nand U13701 (N_13701,N_12991,N_12167);
or U13702 (N_13702,N_12022,N_12093);
nand U13703 (N_13703,N_12169,N_12482);
nor U13704 (N_13704,N_12452,N_12521);
nand U13705 (N_13705,N_12232,N_12383);
and U13706 (N_13706,N_12942,N_12152);
nand U13707 (N_13707,N_12682,N_12482);
nor U13708 (N_13708,N_12017,N_12094);
nor U13709 (N_13709,N_12755,N_12948);
nand U13710 (N_13710,N_12596,N_12318);
xor U13711 (N_13711,N_12693,N_12243);
or U13712 (N_13712,N_12138,N_12816);
xnor U13713 (N_13713,N_12665,N_12570);
or U13714 (N_13714,N_12447,N_12096);
nor U13715 (N_13715,N_12377,N_12079);
xnor U13716 (N_13716,N_12914,N_12986);
nand U13717 (N_13717,N_12180,N_12165);
nand U13718 (N_13718,N_12607,N_12133);
or U13719 (N_13719,N_12007,N_12021);
and U13720 (N_13720,N_12575,N_12830);
xor U13721 (N_13721,N_12672,N_12063);
xnor U13722 (N_13722,N_12536,N_12548);
and U13723 (N_13723,N_12122,N_12293);
xnor U13724 (N_13724,N_12787,N_12026);
or U13725 (N_13725,N_12266,N_12798);
xor U13726 (N_13726,N_12343,N_12471);
nor U13727 (N_13727,N_12558,N_12530);
xnor U13728 (N_13728,N_12477,N_12709);
and U13729 (N_13729,N_12326,N_12917);
nor U13730 (N_13730,N_12784,N_12902);
xor U13731 (N_13731,N_12700,N_12490);
nor U13732 (N_13732,N_12809,N_12620);
xnor U13733 (N_13733,N_12579,N_12663);
and U13734 (N_13734,N_12845,N_12046);
nor U13735 (N_13735,N_12837,N_12568);
and U13736 (N_13736,N_12169,N_12264);
and U13737 (N_13737,N_12524,N_12532);
xor U13738 (N_13738,N_12333,N_12475);
nor U13739 (N_13739,N_12935,N_12221);
xnor U13740 (N_13740,N_12992,N_12511);
nor U13741 (N_13741,N_12170,N_12592);
or U13742 (N_13742,N_12903,N_12943);
xnor U13743 (N_13743,N_12738,N_12670);
and U13744 (N_13744,N_12282,N_12545);
or U13745 (N_13745,N_12771,N_12726);
or U13746 (N_13746,N_12049,N_12560);
or U13747 (N_13747,N_12551,N_12403);
nor U13748 (N_13748,N_12206,N_12520);
nor U13749 (N_13749,N_12800,N_12664);
nand U13750 (N_13750,N_12856,N_12275);
xor U13751 (N_13751,N_12915,N_12068);
nor U13752 (N_13752,N_12131,N_12387);
xor U13753 (N_13753,N_12888,N_12763);
or U13754 (N_13754,N_12572,N_12416);
nor U13755 (N_13755,N_12022,N_12670);
nor U13756 (N_13756,N_12469,N_12197);
and U13757 (N_13757,N_12243,N_12119);
nor U13758 (N_13758,N_12615,N_12862);
and U13759 (N_13759,N_12091,N_12790);
nor U13760 (N_13760,N_12294,N_12612);
nand U13761 (N_13761,N_12985,N_12306);
or U13762 (N_13762,N_12096,N_12195);
nor U13763 (N_13763,N_12293,N_12955);
xnor U13764 (N_13764,N_12388,N_12712);
nor U13765 (N_13765,N_12522,N_12906);
and U13766 (N_13766,N_12254,N_12088);
xnor U13767 (N_13767,N_12820,N_12234);
and U13768 (N_13768,N_12907,N_12862);
nand U13769 (N_13769,N_12947,N_12369);
nand U13770 (N_13770,N_12719,N_12259);
nand U13771 (N_13771,N_12476,N_12344);
nand U13772 (N_13772,N_12829,N_12453);
or U13773 (N_13773,N_12036,N_12938);
or U13774 (N_13774,N_12428,N_12816);
xor U13775 (N_13775,N_12804,N_12948);
nor U13776 (N_13776,N_12827,N_12940);
nor U13777 (N_13777,N_12111,N_12844);
or U13778 (N_13778,N_12700,N_12591);
and U13779 (N_13779,N_12131,N_12946);
or U13780 (N_13780,N_12509,N_12068);
and U13781 (N_13781,N_12465,N_12157);
nor U13782 (N_13782,N_12052,N_12602);
xnor U13783 (N_13783,N_12214,N_12414);
xnor U13784 (N_13784,N_12351,N_12057);
and U13785 (N_13785,N_12440,N_12753);
nor U13786 (N_13786,N_12822,N_12616);
and U13787 (N_13787,N_12616,N_12595);
and U13788 (N_13788,N_12940,N_12666);
xor U13789 (N_13789,N_12194,N_12807);
nand U13790 (N_13790,N_12921,N_12795);
xor U13791 (N_13791,N_12855,N_12359);
xnor U13792 (N_13792,N_12109,N_12481);
nor U13793 (N_13793,N_12776,N_12174);
nor U13794 (N_13794,N_12485,N_12047);
and U13795 (N_13795,N_12003,N_12984);
nand U13796 (N_13796,N_12600,N_12028);
or U13797 (N_13797,N_12664,N_12376);
or U13798 (N_13798,N_12870,N_12093);
nand U13799 (N_13799,N_12022,N_12658);
nand U13800 (N_13800,N_12417,N_12186);
and U13801 (N_13801,N_12941,N_12512);
xor U13802 (N_13802,N_12563,N_12304);
nor U13803 (N_13803,N_12364,N_12968);
or U13804 (N_13804,N_12743,N_12968);
or U13805 (N_13805,N_12252,N_12853);
and U13806 (N_13806,N_12131,N_12455);
nand U13807 (N_13807,N_12928,N_12451);
nor U13808 (N_13808,N_12650,N_12685);
nor U13809 (N_13809,N_12985,N_12287);
and U13810 (N_13810,N_12095,N_12445);
and U13811 (N_13811,N_12217,N_12541);
xnor U13812 (N_13812,N_12641,N_12377);
or U13813 (N_13813,N_12467,N_12548);
xor U13814 (N_13814,N_12549,N_12140);
nand U13815 (N_13815,N_12090,N_12641);
nand U13816 (N_13816,N_12976,N_12292);
xor U13817 (N_13817,N_12284,N_12976);
and U13818 (N_13818,N_12557,N_12978);
xnor U13819 (N_13819,N_12175,N_12769);
and U13820 (N_13820,N_12887,N_12601);
or U13821 (N_13821,N_12641,N_12327);
nor U13822 (N_13822,N_12270,N_12097);
and U13823 (N_13823,N_12835,N_12692);
nand U13824 (N_13824,N_12035,N_12177);
and U13825 (N_13825,N_12144,N_12695);
xnor U13826 (N_13826,N_12099,N_12914);
or U13827 (N_13827,N_12207,N_12851);
nand U13828 (N_13828,N_12207,N_12708);
xor U13829 (N_13829,N_12638,N_12257);
and U13830 (N_13830,N_12318,N_12018);
or U13831 (N_13831,N_12932,N_12302);
nand U13832 (N_13832,N_12251,N_12741);
xnor U13833 (N_13833,N_12963,N_12135);
and U13834 (N_13834,N_12563,N_12530);
and U13835 (N_13835,N_12350,N_12205);
or U13836 (N_13836,N_12661,N_12471);
nor U13837 (N_13837,N_12794,N_12236);
and U13838 (N_13838,N_12230,N_12192);
or U13839 (N_13839,N_12377,N_12235);
and U13840 (N_13840,N_12374,N_12606);
nand U13841 (N_13841,N_12813,N_12477);
or U13842 (N_13842,N_12707,N_12077);
xor U13843 (N_13843,N_12591,N_12884);
xor U13844 (N_13844,N_12909,N_12029);
or U13845 (N_13845,N_12644,N_12882);
xor U13846 (N_13846,N_12861,N_12454);
nor U13847 (N_13847,N_12280,N_12935);
or U13848 (N_13848,N_12310,N_12761);
nand U13849 (N_13849,N_12384,N_12178);
and U13850 (N_13850,N_12450,N_12060);
xor U13851 (N_13851,N_12511,N_12123);
and U13852 (N_13852,N_12360,N_12726);
nand U13853 (N_13853,N_12268,N_12039);
and U13854 (N_13854,N_12802,N_12923);
nor U13855 (N_13855,N_12448,N_12598);
and U13856 (N_13856,N_12741,N_12419);
xor U13857 (N_13857,N_12028,N_12458);
or U13858 (N_13858,N_12107,N_12314);
and U13859 (N_13859,N_12380,N_12727);
nand U13860 (N_13860,N_12359,N_12847);
or U13861 (N_13861,N_12920,N_12536);
nand U13862 (N_13862,N_12303,N_12982);
nand U13863 (N_13863,N_12259,N_12701);
nand U13864 (N_13864,N_12857,N_12115);
nor U13865 (N_13865,N_12175,N_12306);
and U13866 (N_13866,N_12263,N_12311);
nand U13867 (N_13867,N_12567,N_12963);
and U13868 (N_13868,N_12361,N_12343);
xor U13869 (N_13869,N_12965,N_12990);
and U13870 (N_13870,N_12618,N_12794);
nor U13871 (N_13871,N_12522,N_12872);
and U13872 (N_13872,N_12549,N_12814);
nand U13873 (N_13873,N_12445,N_12868);
nand U13874 (N_13874,N_12437,N_12596);
xnor U13875 (N_13875,N_12382,N_12122);
nand U13876 (N_13876,N_12800,N_12763);
nand U13877 (N_13877,N_12244,N_12168);
xor U13878 (N_13878,N_12299,N_12143);
nor U13879 (N_13879,N_12187,N_12415);
nor U13880 (N_13880,N_12251,N_12567);
xnor U13881 (N_13881,N_12107,N_12394);
nand U13882 (N_13882,N_12907,N_12354);
nor U13883 (N_13883,N_12669,N_12962);
and U13884 (N_13884,N_12365,N_12375);
nand U13885 (N_13885,N_12739,N_12905);
xor U13886 (N_13886,N_12848,N_12247);
nand U13887 (N_13887,N_12833,N_12503);
nor U13888 (N_13888,N_12975,N_12629);
or U13889 (N_13889,N_12072,N_12586);
and U13890 (N_13890,N_12433,N_12876);
xor U13891 (N_13891,N_12854,N_12146);
and U13892 (N_13892,N_12731,N_12018);
nor U13893 (N_13893,N_12282,N_12479);
nor U13894 (N_13894,N_12684,N_12757);
or U13895 (N_13895,N_12686,N_12964);
xor U13896 (N_13896,N_12457,N_12630);
nor U13897 (N_13897,N_12632,N_12116);
nor U13898 (N_13898,N_12751,N_12157);
nand U13899 (N_13899,N_12593,N_12622);
nor U13900 (N_13900,N_12673,N_12638);
and U13901 (N_13901,N_12013,N_12399);
or U13902 (N_13902,N_12172,N_12277);
xnor U13903 (N_13903,N_12025,N_12725);
nor U13904 (N_13904,N_12453,N_12476);
xnor U13905 (N_13905,N_12266,N_12177);
nand U13906 (N_13906,N_12592,N_12735);
and U13907 (N_13907,N_12528,N_12374);
or U13908 (N_13908,N_12597,N_12026);
nor U13909 (N_13909,N_12339,N_12794);
and U13910 (N_13910,N_12646,N_12982);
xnor U13911 (N_13911,N_12339,N_12341);
nor U13912 (N_13912,N_12448,N_12300);
xor U13913 (N_13913,N_12693,N_12045);
and U13914 (N_13914,N_12036,N_12081);
or U13915 (N_13915,N_12984,N_12976);
or U13916 (N_13916,N_12847,N_12760);
nand U13917 (N_13917,N_12396,N_12584);
xnor U13918 (N_13918,N_12636,N_12736);
xor U13919 (N_13919,N_12061,N_12089);
xor U13920 (N_13920,N_12795,N_12306);
or U13921 (N_13921,N_12640,N_12280);
nand U13922 (N_13922,N_12097,N_12094);
nor U13923 (N_13923,N_12577,N_12310);
xnor U13924 (N_13924,N_12386,N_12424);
xnor U13925 (N_13925,N_12699,N_12894);
xnor U13926 (N_13926,N_12221,N_12733);
xnor U13927 (N_13927,N_12749,N_12020);
or U13928 (N_13928,N_12099,N_12722);
nor U13929 (N_13929,N_12356,N_12099);
xnor U13930 (N_13930,N_12088,N_12018);
nand U13931 (N_13931,N_12295,N_12548);
xor U13932 (N_13932,N_12671,N_12366);
or U13933 (N_13933,N_12430,N_12478);
nor U13934 (N_13934,N_12418,N_12055);
nor U13935 (N_13935,N_12731,N_12052);
xnor U13936 (N_13936,N_12693,N_12387);
nand U13937 (N_13937,N_12059,N_12273);
nor U13938 (N_13938,N_12439,N_12620);
nor U13939 (N_13939,N_12413,N_12838);
nor U13940 (N_13940,N_12294,N_12007);
xor U13941 (N_13941,N_12459,N_12507);
nor U13942 (N_13942,N_12458,N_12917);
and U13943 (N_13943,N_12234,N_12861);
and U13944 (N_13944,N_12768,N_12985);
nand U13945 (N_13945,N_12907,N_12521);
nor U13946 (N_13946,N_12146,N_12145);
or U13947 (N_13947,N_12832,N_12590);
or U13948 (N_13948,N_12085,N_12821);
xnor U13949 (N_13949,N_12725,N_12433);
nand U13950 (N_13950,N_12273,N_12991);
nor U13951 (N_13951,N_12489,N_12112);
xnor U13952 (N_13952,N_12139,N_12828);
and U13953 (N_13953,N_12866,N_12743);
xnor U13954 (N_13954,N_12548,N_12833);
xnor U13955 (N_13955,N_12604,N_12771);
nor U13956 (N_13956,N_12537,N_12618);
nand U13957 (N_13957,N_12180,N_12941);
xor U13958 (N_13958,N_12908,N_12903);
nor U13959 (N_13959,N_12623,N_12130);
and U13960 (N_13960,N_12444,N_12538);
xor U13961 (N_13961,N_12574,N_12652);
and U13962 (N_13962,N_12267,N_12658);
or U13963 (N_13963,N_12957,N_12831);
and U13964 (N_13964,N_12189,N_12870);
and U13965 (N_13965,N_12696,N_12780);
nor U13966 (N_13966,N_12281,N_12855);
nor U13967 (N_13967,N_12609,N_12698);
or U13968 (N_13968,N_12458,N_12710);
and U13969 (N_13969,N_12977,N_12746);
nor U13970 (N_13970,N_12288,N_12063);
nor U13971 (N_13971,N_12178,N_12957);
nand U13972 (N_13972,N_12386,N_12670);
nor U13973 (N_13973,N_12544,N_12626);
nand U13974 (N_13974,N_12364,N_12471);
nand U13975 (N_13975,N_12435,N_12745);
and U13976 (N_13976,N_12316,N_12482);
nand U13977 (N_13977,N_12770,N_12985);
and U13978 (N_13978,N_12412,N_12968);
or U13979 (N_13979,N_12927,N_12319);
or U13980 (N_13980,N_12486,N_12550);
nand U13981 (N_13981,N_12546,N_12566);
or U13982 (N_13982,N_12830,N_12260);
nor U13983 (N_13983,N_12037,N_12840);
and U13984 (N_13984,N_12416,N_12877);
and U13985 (N_13985,N_12570,N_12660);
nand U13986 (N_13986,N_12623,N_12923);
or U13987 (N_13987,N_12147,N_12537);
and U13988 (N_13988,N_12300,N_12931);
xnor U13989 (N_13989,N_12671,N_12003);
nand U13990 (N_13990,N_12974,N_12895);
nor U13991 (N_13991,N_12178,N_12903);
xnor U13992 (N_13992,N_12968,N_12107);
and U13993 (N_13993,N_12064,N_12074);
xnor U13994 (N_13994,N_12436,N_12070);
xor U13995 (N_13995,N_12468,N_12420);
and U13996 (N_13996,N_12987,N_12272);
nor U13997 (N_13997,N_12348,N_12180);
xnor U13998 (N_13998,N_12826,N_12801);
and U13999 (N_13999,N_12044,N_12644);
or U14000 (N_14000,N_13700,N_13562);
or U14001 (N_14001,N_13420,N_13231);
nand U14002 (N_14002,N_13290,N_13792);
and U14003 (N_14003,N_13873,N_13026);
and U14004 (N_14004,N_13281,N_13378);
xor U14005 (N_14005,N_13244,N_13286);
nor U14006 (N_14006,N_13314,N_13411);
and U14007 (N_14007,N_13487,N_13796);
nor U14008 (N_14008,N_13850,N_13312);
xor U14009 (N_14009,N_13085,N_13391);
nand U14010 (N_14010,N_13564,N_13886);
and U14011 (N_14011,N_13777,N_13876);
and U14012 (N_14012,N_13227,N_13473);
nand U14013 (N_14013,N_13406,N_13058);
nand U14014 (N_14014,N_13545,N_13152);
and U14015 (N_14015,N_13889,N_13456);
and U14016 (N_14016,N_13495,N_13797);
nand U14017 (N_14017,N_13134,N_13121);
or U14018 (N_14018,N_13900,N_13968);
nand U14019 (N_14019,N_13424,N_13434);
and U14020 (N_14020,N_13100,N_13809);
or U14021 (N_14021,N_13270,N_13893);
nand U14022 (N_14022,N_13661,N_13831);
and U14023 (N_14023,N_13385,N_13051);
nor U14024 (N_14024,N_13083,N_13645);
or U14025 (N_14025,N_13352,N_13032);
xor U14026 (N_14026,N_13490,N_13945);
nor U14027 (N_14027,N_13128,N_13158);
xnor U14028 (N_14028,N_13526,N_13810);
nor U14029 (N_14029,N_13961,N_13239);
and U14030 (N_14030,N_13366,N_13885);
nand U14031 (N_14031,N_13933,N_13837);
nand U14032 (N_14032,N_13834,N_13301);
or U14033 (N_14033,N_13588,N_13811);
nor U14034 (N_14034,N_13872,N_13418);
nand U14035 (N_14035,N_13108,N_13828);
xor U14036 (N_14036,N_13416,N_13899);
nor U14037 (N_14037,N_13536,N_13113);
and U14038 (N_14038,N_13677,N_13095);
xnor U14039 (N_14039,N_13435,N_13868);
nand U14040 (N_14040,N_13496,N_13116);
xor U14041 (N_14041,N_13742,N_13660);
nand U14042 (N_14042,N_13068,N_13315);
or U14043 (N_14043,N_13909,N_13120);
and U14044 (N_14044,N_13402,N_13842);
nor U14045 (N_14045,N_13171,N_13199);
nand U14046 (N_14046,N_13010,N_13392);
nor U14047 (N_14047,N_13519,N_13360);
nand U14048 (N_14048,N_13729,N_13617);
and U14049 (N_14049,N_13864,N_13509);
or U14050 (N_14050,N_13303,N_13350);
xnor U14051 (N_14051,N_13801,N_13339);
nor U14052 (N_14052,N_13881,N_13691);
xor U14053 (N_14053,N_13566,N_13727);
or U14054 (N_14054,N_13537,N_13400);
or U14055 (N_14055,N_13821,N_13606);
and U14056 (N_14056,N_13305,N_13017);
or U14057 (N_14057,N_13274,N_13920);
nand U14058 (N_14058,N_13813,N_13266);
and U14059 (N_14059,N_13141,N_13963);
nor U14060 (N_14060,N_13527,N_13877);
and U14061 (N_14061,N_13468,N_13452);
nand U14062 (N_14062,N_13501,N_13135);
nand U14063 (N_14063,N_13553,N_13043);
nor U14064 (N_14064,N_13084,N_13443);
nor U14065 (N_14065,N_13294,N_13172);
and U14066 (N_14066,N_13322,N_13634);
and U14067 (N_14067,N_13369,N_13637);
or U14068 (N_14068,N_13150,N_13246);
xor U14069 (N_14069,N_13204,N_13164);
xnor U14070 (N_14070,N_13169,N_13160);
xnor U14071 (N_14071,N_13410,N_13380);
xnor U14072 (N_14072,N_13200,N_13919);
nand U14073 (N_14073,N_13803,N_13089);
xor U14074 (N_14074,N_13897,N_13181);
or U14075 (N_14075,N_13002,N_13829);
or U14076 (N_14076,N_13975,N_13052);
and U14077 (N_14077,N_13447,N_13869);
or U14078 (N_14078,N_13003,N_13917);
xor U14079 (N_14079,N_13672,N_13236);
nor U14080 (N_14080,N_13093,N_13823);
and U14081 (N_14081,N_13921,N_13977);
and U14082 (N_14082,N_13067,N_13623);
nor U14083 (N_14083,N_13336,N_13839);
and U14084 (N_14084,N_13060,N_13870);
nand U14085 (N_14085,N_13807,N_13081);
xnor U14086 (N_14086,N_13958,N_13460);
nor U14087 (N_14087,N_13875,N_13138);
nor U14088 (N_14088,N_13604,N_13764);
xor U14089 (N_14089,N_13163,N_13191);
nand U14090 (N_14090,N_13551,N_13583);
or U14091 (N_14091,N_13155,N_13388);
nor U14092 (N_14092,N_13959,N_13636);
or U14093 (N_14093,N_13795,N_13210);
xnor U14094 (N_14094,N_13702,N_13770);
or U14095 (N_14095,N_13767,N_13045);
and U14096 (N_14096,N_13302,N_13678);
or U14097 (N_14097,N_13934,N_13321);
or U14098 (N_14098,N_13852,N_13642);
and U14099 (N_14099,N_13329,N_13653);
xor U14100 (N_14100,N_13713,N_13944);
nand U14101 (N_14101,N_13507,N_13820);
or U14102 (N_14102,N_13655,N_13215);
nor U14103 (N_14103,N_13405,N_13709);
nor U14104 (N_14104,N_13334,N_13225);
or U14105 (N_14105,N_13865,N_13034);
or U14106 (N_14106,N_13001,N_13086);
nand U14107 (N_14107,N_13912,N_13728);
and U14108 (N_14108,N_13048,N_13379);
xnor U14109 (N_14109,N_13656,N_13791);
nor U14110 (N_14110,N_13752,N_13976);
or U14111 (N_14111,N_13450,N_13166);
nand U14112 (N_14112,N_13740,N_13037);
nor U14113 (N_14113,N_13387,N_13457);
nor U14114 (N_14114,N_13162,N_13114);
and U14115 (N_14115,N_13620,N_13187);
xnor U14116 (N_14116,N_13768,N_13860);
nand U14117 (N_14117,N_13679,N_13971);
or U14118 (N_14118,N_13479,N_13466);
or U14119 (N_14119,N_13987,N_13218);
or U14120 (N_14120,N_13178,N_13065);
xor U14121 (N_14121,N_13248,N_13836);
nand U14122 (N_14122,N_13573,N_13408);
or U14123 (N_14123,N_13330,N_13287);
and U14124 (N_14124,N_13265,N_13147);
xor U14125 (N_14125,N_13586,N_13421);
and U14126 (N_14126,N_13039,N_13111);
nand U14127 (N_14127,N_13448,N_13070);
or U14128 (N_14128,N_13066,N_13716);
or U14129 (N_14129,N_13332,N_13175);
nor U14130 (N_14130,N_13931,N_13733);
or U14131 (N_14131,N_13597,N_13608);
nand U14132 (N_14132,N_13080,N_13861);
or U14133 (N_14133,N_13538,N_13982);
xnor U14134 (N_14134,N_13318,N_13022);
or U14135 (N_14135,N_13626,N_13619);
nor U14136 (N_14136,N_13185,N_13932);
xor U14137 (N_14137,N_13442,N_13346);
xor U14138 (N_14138,N_13962,N_13401);
or U14139 (N_14139,N_13041,N_13470);
and U14140 (N_14140,N_13947,N_13370);
or U14141 (N_14141,N_13874,N_13072);
nor U14142 (N_14142,N_13590,N_13396);
and U14143 (N_14143,N_13990,N_13296);
nand U14144 (N_14144,N_13168,N_13751);
and U14145 (N_14145,N_13485,N_13628);
and U14146 (N_14146,N_13004,N_13585);
nand U14147 (N_14147,N_13746,N_13433);
xnor U14148 (N_14148,N_13324,N_13698);
nand U14149 (N_14149,N_13109,N_13974);
nand U14150 (N_14150,N_13785,N_13731);
and U14151 (N_14151,N_13477,N_13295);
or U14152 (N_14152,N_13409,N_13146);
or U14153 (N_14153,N_13057,N_13983);
or U14154 (N_14154,N_13769,N_13725);
nor U14155 (N_14155,N_13474,N_13625);
nor U14156 (N_14156,N_13220,N_13841);
or U14157 (N_14157,N_13394,N_13825);
or U14158 (N_14158,N_13489,N_13510);
nor U14159 (N_14159,N_13614,N_13078);
xnor U14160 (N_14160,N_13978,N_13844);
and U14161 (N_14161,N_13595,N_13046);
xnor U14162 (N_14162,N_13268,N_13908);
and U14163 (N_14163,N_13613,N_13719);
nand U14164 (N_14164,N_13758,N_13923);
xor U14165 (N_14165,N_13817,N_13705);
nand U14166 (N_14166,N_13883,N_13596);
and U14167 (N_14167,N_13670,N_13224);
nor U14168 (N_14168,N_13355,N_13455);
or U14169 (N_14169,N_13822,N_13622);
and U14170 (N_14170,N_13542,N_13389);
and U14171 (N_14171,N_13759,N_13439);
or U14172 (N_14172,N_13251,N_13800);
or U14173 (N_14173,N_13998,N_13087);
xnor U14174 (N_14174,N_13621,N_13748);
or U14175 (N_14175,N_13763,N_13140);
and U14176 (N_14176,N_13079,N_13300);
and U14177 (N_14177,N_13565,N_13543);
nor U14178 (N_14178,N_13269,N_13518);
and U14179 (N_14179,N_13955,N_13319);
xor U14180 (N_14180,N_13765,N_13130);
and U14181 (N_14181,N_13571,N_13425);
and U14182 (N_14182,N_13694,N_13031);
xnor U14183 (N_14183,N_13690,N_13730);
xor U14184 (N_14184,N_13423,N_13560);
and U14185 (N_14185,N_13532,N_13640);
xnor U14186 (N_14186,N_13042,N_13833);
nor U14187 (N_14187,N_13107,N_13890);
xnor U14188 (N_14188,N_13991,N_13643);
nor U14189 (N_14189,N_13345,N_13972);
nor U14190 (N_14190,N_13309,N_13371);
nor U14191 (N_14191,N_13144,N_13522);
nor U14192 (N_14192,N_13292,N_13780);
nand U14193 (N_14193,N_13050,N_13584);
xor U14194 (N_14194,N_13009,N_13547);
or U14195 (N_14195,N_13372,N_13011);
or U14196 (N_14196,N_13335,N_13880);
nor U14197 (N_14197,N_13687,N_13040);
nor U14198 (N_14198,N_13732,N_13652);
nor U14199 (N_14199,N_13697,N_13206);
or U14200 (N_14200,N_13493,N_13232);
nand U14201 (N_14201,N_13126,N_13854);
nand U14202 (N_14202,N_13238,N_13271);
nand U14203 (N_14203,N_13465,N_13910);
or U14204 (N_14204,N_13024,N_13717);
and U14205 (N_14205,N_13306,N_13816);
nor U14206 (N_14206,N_13417,N_13293);
nor U14207 (N_14207,N_13013,N_13578);
nand U14208 (N_14208,N_13517,N_13341);
xnor U14209 (N_14209,N_13182,N_13307);
xnor U14210 (N_14210,N_13946,N_13888);
xor U14211 (N_14211,N_13985,N_13285);
nand U14212 (N_14212,N_13049,N_13170);
or U14213 (N_14213,N_13631,N_13499);
or U14214 (N_14214,N_13279,N_13895);
nand U14215 (N_14215,N_13221,N_13263);
nand U14216 (N_14216,N_13505,N_13942);
xnor U14217 (N_14217,N_13649,N_13407);
xnor U14218 (N_14218,N_13289,N_13283);
or U14219 (N_14219,N_13480,N_13139);
nand U14220 (N_14220,N_13815,N_13775);
and U14221 (N_14221,N_13374,N_13131);
or U14222 (N_14222,N_13119,N_13444);
or U14223 (N_14223,N_13761,N_13937);
nor U14224 (N_14224,N_13094,N_13217);
nor U14225 (N_14225,N_13514,N_13960);
nand U14226 (N_14226,N_13602,N_13755);
nand U14227 (N_14227,N_13552,N_13124);
xor U14228 (N_14228,N_13384,N_13711);
nand U14229 (N_14229,N_13824,N_13484);
nor U14230 (N_14230,N_13581,N_13249);
or U14231 (N_14231,N_13241,N_13492);
nor U14232 (N_14232,N_13927,N_13849);
and U14233 (N_14233,N_13575,N_13115);
and U14234 (N_14234,N_13007,N_13704);
nor U14235 (N_14235,N_13952,N_13062);
nor U14236 (N_14236,N_13667,N_13528);
nor U14237 (N_14237,N_13794,N_13282);
xnor U14238 (N_14238,N_13255,N_13964);
or U14239 (N_14239,N_13063,N_13659);
nor U14240 (N_14240,N_13530,N_13938);
nor U14241 (N_14241,N_13710,N_13390);
and U14242 (N_14242,N_13806,N_13340);
xnor U14243 (N_14243,N_13277,N_13627);
nor U14244 (N_14244,N_13999,N_13102);
nand U14245 (N_14245,N_13524,N_13023);
nor U14246 (N_14246,N_13356,N_13074);
nand U14247 (N_14247,N_13386,N_13859);
xor U14248 (N_14248,N_13563,N_13230);
xnor U14249 (N_14249,N_13110,N_13398);
xnor U14250 (N_14250,N_13061,N_13894);
nor U14251 (N_14251,N_13237,N_13592);
xnor U14252 (N_14252,N_13245,N_13579);
nor U14253 (N_14253,N_13684,N_13123);
and U14254 (N_14254,N_13980,N_13183);
and U14255 (N_14255,N_13916,N_13304);
and U14256 (N_14256,N_13475,N_13106);
and U14257 (N_14257,N_13438,N_13601);
nand U14258 (N_14258,N_13663,N_13478);
and U14259 (N_14259,N_13568,N_13205);
and U14260 (N_14260,N_13056,N_13903);
xnor U14261 (N_14261,N_13981,N_13097);
xor U14262 (N_14262,N_13202,N_13706);
nand U14263 (N_14263,N_13342,N_13539);
xor U14264 (N_14264,N_13789,N_13951);
or U14265 (N_14265,N_13693,N_13646);
or U14266 (N_14266,N_13317,N_13762);
nand U14267 (N_14267,N_13088,N_13979);
xor U14268 (N_14268,N_13574,N_13924);
xnor U14269 (N_14269,N_13272,N_13735);
nand U14270 (N_14270,N_13871,N_13177);
nor U14271 (N_14271,N_13949,N_13741);
and U14272 (N_14272,N_13472,N_13252);
nand U14273 (N_14273,N_13453,N_13898);
and U14274 (N_14274,N_13494,N_13149);
and U14275 (N_14275,N_13805,N_13207);
nand U14276 (N_14276,N_13180,N_13362);
nor U14277 (N_14277,N_13432,N_13257);
xor U14278 (N_14278,N_13544,N_13556);
xor U14279 (N_14279,N_13750,N_13333);
or U14280 (N_14280,N_13624,N_13887);
and U14281 (N_14281,N_13686,N_13683);
and U14282 (N_14282,N_13882,N_13772);
and U14283 (N_14283,N_13892,N_13491);
xor U14284 (N_14284,N_13075,N_13488);
or U14285 (N_14285,N_13462,N_13722);
and U14286 (N_14286,N_13261,N_13688);
nand U14287 (N_14287,N_13047,N_13243);
xor U14288 (N_14288,N_13993,N_13753);
nand U14289 (N_14289,N_13853,N_13469);
nand U14290 (N_14290,N_13776,N_13657);
and U14291 (N_14291,N_13373,N_13591);
nand U14292 (N_14292,N_13593,N_13577);
nand U14293 (N_14293,N_13395,N_13743);
and U14294 (N_14294,N_13662,N_13749);
xnor U14295 (N_14295,N_13630,N_13576);
xor U14296 (N_14296,N_13000,N_13965);
or U14297 (N_14297,N_13724,N_13835);
nand U14298 (N_14298,N_13328,N_13846);
and U14299 (N_14299,N_13142,N_13414);
nand U14300 (N_14300,N_13316,N_13830);
and U14301 (N_14301,N_13464,N_13648);
nand U14302 (N_14302,N_13349,N_13441);
and U14303 (N_14303,N_13254,N_13726);
or U14304 (N_14304,N_13471,N_13913);
nand U14305 (N_14305,N_13219,N_13941);
nand U14306 (N_14306,N_13247,N_13504);
or U14307 (N_14307,N_13012,N_13918);
or U14308 (N_14308,N_13523,N_13550);
or U14309 (N_14309,N_13943,N_13020);
nand U14310 (N_14310,N_13159,N_13760);
nand U14311 (N_14311,N_13548,N_13629);
nand U14312 (N_14312,N_13969,N_13610);
and U14313 (N_14313,N_13773,N_13914);
xnor U14314 (N_14314,N_13132,N_13071);
nand U14315 (N_14315,N_13612,N_13666);
and U14316 (N_14316,N_13156,N_13555);
or U14317 (N_14317,N_13264,N_13189);
nand U14318 (N_14318,N_13154,N_13481);
nand U14319 (N_14319,N_13165,N_13173);
nand U14320 (N_14320,N_13192,N_13745);
or U14321 (N_14321,N_13229,N_13174);
nor U14322 (N_14322,N_13896,N_13511);
nand U14323 (N_14323,N_13233,N_13948);
or U14324 (N_14324,N_13069,N_13615);
and U14325 (N_14325,N_13008,N_13073);
xor U14326 (N_14326,N_13779,N_13638);
or U14327 (N_14327,N_13436,N_13476);
nor U14328 (N_14328,N_13506,N_13720);
xnor U14329 (N_14329,N_13044,N_13025);
xor U14330 (N_14330,N_13325,N_13297);
nor U14331 (N_14331,N_13699,N_13580);
nor U14332 (N_14332,N_13734,N_13953);
or U14333 (N_14333,N_13376,N_13950);
or U14334 (N_14334,N_13611,N_13814);
nor U14335 (N_14335,N_13299,N_13879);
nor U14336 (N_14336,N_13430,N_13546);
xor U14337 (N_14337,N_13689,N_13675);
nor U14338 (N_14338,N_13736,N_13127);
xor U14339 (N_14339,N_13654,N_13320);
nand U14340 (N_14340,N_13226,N_13122);
xnor U14341 (N_14341,N_13925,N_13323);
or U14342 (N_14342,N_13030,N_13015);
xor U14343 (N_14343,N_13104,N_13862);
and U14344 (N_14344,N_13167,N_13313);
xor U14345 (N_14345,N_13529,N_13907);
and U14346 (N_14346,N_13808,N_13059);
nand U14347 (N_14347,N_13018,N_13723);
and U14348 (N_14348,N_13076,N_13184);
nor U14349 (N_14349,N_13367,N_13454);
nand U14350 (N_14350,N_13036,N_13714);
nand U14351 (N_14351,N_13996,N_13603);
xnor U14352 (N_14352,N_13804,N_13148);
nand U14353 (N_14353,N_13739,N_13747);
or U14354 (N_14354,N_13929,N_13354);
and U14355 (N_14355,N_13771,N_13326);
nor U14356 (N_14356,N_13639,N_13188);
nand U14357 (N_14357,N_13520,N_13599);
or U14358 (N_14358,N_13458,N_13533);
nand U14359 (N_14359,N_13103,N_13431);
xor U14360 (N_14360,N_13055,N_13812);
and U14361 (N_14361,N_13195,N_13486);
nor U14362 (N_14362,N_13682,N_13446);
and U14363 (N_14363,N_13014,N_13954);
nand U14364 (N_14364,N_13415,N_13117);
nand U14365 (N_14365,N_13926,N_13644);
nand U14366 (N_14366,N_13383,N_13358);
xor U14367 (N_14367,N_13905,N_13098);
and U14368 (N_14368,N_13557,N_13203);
or U14369 (N_14369,N_13549,N_13213);
xnor U14370 (N_14370,N_13701,N_13651);
or U14371 (N_14371,N_13986,N_13818);
nand U14372 (N_14372,N_13940,N_13695);
xor U14373 (N_14373,N_13449,N_13179);
or U14374 (N_14374,N_13005,N_13242);
xnor U14375 (N_14375,N_13368,N_13855);
nor U14376 (N_14376,N_13570,N_13344);
nor U14377 (N_14377,N_13534,N_13848);
nand U14378 (N_14378,N_13404,N_13778);
xor U14379 (N_14379,N_13228,N_13658);
or U14380 (N_14380,N_13176,N_13193);
nor U14381 (N_14381,N_13253,N_13482);
xnor U14382 (N_14382,N_13680,N_13561);
xnor U14383 (N_14383,N_13664,N_13707);
and U14384 (N_14384,N_13381,N_13754);
and U14385 (N_14385,N_13558,N_13559);
nand U14386 (N_14386,N_13145,N_13508);
nor U14387 (N_14387,N_13632,N_13463);
nand U14388 (N_14388,N_13994,N_13118);
xnor U14389 (N_14389,N_13647,N_13856);
or U14390 (N_14390,N_13311,N_13826);
and U14391 (N_14391,N_13607,N_13737);
nand U14392 (N_14392,N_13092,N_13708);
nor U14393 (N_14393,N_13721,N_13082);
nor U14394 (N_14394,N_13669,N_13798);
nand U14395 (N_14395,N_13851,N_13715);
nand U14396 (N_14396,N_13413,N_13609);
and U14397 (N_14397,N_13676,N_13525);
nor U14398 (N_14398,N_13382,N_13957);
xor U14399 (N_14399,N_13359,N_13995);
nor U14400 (N_14400,N_13194,N_13461);
or U14401 (N_14401,N_13250,N_13054);
nand U14402 (N_14402,N_13437,N_13766);
and U14403 (N_14403,N_13426,N_13594);
and U14404 (N_14404,N_13939,N_13616);
xnor U14405 (N_14405,N_13867,N_13930);
and U14406 (N_14406,N_13992,N_13989);
or U14407 (N_14407,N_13671,N_13674);
or U14408 (N_14408,N_13703,N_13902);
nor U14409 (N_14409,N_13275,N_13541);
nor U14410 (N_14410,N_13858,N_13567);
xnor U14411 (N_14411,N_13685,N_13211);
nand U14412 (N_14412,N_13845,N_13535);
nor U14413 (N_14413,N_13019,N_13515);
nand U14414 (N_14414,N_13832,N_13967);
xor U14415 (N_14415,N_13847,N_13774);
xnor U14416 (N_14416,N_13582,N_13235);
nand U14417 (N_14417,N_13668,N_13513);
and U14418 (N_14418,N_13936,N_13997);
nand U14419 (N_14419,N_13353,N_13214);
nor U14420 (N_14420,N_13337,N_13133);
nor U14421 (N_14421,N_13365,N_13298);
and U14422 (N_14422,N_13161,N_13310);
nand U14423 (N_14423,N_13006,N_13357);
nor U14424 (N_14424,N_13393,N_13222);
and U14425 (N_14425,N_13956,N_13843);
xor U14426 (N_14426,N_13459,N_13445);
or U14427 (N_14427,N_13273,N_13863);
or U14428 (N_14428,N_13331,N_13712);
nand U14429 (N_14429,N_13101,N_13276);
and U14430 (N_14430,N_13451,N_13259);
nor U14431 (N_14431,N_13572,N_13598);
xnor U14432 (N_14432,N_13665,N_13641);
nor U14433 (N_14433,N_13827,N_13600);
and U14434 (N_14434,N_13212,N_13738);
xnor U14435 (N_14435,N_13403,N_13267);
or U14436 (N_14436,N_13223,N_13799);
nor U14437 (N_14437,N_13467,N_13260);
nor U14438 (N_14438,N_13589,N_13428);
nand U14439 (N_14439,N_13531,N_13483);
or U14440 (N_14440,N_13540,N_13077);
and U14441 (N_14441,N_13209,N_13696);
nor U14442 (N_14442,N_13397,N_13338);
nor U14443 (N_14443,N_13783,N_13129);
and U14444 (N_14444,N_13064,N_13399);
nand U14445 (N_14445,N_13125,N_13099);
nor U14446 (N_14446,N_13096,N_13915);
nor U14447 (N_14447,N_13284,N_13198);
nand U14448 (N_14448,N_13197,N_13347);
nand U14449 (N_14449,N_13635,N_13262);
and U14450 (N_14450,N_13840,N_13970);
and U14451 (N_14451,N_13866,N_13819);
or U14452 (N_14452,N_13343,N_13498);
xor U14453 (N_14453,N_13419,N_13718);
and U14454 (N_14454,N_13053,N_13878);
and U14455 (N_14455,N_13781,N_13136);
nor U14456 (N_14456,N_13793,N_13802);
and U14457 (N_14457,N_13258,N_13891);
xnor U14458 (N_14458,N_13157,N_13782);
xor U14459 (N_14459,N_13605,N_13857);
nor U14460 (N_14460,N_13029,N_13928);
or U14461 (N_14461,N_13681,N_13935);
nor U14462 (N_14462,N_13966,N_13143);
xnor U14463 (N_14463,N_13786,N_13153);
xnor U14464 (N_14464,N_13105,N_13090);
xor U14465 (N_14465,N_13884,N_13633);
nor U14466 (N_14466,N_13911,N_13901);
or U14467 (N_14467,N_13650,N_13784);
nor U14468 (N_14468,N_13412,N_13502);
nor U14469 (N_14469,N_13521,N_13038);
and U14470 (N_14470,N_13240,N_13587);
and U14471 (N_14471,N_13035,N_13904);
nor U14472 (N_14472,N_13500,N_13692);
nand U14473 (N_14473,N_13351,N_13375);
and U14474 (N_14474,N_13363,N_13569);
nand U14475 (N_14475,N_13256,N_13137);
or U14476 (N_14476,N_13377,N_13196);
or U14477 (N_14477,N_13021,N_13278);
nand U14478 (N_14478,N_13922,N_13364);
and U14479 (N_14479,N_13757,N_13234);
nand U14480 (N_14480,N_13348,N_13288);
and U14481 (N_14481,N_13973,N_13790);
or U14482 (N_14482,N_13112,N_13216);
or U14483 (N_14483,N_13788,N_13091);
or U14484 (N_14484,N_13984,N_13673);
xnor U14485 (N_14485,N_13756,N_13201);
nor U14486 (N_14486,N_13186,N_13497);
and U14487 (N_14487,N_13033,N_13291);
nand U14488 (N_14488,N_13516,N_13838);
and U14489 (N_14489,N_13308,N_13988);
and U14490 (N_14490,N_13016,N_13208);
nand U14491 (N_14491,N_13440,N_13028);
nor U14492 (N_14492,N_13190,N_13280);
nand U14493 (N_14493,N_13429,N_13787);
and U14494 (N_14494,N_13151,N_13327);
or U14495 (N_14495,N_13422,N_13906);
xor U14496 (N_14496,N_13427,N_13027);
nor U14497 (N_14497,N_13554,N_13744);
nand U14498 (N_14498,N_13361,N_13503);
nand U14499 (N_14499,N_13512,N_13618);
nor U14500 (N_14500,N_13619,N_13200);
xor U14501 (N_14501,N_13460,N_13990);
or U14502 (N_14502,N_13200,N_13216);
and U14503 (N_14503,N_13339,N_13783);
nand U14504 (N_14504,N_13058,N_13417);
and U14505 (N_14505,N_13409,N_13089);
nand U14506 (N_14506,N_13951,N_13502);
and U14507 (N_14507,N_13413,N_13396);
and U14508 (N_14508,N_13269,N_13235);
nand U14509 (N_14509,N_13144,N_13652);
or U14510 (N_14510,N_13573,N_13491);
and U14511 (N_14511,N_13130,N_13329);
nor U14512 (N_14512,N_13179,N_13777);
nor U14513 (N_14513,N_13126,N_13539);
or U14514 (N_14514,N_13441,N_13763);
nor U14515 (N_14515,N_13189,N_13895);
or U14516 (N_14516,N_13251,N_13021);
and U14517 (N_14517,N_13055,N_13002);
xor U14518 (N_14518,N_13468,N_13554);
xor U14519 (N_14519,N_13886,N_13372);
nand U14520 (N_14520,N_13176,N_13136);
or U14521 (N_14521,N_13001,N_13333);
nor U14522 (N_14522,N_13929,N_13762);
xor U14523 (N_14523,N_13157,N_13623);
nor U14524 (N_14524,N_13700,N_13118);
xnor U14525 (N_14525,N_13670,N_13880);
nor U14526 (N_14526,N_13060,N_13339);
or U14527 (N_14527,N_13534,N_13753);
xnor U14528 (N_14528,N_13239,N_13528);
nor U14529 (N_14529,N_13656,N_13895);
and U14530 (N_14530,N_13104,N_13329);
xnor U14531 (N_14531,N_13588,N_13686);
or U14532 (N_14532,N_13212,N_13870);
and U14533 (N_14533,N_13117,N_13243);
nor U14534 (N_14534,N_13211,N_13897);
xor U14535 (N_14535,N_13839,N_13406);
or U14536 (N_14536,N_13169,N_13250);
nor U14537 (N_14537,N_13419,N_13774);
or U14538 (N_14538,N_13861,N_13621);
and U14539 (N_14539,N_13220,N_13604);
nand U14540 (N_14540,N_13077,N_13942);
and U14541 (N_14541,N_13363,N_13338);
nor U14542 (N_14542,N_13058,N_13519);
nand U14543 (N_14543,N_13294,N_13971);
or U14544 (N_14544,N_13519,N_13109);
nor U14545 (N_14545,N_13827,N_13966);
nor U14546 (N_14546,N_13078,N_13900);
nor U14547 (N_14547,N_13726,N_13748);
nor U14548 (N_14548,N_13684,N_13390);
nor U14549 (N_14549,N_13365,N_13542);
nand U14550 (N_14550,N_13053,N_13439);
nand U14551 (N_14551,N_13205,N_13169);
and U14552 (N_14552,N_13634,N_13255);
nor U14553 (N_14553,N_13391,N_13771);
or U14554 (N_14554,N_13451,N_13872);
xnor U14555 (N_14555,N_13528,N_13513);
and U14556 (N_14556,N_13669,N_13558);
nor U14557 (N_14557,N_13057,N_13490);
or U14558 (N_14558,N_13680,N_13757);
nand U14559 (N_14559,N_13300,N_13548);
and U14560 (N_14560,N_13193,N_13904);
nand U14561 (N_14561,N_13051,N_13371);
and U14562 (N_14562,N_13400,N_13912);
and U14563 (N_14563,N_13164,N_13324);
and U14564 (N_14564,N_13842,N_13807);
or U14565 (N_14565,N_13692,N_13843);
and U14566 (N_14566,N_13725,N_13045);
or U14567 (N_14567,N_13536,N_13588);
nor U14568 (N_14568,N_13043,N_13332);
and U14569 (N_14569,N_13493,N_13696);
nand U14570 (N_14570,N_13855,N_13397);
xnor U14571 (N_14571,N_13147,N_13109);
and U14572 (N_14572,N_13264,N_13918);
nor U14573 (N_14573,N_13569,N_13884);
or U14574 (N_14574,N_13568,N_13831);
or U14575 (N_14575,N_13503,N_13804);
and U14576 (N_14576,N_13909,N_13847);
and U14577 (N_14577,N_13969,N_13604);
or U14578 (N_14578,N_13739,N_13734);
nand U14579 (N_14579,N_13030,N_13119);
or U14580 (N_14580,N_13308,N_13544);
and U14581 (N_14581,N_13071,N_13964);
or U14582 (N_14582,N_13949,N_13721);
or U14583 (N_14583,N_13126,N_13026);
nand U14584 (N_14584,N_13643,N_13572);
nand U14585 (N_14585,N_13864,N_13230);
nor U14586 (N_14586,N_13114,N_13510);
or U14587 (N_14587,N_13613,N_13726);
nand U14588 (N_14588,N_13556,N_13070);
nand U14589 (N_14589,N_13004,N_13979);
or U14590 (N_14590,N_13168,N_13701);
nor U14591 (N_14591,N_13732,N_13830);
nand U14592 (N_14592,N_13248,N_13796);
xor U14593 (N_14593,N_13270,N_13945);
xor U14594 (N_14594,N_13411,N_13067);
xor U14595 (N_14595,N_13330,N_13875);
or U14596 (N_14596,N_13363,N_13398);
nor U14597 (N_14597,N_13069,N_13712);
and U14598 (N_14598,N_13346,N_13386);
nor U14599 (N_14599,N_13623,N_13946);
nand U14600 (N_14600,N_13497,N_13927);
or U14601 (N_14601,N_13510,N_13553);
xnor U14602 (N_14602,N_13785,N_13240);
or U14603 (N_14603,N_13669,N_13323);
nor U14604 (N_14604,N_13397,N_13889);
or U14605 (N_14605,N_13325,N_13601);
nor U14606 (N_14606,N_13160,N_13768);
xnor U14607 (N_14607,N_13663,N_13044);
and U14608 (N_14608,N_13242,N_13663);
or U14609 (N_14609,N_13911,N_13661);
nor U14610 (N_14610,N_13003,N_13204);
and U14611 (N_14611,N_13421,N_13797);
nor U14612 (N_14612,N_13122,N_13174);
nor U14613 (N_14613,N_13708,N_13583);
and U14614 (N_14614,N_13677,N_13348);
nor U14615 (N_14615,N_13730,N_13254);
xor U14616 (N_14616,N_13248,N_13562);
nor U14617 (N_14617,N_13637,N_13866);
and U14618 (N_14618,N_13326,N_13007);
and U14619 (N_14619,N_13747,N_13108);
nor U14620 (N_14620,N_13584,N_13301);
nor U14621 (N_14621,N_13933,N_13447);
or U14622 (N_14622,N_13085,N_13591);
and U14623 (N_14623,N_13576,N_13870);
nand U14624 (N_14624,N_13572,N_13498);
nand U14625 (N_14625,N_13929,N_13317);
nor U14626 (N_14626,N_13204,N_13749);
or U14627 (N_14627,N_13527,N_13766);
xor U14628 (N_14628,N_13532,N_13539);
nand U14629 (N_14629,N_13302,N_13125);
and U14630 (N_14630,N_13996,N_13238);
or U14631 (N_14631,N_13277,N_13842);
and U14632 (N_14632,N_13202,N_13494);
nor U14633 (N_14633,N_13561,N_13292);
or U14634 (N_14634,N_13620,N_13279);
and U14635 (N_14635,N_13854,N_13736);
and U14636 (N_14636,N_13127,N_13808);
xor U14637 (N_14637,N_13729,N_13615);
nand U14638 (N_14638,N_13941,N_13787);
or U14639 (N_14639,N_13219,N_13340);
or U14640 (N_14640,N_13351,N_13986);
nor U14641 (N_14641,N_13058,N_13197);
and U14642 (N_14642,N_13823,N_13970);
and U14643 (N_14643,N_13112,N_13110);
xnor U14644 (N_14644,N_13192,N_13875);
xnor U14645 (N_14645,N_13129,N_13516);
or U14646 (N_14646,N_13690,N_13149);
or U14647 (N_14647,N_13084,N_13844);
and U14648 (N_14648,N_13409,N_13291);
nor U14649 (N_14649,N_13948,N_13405);
or U14650 (N_14650,N_13978,N_13152);
and U14651 (N_14651,N_13877,N_13021);
or U14652 (N_14652,N_13520,N_13472);
or U14653 (N_14653,N_13782,N_13406);
and U14654 (N_14654,N_13309,N_13976);
and U14655 (N_14655,N_13660,N_13987);
nand U14656 (N_14656,N_13349,N_13635);
nand U14657 (N_14657,N_13526,N_13120);
and U14658 (N_14658,N_13749,N_13759);
nand U14659 (N_14659,N_13056,N_13062);
nand U14660 (N_14660,N_13536,N_13827);
nor U14661 (N_14661,N_13608,N_13134);
xor U14662 (N_14662,N_13265,N_13119);
nor U14663 (N_14663,N_13873,N_13913);
and U14664 (N_14664,N_13283,N_13019);
or U14665 (N_14665,N_13664,N_13858);
xor U14666 (N_14666,N_13752,N_13967);
xor U14667 (N_14667,N_13107,N_13899);
or U14668 (N_14668,N_13500,N_13298);
xnor U14669 (N_14669,N_13642,N_13557);
nand U14670 (N_14670,N_13386,N_13331);
nand U14671 (N_14671,N_13131,N_13375);
xor U14672 (N_14672,N_13776,N_13304);
or U14673 (N_14673,N_13316,N_13359);
xor U14674 (N_14674,N_13368,N_13886);
or U14675 (N_14675,N_13799,N_13710);
and U14676 (N_14676,N_13626,N_13640);
nand U14677 (N_14677,N_13137,N_13470);
xnor U14678 (N_14678,N_13303,N_13500);
nor U14679 (N_14679,N_13633,N_13092);
xnor U14680 (N_14680,N_13199,N_13570);
or U14681 (N_14681,N_13772,N_13341);
or U14682 (N_14682,N_13845,N_13589);
and U14683 (N_14683,N_13830,N_13960);
or U14684 (N_14684,N_13451,N_13382);
or U14685 (N_14685,N_13880,N_13743);
or U14686 (N_14686,N_13093,N_13367);
or U14687 (N_14687,N_13730,N_13349);
xor U14688 (N_14688,N_13030,N_13856);
xor U14689 (N_14689,N_13991,N_13306);
nor U14690 (N_14690,N_13083,N_13133);
nand U14691 (N_14691,N_13078,N_13757);
or U14692 (N_14692,N_13738,N_13981);
or U14693 (N_14693,N_13472,N_13611);
or U14694 (N_14694,N_13081,N_13784);
and U14695 (N_14695,N_13557,N_13872);
nand U14696 (N_14696,N_13943,N_13501);
and U14697 (N_14697,N_13288,N_13510);
xor U14698 (N_14698,N_13480,N_13957);
or U14699 (N_14699,N_13137,N_13797);
and U14700 (N_14700,N_13322,N_13298);
nor U14701 (N_14701,N_13855,N_13270);
xnor U14702 (N_14702,N_13321,N_13542);
xor U14703 (N_14703,N_13475,N_13163);
nand U14704 (N_14704,N_13866,N_13075);
nand U14705 (N_14705,N_13774,N_13413);
xnor U14706 (N_14706,N_13725,N_13920);
and U14707 (N_14707,N_13622,N_13497);
nor U14708 (N_14708,N_13942,N_13244);
nor U14709 (N_14709,N_13754,N_13944);
or U14710 (N_14710,N_13250,N_13678);
nor U14711 (N_14711,N_13982,N_13883);
and U14712 (N_14712,N_13054,N_13838);
or U14713 (N_14713,N_13642,N_13734);
or U14714 (N_14714,N_13312,N_13774);
or U14715 (N_14715,N_13284,N_13197);
and U14716 (N_14716,N_13565,N_13025);
nor U14717 (N_14717,N_13183,N_13533);
xnor U14718 (N_14718,N_13986,N_13534);
xnor U14719 (N_14719,N_13423,N_13557);
nand U14720 (N_14720,N_13387,N_13553);
nand U14721 (N_14721,N_13356,N_13927);
xnor U14722 (N_14722,N_13893,N_13479);
or U14723 (N_14723,N_13717,N_13639);
or U14724 (N_14724,N_13055,N_13411);
and U14725 (N_14725,N_13632,N_13147);
or U14726 (N_14726,N_13345,N_13484);
or U14727 (N_14727,N_13461,N_13292);
nand U14728 (N_14728,N_13054,N_13976);
nand U14729 (N_14729,N_13486,N_13184);
nor U14730 (N_14730,N_13483,N_13709);
xnor U14731 (N_14731,N_13576,N_13189);
and U14732 (N_14732,N_13190,N_13167);
nand U14733 (N_14733,N_13866,N_13844);
nand U14734 (N_14734,N_13941,N_13312);
xor U14735 (N_14735,N_13368,N_13363);
xor U14736 (N_14736,N_13316,N_13449);
and U14737 (N_14737,N_13295,N_13930);
xnor U14738 (N_14738,N_13273,N_13274);
or U14739 (N_14739,N_13589,N_13947);
nor U14740 (N_14740,N_13156,N_13545);
nand U14741 (N_14741,N_13926,N_13622);
nand U14742 (N_14742,N_13442,N_13901);
and U14743 (N_14743,N_13839,N_13716);
nand U14744 (N_14744,N_13647,N_13681);
xor U14745 (N_14745,N_13063,N_13409);
xor U14746 (N_14746,N_13575,N_13080);
or U14747 (N_14747,N_13428,N_13171);
nand U14748 (N_14748,N_13484,N_13892);
nor U14749 (N_14749,N_13701,N_13532);
and U14750 (N_14750,N_13118,N_13841);
xor U14751 (N_14751,N_13077,N_13987);
xnor U14752 (N_14752,N_13018,N_13974);
xor U14753 (N_14753,N_13720,N_13570);
xnor U14754 (N_14754,N_13609,N_13561);
or U14755 (N_14755,N_13922,N_13173);
and U14756 (N_14756,N_13321,N_13666);
or U14757 (N_14757,N_13510,N_13882);
or U14758 (N_14758,N_13326,N_13293);
nand U14759 (N_14759,N_13835,N_13508);
nor U14760 (N_14760,N_13060,N_13370);
xor U14761 (N_14761,N_13458,N_13679);
nor U14762 (N_14762,N_13748,N_13361);
nor U14763 (N_14763,N_13483,N_13327);
xor U14764 (N_14764,N_13439,N_13648);
xor U14765 (N_14765,N_13687,N_13134);
xor U14766 (N_14766,N_13683,N_13367);
xnor U14767 (N_14767,N_13675,N_13327);
nor U14768 (N_14768,N_13323,N_13133);
and U14769 (N_14769,N_13488,N_13696);
nand U14770 (N_14770,N_13113,N_13891);
and U14771 (N_14771,N_13377,N_13447);
nand U14772 (N_14772,N_13313,N_13246);
xnor U14773 (N_14773,N_13567,N_13989);
nor U14774 (N_14774,N_13240,N_13768);
nor U14775 (N_14775,N_13222,N_13213);
nand U14776 (N_14776,N_13131,N_13102);
xor U14777 (N_14777,N_13208,N_13825);
and U14778 (N_14778,N_13409,N_13785);
nand U14779 (N_14779,N_13975,N_13895);
nand U14780 (N_14780,N_13459,N_13871);
nand U14781 (N_14781,N_13951,N_13464);
and U14782 (N_14782,N_13435,N_13756);
and U14783 (N_14783,N_13744,N_13392);
nor U14784 (N_14784,N_13215,N_13410);
nand U14785 (N_14785,N_13011,N_13916);
xor U14786 (N_14786,N_13066,N_13897);
nand U14787 (N_14787,N_13330,N_13756);
nand U14788 (N_14788,N_13613,N_13286);
nand U14789 (N_14789,N_13505,N_13221);
and U14790 (N_14790,N_13275,N_13908);
nor U14791 (N_14791,N_13701,N_13000);
or U14792 (N_14792,N_13920,N_13910);
nor U14793 (N_14793,N_13499,N_13371);
and U14794 (N_14794,N_13250,N_13106);
or U14795 (N_14795,N_13888,N_13443);
or U14796 (N_14796,N_13160,N_13024);
xor U14797 (N_14797,N_13945,N_13032);
and U14798 (N_14798,N_13189,N_13065);
and U14799 (N_14799,N_13421,N_13347);
and U14800 (N_14800,N_13110,N_13632);
and U14801 (N_14801,N_13763,N_13459);
or U14802 (N_14802,N_13648,N_13009);
or U14803 (N_14803,N_13604,N_13861);
xor U14804 (N_14804,N_13925,N_13555);
nor U14805 (N_14805,N_13097,N_13226);
or U14806 (N_14806,N_13425,N_13528);
and U14807 (N_14807,N_13062,N_13265);
or U14808 (N_14808,N_13193,N_13625);
and U14809 (N_14809,N_13204,N_13736);
nand U14810 (N_14810,N_13556,N_13482);
xnor U14811 (N_14811,N_13423,N_13823);
nand U14812 (N_14812,N_13041,N_13894);
and U14813 (N_14813,N_13084,N_13690);
or U14814 (N_14814,N_13485,N_13949);
nor U14815 (N_14815,N_13699,N_13530);
and U14816 (N_14816,N_13818,N_13684);
xor U14817 (N_14817,N_13551,N_13595);
and U14818 (N_14818,N_13045,N_13294);
xor U14819 (N_14819,N_13295,N_13667);
and U14820 (N_14820,N_13297,N_13191);
nor U14821 (N_14821,N_13404,N_13371);
nand U14822 (N_14822,N_13935,N_13369);
or U14823 (N_14823,N_13893,N_13601);
nor U14824 (N_14824,N_13110,N_13661);
and U14825 (N_14825,N_13394,N_13803);
xor U14826 (N_14826,N_13616,N_13341);
and U14827 (N_14827,N_13989,N_13036);
and U14828 (N_14828,N_13717,N_13753);
and U14829 (N_14829,N_13009,N_13021);
and U14830 (N_14830,N_13438,N_13572);
xnor U14831 (N_14831,N_13535,N_13331);
nand U14832 (N_14832,N_13013,N_13605);
or U14833 (N_14833,N_13983,N_13961);
or U14834 (N_14834,N_13181,N_13433);
xor U14835 (N_14835,N_13557,N_13301);
xor U14836 (N_14836,N_13905,N_13764);
and U14837 (N_14837,N_13504,N_13602);
and U14838 (N_14838,N_13036,N_13230);
nand U14839 (N_14839,N_13273,N_13377);
nor U14840 (N_14840,N_13221,N_13770);
and U14841 (N_14841,N_13480,N_13964);
nor U14842 (N_14842,N_13827,N_13457);
or U14843 (N_14843,N_13934,N_13562);
or U14844 (N_14844,N_13121,N_13054);
and U14845 (N_14845,N_13091,N_13889);
nor U14846 (N_14846,N_13818,N_13526);
nand U14847 (N_14847,N_13205,N_13678);
and U14848 (N_14848,N_13160,N_13533);
nor U14849 (N_14849,N_13560,N_13186);
and U14850 (N_14850,N_13491,N_13431);
xor U14851 (N_14851,N_13256,N_13558);
nor U14852 (N_14852,N_13927,N_13899);
nand U14853 (N_14853,N_13439,N_13548);
nand U14854 (N_14854,N_13768,N_13652);
nand U14855 (N_14855,N_13402,N_13333);
nand U14856 (N_14856,N_13022,N_13641);
nor U14857 (N_14857,N_13324,N_13145);
nand U14858 (N_14858,N_13349,N_13454);
xnor U14859 (N_14859,N_13477,N_13327);
nor U14860 (N_14860,N_13665,N_13238);
nor U14861 (N_14861,N_13405,N_13876);
xnor U14862 (N_14862,N_13030,N_13037);
or U14863 (N_14863,N_13399,N_13243);
or U14864 (N_14864,N_13875,N_13063);
nor U14865 (N_14865,N_13938,N_13634);
xor U14866 (N_14866,N_13724,N_13320);
nand U14867 (N_14867,N_13768,N_13834);
nand U14868 (N_14868,N_13551,N_13990);
nor U14869 (N_14869,N_13368,N_13584);
xor U14870 (N_14870,N_13327,N_13824);
nor U14871 (N_14871,N_13473,N_13583);
xor U14872 (N_14872,N_13279,N_13002);
xnor U14873 (N_14873,N_13149,N_13951);
or U14874 (N_14874,N_13422,N_13914);
xnor U14875 (N_14875,N_13894,N_13966);
xor U14876 (N_14876,N_13728,N_13413);
nor U14877 (N_14877,N_13405,N_13691);
or U14878 (N_14878,N_13187,N_13405);
and U14879 (N_14879,N_13419,N_13783);
and U14880 (N_14880,N_13588,N_13998);
nor U14881 (N_14881,N_13964,N_13914);
nand U14882 (N_14882,N_13494,N_13316);
and U14883 (N_14883,N_13200,N_13156);
nor U14884 (N_14884,N_13118,N_13532);
or U14885 (N_14885,N_13123,N_13278);
and U14886 (N_14886,N_13253,N_13599);
or U14887 (N_14887,N_13443,N_13464);
nand U14888 (N_14888,N_13098,N_13735);
nand U14889 (N_14889,N_13700,N_13993);
nor U14890 (N_14890,N_13610,N_13290);
and U14891 (N_14891,N_13082,N_13209);
and U14892 (N_14892,N_13616,N_13121);
nand U14893 (N_14893,N_13766,N_13929);
xnor U14894 (N_14894,N_13380,N_13444);
or U14895 (N_14895,N_13647,N_13966);
nor U14896 (N_14896,N_13470,N_13784);
nand U14897 (N_14897,N_13071,N_13740);
or U14898 (N_14898,N_13391,N_13198);
and U14899 (N_14899,N_13113,N_13780);
nand U14900 (N_14900,N_13072,N_13480);
xor U14901 (N_14901,N_13424,N_13671);
nor U14902 (N_14902,N_13419,N_13225);
or U14903 (N_14903,N_13660,N_13195);
nand U14904 (N_14904,N_13610,N_13271);
and U14905 (N_14905,N_13864,N_13520);
nor U14906 (N_14906,N_13290,N_13896);
nand U14907 (N_14907,N_13336,N_13752);
nand U14908 (N_14908,N_13650,N_13639);
nor U14909 (N_14909,N_13330,N_13250);
and U14910 (N_14910,N_13033,N_13544);
or U14911 (N_14911,N_13917,N_13757);
or U14912 (N_14912,N_13610,N_13949);
xnor U14913 (N_14913,N_13552,N_13455);
or U14914 (N_14914,N_13687,N_13630);
nor U14915 (N_14915,N_13332,N_13294);
nor U14916 (N_14916,N_13349,N_13947);
xnor U14917 (N_14917,N_13993,N_13163);
nor U14918 (N_14918,N_13507,N_13693);
nand U14919 (N_14919,N_13023,N_13009);
xor U14920 (N_14920,N_13137,N_13435);
and U14921 (N_14921,N_13352,N_13106);
nor U14922 (N_14922,N_13510,N_13191);
nand U14923 (N_14923,N_13005,N_13851);
nand U14924 (N_14924,N_13439,N_13086);
nand U14925 (N_14925,N_13054,N_13178);
and U14926 (N_14926,N_13359,N_13825);
and U14927 (N_14927,N_13953,N_13774);
or U14928 (N_14928,N_13791,N_13465);
xor U14929 (N_14929,N_13067,N_13542);
nand U14930 (N_14930,N_13771,N_13353);
nor U14931 (N_14931,N_13869,N_13436);
or U14932 (N_14932,N_13576,N_13531);
nor U14933 (N_14933,N_13975,N_13775);
xnor U14934 (N_14934,N_13647,N_13304);
nand U14935 (N_14935,N_13542,N_13469);
or U14936 (N_14936,N_13343,N_13226);
or U14937 (N_14937,N_13778,N_13553);
xnor U14938 (N_14938,N_13483,N_13611);
nand U14939 (N_14939,N_13474,N_13772);
or U14940 (N_14940,N_13525,N_13793);
and U14941 (N_14941,N_13826,N_13467);
xnor U14942 (N_14942,N_13436,N_13318);
and U14943 (N_14943,N_13659,N_13135);
nor U14944 (N_14944,N_13264,N_13708);
or U14945 (N_14945,N_13393,N_13806);
nand U14946 (N_14946,N_13555,N_13910);
xor U14947 (N_14947,N_13719,N_13240);
and U14948 (N_14948,N_13630,N_13269);
nand U14949 (N_14949,N_13676,N_13722);
and U14950 (N_14950,N_13864,N_13396);
and U14951 (N_14951,N_13775,N_13848);
or U14952 (N_14952,N_13381,N_13542);
or U14953 (N_14953,N_13427,N_13686);
and U14954 (N_14954,N_13016,N_13259);
nand U14955 (N_14955,N_13376,N_13363);
xor U14956 (N_14956,N_13549,N_13918);
and U14957 (N_14957,N_13963,N_13430);
nor U14958 (N_14958,N_13171,N_13004);
or U14959 (N_14959,N_13222,N_13085);
nand U14960 (N_14960,N_13391,N_13924);
and U14961 (N_14961,N_13469,N_13823);
xnor U14962 (N_14962,N_13366,N_13382);
nand U14963 (N_14963,N_13403,N_13273);
nand U14964 (N_14964,N_13570,N_13355);
and U14965 (N_14965,N_13834,N_13529);
and U14966 (N_14966,N_13714,N_13441);
nor U14967 (N_14967,N_13213,N_13707);
and U14968 (N_14968,N_13740,N_13091);
or U14969 (N_14969,N_13984,N_13270);
nand U14970 (N_14970,N_13638,N_13843);
xnor U14971 (N_14971,N_13202,N_13734);
or U14972 (N_14972,N_13963,N_13039);
and U14973 (N_14973,N_13232,N_13736);
xnor U14974 (N_14974,N_13136,N_13435);
xnor U14975 (N_14975,N_13682,N_13575);
nor U14976 (N_14976,N_13016,N_13705);
or U14977 (N_14977,N_13853,N_13744);
and U14978 (N_14978,N_13865,N_13347);
nor U14979 (N_14979,N_13083,N_13538);
nand U14980 (N_14980,N_13338,N_13023);
nor U14981 (N_14981,N_13093,N_13644);
xnor U14982 (N_14982,N_13821,N_13879);
nand U14983 (N_14983,N_13452,N_13731);
nor U14984 (N_14984,N_13084,N_13995);
xnor U14985 (N_14985,N_13591,N_13339);
or U14986 (N_14986,N_13474,N_13393);
or U14987 (N_14987,N_13834,N_13784);
xnor U14988 (N_14988,N_13353,N_13618);
nor U14989 (N_14989,N_13487,N_13648);
nor U14990 (N_14990,N_13458,N_13465);
nor U14991 (N_14991,N_13464,N_13274);
nand U14992 (N_14992,N_13513,N_13359);
and U14993 (N_14993,N_13971,N_13677);
nor U14994 (N_14994,N_13780,N_13065);
nor U14995 (N_14995,N_13450,N_13858);
or U14996 (N_14996,N_13273,N_13351);
nor U14997 (N_14997,N_13597,N_13540);
nor U14998 (N_14998,N_13293,N_13155);
or U14999 (N_14999,N_13761,N_13664);
xnor U15000 (N_15000,N_14757,N_14529);
nor U15001 (N_15001,N_14052,N_14148);
and U15002 (N_15002,N_14895,N_14259);
nand U15003 (N_15003,N_14696,N_14044);
xor U15004 (N_15004,N_14103,N_14745);
nor U15005 (N_15005,N_14706,N_14087);
nor U15006 (N_15006,N_14917,N_14024);
nand U15007 (N_15007,N_14976,N_14017);
or U15008 (N_15008,N_14955,N_14187);
xnor U15009 (N_15009,N_14786,N_14344);
nor U15010 (N_15010,N_14340,N_14758);
and U15011 (N_15011,N_14799,N_14514);
nor U15012 (N_15012,N_14948,N_14824);
xor U15013 (N_15013,N_14361,N_14167);
and U15014 (N_15014,N_14082,N_14375);
and U15015 (N_15015,N_14847,N_14715);
and U15016 (N_15016,N_14341,N_14887);
nand U15017 (N_15017,N_14343,N_14671);
or U15018 (N_15018,N_14525,N_14518);
or U15019 (N_15019,N_14694,N_14399);
nor U15020 (N_15020,N_14284,N_14446);
nor U15021 (N_15021,N_14179,N_14865);
and U15022 (N_15022,N_14538,N_14803);
nor U15023 (N_15023,N_14633,N_14337);
xnor U15024 (N_15024,N_14703,N_14926);
xnor U15025 (N_15025,N_14606,N_14330);
nor U15026 (N_15026,N_14669,N_14235);
xor U15027 (N_15027,N_14198,N_14298);
or U15028 (N_15028,N_14062,N_14873);
nand U15029 (N_15029,N_14989,N_14688);
nor U15030 (N_15030,N_14624,N_14582);
nor U15031 (N_15031,N_14831,N_14505);
nor U15032 (N_15032,N_14072,N_14580);
nand U15033 (N_15033,N_14031,N_14933);
nor U15034 (N_15034,N_14921,N_14172);
nor U15035 (N_15035,N_14697,N_14982);
nor U15036 (N_15036,N_14101,N_14882);
nor U15037 (N_15037,N_14060,N_14117);
or U15038 (N_15038,N_14675,N_14796);
nor U15039 (N_15039,N_14281,N_14137);
xnor U15040 (N_15040,N_14025,N_14480);
xnor U15041 (N_15041,N_14422,N_14490);
xnor U15042 (N_15042,N_14618,N_14195);
and U15043 (N_15043,N_14682,N_14864);
or U15044 (N_15044,N_14977,N_14056);
or U15045 (N_15045,N_14731,N_14540);
xnor U15046 (N_15046,N_14720,N_14637);
xor U15047 (N_15047,N_14849,N_14829);
or U15048 (N_15048,N_14738,N_14274);
xor U15049 (N_15049,N_14070,N_14657);
nand U15050 (N_15050,N_14171,N_14838);
xor U15051 (N_15051,N_14477,N_14109);
xnor U15052 (N_15052,N_14812,N_14810);
xnor U15053 (N_15053,N_14635,N_14748);
nand U15054 (N_15054,N_14861,N_14742);
nand U15055 (N_15055,N_14627,N_14462);
nand U15056 (N_15056,N_14068,N_14604);
or U15057 (N_15057,N_14503,N_14793);
xor U15058 (N_15058,N_14721,N_14150);
nor U15059 (N_15059,N_14862,N_14196);
or U15060 (N_15060,N_14636,N_14572);
nand U15061 (N_15061,N_14750,N_14765);
or U15062 (N_15062,N_14863,N_14647);
xnor U15063 (N_15063,N_14037,N_14941);
and U15064 (N_15064,N_14421,N_14692);
xnor U15065 (N_15065,N_14248,N_14419);
xor U15066 (N_15066,N_14869,N_14559);
nor U15067 (N_15067,N_14183,N_14632);
nand U15068 (N_15068,N_14276,N_14913);
xor U15069 (N_15069,N_14549,N_14766);
nor U15070 (N_15070,N_14412,N_14759);
and U15071 (N_15071,N_14231,N_14883);
nor U15072 (N_15072,N_14186,N_14565);
and U15073 (N_15073,N_14079,N_14428);
xnor U15074 (N_15074,N_14224,N_14468);
or U15075 (N_15075,N_14752,N_14764);
nor U15076 (N_15076,N_14992,N_14312);
nand U15077 (N_15077,N_14270,N_14612);
nand U15078 (N_15078,N_14794,N_14979);
xnor U15079 (N_15079,N_14147,N_14449);
or U15080 (N_15080,N_14719,N_14656);
nand U15081 (N_15081,N_14489,N_14120);
or U15082 (N_15082,N_14563,N_14176);
xor U15083 (N_15083,N_14965,N_14386);
nor U15084 (N_15084,N_14725,N_14564);
xnor U15085 (N_15085,N_14999,N_14493);
or U15086 (N_15086,N_14896,N_14839);
and U15087 (N_15087,N_14121,N_14322);
xor U15088 (N_15088,N_14980,N_14436);
nor U15089 (N_15089,N_14767,N_14324);
nor U15090 (N_15090,N_14676,N_14755);
nand U15091 (N_15091,N_14258,N_14374);
nand U15092 (N_15092,N_14389,N_14901);
xnor U15093 (N_15093,N_14283,N_14491);
xor U15094 (N_15094,N_14294,N_14898);
nor U15095 (N_15095,N_14732,N_14910);
xnor U15096 (N_15096,N_14275,N_14333);
xnor U15097 (N_15097,N_14830,N_14492);
nand U15098 (N_15098,N_14516,N_14100);
nand U15099 (N_15099,N_14026,N_14202);
xor U15100 (N_15100,N_14640,N_14645);
or U15101 (N_15101,N_14634,N_14095);
nand U15102 (N_15102,N_14879,N_14194);
and U15103 (N_15103,N_14140,N_14570);
or U15104 (N_15104,N_14153,N_14049);
and U15105 (N_15105,N_14097,N_14825);
and U15106 (N_15106,N_14304,N_14860);
nor U15107 (N_15107,N_14139,N_14032);
nand U15108 (N_15108,N_14008,N_14951);
xnor U15109 (N_15109,N_14596,N_14236);
xnor U15110 (N_15110,N_14465,N_14030);
xnor U15111 (N_15111,N_14173,N_14833);
xor U15112 (N_15112,N_14997,N_14456);
nor U15113 (N_15113,N_14016,N_14295);
or U15114 (N_15114,N_14351,N_14573);
nor U15115 (N_15115,N_14502,N_14408);
nand U15116 (N_15116,N_14190,N_14963);
nand U15117 (N_15117,N_14401,N_14940);
nor U15118 (N_15118,N_14978,N_14042);
or U15119 (N_15119,N_14850,N_14650);
nor U15120 (N_15120,N_14553,N_14654);
xnor U15121 (N_15121,N_14218,N_14223);
nand U15122 (N_15122,N_14728,N_14558);
xnor U15123 (N_15123,N_14835,N_14648);
xnor U15124 (N_15124,N_14729,N_14402);
nor U15125 (N_15125,N_14968,N_14497);
or U15126 (N_15126,N_14617,N_14157);
or U15127 (N_15127,N_14945,N_14667);
xnor U15128 (N_15128,N_14858,N_14473);
xor U15129 (N_15129,N_14433,N_14006);
nand U15130 (N_15130,N_14046,N_14601);
xnor U15131 (N_15131,N_14054,N_14000);
and U15132 (N_15132,N_14585,N_14717);
xor U15133 (N_15133,N_14791,N_14746);
or U15134 (N_15134,N_14893,N_14944);
nor U15135 (N_15135,N_14819,N_14615);
and U15136 (N_15136,N_14110,N_14439);
nor U15137 (N_15137,N_14081,N_14301);
xor U15138 (N_15138,N_14498,N_14916);
and U15139 (N_15139,N_14271,N_14028);
xor U15140 (N_15140,N_14990,N_14364);
xnor U15141 (N_15141,N_14760,N_14486);
and U15142 (N_15142,N_14774,N_14821);
and U15143 (N_15143,N_14614,N_14009);
nand U15144 (N_15144,N_14407,N_14923);
xor U15145 (N_15145,N_14321,N_14372);
and U15146 (N_15146,N_14785,N_14924);
xor U15147 (N_15147,N_14711,N_14909);
nor U15148 (N_15148,N_14180,N_14960);
nand U15149 (N_15149,N_14464,N_14434);
xnor U15150 (N_15150,N_14929,N_14643);
and U15151 (N_15151,N_14149,N_14841);
xor U15152 (N_15152,N_14685,N_14504);
nand U15153 (N_15153,N_14797,N_14286);
xnor U15154 (N_15154,N_14158,N_14423);
and U15155 (N_15155,N_14957,N_14519);
and U15156 (N_15156,N_14219,N_14613);
nand U15157 (N_15157,N_14023,N_14851);
xnor U15158 (N_15158,N_14975,N_14175);
xnor U15159 (N_15159,N_14561,N_14946);
and U15160 (N_15160,N_14619,N_14466);
xor U15161 (N_15161,N_14602,N_14253);
xnor U15162 (N_15162,N_14133,N_14903);
nand U15163 (N_15163,N_14693,N_14802);
nand U15164 (N_15164,N_14378,N_14953);
nor U15165 (N_15165,N_14469,N_14775);
and U15166 (N_15166,N_14328,N_14096);
or U15167 (N_15167,N_14954,N_14047);
and U15168 (N_15168,N_14652,N_14297);
xor U15169 (N_15169,N_14155,N_14943);
nor U15170 (N_15170,N_14528,N_14307);
nand U15171 (N_15171,N_14994,N_14868);
and U15172 (N_15172,N_14735,N_14078);
and U15173 (N_15173,N_14457,N_14192);
nand U15174 (N_15174,N_14085,N_14151);
nor U15175 (N_15175,N_14826,N_14162);
nor U15176 (N_15176,N_14059,N_14368);
xnor U15177 (N_15177,N_14988,N_14201);
or U15178 (N_15178,N_14288,N_14416);
nor U15179 (N_15179,N_14291,N_14554);
nand U15180 (N_15180,N_14754,N_14138);
and U15181 (N_15181,N_14327,N_14279);
or U15182 (N_15182,N_14885,N_14126);
or U15183 (N_15183,N_14418,N_14273);
or U15184 (N_15184,N_14232,N_14984);
nand U15185 (N_15185,N_14744,N_14845);
nor U15186 (N_15186,N_14673,N_14567);
xnor U15187 (N_15187,N_14934,N_14672);
nor U15188 (N_15188,N_14107,N_14130);
or U15189 (N_15189,N_14217,N_14471);
nand U15190 (N_15190,N_14228,N_14890);
nand U15191 (N_15191,N_14427,N_14598);
and U15192 (N_15192,N_14914,N_14323);
nor U15193 (N_15193,N_14413,N_14816);
xnor U15194 (N_15194,N_14022,N_14680);
nand U15195 (N_15195,N_14296,N_14781);
and U15196 (N_15196,N_14355,N_14702);
and U15197 (N_15197,N_14369,N_14114);
or U15198 (N_15198,N_14250,N_14973);
and U15199 (N_15199,N_14302,N_14512);
nand U15200 (N_15200,N_14445,N_14161);
nor U15201 (N_15201,N_14737,N_14533);
nand U15202 (N_15202,N_14277,N_14993);
and U15203 (N_15203,N_14808,N_14531);
and U15204 (N_15204,N_14779,N_14560);
xnor U15205 (N_15205,N_14952,N_14991);
xnor U15206 (N_15206,N_14257,N_14552);
nor U15207 (N_15207,N_14393,N_14320);
xnor U15208 (N_15208,N_14391,N_14677);
nor U15209 (N_15209,N_14790,N_14181);
xnor U15210 (N_15210,N_14818,N_14638);
or U15211 (N_15211,N_14964,N_14623);
or U15212 (N_15212,N_14144,N_14390);
and U15213 (N_15213,N_14678,N_14691);
xnor U15214 (N_15214,N_14429,N_14641);
and U15215 (N_15215,N_14145,N_14747);
and U15216 (N_15216,N_14420,N_14484);
xnor U15217 (N_15217,N_14542,N_14244);
or U15218 (N_15218,N_14783,N_14255);
xor U15219 (N_15219,N_14911,N_14050);
or U15220 (N_15220,N_14524,N_14629);
and U15221 (N_15221,N_14463,N_14170);
nor U15222 (N_15222,N_14592,N_14756);
nand U15223 (N_15223,N_14319,N_14937);
nor U15224 (N_15224,N_14018,N_14712);
nand U15225 (N_15225,N_14003,N_14545);
nor U15226 (N_15226,N_14451,N_14125);
nand U15227 (N_15227,N_14537,N_14058);
nor U15228 (N_15228,N_14844,N_14156);
or U15229 (N_15229,N_14460,N_14905);
and U15230 (N_15230,N_14185,N_14986);
nor U15231 (N_15231,N_14143,N_14398);
xor U15232 (N_15232,N_14315,N_14132);
xnor U15233 (N_15233,N_14285,N_14290);
nand U15234 (N_15234,N_14483,N_14071);
and U15235 (N_15235,N_14091,N_14772);
nor U15236 (N_15236,N_14718,N_14662);
nor U15237 (N_15237,N_14350,N_14448);
or U15238 (N_15238,N_14383,N_14777);
or U15239 (N_15239,N_14316,N_14246);
nand U15240 (N_15240,N_14400,N_14740);
xnor U15241 (N_15241,N_14251,N_14699);
and U15242 (N_15242,N_14814,N_14900);
xor U15243 (N_15243,N_14608,N_14266);
or U15244 (N_15244,N_14012,N_14690);
nand U15245 (N_15245,N_14247,N_14043);
nand U15246 (N_15246,N_14949,N_14005);
or U15247 (N_15247,N_14931,N_14588);
or U15248 (N_15248,N_14878,N_14809);
xor U15249 (N_15249,N_14041,N_14090);
and U15250 (N_15250,N_14122,N_14532);
nor U15251 (N_15251,N_14587,N_14204);
nor U15252 (N_15252,N_14800,N_14189);
nand U15253 (N_15253,N_14222,N_14888);
nor U15254 (N_15254,N_14123,N_14015);
or U15255 (N_15255,N_14751,N_14356);
nand U15256 (N_15256,N_14723,N_14063);
nand U15257 (N_15257,N_14543,N_14238);
nor U15258 (N_15258,N_14568,N_14891);
xnor U15259 (N_15259,N_14622,N_14551);
xor U15260 (N_15260,N_14621,N_14211);
or U15261 (N_15261,N_14184,N_14045);
nand U15262 (N_15262,N_14792,N_14987);
nand U15263 (N_15263,N_14264,N_14971);
nand U15264 (N_15264,N_14007,N_14876);
nor U15265 (N_15265,N_14942,N_14507);
or U15266 (N_15266,N_14763,N_14713);
nor U15267 (N_15267,N_14104,N_14761);
nor U15268 (N_15268,N_14405,N_14415);
or U15269 (N_15269,N_14983,N_14245);
nor U15270 (N_15270,N_14472,N_14523);
and U15271 (N_15271,N_14013,N_14021);
nor U15272 (N_15272,N_14256,N_14334);
nand U15273 (N_15273,N_14762,N_14267);
or U15274 (N_15274,N_14010,N_14075);
and U15275 (N_15275,N_14787,N_14730);
or U15276 (N_15276,N_14443,N_14293);
xor U15277 (N_15277,N_14660,N_14578);
xnor U15278 (N_15278,N_14135,N_14426);
nand U15279 (N_15279,N_14292,N_14912);
or U15280 (N_15280,N_14020,N_14438);
and U15281 (N_15281,N_14628,N_14159);
nor U15282 (N_15282,N_14546,N_14169);
or U15283 (N_15283,N_14842,N_14789);
nand U15284 (N_15284,N_14102,N_14033);
or U15285 (N_15285,N_14778,N_14115);
nand U15286 (N_15286,N_14630,N_14877);
xnor U15287 (N_15287,N_14425,N_14659);
nand U15288 (N_15288,N_14859,N_14379);
or U15289 (N_15289,N_14265,N_14057);
and U15290 (N_15290,N_14521,N_14481);
nor U15291 (N_15291,N_14233,N_14128);
nand U15292 (N_15292,N_14146,N_14499);
and U15293 (N_15293,N_14739,N_14855);
or U15294 (N_15294,N_14846,N_14708);
nand U15295 (N_15295,N_14575,N_14919);
nor U15296 (N_15296,N_14331,N_14208);
or U15297 (N_15297,N_14225,N_14626);
nor U15298 (N_15298,N_14881,N_14611);
or U15299 (N_15299,N_14874,N_14930);
xnor U15300 (N_15300,N_14589,N_14653);
and U15301 (N_15301,N_14177,N_14593);
and U15302 (N_15302,N_14452,N_14639);
nand U15303 (N_15303,N_14773,N_14313);
nor U15304 (N_15304,N_14925,N_14674);
or U15305 (N_15305,N_14679,N_14666);
and U15306 (N_15306,N_14741,N_14616);
nor U15307 (N_15307,N_14458,N_14303);
and U15308 (N_15308,N_14476,N_14113);
xnor U15309 (N_15309,N_14834,N_14029);
or U15310 (N_15310,N_14127,N_14396);
nor U15311 (N_15311,N_14958,N_14815);
nor U15312 (N_15312,N_14406,N_14707);
or U15313 (N_15313,N_14371,N_14182);
or U15314 (N_15314,N_14394,N_14093);
and U15315 (N_15315,N_14430,N_14557);
nor U15316 (N_15316,N_14928,N_14820);
nand U15317 (N_15317,N_14280,N_14366);
or U15318 (N_15318,N_14506,N_14178);
or U15319 (N_15319,N_14482,N_14387);
nand U15320 (N_15320,N_14642,N_14875);
nand U15321 (N_15321,N_14547,N_14160);
or U15322 (N_15322,N_14510,N_14088);
xnor U15323 (N_15323,N_14681,N_14376);
nor U15324 (N_15324,N_14348,N_14590);
nor U15325 (N_15325,N_14335,N_14727);
nand U15326 (N_15326,N_14444,N_14969);
and U15327 (N_15327,N_14695,N_14154);
and U15328 (N_15328,N_14716,N_14210);
and U15329 (N_15329,N_14134,N_14237);
and U15330 (N_15330,N_14254,N_14966);
nor U15331 (N_15331,N_14530,N_14262);
xor U15332 (N_15332,N_14048,N_14522);
nor U15333 (N_15333,N_14431,N_14311);
nand U15334 (N_15334,N_14437,N_14065);
and U15335 (N_15335,N_14207,N_14584);
nand U15336 (N_15336,N_14474,N_14795);
nand U15337 (N_15337,N_14019,N_14804);
xnor U15338 (N_15338,N_14440,N_14241);
nand U15339 (N_15339,N_14535,N_14668);
and U15340 (N_15340,N_14603,N_14347);
xor U15341 (N_15341,N_14105,N_14329);
xnor U15342 (N_15342,N_14705,N_14907);
xnor U15343 (N_15343,N_14947,N_14594);
and U15344 (N_15344,N_14866,N_14004);
and U15345 (N_15345,N_14768,N_14487);
nor U15346 (N_15346,N_14574,N_14282);
or U15347 (N_15347,N_14962,N_14827);
nand U15348 (N_15348,N_14698,N_14252);
or U15349 (N_15349,N_14141,N_14597);
nor U15350 (N_15350,N_14508,N_14166);
nand U15351 (N_15351,N_14395,N_14388);
nor U15352 (N_15352,N_14308,N_14897);
or U15353 (N_15353,N_14899,N_14577);
xnor U15354 (N_15354,N_14817,N_14360);
or U15355 (N_15355,N_14035,N_14209);
and U15356 (N_15356,N_14520,N_14509);
nand U15357 (N_15357,N_14664,N_14336);
xor U15358 (N_15358,N_14541,N_14870);
or U15359 (N_15359,N_14011,N_14788);
and U15360 (N_15360,N_14345,N_14724);
nand U15361 (N_15361,N_14357,N_14129);
and U15362 (N_15362,N_14205,N_14260);
nor U15363 (N_15363,N_14769,N_14722);
or U15364 (N_15364,N_14089,N_14411);
or U15365 (N_15365,N_14142,N_14927);
nand U15366 (N_15366,N_14432,N_14961);
nor U15367 (N_15367,N_14461,N_14467);
or U15368 (N_15368,N_14956,N_14488);
nand U15369 (N_15369,N_14039,N_14073);
nand U15370 (N_15370,N_14872,N_14950);
nor U15371 (N_15371,N_14555,N_14014);
nor U15372 (N_15372,N_14556,N_14871);
or U15373 (N_15373,N_14811,N_14995);
nor U15374 (N_15374,N_14338,N_14922);
or U15375 (N_15375,N_14749,N_14414);
or U15376 (N_15376,N_14714,N_14981);
nand U15377 (N_15377,N_14342,N_14583);
and U15378 (N_15378,N_14197,N_14736);
and U15379 (N_15379,N_14700,N_14098);
nand U15380 (N_15380,N_14548,N_14188);
nor U15381 (N_15381,N_14848,N_14500);
nand U15382 (N_15382,N_14972,N_14397);
or U15383 (N_15383,N_14309,N_14212);
xor U15384 (N_15384,N_14889,N_14136);
nand U15385 (N_15385,N_14417,N_14805);
nand U15386 (N_15386,N_14036,N_14892);
and U15387 (N_15387,N_14726,N_14111);
xor U15388 (N_15388,N_14243,N_14268);
and U15389 (N_15389,N_14579,N_14261);
nor U15390 (N_15390,N_14447,N_14353);
xor U15391 (N_15391,N_14119,N_14689);
nor U15392 (N_15392,N_14027,N_14517);
xor U15393 (N_15393,N_14663,N_14665);
nor U15394 (N_15394,N_14441,N_14600);
nand U15395 (N_15395,N_14852,N_14403);
nand U15396 (N_15396,N_14226,N_14683);
or U15397 (N_15397,N_14346,N_14959);
nor U15398 (N_15398,N_14116,N_14479);
nor U15399 (N_15399,N_14936,N_14470);
nor U15400 (N_15400,N_14455,N_14806);
or U15401 (N_15401,N_14227,N_14040);
and U15402 (N_15402,N_14263,N_14687);
nor U15403 (N_15403,N_14658,N_14733);
nand U15404 (N_15404,N_14239,N_14822);
xor U15405 (N_15405,N_14475,N_14220);
xnor U15406 (N_15406,N_14782,N_14801);
nand U15407 (N_15407,N_14813,N_14099);
and U15408 (N_15408,N_14974,N_14191);
or U15409 (N_15409,N_14832,N_14435);
or U15410 (N_15410,N_14174,N_14365);
and U15411 (N_15411,N_14074,N_14527);
or U15412 (N_15412,N_14501,N_14215);
xor U15413 (N_15413,N_14938,N_14843);
nor U15414 (N_15414,N_14534,N_14620);
nor U15415 (N_15415,N_14780,N_14106);
xor U15416 (N_15416,N_14646,N_14591);
xnor U15417 (N_15417,N_14837,N_14609);
nand U15418 (N_15418,N_14373,N_14055);
and U15419 (N_15419,N_14478,N_14358);
and U15420 (N_15420,N_14539,N_14840);
and U15421 (N_15421,N_14234,N_14287);
xor U15422 (N_15422,N_14884,N_14701);
or U15423 (N_15423,N_14670,N_14569);
nor U15424 (N_15424,N_14310,N_14001);
nand U15425 (N_15425,N_14576,N_14515);
nand U15426 (N_15426,N_14908,N_14453);
or U15427 (N_15427,N_14038,N_14200);
or U15428 (N_15428,N_14526,N_14272);
nor U15429 (N_15429,N_14536,N_14199);
and U15430 (N_15430,N_14249,N_14124);
or U15431 (N_15431,N_14454,N_14828);
and U15432 (N_15432,N_14318,N_14203);
xnor U15433 (N_15433,N_14332,N_14240);
and U15434 (N_15434,N_14108,N_14352);
nor U15435 (N_15435,N_14051,N_14325);
and U15436 (N_15436,N_14242,N_14970);
or U15437 (N_15437,N_14867,N_14339);
nor U15438 (N_15438,N_14362,N_14998);
nor U15439 (N_15439,N_14354,N_14915);
and U15440 (N_15440,N_14743,N_14661);
nand U15441 (N_15441,N_14599,N_14807);
nor U15442 (N_15442,N_14305,N_14625);
and U15443 (N_15443,N_14216,N_14776);
nand U15444 (N_15444,N_14034,N_14306);
nand U15445 (N_15445,N_14083,N_14392);
xor U15446 (N_15446,N_14770,N_14230);
nand U15447 (N_15447,N_14076,N_14857);
or U15448 (N_15448,N_14513,N_14077);
or U15449 (N_15449,N_14385,N_14798);
or U15450 (N_15450,N_14384,N_14326);
nor U15451 (N_15451,N_14967,N_14442);
xnor U15452 (N_15452,N_14586,N_14300);
or U15453 (N_15453,N_14734,N_14382);
and U15454 (N_15454,N_14080,N_14061);
or U15455 (N_15455,N_14880,N_14644);
or U15456 (N_15456,N_14562,N_14686);
and U15457 (N_15457,N_14086,N_14314);
nor U15458 (N_15458,N_14886,N_14064);
xor U15459 (N_15459,N_14985,N_14152);
or U15460 (N_15460,N_14289,N_14649);
or U15461 (N_15461,N_14495,N_14363);
and U15462 (N_15462,N_14709,N_14380);
or U15463 (N_15463,N_14377,N_14094);
or U15464 (N_15464,N_14317,N_14823);
xor U15465 (N_15465,N_14655,N_14206);
or U15466 (N_15466,N_14902,N_14168);
and U15467 (N_15467,N_14996,N_14404);
xnor U15468 (N_15468,N_14084,N_14450);
nor U15469 (N_15469,N_14367,N_14067);
and U15470 (N_15470,N_14494,N_14581);
or U15471 (N_15471,N_14854,N_14894);
xor U15472 (N_15472,N_14651,N_14213);
or U15473 (N_15473,N_14370,N_14710);
xnor U15474 (N_15474,N_14836,N_14939);
and U15475 (N_15475,N_14299,N_14544);
and U15476 (N_15476,N_14278,N_14410);
nand U15477 (N_15477,N_14118,N_14607);
or U15478 (N_15478,N_14853,N_14349);
xnor U15479 (N_15479,N_14221,N_14904);
and U15480 (N_15480,N_14229,N_14112);
xor U15481 (N_15481,N_14935,N_14485);
nor U15482 (N_15482,N_14269,N_14771);
nand U15483 (N_15483,N_14066,N_14359);
nor U15484 (N_15484,N_14496,N_14595);
nand U15485 (N_15485,N_14753,N_14684);
nand U15486 (N_15486,N_14918,N_14409);
or U15487 (N_15487,N_14631,N_14856);
nor U15488 (N_15488,N_14459,N_14214);
xor U15489 (N_15489,N_14610,N_14550);
and U15490 (N_15490,N_14424,N_14932);
xnor U15491 (N_15491,N_14571,N_14002);
xnor U15492 (N_15492,N_14092,N_14920);
xor U15493 (N_15493,N_14193,N_14381);
or U15494 (N_15494,N_14163,N_14069);
nand U15495 (N_15495,N_14605,N_14164);
or U15496 (N_15496,N_14165,N_14784);
or U15497 (N_15497,N_14053,N_14906);
nor U15498 (N_15498,N_14566,N_14704);
or U15499 (N_15499,N_14511,N_14131);
nor U15500 (N_15500,N_14449,N_14864);
nand U15501 (N_15501,N_14967,N_14112);
nand U15502 (N_15502,N_14350,N_14723);
nor U15503 (N_15503,N_14713,N_14338);
xnor U15504 (N_15504,N_14968,N_14966);
or U15505 (N_15505,N_14695,N_14531);
or U15506 (N_15506,N_14042,N_14011);
and U15507 (N_15507,N_14601,N_14918);
or U15508 (N_15508,N_14196,N_14820);
or U15509 (N_15509,N_14329,N_14368);
nor U15510 (N_15510,N_14929,N_14168);
nor U15511 (N_15511,N_14567,N_14022);
xnor U15512 (N_15512,N_14158,N_14683);
xor U15513 (N_15513,N_14855,N_14780);
xor U15514 (N_15514,N_14729,N_14216);
xnor U15515 (N_15515,N_14318,N_14726);
or U15516 (N_15516,N_14080,N_14024);
nand U15517 (N_15517,N_14521,N_14143);
or U15518 (N_15518,N_14862,N_14150);
or U15519 (N_15519,N_14498,N_14828);
xor U15520 (N_15520,N_14031,N_14380);
xnor U15521 (N_15521,N_14668,N_14253);
nand U15522 (N_15522,N_14281,N_14291);
nor U15523 (N_15523,N_14851,N_14980);
nor U15524 (N_15524,N_14887,N_14672);
xnor U15525 (N_15525,N_14068,N_14232);
and U15526 (N_15526,N_14119,N_14893);
or U15527 (N_15527,N_14529,N_14611);
nor U15528 (N_15528,N_14756,N_14451);
xor U15529 (N_15529,N_14312,N_14390);
or U15530 (N_15530,N_14556,N_14968);
nand U15531 (N_15531,N_14764,N_14454);
and U15532 (N_15532,N_14312,N_14035);
or U15533 (N_15533,N_14749,N_14090);
and U15534 (N_15534,N_14473,N_14212);
nand U15535 (N_15535,N_14285,N_14820);
nand U15536 (N_15536,N_14135,N_14698);
nor U15537 (N_15537,N_14459,N_14667);
xnor U15538 (N_15538,N_14605,N_14822);
xnor U15539 (N_15539,N_14323,N_14283);
and U15540 (N_15540,N_14072,N_14946);
nand U15541 (N_15541,N_14848,N_14126);
nand U15542 (N_15542,N_14216,N_14936);
and U15543 (N_15543,N_14003,N_14438);
or U15544 (N_15544,N_14996,N_14084);
and U15545 (N_15545,N_14834,N_14471);
nand U15546 (N_15546,N_14951,N_14934);
or U15547 (N_15547,N_14788,N_14905);
or U15548 (N_15548,N_14107,N_14569);
nand U15549 (N_15549,N_14342,N_14869);
nand U15550 (N_15550,N_14311,N_14252);
nand U15551 (N_15551,N_14997,N_14036);
nor U15552 (N_15552,N_14985,N_14651);
nand U15553 (N_15553,N_14083,N_14831);
xnor U15554 (N_15554,N_14426,N_14606);
xnor U15555 (N_15555,N_14208,N_14735);
nand U15556 (N_15556,N_14057,N_14091);
and U15557 (N_15557,N_14717,N_14256);
or U15558 (N_15558,N_14560,N_14801);
nor U15559 (N_15559,N_14066,N_14264);
or U15560 (N_15560,N_14726,N_14226);
xor U15561 (N_15561,N_14471,N_14406);
nor U15562 (N_15562,N_14899,N_14428);
nor U15563 (N_15563,N_14093,N_14883);
xnor U15564 (N_15564,N_14648,N_14846);
and U15565 (N_15565,N_14214,N_14809);
and U15566 (N_15566,N_14621,N_14431);
and U15567 (N_15567,N_14443,N_14877);
or U15568 (N_15568,N_14409,N_14100);
and U15569 (N_15569,N_14071,N_14664);
and U15570 (N_15570,N_14379,N_14858);
and U15571 (N_15571,N_14345,N_14697);
nor U15572 (N_15572,N_14366,N_14242);
nor U15573 (N_15573,N_14513,N_14483);
xnor U15574 (N_15574,N_14719,N_14614);
and U15575 (N_15575,N_14220,N_14218);
and U15576 (N_15576,N_14491,N_14423);
and U15577 (N_15577,N_14900,N_14893);
nand U15578 (N_15578,N_14755,N_14222);
and U15579 (N_15579,N_14252,N_14219);
nor U15580 (N_15580,N_14766,N_14545);
or U15581 (N_15581,N_14893,N_14454);
or U15582 (N_15582,N_14818,N_14902);
or U15583 (N_15583,N_14976,N_14003);
or U15584 (N_15584,N_14878,N_14596);
xnor U15585 (N_15585,N_14720,N_14572);
nand U15586 (N_15586,N_14025,N_14076);
nand U15587 (N_15587,N_14774,N_14420);
or U15588 (N_15588,N_14892,N_14073);
and U15589 (N_15589,N_14683,N_14880);
or U15590 (N_15590,N_14711,N_14443);
nand U15591 (N_15591,N_14698,N_14518);
and U15592 (N_15592,N_14879,N_14326);
and U15593 (N_15593,N_14773,N_14415);
nand U15594 (N_15594,N_14558,N_14914);
and U15595 (N_15595,N_14668,N_14633);
xnor U15596 (N_15596,N_14096,N_14320);
or U15597 (N_15597,N_14866,N_14432);
xor U15598 (N_15598,N_14801,N_14742);
nor U15599 (N_15599,N_14217,N_14106);
nor U15600 (N_15600,N_14503,N_14776);
and U15601 (N_15601,N_14827,N_14239);
and U15602 (N_15602,N_14367,N_14657);
nor U15603 (N_15603,N_14652,N_14228);
xor U15604 (N_15604,N_14688,N_14620);
nor U15605 (N_15605,N_14736,N_14112);
or U15606 (N_15606,N_14569,N_14343);
or U15607 (N_15607,N_14803,N_14517);
nor U15608 (N_15608,N_14692,N_14694);
or U15609 (N_15609,N_14943,N_14001);
or U15610 (N_15610,N_14321,N_14476);
nand U15611 (N_15611,N_14665,N_14493);
nor U15612 (N_15612,N_14112,N_14431);
nand U15613 (N_15613,N_14399,N_14300);
xor U15614 (N_15614,N_14625,N_14615);
or U15615 (N_15615,N_14360,N_14208);
nand U15616 (N_15616,N_14714,N_14328);
or U15617 (N_15617,N_14261,N_14835);
and U15618 (N_15618,N_14318,N_14299);
nor U15619 (N_15619,N_14186,N_14830);
and U15620 (N_15620,N_14752,N_14411);
nand U15621 (N_15621,N_14556,N_14960);
nor U15622 (N_15622,N_14963,N_14037);
and U15623 (N_15623,N_14059,N_14969);
or U15624 (N_15624,N_14323,N_14699);
nand U15625 (N_15625,N_14386,N_14391);
xor U15626 (N_15626,N_14268,N_14682);
and U15627 (N_15627,N_14551,N_14708);
nand U15628 (N_15628,N_14001,N_14229);
or U15629 (N_15629,N_14266,N_14789);
or U15630 (N_15630,N_14527,N_14160);
or U15631 (N_15631,N_14344,N_14859);
xor U15632 (N_15632,N_14123,N_14710);
nand U15633 (N_15633,N_14091,N_14997);
nor U15634 (N_15634,N_14982,N_14003);
xor U15635 (N_15635,N_14363,N_14135);
nand U15636 (N_15636,N_14904,N_14656);
or U15637 (N_15637,N_14727,N_14824);
nand U15638 (N_15638,N_14241,N_14028);
or U15639 (N_15639,N_14293,N_14012);
or U15640 (N_15640,N_14910,N_14513);
and U15641 (N_15641,N_14113,N_14429);
nand U15642 (N_15642,N_14238,N_14126);
or U15643 (N_15643,N_14412,N_14918);
xnor U15644 (N_15644,N_14586,N_14480);
xnor U15645 (N_15645,N_14771,N_14663);
and U15646 (N_15646,N_14371,N_14529);
nand U15647 (N_15647,N_14664,N_14800);
or U15648 (N_15648,N_14509,N_14980);
nor U15649 (N_15649,N_14856,N_14889);
nor U15650 (N_15650,N_14644,N_14004);
and U15651 (N_15651,N_14073,N_14141);
and U15652 (N_15652,N_14879,N_14289);
nand U15653 (N_15653,N_14167,N_14819);
and U15654 (N_15654,N_14489,N_14909);
xnor U15655 (N_15655,N_14558,N_14534);
xnor U15656 (N_15656,N_14637,N_14518);
xor U15657 (N_15657,N_14569,N_14491);
nand U15658 (N_15658,N_14431,N_14594);
nor U15659 (N_15659,N_14401,N_14742);
xnor U15660 (N_15660,N_14085,N_14247);
or U15661 (N_15661,N_14035,N_14279);
nor U15662 (N_15662,N_14793,N_14807);
nand U15663 (N_15663,N_14790,N_14851);
and U15664 (N_15664,N_14596,N_14131);
nor U15665 (N_15665,N_14597,N_14900);
or U15666 (N_15666,N_14601,N_14473);
or U15667 (N_15667,N_14443,N_14499);
nand U15668 (N_15668,N_14608,N_14892);
and U15669 (N_15669,N_14579,N_14885);
nand U15670 (N_15670,N_14213,N_14446);
xnor U15671 (N_15671,N_14281,N_14855);
xnor U15672 (N_15672,N_14908,N_14318);
nor U15673 (N_15673,N_14558,N_14452);
nand U15674 (N_15674,N_14298,N_14177);
nand U15675 (N_15675,N_14098,N_14386);
and U15676 (N_15676,N_14428,N_14169);
xnor U15677 (N_15677,N_14249,N_14264);
nand U15678 (N_15678,N_14870,N_14142);
nand U15679 (N_15679,N_14689,N_14447);
nand U15680 (N_15680,N_14324,N_14340);
or U15681 (N_15681,N_14565,N_14230);
and U15682 (N_15682,N_14654,N_14623);
xnor U15683 (N_15683,N_14624,N_14999);
nor U15684 (N_15684,N_14963,N_14283);
and U15685 (N_15685,N_14555,N_14678);
nand U15686 (N_15686,N_14607,N_14608);
xnor U15687 (N_15687,N_14581,N_14075);
or U15688 (N_15688,N_14372,N_14508);
or U15689 (N_15689,N_14257,N_14635);
nand U15690 (N_15690,N_14539,N_14704);
and U15691 (N_15691,N_14878,N_14843);
nand U15692 (N_15692,N_14110,N_14153);
nor U15693 (N_15693,N_14422,N_14791);
or U15694 (N_15694,N_14734,N_14585);
and U15695 (N_15695,N_14935,N_14255);
xor U15696 (N_15696,N_14811,N_14088);
and U15697 (N_15697,N_14134,N_14100);
nor U15698 (N_15698,N_14155,N_14755);
and U15699 (N_15699,N_14244,N_14184);
nand U15700 (N_15700,N_14512,N_14920);
xnor U15701 (N_15701,N_14619,N_14046);
or U15702 (N_15702,N_14938,N_14587);
or U15703 (N_15703,N_14025,N_14597);
or U15704 (N_15704,N_14223,N_14250);
and U15705 (N_15705,N_14204,N_14194);
and U15706 (N_15706,N_14659,N_14176);
and U15707 (N_15707,N_14540,N_14359);
nor U15708 (N_15708,N_14064,N_14761);
nor U15709 (N_15709,N_14278,N_14987);
or U15710 (N_15710,N_14676,N_14825);
or U15711 (N_15711,N_14281,N_14374);
nand U15712 (N_15712,N_14965,N_14711);
or U15713 (N_15713,N_14280,N_14499);
and U15714 (N_15714,N_14854,N_14579);
nand U15715 (N_15715,N_14404,N_14365);
xnor U15716 (N_15716,N_14712,N_14176);
nand U15717 (N_15717,N_14976,N_14636);
and U15718 (N_15718,N_14966,N_14962);
nand U15719 (N_15719,N_14209,N_14310);
nand U15720 (N_15720,N_14023,N_14252);
or U15721 (N_15721,N_14554,N_14464);
nand U15722 (N_15722,N_14264,N_14228);
nand U15723 (N_15723,N_14698,N_14120);
nor U15724 (N_15724,N_14484,N_14049);
nor U15725 (N_15725,N_14500,N_14838);
or U15726 (N_15726,N_14894,N_14402);
and U15727 (N_15727,N_14060,N_14201);
or U15728 (N_15728,N_14058,N_14170);
or U15729 (N_15729,N_14158,N_14690);
nand U15730 (N_15730,N_14088,N_14574);
and U15731 (N_15731,N_14935,N_14572);
and U15732 (N_15732,N_14306,N_14721);
nor U15733 (N_15733,N_14301,N_14439);
or U15734 (N_15734,N_14359,N_14566);
nand U15735 (N_15735,N_14405,N_14610);
xor U15736 (N_15736,N_14429,N_14970);
xnor U15737 (N_15737,N_14995,N_14989);
xnor U15738 (N_15738,N_14865,N_14022);
and U15739 (N_15739,N_14886,N_14915);
or U15740 (N_15740,N_14914,N_14136);
or U15741 (N_15741,N_14196,N_14971);
and U15742 (N_15742,N_14259,N_14108);
and U15743 (N_15743,N_14773,N_14890);
and U15744 (N_15744,N_14799,N_14899);
and U15745 (N_15745,N_14355,N_14653);
or U15746 (N_15746,N_14084,N_14562);
or U15747 (N_15747,N_14318,N_14914);
and U15748 (N_15748,N_14043,N_14744);
and U15749 (N_15749,N_14748,N_14711);
xor U15750 (N_15750,N_14371,N_14092);
nand U15751 (N_15751,N_14084,N_14031);
nand U15752 (N_15752,N_14684,N_14878);
nor U15753 (N_15753,N_14821,N_14847);
xnor U15754 (N_15754,N_14963,N_14321);
or U15755 (N_15755,N_14972,N_14672);
and U15756 (N_15756,N_14960,N_14464);
and U15757 (N_15757,N_14327,N_14767);
nand U15758 (N_15758,N_14356,N_14615);
and U15759 (N_15759,N_14285,N_14681);
nand U15760 (N_15760,N_14139,N_14252);
nand U15761 (N_15761,N_14344,N_14752);
xnor U15762 (N_15762,N_14958,N_14007);
and U15763 (N_15763,N_14234,N_14913);
xnor U15764 (N_15764,N_14081,N_14641);
nand U15765 (N_15765,N_14733,N_14527);
nand U15766 (N_15766,N_14907,N_14839);
nor U15767 (N_15767,N_14372,N_14831);
or U15768 (N_15768,N_14253,N_14644);
xor U15769 (N_15769,N_14388,N_14358);
and U15770 (N_15770,N_14347,N_14494);
and U15771 (N_15771,N_14521,N_14236);
nand U15772 (N_15772,N_14961,N_14969);
nand U15773 (N_15773,N_14969,N_14405);
and U15774 (N_15774,N_14119,N_14605);
and U15775 (N_15775,N_14616,N_14842);
and U15776 (N_15776,N_14014,N_14600);
xor U15777 (N_15777,N_14065,N_14479);
and U15778 (N_15778,N_14458,N_14625);
nand U15779 (N_15779,N_14227,N_14142);
and U15780 (N_15780,N_14093,N_14534);
nor U15781 (N_15781,N_14692,N_14125);
or U15782 (N_15782,N_14254,N_14843);
nor U15783 (N_15783,N_14166,N_14577);
and U15784 (N_15784,N_14121,N_14425);
nand U15785 (N_15785,N_14743,N_14210);
xnor U15786 (N_15786,N_14162,N_14638);
nand U15787 (N_15787,N_14300,N_14598);
xor U15788 (N_15788,N_14052,N_14800);
nand U15789 (N_15789,N_14570,N_14417);
nor U15790 (N_15790,N_14694,N_14982);
or U15791 (N_15791,N_14660,N_14750);
nor U15792 (N_15792,N_14239,N_14954);
nor U15793 (N_15793,N_14775,N_14127);
xnor U15794 (N_15794,N_14406,N_14281);
and U15795 (N_15795,N_14490,N_14081);
nand U15796 (N_15796,N_14630,N_14369);
or U15797 (N_15797,N_14949,N_14872);
and U15798 (N_15798,N_14155,N_14940);
nand U15799 (N_15799,N_14232,N_14445);
or U15800 (N_15800,N_14282,N_14178);
or U15801 (N_15801,N_14045,N_14961);
xnor U15802 (N_15802,N_14004,N_14127);
nor U15803 (N_15803,N_14937,N_14388);
nor U15804 (N_15804,N_14582,N_14491);
nor U15805 (N_15805,N_14897,N_14840);
or U15806 (N_15806,N_14549,N_14494);
nor U15807 (N_15807,N_14318,N_14502);
xor U15808 (N_15808,N_14358,N_14574);
and U15809 (N_15809,N_14729,N_14202);
nor U15810 (N_15810,N_14264,N_14061);
or U15811 (N_15811,N_14329,N_14970);
xor U15812 (N_15812,N_14441,N_14985);
xor U15813 (N_15813,N_14217,N_14712);
xnor U15814 (N_15814,N_14649,N_14870);
xnor U15815 (N_15815,N_14675,N_14517);
nand U15816 (N_15816,N_14757,N_14554);
nand U15817 (N_15817,N_14642,N_14386);
nor U15818 (N_15818,N_14346,N_14645);
and U15819 (N_15819,N_14514,N_14907);
nand U15820 (N_15820,N_14516,N_14643);
xnor U15821 (N_15821,N_14444,N_14646);
nor U15822 (N_15822,N_14857,N_14867);
and U15823 (N_15823,N_14457,N_14923);
or U15824 (N_15824,N_14055,N_14968);
xnor U15825 (N_15825,N_14936,N_14778);
xnor U15826 (N_15826,N_14489,N_14857);
or U15827 (N_15827,N_14553,N_14727);
or U15828 (N_15828,N_14832,N_14055);
nand U15829 (N_15829,N_14141,N_14405);
and U15830 (N_15830,N_14681,N_14808);
xor U15831 (N_15831,N_14599,N_14863);
and U15832 (N_15832,N_14670,N_14911);
nor U15833 (N_15833,N_14038,N_14656);
nand U15834 (N_15834,N_14267,N_14914);
or U15835 (N_15835,N_14405,N_14323);
xnor U15836 (N_15836,N_14357,N_14837);
and U15837 (N_15837,N_14203,N_14681);
nand U15838 (N_15838,N_14154,N_14241);
and U15839 (N_15839,N_14062,N_14663);
and U15840 (N_15840,N_14985,N_14524);
nor U15841 (N_15841,N_14183,N_14073);
nand U15842 (N_15842,N_14921,N_14134);
nor U15843 (N_15843,N_14971,N_14928);
nand U15844 (N_15844,N_14094,N_14313);
nor U15845 (N_15845,N_14328,N_14912);
nor U15846 (N_15846,N_14408,N_14255);
xor U15847 (N_15847,N_14346,N_14536);
nand U15848 (N_15848,N_14159,N_14994);
nor U15849 (N_15849,N_14695,N_14289);
xor U15850 (N_15850,N_14624,N_14788);
nand U15851 (N_15851,N_14721,N_14915);
or U15852 (N_15852,N_14051,N_14230);
and U15853 (N_15853,N_14983,N_14168);
or U15854 (N_15854,N_14477,N_14240);
or U15855 (N_15855,N_14896,N_14407);
xnor U15856 (N_15856,N_14288,N_14411);
xnor U15857 (N_15857,N_14769,N_14002);
or U15858 (N_15858,N_14354,N_14882);
and U15859 (N_15859,N_14661,N_14827);
xor U15860 (N_15860,N_14196,N_14079);
nor U15861 (N_15861,N_14232,N_14847);
xnor U15862 (N_15862,N_14536,N_14099);
or U15863 (N_15863,N_14283,N_14450);
nor U15864 (N_15864,N_14725,N_14204);
xnor U15865 (N_15865,N_14000,N_14567);
and U15866 (N_15866,N_14513,N_14832);
nand U15867 (N_15867,N_14835,N_14170);
nand U15868 (N_15868,N_14236,N_14197);
nor U15869 (N_15869,N_14480,N_14374);
nand U15870 (N_15870,N_14902,N_14660);
nor U15871 (N_15871,N_14810,N_14740);
nand U15872 (N_15872,N_14354,N_14780);
and U15873 (N_15873,N_14860,N_14294);
or U15874 (N_15874,N_14941,N_14480);
or U15875 (N_15875,N_14985,N_14768);
nor U15876 (N_15876,N_14502,N_14422);
or U15877 (N_15877,N_14072,N_14224);
or U15878 (N_15878,N_14285,N_14988);
nand U15879 (N_15879,N_14544,N_14060);
and U15880 (N_15880,N_14067,N_14492);
nor U15881 (N_15881,N_14914,N_14618);
nand U15882 (N_15882,N_14690,N_14691);
and U15883 (N_15883,N_14248,N_14467);
nand U15884 (N_15884,N_14421,N_14171);
and U15885 (N_15885,N_14341,N_14038);
or U15886 (N_15886,N_14282,N_14461);
xnor U15887 (N_15887,N_14671,N_14178);
and U15888 (N_15888,N_14620,N_14711);
or U15889 (N_15889,N_14192,N_14788);
nor U15890 (N_15890,N_14060,N_14611);
and U15891 (N_15891,N_14739,N_14749);
or U15892 (N_15892,N_14564,N_14596);
xnor U15893 (N_15893,N_14727,N_14632);
and U15894 (N_15894,N_14844,N_14202);
nor U15895 (N_15895,N_14070,N_14883);
nor U15896 (N_15896,N_14043,N_14629);
nor U15897 (N_15897,N_14729,N_14129);
nor U15898 (N_15898,N_14694,N_14782);
nor U15899 (N_15899,N_14865,N_14793);
or U15900 (N_15900,N_14961,N_14556);
xor U15901 (N_15901,N_14815,N_14850);
nor U15902 (N_15902,N_14628,N_14609);
nand U15903 (N_15903,N_14624,N_14679);
nand U15904 (N_15904,N_14171,N_14566);
xor U15905 (N_15905,N_14776,N_14068);
or U15906 (N_15906,N_14094,N_14433);
and U15907 (N_15907,N_14417,N_14318);
or U15908 (N_15908,N_14907,N_14097);
xnor U15909 (N_15909,N_14384,N_14475);
xnor U15910 (N_15910,N_14140,N_14034);
and U15911 (N_15911,N_14540,N_14264);
xor U15912 (N_15912,N_14584,N_14209);
nor U15913 (N_15913,N_14669,N_14062);
nor U15914 (N_15914,N_14684,N_14499);
nor U15915 (N_15915,N_14053,N_14817);
or U15916 (N_15916,N_14894,N_14249);
or U15917 (N_15917,N_14452,N_14495);
xnor U15918 (N_15918,N_14052,N_14884);
and U15919 (N_15919,N_14894,N_14056);
or U15920 (N_15920,N_14425,N_14212);
nand U15921 (N_15921,N_14655,N_14293);
nand U15922 (N_15922,N_14240,N_14898);
nor U15923 (N_15923,N_14100,N_14292);
and U15924 (N_15924,N_14748,N_14895);
or U15925 (N_15925,N_14570,N_14475);
nand U15926 (N_15926,N_14466,N_14695);
or U15927 (N_15927,N_14254,N_14981);
xor U15928 (N_15928,N_14047,N_14528);
and U15929 (N_15929,N_14520,N_14899);
nor U15930 (N_15930,N_14836,N_14246);
or U15931 (N_15931,N_14493,N_14032);
nand U15932 (N_15932,N_14774,N_14304);
nor U15933 (N_15933,N_14225,N_14763);
xor U15934 (N_15934,N_14397,N_14055);
nor U15935 (N_15935,N_14836,N_14994);
or U15936 (N_15936,N_14258,N_14913);
and U15937 (N_15937,N_14489,N_14801);
nand U15938 (N_15938,N_14802,N_14516);
nor U15939 (N_15939,N_14524,N_14777);
nor U15940 (N_15940,N_14423,N_14996);
and U15941 (N_15941,N_14338,N_14706);
and U15942 (N_15942,N_14793,N_14296);
xor U15943 (N_15943,N_14210,N_14409);
nor U15944 (N_15944,N_14357,N_14716);
nor U15945 (N_15945,N_14959,N_14343);
and U15946 (N_15946,N_14344,N_14317);
or U15947 (N_15947,N_14611,N_14719);
nand U15948 (N_15948,N_14420,N_14278);
xor U15949 (N_15949,N_14331,N_14277);
nand U15950 (N_15950,N_14660,N_14256);
nand U15951 (N_15951,N_14882,N_14276);
xnor U15952 (N_15952,N_14953,N_14003);
xor U15953 (N_15953,N_14819,N_14071);
nand U15954 (N_15954,N_14348,N_14506);
xnor U15955 (N_15955,N_14019,N_14037);
nand U15956 (N_15956,N_14136,N_14626);
and U15957 (N_15957,N_14481,N_14110);
or U15958 (N_15958,N_14316,N_14119);
and U15959 (N_15959,N_14448,N_14714);
xnor U15960 (N_15960,N_14863,N_14532);
or U15961 (N_15961,N_14863,N_14048);
and U15962 (N_15962,N_14895,N_14490);
nor U15963 (N_15963,N_14016,N_14185);
xnor U15964 (N_15964,N_14146,N_14162);
nor U15965 (N_15965,N_14401,N_14345);
or U15966 (N_15966,N_14030,N_14965);
xor U15967 (N_15967,N_14634,N_14329);
or U15968 (N_15968,N_14536,N_14080);
and U15969 (N_15969,N_14199,N_14831);
or U15970 (N_15970,N_14782,N_14664);
and U15971 (N_15971,N_14809,N_14724);
xor U15972 (N_15972,N_14904,N_14219);
nor U15973 (N_15973,N_14857,N_14724);
xor U15974 (N_15974,N_14259,N_14812);
nor U15975 (N_15975,N_14749,N_14960);
nor U15976 (N_15976,N_14253,N_14688);
and U15977 (N_15977,N_14350,N_14128);
or U15978 (N_15978,N_14988,N_14165);
and U15979 (N_15979,N_14984,N_14283);
nand U15980 (N_15980,N_14555,N_14650);
nand U15981 (N_15981,N_14584,N_14710);
nor U15982 (N_15982,N_14988,N_14610);
xor U15983 (N_15983,N_14982,N_14826);
or U15984 (N_15984,N_14910,N_14350);
and U15985 (N_15985,N_14552,N_14106);
nor U15986 (N_15986,N_14415,N_14824);
or U15987 (N_15987,N_14488,N_14220);
nor U15988 (N_15988,N_14505,N_14865);
and U15989 (N_15989,N_14063,N_14074);
nand U15990 (N_15990,N_14209,N_14300);
nor U15991 (N_15991,N_14607,N_14701);
nand U15992 (N_15992,N_14371,N_14054);
nor U15993 (N_15993,N_14768,N_14512);
and U15994 (N_15994,N_14640,N_14928);
and U15995 (N_15995,N_14316,N_14394);
xor U15996 (N_15996,N_14164,N_14118);
xor U15997 (N_15997,N_14109,N_14177);
or U15998 (N_15998,N_14004,N_14197);
and U15999 (N_15999,N_14391,N_14665);
nor U16000 (N_16000,N_15048,N_15663);
xnor U16001 (N_16001,N_15806,N_15608);
nor U16002 (N_16002,N_15648,N_15639);
or U16003 (N_16003,N_15547,N_15548);
and U16004 (N_16004,N_15029,N_15749);
or U16005 (N_16005,N_15607,N_15817);
and U16006 (N_16006,N_15978,N_15732);
nor U16007 (N_16007,N_15559,N_15613);
nor U16008 (N_16008,N_15763,N_15595);
or U16009 (N_16009,N_15569,N_15687);
xor U16010 (N_16010,N_15249,N_15254);
nor U16011 (N_16011,N_15622,N_15138);
nand U16012 (N_16012,N_15717,N_15565);
xnor U16013 (N_16013,N_15344,N_15491);
nor U16014 (N_16014,N_15268,N_15426);
nand U16015 (N_16015,N_15073,N_15477);
nor U16016 (N_16016,N_15093,N_15352);
and U16017 (N_16017,N_15362,N_15366);
nand U16018 (N_16018,N_15996,N_15417);
xnor U16019 (N_16019,N_15606,N_15970);
and U16020 (N_16020,N_15302,N_15780);
xnor U16021 (N_16021,N_15348,N_15209);
nor U16022 (N_16022,N_15112,N_15079);
and U16023 (N_16023,N_15785,N_15200);
nor U16024 (N_16024,N_15310,N_15410);
xor U16025 (N_16025,N_15217,N_15272);
nor U16026 (N_16026,N_15767,N_15891);
or U16027 (N_16027,N_15974,N_15598);
xnor U16028 (N_16028,N_15419,N_15935);
nand U16029 (N_16029,N_15792,N_15975);
nand U16030 (N_16030,N_15218,N_15945);
or U16031 (N_16031,N_15405,N_15323);
nor U16032 (N_16032,N_15962,N_15810);
or U16033 (N_16033,N_15492,N_15528);
xnor U16034 (N_16034,N_15279,N_15508);
nand U16035 (N_16035,N_15504,N_15852);
nand U16036 (N_16036,N_15241,N_15679);
or U16037 (N_16037,N_15418,N_15034);
nor U16038 (N_16038,N_15447,N_15963);
or U16039 (N_16039,N_15692,N_15585);
xnor U16040 (N_16040,N_15427,N_15737);
and U16041 (N_16041,N_15246,N_15248);
xnor U16042 (N_16042,N_15311,N_15726);
nand U16043 (N_16043,N_15016,N_15158);
and U16044 (N_16044,N_15425,N_15846);
nor U16045 (N_16045,N_15818,N_15681);
xor U16046 (N_16046,N_15252,N_15142);
and U16047 (N_16047,N_15951,N_15683);
nand U16048 (N_16048,N_15519,N_15887);
or U16049 (N_16049,N_15855,N_15873);
and U16050 (N_16050,N_15910,N_15654);
nor U16051 (N_16051,N_15037,N_15345);
or U16052 (N_16052,N_15295,N_15965);
nor U16053 (N_16053,N_15959,N_15340);
and U16054 (N_16054,N_15153,N_15729);
nand U16055 (N_16055,N_15214,N_15777);
nand U16056 (N_16056,N_15495,N_15986);
or U16057 (N_16057,N_15857,N_15320);
or U16058 (N_16058,N_15605,N_15004);
xnor U16059 (N_16059,N_15771,N_15721);
xnor U16060 (N_16060,N_15733,N_15841);
nor U16061 (N_16061,N_15532,N_15007);
xor U16062 (N_16062,N_15778,N_15713);
nor U16063 (N_16063,N_15646,N_15064);
nand U16064 (N_16064,N_15828,N_15616);
and U16065 (N_16065,N_15830,N_15800);
nand U16066 (N_16066,N_15689,N_15160);
and U16067 (N_16067,N_15682,N_15239);
nand U16068 (N_16068,N_15403,N_15333);
and U16069 (N_16069,N_15637,N_15432);
or U16070 (N_16070,N_15497,N_15210);
and U16071 (N_16071,N_15437,N_15757);
nor U16072 (N_16072,N_15961,N_15515);
and U16073 (N_16073,N_15745,N_15013);
and U16074 (N_16074,N_15998,N_15601);
or U16075 (N_16075,N_15191,N_15521);
or U16076 (N_16076,N_15304,N_15206);
xnor U16077 (N_16077,N_15152,N_15168);
xnor U16078 (N_16078,N_15240,N_15411);
nand U16079 (N_16079,N_15286,N_15627);
and U16080 (N_16080,N_15014,N_15898);
nand U16081 (N_16081,N_15434,N_15995);
nand U16082 (N_16082,N_15851,N_15151);
and U16083 (N_16083,N_15523,N_15685);
or U16084 (N_16084,N_15849,N_15065);
or U16085 (N_16085,N_15185,N_15212);
or U16086 (N_16086,N_15154,N_15061);
xor U16087 (N_16087,N_15755,N_15883);
nor U16088 (N_16088,N_15581,N_15102);
and U16089 (N_16089,N_15084,N_15072);
or U16090 (N_16090,N_15502,N_15439);
nor U16091 (N_16091,N_15619,N_15827);
nand U16092 (N_16092,N_15026,N_15522);
xor U16093 (N_16093,N_15047,N_15002);
nor U16094 (N_16094,N_15489,N_15364);
xnor U16095 (N_16095,N_15141,N_15285);
nand U16096 (N_16096,N_15269,N_15629);
xnor U16097 (N_16097,N_15558,N_15402);
nor U16098 (N_16098,N_15586,N_15696);
nor U16099 (N_16099,N_15684,N_15588);
and U16100 (N_16100,N_15609,N_15162);
and U16101 (N_16101,N_15174,N_15602);
nand U16102 (N_16102,N_15924,N_15095);
nand U16103 (N_16103,N_15464,N_15886);
nor U16104 (N_16104,N_15190,N_15894);
xnor U16105 (N_16105,N_15021,N_15087);
xnor U16106 (N_16106,N_15300,N_15155);
nand U16107 (N_16107,N_15568,N_15574);
and U16108 (N_16108,N_15336,N_15308);
and U16109 (N_16109,N_15135,N_15474);
nor U16110 (N_16110,N_15298,N_15765);
nand U16111 (N_16111,N_15401,N_15049);
or U16112 (N_16112,N_15005,N_15186);
xor U16113 (N_16113,N_15435,N_15192);
and U16114 (N_16114,N_15531,N_15723);
nand U16115 (N_16115,N_15150,N_15165);
nor U16116 (N_16116,N_15768,N_15372);
or U16117 (N_16117,N_15416,N_15808);
xnor U16118 (N_16118,N_15059,N_15621);
or U16119 (N_16119,N_15670,N_15467);
xnor U16120 (N_16120,N_15864,N_15707);
nand U16121 (N_16121,N_15554,N_15664);
xnor U16122 (N_16122,N_15255,N_15754);
xor U16123 (N_16123,N_15913,N_15315);
or U16124 (N_16124,N_15660,N_15843);
and U16125 (N_16125,N_15111,N_15144);
xor U16126 (N_16126,N_15469,N_15566);
nor U16127 (N_16127,N_15273,N_15727);
and U16128 (N_16128,N_15899,N_15460);
nand U16129 (N_16129,N_15100,N_15736);
nand U16130 (N_16130,N_15098,N_15573);
xor U16131 (N_16131,N_15947,N_15674);
or U16132 (N_16132,N_15067,N_15258);
nor U16133 (N_16133,N_15916,N_15261);
or U16134 (N_16134,N_15119,N_15114);
nand U16135 (N_16135,N_15475,N_15433);
nor U16136 (N_16136,N_15977,N_15610);
and U16137 (N_16137,N_15139,N_15706);
or U16138 (N_16138,N_15159,N_15739);
xor U16139 (N_16139,N_15611,N_15445);
xnor U16140 (N_16140,N_15690,N_15710);
nand U16141 (N_16141,N_15571,N_15484);
and U16142 (N_16142,N_15695,N_15866);
xor U16143 (N_16143,N_15931,N_15539);
and U16144 (N_16144,N_15888,N_15889);
or U16145 (N_16145,N_15716,N_15176);
xor U16146 (N_16146,N_15688,N_15090);
xnor U16147 (N_16147,N_15507,N_15636);
nor U16148 (N_16148,N_15877,N_15099);
nor U16149 (N_16149,N_15053,N_15546);
nor U16150 (N_16150,N_15809,N_15089);
nand U16151 (N_16151,N_15166,N_15035);
nand U16152 (N_16152,N_15537,N_15494);
nor U16153 (N_16153,N_15589,N_15872);
nor U16154 (N_16154,N_15193,N_15381);
nand U16155 (N_16155,N_15337,N_15587);
nor U16156 (N_16156,N_15413,N_15634);
nand U16157 (N_16157,N_15431,N_15786);
nor U16158 (N_16158,N_15705,N_15329);
or U16159 (N_16159,N_15902,N_15980);
nand U16160 (N_16160,N_15594,N_15057);
nand U16161 (N_16161,N_15673,N_15700);
or U16162 (N_16162,N_15972,N_15470);
nor U16163 (N_16163,N_15094,N_15330);
nor U16164 (N_16164,N_15908,N_15997);
and U16165 (N_16165,N_15450,N_15224);
xor U16166 (N_16166,N_15526,N_15031);
xor U16167 (N_16167,N_15911,N_15371);
xor U16168 (N_16168,N_15010,N_15479);
nor U16169 (N_16169,N_15487,N_15488);
and U16170 (N_16170,N_15271,N_15291);
xor U16171 (N_16171,N_15844,N_15867);
xor U16172 (N_16172,N_15243,N_15283);
nor U16173 (N_16173,N_15208,N_15836);
xor U16174 (N_16174,N_15422,N_15562);
nor U16175 (N_16175,N_15091,N_15143);
xnor U16176 (N_16176,N_15884,N_15868);
nand U16177 (N_16177,N_15436,N_15615);
and U16178 (N_16178,N_15661,N_15046);
nand U16179 (N_16179,N_15979,N_15576);
nand U16180 (N_16180,N_15990,N_15245);
nand U16181 (N_16181,N_15604,N_15787);
and U16182 (N_16182,N_15288,N_15630);
xnor U16183 (N_16183,N_15060,N_15443);
and U16184 (N_16184,N_15327,N_15544);
nor U16185 (N_16185,N_15582,N_15761);
or U16186 (N_16186,N_15662,N_15989);
nor U16187 (N_16187,N_15070,N_15938);
xnor U16188 (N_16188,N_15472,N_15505);
nor U16189 (N_16189,N_15205,N_15038);
xnor U16190 (N_16190,N_15635,N_15770);
or U16191 (N_16191,N_15612,N_15735);
nor U16192 (N_16192,N_15213,N_15316);
and U16193 (N_16193,N_15032,N_15314);
or U16194 (N_16194,N_15944,N_15398);
nand U16195 (N_16195,N_15306,N_15369);
or U16196 (N_16196,N_15878,N_15642);
nand U16197 (N_16197,N_15317,N_15077);
nor U16198 (N_16198,N_15517,N_15510);
and U16199 (N_16199,N_15753,N_15033);
and U16200 (N_16200,N_15686,N_15772);
xnor U16201 (N_16201,N_15137,N_15386);
nor U16202 (N_16202,N_15197,N_15179);
nand U16203 (N_16203,N_15365,N_15578);
nand U16204 (N_16204,N_15628,N_15313);
nand U16205 (N_16205,N_15698,N_15506);
and U16206 (N_16206,N_15232,N_15359);
nand U16207 (N_16207,N_15549,N_15912);
nor U16208 (N_16208,N_15744,N_15020);
nor U16209 (N_16209,N_15062,N_15019);
nor U16210 (N_16210,N_15861,N_15430);
nand U16211 (N_16211,N_15027,N_15643);
nand U16212 (N_16212,N_15829,N_15129);
xnor U16213 (N_16213,N_15001,N_15096);
nor U16214 (N_16214,N_15927,N_15764);
nor U16215 (N_16215,N_15535,N_15242);
xor U16216 (N_16216,N_15520,N_15292);
or U16217 (N_16217,N_15324,N_15882);
nor U16218 (N_16218,N_15069,N_15983);
or U16219 (N_16219,N_15968,N_15379);
nor U16220 (N_16220,N_15950,N_15260);
or U16221 (N_16221,N_15584,N_15534);
and U16222 (N_16222,N_15921,N_15455);
nand U16223 (N_16223,N_15363,N_15335);
xor U16224 (N_16224,N_15025,N_15656);
and U16225 (N_16225,N_15711,N_15804);
xor U16226 (N_16226,N_15383,N_15428);
nor U16227 (N_16227,N_15188,N_15955);
and U16228 (N_16228,N_15473,N_15513);
nor U16229 (N_16229,N_15332,N_15967);
xnor U16230 (N_16230,N_15115,N_15468);
nand U16231 (N_16231,N_15361,N_15597);
nor U16232 (N_16232,N_15650,N_15390);
and U16233 (N_16233,N_15774,N_15697);
nor U16234 (N_16234,N_15550,N_15189);
or U16235 (N_16235,N_15287,N_15238);
xnor U16236 (N_16236,N_15555,N_15799);
nand U16237 (N_16237,N_15540,N_15408);
nand U16238 (N_16238,N_15230,N_15264);
or U16239 (N_16239,N_15915,N_15126);
or U16240 (N_16240,N_15703,N_15058);
nand U16241 (N_16241,N_15227,N_15655);
nand U16242 (N_16242,N_15907,N_15498);
nor U16243 (N_16243,N_15766,N_15220);
xnor U16244 (N_16244,N_15922,N_15929);
nand U16245 (N_16245,N_15044,N_15590);
or U16246 (N_16246,N_15175,N_15824);
nand U16247 (N_16247,N_15395,N_15163);
nand U16248 (N_16248,N_15815,N_15463);
xnor U16249 (N_16249,N_15665,N_15346);
nor U16250 (N_16250,N_15625,N_15109);
nor U16251 (N_16251,N_15719,N_15368);
nor U16252 (N_16252,N_15458,N_15853);
nor U16253 (N_16253,N_15832,N_15219);
or U16254 (N_16254,N_15904,N_15042);
nand U16255 (N_16255,N_15600,N_15289);
or U16256 (N_16256,N_15842,N_15128);
nand U16257 (N_16257,N_15712,N_15040);
nor U16258 (N_16258,N_15518,N_15149);
xor U16259 (N_16259,N_15134,N_15483);
xor U16260 (N_16260,N_15876,N_15577);
nor U16261 (N_16261,N_15274,N_15860);
and U16262 (N_16262,N_15409,N_15028);
nand U16263 (N_16263,N_15756,N_15747);
and U16264 (N_16264,N_15869,N_15400);
or U16265 (N_16265,N_15708,N_15840);
or U16266 (N_16266,N_15805,N_15167);
xor U16267 (N_16267,N_15415,N_15850);
xnor U16268 (N_16268,N_15294,N_15941);
nor U16269 (N_16269,N_15451,N_15375);
nand U16270 (N_16270,N_15082,N_15543);
nor U16271 (N_16271,N_15669,N_15797);
nand U16272 (N_16272,N_15045,N_15183);
nor U16273 (N_16273,N_15976,N_15798);
or U16274 (N_16274,N_15136,N_15837);
xnor U16275 (N_16275,N_15303,N_15516);
nor U16276 (N_16276,N_15956,N_15318);
and U16277 (N_16277,N_15811,N_15078);
nand U16278 (N_16278,N_15389,N_15652);
nand U16279 (N_16279,N_15934,N_15351);
or U16280 (N_16280,N_15056,N_15457);
nand U16281 (N_16281,N_15591,N_15856);
nand U16282 (N_16282,N_15448,N_15377);
nand U16283 (N_16283,N_15958,N_15380);
nor U16284 (N_16284,N_15299,N_15592);
xnor U16285 (N_16285,N_15404,N_15216);
and U16286 (N_16286,N_15942,N_15130);
and U16287 (N_16287,N_15552,N_15499);
nor U16288 (N_16288,N_15795,N_15501);
nand U16289 (N_16289,N_15617,N_15834);
xor U16290 (N_16290,N_15985,N_15266);
nor U16291 (N_16291,N_15940,N_15406);
nor U16292 (N_16292,N_15131,N_15339);
nor U16293 (N_16293,N_15527,N_15235);
nand U16294 (N_16294,N_15341,N_15905);
nand U16295 (N_16295,N_15123,N_15715);
and U16296 (N_16296,N_15080,N_15229);
nand U16297 (N_16297,N_15847,N_15357);
xor U16298 (N_16298,N_15181,N_15781);
nand U16299 (N_16299,N_15171,N_15999);
xor U16300 (N_16300,N_15953,N_15113);
nor U16301 (N_16301,N_15140,N_15796);
nor U16302 (N_16302,N_15890,N_15125);
xor U16303 (N_16303,N_15909,N_15831);
nor U16304 (N_16304,N_15173,N_15728);
and U16305 (N_16305,N_15259,N_15897);
nand U16306 (N_16306,N_15741,N_15250);
xor U16307 (N_16307,N_15257,N_15374);
nor U16308 (N_16308,N_15807,N_15453);
nand U16309 (N_16309,N_15691,N_15305);
nand U16310 (N_16310,N_15036,N_15881);
nand U16311 (N_16311,N_15462,N_15478);
nand U16312 (N_16312,N_15752,N_15184);
nand U16313 (N_16313,N_15788,N_15482);
and U16314 (N_16314,N_15465,N_15172);
xnor U16315 (N_16315,N_15511,N_15039);
or U16316 (N_16316,N_15790,N_15023);
or U16317 (N_16317,N_15182,N_15969);
nand U16318 (N_16318,N_15440,N_15814);
or U16319 (N_16319,N_15066,N_15006);
and U16320 (N_16320,N_15759,N_15120);
xnor U16321 (N_16321,N_15812,N_15743);
nand U16322 (N_16322,N_15496,N_15903);
xor U16323 (N_16323,N_15614,N_15525);
nor U16324 (N_16324,N_15760,N_15164);
xnor U16325 (N_16325,N_15122,N_15370);
xnor U16326 (N_16326,N_15821,N_15018);
nand U16327 (N_16327,N_15981,N_15051);
and U16328 (N_16328,N_15012,N_15097);
xnor U16329 (N_16329,N_15791,N_15349);
nand U16330 (N_16330,N_15966,N_15423);
nand U16331 (N_16331,N_15068,N_15284);
and U16332 (N_16332,N_15694,N_15226);
nor U16333 (N_16333,N_15680,N_15993);
and U16334 (N_16334,N_15008,N_15776);
xnor U16335 (N_16335,N_15623,N_15071);
nor U16336 (N_16336,N_15748,N_15009);
and U16337 (N_16337,N_15557,N_15750);
and U16338 (N_16338,N_15542,N_15177);
nand U16339 (N_16339,N_15461,N_15917);
xor U16340 (N_16340,N_15347,N_15301);
and U16341 (N_16341,N_15533,N_15223);
xnor U16342 (N_16342,N_15514,N_15678);
nor U16343 (N_16343,N_15987,N_15251);
nor U16344 (N_16344,N_15848,N_15107);
nand U16345 (N_16345,N_15822,N_15399);
nand U16346 (N_16346,N_15724,N_15074);
nand U16347 (N_16347,N_15180,N_15024);
xor U16348 (N_16348,N_15353,N_15556);
nor U16349 (N_16349,N_15309,N_15823);
nand U16350 (N_16350,N_15011,N_15378);
and U16351 (N_16351,N_15281,N_15454);
xor U16352 (N_16352,N_15722,N_15263);
xnor U16353 (N_16353,N_15593,N_15779);
xor U16354 (N_16354,N_15041,N_15936);
nor U16355 (N_16355,N_15971,N_15198);
xnor U16356 (N_16356,N_15338,N_15839);
and U16357 (N_16357,N_15992,N_15561);
xor U16358 (N_16358,N_15580,N_15476);
xor U16359 (N_16359,N_15793,N_15367);
or U16360 (N_16360,N_15933,N_15503);
or U16361 (N_16361,N_15196,N_15355);
nand U16362 (N_16362,N_15480,N_15833);
xnor U16363 (N_16363,N_15896,N_15657);
nand U16364 (N_16364,N_15782,N_15583);
and U16365 (N_16365,N_15276,N_15645);
xnor U16366 (N_16366,N_15485,N_15106);
nand U16367 (N_16367,N_15512,N_15148);
or U16368 (N_16368,N_15858,N_15730);
xnor U16369 (N_16369,N_15826,N_15414);
nand U16370 (N_16370,N_15994,N_15030);
xor U16371 (N_16371,N_15412,N_15396);
xor U16372 (N_16372,N_15862,N_15343);
xnor U16373 (N_16373,N_15640,N_15803);
and U16374 (N_16374,N_15043,N_15704);
or U16375 (N_16375,N_15820,N_15603);
and U16376 (N_16376,N_15222,N_15170);
xnor U16377 (N_16377,N_15215,N_15874);
xnor U16378 (N_16378,N_15000,N_15638);
nand U16379 (N_16379,N_15957,N_15802);
or U16380 (N_16380,N_15221,N_15575);
nand U16381 (N_16381,N_15354,N_15312);
and U16382 (N_16382,N_15734,N_15784);
or U16383 (N_16383,N_15199,N_15247);
nor U16384 (N_16384,N_15675,N_15751);
xor U16385 (N_16385,N_15509,N_15262);
nand U16386 (N_16386,N_15919,N_15863);
or U16387 (N_16387,N_15233,N_15725);
nand U16388 (N_16388,N_15103,N_15659);
or U16389 (N_16389,N_15178,N_15564);
nand U16390 (N_16390,N_15195,N_15923);
and U16391 (N_16391,N_15988,N_15816);
nor U16392 (N_16392,N_15421,N_15157);
and U16393 (N_16393,N_15668,N_15373);
nand U16394 (N_16394,N_15438,N_15277);
or U16395 (N_16395,N_15105,N_15169);
xnor U16396 (N_16396,N_15116,N_15702);
or U16397 (N_16397,N_15641,N_15633);
or U16398 (N_16398,N_15649,N_15948);
and U16399 (N_16399,N_15892,N_15296);
or U16400 (N_16400,N_15536,N_15083);
nor U16401 (N_16401,N_15901,N_15081);
or U16402 (N_16402,N_15859,N_15388);
or U16403 (N_16403,N_15146,N_15937);
xnor U16404 (N_16404,N_15570,N_15984);
nor U16405 (N_16405,N_15393,N_15783);
nor U16406 (N_16406,N_15290,N_15356);
or U16407 (N_16407,N_15456,N_15775);
and U16408 (N_16408,N_15110,N_15572);
nor U16409 (N_16409,N_15328,N_15845);
nor U16410 (N_16410,N_15055,N_15088);
xnor U16411 (N_16411,N_15202,N_15444);
nand U16412 (N_16412,N_15651,N_15325);
or U16413 (N_16413,N_15054,N_15631);
nand U16414 (N_16414,N_15677,N_15086);
or U16415 (N_16415,N_15397,N_15231);
xnor U16416 (N_16416,N_15553,N_15236);
nand U16417 (N_16417,N_15579,N_15762);
nand U16418 (N_16418,N_15376,N_15280);
or U16419 (N_16419,N_15321,N_15709);
xor U16420 (N_16420,N_15865,N_15121);
nor U16421 (N_16421,N_15420,N_15952);
nand U16422 (N_16422,N_15746,N_15538);
nand U16423 (N_16423,N_15854,N_15441);
nand U16424 (N_16424,N_15334,N_15392);
or U16425 (N_16425,N_15391,N_15204);
xor U16426 (N_16426,N_15265,N_15900);
or U16427 (N_16427,N_15738,N_15201);
xor U16428 (N_16428,N_15145,N_15560);
nand U16429 (N_16429,N_15124,N_15835);
and U16430 (N_16430,N_15253,N_15319);
and U16431 (N_16431,N_15358,N_15740);
or U16432 (N_16432,N_15893,N_15331);
or U16433 (N_16433,N_15267,N_15914);
or U16434 (N_16434,N_15880,N_15599);
nor U16435 (N_16435,N_15644,N_15949);
nor U16436 (N_16436,N_15085,N_15161);
nand U16437 (N_16437,N_15524,N_15672);
or U16438 (N_16438,N_15714,N_15187);
nand U16439 (N_16439,N_15667,N_15234);
and U16440 (N_16440,N_15943,N_15394);
and U16441 (N_16441,N_15108,N_15132);
nand U16442 (N_16442,N_15076,N_15307);
nand U16443 (N_16443,N_15449,N_15466);
nor U16444 (N_16444,N_15228,N_15282);
and U16445 (N_16445,N_15720,N_15838);
xor U16446 (N_16446,N_15493,N_15819);
and U16447 (N_16447,N_15015,N_15481);
nand U16448 (N_16448,N_15442,N_15211);
and U16449 (N_16449,N_15275,N_15147);
nand U16450 (N_16450,N_15954,N_15742);
and U16451 (N_16451,N_15063,N_15794);
and U16452 (N_16452,N_15384,N_15666);
or U16453 (N_16453,N_15133,N_15022);
and U16454 (N_16454,N_15701,N_15278);
xnor U16455 (N_16455,N_15789,N_15541);
or U16456 (N_16456,N_15671,N_15926);
and U16457 (N_16457,N_15939,N_15885);
nor U16458 (N_16458,N_15075,N_15237);
or U16459 (N_16459,N_15156,N_15429);
xor U16460 (N_16460,N_15471,N_15567);
and U16461 (N_16461,N_15870,N_15117);
nor U16462 (N_16462,N_15653,N_15459);
and U16463 (N_16463,N_15626,N_15387);
nor U16464 (N_16464,N_15407,N_15446);
and U16465 (N_16465,N_15932,N_15946);
or U16466 (N_16466,N_15385,N_15293);
nor U16467 (N_16467,N_15925,N_15530);
xnor U16468 (N_16468,N_15693,N_15326);
nand U16469 (N_16469,N_15101,N_15297);
xnor U16470 (N_16470,N_15825,N_15194);
or U16471 (N_16471,N_15930,N_15982);
xor U16472 (N_16472,N_15871,N_15928);
or U16473 (N_16473,N_15382,N_15813);
nor U16474 (N_16474,N_15017,N_15960);
nor U16475 (N_16475,N_15973,N_15624);
xor U16476 (N_16476,N_15225,N_15991);
nor U16477 (N_16477,N_15875,N_15906);
and U16478 (N_16478,N_15127,N_15207);
nand U16479 (N_16479,N_15879,N_15244);
xnor U16480 (N_16480,N_15529,N_15658);
and U16481 (N_16481,N_15203,N_15104);
and U16482 (N_16482,N_15270,N_15632);
and U16483 (N_16483,N_15256,N_15773);
or U16484 (N_16484,N_15003,N_15731);
xor U16485 (N_16485,N_15118,N_15758);
xnor U16486 (N_16486,N_15052,N_15500);
nor U16487 (N_16487,N_15647,N_15050);
nor U16488 (N_16488,N_15486,N_15342);
and U16489 (N_16489,N_15769,N_15596);
xor U16490 (N_16490,N_15322,N_15563);
and U16491 (N_16491,N_15699,N_15092);
or U16492 (N_16492,N_15895,N_15360);
xor U16493 (N_16493,N_15545,N_15801);
nor U16494 (N_16494,N_15452,N_15350);
or U16495 (N_16495,N_15918,N_15718);
and U16496 (N_16496,N_15620,N_15920);
or U16497 (N_16497,N_15676,N_15618);
nand U16498 (N_16498,N_15551,N_15964);
nand U16499 (N_16499,N_15424,N_15490);
nor U16500 (N_16500,N_15670,N_15292);
nand U16501 (N_16501,N_15969,N_15082);
xor U16502 (N_16502,N_15399,N_15191);
nor U16503 (N_16503,N_15958,N_15536);
nor U16504 (N_16504,N_15459,N_15463);
nand U16505 (N_16505,N_15387,N_15207);
and U16506 (N_16506,N_15231,N_15128);
and U16507 (N_16507,N_15688,N_15739);
nor U16508 (N_16508,N_15063,N_15500);
and U16509 (N_16509,N_15984,N_15373);
xnor U16510 (N_16510,N_15746,N_15837);
xnor U16511 (N_16511,N_15773,N_15778);
xor U16512 (N_16512,N_15250,N_15764);
nand U16513 (N_16513,N_15473,N_15297);
and U16514 (N_16514,N_15772,N_15768);
nor U16515 (N_16515,N_15443,N_15681);
nor U16516 (N_16516,N_15208,N_15546);
nor U16517 (N_16517,N_15132,N_15250);
and U16518 (N_16518,N_15428,N_15029);
xnor U16519 (N_16519,N_15672,N_15586);
and U16520 (N_16520,N_15865,N_15460);
and U16521 (N_16521,N_15540,N_15905);
nand U16522 (N_16522,N_15912,N_15141);
or U16523 (N_16523,N_15662,N_15890);
xnor U16524 (N_16524,N_15933,N_15320);
xor U16525 (N_16525,N_15584,N_15347);
nor U16526 (N_16526,N_15828,N_15609);
xnor U16527 (N_16527,N_15031,N_15992);
nor U16528 (N_16528,N_15936,N_15306);
and U16529 (N_16529,N_15177,N_15594);
nor U16530 (N_16530,N_15595,N_15133);
or U16531 (N_16531,N_15172,N_15398);
xnor U16532 (N_16532,N_15886,N_15563);
and U16533 (N_16533,N_15917,N_15396);
or U16534 (N_16534,N_15523,N_15299);
and U16535 (N_16535,N_15335,N_15459);
and U16536 (N_16536,N_15425,N_15754);
and U16537 (N_16537,N_15543,N_15207);
and U16538 (N_16538,N_15688,N_15413);
nand U16539 (N_16539,N_15186,N_15954);
xor U16540 (N_16540,N_15881,N_15972);
or U16541 (N_16541,N_15396,N_15893);
or U16542 (N_16542,N_15473,N_15824);
nor U16543 (N_16543,N_15072,N_15223);
nand U16544 (N_16544,N_15044,N_15071);
xor U16545 (N_16545,N_15890,N_15101);
or U16546 (N_16546,N_15138,N_15552);
xor U16547 (N_16547,N_15421,N_15166);
or U16548 (N_16548,N_15298,N_15166);
nor U16549 (N_16549,N_15787,N_15629);
nor U16550 (N_16550,N_15058,N_15701);
nand U16551 (N_16551,N_15468,N_15280);
or U16552 (N_16552,N_15861,N_15265);
nor U16553 (N_16553,N_15213,N_15085);
xnor U16554 (N_16554,N_15711,N_15098);
nand U16555 (N_16555,N_15890,N_15881);
nor U16556 (N_16556,N_15340,N_15105);
nand U16557 (N_16557,N_15349,N_15150);
xnor U16558 (N_16558,N_15849,N_15018);
or U16559 (N_16559,N_15444,N_15770);
nand U16560 (N_16560,N_15216,N_15277);
or U16561 (N_16561,N_15509,N_15543);
xnor U16562 (N_16562,N_15226,N_15039);
nor U16563 (N_16563,N_15792,N_15746);
nor U16564 (N_16564,N_15546,N_15891);
nand U16565 (N_16565,N_15648,N_15924);
and U16566 (N_16566,N_15871,N_15555);
nand U16567 (N_16567,N_15422,N_15594);
nand U16568 (N_16568,N_15482,N_15447);
xnor U16569 (N_16569,N_15834,N_15623);
xnor U16570 (N_16570,N_15185,N_15443);
nand U16571 (N_16571,N_15891,N_15172);
xor U16572 (N_16572,N_15048,N_15830);
and U16573 (N_16573,N_15020,N_15796);
or U16574 (N_16574,N_15116,N_15046);
and U16575 (N_16575,N_15294,N_15367);
or U16576 (N_16576,N_15398,N_15049);
or U16577 (N_16577,N_15836,N_15017);
nand U16578 (N_16578,N_15771,N_15637);
or U16579 (N_16579,N_15514,N_15624);
nor U16580 (N_16580,N_15120,N_15442);
or U16581 (N_16581,N_15747,N_15014);
nor U16582 (N_16582,N_15804,N_15933);
nor U16583 (N_16583,N_15258,N_15702);
xnor U16584 (N_16584,N_15014,N_15457);
and U16585 (N_16585,N_15686,N_15774);
nand U16586 (N_16586,N_15242,N_15578);
xnor U16587 (N_16587,N_15661,N_15277);
and U16588 (N_16588,N_15091,N_15249);
and U16589 (N_16589,N_15948,N_15121);
nand U16590 (N_16590,N_15672,N_15650);
nand U16591 (N_16591,N_15270,N_15406);
and U16592 (N_16592,N_15440,N_15001);
nand U16593 (N_16593,N_15491,N_15872);
nand U16594 (N_16594,N_15389,N_15169);
nor U16595 (N_16595,N_15893,N_15546);
nor U16596 (N_16596,N_15612,N_15704);
and U16597 (N_16597,N_15621,N_15492);
or U16598 (N_16598,N_15209,N_15819);
xor U16599 (N_16599,N_15870,N_15951);
xnor U16600 (N_16600,N_15744,N_15959);
nand U16601 (N_16601,N_15628,N_15695);
nor U16602 (N_16602,N_15716,N_15744);
nor U16603 (N_16603,N_15262,N_15638);
or U16604 (N_16604,N_15596,N_15870);
or U16605 (N_16605,N_15385,N_15816);
xor U16606 (N_16606,N_15694,N_15531);
xor U16607 (N_16607,N_15265,N_15130);
nand U16608 (N_16608,N_15242,N_15968);
nor U16609 (N_16609,N_15451,N_15163);
xor U16610 (N_16610,N_15616,N_15815);
xnor U16611 (N_16611,N_15752,N_15420);
nand U16612 (N_16612,N_15686,N_15529);
nor U16613 (N_16613,N_15305,N_15993);
xnor U16614 (N_16614,N_15855,N_15971);
or U16615 (N_16615,N_15464,N_15893);
xnor U16616 (N_16616,N_15212,N_15828);
and U16617 (N_16617,N_15040,N_15323);
nand U16618 (N_16618,N_15985,N_15458);
xnor U16619 (N_16619,N_15654,N_15608);
nand U16620 (N_16620,N_15381,N_15574);
nand U16621 (N_16621,N_15513,N_15936);
nor U16622 (N_16622,N_15266,N_15102);
and U16623 (N_16623,N_15901,N_15856);
and U16624 (N_16624,N_15719,N_15911);
nand U16625 (N_16625,N_15483,N_15664);
nor U16626 (N_16626,N_15047,N_15568);
nor U16627 (N_16627,N_15143,N_15088);
nand U16628 (N_16628,N_15557,N_15053);
and U16629 (N_16629,N_15621,N_15400);
nand U16630 (N_16630,N_15080,N_15671);
and U16631 (N_16631,N_15520,N_15101);
nor U16632 (N_16632,N_15716,N_15907);
or U16633 (N_16633,N_15307,N_15638);
nor U16634 (N_16634,N_15195,N_15001);
and U16635 (N_16635,N_15658,N_15128);
and U16636 (N_16636,N_15329,N_15954);
and U16637 (N_16637,N_15415,N_15248);
or U16638 (N_16638,N_15122,N_15810);
and U16639 (N_16639,N_15439,N_15648);
and U16640 (N_16640,N_15437,N_15512);
xor U16641 (N_16641,N_15976,N_15605);
or U16642 (N_16642,N_15338,N_15585);
xnor U16643 (N_16643,N_15876,N_15097);
xnor U16644 (N_16644,N_15898,N_15037);
nor U16645 (N_16645,N_15984,N_15324);
nand U16646 (N_16646,N_15478,N_15489);
and U16647 (N_16647,N_15952,N_15991);
nand U16648 (N_16648,N_15842,N_15168);
nand U16649 (N_16649,N_15090,N_15093);
or U16650 (N_16650,N_15730,N_15056);
or U16651 (N_16651,N_15440,N_15100);
xnor U16652 (N_16652,N_15432,N_15782);
nand U16653 (N_16653,N_15274,N_15102);
xnor U16654 (N_16654,N_15075,N_15209);
xor U16655 (N_16655,N_15537,N_15892);
nor U16656 (N_16656,N_15580,N_15018);
nor U16657 (N_16657,N_15553,N_15244);
nor U16658 (N_16658,N_15673,N_15760);
or U16659 (N_16659,N_15749,N_15887);
and U16660 (N_16660,N_15603,N_15178);
or U16661 (N_16661,N_15310,N_15039);
or U16662 (N_16662,N_15899,N_15642);
nor U16663 (N_16663,N_15279,N_15385);
and U16664 (N_16664,N_15842,N_15929);
nor U16665 (N_16665,N_15081,N_15289);
xnor U16666 (N_16666,N_15723,N_15501);
nand U16667 (N_16667,N_15531,N_15422);
nor U16668 (N_16668,N_15287,N_15519);
and U16669 (N_16669,N_15903,N_15295);
or U16670 (N_16670,N_15592,N_15745);
nor U16671 (N_16671,N_15406,N_15932);
nand U16672 (N_16672,N_15025,N_15620);
or U16673 (N_16673,N_15476,N_15061);
nand U16674 (N_16674,N_15224,N_15552);
or U16675 (N_16675,N_15465,N_15650);
xnor U16676 (N_16676,N_15493,N_15381);
xnor U16677 (N_16677,N_15324,N_15808);
nor U16678 (N_16678,N_15575,N_15725);
and U16679 (N_16679,N_15201,N_15253);
xor U16680 (N_16680,N_15708,N_15439);
nand U16681 (N_16681,N_15107,N_15270);
nor U16682 (N_16682,N_15889,N_15267);
xnor U16683 (N_16683,N_15265,N_15009);
xnor U16684 (N_16684,N_15813,N_15882);
xor U16685 (N_16685,N_15277,N_15904);
nand U16686 (N_16686,N_15896,N_15856);
nor U16687 (N_16687,N_15139,N_15464);
nand U16688 (N_16688,N_15505,N_15594);
and U16689 (N_16689,N_15279,N_15365);
or U16690 (N_16690,N_15336,N_15785);
xnor U16691 (N_16691,N_15825,N_15480);
nand U16692 (N_16692,N_15900,N_15114);
nor U16693 (N_16693,N_15496,N_15241);
nor U16694 (N_16694,N_15206,N_15309);
or U16695 (N_16695,N_15809,N_15146);
and U16696 (N_16696,N_15093,N_15468);
nor U16697 (N_16697,N_15691,N_15898);
xor U16698 (N_16698,N_15205,N_15917);
nand U16699 (N_16699,N_15621,N_15722);
nand U16700 (N_16700,N_15169,N_15321);
and U16701 (N_16701,N_15077,N_15160);
and U16702 (N_16702,N_15189,N_15185);
and U16703 (N_16703,N_15464,N_15737);
nand U16704 (N_16704,N_15060,N_15451);
or U16705 (N_16705,N_15962,N_15498);
xnor U16706 (N_16706,N_15312,N_15965);
nand U16707 (N_16707,N_15519,N_15546);
and U16708 (N_16708,N_15657,N_15820);
nand U16709 (N_16709,N_15572,N_15124);
nand U16710 (N_16710,N_15561,N_15278);
nor U16711 (N_16711,N_15437,N_15150);
nand U16712 (N_16712,N_15462,N_15327);
nand U16713 (N_16713,N_15606,N_15889);
or U16714 (N_16714,N_15585,N_15751);
nor U16715 (N_16715,N_15739,N_15231);
nor U16716 (N_16716,N_15732,N_15690);
and U16717 (N_16717,N_15870,N_15860);
or U16718 (N_16718,N_15580,N_15114);
or U16719 (N_16719,N_15285,N_15213);
nand U16720 (N_16720,N_15383,N_15823);
nand U16721 (N_16721,N_15976,N_15392);
or U16722 (N_16722,N_15069,N_15450);
nand U16723 (N_16723,N_15735,N_15729);
nand U16724 (N_16724,N_15559,N_15301);
nor U16725 (N_16725,N_15781,N_15962);
nand U16726 (N_16726,N_15103,N_15988);
xnor U16727 (N_16727,N_15728,N_15180);
nand U16728 (N_16728,N_15049,N_15662);
or U16729 (N_16729,N_15045,N_15853);
or U16730 (N_16730,N_15588,N_15696);
and U16731 (N_16731,N_15247,N_15532);
or U16732 (N_16732,N_15584,N_15626);
or U16733 (N_16733,N_15518,N_15420);
nand U16734 (N_16734,N_15866,N_15822);
nand U16735 (N_16735,N_15140,N_15450);
xor U16736 (N_16736,N_15576,N_15733);
or U16737 (N_16737,N_15109,N_15631);
or U16738 (N_16738,N_15970,N_15019);
nand U16739 (N_16739,N_15528,N_15790);
nand U16740 (N_16740,N_15997,N_15160);
nor U16741 (N_16741,N_15881,N_15693);
and U16742 (N_16742,N_15481,N_15676);
nand U16743 (N_16743,N_15922,N_15836);
xnor U16744 (N_16744,N_15666,N_15146);
nand U16745 (N_16745,N_15815,N_15409);
nor U16746 (N_16746,N_15968,N_15766);
or U16747 (N_16747,N_15154,N_15308);
nand U16748 (N_16748,N_15319,N_15065);
nor U16749 (N_16749,N_15770,N_15477);
or U16750 (N_16750,N_15399,N_15234);
nand U16751 (N_16751,N_15522,N_15751);
and U16752 (N_16752,N_15186,N_15143);
nand U16753 (N_16753,N_15791,N_15640);
and U16754 (N_16754,N_15318,N_15458);
nor U16755 (N_16755,N_15876,N_15015);
nor U16756 (N_16756,N_15462,N_15755);
nand U16757 (N_16757,N_15384,N_15104);
nor U16758 (N_16758,N_15437,N_15462);
and U16759 (N_16759,N_15245,N_15740);
nor U16760 (N_16760,N_15193,N_15661);
nand U16761 (N_16761,N_15172,N_15083);
and U16762 (N_16762,N_15817,N_15935);
xnor U16763 (N_16763,N_15990,N_15178);
nor U16764 (N_16764,N_15893,N_15403);
and U16765 (N_16765,N_15601,N_15868);
xor U16766 (N_16766,N_15520,N_15699);
xor U16767 (N_16767,N_15345,N_15678);
nand U16768 (N_16768,N_15556,N_15641);
nor U16769 (N_16769,N_15837,N_15743);
nor U16770 (N_16770,N_15216,N_15485);
nor U16771 (N_16771,N_15506,N_15284);
nor U16772 (N_16772,N_15804,N_15319);
xnor U16773 (N_16773,N_15283,N_15422);
nand U16774 (N_16774,N_15509,N_15284);
and U16775 (N_16775,N_15445,N_15082);
xnor U16776 (N_16776,N_15237,N_15818);
and U16777 (N_16777,N_15075,N_15322);
or U16778 (N_16778,N_15896,N_15428);
nor U16779 (N_16779,N_15030,N_15115);
and U16780 (N_16780,N_15094,N_15836);
nor U16781 (N_16781,N_15981,N_15437);
xor U16782 (N_16782,N_15993,N_15103);
nor U16783 (N_16783,N_15464,N_15117);
nand U16784 (N_16784,N_15840,N_15357);
or U16785 (N_16785,N_15845,N_15618);
xnor U16786 (N_16786,N_15076,N_15517);
or U16787 (N_16787,N_15207,N_15934);
and U16788 (N_16788,N_15184,N_15930);
nor U16789 (N_16789,N_15267,N_15724);
nand U16790 (N_16790,N_15843,N_15891);
nand U16791 (N_16791,N_15990,N_15256);
or U16792 (N_16792,N_15596,N_15701);
and U16793 (N_16793,N_15126,N_15918);
or U16794 (N_16794,N_15818,N_15398);
xor U16795 (N_16795,N_15190,N_15863);
nor U16796 (N_16796,N_15898,N_15987);
xnor U16797 (N_16797,N_15868,N_15448);
nand U16798 (N_16798,N_15043,N_15016);
or U16799 (N_16799,N_15896,N_15300);
and U16800 (N_16800,N_15178,N_15586);
xnor U16801 (N_16801,N_15821,N_15703);
and U16802 (N_16802,N_15939,N_15886);
and U16803 (N_16803,N_15944,N_15483);
or U16804 (N_16804,N_15127,N_15612);
nor U16805 (N_16805,N_15633,N_15380);
xnor U16806 (N_16806,N_15596,N_15084);
or U16807 (N_16807,N_15436,N_15348);
xnor U16808 (N_16808,N_15179,N_15065);
nor U16809 (N_16809,N_15507,N_15883);
and U16810 (N_16810,N_15288,N_15685);
and U16811 (N_16811,N_15311,N_15742);
and U16812 (N_16812,N_15439,N_15249);
or U16813 (N_16813,N_15211,N_15293);
or U16814 (N_16814,N_15106,N_15216);
and U16815 (N_16815,N_15504,N_15618);
xor U16816 (N_16816,N_15477,N_15354);
nor U16817 (N_16817,N_15195,N_15824);
nand U16818 (N_16818,N_15644,N_15301);
nand U16819 (N_16819,N_15311,N_15675);
nand U16820 (N_16820,N_15454,N_15129);
nand U16821 (N_16821,N_15192,N_15930);
nand U16822 (N_16822,N_15389,N_15375);
and U16823 (N_16823,N_15002,N_15597);
nor U16824 (N_16824,N_15456,N_15308);
and U16825 (N_16825,N_15882,N_15104);
nand U16826 (N_16826,N_15274,N_15416);
nor U16827 (N_16827,N_15711,N_15226);
and U16828 (N_16828,N_15071,N_15579);
nor U16829 (N_16829,N_15002,N_15824);
nand U16830 (N_16830,N_15904,N_15921);
nand U16831 (N_16831,N_15164,N_15920);
nor U16832 (N_16832,N_15553,N_15267);
or U16833 (N_16833,N_15475,N_15286);
nand U16834 (N_16834,N_15882,N_15510);
xor U16835 (N_16835,N_15645,N_15469);
xnor U16836 (N_16836,N_15893,N_15273);
xnor U16837 (N_16837,N_15321,N_15876);
nor U16838 (N_16838,N_15621,N_15729);
xnor U16839 (N_16839,N_15609,N_15346);
and U16840 (N_16840,N_15200,N_15484);
nor U16841 (N_16841,N_15313,N_15768);
or U16842 (N_16842,N_15132,N_15624);
nor U16843 (N_16843,N_15743,N_15727);
xnor U16844 (N_16844,N_15277,N_15670);
nand U16845 (N_16845,N_15218,N_15257);
nand U16846 (N_16846,N_15054,N_15022);
or U16847 (N_16847,N_15412,N_15737);
xnor U16848 (N_16848,N_15879,N_15202);
and U16849 (N_16849,N_15631,N_15065);
or U16850 (N_16850,N_15390,N_15972);
nor U16851 (N_16851,N_15939,N_15042);
and U16852 (N_16852,N_15133,N_15497);
nor U16853 (N_16853,N_15089,N_15928);
nand U16854 (N_16854,N_15108,N_15649);
nor U16855 (N_16855,N_15951,N_15997);
xnor U16856 (N_16856,N_15110,N_15397);
or U16857 (N_16857,N_15202,N_15313);
or U16858 (N_16858,N_15336,N_15488);
and U16859 (N_16859,N_15668,N_15182);
nor U16860 (N_16860,N_15506,N_15709);
xnor U16861 (N_16861,N_15710,N_15033);
or U16862 (N_16862,N_15190,N_15836);
nor U16863 (N_16863,N_15658,N_15493);
nand U16864 (N_16864,N_15573,N_15066);
or U16865 (N_16865,N_15776,N_15248);
xor U16866 (N_16866,N_15485,N_15981);
or U16867 (N_16867,N_15582,N_15543);
or U16868 (N_16868,N_15023,N_15461);
xnor U16869 (N_16869,N_15005,N_15172);
or U16870 (N_16870,N_15872,N_15667);
nand U16871 (N_16871,N_15255,N_15604);
and U16872 (N_16872,N_15310,N_15323);
xor U16873 (N_16873,N_15513,N_15359);
nor U16874 (N_16874,N_15472,N_15986);
and U16875 (N_16875,N_15205,N_15172);
xnor U16876 (N_16876,N_15535,N_15757);
xor U16877 (N_16877,N_15744,N_15482);
and U16878 (N_16878,N_15665,N_15237);
and U16879 (N_16879,N_15868,N_15511);
and U16880 (N_16880,N_15028,N_15852);
nand U16881 (N_16881,N_15643,N_15984);
xor U16882 (N_16882,N_15382,N_15195);
nor U16883 (N_16883,N_15599,N_15662);
xnor U16884 (N_16884,N_15257,N_15937);
or U16885 (N_16885,N_15068,N_15971);
nand U16886 (N_16886,N_15723,N_15933);
nor U16887 (N_16887,N_15110,N_15368);
nand U16888 (N_16888,N_15048,N_15012);
nor U16889 (N_16889,N_15544,N_15187);
nand U16890 (N_16890,N_15595,N_15520);
and U16891 (N_16891,N_15697,N_15918);
xnor U16892 (N_16892,N_15974,N_15968);
nand U16893 (N_16893,N_15218,N_15882);
nor U16894 (N_16894,N_15246,N_15566);
nand U16895 (N_16895,N_15678,N_15196);
nand U16896 (N_16896,N_15708,N_15179);
nor U16897 (N_16897,N_15744,N_15148);
or U16898 (N_16898,N_15354,N_15883);
or U16899 (N_16899,N_15130,N_15482);
and U16900 (N_16900,N_15350,N_15454);
and U16901 (N_16901,N_15303,N_15741);
nand U16902 (N_16902,N_15775,N_15320);
and U16903 (N_16903,N_15688,N_15306);
nand U16904 (N_16904,N_15221,N_15019);
xnor U16905 (N_16905,N_15907,N_15090);
xnor U16906 (N_16906,N_15229,N_15390);
nand U16907 (N_16907,N_15869,N_15496);
xor U16908 (N_16908,N_15362,N_15131);
xor U16909 (N_16909,N_15974,N_15724);
and U16910 (N_16910,N_15901,N_15387);
or U16911 (N_16911,N_15475,N_15046);
nand U16912 (N_16912,N_15271,N_15322);
nor U16913 (N_16913,N_15762,N_15811);
nor U16914 (N_16914,N_15605,N_15730);
and U16915 (N_16915,N_15786,N_15466);
xor U16916 (N_16916,N_15924,N_15135);
nor U16917 (N_16917,N_15230,N_15329);
xor U16918 (N_16918,N_15003,N_15475);
nand U16919 (N_16919,N_15562,N_15091);
nor U16920 (N_16920,N_15587,N_15088);
xor U16921 (N_16921,N_15148,N_15542);
nand U16922 (N_16922,N_15103,N_15465);
nor U16923 (N_16923,N_15265,N_15196);
and U16924 (N_16924,N_15400,N_15000);
nand U16925 (N_16925,N_15058,N_15826);
or U16926 (N_16926,N_15177,N_15240);
or U16927 (N_16927,N_15507,N_15388);
or U16928 (N_16928,N_15947,N_15483);
nand U16929 (N_16929,N_15370,N_15210);
nand U16930 (N_16930,N_15176,N_15804);
nand U16931 (N_16931,N_15859,N_15131);
and U16932 (N_16932,N_15332,N_15709);
nor U16933 (N_16933,N_15349,N_15395);
and U16934 (N_16934,N_15727,N_15647);
xor U16935 (N_16935,N_15886,N_15976);
xor U16936 (N_16936,N_15606,N_15250);
or U16937 (N_16937,N_15713,N_15772);
nand U16938 (N_16938,N_15266,N_15955);
nor U16939 (N_16939,N_15950,N_15862);
xnor U16940 (N_16940,N_15629,N_15785);
nand U16941 (N_16941,N_15367,N_15425);
nor U16942 (N_16942,N_15396,N_15762);
xnor U16943 (N_16943,N_15042,N_15369);
and U16944 (N_16944,N_15505,N_15342);
xor U16945 (N_16945,N_15669,N_15473);
nand U16946 (N_16946,N_15190,N_15326);
nor U16947 (N_16947,N_15073,N_15377);
xor U16948 (N_16948,N_15392,N_15269);
or U16949 (N_16949,N_15944,N_15230);
and U16950 (N_16950,N_15715,N_15004);
nor U16951 (N_16951,N_15449,N_15792);
or U16952 (N_16952,N_15028,N_15670);
nand U16953 (N_16953,N_15484,N_15169);
nor U16954 (N_16954,N_15495,N_15778);
nand U16955 (N_16955,N_15986,N_15118);
nand U16956 (N_16956,N_15544,N_15485);
and U16957 (N_16957,N_15524,N_15498);
nor U16958 (N_16958,N_15389,N_15919);
or U16959 (N_16959,N_15293,N_15054);
xor U16960 (N_16960,N_15471,N_15988);
xnor U16961 (N_16961,N_15572,N_15478);
nor U16962 (N_16962,N_15762,N_15894);
nor U16963 (N_16963,N_15884,N_15601);
xnor U16964 (N_16964,N_15528,N_15322);
and U16965 (N_16965,N_15796,N_15022);
xnor U16966 (N_16966,N_15067,N_15551);
or U16967 (N_16967,N_15382,N_15519);
and U16968 (N_16968,N_15940,N_15834);
xnor U16969 (N_16969,N_15817,N_15876);
and U16970 (N_16970,N_15047,N_15800);
nand U16971 (N_16971,N_15278,N_15115);
and U16972 (N_16972,N_15816,N_15755);
nand U16973 (N_16973,N_15160,N_15548);
nand U16974 (N_16974,N_15865,N_15386);
xor U16975 (N_16975,N_15960,N_15271);
xor U16976 (N_16976,N_15592,N_15234);
or U16977 (N_16977,N_15793,N_15402);
xnor U16978 (N_16978,N_15162,N_15627);
xor U16979 (N_16979,N_15367,N_15355);
nor U16980 (N_16980,N_15566,N_15165);
nand U16981 (N_16981,N_15621,N_15772);
and U16982 (N_16982,N_15096,N_15366);
xor U16983 (N_16983,N_15772,N_15850);
and U16984 (N_16984,N_15954,N_15407);
nand U16985 (N_16985,N_15058,N_15829);
and U16986 (N_16986,N_15361,N_15951);
xor U16987 (N_16987,N_15948,N_15832);
xor U16988 (N_16988,N_15709,N_15449);
and U16989 (N_16989,N_15688,N_15390);
or U16990 (N_16990,N_15685,N_15497);
and U16991 (N_16991,N_15943,N_15455);
and U16992 (N_16992,N_15790,N_15897);
and U16993 (N_16993,N_15912,N_15166);
xor U16994 (N_16994,N_15257,N_15072);
nand U16995 (N_16995,N_15778,N_15173);
nand U16996 (N_16996,N_15763,N_15460);
nand U16997 (N_16997,N_15137,N_15650);
nand U16998 (N_16998,N_15865,N_15049);
nand U16999 (N_16999,N_15125,N_15132);
nor U17000 (N_17000,N_16343,N_16240);
or U17001 (N_17001,N_16964,N_16219);
xor U17002 (N_17002,N_16027,N_16991);
and U17003 (N_17003,N_16420,N_16811);
nor U17004 (N_17004,N_16212,N_16855);
nand U17005 (N_17005,N_16138,N_16531);
nand U17006 (N_17006,N_16644,N_16398);
nand U17007 (N_17007,N_16617,N_16028);
xor U17008 (N_17008,N_16649,N_16361);
or U17009 (N_17009,N_16836,N_16320);
and U17010 (N_17010,N_16423,N_16456);
and U17011 (N_17011,N_16419,N_16498);
nor U17012 (N_17012,N_16656,N_16799);
and U17013 (N_17013,N_16401,N_16141);
and U17014 (N_17014,N_16198,N_16001);
and U17015 (N_17015,N_16695,N_16618);
or U17016 (N_17016,N_16332,N_16462);
nand U17017 (N_17017,N_16099,N_16155);
nand U17018 (N_17018,N_16019,N_16190);
xnor U17019 (N_17019,N_16402,N_16534);
or U17020 (N_17020,N_16747,N_16338);
xnor U17021 (N_17021,N_16205,N_16725);
and U17022 (N_17022,N_16907,N_16117);
nor U17023 (N_17023,N_16951,N_16354);
or U17024 (N_17024,N_16283,N_16153);
and U17025 (N_17025,N_16883,N_16102);
nand U17026 (N_17026,N_16200,N_16700);
xor U17027 (N_17027,N_16773,N_16584);
nor U17028 (N_17028,N_16378,N_16193);
and U17029 (N_17029,N_16095,N_16923);
nor U17030 (N_17030,N_16363,N_16480);
nor U17031 (N_17031,N_16229,N_16986);
and U17032 (N_17032,N_16582,N_16526);
xnor U17033 (N_17033,N_16768,N_16552);
nand U17034 (N_17034,N_16581,N_16559);
nor U17035 (N_17035,N_16786,N_16231);
and U17036 (N_17036,N_16172,N_16440);
nor U17037 (N_17037,N_16962,N_16673);
xor U17038 (N_17038,N_16350,N_16958);
nand U17039 (N_17039,N_16566,N_16202);
nor U17040 (N_17040,N_16137,N_16128);
nand U17041 (N_17041,N_16548,N_16011);
or U17042 (N_17042,N_16988,N_16220);
nand U17043 (N_17043,N_16287,N_16792);
and U17044 (N_17044,N_16689,N_16379);
and U17045 (N_17045,N_16922,N_16245);
xnor U17046 (N_17046,N_16318,N_16371);
xor U17047 (N_17047,N_16921,N_16258);
xor U17048 (N_17048,N_16391,N_16334);
nor U17049 (N_17049,N_16643,N_16234);
nand U17050 (N_17050,N_16623,N_16632);
nand U17051 (N_17051,N_16347,N_16140);
or U17052 (N_17052,N_16262,N_16238);
nand U17053 (N_17053,N_16930,N_16257);
nand U17054 (N_17054,N_16024,N_16443);
xor U17055 (N_17055,N_16676,N_16603);
xnor U17056 (N_17056,N_16506,N_16943);
nand U17057 (N_17057,N_16520,N_16741);
nand U17058 (N_17058,N_16299,N_16235);
and U17059 (N_17059,N_16984,N_16165);
and U17060 (N_17060,N_16933,N_16226);
or U17061 (N_17061,N_16448,N_16681);
and U17062 (N_17062,N_16110,N_16939);
nor U17063 (N_17063,N_16062,N_16715);
and U17064 (N_17064,N_16641,N_16166);
or U17065 (N_17065,N_16665,N_16625);
and U17066 (N_17066,N_16090,N_16291);
xnor U17067 (N_17067,N_16055,N_16032);
nand U17068 (N_17068,N_16982,N_16216);
and U17069 (N_17069,N_16455,N_16495);
nand U17070 (N_17070,N_16127,N_16732);
nand U17071 (N_17071,N_16908,N_16413);
and U17072 (N_17072,N_16784,N_16176);
nand U17073 (N_17073,N_16282,N_16187);
nor U17074 (N_17074,N_16749,N_16123);
nand U17075 (N_17075,N_16454,N_16653);
nor U17076 (N_17076,N_16931,N_16429);
nand U17077 (N_17077,N_16453,N_16040);
nor U17078 (N_17078,N_16727,N_16925);
and U17079 (N_17079,N_16758,N_16514);
and U17080 (N_17080,N_16738,N_16094);
or U17081 (N_17081,N_16223,N_16562);
xnor U17082 (N_17082,N_16771,N_16031);
nand U17083 (N_17083,N_16828,N_16859);
or U17084 (N_17084,N_16963,N_16393);
nor U17085 (N_17085,N_16351,N_16563);
nand U17086 (N_17086,N_16979,N_16081);
xnor U17087 (N_17087,N_16913,N_16038);
and U17088 (N_17088,N_16395,N_16645);
xor U17089 (N_17089,N_16210,N_16037);
or U17090 (N_17090,N_16574,N_16048);
and U17091 (N_17091,N_16803,N_16992);
nor U17092 (N_17092,N_16826,N_16909);
nand U17093 (N_17093,N_16415,N_16161);
nand U17094 (N_17094,N_16667,N_16412);
xor U17095 (N_17095,N_16174,N_16766);
nor U17096 (N_17096,N_16899,N_16606);
xor U17097 (N_17097,N_16551,N_16249);
xnor U17098 (N_17098,N_16871,N_16565);
nand U17099 (N_17099,N_16537,N_16146);
nand U17100 (N_17100,N_16060,N_16266);
nor U17101 (N_17101,N_16575,N_16169);
or U17102 (N_17102,N_16598,N_16168);
xor U17103 (N_17103,N_16222,N_16949);
and U17104 (N_17104,N_16898,N_16276);
nand U17105 (N_17105,N_16966,N_16459);
xor U17106 (N_17106,N_16693,N_16634);
xor U17107 (N_17107,N_16724,N_16313);
nand U17108 (N_17108,N_16017,N_16154);
nand U17109 (N_17109,N_16900,N_16466);
nor U17110 (N_17110,N_16564,N_16004);
nor U17111 (N_17111,N_16033,N_16373);
or U17112 (N_17112,N_16678,N_16543);
nand U17113 (N_17113,N_16116,N_16492);
and U17114 (N_17114,N_16630,N_16967);
nor U17115 (N_17115,N_16869,N_16344);
nor U17116 (N_17116,N_16611,N_16906);
nor U17117 (N_17117,N_16449,N_16818);
nand U17118 (N_17118,N_16788,N_16109);
nand U17119 (N_17119,N_16920,N_16845);
nor U17120 (N_17120,N_16330,N_16089);
or U17121 (N_17121,N_16669,N_16701);
xnor U17122 (N_17122,N_16263,N_16853);
xnor U17123 (N_17123,N_16144,N_16542);
xor U17124 (N_17124,N_16185,N_16399);
xnor U17125 (N_17125,N_16787,N_16614);
and U17126 (N_17126,N_16152,N_16721);
and U17127 (N_17127,N_16577,N_16983);
nor U17128 (N_17128,N_16801,N_16971);
nand U17129 (N_17129,N_16252,N_16754);
xor U17130 (N_17130,N_16892,N_16636);
xor U17131 (N_17131,N_16802,N_16135);
nor U17132 (N_17132,N_16328,N_16533);
nand U17133 (N_17133,N_16915,N_16954);
and U17134 (N_17134,N_16477,N_16877);
or U17135 (N_17135,N_16919,N_16195);
nand U17136 (N_17136,N_16184,N_16280);
or U17137 (N_17137,N_16308,N_16126);
or U17138 (N_17138,N_16326,N_16355);
or U17139 (N_17139,N_16389,N_16481);
or U17140 (N_17140,N_16147,N_16905);
nand U17141 (N_17141,N_16647,N_16255);
or U17142 (N_17142,N_16471,N_16854);
or U17143 (N_17143,N_16886,N_16101);
nor U17144 (N_17144,N_16230,N_16006);
nand U17145 (N_17145,N_16894,N_16013);
and U17146 (N_17146,N_16503,N_16160);
and U17147 (N_17147,N_16635,N_16834);
and U17148 (N_17148,N_16705,N_16938);
nand U17149 (N_17149,N_16820,N_16839);
or U17150 (N_17150,N_16627,N_16404);
and U17151 (N_17151,N_16694,N_16056);
and U17152 (N_17152,N_16717,N_16029);
xnor U17153 (N_17153,N_16832,N_16806);
nand U17154 (N_17154,N_16867,N_16528);
nand U17155 (N_17155,N_16163,N_16065);
or U17156 (N_17156,N_16438,N_16122);
and U17157 (N_17157,N_16968,N_16781);
nand U17158 (N_17158,N_16848,N_16484);
xor U17159 (N_17159,N_16396,N_16989);
xor U17160 (N_17160,N_16505,N_16063);
nor U17161 (N_17161,N_16619,N_16868);
nand U17162 (N_17162,N_16596,N_16850);
nand U17163 (N_17163,N_16239,N_16969);
nand U17164 (N_17164,N_16782,N_16622);
nand U17165 (N_17165,N_16458,N_16762);
xor U17166 (N_17166,N_16208,N_16953);
xor U17167 (N_17167,N_16247,N_16586);
nor U17168 (N_17168,N_16433,N_16474);
nor U17169 (N_17169,N_16432,N_16483);
or U17170 (N_17170,N_16544,N_16527);
xnor U17171 (N_17171,N_16279,N_16307);
and U17172 (N_17172,N_16648,N_16324);
xor U17173 (N_17173,N_16881,N_16259);
nand U17174 (N_17174,N_16468,N_16436);
and U17175 (N_17175,N_16446,N_16250);
nand U17176 (N_17176,N_16746,N_16796);
and U17177 (N_17177,N_16382,N_16517);
nand U17178 (N_17178,N_16729,N_16524);
xnor U17179 (N_17179,N_16595,N_16589);
and U17180 (N_17180,N_16192,N_16680);
and U17181 (N_17181,N_16417,N_16134);
xnor U17182 (N_17182,N_16677,N_16772);
nor U17183 (N_17183,N_16713,N_16975);
and U17184 (N_17184,N_16021,N_16815);
nor U17185 (N_17185,N_16639,N_16445);
nor U17186 (N_17186,N_16831,N_16369);
and U17187 (N_17187,N_16692,N_16493);
or U17188 (N_17188,N_16884,N_16604);
nand U17189 (N_17189,N_16108,N_16268);
and U17190 (N_17190,N_16558,N_16740);
xor U17191 (N_17191,N_16366,N_16844);
xnor U17192 (N_17192,N_16149,N_16173);
xnor U17193 (N_17193,N_16421,N_16810);
and U17194 (N_17194,N_16540,N_16856);
xnor U17195 (N_17195,N_16509,N_16360);
or U17196 (N_17196,N_16491,N_16435);
nand U17197 (N_17197,N_16336,N_16197);
and U17198 (N_17198,N_16260,N_16111);
nand U17199 (N_17199,N_16053,N_16057);
nor U17200 (N_17200,N_16388,N_16585);
or U17201 (N_17201,N_16036,N_16182);
nor U17202 (N_17202,N_16816,N_16221);
or U17203 (N_17203,N_16242,N_16698);
nand U17204 (N_17204,N_16916,N_16594);
nor U17205 (N_17205,N_16621,N_16039);
and U17206 (N_17206,N_16885,N_16774);
nor U17207 (N_17207,N_16880,N_16071);
nand U17208 (N_17208,N_16105,N_16025);
and U17209 (N_17209,N_16708,N_16946);
nand U17210 (N_17210,N_16206,N_16246);
or U17211 (N_17211,N_16107,N_16823);
or U17212 (N_17212,N_16339,N_16901);
nand U17213 (N_17213,N_16284,N_16450);
and U17214 (N_17214,N_16115,N_16012);
nor U17215 (N_17215,N_16346,N_16077);
xnor U17216 (N_17216,N_16078,N_16605);
and U17217 (N_17217,N_16007,N_16319);
or U17218 (N_17218,N_16789,N_16191);
nor U17219 (N_17219,N_16237,N_16515);
nand U17220 (N_17220,N_16341,N_16261);
xnor U17221 (N_17221,N_16479,N_16735);
nor U17222 (N_17222,N_16298,N_16325);
nor U17223 (N_17223,N_16858,N_16985);
nand U17224 (N_17224,N_16835,N_16422);
and U17225 (N_17225,N_16857,N_16655);
xor U17226 (N_17226,N_16304,N_16273);
xor U17227 (N_17227,N_16118,N_16322);
nor U17228 (N_17228,N_16893,N_16819);
nand U17229 (N_17229,N_16800,N_16508);
nor U17230 (N_17230,N_16720,N_16935);
xor U17231 (N_17231,N_16485,N_16872);
xnor U17232 (N_17232,N_16306,N_16075);
nor U17233 (N_17233,N_16447,N_16638);
nor U17234 (N_17234,N_16662,N_16164);
nor U17235 (N_17235,N_16996,N_16793);
nor U17236 (N_17236,N_16500,N_16317);
nand U17237 (N_17237,N_16873,N_16403);
nor U17238 (N_17238,N_16797,N_16430);
xnor U17239 (N_17239,N_16532,N_16887);
or U17240 (N_17240,N_16437,N_16312);
and U17241 (N_17241,N_16309,N_16974);
nand U17242 (N_17242,N_16119,N_16794);
and U17243 (N_17243,N_16333,N_16487);
xor U17244 (N_17244,N_16546,N_16947);
xnor U17245 (N_17245,N_16664,N_16241);
and U17246 (N_17246,N_16381,N_16377);
nand U17247 (N_17247,N_16730,N_16757);
and U17248 (N_17248,N_16688,N_16136);
nand U17249 (N_17249,N_16697,N_16442);
or U17250 (N_17250,N_16051,N_16895);
nor U17251 (N_17251,N_16209,N_16156);
xnor U17252 (N_17252,N_16467,N_16215);
or U17253 (N_17253,N_16743,N_16295);
and U17254 (N_17254,N_16650,N_16159);
nand U17255 (N_17255,N_16798,N_16896);
nand U17256 (N_17256,N_16023,N_16386);
xnor U17257 (N_17257,N_16561,N_16504);
and U17258 (N_17258,N_16084,N_16070);
nor U17259 (N_17259,N_16554,N_16568);
nor U17260 (N_17260,N_16670,N_16457);
and U17261 (N_17261,N_16227,N_16349);
nor U17262 (N_17262,N_16271,N_16759);
or U17263 (N_17263,N_16296,N_16890);
nor U17264 (N_17264,N_16671,N_16243);
and U17265 (N_17265,N_16311,N_16960);
nand U17266 (N_17266,N_16726,N_16411);
and U17267 (N_17267,N_16734,N_16936);
or U17268 (N_17268,N_16805,N_16005);
xnor U17269 (N_17269,N_16015,N_16288);
nand U17270 (N_17270,N_16463,N_16008);
and U17271 (N_17271,N_16742,N_16824);
nand U17272 (N_17272,N_16129,N_16876);
and U17273 (N_17273,N_16516,N_16384);
and U17274 (N_17274,N_16218,N_16042);
xor U17275 (N_17275,N_16833,N_16082);
xor U17276 (N_17276,N_16009,N_16994);
or U17277 (N_17277,N_16977,N_16054);
nor U17278 (N_17278,N_16150,N_16602);
xnor U17279 (N_17279,N_16254,N_16633);
and U17280 (N_17280,N_16686,N_16882);
nor U17281 (N_17281,N_16167,N_16668);
xor U17282 (N_17282,N_16593,N_16010);
xnor U17283 (N_17283,N_16764,N_16460);
nor U17284 (N_17284,N_16014,N_16753);
nor U17285 (N_17285,N_16236,N_16583);
xnor U17286 (N_17286,N_16539,N_16264);
nand U17287 (N_17287,N_16244,N_16289);
and U17288 (N_17288,N_16521,N_16934);
nor U17289 (N_17289,N_16225,N_16170);
or U17290 (N_17290,N_16911,N_16426);
xnor U17291 (N_17291,N_16441,N_16745);
xor U17292 (N_17292,N_16512,N_16696);
nand U17293 (N_17293,N_16093,N_16924);
xnor U17294 (N_17294,N_16203,N_16706);
nand U17295 (N_17295,N_16044,N_16294);
xor U17296 (N_17296,N_16874,N_16045);
nor U17297 (N_17297,N_16987,N_16112);
nor U17298 (N_17298,N_16778,N_16470);
and U17299 (N_17299,N_16465,N_16748);
nor U17300 (N_17300,N_16972,N_16059);
nand U17301 (N_17301,N_16702,N_16751);
and U17302 (N_17302,N_16145,N_16875);
and U17303 (N_17303,N_16997,N_16711);
and U17304 (N_17304,N_16494,N_16719);
nor U17305 (N_17305,N_16265,N_16682);
and U17306 (N_17306,N_16385,N_16941);
nand U17307 (N_17307,N_16945,N_16530);
and U17308 (N_17308,N_16770,N_16348);
nand U17309 (N_17309,N_16572,N_16817);
nand U17310 (N_17310,N_16335,N_16612);
nand U17311 (N_17311,N_16106,N_16587);
nand U17312 (N_17312,N_16407,N_16926);
xor U17313 (N_17313,N_16416,N_16502);
xor U17314 (N_17314,N_16376,N_16849);
xnor U17315 (N_17315,N_16124,N_16175);
and U17316 (N_17316,N_16620,N_16889);
nor U17317 (N_17317,N_16529,N_16434);
or U17318 (N_17318,N_16940,N_16590);
nor U17319 (N_17319,N_16808,N_16469);
nor U17320 (N_17320,N_16928,N_16570);
or U17321 (N_17321,N_16651,N_16097);
xor U17322 (N_17322,N_16690,N_16576);
nor U17323 (N_17323,N_16663,N_16121);
or U17324 (N_17324,N_16364,N_16418);
nor U17325 (N_17325,N_16567,N_16478);
xnor U17326 (N_17326,N_16888,N_16684);
nor U17327 (N_17327,N_16660,N_16034);
xnor U17328 (N_17328,N_16948,N_16368);
nand U17329 (N_17329,N_16251,N_16609);
nor U17330 (N_17330,N_16098,N_16879);
nand U17331 (N_17331,N_16253,N_16281);
and U17332 (N_17332,N_16375,N_16973);
nand U17333 (N_17333,N_16113,N_16302);
or U17334 (N_17334,N_16902,N_16327);
nand U17335 (N_17335,N_16813,N_16847);
xor U17336 (N_17336,N_16878,N_16535);
or U17337 (N_17337,N_16995,N_16072);
or U17338 (N_17338,N_16409,N_16359);
nor U17339 (N_17339,N_16672,N_16976);
or U17340 (N_17340,N_16486,N_16091);
nand U17341 (N_17341,N_16511,N_16088);
nor U17342 (N_17342,N_16659,N_16761);
nand U17343 (N_17343,N_16571,N_16917);
nand U17344 (N_17344,N_16016,N_16204);
xnor U17345 (N_17345,N_16750,N_16704);
or U17346 (N_17346,N_16728,N_16536);
nand U17347 (N_17347,N_16104,N_16709);
nand U17348 (N_17348,N_16425,N_16188);
nor U17349 (N_17349,N_16591,N_16497);
or U17350 (N_17350,N_16270,N_16046);
nand U17351 (N_17351,N_16103,N_16840);
nand U17352 (N_17352,N_16523,N_16599);
nor U17353 (N_17353,N_16990,N_16085);
or U17354 (N_17354,N_16980,N_16499);
xor U17355 (N_17355,N_16224,N_16323);
nand U17356 (N_17356,N_16942,N_16999);
or U17357 (N_17357,N_16712,N_16998);
and U17358 (N_17358,N_16356,N_16739);
and U17359 (N_17359,N_16691,N_16353);
and U17360 (N_17360,N_16214,N_16233);
xor U17361 (N_17361,N_16841,N_16130);
and U17362 (N_17362,N_16866,N_16560);
nor U17363 (N_17363,N_16277,N_16052);
nand U17364 (N_17364,N_16944,N_16213);
and U17365 (N_17365,N_16316,N_16358);
and U17366 (N_17366,N_16297,N_16755);
and U17367 (N_17367,N_16143,N_16374);
nor U17368 (N_17368,N_16272,N_16752);
xnor U17369 (N_17369,N_16232,N_16580);
and U17370 (N_17370,N_16707,N_16910);
and U17371 (N_17371,N_16699,N_16079);
or U17372 (N_17372,N_16822,N_16785);
nand U17373 (N_17373,N_16406,N_16020);
nand U17374 (N_17374,N_16870,N_16201);
or U17375 (N_17375,N_16783,N_16763);
nor U17376 (N_17376,N_16362,N_16965);
and U17377 (N_17377,N_16342,N_16380);
nor U17378 (N_17378,N_16452,N_16929);
and U17379 (N_17379,N_16891,N_16613);
nand U17380 (N_17380,N_16600,N_16812);
nor U17381 (N_17381,N_16158,N_16331);
or U17382 (N_17382,N_16597,N_16744);
and U17383 (N_17383,N_16685,N_16439);
and U17384 (N_17384,N_16809,N_16863);
and U17385 (N_17385,N_16714,N_16851);
nor U17386 (N_17386,N_16303,N_16372);
xor U17387 (N_17387,N_16767,N_16186);
xnor U17388 (N_17388,N_16687,N_16838);
xnor U17389 (N_17389,N_16952,N_16675);
xor U17390 (N_17390,N_16357,N_16860);
xor U17391 (N_17391,N_16610,N_16424);
nor U17392 (N_17392,N_16049,N_16776);
xor U17393 (N_17393,N_16657,N_16041);
xor U17394 (N_17394,N_16476,N_16047);
nand U17395 (N_17395,N_16285,N_16189);
nor U17396 (N_17396,N_16064,N_16955);
or U17397 (N_17397,N_16069,N_16628);
xnor U17398 (N_17398,N_16703,N_16807);
or U17399 (N_17399,N_16865,N_16228);
nor U17400 (N_17400,N_16043,N_16067);
and U17401 (N_17401,N_16756,N_16464);
and U17402 (N_17402,N_16179,N_16180);
and U17403 (N_17403,N_16829,N_16427);
xnor U17404 (N_17404,N_16086,N_16557);
nand U17405 (N_17405,N_16092,N_16814);
or U17406 (N_17406,N_16482,N_16646);
and U17407 (N_17407,N_16340,N_16207);
nand U17408 (N_17408,N_16269,N_16821);
nand U17409 (N_17409,N_16181,N_16830);
or U17410 (N_17410,N_16631,N_16003);
and U17411 (N_17411,N_16862,N_16142);
and U17412 (N_17412,N_16337,N_16970);
xor U17413 (N_17413,N_16087,N_16608);
xor U17414 (N_17414,N_16777,N_16300);
xnor U17415 (N_17415,N_16588,N_16837);
and U17416 (N_17416,N_16428,N_16592);
xnor U17417 (N_17417,N_16292,N_16267);
or U17418 (N_17418,N_16733,N_16791);
nand U17419 (N_17419,N_16489,N_16408);
xor U17420 (N_17420,N_16329,N_16932);
nand U17421 (N_17421,N_16274,N_16993);
xnor U17422 (N_17422,N_16293,N_16652);
nand U17423 (N_17423,N_16321,N_16978);
and U17424 (N_17424,N_16400,N_16120);
nor U17425 (N_17425,N_16765,N_16139);
and U17426 (N_17426,N_16654,N_16475);
and U17427 (N_17427,N_16956,N_16914);
or U17428 (N_17428,N_16790,N_16710);
and U17429 (N_17429,N_16780,N_16035);
or U17430 (N_17430,N_16444,N_16278);
nor U17431 (N_17431,N_16513,N_16000);
or U17432 (N_17432,N_16579,N_16405);
or U17433 (N_17433,N_16100,N_16096);
nor U17434 (N_17434,N_16961,N_16125);
or U17435 (N_17435,N_16640,N_16383);
nand U17436 (N_17436,N_16488,N_16177);
or U17437 (N_17437,N_16769,N_16074);
xor U17438 (N_17438,N_16080,N_16301);
and U17439 (N_17439,N_16286,N_16151);
nor U17440 (N_17440,N_16852,N_16957);
nand U17441 (N_17441,N_16083,N_16183);
or U17442 (N_17442,N_16556,N_16666);
xor U17443 (N_17443,N_16199,N_16290);
or U17444 (N_17444,N_16843,N_16629);
nand U17445 (N_17445,N_16392,N_16904);
xnor U17446 (N_17446,N_16981,N_16217);
xor U17447 (N_17447,N_16545,N_16394);
nor U17448 (N_17448,N_16365,N_16553);
and U17449 (N_17449,N_16196,N_16722);
xor U17450 (N_17450,N_16541,N_16737);
xnor U17451 (N_17451,N_16061,N_16842);
nand U17452 (N_17452,N_16736,N_16030);
nor U17453 (N_17453,N_16507,N_16637);
or U17454 (N_17454,N_16148,N_16370);
nand U17455 (N_17455,N_16002,N_16804);
nor U17456 (N_17456,N_16937,N_16194);
or U17457 (N_17457,N_16679,N_16918);
nand U17458 (N_17458,N_16473,N_16133);
nand U17459 (N_17459,N_16731,N_16472);
and U17460 (N_17460,N_16305,N_16315);
xnor U17461 (N_17461,N_16275,N_16518);
nor U17462 (N_17462,N_16601,N_16683);
nand U17463 (N_17463,N_16171,N_16490);
or U17464 (N_17464,N_16775,N_16076);
or U17465 (N_17465,N_16897,N_16397);
xnor U17466 (N_17466,N_16779,N_16626);
or U17467 (N_17467,N_16912,N_16607);
xnor U17468 (N_17468,N_16538,N_16352);
nand U17469 (N_17469,N_16825,N_16018);
nand U17470 (N_17470,N_16861,N_16501);
nor U17471 (N_17471,N_16431,N_16496);
nand U17472 (N_17472,N_16616,N_16624);
or U17473 (N_17473,N_16510,N_16723);
and U17474 (N_17474,N_16959,N_16345);
nor U17475 (N_17475,N_16555,N_16310);
or U17476 (N_17476,N_16950,N_16066);
xnor U17477 (N_17477,N_16795,N_16578);
and U17478 (N_17478,N_16573,N_16314);
or U17479 (N_17479,N_16550,N_16569);
and U17480 (N_17480,N_16927,N_16661);
nor U17481 (N_17481,N_16718,N_16050);
xnor U17482 (N_17482,N_16864,N_16642);
nand U17483 (N_17483,N_16827,N_16451);
nor U17484 (N_17484,N_16525,N_16760);
or U17485 (N_17485,N_16132,N_16615);
and U17486 (N_17486,N_16022,N_16178);
nor U17487 (N_17487,N_16256,N_16461);
or U17488 (N_17488,N_16410,N_16367);
or U17489 (N_17489,N_16549,N_16131);
and U17490 (N_17490,N_16519,N_16157);
nor U17491 (N_17491,N_16846,N_16073);
nor U17492 (N_17492,N_16674,N_16387);
nor U17493 (N_17493,N_16026,N_16068);
nand U17494 (N_17494,N_16658,N_16058);
or U17495 (N_17495,N_16716,N_16162);
nor U17496 (N_17496,N_16114,N_16547);
xnor U17497 (N_17497,N_16903,N_16522);
or U17498 (N_17498,N_16248,N_16211);
xor U17499 (N_17499,N_16414,N_16390);
nand U17500 (N_17500,N_16649,N_16552);
xor U17501 (N_17501,N_16224,N_16052);
xnor U17502 (N_17502,N_16842,N_16253);
xor U17503 (N_17503,N_16168,N_16328);
nor U17504 (N_17504,N_16040,N_16238);
and U17505 (N_17505,N_16733,N_16859);
or U17506 (N_17506,N_16855,N_16108);
nor U17507 (N_17507,N_16881,N_16116);
nor U17508 (N_17508,N_16316,N_16836);
or U17509 (N_17509,N_16002,N_16319);
nand U17510 (N_17510,N_16657,N_16000);
and U17511 (N_17511,N_16259,N_16857);
nor U17512 (N_17512,N_16426,N_16470);
xor U17513 (N_17513,N_16294,N_16076);
nand U17514 (N_17514,N_16134,N_16075);
nand U17515 (N_17515,N_16392,N_16469);
nand U17516 (N_17516,N_16012,N_16680);
xor U17517 (N_17517,N_16165,N_16215);
xor U17518 (N_17518,N_16078,N_16069);
nor U17519 (N_17519,N_16292,N_16328);
nand U17520 (N_17520,N_16222,N_16786);
xor U17521 (N_17521,N_16391,N_16312);
xor U17522 (N_17522,N_16926,N_16607);
nor U17523 (N_17523,N_16374,N_16773);
nor U17524 (N_17524,N_16953,N_16369);
nand U17525 (N_17525,N_16258,N_16164);
nor U17526 (N_17526,N_16012,N_16344);
xnor U17527 (N_17527,N_16733,N_16634);
xnor U17528 (N_17528,N_16045,N_16721);
nor U17529 (N_17529,N_16992,N_16851);
and U17530 (N_17530,N_16621,N_16209);
nor U17531 (N_17531,N_16554,N_16582);
or U17532 (N_17532,N_16049,N_16469);
or U17533 (N_17533,N_16243,N_16093);
and U17534 (N_17534,N_16106,N_16363);
or U17535 (N_17535,N_16508,N_16598);
xor U17536 (N_17536,N_16485,N_16315);
nor U17537 (N_17537,N_16650,N_16936);
nand U17538 (N_17538,N_16540,N_16329);
nand U17539 (N_17539,N_16902,N_16058);
nand U17540 (N_17540,N_16618,N_16357);
or U17541 (N_17541,N_16992,N_16282);
or U17542 (N_17542,N_16458,N_16447);
nand U17543 (N_17543,N_16193,N_16089);
nor U17544 (N_17544,N_16608,N_16835);
and U17545 (N_17545,N_16769,N_16869);
nor U17546 (N_17546,N_16281,N_16154);
nor U17547 (N_17547,N_16418,N_16221);
nor U17548 (N_17548,N_16738,N_16588);
and U17549 (N_17549,N_16473,N_16598);
or U17550 (N_17550,N_16926,N_16340);
xor U17551 (N_17551,N_16401,N_16368);
xnor U17552 (N_17552,N_16409,N_16328);
nand U17553 (N_17553,N_16073,N_16472);
xor U17554 (N_17554,N_16463,N_16855);
or U17555 (N_17555,N_16767,N_16172);
and U17556 (N_17556,N_16061,N_16106);
and U17557 (N_17557,N_16977,N_16985);
xnor U17558 (N_17558,N_16476,N_16930);
or U17559 (N_17559,N_16351,N_16524);
and U17560 (N_17560,N_16629,N_16251);
and U17561 (N_17561,N_16507,N_16719);
and U17562 (N_17562,N_16832,N_16011);
or U17563 (N_17563,N_16151,N_16751);
nor U17564 (N_17564,N_16673,N_16943);
and U17565 (N_17565,N_16253,N_16919);
nand U17566 (N_17566,N_16544,N_16845);
xor U17567 (N_17567,N_16753,N_16824);
or U17568 (N_17568,N_16605,N_16178);
or U17569 (N_17569,N_16994,N_16482);
or U17570 (N_17570,N_16237,N_16045);
nor U17571 (N_17571,N_16882,N_16710);
xnor U17572 (N_17572,N_16168,N_16860);
or U17573 (N_17573,N_16675,N_16153);
nand U17574 (N_17574,N_16651,N_16666);
or U17575 (N_17575,N_16029,N_16371);
and U17576 (N_17576,N_16318,N_16605);
xnor U17577 (N_17577,N_16649,N_16631);
nand U17578 (N_17578,N_16186,N_16655);
or U17579 (N_17579,N_16747,N_16830);
nand U17580 (N_17580,N_16604,N_16874);
and U17581 (N_17581,N_16463,N_16579);
or U17582 (N_17582,N_16944,N_16867);
nor U17583 (N_17583,N_16991,N_16901);
and U17584 (N_17584,N_16660,N_16402);
nor U17585 (N_17585,N_16008,N_16777);
nand U17586 (N_17586,N_16495,N_16769);
nor U17587 (N_17587,N_16881,N_16068);
nor U17588 (N_17588,N_16095,N_16364);
nor U17589 (N_17589,N_16063,N_16081);
or U17590 (N_17590,N_16125,N_16068);
nand U17591 (N_17591,N_16368,N_16295);
or U17592 (N_17592,N_16438,N_16777);
and U17593 (N_17593,N_16080,N_16276);
or U17594 (N_17594,N_16935,N_16822);
and U17595 (N_17595,N_16012,N_16510);
nand U17596 (N_17596,N_16125,N_16562);
or U17597 (N_17597,N_16806,N_16293);
nand U17598 (N_17598,N_16138,N_16095);
nand U17599 (N_17599,N_16397,N_16052);
nor U17600 (N_17600,N_16558,N_16791);
nor U17601 (N_17601,N_16069,N_16117);
or U17602 (N_17602,N_16330,N_16226);
or U17603 (N_17603,N_16215,N_16306);
or U17604 (N_17604,N_16193,N_16985);
or U17605 (N_17605,N_16026,N_16491);
nand U17606 (N_17606,N_16195,N_16713);
nor U17607 (N_17607,N_16287,N_16867);
or U17608 (N_17608,N_16202,N_16494);
nor U17609 (N_17609,N_16827,N_16020);
or U17610 (N_17610,N_16676,N_16293);
or U17611 (N_17611,N_16005,N_16273);
xor U17612 (N_17612,N_16281,N_16606);
and U17613 (N_17613,N_16784,N_16229);
and U17614 (N_17614,N_16625,N_16461);
or U17615 (N_17615,N_16907,N_16865);
nand U17616 (N_17616,N_16095,N_16341);
nand U17617 (N_17617,N_16118,N_16008);
xnor U17618 (N_17618,N_16548,N_16119);
nor U17619 (N_17619,N_16513,N_16691);
or U17620 (N_17620,N_16324,N_16413);
nor U17621 (N_17621,N_16983,N_16151);
nor U17622 (N_17622,N_16203,N_16449);
or U17623 (N_17623,N_16354,N_16861);
xnor U17624 (N_17624,N_16826,N_16699);
nor U17625 (N_17625,N_16162,N_16980);
nor U17626 (N_17626,N_16365,N_16603);
or U17627 (N_17627,N_16656,N_16768);
nand U17628 (N_17628,N_16324,N_16063);
and U17629 (N_17629,N_16251,N_16431);
and U17630 (N_17630,N_16690,N_16694);
nor U17631 (N_17631,N_16902,N_16224);
nand U17632 (N_17632,N_16120,N_16428);
or U17633 (N_17633,N_16828,N_16474);
nor U17634 (N_17634,N_16660,N_16700);
xor U17635 (N_17635,N_16163,N_16352);
nor U17636 (N_17636,N_16421,N_16744);
nor U17637 (N_17637,N_16822,N_16720);
nand U17638 (N_17638,N_16523,N_16441);
nand U17639 (N_17639,N_16378,N_16329);
nand U17640 (N_17640,N_16206,N_16885);
xor U17641 (N_17641,N_16548,N_16490);
or U17642 (N_17642,N_16999,N_16680);
or U17643 (N_17643,N_16648,N_16880);
or U17644 (N_17644,N_16353,N_16431);
xor U17645 (N_17645,N_16647,N_16898);
xor U17646 (N_17646,N_16497,N_16058);
nor U17647 (N_17647,N_16929,N_16010);
xor U17648 (N_17648,N_16028,N_16411);
nor U17649 (N_17649,N_16483,N_16036);
or U17650 (N_17650,N_16516,N_16716);
or U17651 (N_17651,N_16055,N_16976);
nor U17652 (N_17652,N_16340,N_16391);
and U17653 (N_17653,N_16813,N_16124);
nand U17654 (N_17654,N_16206,N_16111);
or U17655 (N_17655,N_16114,N_16253);
or U17656 (N_17656,N_16831,N_16005);
xor U17657 (N_17657,N_16237,N_16131);
or U17658 (N_17658,N_16666,N_16047);
or U17659 (N_17659,N_16391,N_16637);
nor U17660 (N_17660,N_16307,N_16206);
xor U17661 (N_17661,N_16622,N_16114);
or U17662 (N_17662,N_16808,N_16491);
xnor U17663 (N_17663,N_16674,N_16618);
nand U17664 (N_17664,N_16695,N_16057);
nor U17665 (N_17665,N_16255,N_16803);
and U17666 (N_17666,N_16211,N_16022);
xor U17667 (N_17667,N_16904,N_16453);
nor U17668 (N_17668,N_16895,N_16614);
xnor U17669 (N_17669,N_16948,N_16852);
nor U17670 (N_17670,N_16756,N_16151);
and U17671 (N_17671,N_16293,N_16386);
or U17672 (N_17672,N_16054,N_16940);
or U17673 (N_17673,N_16554,N_16669);
xor U17674 (N_17674,N_16351,N_16750);
and U17675 (N_17675,N_16293,N_16232);
and U17676 (N_17676,N_16514,N_16512);
xnor U17677 (N_17677,N_16386,N_16588);
nand U17678 (N_17678,N_16644,N_16956);
and U17679 (N_17679,N_16986,N_16057);
or U17680 (N_17680,N_16994,N_16786);
xor U17681 (N_17681,N_16147,N_16451);
nand U17682 (N_17682,N_16608,N_16526);
and U17683 (N_17683,N_16854,N_16959);
and U17684 (N_17684,N_16215,N_16976);
nor U17685 (N_17685,N_16048,N_16866);
nand U17686 (N_17686,N_16572,N_16779);
xnor U17687 (N_17687,N_16420,N_16674);
or U17688 (N_17688,N_16969,N_16613);
nor U17689 (N_17689,N_16220,N_16086);
and U17690 (N_17690,N_16263,N_16233);
xor U17691 (N_17691,N_16398,N_16524);
nand U17692 (N_17692,N_16014,N_16790);
xnor U17693 (N_17693,N_16642,N_16046);
xnor U17694 (N_17694,N_16962,N_16787);
nand U17695 (N_17695,N_16262,N_16081);
nor U17696 (N_17696,N_16101,N_16304);
xor U17697 (N_17697,N_16814,N_16981);
and U17698 (N_17698,N_16122,N_16047);
nor U17699 (N_17699,N_16020,N_16246);
nand U17700 (N_17700,N_16652,N_16018);
or U17701 (N_17701,N_16849,N_16802);
nand U17702 (N_17702,N_16027,N_16941);
nand U17703 (N_17703,N_16549,N_16995);
and U17704 (N_17704,N_16296,N_16216);
xor U17705 (N_17705,N_16514,N_16701);
nand U17706 (N_17706,N_16908,N_16525);
or U17707 (N_17707,N_16656,N_16262);
nor U17708 (N_17708,N_16500,N_16072);
nor U17709 (N_17709,N_16620,N_16078);
or U17710 (N_17710,N_16954,N_16221);
or U17711 (N_17711,N_16227,N_16650);
xnor U17712 (N_17712,N_16727,N_16340);
or U17713 (N_17713,N_16544,N_16139);
nor U17714 (N_17714,N_16005,N_16724);
xor U17715 (N_17715,N_16873,N_16028);
or U17716 (N_17716,N_16285,N_16240);
nand U17717 (N_17717,N_16110,N_16897);
and U17718 (N_17718,N_16805,N_16213);
or U17719 (N_17719,N_16195,N_16292);
nor U17720 (N_17720,N_16001,N_16221);
xor U17721 (N_17721,N_16518,N_16837);
or U17722 (N_17722,N_16677,N_16417);
and U17723 (N_17723,N_16579,N_16114);
nor U17724 (N_17724,N_16584,N_16281);
xor U17725 (N_17725,N_16442,N_16666);
nand U17726 (N_17726,N_16507,N_16762);
or U17727 (N_17727,N_16457,N_16775);
nand U17728 (N_17728,N_16713,N_16742);
nor U17729 (N_17729,N_16051,N_16306);
nor U17730 (N_17730,N_16085,N_16177);
and U17731 (N_17731,N_16333,N_16039);
or U17732 (N_17732,N_16443,N_16576);
nor U17733 (N_17733,N_16653,N_16849);
nand U17734 (N_17734,N_16599,N_16921);
and U17735 (N_17735,N_16768,N_16758);
nand U17736 (N_17736,N_16971,N_16552);
nand U17737 (N_17737,N_16893,N_16897);
nand U17738 (N_17738,N_16838,N_16362);
xnor U17739 (N_17739,N_16064,N_16740);
nor U17740 (N_17740,N_16242,N_16894);
or U17741 (N_17741,N_16483,N_16008);
and U17742 (N_17742,N_16098,N_16910);
nand U17743 (N_17743,N_16709,N_16434);
xor U17744 (N_17744,N_16608,N_16338);
xnor U17745 (N_17745,N_16574,N_16879);
and U17746 (N_17746,N_16507,N_16737);
and U17747 (N_17747,N_16111,N_16239);
nand U17748 (N_17748,N_16312,N_16633);
nor U17749 (N_17749,N_16481,N_16554);
nor U17750 (N_17750,N_16835,N_16960);
or U17751 (N_17751,N_16451,N_16590);
or U17752 (N_17752,N_16828,N_16440);
nor U17753 (N_17753,N_16286,N_16528);
or U17754 (N_17754,N_16853,N_16460);
nand U17755 (N_17755,N_16907,N_16823);
and U17756 (N_17756,N_16384,N_16315);
and U17757 (N_17757,N_16074,N_16505);
xor U17758 (N_17758,N_16592,N_16065);
xnor U17759 (N_17759,N_16472,N_16981);
nand U17760 (N_17760,N_16053,N_16626);
and U17761 (N_17761,N_16239,N_16306);
and U17762 (N_17762,N_16553,N_16035);
nor U17763 (N_17763,N_16373,N_16395);
or U17764 (N_17764,N_16394,N_16188);
nand U17765 (N_17765,N_16770,N_16411);
nor U17766 (N_17766,N_16985,N_16719);
or U17767 (N_17767,N_16984,N_16595);
and U17768 (N_17768,N_16662,N_16466);
nor U17769 (N_17769,N_16927,N_16083);
and U17770 (N_17770,N_16937,N_16849);
nand U17771 (N_17771,N_16102,N_16494);
nand U17772 (N_17772,N_16945,N_16018);
nor U17773 (N_17773,N_16400,N_16822);
nand U17774 (N_17774,N_16769,N_16337);
or U17775 (N_17775,N_16119,N_16785);
and U17776 (N_17776,N_16838,N_16134);
nor U17777 (N_17777,N_16757,N_16512);
nor U17778 (N_17778,N_16608,N_16486);
or U17779 (N_17779,N_16937,N_16325);
and U17780 (N_17780,N_16676,N_16645);
nand U17781 (N_17781,N_16013,N_16730);
nand U17782 (N_17782,N_16188,N_16416);
and U17783 (N_17783,N_16789,N_16268);
or U17784 (N_17784,N_16714,N_16589);
xor U17785 (N_17785,N_16231,N_16395);
nand U17786 (N_17786,N_16640,N_16820);
and U17787 (N_17787,N_16774,N_16249);
nor U17788 (N_17788,N_16051,N_16795);
and U17789 (N_17789,N_16125,N_16965);
nor U17790 (N_17790,N_16921,N_16894);
nand U17791 (N_17791,N_16329,N_16708);
nor U17792 (N_17792,N_16755,N_16302);
nor U17793 (N_17793,N_16687,N_16805);
xnor U17794 (N_17794,N_16285,N_16482);
nor U17795 (N_17795,N_16633,N_16852);
nor U17796 (N_17796,N_16216,N_16657);
and U17797 (N_17797,N_16267,N_16286);
nand U17798 (N_17798,N_16441,N_16419);
or U17799 (N_17799,N_16364,N_16126);
nor U17800 (N_17800,N_16176,N_16726);
and U17801 (N_17801,N_16139,N_16211);
xor U17802 (N_17802,N_16413,N_16029);
xnor U17803 (N_17803,N_16788,N_16542);
nor U17804 (N_17804,N_16226,N_16513);
and U17805 (N_17805,N_16858,N_16399);
xnor U17806 (N_17806,N_16212,N_16124);
nand U17807 (N_17807,N_16389,N_16425);
nor U17808 (N_17808,N_16067,N_16209);
and U17809 (N_17809,N_16833,N_16738);
xnor U17810 (N_17810,N_16633,N_16794);
and U17811 (N_17811,N_16327,N_16204);
or U17812 (N_17812,N_16228,N_16394);
or U17813 (N_17813,N_16318,N_16742);
xor U17814 (N_17814,N_16834,N_16300);
nand U17815 (N_17815,N_16275,N_16485);
or U17816 (N_17816,N_16147,N_16589);
nand U17817 (N_17817,N_16041,N_16826);
nor U17818 (N_17818,N_16979,N_16988);
nand U17819 (N_17819,N_16772,N_16874);
or U17820 (N_17820,N_16434,N_16947);
nor U17821 (N_17821,N_16544,N_16496);
or U17822 (N_17822,N_16769,N_16585);
nand U17823 (N_17823,N_16554,N_16699);
nor U17824 (N_17824,N_16298,N_16123);
nor U17825 (N_17825,N_16846,N_16871);
and U17826 (N_17826,N_16943,N_16699);
and U17827 (N_17827,N_16071,N_16688);
nand U17828 (N_17828,N_16962,N_16557);
and U17829 (N_17829,N_16183,N_16629);
and U17830 (N_17830,N_16372,N_16711);
and U17831 (N_17831,N_16757,N_16417);
nand U17832 (N_17832,N_16677,N_16282);
nor U17833 (N_17833,N_16203,N_16320);
nor U17834 (N_17834,N_16795,N_16645);
nor U17835 (N_17835,N_16959,N_16328);
or U17836 (N_17836,N_16235,N_16270);
xnor U17837 (N_17837,N_16776,N_16791);
and U17838 (N_17838,N_16188,N_16136);
or U17839 (N_17839,N_16659,N_16119);
nand U17840 (N_17840,N_16052,N_16489);
nand U17841 (N_17841,N_16918,N_16427);
and U17842 (N_17842,N_16825,N_16166);
nand U17843 (N_17843,N_16687,N_16157);
nor U17844 (N_17844,N_16554,N_16557);
or U17845 (N_17845,N_16112,N_16590);
nor U17846 (N_17846,N_16728,N_16320);
xnor U17847 (N_17847,N_16457,N_16683);
nand U17848 (N_17848,N_16433,N_16839);
and U17849 (N_17849,N_16682,N_16350);
or U17850 (N_17850,N_16886,N_16005);
or U17851 (N_17851,N_16054,N_16504);
xnor U17852 (N_17852,N_16112,N_16207);
xnor U17853 (N_17853,N_16332,N_16406);
xor U17854 (N_17854,N_16207,N_16750);
nand U17855 (N_17855,N_16921,N_16784);
xnor U17856 (N_17856,N_16612,N_16750);
nand U17857 (N_17857,N_16055,N_16661);
xor U17858 (N_17858,N_16139,N_16793);
xor U17859 (N_17859,N_16081,N_16717);
and U17860 (N_17860,N_16777,N_16732);
or U17861 (N_17861,N_16598,N_16286);
or U17862 (N_17862,N_16275,N_16883);
or U17863 (N_17863,N_16151,N_16792);
nand U17864 (N_17864,N_16264,N_16148);
xor U17865 (N_17865,N_16553,N_16078);
xnor U17866 (N_17866,N_16898,N_16570);
nor U17867 (N_17867,N_16175,N_16252);
xnor U17868 (N_17868,N_16263,N_16349);
nor U17869 (N_17869,N_16023,N_16741);
nand U17870 (N_17870,N_16271,N_16672);
or U17871 (N_17871,N_16507,N_16084);
xor U17872 (N_17872,N_16001,N_16477);
or U17873 (N_17873,N_16895,N_16526);
nand U17874 (N_17874,N_16512,N_16476);
xnor U17875 (N_17875,N_16891,N_16437);
nand U17876 (N_17876,N_16973,N_16682);
nor U17877 (N_17877,N_16921,N_16611);
and U17878 (N_17878,N_16483,N_16441);
xor U17879 (N_17879,N_16706,N_16951);
nand U17880 (N_17880,N_16199,N_16621);
and U17881 (N_17881,N_16945,N_16813);
and U17882 (N_17882,N_16574,N_16274);
nand U17883 (N_17883,N_16533,N_16180);
nand U17884 (N_17884,N_16891,N_16706);
xor U17885 (N_17885,N_16529,N_16096);
xor U17886 (N_17886,N_16973,N_16252);
xor U17887 (N_17887,N_16097,N_16975);
nor U17888 (N_17888,N_16051,N_16392);
and U17889 (N_17889,N_16777,N_16699);
or U17890 (N_17890,N_16221,N_16386);
nor U17891 (N_17891,N_16436,N_16711);
or U17892 (N_17892,N_16506,N_16158);
or U17893 (N_17893,N_16056,N_16161);
nor U17894 (N_17894,N_16942,N_16943);
xnor U17895 (N_17895,N_16969,N_16286);
nor U17896 (N_17896,N_16304,N_16192);
nor U17897 (N_17897,N_16223,N_16199);
nor U17898 (N_17898,N_16790,N_16648);
nor U17899 (N_17899,N_16006,N_16979);
nor U17900 (N_17900,N_16957,N_16660);
xnor U17901 (N_17901,N_16723,N_16303);
and U17902 (N_17902,N_16539,N_16989);
nand U17903 (N_17903,N_16058,N_16012);
xnor U17904 (N_17904,N_16258,N_16212);
or U17905 (N_17905,N_16660,N_16789);
or U17906 (N_17906,N_16143,N_16829);
xnor U17907 (N_17907,N_16753,N_16377);
or U17908 (N_17908,N_16300,N_16233);
nor U17909 (N_17909,N_16568,N_16757);
nor U17910 (N_17910,N_16720,N_16866);
nand U17911 (N_17911,N_16329,N_16165);
xnor U17912 (N_17912,N_16620,N_16179);
xnor U17913 (N_17913,N_16792,N_16676);
xor U17914 (N_17914,N_16342,N_16334);
and U17915 (N_17915,N_16499,N_16835);
or U17916 (N_17916,N_16431,N_16848);
and U17917 (N_17917,N_16613,N_16831);
xnor U17918 (N_17918,N_16148,N_16492);
and U17919 (N_17919,N_16723,N_16504);
nand U17920 (N_17920,N_16381,N_16655);
nand U17921 (N_17921,N_16849,N_16238);
nor U17922 (N_17922,N_16932,N_16980);
nand U17923 (N_17923,N_16202,N_16058);
nand U17924 (N_17924,N_16184,N_16049);
nand U17925 (N_17925,N_16977,N_16905);
or U17926 (N_17926,N_16247,N_16989);
and U17927 (N_17927,N_16933,N_16784);
nand U17928 (N_17928,N_16119,N_16660);
nor U17929 (N_17929,N_16545,N_16863);
nor U17930 (N_17930,N_16086,N_16707);
or U17931 (N_17931,N_16556,N_16299);
nor U17932 (N_17932,N_16692,N_16148);
xnor U17933 (N_17933,N_16226,N_16301);
or U17934 (N_17934,N_16556,N_16725);
or U17935 (N_17935,N_16551,N_16847);
xnor U17936 (N_17936,N_16601,N_16924);
nand U17937 (N_17937,N_16685,N_16064);
nand U17938 (N_17938,N_16593,N_16768);
or U17939 (N_17939,N_16662,N_16199);
or U17940 (N_17940,N_16245,N_16955);
and U17941 (N_17941,N_16082,N_16134);
nand U17942 (N_17942,N_16598,N_16471);
nor U17943 (N_17943,N_16737,N_16991);
or U17944 (N_17944,N_16090,N_16031);
nand U17945 (N_17945,N_16107,N_16543);
nand U17946 (N_17946,N_16949,N_16049);
xnor U17947 (N_17947,N_16707,N_16533);
nand U17948 (N_17948,N_16897,N_16172);
nand U17949 (N_17949,N_16677,N_16504);
and U17950 (N_17950,N_16005,N_16444);
nand U17951 (N_17951,N_16226,N_16136);
xnor U17952 (N_17952,N_16490,N_16520);
xnor U17953 (N_17953,N_16250,N_16553);
nand U17954 (N_17954,N_16152,N_16244);
nand U17955 (N_17955,N_16666,N_16808);
xor U17956 (N_17956,N_16629,N_16476);
xor U17957 (N_17957,N_16474,N_16057);
and U17958 (N_17958,N_16351,N_16508);
or U17959 (N_17959,N_16726,N_16388);
nor U17960 (N_17960,N_16301,N_16070);
nand U17961 (N_17961,N_16485,N_16476);
and U17962 (N_17962,N_16250,N_16423);
nor U17963 (N_17963,N_16163,N_16912);
nor U17964 (N_17964,N_16033,N_16997);
nand U17965 (N_17965,N_16801,N_16746);
nand U17966 (N_17966,N_16805,N_16609);
xor U17967 (N_17967,N_16512,N_16704);
xnor U17968 (N_17968,N_16831,N_16936);
xor U17969 (N_17969,N_16599,N_16475);
and U17970 (N_17970,N_16446,N_16043);
and U17971 (N_17971,N_16570,N_16017);
nand U17972 (N_17972,N_16415,N_16880);
xnor U17973 (N_17973,N_16438,N_16214);
and U17974 (N_17974,N_16070,N_16300);
nor U17975 (N_17975,N_16321,N_16108);
nand U17976 (N_17976,N_16553,N_16891);
nor U17977 (N_17977,N_16390,N_16977);
nor U17978 (N_17978,N_16543,N_16444);
nor U17979 (N_17979,N_16184,N_16952);
nand U17980 (N_17980,N_16760,N_16085);
nand U17981 (N_17981,N_16943,N_16301);
and U17982 (N_17982,N_16451,N_16640);
nor U17983 (N_17983,N_16798,N_16655);
xnor U17984 (N_17984,N_16357,N_16368);
nor U17985 (N_17985,N_16955,N_16212);
nand U17986 (N_17986,N_16776,N_16294);
and U17987 (N_17987,N_16067,N_16360);
nor U17988 (N_17988,N_16639,N_16103);
or U17989 (N_17989,N_16397,N_16521);
nor U17990 (N_17990,N_16717,N_16300);
xnor U17991 (N_17991,N_16952,N_16783);
and U17992 (N_17992,N_16150,N_16429);
xor U17993 (N_17993,N_16777,N_16484);
nor U17994 (N_17994,N_16835,N_16515);
nor U17995 (N_17995,N_16001,N_16807);
nor U17996 (N_17996,N_16802,N_16050);
xnor U17997 (N_17997,N_16558,N_16967);
xnor U17998 (N_17998,N_16232,N_16695);
and U17999 (N_17999,N_16185,N_16494);
or U18000 (N_18000,N_17923,N_17579);
and U18001 (N_18001,N_17120,N_17224);
nand U18002 (N_18002,N_17740,N_17123);
or U18003 (N_18003,N_17532,N_17915);
and U18004 (N_18004,N_17194,N_17349);
and U18005 (N_18005,N_17616,N_17651);
xnor U18006 (N_18006,N_17515,N_17784);
xor U18007 (N_18007,N_17965,N_17030);
nand U18008 (N_18008,N_17434,N_17510);
nor U18009 (N_18009,N_17960,N_17011);
or U18010 (N_18010,N_17757,N_17792);
or U18011 (N_18011,N_17004,N_17537);
nand U18012 (N_18012,N_17936,N_17296);
nand U18013 (N_18013,N_17855,N_17441);
nor U18014 (N_18014,N_17043,N_17594);
nor U18015 (N_18015,N_17967,N_17481);
nor U18016 (N_18016,N_17014,N_17648);
nor U18017 (N_18017,N_17061,N_17478);
and U18018 (N_18018,N_17169,N_17225);
xnor U18019 (N_18019,N_17955,N_17804);
or U18020 (N_18020,N_17362,N_17139);
nor U18021 (N_18021,N_17674,N_17426);
and U18022 (N_18022,N_17914,N_17494);
and U18023 (N_18023,N_17642,N_17581);
or U18024 (N_18024,N_17228,N_17365);
or U18025 (N_18025,N_17237,N_17896);
nor U18026 (N_18026,N_17111,N_17096);
or U18027 (N_18027,N_17591,N_17078);
nor U18028 (N_18028,N_17844,N_17099);
and U18029 (N_18029,N_17003,N_17779);
and U18030 (N_18030,N_17466,N_17387);
or U18031 (N_18031,N_17356,N_17005);
and U18032 (N_18032,N_17793,N_17089);
xnor U18033 (N_18033,N_17649,N_17333);
and U18034 (N_18034,N_17791,N_17271);
and U18035 (N_18035,N_17673,N_17538);
xor U18036 (N_18036,N_17599,N_17427);
nand U18037 (N_18037,N_17605,N_17530);
or U18038 (N_18038,N_17145,N_17208);
and U18039 (N_18039,N_17385,N_17761);
xor U18040 (N_18040,N_17430,N_17545);
and U18041 (N_18041,N_17406,N_17637);
nor U18042 (N_18042,N_17920,N_17662);
nand U18043 (N_18043,N_17218,N_17968);
or U18044 (N_18044,N_17289,N_17108);
nand U18045 (N_18045,N_17308,N_17009);
or U18046 (N_18046,N_17910,N_17116);
or U18047 (N_18047,N_17253,N_17195);
and U18048 (N_18048,N_17879,N_17025);
nor U18049 (N_18049,N_17068,N_17925);
xor U18050 (N_18050,N_17128,N_17277);
nor U18051 (N_18051,N_17344,N_17200);
nor U18052 (N_18052,N_17322,N_17058);
xnor U18053 (N_18053,N_17389,N_17683);
nand U18054 (N_18054,N_17611,N_17557);
xnor U18055 (N_18055,N_17086,N_17475);
or U18056 (N_18056,N_17191,N_17807);
xnor U18057 (N_18057,N_17613,N_17379);
nand U18058 (N_18058,N_17205,N_17847);
nand U18059 (N_18059,N_17511,N_17580);
nand U18060 (N_18060,N_17718,N_17703);
nand U18061 (N_18061,N_17549,N_17760);
nand U18062 (N_18062,N_17653,N_17996);
xnor U18063 (N_18063,N_17340,N_17608);
and U18064 (N_18064,N_17629,N_17382);
and U18065 (N_18065,N_17449,N_17564);
nand U18066 (N_18066,N_17464,N_17363);
xnor U18067 (N_18067,N_17026,N_17242);
and U18068 (N_18068,N_17047,N_17937);
nor U18069 (N_18069,N_17492,N_17151);
or U18070 (N_18070,N_17882,N_17552);
nand U18071 (N_18071,N_17971,N_17425);
nor U18072 (N_18072,N_17768,N_17186);
nor U18073 (N_18073,N_17725,N_17754);
and U18074 (N_18074,N_17626,N_17493);
or U18075 (N_18075,N_17583,N_17358);
nor U18076 (N_18076,N_17023,N_17395);
or U18077 (N_18077,N_17508,N_17459);
or U18078 (N_18078,N_17403,N_17097);
nand U18079 (N_18079,N_17122,N_17721);
and U18080 (N_18080,N_17782,N_17229);
nand U18081 (N_18081,N_17498,N_17269);
and U18082 (N_18082,N_17317,N_17342);
or U18083 (N_18083,N_17364,N_17748);
or U18084 (N_18084,N_17243,N_17990);
or U18085 (N_18085,N_17963,N_17625);
nor U18086 (N_18086,N_17874,N_17627);
nor U18087 (N_18087,N_17331,N_17708);
and U18088 (N_18088,N_17540,N_17315);
or U18089 (N_18089,N_17534,N_17823);
nor U18090 (N_18090,N_17446,N_17590);
xnor U18091 (N_18091,N_17067,N_17873);
nor U18092 (N_18092,N_17696,N_17070);
or U18093 (N_18093,N_17911,N_17343);
and U18094 (N_18094,N_17057,N_17739);
nor U18095 (N_18095,N_17077,N_17885);
nor U18096 (N_18096,N_17150,N_17053);
nor U18097 (N_18097,N_17082,N_17719);
or U18098 (N_18098,N_17869,N_17084);
and U18099 (N_18099,N_17726,N_17856);
xor U18100 (N_18100,N_17659,N_17692);
nand U18101 (N_18101,N_17094,N_17109);
xor U18102 (N_18102,N_17350,N_17360);
xnor U18103 (N_18103,N_17119,N_17815);
xnor U18104 (N_18104,N_17368,N_17972);
and U18105 (N_18105,N_17558,N_17973);
nand U18106 (N_18106,N_17908,N_17482);
nand U18107 (N_18107,N_17222,N_17341);
nand U18108 (N_18108,N_17531,N_17215);
nand U18109 (N_18109,N_17671,N_17774);
nor U18110 (N_18110,N_17802,N_17861);
nor U18111 (N_18111,N_17687,N_17201);
and U18112 (N_18112,N_17268,N_17091);
xnor U18113 (N_18113,N_17130,N_17589);
or U18114 (N_18114,N_17049,N_17704);
xnor U18115 (N_18115,N_17985,N_17541);
nor U18116 (N_18116,N_17016,N_17623);
xnor U18117 (N_18117,N_17255,N_17007);
nor U18118 (N_18118,N_17100,N_17560);
nand U18119 (N_18119,N_17448,N_17926);
nand U18120 (N_18120,N_17307,N_17993);
or U18121 (N_18121,N_17773,N_17431);
nor U18122 (N_18122,N_17886,N_17713);
and U18123 (N_18123,N_17414,N_17104);
xor U18124 (N_18124,N_17880,N_17313);
or U18125 (N_18125,N_17180,N_17079);
xnor U18126 (N_18126,N_17989,N_17176);
nand U18127 (N_18127,N_17216,N_17311);
xnor U18128 (N_18128,N_17036,N_17747);
nand U18129 (N_18129,N_17080,N_17593);
nand U18130 (N_18130,N_17232,N_17376);
xnor U18131 (N_18131,N_17612,N_17592);
and U18132 (N_18132,N_17320,N_17859);
and U18133 (N_18133,N_17889,N_17716);
or U18134 (N_18134,N_17756,N_17428);
xnor U18135 (N_18135,N_17957,N_17845);
or U18136 (N_18136,N_17790,N_17931);
or U18137 (N_18137,N_17249,N_17283);
or U18138 (N_18138,N_17744,N_17789);
xnor U18139 (N_18139,N_17676,N_17470);
xor U18140 (N_18140,N_17285,N_17155);
nand U18141 (N_18141,N_17633,N_17121);
nand U18142 (N_18142,N_17477,N_17520);
nor U18143 (N_18143,N_17574,N_17468);
nand U18144 (N_18144,N_17240,N_17894);
and U18145 (N_18145,N_17338,N_17125);
xnor U18146 (N_18146,N_17234,N_17359);
and U18147 (N_18147,N_17083,N_17691);
nand U18148 (N_18148,N_17219,N_17614);
or U18149 (N_18149,N_17962,N_17286);
or U18150 (N_18150,N_17452,N_17055);
nand U18151 (N_18151,N_17330,N_17752);
xor U18152 (N_18152,N_17717,N_17033);
nor U18153 (N_18153,N_17185,N_17213);
and U18154 (N_18154,N_17413,N_17546);
nand U18155 (N_18155,N_17987,N_17136);
nor U18156 (N_18156,N_17354,N_17245);
or U18157 (N_18157,N_17361,N_17897);
xor U18158 (N_18158,N_17995,N_17597);
nand U18159 (N_18159,N_17293,N_17034);
xor U18160 (N_18160,N_17404,N_17827);
xnor U18161 (N_18161,N_17841,N_17550);
xnor U18162 (N_18162,N_17974,N_17012);
nand U18163 (N_18163,N_17019,N_17595);
or U18164 (N_18164,N_17071,N_17573);
and U18165 (N_18165,N_17472,N_17586);
nor U18166 (N_18166,N_17017,N_17453);
nor U18167 (N_18167,N_17497,N_17115);
nor U18168 (N_18168,N_17235,N_17536);
nand U18169 (N_18169,N_17876,N_17852);
nor U18170 (N_18170,N_17835,N_17667);
nor U18171 (N_18171,N_17027,N_17266);
and U18172 (N_18172,N_17298,N_17887);
nor U18173 (N_18173,N_17838,N_17165);
or U18174 (N_18174,N_17064,N_17276);
and U18175 (N_18175,N_17321,N_17037);
and U18176 (N_18176,N_17352,N_17621);
xor U18177 (N_18177,N_17101,N_17143);
nand U18178 (N_18178,N_17433,N_17471);
nor U18179 (N_18179,N_17603,N_17863);
and U18180 (N_18180,N_17217,N_17295);
nand U18181 (N_18181,N_17429,N_17110);
nand U18182 (N_18182,N_17578,N_17417);
nor U18183 (N_18183,N_17056,N_17450);
and U18184 (N_18184,N_17762,N_17959);
and U18185 (N_18185,N_17800,N_17373);
xor U18186 (N_18186,N_17198,N_17206);
nand U18187 (N_18187,N_17712,N_17465);
xnor U18188 (N_18188,N_17875,N_17436);
or U18189 (N_18189,N_17476,N_17418);
and U18190 (N_18190,N_17275,N_17551);
or U18191 (N_18191,N_17256,N_17178);
nand U18192 (N_18192,N_17502,N_17854);
and U18193 (N_18193,N_17484,N_17930);
xnor U18194 (N_18194,N_17107,N_17357);
or U18195 (N_18195,N_17173,N_17786);
or U18196 (N_18196,N_17265,N_17817);
and U18197 (N_18197,N_17644,N_17624);
nand U18198 (N_18198,N_17575,N_17862);
nor U18199 (N_18199,N_17327,N_17826);
nor U18200 (N_18200,N_17144,N_17187);
xnor U18201 (N_18201,N_17830,N_17542);
or U18202 (N_18202,N_17252,N_17678);
nand U18203 (N_18203,N_17775,N_17851);
and U18204 (N_18204,N_17939,N_17035);
and U18205 (N_18205,N_17867,N_17374);
nor U18206 (N_18206,N_17951,N_17733);
nor U18207 (N_18207,N_17730,N_17399);
or U18208 (N_18208,N_17260,N_17190);
nor U18209 (N_18209,N_17246,N_17044);
and U18210 (N_18210,N_17188,N_17263);
nand U18211 (N_18211,N_17183,N_17182);
or U18212 (N_18212,N_17505,N_17038);
and U18213 (N_18213,N_17239,N_17149);
xnor U18214 (N_18214,N_17961,N_17656);
or U18215 (N_18215,N_17309,N_17698);
and U18216 (N_18216,N_17416,N_17022);
xnor U18217 (N_18217,N_17102,N_17073);
and U18218 (N_18218,N_17457,N_17400);
nor U18219 (N_18219,N_17607,N_17525);
and U18220 (N_18220,N_17443,N_17864);
xnor U18221 (N_18221,N_17474,N_17158);
nand U18222 (N_18222,N_17447,N_17041);
or U18223 (N_18223,N_17600,N_17689);
xor U18224 (N_18224,N_17000,N_17688);
nand U18225 (N_18225,N_17290,N_17829);
and U18226 (N_18226,N_17170,N_17619);
xor U18227 (N_18227,N_17646,N_17634);
xor U18228 (N_18228,N_17986,N_17378);
or U18229 (N_18229,N_17813,N_17615);
nand U18230 (N_18230,N_17977,N_17189);
xor U18231 (N_18231,N_17456,N_17112);
or U18232 (N_18232,N_17334,N_17780);
xor U18233 (N_18233,N_17172,N_17715);
xnor U18234 (N_18234,N_17883,N_17919);
nor U18235 (N_18235,N_17566,N_17390);
nor U18236 (N_18236,N_17212,N_17556);
xnor U18237 (N_18237,N_17741,N_17682);
or U18238 (N_18238,N_17500,N_17280);
and U18239 (N_18239,N_17927,N_17893);
and U18240 (N_18240,N_17522,N_17632);
or U18241 (N_18241,N_17749,N_17154);
or U18242 (N_18242,N_17994,N_17148);
nor U18243 (N_18243,N_17628,N_17720);
or U18244 (N_18244,N_17010,N_17496);
xor U18245 (N_18245,N_17895,N_17103);
and U18246 (N_18246,N_17814,N_17164);
nor U18247 (N_18247,N_17846,N_17300);
xnor U18248 (N_18248,N_17337,N_17060);
xnor U18249 (N_18249,N_17024,N_17346);
xor U18250 (N_18250,N_17901,N_17942);
nor U18251 (N_18251,N_17833,N_17710);
nand U18252 (N_18252,N_17066,N_17236);
or U18253 (N_18253,N_17348,N_17964);
nand U18254 (N_18254,N_17527,N_17998);
nand U18255 (N_18255,N_17559,N_17788);
nand U18256 (N_18256,N_17891,N_17900);
or U18257 (N_18257,N_17287,N_17432);
xnor U18258 (N_18258,N_17906,N_17743);
xor U18259 (N_18259,N_17764,N_17031);
nand U18260 (N_18260,N_17162,N_17909);
nand U18261 (N_18261,N_17132,N_17902);
or U18262 (N_18262,N_17650,N_17709);
xnor U18263 (N_18263,N_17383,N_17604);
xor U18264 (N_18264,N_17226,N_17439);
nor U18265 (N_18265,N_17798,N_17495);
nor U18266 (N_18266,N_17196,N_17654);
nor U18267 (N_18267,N_17291,N_17938);
and U18268 (N_18268,N_17618,N_17455);
or U18269 (N_18269,N_17622,N_17199);
nor U18270 (N_18270,N_17167,N_17763);
or U18271 (N_18271,N_17655,N_17489);
nor U18272 (N_18272,N_17904,N_17858);
nand U18273 (N_18273,N_17402,N_17272);
nand U18274 (N_18274,N_17072,N_17680);
nor U18275 (N_18275,N_17577,N_17701);
nand U18276 (N_18276,N_17140,N_17587);
and U18277 (N_18277,N_17606,N_17585);
nor U18278 (N_18278,N_17588,N_17778);
and U18279 (N_18279,N_17127,N_17948);
xor U18280 (N_18280,N_17842,N_17811);
and U18281 (N_18281,N_17137,N_17694);
xnor U18282 (N_18282,N_17419,N_17048);
and U18283 (N_18283,N_17746,N_17421);
xnor U18284 (N_18284,N_17281,N_17569);
and U18285 (N_18285,N_17576,N_17799);
xor U18286 (N_18286,N_17705,N_17685);
nand U18287 (N_18287,N_17535,N_17943);
or U18288 (N_18288,N_17405,N_17202);
nor U18289 (N_18289,N_17670,N_17160);
nand U18290 (N_18290,N_17503,N_17991);
or U18291 (N_18291,N_17770,N_17772);
xnor U18292 (N_18292,N_17020,N_17166);
nand U18293 (N_18293,N_17001,N_17257);
or U18294 (N_18294,N_17918,N_17840);
and U18295 (N_18295,N_17513,N_17050);
xnor U18296 (N_18296,N_17881,N_17485);
nor U18297 (N_18297,N_17988,N_17345);
or U18298 (N_18298,N_17582,N_17984);
nand U18299 (N_18299,N_17658,N_17220);
xnor U18300 (N_18300,N_17401,N_17602);
and U18301 (N_18301,N_17254,N_17509);
and U18302 (N_18302,N_17735,N_17533);
nand U18303 (N_18303,N_17843,N_17490);
or U18304 (N_18304,N_17258,N_17098);
nand U18305 (N_18305,N_17193,N_17380);
or U18306 (N_18306,N_17516,N_17052);
or U18307 (N_18307,N_17803,N_17442);
or U18308 (N_18308,N_17244,N_17381);
or U18309 (N_18309,N_17714,N_17711);
or U18310 (N_18310,N_17640,N_17106);
and U18311 (N_18311,N_17983,N_17042);
nor U18312 (N_18312,N_17006,N_17386);
nand U18313 (N_18313,N_17051,N_17652);
nor U18314 (N_18314,N_17877,N_17999);
nand U18315 (N_18315,N_17437,N_17131);
xnor U18316 (N_18316,N_17323,N_17335);
xor U18317 (N_18317,N_17250,N_17529);
xor U18318 (N_18318,N_17736,N_17241);
nor U18319 (N_18319,N_17928,N_17002);
or U18320 (N_18320,N_17828,N_17737);
or U18321 (N_18321,N_17572,N_17848);
and U18322 (N_18322,N_17903,N_17227);
xnor U18323 (N_18323,N_17913,N_17370);
nand U18324 (N_18324,N_17458,N_17539);
xor U18325 (N_18325,N_17684,N_17562);
or U18326 (N_18326,N_17324,N_17328);
nand U18327 (N_18327,N_17554,N_17561);
nand U18328 (N_18328,N_17114,N_17018);
xnor U18329 (N_18329,N_17620,N_17221);
nor U18330 (N_18330,N_17636,N_17675);
nor U18331 (N_18331,N_17781,N_17074);
or U18332 (N_18332,N_17565,N_17679);
nand U18333 (N_18333,N_17506,N_17105);
and U18334 (N_18334,N_17932,N_17231);
nand U18335 (N_18335,N_17367,N_17392);
xnor U18336 (N_18336,N_17865,N_17722);
xor U18337 (N_18337,N_17917,N_17398);
nor U18338 (N_18338,N_17032,N_17273);
nand U18339 (N_18339,N_17980,N_17617);
and U18340 (N_18340,N_17785,N_17821);
nor U18341 (N_18341,N_17059,N_17934);
xor U18342 (N_18342,N_17075,N_17021);
nor U18343 (N_18343,N_17366,N_17161);
nand U18344 (N_18344,N_17204,N_17157);
and U18345 (N_18345,N_17301,N_17734);
and U18346 (N_18346,N_17944,N_17796);
or U18347 (N_18347,N_17953,N_17794);
nand U18348 (N_18348,N_17647,N_17767);
or U18349 (N_18349,N_17677,N_17635);
or U18350 (N_18350,N_17029,N_17898);
xor U18351 (N_18351,N_17299,N_17069);
xor U18352 (N_18352,N_17834,N_17469);
nand U18353 (N_18353,N_17142,N_17134);
nor U18354 (N_18354,N_17251,N_17480);
xor U18355 (N_18355,N_17753,N_17092);
nor U18356 (N_18356,N_17093,N_17818);
nor U18357 (N_18357,N_17415,N_17504);
nand U18358 (N_18358,N_17325,N_17755);
and U18359 (N_18359,N_17871,N_17921);
nor U18360 (N_18360,N_17878,N_17292);
xor U18361 (N_18361,N_17982,N_17270);
and U18362 (N_18362,N_17384,N_17601);
and U18363 (N_18363,N_17488,N_17553);
nand U18364 (N_18364,N_17372,N_17526);
nand U18365 (N_18365,N_17375,N_17949);
nor U18366 (N_18366,N_17393,N_17126);
nor U18367 (N_18367,N_17806,N_17090);
xor U18368 (N_18368,N_17259,N_17700);
xnor U18369 (N_18369,N_17888,N_17669);
or U18370 (N_18370,N_17284,N_17312);
or U18371 (N_18371,N_17046,N_17750);
xnor U18372 (N_18372,N_17661,N_17336);
or U18373 (N_18373,N_17423,N_17769);
nor U18374 (N_18374,N_17810,N_17702);
or U18375 (N_18375,N_17391,N_17302);
or U18376 (N_18376,N_17727,N_17641);
or U18377 (N_18377,N_17435,N_17638);
or U18378 (N_18378,N_17849,N_17831);
xnor U18379 (N_18379,N_17454,N_17732);
and U18380 (N_18380,N_17521,N_17945);
nand U18381 (N_18381,N_17795,N_17808);
nand U18382 (N_18382,N_17728,N_17141);
xnor U18383 (N_18383,N_17866,N_17184);
xnor U18384 (N_18384,N_17825,N_17451);
and U18385 (N_18385,N_17668,N_17933);
nand U18386 (N_18386,N_17440,N_17054);
nand U18387 (N_18387,N_17460,N_17486);
nor U18388 (N_18388,N_17979,N_17820);
or U18389 (N_18389,N_17230,N_17279);
or U18390 (N_18390,N_17868,N_17326);
nand U18391 (N_18391,N_17063,N_17639);
nor U18392 (N_18392,N_17935,N_17095);
nand U18393 (N_18393,N_17135,N_17210);
xnor U18394 (N_18394,N_17666,N_17339);
xnor U18395 (N_18395,N_17304,N_17518);
xor U18396 (N_18396,N_17822,N_17267);
nor U18397 (N_18397,N_17015,N_17444);
nor U18398 (N_18398,N_17407,N_17872);
nand U18399 (N_18399,N_17347,N_17197);
nand U18400 (N_18400,N_17233,N_17870);
and U18401 (N_18401,N_17355,N_17524);
nor U18402 (N_18402,N_17514,N_17660);
or U18403 (N_18403,N_17706,N_17129);
and U18404 (N_18404,N_17956,N_17610);
xor U18405 (N_18405,N_17351,N_17462);
or U18406 (N_18406,N_17420,N_17596);
xor U18407 (N_18407,N_17681,N_17801);
nor U18408 (N_18408,N_17969,N_17742);
or U18409 (N_18409,N_17805,N_17922);
nand U18410 (N_18410,N_17517,N_17118);
nor U18411 (N_18411,N_17318,N_17411);
nand U18412 (N_18412,N_17174,N_17146);
and U18413 (N_18413,N_17329,N_17065);
nand U18414 (N_18414,N_17013,N_17777);
or U18415 (N_18415,N_17223,N_17238);
nand U18416 (N_18416,N_17857,N_17479);
or U18417 (N_18417,N_17377,N_17288);
or U18418 (N_18418,N_17631,N_17528);
nor U18419 (N_18419,N_17759,N_17463);
xor U18420 (N_18420,N_17584,N_17975);
xnor U18421 (N_18421,N_17907,N_17499);
or U18422 (N_18422,N_17081,N_17211);
or U18423 (N_18423,N_17396,N_17853);
xor U18424 (N_18424,N_17693,N_17181);
or U18425 (N_18425,N_17179,N_17899);
nand U18426 (N_18426,N_17369,N_17690);
and U18427 (N_18427,N_17563,N_17954);
and U18428 (N_18428,N_17353,N_17422);
nand U18429 (N_18429,N_17997,N_17214);
or U18430 (N_18430,N_17424,N_17306);
nand U18431 (N_18431,N_17850,N_17837);
and U18432 (N_18432,N_17207,N_17787);
nor U18433 (N_18433,N_17316,N_17905);
nor U18434 (N_18434,N_17643,N_17766);
xnor U18435 (N_18435,N_17085,N_17297);
nand U18436 (N_18436,N_17570,N_17394);
and U18437 (N_18437,N_17745,N_17410);
nand U18438 (N_18438,N_17209,N_17812);
and U18439 (N_18439,N_17156,N_17751);
or U18440 (N_18440,N_17133,N_17797);
or U18441 (N_18441,N_17159,N_17916);
nand U18442 (N_18442,N_17177,N_17758);
nor U18443 (N_18443,N_17783,N_17731);
and U18444 (N_18444,N_17672,N_17890);
nor U18445 (N_18445,N_17028,N_17117);
nor U18446 (N_18446,N_17824,N_17548);
xor U18447 (N_18447,N_17487,N_17147);
nand U18448 (N_18448,N_17892,N_17203);
nand U18449 (N_18449,N_17664,N_17809);
xnor U18450 (N_18450,N_17388,N_17819);
xnor U18451 (N_18451,N_17473,N_17630);
xnor U18452 (N_18452,N_17408,N_17941);
nand U18453 (N_18453,N_17319,N_17138);
nor U18454 (N_18454,N_17153,N_17884);
or U18455 (N_18455,N_17294,N_17519);
or U18456 (N_18456,N_17568,N_17924);
and U18457 (N_18457,N_17567,N_17771);
or U18458 (N_18458,N_17729,N_17571);
xnor U18459 (N_18459,N_17461,N_17278);
or U18460 (N_18460,N_17305,N_17978);
or U18461 (N_18461,N_17501,N_17929);
or U18462 (N_18462,N_17832,N_17697);
and U18463 (N_18463,N_17952,N_17609);
or U18464 (N_18464,N_17836,N_17547);
nor U18465 (N_18465,N_17310,N_17738);
or U18466 (N_18466,N_17657,N_17839);
xor U18467 (N_18467,N_17332,N_17045);
nand U18468 (N_18468,N_17543,N_17544);
xor U18469 (N_18469,N_17303,N_17724);
and U18470 (N_18470,N_17152,N_17171);
nor U18471 (N_18471,N_17765,N_17371);
nor U18472 (N_18472,N_17412,N_17282);
and U18473 (N_18473,N_17695,N_17088);
xor U18474 (N_18474,N_17512,N_17946);
or U18475 (N_18475,N_17663,N_17248);
nand U18476 (N_18476,N_17113,N_17966);
xor U18477 (N_18477,N_17723,N_17950);
nor U18478 (N_18478,N_17438,N_17491);
or U18479 (N_18479,N_17686,N_17555);
nand U18480 (N_18480,N_17992,N_17981);
and U18481 (N_18481,N_17262,N_17645);
nor U18482 (N_18482,N_17483,N_17665);
xor U18483 (N_18483,N_17409,N_17940);
and U18484 (N_18484,N_17860,N_17816);
or U18485 (N_18485,N_17039,N_17314);
nor U18486 (N_18486,N_17445,N_17168);
xnor U18487 (N_18487,N_17523,N_17947);
or U18488 (N_18488,N_17707,N_17958);
xnor U18489 (N_18489,N_17776,N_17264);
xor U18490 (N_18490,N_17912,N_17076);
nor U18491 (N_18491,N_17040,N_17507);
xnor U18492 (N_18492,N_17970,N_17467);
nand U18493 (N_18493,N_17247,N_17976);
nand U18494 (N_18494,N_17175,N_17192);
or U18495 (N_18495,N_17397,N_17598);
nand U18496 (N_18496,N_17087,N_17008);
and U18497 (N_18497,N_17124,N_17261);
and U18498 (N_18498,N_17062,N_17699);
xor U18499 (N_18499,N_17163,N_17274);
and U18500 (N_18500,N_17482,N_17625);
xor U18501 (N_18501,N_17503,N_17484);
xor U18502 (N_18502,N_17634,N_17278);
or U18503 (N_18503,N_17547,N_17940);
nand U18504 (N_18504,N_17469,N_17248);
xnor U18505 (N_18505,N_17926,N_17886);
nand U18506 (N_18506,N_17563,N_17813);
nand U18507 (N_18507,N_17937,N_17346);
and U18508 (N_18508,N_17483,N_17802);
nand U18509 (N_18509,N_17530,N_17033);
nor U18510 (N_18510,N_17892,N_17871);
or U18511 (N_18511,N_17019,N_17671);
nor U18512 (N_18512,N_17599,N_17679);
nand U18513 (N_18513,N_17502,N_17811);
or U18514 (N_18514,N_17193,N_17489);
and U18515 (N_18515,N_17034,N_17695);
nand U18516 (N_18516,N_17810,N_17253);
and U18517 (N_18517,N_17726,N_17512);
xor U18518 (N_18518,N_17662,N_17202);
nand U18519 (N_18519,N_17333,N_17432);
or U18520 (N_18520,N_17409,N_17923);
nand U18521 (N_18521,N_17983,N_17027);
or U18522 (N_18522,N_17260,N_17181);
or U18523 (N_18523,N_17782,N_17208);
nand U18524 (N_18524,N_17634,N_17828);
nor U18525 (N_18525,N_17726,N_17900);
or U18526 (N_18526,N_17536,N_17049);
or U18527 (N_18527,N_17986,N_17692);
or U18528 (N_18528,N_17173,N_17848);
nor U18529 (N_18529,N_17300,N_17572);
nand U18530 (N_18530,N_17394,N_17277);
nor U18531 (N_18531,N_17485,N_17604);
xnor U18532 (N_18532,N_17587,N_17291);
nand U18533 (N_18533,N_17668,N_17148);
nand U18534 (N_18534,N_17651,N_17938);
nor U18535 (N_18535,N_17986,N_17971);
nor U18536 (N_18536,N_17881,N_17738);
and U18537 (N_18537,N_17595,N_17349);
nor U18538 (N_18538,N_17485,N_17600);
xnor U18539 (N_18539,N_17944,N_17212);
nor U18540 (N_18540,N_17515,N_17363);
and U18541 (N_18541,N_17427,N_17606);
and U18542 (N_18542,N_17381,N_17723);
nand U18543 (N_18543,N_17238,N_17111);
or U18544 (N_18544,N_17638,N_17199);
nand U18545 (N_18545,N_17231,N_17255);
nand U18546 (N_18546,N_17179,N_17729);
nand U18547 (N_18547,N_17033,N_17655);
nor U18548 (N_18548,N_17003,N_17776);
nand U18549 (N_18549,N_17635,N_17908);
xnor U18550 (N_18550,N_17495,N_17041);
xor U18551 (N_18551,N_17032,N_17751);
and U18552 (N_18552,N_17081,N_17050);
and U18553 (N_18553,N_17176,N_17876);
xnor U18554 (N_18554,N_17494,N_17168);
xor U18555 (N_18555,N_17551,N_17128);
and U18556 (N_18556,N_17416,N_17822);
xnor U18557 (N_18557,N_17353,N_17579);
and U18558 (N_18558,N_17031,N_17669);
nand U18559 (N_18559,N_17806,N_17468);
and U18560 (N_18560,N_17885,N_17949);
nor U18561 (N_18561,N_17872,N_17502);
nand U18562 (N_18562,N_17728,N_17972);
or U18563 (N_18563,N_17121,N_17672);
nand U18564 (N_18564,N_17718,N_17756);
or U18565 (N_18565,N_17606,N_17506);
xnor U18566 (N_18566,N_17434,N_17542);
nand U18567 (N_18567,N_17759,N_17241);
nand U18568 (N_18568,N_17030,N_17273);
nand U18569 (N_18569,N_17677,N_17533);
or U18570 (N_18570,N_17828,N_17534);
xnor U18571 (N_18571,N_17450,N_17628);
or U18572 (N_18572,N_17792,N_17094);
and U18573 (N_18573,N_17317,N_17013);
and U18574 (N_18574,N_17075,N_17138);
nor U18575 (N_18575,N_17392,N_17839);
nor U18576 (N_18576,N_17053,N_17691);
nand U18577 (N_18577,N_17072,N_17002);
and U18578 (N_18578,N_17666,N_17902);
nand U18579 (N_18579,N_17044,N_17487);
or U18580 (N_18580,N_17239,N_17640);
nor U18581 (N_18581,N_17052,N_17075);
nor U18582 (N_18582,N_17827,N_17783);
or U18583 (N_18583,N_17835,N_17666);
or U18584 (N_18584,N_17200,N_17675);
nor U18585 (N_18585,N_17372,N_17520);
and U18586 (N_18586,N_17334,N_17538);
nand U18587 (N_18587,N_17511,N_17178);
and U18588 (N_18588,N_17495,N_17212);
and U18589 (N_18589,N_17238,N_17251);
xor U18590 (N_18590,N_17089,N_17712);
xnor U18591 (N_18591,N_17096,N_17050);
xor U18592 (N_18592,N_17028,N_17119);
and U18593 (N_18593,N_17968,N_17001);
nand U18594 (N_18594,N_17973,N_17099);
and U18595 (N_18595,N_17162,N_17194);
nand U18596 (N_18596,N_17191,N_17599);
and U18597 (N_18597,N_17394,N_17296);
or U18598 (N_18598,N_17202,N_17856);
nand U18599 (N_18599,N_17260,N_17751);
nor U18600 (N_18600,N_17755,N_17868);
xor U18601 (N_18601,N_17785,N_17539);
nand U18602 (N_18602,N_17706,N_17598);
or U18603 (N_18603,N_17392,N_17818);
nor U18604 (N_18604,N_17158,N_17643);
or U18605 (N_18605,N_17022,N_17640);
nor U18606 (N_18606,N_17812,N_17666);
and U18607 (N_18607,N_17628,N_17907);
xnor U18608 (N_18608,N_17115,N_17795);
nand U18609 (N_18609,N_17426,N_17594);
nand U18610 (N_18610,N_17158,N_17672);
or U18611 (N_18611,N_17695,N_17037);
nand U18612 (N_18612,N_17187,N_17448);
nand U18613 (N_18613,N_17065,N_17047);
nand U18614 (N_18614,N_17662,N_17770);
or U18615 (N_18615,N_17605,N_17204);
xnor U18616 (N_18616,N_17357,N_17920);
xnor U18617 (N_18617,N_17807,N_17240);
nor U18618 (N_18618,N_17074,N_17338);
or U18619 (N_18619,N_17400,N_17997);
xor U18620 (N_18620,N_17282,N_17898);
and U18621 (N_18621,N_17303,N_17919);
and U18622 (N_18622,N_17575,N_17415);
or U18623 (N_18623,N_17013,N_17202);
xor U18624 (N_18624,N_17276,N_17731);
nor U18625 (N_18625,N_17239,N_17213);
or U18626 (N_18626,N_17256,N_17433);
nor U18627 (N_18627,N_17080,N_17992);
nand U18628 (N_18628,N_17895,N_17440);
nand U18629 (N_18629,N_17213,N_17119);
xor U18630 (N_18630,N_17015,N_17130);
and U18631 (N_18631,N_17744,N_17364);
and U18632 (N_18632,N_17798,N_17145);
and U18633 (N_18633,N_17984,N_17449);
nor U18634 (N_18634,N_17458,N_17255);
and U18635 (N_18635,N_17562,N_17447);
and U18636 (N_18636,N_17622,N_17296);
xor U18637 (N_18637,N_17731,N_17045);
or U18638 (N_18638,N_17805,N_17088);
or U18639 (N_18639,N_17760,N_17327);
nor U18640 (N_18640,N_17285,N_17385);
and U18641 (N_18641,N_17874,N_17653);
nand U18642 (N_18642,N_17472,N_17650);
nand U18643 (N_18643,N_17840,N_17545);
or U18644 (N_18644,N_17891,N_17550);
and U18645 (N_18645,N_17457,N_17480);
xnor U18646 (N_18646,N_17905,N_17286);
and U18647 (N_18647,N_17485,N_17260);
nand U18648 (N_18648,N_17933,N_17070);
and U18649 (N_18649,N_17318,N_17049);
and U18650 (N_18650,N_17873,N_17915);
and U18651 (N_18651,N_17946,N_17394);
or U18652 (N_18652,N_17899,N_17688);
or U18653 (N_18653,N_17821,N_17339);
or U18654 (N_18654,N_17660,N_17710);
and U18655 (N_18655,N_17248,N_17890);
xor U18656 (N_18656,N_17533,N_17725);
xnor U18657 (N_18657,N_17680,N_17452);
nor U18658 (N_18658,N_17969,N_17794);
nor U18659 (N_18659,N_17355,N_17096);
nand U18660 (N_18660,N_17733,N_17404);
nor U18661 (N_18661,N_17642,N_17410);
xor U18662 (N_18662,N_17988,N_17751);
nor U18663 (N_18663,N_17763,N_17115);
nand U18664 (N_18664,N_17604,N_17650);
or U18665 (N_18665,N_17546,N_17007);
xor U18666 (N_18666,N_17079,N_17892);
xor U18667 (N_18667,N_17174,N_17201);
nand U18668 (N_18668,N_17763,N_17635);
or U18669 (N_18669,N_17954,N_17889);
or U18670 (N_18670,N_17183,N_17038);
nand U18671 (N_18671,N_17655,N_17549);
nor U18672 (N_18672,N_17517,N_17349);
or U18673 (N_18673,N_17620,N_17489);
or U18674 (N_18674,N_17823,N_17194);
or U18675 (N_18675,N_17357,N_17002);
nor U18676 (N_18676,N_17015,N_17859);
xor U18677 (N_18677,N_17874,N_17105);
and U18678 (N_18678,N_17153,N_17080);
xnor U18679 (N_18679,N_17597,N_17138);
nor U18680 (N_18680,N_17256,N_17780);
or U18681 (N_18681,N_17001,N_17961);
xnor U18682 (N_18682,N_17744,N_17997);
nor U18683 (N_18683,N_17522,N_17110);
and U18684 (N_18684,N_17082,N_17231);
nor U18685 (N_18685,N_17823,N_17032);
nand U18686 (N_18686,N_17356,N_17333);
nor U18687 (N_18687,N_17116,N_17314);
nand U18688 (N_18688,N_17085,N_17025);
nand U18689 (N_18689,N_17253,N_17753);
and U18690 (N_18690,N_17056,N_17851);
and U18691 (N_18691,N_17844,N_17268);
nand U18692 (N_18692,N_17606,N_17647);
xnor U18693 (N_18693,N_17073,N_17330);
and U18694 (N_18694,N_17042,N_17548);
nand U18695 (N_18695,N_17368,N_17455);
nor U18696 (N_18696,N_17766,N_17601);
and U18697 (N_18697,N_17784,N_17634);
nand U18698 (N_18698,N_17546,N_17217);
nor U18699 (N_18699,N_17904,N_17859);
xor U18700 (N_18700,N_17758,N_17123);
and U18701 (N_18701,N_17092,N_17750);
and U18702 (N_18702,N_17714,N_17404);
or U18703 (N_18703,N_17814,N_17877);
and U18704 (N_18704,N_17219,N_17995);
nor U18705 (N_18705,N_17282,N_17409);
and U18706 (N_18706,N_17501,N_17407);
and U18707 (N_18707,N_17123,N_17780);
or U18708 (N_18708,N_17718,N_17014);
or U18709 (N_18709,N_17139,N_17273);
nor U18710 (N_18710,N_17575,N_17048);
or U18711 (N_18711,N_17867,N_17714);
and U18712 (N_18712,N_17446,N_17584);
and U18713 (N_18713,N_17346,N_17526);
and U18714 (N_18714,N_17291,N_17840);
nor U18715 (N_18715,N_17165,N_17989);
or U18716 (N_18716,N_17848,N_17522);
nand U18717 (N_18717,N_17606,N_17658);
xor U18718 (N_18718,N_17155,N_17334);
and U18719 (N_18719,N_17344,N_17490);
nor U18720 (N_18720,N_17877,N_17825);
or U18721 (N_18721,N_17369,N_17337);
nand U18722 (N_18722,N_17694,N_17251);
nor U18723 (N_18723,N_17193,N_17059);
nor U18724 (N_18724,N_17713,N_17342);
or U18725 (N_18725,N_17111,N_17159);
nor U18726 (N_18726,N_17576,N_17246);
and U18727 (N_18727,N_17873,N_17096);
or U18728 (N_18728,N_17408,N_17135);
xor U18729 (N_18729,N_17301,N_17680);
nor U18730 (N_18730,N_17097,N_17152);
nor U18731 (N_18731,N_17166,N_17205);
and U18732 (N_18732,N_17024,N_17793);
xor U18733 (N_18733,N_17690,N_17384);
nand U18734 (N_18734,N_17924,N_17127);
xor U18735 (N_18735,N_17979,N_17325);
nor U18736 (N_18736,N_17269,N_17403);
nor U18737 (N_18737,N_17768,N_17115);
nand U18738 (N_18738,N_17816,N_17786);
nand U18739 (N_18739,N_17918,N_17650);
nor U18740 (N_18740,N_17217,N_17247);
and U18741 (N_18741,N_17944,N_17684);
xnor U18742 (N_18742,N_17218,N_17571);
or U18743 (N_18743,N_17496,N_17488);
nor U18744 (N_18744,N_17977,N_17292);
nand U18745 (N_18745,N_17042,N_17473);
nor U18746 (N_18746,N_17123,N_17590);
xnor U18747 (N_18747,N_17258,N_17668);
and U18748 (N_18748,N_17147,N_17094);
nand U18749 (N_18749,N_17847,N_17263);
nor U18750 (N_18750,N_17192,N_17194);
xnor U18751 (N_18751,N_17653,N_17651);
xnor U18752 (N_18752,N_17359,N_17309);
or U18753 (N_18753,N_17815,N_17738);
nor U18754 (N_18754,N_17567,N_17625);
xnor U18755 (N_18755,N_17135,N_17087);
xor U18756 (N_18756,N_17008,N_17695);
or U18757 (N_18757,N_17658,N_17460);
nand U18758 (N_18758,N_17842,N_17829);
xnor U18759 (N_18759,N_17190,N_17168);
nand U18760 (N_18760,N_17248,N_17839);
xnor U18761 (N_18761,N_17506,N_17651);
nor U18762 (N_18762,N_17337,N_17205);
and U18763 (N_18763,N_17503,N_17407);
or U18764 (N_18764,N_17631,N_17582);
nand U18765 (N_18765,N_17159,N_17928);
or U18766 (N_18766,N_17989,N_17451);
xnor U18767 (N_18767,N_17465,N_17410);
and U18768 (N_18768,N_17041,N_17302);
nand U18769 (N_18769,N_17671,N_17178);
nor U18770 (N_18770,N_17874,N_17992);
nand U18771 (N_18771,N_17882,N_17586);
or U18772 (N_18772,N_17395,N_17096);
and U18773 (N_18773,N_17257,N_17593);
and U18774 (N_18774,N_17302,N_17347);
nor U18775 (N_18775,N_17994,N_17701);
nor U18776 (N_18776,N_17832,N_17213);
nand U18777 (N_18777,N_17571,N_17850);
nand U18778 (N_18778,N_17078,N_17021);
xor U18779 (N_18779,N_17045,N_17968);
and U18780 (N_18780,N_17208,N_17099);
nor U18781 (N_18781,N_17261,N_17622);
nand U18782 (N_18782,N_17201,N_17607);
xnor U18783 (N_18783,N_17174,N_17735);
nor U18784 (N_18784,N_17432,N_17342);
or U18785 (N_18785,N_17440,N_17799);
or U18786 (N_18786,N_17965,N_17199);
nand U18787 (N_18787,N_17976,N_17724);
and U18788 (N_18788,N_17928,N_17040);
xor U18789 (N_18789,N_17007,N_17455);
and U18790 (N_18790,N_17220,N_17523);
xor U18791 (N_18791,N_17823,N_17605);
and U18792 (N_18792,N_17609,N_17936);
nor U18793 (N_18793,N_17576,N_17577);
xor U18794 (N_18794,N_17385,N_17848);
xor U18795 (N_18795,N_17808,N_17287);
nor U18796 (N_18796,N_17126,N_17553);
xor U18797 (N_18797,N_17079,N_17846);
nand U18798 (N_18798,N_17160,N_17526);
nand U18799 (N_18799,N_17953,N_17992);
xnor U18800 (N_18800,N_17422,N_17432);
xnor U18801 (N_18801,N_17450,N_17349);
xor U18802 (N_18802,N_17647,N_17339);
or U18803 (N_18803,N_17009,N_17685);
or U18804 (N_18804,N_17080,N_17285);
xnor U18805 (N_18805,N_17187,N_17269);
nor U18806 (N_18806,N_17195,N_17327);
or U18807 (N_18807,N_17097,N_17525);
xnor U18808 (N_18808,N_17078,N_17939);
nor U18809 (N_18809,N_17523,N_17790);
and U18810 (N_18810,N_17721,N_17623);
xnor U18811 (N_18811,N_17812,N_17054);
nor U18812 (N_18812,N_17647,N_17981);
nand U18813 (N_18813,N_17243,N_17389);
and U18814 (N_18814,N_17197,N_17427);
or U18815 (N_18815,N_17829,N_17225);
xnor U18816 (N_18816,N_17370,N_17290);
or U18817 (N_18817,N_17175,N_17622);
nor U18818 (N_18818,N_17709,N_17624);
or U18819 (N_18819,N_17413,N_17342);
and U18820 (N_18820,N_17262,N_17560);
or U18821 (N_18821,N_17713,N_17480);
xnor U18822 (N_18822,N_17750,N_17542);
xnor U18823 (N_18823,N_17424,N_17574);
xor U18824 (N_18824,N_17642,N_17341);
xnor U18825 (N_18825,N_17072,N_17177);
and U18826 (N_18826,N_17834,N_17653);
or U18827 (N_18827,N_17957,N_17774);
xnor U18828 (N_18828,N_17586,N_17244);
nand U18829 (N_18829,N_17779,N_17957);
xor U18830 (N_18830,N_17085,N_17750);
nand U18831 (N_18831,N_17016,N_17580);
nor U18832 (N_18832,N_17132,N_17740);
nand U18833 (N_18833,N_17287,N_17595);
nand U18834 (N_18834,N_17158,N_17784);
and U18835 (N_18835,N_17466,N_17896);
or U18836 (N_18836,N_17489,N_17384);
nor U18837 (N_18837,N_17634,N_17279);
xor U18838 (N_18838,N_17252,N_17339);
or U18839 (N_18839,N_17995,N_17551);
nor U18840 (N_18840,N_17875,N_17059);
nand U18841 (N_18841,N_17249,N_17939);
or U18842 (N_18842,N_17643,N_17392);
nand U18843 (N_18843,N_17278,N_17918);
nand U18844 (N_18844,N_17235,N_17099);
nor U18845 (N_18845,N_17636,N_17442);
nand U18846 (N_18846,N_17962,N_17789);
or U18847 (N_18847,N_17732,N_17980);
and U18848 (N_18848,N_17343,N_17807);
xor U18849 (N_18849,N_17605,N_17968);
or U18850 (N_18850,N_17003,N_17836);
nor U18851 (N_18851,N_17422,N_17652);
nand U18852 (N_18852,N_17344,N_17161);
nor U18853 (N_18853,N_17185,N_17962);
nor U18854 (N_18854,N_17393,N_17528);
xor U18855 (N_18855,N_17535,N_17945);
nand U18856 (N_18856,N_17604,N_17042);
nand U18857 (N_18857,N_17441,N_17305);
and U18858 (N_18858,N_17381,N_17508);
or U18859 (N_18859,N_17080,N_17820);
and U18860 (N_18860,N_17750,N_17489);
or U18861 (N_18861,N_17788,N_17636);
or U18862 (N_18862,N_17915,N_17068);
and U18863 (N_18863,N_17808,N_17425);
or U18864 (N_18864,N_17558,N_17351);
or U18865 (N_18865,N_17732,N_17104);
nand U18866 (N_18866,N_17659,N_17490);
nor U18867 (N_18867,N_17002,N_17554);
xor U18868 (N_18868,N_17017,N_17807);
nor U18869 (N_18869,N_17961,N_17297);
nor U18870 (N_18870,N_17380,N_17815);
nor U18871 (N_18871,N_17152,N_17235);
nand U18872 (N_18872,N_17400,N_17275);
or U18873 (N_18873,N_17798,N_17118);
xor U18874 (N_18874,N_17251,N_17164);
or U18875 (N_18875,N_17086,N_17714);
xor U18876 (N_18876,N_17518,N_17452);
nor U18877 (N_18877,N_17623,N_17944);
xnor U18878 (N_18878,N_17897,N_17265);
or U18879 (N_18879,N_17493,N_17633);
and U18880 (N_18880,N_17865,N_17471);
and U18881 (N_18881,N_17341,N_17078);
and U18882 (N_18882,N_17924,N_17227);
xnor U18883 (N_18883,N_17668,N_17935);
nor U18884 (N_18884,N_17836,N_17168);
and U18885 (N_18885,N_17659,N_17298);
nand U18886 (N_18886,N_17380,N_17381);
or U18887 (N_18887,N_17092,N_17874);
xnor U18888 (N_18888,N_17105,N_17412);
xor U18889 (N_18889,N_17808,N_17939);
or U18890 (N_18890,N_17996,N_17498);
xor U18891 (N_18891,N_17875,N_17778);
or U18892 (N_18892,N_17062,N_17204);
nand U18893 (N_18893,N_17818,N_17146);
xnor U18894 (N_18894,N_17359,N_17555);
xor U18895 (N_18895,N_17515,N_17200);
and U18896 (N_18896,N_17492,N_17825);
and U18897 (N_18897,N_17166,N_17411);
nand U18898 (N_18898,N_17782,N_17369);
xor U18899 (N_18899,N_17931,N_17632);
nor U18900 (N_18900,N_17307,N_17804);
nor U18901 (N_18901,N_17476,N_17364);
nand U18902 (N_18902,N_17389,N_17309);
or U18903 (N_18903,N_17558,N_17836);
nor U18904 (N_18904,N_17424,N_17983);
nand U18905 (N_18905,N_17380,N_17450);
nand U18906 (N_18906,N_17305,N_17404);
and U18907 (N_18907,N_17667,N_17525);
and U18908 (N_18908,N_17968,N_17039);
or U18909 (N_18909,N_17509,N_17290);
or U18910 (N_18910,N_17425,N_17833);
or U18911 (N_18911,N_17919,N_17097);
and U18912 (N_18912,N_17290,N_17532);
nand U18913 (N_18913,N_17553,N_17690);
nand U18914 (N_18914,N_17455,N_17298);
xnor U18915 (N_18915,N_17140,N_17005);
nand U18916 (N_18916,N_17612,N_17457);
nor U18917 (N_18917,N_17282,N_17582);
or U18918 (N_18918,N_17154,N_17458);
xnor U18919 (N_18919,N_17393,N_17098);
nor U18920 (N_18920,N_17837,N_17384);
and U18921 (N_18921,N_17190,N_17030);
nand U18922 (N_18922,N_17887,N_17878);
and U18923 (N_18923,N_17645,N_17183);
and U18924 (N_18924,N_17942,N_17333);
or U18925 (N_18925,N_17065,N_17371);
nand U18926 (N_18926,N_17672,N_17746);
xnor U18927 (N_18927,N_17938,N_17181);
nand U18928 (N_18928,N_17979,N_17592);
nand U18929 (N_18929,N_17611,N_17757);
xnor U18930 (N_18930,N_17783,N_17238);
or U18931 (N_18931,N_17374,N_17837);
xor U18932 (N_18932,N_17457,N_17898);
nand U18933 (N_18933,N_17772,N_17464);
nor U18934 (N_18934,N_17836,N_17152);
xnor U18935 (N_18935,N_17412,N_17948);
and U18936 (N_18936,N_17057,N_17734);
or U18937 (N_18937,N_17340,N_17786);
nand U18938 (N_18938,N_17503,N_17801);
nand U18939 (N_18939,N_17627,N_17026);
nand U18940 (N_18940,N_17470,N_17079);
nor U18941 (N_18941,N_17340,N_17118);
nor U18942 (N_18942,N_17082,N_17767);
or U18943 (N_18943,N_17927,N_17186);
and U18944 (N_18944,N_17339,N_17396);
nor U18945 (N_18945,N_17459,N_17341);
or U18946 (N_18946,N_17894,N_17142);
and U18947 (N_18947,N_17358,N_17124);
xor U18948 (N_18948,N_17924,N_17652);
nand U18949 (N_18949,N_17204,N_17673);
nand U18950 (N_18950,N_17355,N_17287);
nand U18951 (N_18951,N_17891,N_17578);
or U18952 (N_18952,N_17705,N_17815);
or U18953 (N_18953,N_17581,N_17232);
and U18954 (N_18954,N_17764,N_17854);
and U18955 (N_18955,N_17747,N_17073);
nand U18956 (N_18956,N_17956,N_17047);
nand U18957 (N_18957,N_17837,N_17997);
xnor U18958 (N_18958,N_17056,N_17264);
or U18959 (N_18959,N_17792,N_17933);
or U18960 (N_18960,N_17654,N_17657);
nand U18961 (N_18961,N_17341,N_17811);
and U18962 (N_18962,N_17285,N_17421);
nand U18963 (N_18963,N_17092,N_17553);
or U18964 (N_18964,N_17301,N_17372);
xnor U18965 (N_18965,N_17643,N_17890);
or U18966 (N_18966,N_17565,N_17466);
or U18967 (N_18967,N_17956,N_17814);
and U18968 (N_18968,N_17292,N_17291);
and U18969 (N_18969,N_17703,N_17240);
xnor U18970 (N_18970,N_17124,N_17435);
xor U18971 (N_18971,N_17735,N_17064);
nand U18972 (N_18972,N_17762,N_17901);
xor U18973 (N_18973,N_17528,N_17521);
or U18974 (N_18974,N_17078,N_17457);
nand U18975 (N_18975,N_17618,N_17389);
nor U18976 (N_18976,N_17017,N_17758);
xnor U18977 (N_18977,N_17470,N_17113);
nand U18978 (N_18978,N_17565,N_17944);
xnor U18979 (N_18979,N_17500,N_17821);
and U18980 (N_18980,N_17048,N_17982);
xor U18981 (N_18981,N_17249,N_17164);
or U18982 (N_18982,N_17174,N_17383);
xor U18983 (N_18983,N_17451,N_17588);
nand U18984 (N_18984,N_17195,N_17913);
or U18985 (N_18985,N_17687,N_17022);
nand U18986 (N_18986,N_17871,N_17519);
and U18987 (N_18987,N_17426,N_17136);
xor U18988 (N_18988,N_17001,N_17356);
nand U18989 (N_18989,N_17362,N_17246);
nor U18990 (N_18990,N_17775,N_17178);
and U18991 (N_18991,N_17899,N_17593);
nand U18992 (N_18992,N_17922,N_17916);
nand U18993 (N_18993,N_17146,N_17589);
nor U18994 (N_18994,N_17263,N_17938);
and U18995 (N_18995,N_17884,N_17266);
and U18996 (N_18996,N_17484,N_17708);
xnor U18997 (N_18997,N_17714,N_17847);
xnor U18998 (N_18998,N_17614,N_17885);
or U18999 (N_18999,N_17520,N_17028);
or U19000 (N_19000,N_18577,N_18563);
and U19001 (N_19001,N_18900,N_18239);
or U19002 (N_19002,N_18150,N_18605);
nor U19003 (N_19003,N_18041,N_18879);
nand U19004 (N_19004,N_18917,N_18462);
nand U19005 (N_19005,N_18548,N_18007);
or U19006 (N_19006,N_18358,N_18293);
xor U19007 (N_19007,N_18641,N_18770);
nor U19008 (N_19008,N_18314,N_18649);
nand U19009 (N_19009,N_18196,N_18801);
nor U19010 (N_19010,N_18178,N_18846);
nand U19011 (N_19011,N_18613,N_18591);
nand U19012 (N_19012,N_18315,N_18416);
xnor U19013 (N_19013,N_18124,N_18505);
nand U19014 (N_19014,N_18513,N_18109);
xor U19015 (N_19015,N_18881,N_18869);
and U19016 (N_19016,N_18834,N_18222);
xnor U19017 (N_19017,N_18495,N_18086);
nor U19018 (N_19018,N_18257,N_18687);
nand U19019 (N_19019,N_18515,N_18108);
and U19020 (N_19020,N_18956,N_18854);
nand U19021 (N_19021,N_18389,N_18087);
nor U19022 (N_19022,N_18329,N_18633);
xor U19023 (N_19023,N_18324,N_18964);
or U19024 (N_19024,N_18866,N_18403);
nor U19025 (N_19025,N_18494,N_18247);
nand U19026 (N_19026,N_18394,N_18910);
or U19027 (N_19027,N_18374,N_18698);
and U19028 (N_19028,N_18837,N_18651);
nor U19029 (N_19029,N_18249,N_18119);
nand U19030 (N_19030,N_18382,N_18506);
xor U19031 (N_19031,N_18053,N_18221);
nor U19032 (N_19032,N_18711,N_18231);
nor U19033 (N_19033,N_18372,N_18901);
or U19034 (N_19034,N_18559,N_18212);
or U19035 (N_19035,N_18012,N_18820);
nand U19036 (N_19036,N_18427,N_18502);
nor U19037 (N_19037,N_18682,N_18552);
nand U19038 (N_19038,N_18530,N_18233);
xor U19039 (N_19039,N_18617,N_18159);
and U19040 (N_19040,N_18156,N_18670);
or U19041 (N_19041,N_18180,N_18570);
and U19042 (N_19042,N_18798,N_18772);
and U19043 (N_19043,N_18133,N_18242);
and U19044 (N_19044,N_18479,N_18839);
nand U19045 (N_19045,N_18767,N_18807);
and U19046 (N_19046,N_18415,N_18726);
and U19047 (N_19047,N_18323,N_18840);
and U19048 (N_19048,N_18256,N_18643);
nand U19049 (N_19049,N_18349,N_18569);
nor U19050 (N_19050,N_18013,N_18624);
nand U19051 (N_19051,N_18457,N_18622);
and U19052 (N_19052,N_18052,N_18824);
or U19053 (N_19053,N_18134,N_18896);
nor U19054 (N_19054,N_18568,N_18011);
nand U19055 (N_19055,N_18929,N_18113);
nand U19056 (N_19056,N_18948,N_18520);
and U19057 (N_19057,N_18606,N_18432);
xor U19058 (N_19058,N_18688,N_18655);
or U19059 (N_19059,N_18126,N_18939);
nor U19060 (N_19060,N_18952,N_18173);
xnor U19061 (N_19061,N_18276,N_18386);
and U19062 (N_19062,N_18344,N_18650);
or U19063 (N_19063,N_18867,N_18312);
nand U19064 (N_19064,N_18618,N_18240);
nor U19065 (N_19065,N_18456,N_18877);
nand U19066 (N_19066,N_18454,N_18678);
and U19067 (N_19067,N_18431,N_18665);
xor U19068 (N_19068,N_18756,N_18683);
nor U19069 (N_19069,N_18627,N_18561);
nand U19070 (N_19070,N_18850,N_18458);
nand U19071 (N_19071,N_18923,N_18201);
and U19072 (N_19072,N_18039,N_18499);
nand U19073 (N_19073,N_18700,N_18593);
nor U19074 (N_19074,N_18521,N_18773);
xor U19075 (N_19075,N_18294,N_18465);
and U19076 (N_19076,N_18355,N_18288);
or U19077 (N_19077,N_18712,N_18895);
nor U19078 (N_19078,N_18913,N_18400);
nand U19079 (N_19079,N_18657,N_18528);
and U19080 (N_19080,N_18849,N_18414);
nor U19081 (N_19081,N_18885,N_18009);
or U19082 (N_19082,N_18006,N_18601);
xnor U19083 (N_19083,N_18790,N_18610);
xnor U19084 (N_19084,N_18171,N_18341);
nor U19085 (N_19085,N_18958,N_18460);
or U19086 (N_19086,N_18793,N_18645);
and U19087 (N_19087,N_18275,N_18061);
and U19088 (N_19088,N_18940,N_18283);
and U19089 (N_19089,N_18120,N_18220);
or U19090 (N_19090,N_18567,N_18851);
nand U19091 (N_19091,N_18174,N_18626);
nand U19092 (N_19092,N_18042,N_18640);
xnor U19093 (N_19093,N_18704,N_18269);
and U19094 (N_19094,N_18304,N_18959);
nor U19095 (N_19095,N_18379,N_18997);
and U19096 (N_19096,N_18906,N_18821);
or U19097 (N_19097,N_18290,N_18144);
or U19098 (N_19098,N_18830,N_18365);
nor U19099 (N_19099,N_18153,N_18518);
nand U19100 (N_19100,N_18788,N_18535);
and U19101 (N_19101,N_18463,N_18122);
and U19102 (N_19102,N_18031,N_18017);
nor U19103 (N_19103,N_18320,N_18916);
or U19104 (N_19104,N_18966,N_18861);
xnor U19105 (N_19105,N_18614,N_18067);
xor U19106 (N_19106,N_18470,N_18504);
nand U19107 (N_19107,N_18097,N_18746);
nand U19108 (N_19108,N_18918,N_18182);
or U19109 (N_19109,N_18048,N_18533);
nor U19110 (N_19110,N_18181,N_18326);
nand U19111 (N_19111,N_18538,N_18080);
nor U19112 (N_19112,N_18782,N_18160);
or U19113 (N_19113,N_18443,N_18975);
nand U19114 (N_19114,N_18003,N_18090);
or U19115 (N_19115,N_18033,N_18914);
nor U19116 (N_19116,N_18537,N_18440);
nand U19117 (N_19117,N_18101,N_18663);
xor U19118 (N_19118,N_18436,N_18799);
and U19119 (N_19119,N_18378,N_18168);
nand U19120 (N_19120,N_18322,N_18066);
nand U19121 (N_19121,N_18628,N_18500);
or U19122 (N_19122,N_18638,N_18448);
xor U19123 (N_19123,N_18576,N_18217);
or U19124 (N_19124,N_18919,N_18232);
and U19125 (N_19125,N_18703,N_18352);
and U19126 (N_19126,N_18699,N_18833);
and U19127 (N_19127,N_18862,N_18282);
xnor U19128 (N_19128,N_18478,N_18921);
nand U19129 (N_19129,N_18564,N_18104);
xnor U19130 (N_19130,N_18350,N_18556);
and U19131 (N_19131,N_18371,N_18037);
nand U19132 (N_19132,N_18313,N_18864);
nand U19133 (N_19133,N_18803,N_18169);
nor U19134 (N_19134,N_18207,N_18077);
nand U19135 (N_19135,N_18199,N_18811);
nor U19136 (N_19136,N_18656,N_18238);
or U19137 (N_19137,N_18004,N_18795);
or U19138 (N_19138,N_18765,N_18370);
nor U19139 (N_19139,N_18707,N_18865);
nand U19140 (N_19140,N_18875,N_18301);
or U19141 (N_19141,N_18999,N_18486);
or U19142 (N_19142,N_18511,N_18105);
nand U19143 (N_19143,N_18493,N_18955);
nand U19144 (N_19144,N_18482,N_18620);
nand U19145 (N_19145,N_18646,N_18557);
and U19146 (N_19146,N_18008,N_18029);
or U19147 (N_19147,N_18059,N_18010);
nand U19148 (N_19148,N_18198,N_18095);
nand U19149 (N_19149,N_18058,N_18945);
xnor U19150 (N_19150,N_18551,N_18084);
nand U19151 (N_19151,N_18353,N_18904);
or U19152 (N_19152,N_18596,N_18298);
xor U19153 (N_19153,N_18366,N_18377);
or U19154 (N_19154,N_18447,N_18580);
nor U19155 (N_19155,N_18225,N_18068);
and U19156 (N_19156,N_18884,N_18550);
and U19157 (N_19157,N_18021,N_18244);
nor U19158 (N_19158,N_18155,N_18000);
nor U19159 (N_19159,N_18481,N_18994);
and U19160 (N_19160,N_18229,N_18719);
or U19161 (N_19161,N_18438,N_18536);
nor U19162 (N_19162,N_18045,N_18336);
nor U19163 (N_19163,N_18965,N_18780);
nand U19164 (N_19164,N_18855,N_18760);
nand U19165 (N_19165,N_18951,N_18297);
or U19166 (N_19166,N_18743,N_18594);
and U19167 (N_19167,N_18270,N_18998);
and U19168 (N_19168,N_18762,N_18903);
xor U19169 (N_19169,N_18843,N_18206);
nor U19170 (N_19170,N_18608,N_18075);
nor U19171 (N_19171,N_18211,N_18475);
xnor U19172 (N_19172,N_18453,N_18020);
or U19173 (N_19173,N_18744,N_18176);
nor U19174 (N_19174,N_18727,N_18979);
xnor U19175 (N_19175,N_18857,N_18736);
or U19176 (N_19176,N_18183,N_18510);
xnor U19177 (N_19177,N_18532,N_18946);
nand U19178 (N_19178,N_18674,N_18092);
and U19179 (N_19179,N_18410,N_18963);
and U19180 (N_19180,N_18652,N_18339);
nand U19181 (N_19181,N_18328,N_18469);
and U19182 (N_19182,N_18433,N_18615);
xnor U19183 (N_19183,N_18747,N_18026);
nand U19184 (N_19184,N_18632,N_18209);
nand U19185 (N_19185,N_18060,N_18118);
or U19186 (N_19186,N_18934,N_18194);
nand U19187 (N_19187,N_18716,N_18452);
or U19188 (N_19188,N_18348,N_18172);
or U19189 (N_19189,N_18188,N_18985);
nand U19190 (N_19190,N_18630,N_18274);
xnor U19191 (N_19191,N_18996,N_18303);
xnor U19192 (N_19192,N_18404,N_18942);
and U19193 (N_19193,N_18295,N_18709);
xor U19194 (N_19194,N_18123,N_18391);
nand U19195 (N_19195,N_18592,N_18741);
xor U19196 (N_19196,N_18990,N_18920);
xnor U19197 (N_19197,N_18325,N_18125);
nor U19198 (N_19198,N_18813,N_18316);
xnor U19199 (N_19199,N_18149,N_18891);
xnor U19200 (N_19200,N_18546,N_18897);
nor U19201 (N_19201,N_18035,N_18284);
or U19202 (N_19202,N_18056,N_18573);
or U19203 (N_19203,N_18733,N_18730);
nor U19204 (N_19204,N_18018,N_18305);
xnor U19205 (N_19205,N_18944,N_18356);
and U19206 (N_19206,N_18468,N_18572);
nor U19207 (N_19207,N_18337,N_18675);
xnor U19208 (N_19208,N_18319,N_18602);
and U19209 (N_19209,N_18291,N_18005);
or U19210 (N_19210,N_18783,N_18406);
and U19211 (N_19211,N_18445,N_18265);
and U19212 (N_19212,N_18278,N_18096);
nor U19213 (N_19213,N_18986,N_18749);
nand U19214 (N_19214,N_18729,N_18525);
or U19215 (N_19215,N_18697,N_18634);
or U19216 (N_19216,N_18272,N_18128);
xnor U19217 (N_19217,N_18995,N_18589);
xor U19218 (N_19218,N_18794,N_18132);
xor U19219 (N_19219,N_18519,N_18595);
or U19220 (N_19220,N_18425,N_18260);
or U19221 (N_19221,N_18387,N_18512);
and U19222 (N_19222,N_18681,N_18116);
nand U19223 (N_19223,N_18507,N_18930);
or U19224 (N_19224,N_18516,N_18876);
and U19225 (N_19225,N_18720,N_18937);
or U19226 (N_19226,N_18190,N_18088);
nand U19227 (N_19227,N_18040,N_18714);
nor U19228 (N_19228,N_18822,N_18886);
or U19229 (N_19229,N_18079,N_18642);
or U19230 (N_19230,N_18145,N_18899);
nand U19231 (N_19231,N_18543,N_18841);
nand U19232 (N_19232,N_18664,N_18385);
nand U19233 (N_19233,N_18488,N_18828);
or U19234 (N_19234,N_18922,N_18070);
nand U19235 (N_19235,N_18393,N_18091);
nand U19236 (N_19236,N_18069,N_18737);
or U19237 (N_19237,N_18676,N_18338);
nor U19238 (N_19238,N_18263,N_18024);
xor U19239 (N_19239,N_18083,N_18361);
xnor U19240 (N_19240,N_18781,N_18562);
nand U19241 (N_19241,N_18390,N_18115);
or U19242 (N_19242,N_18107,N_18566);
xor U19243 (N_19243,N_18311,N_18332);
nor U19244 (N_19244,N_18420,N_18223);
or U19245 (N_19245,N_18451,N_18342);
xnor U19246 (N_19246,N_18299,N_18832);
or U19247 (N_19247,N_18635,N_18871);
nor U19248 (N_19248,N_18476,N_18555);
or U19249 (N_19249,N_18582,N_18166);
nand U19250 (N_19250,N_18976,N_18960);
nand U19251 (N_19251,N_18870,N_18838);
xnor U19252 (N_19252,N_18364,N_18637);
xor U19253 (N_19253,N_18384,N_18292);
and U19254 (N_19254,N_18074,N_18597);
nand U19255 (N_19255,N_18926,N_18581);
or U19256 (N_19256,N_18522,N_18752);
nor U19257 (N_19257,N_18738,N_18763);
or U19258 (N_19258,N_18245,N_18185);
xor U19259 (N_19259,N_18883,N_18197);
and U19260 (N_19260,N_18915,N_18224);
nand U19261 (N_19261,N_18271,N_18474);
xnor U19262 (N_19262,N_18192,N_18836);
or U19263 (N_19263,N_18397,N_18137);
xnor U19264 (N_19264,N_18131,N_18205);
xnor U19265 (N_19265,N_18121,N_18140);
xnor U19266 (N_19266,N_18873,N_18887);
xnor U19267 (N_19267,N_18027,N_18732);
xnor U19268 (N_19268,N_18847,N_18019);
nand U19269 (N_19269,N_18127,N_18014);
xnor U19270 (N_19270,N_18280,N_18015);
xor U19271 (N_19271,N_18829,N_18503);
or U19272 (N_19272,N_18739,N_18671);
nand U19273 (N_19273,N_18164,N_18255);
nand U19274 (N_19274,N_18351,N_18742);
or U19275 (N_19275,N_18179,N_18446);
and U19276 (N_19276,N_18842,N_18193);
and U19277 (N_19277,N_18234,N_18947);
and U19278 (N_19278,N_18653,N_18565);
and U19279 (N_19279,N_18286,N_18191);
or U19280 (N_19280,N_18983,N_18508);
nand U19281 (N_19281,N_18327,N_18340);
and U19282 (N_19282,N_18187,N_18266);
and U19283 (N_19283,N_18785,N_18310);
nand U19284 (N_19284,N_18514,N_18970);
or U19285 (N_19285,N_18129,N_18208);
or U19286 (N_19286,N_18442,N_18542);
nand U19287 (N_19287,N_18177,N_18558);
nand U19288 (N_19288,N_18094,N_18151);
or U19289 (N_19289,N_18135,N_18428);
xor U19290 (N_19290,N_18062,N_18775);
xor U19291 (N_19291,N_18954,N_18424);
xor U19292 (N_19292,N_18165,N_18860);
or U19293 (N_19293,N_18778,N_18710);
and U19294 (N_19294,N_18689,N_18808);
or U19295 (N_19295,N_18189,N_18072);
nand U19296 (N_19296,N_18631,N_18523);
nor U19297 (N_19297,N_18680,N_18421);
xor U19298 (N_19298,N_18784,N_18235);
xnor U19299 (N_19299,N_18334,N_18932);
or U19300 (N_19300,N_18654,N_18611);
xnor U19301 (N_19301,N_18418,N_18335);
and U19302 (N_19302,N_18435,N_18531);
xor U19303 (N_19303,N_18574,N_18363);
xnor U19304 (N_19304,N_18529,N_18912);
and U19305 (N_19305,N_18089,N_18441);
or U19306 (N_19306,N_18735,N_18677);
nand U19307 (N_19307,N_18471,N_18667);
nor U19308 (N_19308,N_18175,N_18152);
nor U19309 (N_19309,N_18872,N_18057);
xnor U19310 (N_19310,N_18988,N_18085);
xnor U19311 (N_19311,N_18599,N_18241);
nor U19312 (N_19312,N_18243,N_18973);
xor U19313 (N_19313,N_18740,N_18962);
or U19314 (N_19314,N_18941,N_18268);
nor U19315 (N_19315,N_18713,N_18868);
xor U19316 (N_19316,N_18658,N_18810);
xor U19317 (N_19317,N_18544,N_18022);
xnor U19318 (N_19318,N_18554,N_18974);
nor U19319 (N_19319,N_18405,N_18309);
and U19320 (N_19320,N_18686,N_18787);
and U19321 (N_19321,N_18831,N_18981);
nand U19322 (N_19322,N_18484,N_18691);
nor U19323 (N_19323,N_18660,N_18413);
or U19324 (N_19324,N_18219,N_18526);
xor U19325 (N_19325,N_18585,N_18844);
xor U19326 (N_19326,N_18859,N_18882);
and U19327 (N_19327,N_18203,N_18411);
nor U19328 (N_19328,N_18236,N_18501);
nand U19329 (N_19329,N_18705,N_18874);
nor U19330 (N_19330,N_18202,N_18321);
nor U19331 (N_19331,N_18750,N_18819);
nor U19332 (N_19332,N_18464,N_18267);
nor U19333 (N_19333,N_18950,N_18647);
or U19334 (N_19334,N_18967,N_18002);
nand U19335 (N_19335,N_18430,N_18722);
or U19336 (N_19336,N_18258,N_18724);
nand U19337 (N_19337,N_18991,N_18215);
nand U19338 (N_19338,N_18496,N_18346);
or U19339 (N_19339,N_18971,N_18110);
and U19340 (N_19340,N_18845,N_18163);
xor U19341 (N_19341,N_18890,N_18993);
nor U19342 (N_19342,N_18330,N_18685);
nand U19343 (N_19343,N_18791,N_18343);
or U19344 (N_19344,N_18143,N_18911);
or U19345 (N_19345,N_18666,N_18226);
and U19346 (N_19346,N_18717,N_18081);
and U19347 (N_19347,N_18114,N_18745);
and U19348 (N_19348,N_18186,N_18804);
and U19349 (N_19349,N_18708,N_18786);
or U19350 (N_19350,N_18306,N_18806);
and U19351 (N_19351,N_18603,N_18401);
or U19352 (N_19352,N_18333,N_18761);
nand U19353 (N_19353,N_18961,N_18982);
and U19354 (N_19354,N_18373,N_18672);
nor U19355 (N_19355,N_18277,N_18139);
xnor U19356 (N_19356,N_18639,N_18036);
or U19357 (N_19357,N_18908,N_18909);
xnor U19358 (N_19358,N_18560,N_18034);
xnor U19359 (N_19359,N_18853,N_18972);
and U19360 (N_19360,N_18753,N_18461);
nand U19361 (N_19361,N_18751,N_18308);
xor U19362 (N_19362,N_18136,N_18905);
and U19363 (N_19363,N_18099,N_18583);
xor U19364 (N_19364,N_18823,N_18025);
nand U19365 (N_19365,N_18578,N_18376);
or U19366 (N_19366,N_18130,N_18422);
or U19367 (N_19367,N_18409,N_18898);
nand U19368 (N_19368,N_18644,N_18809);
nand U19369 (N_19369,N_18759,N_18927);
nor U19370 (N_19370,N_18345,N_18038);
nor U19371 (N_19371,N_18586,N_18388);
nand U19372 (N_19372,N_18587,N_18792);
nor U19373 (N_19373,N_18210,N_18281);
and U19374 (N_19374,N_18623,N_18609);
and U19375 (N_19375,N_18835,N_18547);
and U19376 (N_19376,N_18769,N_18093);
or U19377 (N_19377,N_18987,N_18046);
nor U19378 (N_19378,N_18398,N_18734);
or U19379 (N_19379,N_18073,N_18098);
nor U19380 (N_19380,N_18318,N_18112);
xnor U19381 (N_19381,N_18103,N_18213);
xnor U19382 (N_19382,N_18827,N_18158);
and U19383 (N_19383,N_18980,N_18357);
xnor U19384 (N_19384,N_18362,N_18147);
and U19385 (N_19385,N_18978,N_18148);
nand U19386 (N_19386,N_18774,N_18032);
nor U19387 (N_19387,N_18047,N_18584);
nor U19388 (N_19388,N_18489,N_18858);
xnor U19389 (N_19389,N_18287,N_18161);
nand U19390 (N_19390,N_18279,N_18779);
nand U19391 (N_19391,N_18977,N_18050);
or U19392 (N_19392,N_18162,N_18368);
xor U19393 (N_19393,N_18679,N_18396);
nand U19394 (N_19394,N_18417,N_18359);
nor U19395 (N_19395,N_18553,N_18619);
and U19396 (N_19396,N_18648,N_18467);
or U19397 (N_19397,N_18216,N_18659);
nand U19398 (N_19398,N_18549,N_18360);
nor U19399 (N_19399,N_18517,N_18579);
nand U19400 (N_19400,N_18204,N_18931);
nand U19401 (N_19401,N_18138,N_18625);
xnor U19402 (N_19402,N_18826,N_18285);
nor U19403 (N_19403,N_18814,N_18825);
xor U19404 (N_19404,N_18369,N_18616);
nor U19405 (N_19405,N_18170,N_18100);
nor U19406 (N_19406,N_18662,N_18629);
nand U19407 (N_19407,N_18117,N_18262);
and U19408 (N_19408,N_18264,N_18771);
or U19409 (N_19409,N_18071,N_18218);
and U19410 (N_19410,N_18273,N_18102);
and U19411 (N_19411,N_18802,N_18848);
nor U19412 (N_19412,N_18450,N_18925);
nand U19413 (N_19413,N_18111,N_18483);
nor U19414 (N_19414,N_18383,N_18852);
or U19415 (N_19415,N_18706,N_18141);
nor U19416 (N_19416,N_18892,N_18612);
xnor U19417 (N_19417,N_18049,N_18289);
or U19418 (N_19418,N_18228,N_18894);
nor U19419 (N_19419,N_18758,N_18856);
nor U19420 (N_19420,N_18943,N_18661);
and U19421 (N_19421,N_18195,N_18701);
nand U19422 (N_19422,N_18001,N_18527);
and U19423 (N_19423,N_18969,N_18146);
nand U19424 (N_19424,N_18902,N_18480);
nor U19425 (N_19425,N_18254,N_18347);
or U19426 (N_19426,N_18694,N_18076);
xor U19427 (N_19427,N_18055,N_18796);
nand U19428 (N_19428,N_18251,N_18466);
and U19429 (N_19429,N_18472,N_18167);
or U19430 (N_19430,N_18721,N_18936);
nand U19431 (N_19431,N_18434,N_18261);
or U19432 (N_19432,N_18491,N_18755);
xnor U19433 (N_19433,N_18296,N_18968);
nor U19434 (N_19434,N_18317,N_18246);
and U19435 (N_19435,N_18395,N_18636);
nand U19436 (N_19436,N_18230,N_18789);
or U19437 (N_19437,N_18805,N_18375);
and U19438 (N_19438,N_18907,N_18728);
or U19439 (N_19439,N_18816,N_18030);
nor U19440 (N_19440,N_18777,N_18399);
nand U19441 (N_19441,N_18725,N_18889);
or U19442 (N_19442,N_18429,N_18754);
or U19443 (N_19443,N_18723,N_18490);
nor U19444 (N_19444,N_18142,N_18065);
and U19445 (N_19445,N_18764,N_18957);
nor U19446 (N_19446,N_18668,N_18419);
and U19447 (N_19447,N_18992,N_18541);
xor U19448 (N_19448,N_18184,N_18757);
nor U19449 (N_19449,N_18540,N_18815);
nand U19450 (N_19450,N_18227,N_18082);
xor U19451 (N_19451,N_18695,N_18354);
and U19452 (N_19452,N_18307,N_18439);
nor U19453 (N_19453,N_18078,N_18455);
or U19454 (N_19454,N_18539,N_18051);
and U19455 (N_19455,N_18485,N_18253);
nand U19456 (N_19456,N_18043,N_18449);
and U19457 (N_19457,N_18367,N_18669);
nand U19458 (N_19458,N_18016,N_18380);
nand U19459 (N_19459,N_18953,N_18818);
and U19460 (N_19460,N_18800,N_18673);
or U19461 (N_19461,N_18766,N_18473);
nand U19462 (N_19462,N_18302,N_18598);
and U19463 (N_19463,N_18492,N_18402);
or U19464 (N_19464,N_18702,N_18237);
nor U19465 (N_19465,N_18259,N_18878);
nor U19466 (N_19466,N_18407,N_18381);
or U19467 (N_19467,N_18028,N_18600);
nor U19468 (N_19468,N_18621,N_18863);
nand U19469 (N_19469,N_18604,N_18938);
nor U19470 (N_19470,N_18888,N_18933);
or U19471 (N_19471,N_18392,N_18064);
or U19472 (N_19472,N_18748,N_18693);
nand U19473 (N_19473,N_18509,N_18524);
nand U19474 (N_19474,N_18252,N_18154);
or U19475 (N_19475,N_18590,N_18588);
or U19476 (N_19476,N_18444,N_18928);
nor U19477 (N_19477,N_18812,N_18718);
and U19478 (N_19478,N_18063,N_18248);
nand U19479 (N_19479,N_18817,N_18534);
and U19480 (N_19480,N_18331,N_18696);
and U19481 (N_19481,N_18044,N_18776);
and U19482 (N_19482,N_18459,N_18426);
and U19483 (N_19483,N_18487,N_18054);
nor U19484 (N_19484,N_18571,N_18731);
and U19485 (N_19485,N_18545,N_18797);
nor U19486 (N_19486,N_18989,N_18250);
nor U19487 (N_19487,N_18984,N_18437);
nor U19488 (N_19488,N_18497,N_18157);
nor U19489 (N_19489,N_18498,N_18924);
or U19490 (N_19490,N_18477,N_18935);
or U19491 (N_19491,N_18200,N_18949);
nor U19492 (N_19492,N_18214,N_18690);
or U19493 (N_19493,N_18023,N_18893);
xnor U19494 (N_19494,N_18412,N_18575);
or U19495 (N_19495,N_18300,N_18692);
nand U19496 (N_19496,N_18684,N_18423);
nand U19497 (N_19497,N_18408,N_18106);
nand U19498 (N_19498,N_18880,N_18715);
xor U19499 (N_19499,N_18607,N_18768);
or U19500 (N_19500,N_18570,N_18397);
nand U19501 (N_19501,N_18691,N_18405);
xor U19502 (N_19502,N_18880,N_18927);
xor U19503 (N_19503,N_18779,N_18292);
nor U19504 (N_19504,N_18726,N_18709);
xnor U19505 (N_19505,N_18724,N_18487);
xnor U19506 (N_19506,N_18580,N_18614);
nand U19507 (N_19507,N_18011,N_18537);
and U19508 (N_19508,N_18524,N_18414);
xor U19509 (N_19509,N_18050,N_18513);
and U19510 (N_19510,N_18333,N_18862);
nand U19511 (N_19511,N_18969,N_18669);
and U19512 (N_19512,N_18013,N_18833);
nand U19513 (N_19513,N_18438,N_18019);
xor U19514 (N_19514,N_18234,N_18782);
xor U19515 (N_19515,N_18505,N_18070);
nand U19516 (N_19516,N_18990,N_18998);
and U19517 (N_19517,N_18165,N_18305);
xnor U19518 (N_19518,N_18180,N_18589);
xnor U19519 (N_19519,N_18048,N_18254);
and U19520 (N_19520,N_18443,N_18598);
nand U19521 (N_19521,N_18535,N_18110);
nand U19522 (N_19522,N_18397,N_18564);
or U19523 (N_19523,N_18718,N_18093);
and U19524 (N_19524,N_18131,N_18632);
nand U19525 (N_19525,N_18279,N_18987);
xnor U19526 (N_19526,N_18150,N_18537);
and U19527 (N_19527,N_18875,N_18391);
or U19528 (N_19528,N_18974,N_18526);
or U19529 (N_19529,N_18252,N_18828);
nand U19530 (N_19530,N_18524,N_18018);
and U19531 (N_19531,N_18029,N_18700);
xnor U19532 (N_19532,N_18286,N_18847);
nor U19533 (N_19533,N_18865,N_18772);
and U19534 (N_19534,N_18191,N_18644);
and U19535 (N_19535,N_18813,N_18851);
nor U19536 (N_19536,N_18688,N_18686);
nor U19537 (N_19537,N_18126,N_18058);
nor U19538 (N_19538,N_18313,N_18591);
nor U19539 (N_19539,N_18084,N_18033);
xnor U19540 (N_19540,N_18577,N_18179);
nor U19541 (N_19541,N_18369,N_18308);
or U19542 (N_19542,N_18257,N_18376);
nor U19543 (N_19543,N_18559,N_18950);
nor U19544 (N_19544,N_18192,N_18996);
or U19545 (N_19545,N_18341,N_18090);
nand U19546 (N_19546,N_18612,N_18848);
or U19547 (N_19547,N_18528,N_18252);
and U19548 (N_19548,N_18746,N_18838);
or U19549 (N_19549,N_18301,N_18569);
nor U19550 (N_19550,N_18753,N_18017);
or U19551 (N_19551,N_18058,N_18642);
nor U19552 (N_19552,N_18739,N_18685);
and U19553 (N_19553,N_18683,N_18875);
and U19554 (N_19554,N_18991,N_18483);
xnor U19555 (N_19555,N_18081,N_18847);
xnor U19556 (N_19556,N_18532,N_18081);
or U19557 (N_19557,N_18265,N_18471);
and U19558 (N_19558,N_18960,N_18407);
or U19559 (N_19559,N_18344,N_18616);
nand U19560 (N_19560,N_18051,N_18669);
nor U19561 (N_19561,N_18590,N_18657);
or U19562 (N_19562,N_18144,N_18616);
nand U19563 (N_19563,N_18460,N_18468);
nand U19564 (N_19564,N_18154,N_18241);
nor U19565 (N_19565,N_18450,N_18273);
nor U19566 (N_19566,N_18896,N_18030);
or U19567 (N_19567,N_18289,N_18499);
and U19568 (N_19568,N_18073,N_18488);
or U19569 (N_19569,N_18429,N_18466);
nor U19570 (N_19570,N_18985,N_18911);
or U19571 (N_19571,N_18015,N_18873);
nor U19572 (N_19572,N_18156,N_18560);
xor U19573 (N_19573,N_18785,N_18745);
or U19574 (N_19574,N_18928,N_18786);
xor U19575 (N_19575,N_18851,N_18049);
nand U19576 (N_19576,N_18340,N_18256);
or U19577 (N_19577,N_18800,N_18385);
nand U19578 (N_19578,N_18613,N_18010);
nor U19579 (N_19579,N_18029,N_18638);
nand U19580 (N_19580,N_18497,N_18629);
and U19581 (N_19581,N_18610,N_18717);
and U19582 (N_19582,N_18361,N_18218);
nor U19583 (N_19583,N_18408,N_18630);
and U19584 (N_19584,N_18858,N_18290);
nand U19585 (N_19585,N_18369,N_18584);
nand U19586 (N_19586,N_18046,N_18552);
nand U19587 (N_19587,N_18063,N_18503);
and U19588 (N_19588,N_18502,N_18078);
or U19589 (N_19589,N_18182,N_18192);
nand U19590 (N_19590,N_18150,N_18789);
or U19591 (N_19591,N_18470,N_18076);
xnor U19592 (N_19592,N_18041,N_18272);
or U19593 (N_19593,N_18429,N_18820);
or U19594 (N_19594,N_18507,N_18227);
nand U19595 (N_19595,N_18788,N_18689);
and U19596 (N_19596,N_18370,N_18715);
or U19597 (N_19597,N_18050,N_18539);
or U19598 (N_19598,N_18537,N_18516);
nand U19599 (N_19599,N_18634,N_18748);
nand U19600 (N_19600,N_18368,N_18239);
or U19601 (N_19601,N_18834,N_18479);
nor U19602 (N_19602,N_18252,N_18474);
nor U19603 (N_19603,N_18527,N_18790);
and U19604 (N_19604,N_18482,N_18377);
xnor U19605 (N_19605,N_18623,N_18963);
xor U19606 (N_19606,N_18814,N_18771);
and U19607 (N_19607,N_18622,N_18135);
and U19608 (N_19608,N_18402,N_18060);
nor U19609 (N_19609,N_18330,N_18577);
nor U19610 (N_19610,N_18783,N_18645);
xnor U19611 (N_19611,N_18970,N_18897);
or U19612 (N_19612,N_18407,N_18091);
xnor U19613 (N_19613,N_18137,N_18813);
nor U19614 (N_19614,N_18941,N_18465);
nand U19615 (N_19615,N_18627,N_18819);
and U19616 (N_19616,N_18951,N_18716);
nand U19617 (N_19617,N_18533,N_18178);
and U19618 (N_19618,N_18369,N_18328);
xor U19619 (N_19619,N_18020,N_18602);
nand U19620 (N_19620,N_18046,N_18865);
nand U19621 (N_19621,N_18877,N_18938);
nand U19622 (N_19622,N_18389,N_18688);
and U19623 (N_19623,N_18637,N_18123);
nand U19624 (N_19624,N_18722,N_18759);
and U19625 (N_19625,N_18352,N_18142);
or U19626 (N_19626,N_18731,N_18451);
or U19627 (N_19627,N_18266,N_18356);
nor U19628 (N_19628,N_18872,N_18935);
xnor U19629 (N_19629,N_18333,N_18758);
nor U19630 (N_19630,N_18191,N_18214);
and U19631 (N_19631,N_18451,N_18624);
nor U19632 (N_19632,N_18847,N_18900);
nand U19633 (N_19633,N_18089,N_18533);
nand U19634 (N_19634,N_18414,N_18880);
nor U19635 (N_19635,N_18036,N_18017);
xnor U19636 (N_19636,N_18148,N_18572);
nand U19637 (N_19637,N_18986,N_18109);
nand U19638 (N_19638,N_18453,N_18908);
xnor U19639 (N_19639,N_18180,N_18101);
and U19640 (N_19640,N_18620,N_18686);
nand U19641 (N_19641,N_18093,N_18603);
and U19642 (N_19642,N_18584,N_18571);
or U19643 (N_19643,N_18216,N_18186);
or U19644 (N_19644,N_18365,N_18920);
and U19645 (N_19645,N_18466,N_18615);
xnor U19646 (N_19646,N_18124,N_18015);
nand U19647 (N_19647,N_18710,N_18335);
nand U19648 (N_19648,N_18838,N_18398);
xor U19649 (N_19649,N_18602,N_18367);
xor U19650 (N_19650,N_18775,N_18049);
nor U19651 (N_19651,N_18759,N_18702);
xor U19652 (N_19652,N_18935,N_18775);
and U19653 (N_19653,N_18757,N_18876);
and U19654 (N_19654,N_18993,N_18305);
and U19655 (N_19655,N_18161,N_18744);
or U19656 (N_19656,N_18523,N_18230);
and U19657 (N_19657,N_18621,N_18849);
and U19658 (N_19658,N_18491,N_18886);
and U19659 (N_19659,N_18470,N_18523);
or U19660 (N_19660,N_18897,N_18162);
nor U19661 (N_19661,N_18351,N_18966);
nor U19662 (N_19662,N_18017,N_18084);
xor U19663 (N_19663,N_18903,N_18491);
or U19664 (N_19664,N_18305,N_18493);
nor U19665 (N_19665,N_18954,N_18102);
or U19666 (N_19666,N_18434,N_18457);
nand U19667 (N_19667,N_18924,N_18906);
or U19668 (N_19668,N_18591,N_18893);
nor U19669 (N_19669,N_18638,N_18632);
nor U19670 (N_19670,N_18904,N_18960);
or U19671 (N_19671,N_18392,N_18119);
or U19672 (N_19672,N_18027,N_18687);
nor U19673 (N_19673,N_18428,N_18378);
nand U19674 (N_19674,N_18319,N_18696);
nand U19675 (N_19675,N_18967,N_18457);
and U19676 (N_19676,N_18061,N_18626);
nand U19677 (N_19677,N_18607,N_18788);
and U19678 (N_19678,N_18688,N_18230);
or U19679 (N_19679,N_18839,N_18378);
nand U19680 (N_19680,N_18089,N_18819);
xnor U19681 (N_19681,N_18604,N_18426);
or U19682 (N_19682,N_18559,N_18698);
or U19683 (N_19683,N_18528,N_18561);
or U19684 (N_19684,N_18734,N_18963);
or U19685 (N_19685,N_18951,N_18633);
or U19686 (N_19686,N_18766,N_18085);
nor U19687 (N_19687,N_18287,N_18489);
xnor U19688 (N_19688,N_18721,N_18200);
nand U19689 (N_19689,N_18405,N_18817);
xor U19690 (N_19690,N_18180,N_18584);
nor U19691 (N_19691,N_18292,N_18534);
nand U19692 (N_19692,N_18515,N_18976);
nand U19693 (N_19693,N_18634,N_18378);
or U19694 (N_19694,N_18695,N_18601);
nor U19695 (N_19695,N_18317,N_18235);
nand U19696 (N_19696,N_18973,N_18948);
or U19697 (N_19697,N_18873,N_18343);
xor U19698 (N_19698,N_18639,N_18974);
nand U19699 (N_19699,N_18692,N_18688);
xor U19700 (N_19700,N_18913,N_18202);
or U19701 (N_19701,N_18085,N_18565);
and U19702 (N_19702,N_18475,N_18003);
xnor U19703 (N_19703,N_18200,N_18641);
nor U19704 (N_19704,N_18514,N_18542);
nand U19705 (N_19705,N_18996,N_18527);
nor U19706 (N_19706,N_18684,N_18786);
and U19707 (N_19707,N_18818,N_18028);
and U19708 (N_19708,N_18839,N_18594);
and U19709 (N_19709,N_18602,N_18761);
xor U19710 (N_19710,N_18825,N_18630);
xor U19711 (N_19711,N_18588,N_18369);
xnor U19712 (N_19712,N_18363,N_18039);
nor U19713 (N_19713,N_18401,N_18026);
and U19714 (N_19714,N_18169,N_18281);
nand U19715 (N_19715,N_18381,N_18882);
nor U19716 (N_19716,N_18797,N_18128);
nand U19717 (N_19717,N_18337,N_18898);
nor U19718 (N_19718,N_18193,N_18370);
and U19719 (N_19719,N_18535,N_18892);
nand U19720 (N_19720,N_18067,N_18220);
nor U19721 (N_19721,N_18881,N_18161);
or U19722 (N_19722,N_18657,N_18595);
and U19723 (N_19723,N_18544,N_18783);
nand U19724 (N_19724,N_18997,N_18880);
xor U19725 (N_19725,N_18363,N_18943);
nor U19726 (N_19726,N_18438,N_18503);
nand U19727 (N_19727,N_18254,N_18213);
nand U19728 (N_19728,N_18972,N_18595);
or U19729 (N_19729,N_18211,N_18024);
or U19730 (N_19730,N_18934,N_18709);
xnor U19731 (N_19731,N_18598,N_18753);
and U19732 (N_19732,N_18745,N_18810);
xnor U19733 (N_19733,N_18855,N_18951);
nand U19734 (N_19734,N_18837,N_18912);
or U19735 (N_19735,N_18424,N_18506);
and U19736 (N_19736,N_18582,N_18879);
and U19737 (N_19737,N_18437,N_18192);
nand U19738 (N_19738,N_18820,N_18512);
or U19739 (N_19739,N_18941,N_18786);
xnor U19740 (N_19740,N_18475,N_18764);
nor U19741 (N_19741,N_18394,N_18623);
and U19742 (N_19742,N_18931,N_18384);
nor U19743 (N_19743,N_18588,N_18185);
nand U19744 (N_19744,N_18586,N_18633);
or U19745 (N_19745,N_18888,N_18799);
nand U19746 (N_19746,N_18153,N_18972);
and U19747 (N_19747,N_18920,N_18999);
xor U19748 (N_19748,N_18012,N_18462);
nor U19749 (N_19749,N_18752,N_18158);
and U19750 (N_19750,N_18895,N_18648);
and U19751 (N_19751,N_18997,N_18306);
xnor U19752 (N_19752,N_18373,N_18697);
nand U19753 (N_19753,N_18223,N_18299);
nor U19754 (N_19754,N_18697,N_18449);
nand U19755 (N_19755,N_18347,N_18138);
xnor U19756 (N_19756,N_18417,N_18846);
nor U19757 (N_19757,N_18170,N_18386);
or U19758 (N_19758,N_18440,N_18929);
or U19759 (N_19759,N_18725,N_18171);
nand U19760 (N_19760,N_18704,N_18304);
and U19761 (N_19761,N_18501,N_18725);
or U19762 (N_19762,N_18320,N_18393);
nor U19763 (N_19763,N_18204,N_18338);
xor U19764 (N_19764,N_18845,N_18824);
nor U19765 (N_19765,N_18506,N_18875);
nand U19766 (N_19766,N_18905,N_18460);
nand U19767 (N_19767,N_18482,N_18043);
nor U19768 (N_19768,N_18731,N_18293);
nand U19769 (N_19769,N_18578,N_18724);
nand U19770 (N_19770,N_18717,N_18630);
and U19771 (N_19771,N_18600,N_18782);
or U19772 (N_19772,N_18247,N_18380);
xor U19773 (N_19773,N_18611,N_18696);
or U19774 (N_19774,N_18440,N_18541);
and U19775 (N_19775,N_18753,N_18897);
nand U19776 (N_19776,N_18934,N_18240);
or U19777 (N_19777,N_18256,N_18338);
nor U19778 (N_19778,N_18747,N_18215);
nand U19779 (N_19779,N_18007,N_18445);
or U19780 (N_19780,N_18060,N_18408);
or U19781 (N_19781,N_18742,N_18805);
xnor U19782 (N_19782,N_18322,N_18445);
nor U19783 (N_19783,N_18929,N_18320);
or U19784 (N_19784,N_18159,N_18152);
nand U19785 (N_19785,N_18928,N_18942);
xor U19786 (N_19786,N_18806,N_18116);
and U19787 (N_19787,N_18551,N_18874);
or U19788 (N_19788,N_18044,N_18766);
nor U19789 (N_19789,N_18093,N_18077);
and U19790 (N_19790,N_18735,N_18927);
nand U19791 (N_19791,N_18565,N_18315);
nor U19792 (N_19792,N_18560,N_18328);
and U19793 (N_19793,N_18328,N_18573);
nand U19794 (N_19794,N_18024,N_18516);
nor U19795 (N_19795,N_18093,N_18997);
nand U19796 (N_19796,N_18615,N_18624);
nor U19797 (N_19797,N_18238,N_18983);
or U19798 (N_19798,N_18443,N_18208);
or U19799 (N_19799,N_18864,N_18211);
xor U19800 (N_19800,N_18960,N_18363);
and U19801 (N_19801,N_18330,N_18849);
nand U19802 (N_19802,N_18475,N_18690);
xor U19803 (N_19803,N_18826,N_18559);
xnor U19804 (N_19804,N_18659,N_18672);
nand U19805 (N_19805,N_18261,N_18183);
or U19806 (N_19806,N_18101,N_18424);
and U19807 (N_19807,N_18686,N_18092);
nand U19808 (N_19808,N_18486,N_18897);
xor U19809 (N_19809,N_18711,N_18708);
nor U19810 (N_19810,N_18602,N_18839);
and U19811 (N_19811,N_18391,N_18227);
nand U19812 (N_19812,N_18463,N_18516);
xnor U19813 (N_19813,N_18916,N_18705);
or U19814 (N_19814,N_18335,N_18662);
xor U19815 (N_19815,N_18982,N_18091);
nand U19816 (N_19816,N_18621,N_18082);
nand U19817 (N_19817,N_18267,N_18880);
xor U19818 (N_19818,N_18952,N_18543);
or U19819 (N_19819,N_18313,N_18107);
and U19820 (N_19820,N_18956,N_18341);
nor U19821 (N_19821,N_18026,N_18246);
and U19822 (N_19822,N_18961,N_18611);
nor U19823 (N_19823,N_18542,N_18824);
or U19824 (N_19824,N_18514,N_18258);
and U19825 (N_19825,N_18445,N_18066);
nor U19826 (N_19826,N_18111,N_18175);
and U19827 (N_19827,N_18053,N_18020);
nor U19828 (N_19828,N_18969,N_18210);
xnor U19829 (N_19829,N_18646,N_18473);
nand U19830 (N_19830,N_18045,N_18294);
nor U19831 (N_19831,N_18149,N_18491);
nand U19832 (N_19832,N_18751,N_18197);
and U19833 (N_19833,N_18920,N_18847);
nor U19834 (N_19834,N_18928,N_18790);
xnor U19835 (N_19835,N_18502,N_18149);
nand U19836 (N_19836,N_18989,N_18972);
nand U19837 (N_19837,N_18031,N_18240);
and U19838 (N_19838,N_18880,N_18948);
or U19839 (N_19839,N_18546,N_18544);
xor U19840 (N_19840,N_18265,N_18137);
nor U19841 (N_19841,N_18371,N_18173);
or U19842 (N_19842,N_18263,N_18492);
and U19843 (N_19843,N_18095,N_18950);
xnor U19844 (N_19844,N_18938,N_18283);
nor U19845 (N_19845,N_18537,N_18325);
and U19846 (N_19846,N_18369,N_18054);
nor U19847 (N_19847,N_18060,N_18542);
xnor U19848 (N_19848,N_18693,N_18894);
xnor U19849 (N_19849,N_18439,N_18332);
or U19850 (N_19850,N_18538,N_18574);
xor U19851 (N_19851,N_18444,N_18257);
nor U19852 (N_19852,N_18529,N_18875);
xnor U19853 (N_19853,N_18619,N_18351);
and U19854 (N_19854,N_18610,N_18122);
xnor U19855 (N_19855,N_18814,N_18635);
and U19856 (N_19856,N_18044,N_18638);
nand U19857 (N_19857,N_18142,N_18844);
nor U19858 (N_19858,N_18952,N_18161);
and U19859 (N_19859,N_18204,N_18211);
and U19860 (N_19860,N_18966,N_18934);
nand U19861 (N_19861,N_18208,N_18383);
nor U19862 (N_19862,N_18240,N_18164);
or U19863 (N_19863,N_18984,N_18383);
or U19864 (N_19864,N_18567,N_18392);
or U19865 (N_19865,N_18155,N_18673);
or U19866 (N_19866,N_18074,N_18720);
nand U19867 (N_19867,N_18010,N_18457);
and U19868 (N_19868,N_18392,N_18779);
and U19869 (N_19869,N_18790,N_18856);
or U19870 (N_19870,N_18373,N_18924);
or U19871 (N_19871,N_18254,N_18773);
xnor U19872 (N_19872,N_18124,N_18177);
and U19873 (N_19873,N_18194,N_18560);
or U19874 (N_19874,N_18227,N_18286);
xor U19875 (N_19875,N_18577,N_18328);
and U19876 (N_19876,N_18288,N_18057);
xor U19877 (N_19877,N_18596,N_18462);
xnor U19878 (N_19878,N_18622,N_18806);
nor U19879 (N_19879,N_18334,N_18544);
or U19880 (N_19880,N_18242,N_18484);
xor U19881 (N_19881,N_18846,N_18504);
or U19882 (N_19882,N_18308,N_18090);
xor U19883 (N_19883,N_18697,N_18748);
xor U19884 (N_19884,N_18501,N_18116);
nor U19885 (N_19885,N_18726,N_18520);
or U19886 (N_19886,N_18900,N_18126);
or U19887 (N_19887,N_18376,N_18195);
and U19888 (N_19888,N_18621,N_18899);
and U19889 (N_19889,N_18453,N_18231);
nor U19890 (N_19890,N_18272,N_18449);
nor U19891 (N_19891,N_18516,N_18575);
xor U19892 (N_19892,N_18337,N_18136);
or U19893 (N_19893,N_18229,N_18909);
or U19894 (N_19894,N_18109,N_18882);
or U19895 (N_19895,N_18412,N_18455);
and U19896 (N_19896,N_18818,N_18965);
xnor U19897 (N_19897,N_18508,N_18438);
or U19898 (N_19898,N_18654,N_18270);
nand U19899 (N_19899,N_18114,N_18789);
xor U19900 (N_19900,N_18205,N_18805);
xnor U19901 (N_19901,N_18652,N_18702);
nor U19902 (N_19902,N_18760,N_18184);
nand U19903 (N_19903,N_18905,N_18440);
xor U19904 (N_19904,N_18318,N_18367);
nand U19905 (N_19905,N_18251,N_18593);
and U19906 (N_19906,N_18500,N_18912);
nand U19907 (N_19907,N_18842,N_18138);
and U19908 (N_19908,N_18764,N_18551);
xnor U19909 (N_19909,N_18129,N_18526);
and U19910 (N_19910,N_18930,N_18009);
xnor U19911 (N_19911,N_18708,N_18472);
nand U19912 (N_19912,N_18471,N_18172);
nor U19913 (N_19913,N_18750,N_18640);
nand U19914 (N_19914,N_18977,N_18215);
nand U19915 (N_19915,N_18764,N_18769);
or U19916 (N_19916,N_18762,N_18215);
nor U19917 (N_19917,N_18485,N_18489);
nand U19918 (N_19918,N_18576,N_18810);
nand U19919 (N_19919,N_18890,N_18451);
nor U19920 (N_19920,N_18344,N_18574);
or U19921 (N_19921,N_18465,N_18382);
nand U19922 (N_19922,N_18599,N_18239);
or U19923 (N_19923,N_18584,N_18461);
nand U19924 (N_19924,N_18884,N_18536);
or U19925 (N_19925,N_18376,N_18440);
or U19926 (N_19926,N_18676,N_18562);
and U19927 (N_19927,N_18956,N_18093);
or U19928 (N_19928,N_18448,N_18544);
nor U19929 (N_19929,N_18059,N_18272);
xor U19930 (N_19930,N_18498,N_18051);
nor U19931 (N_19931,N_18161,N_18903);
xnor U19932 (N_19932,N_18434,N_18935);
xnor U19933 (N_19933,N_18392,N_18440);
nand U19934 (N_19934,N_18013,N_18938);
xor U19935 (N_19935,N_18330,N_18168);
xor U19936 (N_19936,N_18829,N_18887);
nor U19937 (N_19937,N_18905,N_18693);
xor U19938 (N_19938,N_18129,N_18774);
or U19939 (N_19939,N_18510,N_18544);
xnor U19940 (N_19940,N_18950,N_18821);
or U19941 (N_19941,N_18854,N_18614);
nor U19942 (N_19942,N_18514,N_18617);
and U19943 (N_19943,N_18578,N_18389);
nand U19944 (N_19944,N_18478,N_18385);
nor U19945 (N_19945,N_18959,N_18826);
xor U19946 (N_19946,N_18449,N_18962);
nor U19947 (N_19947,N_18377,N_18470);
xor U19948 (N_19948,N_18519,N_18587);
nor U19949 (N_19949,N_18507,N_18370);
or U19950 (N_19950,N_18183,N_18248);
or U19951 (N_19951,N_18672,N_18428);
nand U19952 (N_19952,N_18980,N_18316);
xor U19953 (N_19953,N_18379,N_18277);
or U19954 (N_19954,N_18632,N_18811);
or U19955 (N_19955,N_18437,N_18867);
xnor U19956 (N_19956,N_18440,N_18563);
and U19957 (N_19957,N_18171,N_18994);
xnor U19958 (N_19958,N_18729,N_18902);
nand U19959 (N_19959,N_18601,N_18624);
and U19960 (N_19960,N_18776,N_18401);
or U19961 (N_19961,N_18549,N_18140);
and U19962 (N_19962,N_18420,N_18668);
and U19963 (N_19963,N_18942,N_18116);
nand U19964 (N_19964,N_18204,N_18790);
and U19965 (N_19965,N_18855,N_18718);
nor U19966 (N_19966,N_18447,N_18723);
xnor U19967 (N_19967,N_18466,N_18425);
or U19968 (N_19968,N_18222,N_18597);
and U19969 (N_19969,N_18052,N_18283);
nand U19970 (N_19970,N_18527,N_18207);
and U19971 (N_19971,N_18676,N_18349);
nor U19972 (N_19972,N_18312,N_18595);
xnor U19973 (N_19973,N_18525,N_18543);
nor U19974 (N_19974,N_18612,N_18275);
nand U19975 (N_19975,N_18787,N_18615);
nand U19976 (N_19976,N_18762,N_18144);
or U19977 (N_19977,N_18296,N_18439);
xnor U19978 (N_19978,N_18547,N_18443);
or U19979 (N_19979,N_18925,N_18577);
xnor U19980 (N_19980,N_18535,N_18999);
xor U19981 (N_19981,N_18417,N_18555);
xnor U19982 (N_19982,N_18096,N_18121);
xor U19983 (N_19983,N_18065,N_18780);
nand U19984 (N_19984,N_18250,N_18925);
or U19985 (N_19985,N_18628,N_18977);
and U19986 (N_19986,N_18636,N_18706);
and U19987 (N_19987,N_18176,N_18394);
or U19988 (N_19988,N_18730,N_18611);
or U19989 (N_19989,N_18825,N_18739);
or U19990 (N_19990,N_18975,N_18587);
nand U19991 (N_19991,N_18046,N_18023);
and U19992 (N_19992,N_18046,N_18527);
nor U19993 (N_19993,N_18130,N_18887);
xor U19994 (N_19994,N_18385,N_18849);
or U19995 (N_19995,N_18940,N_18148);
xor U19996 (N_19996,N_18699,N_18171);
and U19997 (N_19997,N_18317,N_18016);
nor U19998 (N_19998,N_18946,N_18103);
nand U19999 (N_19999,N_18727,N_18572);
or U20000 (N_20000,N_19069,N_19837);
nand U20001 (N_20001,N_19872,N_19313);
nand U20002 (N_20002,N_19435,N_19421);
or U20003 (N_20003,N_19639,N_19889);
xnor U20004 (N_20004,N_19704,N_19014);
nor U20005 (N_20005,N_19006,N_19991);
nand U20006 (N_20006,N_19992,N_19750);
nand U20007 (N_20007,N_19233,N_19378);
or U20008 (N_20008,N_19795,N_19853);
nand U20009 (N_20009,N_19318,N_19713);
xor U20010 (N_20010,N_19526,N_19434);
or U20011 (N_20011,N_19416,N_19119);
xnor U20012 (N_20012,N_19007,N_19392);
nor U20013 (N_20013,N_19640,N_19855);
and U20014 (N_20014,N_19535,N_19386);
nand U20015 (N_20015,N_19128,N_19338);
and U20016 (N_20016,N_19781,N_19273);
nor U20017 (N_20017,N_19275,N_19624);
nand U20018 (N_20018,N_19364,N_19223);
and U20019 (N_20019,N_19465,N_19210);
or U20020 (N_20020,N_19383,N_19193);
or U20021 (N_20021,N_19179,N_19442);
xor U20022 (N_20022,N_19931,N_19924);
nor U20023 (N_20023,N_19280,N_19057);
xor U20024 (N_20024,N_19360,N_19423);
xor U20025 (N_20025,N_19265,N_19954);
nand U20026 (N_20026,N_19824,N_19212);
nand U20027 (N_20027,N_19870,N_19940);
nor U20028 (N_20028,N_19612,N_19956);
xor U20029 (N_20029,N_19091,N_19946);
nor U20030 (N_20030,N_19926,N_19550);
nand U20031 (N_20031,N_19455,N_19646);
nor U20032 (N_20032,N_19463,N_19860);
nor U20033 (N_20033,N_19437,N_19938);
nor U20034 (N_20034,N_19122,N_19614);
nand U20035 (N_20035,N_19020,N_19753);
and U20036 (N_20036,N_19784,N_19677);
nand U20037 (N_20037,N_19482,N_19089);
nand U20038 (N_20038,N_19398,N_19257);
xor U20039 (N_20039,N_19365,N_19228);
nor U20040 (N_20040,N_19635,N_19008);
xor U20041 (N_20041,N_19335,N_19145);
xnor U20042 (N_20042,N_19272,N_19429);
nor U20043 (N_20043,N_19914,N_19224);
nor U20044 (N_20044,N_19412,N_19654);
nor U20045 (N_20045,N_19552,N_19950);
nor U20046 (N_20046,N_19922,N_19314);
nand U20047 (N_20047,N_19194,N_19116);
nand U20048 (N_20048,N_19137,N_19765);
xnor U20049 (N_20049,N_19984,N_19351);
and U20050 (N_20050,N_19808,N_19969);
xor U20051 (N_20051,N_19915,N_19407);
xnor U20052 (N_20052,N_19250,N_19754);
or U20053 (N_20053,N_19425,N_19086);
nor U20054 (N_20054,N_19447,N_19214);
nand U20055 (N_20055,N_19773,N_19133);
nor U20056 (N_20056,N_19545,N_19177);
xor U20057 (N_20057,N_19740,N_19816);
and U20058 (N_20058,N_19131,N_19221);
and U20059 (N_20059,N_19797,N_19839);
or U20060 (N_20060,N_19592,N_19042);
or U20061 (N_20061,N_19075,N_19655);
xnor U20062 (N_20062,N_19026,N_19236);
and U20063 (N_20063,N_19380,N_19905);
xnor U20064 (N_20064,N_19293,N_19348);
nor U20065 (N_20065,N_19717,N_19032);
or U20066 (N_20066,N_19185,N_19162);
nand U20067 (N_20067,N_19762,N_19722);
and U20068 (N_20068,N_19710,N_19217);
or U20069 (N_20069,N_19671,N_19157);
xnor U20070 (N_20070,N_19589,N_19268);
or U20071 (N_20071,N_19777,N_19166);
or U20072 (N_20072,N_19143,N_19763);
nand U20073 (N_20073,N_19935,N_19325);
or U20074 (N_20074,N_19300,N_19106);
or U20075 (N_20075,N_19527,N_19331);
nor U20076 (N_20076,N_19579,N_19315);
nand U20077 (N_20077,N_19203,N_19319);
xor U20078 (N_20078,N_19323,N_19049);
and U20079 (N_20079,N_19601,N_19670);
nor U20080 (N_20080,N_19349,N_19130);
nor U20081 (N_20081,N_19531,N_19154);
nand U20082 (N_20082,N_19693,N_19522);
xnor U20083 (N_20083,N_19358,N_19947);
nor U20084 (N_20084,N_19818,N_19321);
nor U20085 (N_20085,N_19475,N_19371);
or U20086 (N_20086,N_19517,N_19674);
and U20087 (N_20087,N_19936,N_19793);
and U20088 (N_20088,N_19500,N_19833);
xor U20089 (N_20089,N_19481,N_19381);
nand U20090 (N_20090,N_19827,N_19508);
nand U20091 (N_20091,N_19473,N_19484);
nand U20092 (N_20092,N_19192,N_19735);
or U20093 (N_20093,N_19011,N_19259);
and U20094 (N_20094,N_19172,N_19847);
and U20095 (N_20095,N_19749,N_19974);
and U20096 (N_20096,N_19188,N_19752);
xnor U20097 (N_20097,N_19311,N_19418);
xor U20098 (N_20098,N_19232,N_19714);
xnor U20099 (N_20099,N_19967,N_19189);
nor U20100 (N_20100,N_19397,N_19342);
xnor U20101 (N_20101,N_19098,N_19600);
xnor U20102 (N_20102,N_19852,N_19841);
nor U20103 (N_20103,N_19241,N_19458);
and U20104 (N_20104,N_19685,N_19553);
or U20105 (N_20105,N_19705,N_19389);
or U20106 (N_20106,N_19979,N_19730);
and U20107 (N_20107,N_19766,N_19696);
nand U20108 (N_20108,N_19976,N_19524);
nor U20109 (N_20109,N_19387,N_19151);
xor U20110 (N_20110,N_19316,N_19565);
nand U20111 (N_20111,N_19768,N_19022);
or U20112 (N_20112,N_19863,N_19037);
nor U20113 (N_20113,N_19461,N_19489);
or U20114 (N_20114,N_19448,N_19664);
nand U20115 (N_20115,N_19220,N_19972);
or U20116 (N_20116,N_19453,N_19557);
or U20117 (N_20117,N_19000,N_19549);
and U20118 (N_20118,N_19343,N_19288);
nor U20119 (N_20119,N_19728,N_19799);
or U20120 (N_20120,N_19887,N_19965);
nand U20121 (N_20121,N_19604,N_19650);
xor U20122 (N_20122,N_19875,N_19372);
and U20123 (N_20123,N_19252,N_19046);
nand U20124 (N_20124,N_19541,N_19711);
nand U20125 (N_20125,N_19036,N_19836);
or U20126 (N_20126,N_19138,N_19977);
or U20127 (N_20127,N_19105,N_19809);
nor U20128 (N_20128,N_19647,N_19506);
nor U20129 (N_20129,N_19509,N_19010);
xor U20130 (N_20130,N_19699,N_19480);
xor U20131 (N_20131,N_19227,N_19457);
and U20132 (N_20132,N_19444,N_19814);
xnor U20133 (N_20133,N_19053,N_19634);
xnor U20134 (N_20134,N_19211,N_19216);
xor U20135 (N_20135,N_19230,N_19726);
nand U20136 (N_20136,N_19225,N_19200);
or U20137 (N_20137,N_19487,N_19276);
nand U20138 (N_20138,N_19867,N_19488);
nand U20139 (N_20139,N_19219,N_19174);
nand U20140 (N_20140,N_19414,N_19460);
nand U20141 (N_20141,N_19987,N_19045);
nor U20142 (N_20142,N_19994,N_19708);
xnor U20143 (N_20143,N_19952,N_19433);
nand U20144 (N_20144,N_19208,N_19932);
and U20145 (N_20145,N_19981,N_19783);
nand U20146 (N_20146,N_19663,N_19391);
or U20147 (N_20147,N_19953,N_19761);
xor U20148 (N_20148,N_19238,N_19540);
nand U20149 (N_20149,N_19732,N_19619);
nand U20150 (N_20150,N_19470,N_19377);
nor U20151 (N_20151,N_19408,N_19337);
nand U20152 (N_20152,N_19196,N_19782);
xor U20153 (N_20153,N_19543,N_19874);
and U20154 (N_20154,N_19684,N_19385);
xor U20155 (N_20155,N_19806,N_19001);
xnor U20156 (N_20156,N_19712,N_19110);
xor U20157 (N_20157,N_19755,N_19430);
xnor U20158 (N_20158,N_19747,N_19253);
or U20159 (N_20159,N_19835,N_19111);
xnor U20160 (N_20160,N_19849,N_19563);
and U20161 (N_20161,N_19090,N_19595);
and U20162 (N_20162,N_19529,N_19249);
or U20163 (N_20163,N_19409,N_19577);
and U20164 (N_20164,N_19184,N_19801);
nand U20165 (N_20165,N_19702,N_19082);
and U20166 (N_20166,N_19518,N_19041);
or U20167 (N_20167,N_19993,N_19738);
nor U20168 (N_20168,N_19558,N_19181);
and U20169 (N_20169,N_19050,N_19155);
or U20170 (N_20170,N_19919,N_19842);
nor U20171 (N_20171,N_19477,N_19975);
xor U20172 (N_20172,N_19422,N_19998);
nor U20173 (N_20173,N_19637,N_19132);
and U20174 (N_20174,N_19695,N_19051);
nand U20175 (N_20175,N_19078,N_19024);
nor U20176 (N_20176,N_19396,N_19958);
or U20177 (N_20177,N_19148,N_19995);
or U20178 (N_20178,N_19094,N_19368);
or U20179 (N_20179,N_19725,N_19744);
nor U20180 (N_20180,N_19892,N_19556);
nand U20181 (N_20181,N_19893,N_19894);
and U20182 (N_20182,N_19060,N_19564);
or U20183 (N_20183,N_19403,N_19114);
nand U20184 (N_20184,N_19729,N_19141);
or U20185 (N_20185,N_19301,N_19356);
xnor U20186 (N_20186,N_19811,N_19819);
xor U20187 (N_20187,N_19048,N_19838);
xor U20188 (N_20188,N_19928,N_19978);
and U20189 (N_20189,N_19018,N_19546);
nor U20190 (N_20190,N_19848,N_19679);
or U20191 (N_20191,N_19446,N_19332);
nor U20192 (N_20192,N_19027,N_19675);
nand U20193 (N_20193,N_19017,N_19317);
nand U20194 (N_20194,N_19786,N_19539);
nand U20195 (N_20195,N_19845,N_19617);
nand U20196 (N_20196,N_19748,N_19622);
and U20197 (N_20197,N_19254,N_19247);
nor U20198 (N_20198,N_19582,N_19996);
or U20199 (N_20199,N_19731,N_19873);
nor U20200 (N_20200,N_19350,N_19573);
xnor U20201 (N_20201,N_19034,N_19876);
xor U20202 (N_20202,N_19906,N_19080);
xor U20203 (N_20203,N_19016,N_19913);
or U20204 (N_20204,N_19340,N_19537);
nand U20205 (N_20205,N_19721,N_19469);
nand U20206 (N_20206,N_19934,N_19980);
or U20207 (N_20207,N_19346,N_19633);
xnor U20208 (N_20208,N_19896,N_19339);
xnor U20209 (N_20209,N_19099,N_19333);
nand U20210 (N_20210,N_19596,N_19279);
or U20211 (N_20211,N_19347,N_19180);
nor U20212 (N_20212,N_19511,N_19746);
nor U20213 (N_20213,N_19644,N_19353);
nor U20214 (N_20214,N_19440,N_19419);
nor U20215 (N_20215,N_19076,N_19520);
nand U20216 (N_20216,N_19760,N_19178);
nor U20217 (N_20217,N_19474,N_19160);
xor U20218 (N_20218,N_19191,N_19720);
or U20219 (N_20219,N_19903,N_19941);
nand U20220 (N_20220,N_19400,N_19428);
nand U20221 (N_20221,N_19459,N_19983);
nand U20222 (N_20222,N_19308,N_19052);
or U20223 (N_20223,N_19411,N_19706);
nor U20224 (N_20224,N_19585,N_19124);
and U20225 (N_20225,N_19864,N_19840);
or U20226 (N_20226,N_19395,N_19410);
or U20227 (N_20227,N_19656,N_19108);
and U20228 (N_20228,N_19492,N_19464);
and U20229 (N_20229,N_19576,N_19921);
nand U20230 (N_20230,N_19101,N_19676);
or U20231 (N_20231,N_19070,N_19613);
nor U20232 (N_20232,N_19158,N_19843);
nand U20233 (N_20233,N_19902,N_19586);
nor U20234 (N_20234,N_19569,N_19590);
xnor U20235 (N_20235,N_19519,N_19774);
nor U20236 (N_20236,N_19989,N_19320);
nor U20237 (N_20237,N_19067,N_19112);
nor U20238 (N_20238,N_19190,N_19282);
and U20239 (N_20239,N_19606,N_19496);
or U20240 (N_20240,N_19019,N_19631);
or U20241 (N_20241,N_19528,N_19491);
nor U20242 (N_20242,N_19587,N_19334);
or U20243 (N_20243,N_19013,N_19680);
and U20244 (N_20244,N_19832,N_19466);
nand U20245 (N_20245,N_19575,N_19583);
or U20246 (N_20246,N_19502,N_19697);
nand U20247 (N_20247,N_19248,N_19555);
and U20248 (N_20248,N_19884,N_19891);
and U20249 (N_20249,N_19904,N_19197);
or U20250 (N_20250,N_19206,N_19629);
or U20251 (N_20251,N_19169,N_19035);
nand U20252 (N_20252,N_19649,N_19562);
nor U20253 (N_20253,N_19881,N_19054);
nand U20254 (N_20254,N_19363,N_19431);
nand U20255 (N_20255,N_19739,N_19770);
or U20256 (N_20256,N_19716,N_19719);
and U20257 (N_20257,N_19789,N_19507);
nor U20258 (N_20258,N_19741,N_19426);
nand U20259 (N_20259,N_19957,N_19361);
nor U20260 (N_20260,N_19886,N_19087);
or U20261 (N_20261,N_19767,N_19285);
xor U20262 (N_20262,N_19736,N_19256);
or U20263 (N_20263,N_19682,N_19462);
xnor U20264 (N_20264,N_19805,N_19084);
xnor U20265 (N_20265,N_19305,N_19775);
nor U20266 (N_20266,N_19756,N_19999);
xnor U20267 (N_20267,N_19149,N_19165);
xor U20268 (N_20268,N_19264,N_19287);
nor U20269 (N_20269,N_19689,N_19505);
nand U20270 (N_20270,N_19616,N_19064);
nand U20271 (N_20271,N_19572,N_19261);
nor U20272 (N_20272,N_19375,N_19780);
or U20273 (N_20273,N_19023,N_19794);
xor U20274 (N_20274,N_19910,N_19846);
or U20275 (N_20275,N_19530,N_19943);
or U20276 (N_20276,N_19388,N_19497);
and U20277 (N_20277,N_19907,N_19742);
and U20278 (N_20278,N_19594,N_19115);
xor U20279 (N_20279,N_19439,N_19015);
and U20280 (N_20280,N_19199,N_19127);
xnor U20281 (N_20281,N_19571,N_19504);
nand U20282 (N_20282,N_19501,N_19370);
and U20283 (N_20283,N_19374,N_19920);
xnor U20284 (N_20284,N_19997,N_19289);
nand U20285 (N_20285,N_19503,N_19328);
or U20286 (N_20286,N_19125,N_19865);
nor U20287 (N_20287,N_19290,N_19665);
nand U20288 (N_20288,N_19513,N_19559);
and U20289 (N_20289,N_19605,N_19692);
xor U20290 (N_20290,N_19263,N_19858);
nand U20291 (N_20291,N_19871,N_19669);
nor U20292 (N_20292,N_19204,N_19467);
and U20293 (N_20293,N_19445,N_19142);
xnor U20294 (N_20294,N_19610,N_19869);
xnor U20295 (N_20295,N_19798,N_19175);
nand U20296 (N_20296,N_19608,N_19292);
or U20297 (N_20297,N_19628,N_19945);
and U20298 (N_20298,N_19405,N_19862);
or U20299 (N_20299,N_19703,N_19955);
and U20300 (N_20300,N_19096,N_19698);
or U20301 (N_20301,N_19615,N_19468);
xnor U20302 (N_20302,N_19104,N_19986);
or U20303 (N_20303,N_19866,N_19031);
xnor U20304 (N_20304,N_19415,N_19072);
nand U20305 (N_20305,N_19788,N_19059);
xor U20306 (N_20306,N_19776,N_19183);
or U20307 (N_20307,N_19968,N_19079);
or U20308 (N_20308,N_19927,N_19369);
and U20309 (N_20309,N_19933,N_19146);
nand U20310 (N_20310,N_19578,N_19478);
xnor U20311 (N_20311,N_19345,N_19493);
or U20312 (N_20312,N_19850,N_19456);
nand U20313 (N_20313,N_19909,N_19851);
nor U20314 (N_20314,N_19085,N_19450);
xnor U20315 (N_20315,N_19362,N_19088);
xnor U20316 (N_20316,N_19294,N_19651);
or U20317 (N_20317,N_19299,N_19286);
or U20318 (N_20318,N_19231,N_19771);
nand U20319 (N_20319,N_19690,N_19267);
and U20320 (N_20320,N_19355,N_19427);
nand U20321 (N_20321,N_19802,N_19751);
nand U20322 (N_20322,N_19939,N_19393);
nand U20323 (N_20323,N_19525,N_19964);
or U20324 (N_20324,N_19150,N_19672);
nand U20325 (N_20325,N_19588,N_19218);
or U20326 (N_20326,N_19709,N_19176);
xnor U20327 (N_20327,N_19681,N_19198);
and U20328 (N_20328,N_19658,N_19516);
and U20329 (N_20329,N_19688,N_19718);
nor U20330 (N_20330,N_19260,N_19109);
xor U20331 (N_20331,N_19081,N_19548);
xor U20332 (N_20332,N_19533,N_19195);
nand U20333 (N_20333,N_19973,N_19044);
nor U20334 (N_20334,N_19673,N_19899);
or U20335 (N_20335,N_19630,N_19424);
or U20336 (N_20336,N_19171,N_19170);
or U20337 (N_20337,N_19844,N_19694);
nand U20338 (N_20338,N_19598,N_19376);
nor U20339 (N_20339,N_19599,N_19068);
or U20340 (N_20340,N_19554,N_19187);
xor U20341 (N_20341,N_19215,N_19274);
xnor U20342 (N_20342,N_19800,N_19297);
or U20343 (N_20343,N_19144,N_19560);
or U20344 (N_20344,N_19820,N_19627);
and U20345 (N_20345,N_19542,N_19055);
nor U20346 (N_20346,N_19061,N_19373);
nor U20347 (N_20347,N_19657,N_19164);
nand U20348 (N_20348,N_19944,N_19234);
nand U20349 (N_20349,N_19772,N_19025);
and U20350 (N_20350,N_19226,N_19602);
and U20351 (N_20351,N_19757,N_19514);
or U20352 (N_20352,N_19071,N_19494);
or U20353 (N_20353,N_19004,N_19607);
nand U20354 (N_20354,N_19012,N_19966);
nand U20355 (N_20355,N_19566,N_19161);
and U20356 (N_20356,N_19420,N_19123);
and U20357 (N_20357,N_19399,N_19534);
xor U20358 (N_20358,N_19636,N_19591);
nor U20359 (N_20359,N_19113,N_19344);
nand U20360 (N_20360,N_19073,N_19291);
or U20361 (N_20361,N_19390,N_19406);
xor U20362 (N_20362,N_19003,N_19413);
nand U20363 (N_20363,N_19126,N_19861);
or U20364 (N_20364,N_19483,N_19021);
nand U20365 (N_20365,N_19296,N_19700);
or U20366 (N_20366,N_19538,N_19937);
and U20367 (N_20367,N_19764,N_19618);
nand U20368 (N_20368,N_19173,N_19471);
nor U20369 (N_20369,N_19499,N_19152);
nor U20370 (N_20370,N_19107,N_19322);
and U20371 (N_20371,N_19925,N_19182);
nand U20372 (N_20372,N_19779,N_19120);
nor U20373 (N_20373,N_19402,N_19310);
and U20374 (N_20374,N_19298,N_19597);
nor U20375 (N_20375,N_19923,N_19454);
nand U20376 (N_20376,N_19785,N_19515);
and U20377 (N_20377,N_19336,N_19235);
and U20378 (N_20378,N_19229,N_19822);
nand U20379 (N_20379,N_19312,N_19441);
and U20380 (N_20380,N_19495,N_19118);
xnor U20381 (N_20381,N_19960,N_19643);
xnor U20382 (N_20382,N_19038,N_19258);
nand U20383 (N_20383,N_19401,N_19168);
or U20384 (N_20384,N_19095,N_19666);
nor U20385 (N_20385,N_19568,N_19066);
nand U20386 (N_20386,N_19432,N_19009);
and U20387 (N_20387,N_19813,N_19829);
xnor U20388 (N_20388,N_19417,N_19544);
and U20389 (N_20389,N_19707,N_19790);
and U20390 (N_20390,N_19733,N_19092);
nor U20391 (N_20391,N_19830,N_19240);
or U20392 (N_20392,N_19625,N_19201);
or U20393 (N_20393,N_19859,N_19611);
nand U20394 (N_20394,N_19898,N_19030);
or U20395 (N_20395,N_19567,N_19490);
or U20396 (N_20396,N_19638,N_19367);
xnor U20397 (N_20397,N_19136,N_19683);
nand U20398 (N_20398,N_19277,N_19121);
and U20399 (N_20399,N_19701,N_19498);
or U20400 (N_20400,N_19281,N_19159);
and U20401 (N_20401,N_19948,N_19056);
nand U20402 (N_20402,N_19880,N_19626);
xnor U20403 (N_20403,N_19438,N_19882);
nand U20404 (N_20404,N_19062,N_19510);
nand U20405 (N_20405,N_19737,N_19778);
nor U20406 (N_20406,N_19479,N_19900);
nor U20407 (N_20407,N_19825,N_19352);
nand U20408 (N_20408,N_19834,N_19621);
xor U20409 (N_20409,N_19888,N_19817);
and U20410 (N_20410,N_19959,N_19269);
and U20411 (N_20411,N_19807,N_19942);
xnor U20412 (N_20412,N_19140,N_19270);
nand U20413 (N_20413,N_19584,N_19803);
and U20414 (N_20414,N_19243,N_19202);
or U20415 (N_20415,N_19245,N_19156);
nor U20416 (N_20416,N_19284,N_19890);
and U20417 (N_20417,N_19341,N_19963);
and U20418 (N_20418,N_19662,N_19436);
and U20419 (N_20419,N_19359,N_19603);
or U20420 (N_20420,N_19304,N_19028);
or U20421 (N_20421,N_19758,N_19306);
nand U20422 (N_20422,N_19812,N_19971);
or U20423 (N_20423,N_19970,N_19723);
nor U20424 (N_20424,N_19623,N_19209);
nand U20425 (N_20425,N_19796,N_19961);
nor U20426 (N_20426,N_19828,N_19329);
or U20427 (N_20427,N_19734,N_19632);
xor U20428 (N_20428,N_19661,N_19678);
nand U20429 (N_20429,N_19382,N_19213);
or U20430 (N_20430,N_19951,N_19916);
or U20431 (N_20431,N_19791,N_19384);
or U20432 (N_20432,N_19283,N_19394);
or U20433 (N_20433,N_19033,N_19523);
and U20434 (N_20434,N_19877,N_19854);
and U20435 (N_20435,N_19668,N_19532);
nand U20436 (N_20436,N_19810,N_19574);
nand U20437 (N_20437,N_19404,N_19047);
nand U20438 (N_20438,N_19379,N_19593);
or U20439 (N_20439,N_19687,N_19988);
nor U20440 (N_20440,N_19883,N_19823);
or U20441 (N_20441,N_19911,N_19357);
or U20442 (N_20442,N_19065,N_19645);
and U20443 (N_20443,N_19237,N_19985);
nand U20444 (N_20444,N_19239,N_19485);
and U20445 (N_20445,N_19512,N_19787);
and U20446 (N_20446,N_19135,N_19912);
or U20447 (N_20447,N_19153,N_19759);
nand U20448 (N_20448,N_19570,N_19609);
or U20449 (N_20449,N_19580,N_19255);
and U20450 (N_20450,N_19930,N_19652);
nor U20451 (N_20451,N_19536,N_19354);
nor U20452 (N_20452,N_19100,N_19083);
xor U20453 (N_20453,N_19309,N_19831);
or U20454 (N_20454,N_19648,N_19727);
nand U20455 (N_20455,N_19222,N_19581);
nand U20456 (N_20456,N_19002,N_19792);
xor U20457 (N_20457,N_19908,N_19246);
and U20458 (N_20458,N_19443,N_19660);
nor U20459 (N_20459,N_19163,N_19895);
or U20460 (N_20460,N_19302,N_19029);
or U20461 (N_20461,N_19278,N_19307);
xnor U20462 (N_20462,N_19561,N_19897);
xor U20463 (N_20463,N_19667,N_19366);
nor U20464 (N_20464,N_19005,N_19452);
nand U20465 (N_20465,N_19476,N_19821);
and U20466 (N_20466,N_19074,N_19769);
nand U20467 (N_20467,N_19857,N_19547);
or U20468 (N_20468,N_19917,N_19097);
nand U20469 (N_20469,N_19990,N_19949);
and U20470 (N_20470,N_19326,N_19451);
nand U20471 (N_20471,N_19743,N_19878);
nor U20472 (N_20472,N_19620,N_19167);
and U20473 (N_20473,N_19962,N_19918);
nand U20474 (N_20474,N_19103,N_19521);
nor U20475 (N_20475,N_19129,N_19271);
xnor U20476 (N_20476,N_19885,N_19815);
or U20477 (N_20477,N_19879,N_19244);
nand U20478 (N_20478,N_19826,N_19659);
nand U20479 (N_20479,N_19040,N_19134);
xor U20480 (N_20480,N_19093,N_19686);
nor U20481 (N_20481,N_19868,N_19715);
nand U20482 (N_20482,N_19242,N_19472);
and U20483 (N_20483,N_19186,N_19207);
and U20484 (N_20484,N_19262,N_19295);
or U20485 (N_20485,N_19058,N_19901);
and U20486 (N_20486,N_19691,N_19330);
nand U20487 (N_20487,N_19063,N_19303);
and U20488 (N_20488,N_19724,N_19641);
nand U20489 (N_20489,N_19745,N_19642);
and U20490 (N_20490,N_19139,N_19929);
nor U20491 (N_20491,N_19147,N_19117);
xnor U20492 (N_20492,N_19039,N_19856);
or U20493 (N_20493,N_19043,N_19251);
nand U20494 (N_20494,N_19486,N_19653);
and U20495 (N_20495,N_19102,N_19449);
nor U20496 (N_20496,N_19551,N_19324);
nor U20497 (N_20497,N_19804,N_19327);
nand U20498 (N_20498,N_19205,N_19077);
nand U20499 (N_20499,N_19982,N_19266);
and U20500 (N_20500,N_19074,N_19982);
nor U20501 (N_20501,N_19908,N_19804);
and U20502 (N_20502,N_19414,N_19888);
and U20503 (N_20503,N_19448,N_19568);
nor U20504 (N_20504,N_19575,N_19147);
or U20505 (N_20505,N_19634,N_19756);
nand U20506 (N_20506,N_19369,N_19892);
nand U20507 (N_20507,N_19023,N_19807);
and U20508 (N_20508,N_19051,N_19347);
nand U20509 (N_20509,N_19738,N_19347);
nor U20510 (N_20510,N_19208,N_19164);
nand U20511 (N_20511,N_19546,N_19379);
nand U20512 (N_20512,N_19975,N_19259);
xor U20513 (N_20513,N_19185,N_19175);
xnor U20514 (N_20514,N_19743,N_19273);
and U20515 (N_20515,N_19372,N_19449);
nor U20516 (N_20516,N_19884,N_19735);
or U20517 (N_20517,N_19995,N_19059);
and U20518 (N_20518,N_19329,N_19713);
xor U20519 (N_20519,N_19982,N_19909);
and U20520 (N_20520,N_19772,N_19812);
xnor U20521 (N_20521,N_19157,N_19124);
or U20522 (N_20522,N_19759,N_19848);
or U20523 (N_20523,N_19476,N_19344);
xor U20524 (N_20524,N_19224,N_19155);
or U20525 (N_20525,N_19482,N_19693);
nor U20526 (N_20526,N_19609,N_19630);
and U20527 (N_20527,N_19681,N_19561);
xnor U20528 (N_20528,N_19648,N_19387);
nand U20529 (N_20529,N_19557,N_19369);
nor U20530 (N_20530,N_19786,N_19389);
nand U20531 (N_20531,N_19190,N_19191);
xor U20532 (N_20532,N_19327,N_19782);
xnor U20533 (N_20533,N_19515,N_19327);
or U20534 (N_20534,N_19468,N_19949);
and U20535 (N_20535,N_19948,N_19632);
xnor U20536 (N_20536,N_19460,N_19248);
nor U20537 (N_20537,N_19755,N_19944);
xnor U20538 (N_20538,N_19496,N_19068);
or U20539 (N_20539,N_19754,N_19345);
xnor U20540 (N_20540,N_19929,N_19236);
xnor U20541 (N_20541,N_19030,N_19511);
nor U20542 (N_20542,N_19192,N_19557);
xnor U20543 (N_20543,N_19521,N_19186);
xor U20544 (N_20544,N_19863,N_19991);
and U20545 (N_20545,N_19807,N_19087);
or U20546 (N_20546,N_19505,N_19357);
and U20547 (N_20547,N_19121,N_19182);
nor U20548 (N_20548,N_19555,N_19581);
nand U20549 (N_20549,N_19077,N_19204);
nand U20550 (N_20550,N_19036,N_19237);
nor U20551 (N_20551,N_19188,N_19957);
nand U20552 (N_20552,N_19931,N_19780);
or U20553 (N_20553,N_19612,N_19958);
nand U20554 (N_20554,N_19067,N_19007);
or U20555 (N_20555,N_19319,N_19120);
and U20556 (N_20556,N_19137,N_19309);
and U20557 (N_20557,N_19504,N_19966);
xor U20558 (N_20558,N_19577,N_19478);
or U20559 (N_20559,N_19308,N_19831);
xnor U20560 (N_20560,N_19603,N_19997);
nor U20561 (N_20561,N_19412,N_19786);
or U20562 (N_20562,N_19230,N_19332);
nor U20563 (N_20563,N_19429,N_19706);
or U20564 (N_20564,N_19074,N_19140);
and U20565 (N_20565,N_19359,N_19310);
xnor U20566 (N_20566,N_19290,N_19301);
or U20567 (N_20567,N_19413,N_19641);
or U20568 (N_20568,N_19508,N_19281);
nor U20569 (N_20569,N_19325,N_19728);
and U20570 (N_20570,N_19974,N_19645);
nor U20571 (N_20571,N_19630,N_19927);
nor U20572 (N_20572,N_19471,N_19725);
and U20573 (N_20573,N_19531,N_19606);
nor U20574 (N_20574,N_19105,N_19531);
xor U20575 (N_20575,N_19459,N_19856);
xnor U20576 (N_20576,N_19619,N_19570);
and U20577 (N_20577,N_19029,N_19033);
nand U20578 (N_20578,N_19380,N_19587);
nand U20579 (N_20579,N_19085,N_19411);
or U20580 (N_20580,N_19611,N_19877);
and U20581 (N_20581,N_19278,N_19019);
nor U20582 (N_20582,N_19566,N_19051);
nand U20583 (N_20583,N_19204,N_19303);
nand U20584 (N_20584,N_19783,N_19978);
nand U20585 (N_20585,N_19627,N_19102);
and U20586 (N_20586,N_19615,N_19735);
nor U20587 (N_20587,N_19203,N_19115);
and U20588 (N_20588,N_19583,N_19561);
xor U20589 (N_20589,N_19852,N_19550);
or U20590 (N_20590,N_19213,N_19976);
nor U20591 (N_20591,N_19237,N_19597);
xor U20592 (N_20592,N_19188,N_19637);
and U20593 (N_20593,N_19394,N_19190);
and U20594 (N_20594,N_19902,N_19918);
nand U20595 (N_20595,N_19668,N_19158);
or U20596 (N_20596,N_19079,N_19047);
and U20597 (N_20597,N_19752,N_19758);
and U20598 (N_20598,N_19118,N_19282);
nor U20599 (N_20599,N_19322,N_19997);
or U20600 (N_20600,N_19303,N_19778);
nand U20601 (N_20601,N_19611,N_19678);
or U20602 (N_20602,N_19622,N_19793);
nor U20603 (N_20603,N_19533,N_19683);
and U20604 (N_20604,N_19398,N_19404);
or U20605 (N_20605,N_19622,N_19187);
nor U20606 (N_20606,N_19973,N_19153);
or U20607 (N_20607,N_19287,N_19766);
or U20608 (N_20608,N_19635,N_19007);
nand U20609 (N_20609,N_19157,N_19151);
xor U20610 (N_20610,N_19878,N_19727);
nor U20611 (N_20611,N_19908,N_19220);
and U20612 (N_20612,N_19258,N_19895);
nor U20613 (N_20613,N_19843,N_19029);
xor U20614 (N_20614,N_19380,N_19845);
nor U20615 (N_20615,N_19761,N_19428);
nand U20616 (N_20616,N_19141,N_19333);
and U20617 (N_20617,N_19041,N_19253);
nand U20618 (N_20618,N_19671,N_19878);
xnor U20619 (N_20619,N_19534,N_19915);
nand U20620 (N_20620,N_19174,N_19904);
nand U20621 (N_20621,N_19815,N_19006);
nor U20622 (N_20622,N_19302,N_19487);
nor U20623 (N_20623,N_19907,N_19514);
and U20624 (N_20624,N_19843,N_19969);
and U20625 (N_20625,N_19055,N_19314);
or U20626 (N_20626,N_19601,N_19522);
nand U20627 (N_20627,N_19289,N_19334);
nor U20628 (N_20628,N_19110,N_19473);
nor U20629 (N_20629,N_19752,N_19614);
xnor U20630 (N_20630,N_19849,N_19023);
or U20631 (N_20631,N_19944,N_19388);
nor U20632 (N_20632,N_19269,N_19667);
nand U20633 (N_20633,N_19631,N_19778);
nor U20634 (N_20634,N_19906,N_19133);
and U20635 (N_20635,N_19041,N_19602);
nand U20636 (N_20636,N_19403,N_19589);
and U20637 (N_20637,N_19347,N_19835);
nor U20638 (N_20638,N_19762,N_19988);
xor U20639 (N_20639,N_19054,N_19703);
nand U20640 (N_20640,N_19348,N_19620);
and U20641 (N_20641,N_19429,N_19896);
xor U20642 (N_20642,N_19217,N_19745);
or U20643 (N_20643,N_19211,N_19880);
nor U20644 (N_20644,N_19240,N_19683);
nor U20645 (N_20645,N_19146,N_19910);
xnor U20646 (N_20646,N_19391,N_19180);
or U20647 (N_20647,N_19708,N_19065);
or U20648 (N_20648,N_19606,N_19267);
nor U20649 (N_20649,N_19827,N_19131);
nor U20650 (N_20650,N_19197,N_19146);
and U20651 (N_20651,N_19801,N_19236);
xor U20652 (N_20652,N_19116,N_19887);
or U20653 (N_20653,N_19223,N_19704);
and U20654 (N_20654,N_19965,N_19473);
or U20655 (N_20655,N_19371,N_19584);
xnor U20656 (N_20656,N_19820,N_19422);
or U20657 (N_20657,N_19679,N_19928);
or U20658 (N_20658,N_19253,N_19734);
or U20659 (N_20659,N_19237,N_19365);
and U20660 (N_20660,N_19242,N_19925);
and U20661 (N_20661,N_19786,N_19123);
nor U20662 (N_20662,N_19377,N_19834);
and U20663 (N_20663,N_19973,N_19560);
and U20664 (N_20664,N_19224,N_19505);
xor U20665 (N_20665,N_19723,N_19748);
and U20666 (N_20666,N_19667,N_19599);
nand U20667 (N_20667,N_19486,N_19264);
or U20668 (N_20668,N_19506,N_19976);
or U20669 (N_20669,N_19777,N_19099);
and U20670 (N_20670,N_19388,N_19007);
xnor U20671 (N_20671,N_19460,N_19572);
and U20672 (N_20672,N_19891,N_19710);
nor U20673 (N_20673,N_19810,N_19257);
and U20674 (N_20674,N_19851,N_19726);
xnor U20675 (N_20675,N_19119,N_19797);
and U20676 (N_20676,N_19512,N_19672);
and U20677 (N_20677,N_19173,N_19888);
nor U20678 (N_20678,N_19971,N_19233);
or U20679 (N_20679,N_19216,N_19426);
nor U20680 (N_20680,N_19471,N_19902);
and U20681 (N_20681,N_19570,N_19577);
or U20682 (N_20682,N_19727,N_19628);
xnor U20683 (N_20683,N_19711,N_19625);
and U20684 (N_20684,N_19232,N_19566);
nand U20685 (N_20685,N_19587,N_19427);
xor U20686 (N_20686,N_19713,N_19283);
and U20687 (N_20687,N_19165,N_19710);
or U20688 (N_20688,N_19281,N_19457);
or U20689 (N_20689,N_19011,N_19087);
nand U20690 (N_20690,N_19293,N_19183);
xnor U20691 (N_20691,N_19490,N_19275);
nor U20692 (N_20692,N_19977,N_19399);
nor U20693 (N_20693,N_19177,N_19312);
xnor U20694 (N_20694,N_19931,N_19753);
nand U20695 (N_20695,N_19174,N_19066);
xor U20696 (N_20696,N_19384,N_19008);
and U20697 (N_20697,N_19740,N_19118);
nor U20698 (N_20698,N_19009,N_19282);
nand U20699 (N_20699,N_19024,N_19171);
nor U20700 (N_20700,N_19660,N_19777);
nand U20701 (N_20701,N_19566,N_19434);
nor U20702 (N_20702,N_19225,N_19550);
nor U20703 (N_20703,N_19175,N_19199);
and U20704 (N_20704,N_19602,N_19440);
nor U20705 (N_20705,N_19989,N_19040);
nand U20706 (N_20706,N_19957,N_19091);
nand U20707 (N_20707,N_19248,N_19509);
nor U20708 (N_20708,N_19529,N_19345);
nor U20709 (N_20709,N_19294,N_19837);
and U20710 (N_20710,N_19139,N_19660);
or U20711 (N_20711,N_19654,N_19601);
or U20712 (N_20712,N_19364,N_19602);
and U20713 (N_20713,N_19437,N_19224);
nand U20714 (N_20714,N_19178,N_19889);
nand U20715 (N_20715,N_19844,N_19402);
xnor U20716 (N_20716,N_19652,N_19318);
nor U20717 (N_20717,N_19852,N_19423);
xnor U20718 (N_20718,N_19840,N_19286);
or U20719 (N_20719,N_19607,N_19729);
nand U20720 (N_20720,N_19896,N_19220);
nor U20721 (N_20721,N_19762,N_19376);
or U20722 (N_20722,N_19313,N_19536);
nor U20723 (N_20723,N_19963,N_19371);
nand U20724 (N_20724,N_19478,N_19581);
or U20725 (N_20725,N_19203,N_19124);
nand U20726 (N_20726,N_19722,N_19924);
nor U20727 (N_20727,N_19540,N_19652);
and U20728 (N_20728,N_19538,N_19054);
nor U20729 (N_20729,N_19263,N_19956);
xor U20730 (N_20730,N_19611,N_19361);
xor U20731 (N_20731,N_19582,N_19624);
nand U20732 (N_20732,N_19638,N_19545);
or U20733 (N_20733,N_19128,N_19701);
nor U20734 (N_20734,N_19428,N_19918);
nand U20735 (N_20735,N_19547,N_19862);
or U20736 (N_20736,N_19861,N_19539);
xor U20737 (N_20737,N_19932,N_19736);
nor U20738 (N_20738,N_19458,N_19979);
xnor U20739 (N_20739,N_19936,N_19519);
or U20740 (N_20740,N_19170,N_19626);
or U20741 (N_20741,N_19542,N_19556);
nor U20742 (N_20742,N_19900,N_19776);
xnor U20743 (N_20743,N_19811,N_19897);
nor U20744 (N_20744,N_19616,N_19428);
xor U20745 (N_20745,N_19408,N_19743);
or U20746 (N_20746,N_19510,N_19774);
nand U20747 (N_20747,N_19243,N_19482);
xnor U20748 (N_20748,N_19022,N_19675);
nor U20749 (N_20749,N_19773,N_19150);
nand U20750 (N_20750,N_19298,N_19342);
and U20751 (N_20751,N_19695,N_19124);
or U20752 (N_20752,N_19599,N_19320);
nor U20753 (N_20753,N_19400,N_19637);
nand U20754 (N_20754,N_19844,N_19206);
and U20755 (N_20755,N_19625,N_19952);
nor U20756 (N_20756,N_19796,N_19528);
nand U20757 (N_20757,N_19657,N_19914);
nand U20758 (N_20758,N_19559,N_19306);
and U20759 (N_20759,N_19888,N_19162);
xor U20760 (N_20760,N_19111,N_19883);
or U20761 (N_20761,N_19200,N_19127);
or U20762 (N_20762,N_19717,N_19415);
xnor U20763 (N_20763,N_19976,N_19484);
nor U20764 (N_20764,N_19280,N_19235);
and U20765 (N_20765,N_19903,N_19601);
nor U20766 (N_20766,N_19753,N_19923);
nand U20767 (N_20767,N_19849,N_19167);
nand U20768 (N_20768,N_19562,N_19169);
xnor U20769 (N_20769,N_19085,N_19289);
xor U20770 (N_20770,N_19193,N_19744);
xnor U20771 (N_20771,N_19015,N_19825);
and U20772 (N_20772,N_19021,N_19591);
and U20773 (N_20773,N_19113,N_19815);
nand U20774 (N_20774,N_19818,N_19121);
or U20775 (N_20775,N_19383,N_19039);
or U20776 (N_20776,N_19860,N_19594);
and U20777 (N_20777,N_19867,N_19530);
or U20778 (N_20778,N_19948,N_19275);
nand U20779 (N_20779,N_19535,N_19571);
nor U20780 (N_20780,N_19764,N_19603);
xnor U20781 (N_20781,N_19072,N_19915);
and U20782 (N_20782,N_19937,N_19322);
or U20783 (N_20783,N_19260,N_19107);
nand U20784 (N_20784,N_19706,N_19484);
and U20785 (N_20785,N_19853,N_19554);
or U20786 (N_20786,N_19087,N_19824);
or U20787 (N_20787,N_19631,N_19661);
and U20788 (N_20788,N_19080,N_19935);
nand U20789 (N_20789,N_19284,N_19203);
nand U20790 (N_20790,N_19070,N_19346);
and U20791 (N_20791,N_19005,N_19587);
xor U20792 (N_20792,N_19536,N_19075);
nor U20793 (N_20793,N_19936,N_19351);
xnor U20794 (N_20794,N_19388,N_19439);
or U20795 (N_20795,N_19162,N_19911);
nand U20796 (N_20796,N_19620,N_19846);
and U20797 (N_20797,N_19698,N_19392);
or U20798 (N_20798,N_19083,N_19877);
nor U20799 (N_20799,N_19825,N_19575);
xnor U20800 (N_20800,N_19412,N_19235);
and U20801 (N_20801,N_19604,N_19394);
or U20802 (N_20802,N_19968,N_19734);
xor U20803 (N_20803,N_19004,N_19493);
nand U20804 (N_20804,N_19181,N_19310);
nand U20805 (N_20805,N_19459,N_19904);
or U20806 (N_20806,N_19378,N_19842);
and U20807 (N_20807,N_19122,N_19572);
nor U20808 (N_20808,N_19768,N_19282);
xor U20809 (N_20809,N_19211,N_19183);
xnor U20810 (N_20810,N_19126,N_19537);
nand U20811 (N_20811,N_19567,N_19823);
and U20812 (N_20812,N_19990,N_19158);
or U20813 (N_20813,N_19196,N_19447);
nor U20814 (N_20814,N_19701,N_19385);
nand U20815 (N_20815,N_19575,N_19614);
xnor U20816 (N_20816,N_19891,N_19434);
or U20817 (N_20817,N_19931,N_19030);
or U20818 (N_20818,N_19418,N_19747);
xor U20819 (N_20819,N_19834,N_19719);
or U20820 (N_20820,N_19222,N_19771);
nand U20821 (N_20821,N_19073,N_19132);
and U20822 (N_20822,N_19298,N_19131);
and U20823 (N_20823,N_19427,N_19941);
or U20824 (N_20824,N_19531,N_19061);
nor U20825 (N_20825,N_19050,N_19044);
nand U20826 (N_20826,N_19953,N_19194);
nand U20827 (N_20827,N_19323,N_19451);
nor U20828 (N_20828,N_19864,N_19671);
or U20829 (N_20829,N_19471,N_19485);
or U20830 (N_20830,N_19988,N_19151);
xor U20831 (N_20831,N_19409,N_19570);
xor U20832 (N_20832,N_19730,N_19759);
or U20833 (N_20833,N_19919,N_19395);
nor U20834 (N_20834,N_19933,N_19405);
nor U20835 (N_20835,N_19923,N_19160);
xor U20836 (N_20836,N_19923,N_19770);
nor U20837 (N_20837,N_19193,N_19415);
nor U20838 (N_20838,N_19938,N_19867);
xnor U20839 (N_20839,N_19693,N_19084);
or U20840 (N_20840,N_19201,N_19136);
xor U20841 (N_20841,N_19206,N_19748);
xor U20842 (N_20842,N_19158,N_19938);
or U20843 (N_20843,N_19642,N_19606);
xnor U20844 (N_20844,N_19280,N_19472);
nand U20845 (N_20845,N_19269,N_19109);
or U20846 (N_20846,N_19548,N_19097);
xor U20847 (N_20847,N_19483,N_19238);
or U20848 (N_20848,N_19850,N_19318);
xnor U20849 (N_20849,N_19155,N_19307);
or U20850 (N_20850,N_19882,N_19136);
nand U20851 (N_20851,N_19163,N_19773);
nor U20852 (N_20852,N_19125,N_19976);
or U20853 (N_20853,N_19370,N_19466);
nor U20854 (N_20854,N_19812,N_19581);
and U20855 (N_20855,N_19250,N_19958);
nand U20856 (N_20856,N_19092,N_19484);
and U20857 (N_20857,N_19536,N_19364);
nor U20858 (N_20858,N_19235,N_19975);
xnor U20859 (N_20859,N_19096,N_19493);
and U20860 (N_20860,N_19884,N_19798);
and U20861 (N_20861,N_19736,N_19848);
xor U20862 (N_20862,N_19692,N_19849);
nor U20863 (N_20863,N_19624,N_19419);
nor U20864 (N_20864,N_19787,N_19181);
xnor U20865 (N_20865,N_19033,N_19694);
or U20866 (N_20866,N_19193,N_19365);
nor U20867 (N_20867,N_19233,N_19273);
xnor U20868 (N_20868,N_19561,N_19368);
or U20869 (N_20869,N_19275,N_19914);
or U20870 (N_20870,N_19833,N_19872);
nand U20871 (N_20871,N_19278,N_19794);
or U20872 (N_20872,N_19503,N_19237);
nor U20873 (N_20873,N_19566,N_19593);
or U20874 (N_20874,N_19677,N_19171);
or U20875 (N_20875,N_19398,N_19772);
xor U20876 (N_20876,N_19785,N_19236);
and U20877 (N_20877,N_19864,N_19210);
nand U20878 (N_20878,N_19807,N_19257);
or U20879 (N_20879,N_19950,N_19140);
or U20880 (N_20880,N_19090,N_19911);
and U20881 (N_20881,N_19040,N_19956);
nand U20882 (N_20882,N_19038,N_19125);
and U20883 (N_20883,N_19846,N_19455);
or U20884 (N_20884,N_19065,N_19636);
nor U20885 (N_20885,N_19143,N_19312);
and U20886 (N_20886,N_19179,N_19374);
and U20887 (N_20887,N_19712,N_19664);
nand U20888 (N_20888,N_19852,N_19245);
and U20889 (N_20889,N_19808,N_19441);
nor U20890 (N_20890,N_19266,N_19681);
or U20891 (N_20891,N_19257,N_19612);
nand U20892 (N_20892,N_19954,N_19360);
nand U20893 (N_20893,N_19245,N_19826);
xor U20894 (N_20894,N_19133,N_19585);
and U20895 (N_20895,N_19168,N_19554);
or U20896 (N_20896,N_19869,N_19215);
or U20897 (N_20897,N_19045,N_19546);
and U20898 (N_20898,N_19447,N_19806);
xnor U20899 (N_20899,N_19109,N_19900);
nand U20900 (N_20900,N_19923,N_19519);
nor U20901 (N_20901,N_19651,N_19966);
nor U20902 (N_20902,N_19730,N_19641);
or U20903 (N_20903,N_19205,N_19080);
nor U20904 (N_20904,N_19117,N_19751);
xor U20905 (N_20905,N_19683,N_19369);
and U20906 (N_20906,N_19323,N_19487);
nand U20907 (N_20907,N_19861,N_19374);
nand U20908 (N_20908,N_19508,N_19583);
xnor U20909 (N_20909,N_19032,N_19072);
or U20910 (N_20910,N_19423,N_19581);
and U20911 (N_20911,N_19537,N_19682);
nand U20912 (N_20912,N_19559,N_19725);
and U20913 (N_20913,N_19813,N_19812);
nor U20914 (N_20914,N_19286,N_19859);
and U20915 (N_20915,N_19739,N_19037);
or U20916 (N_20916,N_19964,N_19907);
and U20917 (N_20917,N_19095,N_19577);
or U20918 (N_20918,N_19794,N_19979);
nor U20919 (N_20919,N_19508,N_19734);
nand U20920 (N_20920,N_19664,N_19846);
nor U20921 (N_20921,N_19905,N_19052);
xnor U20922 (N_20922,N_19559,N_19677);
xor U20923 (N_20923,N_19886,N_19656);
and U20924 (N_20924,N_19390,N_19928);
nor U20925 (N_20925,N_19373,N_19996);
nand U20926 (N_20926,N_19868,N_19903);
nor U20927 (N_20927,N_19704,N_19566);
xor U20928 (N_20928,N_19471,N_19713);
nand U20929 (N_20929,N_19564,N_19597);
xor U20930 (N_20930,N_19965,N_19700);
or U20931 (N_20931,N_19174,N_19927);
and U20932 (N_20932,N_19317,N_19422);
or U20933 (N_20933,N_19282,N_19546);
nor U20934 (N_20934,N_19034,N_19805);
nand U20935 (N_20935,N_19971,N_19063);
nor U20936 (N_20936,N_19541,N_19326);
xnor U20937 (N_20937,N_19192,N_19410);
nand U20938 (N_20938,N_19942,N_19642);
and U20939 (N_20939,N_19507,N_19493);
or U20940 (N_20940,N_19169,N_19333);
nor U20941 (N_20941,N_19139,N_19051);
nor U20942 (N_20942,N_19886,N_19489);
xor U20943 (N_20943,N_19522,N_19220);
nand U20944 (N_20944,N_19754,N_19778);
and U20945 (N_20945,N_19053,N_19848);
xnor U20946 (N_20946,N_19899,N_19995);
nand U20947 (N_20947,N_19600,N_19423);
nand U20948 (N_20948,N_19390,N_19116);
or U20949 (N_20949,N_19259,N_19094);
or U20950 (N_20950,N_19283,N_19906);
and U20951 (N_20951,N_19684,N_19085);
or U20952 (N_20952,N_19633,N_19439);
and U20953 (N_20953,N_19538,N_19164);
nor U20954 (N_20954,N_19898,N_19664);
and U20955 (N_20955,N_19675,N_19419);
nand U20956 (N_20956,N_19854,N_19831);
xnor U20957 (N_20957,N_19018,N_19478);
or U20958 (N_20958,N_19133,N_19505);
nand U20959 (N_20959,N_19011,N_19689);
nand U20960 (N_20960,N_19317,N_19367);
nor U20961 (N_20961,N_19182,N_19013);
and U20962 (N_20962,N_19603,N_19950);
xor U20963 (N_20963,N_19285,N_19274);
and U20964 (N_20964,N_19838,N_19973);
nor U20965 (N_20965,N_19387,N_19068);
or U20966 (N_20966,N_19888,N_19789);
nor U20967 (N_20967,N_19183,N_19693);
xnor U20968 (N_20968,N_19091,N_19848);
nor U20969 (N_20969,N_19579,N_19545);
nor U20970 (N_20970,N_19649,N_19844);
xnor U20971 (N_20971,N_19600,N_19553);
xor U20972 (N_20972,N_19849,N_19058);
or U20973 (N_20973,N_19206,N_19441);
nand U20974 (N_20974,N_19554,N_19355);
or U20975 (N_20975,N_19671,N_19272);
nor U20976 (N_20976,N_19077,N_19135);
nand U20977 (N_20977,N_19851,N_19868);
and U20978 (N_20978,N_19493,N_19485);
nand U20979 (N_20979,N_19414,N_19587);
xnor U20980 (N_20980,N_19052,N_19678);
nor U20981 (N_20981,N_19894,N_19644);
or U20982 (N_20982,N_19016,N_19018);
or U20983 (N_20983,N_19195,N_19703);
or U20984 (N_20984,N_19542,N_19283);
and U20985 (N_20985,N_19631,N_19410);
or U20986 (N_20986,N_19331,N_19909);
and U20987 (N_20987,N_19875,N_19601);
and U20988 (N_20988,N_19315,N_19109);
nand U20989 (N_20989,N_19520,N_19672);
nor U20990 (N_20990,N_19355,N_19225);
xnor U20991 (N_20991,N_19048,N_19811);
or U20992 (N_20992,N_19802,N_19892);
or U20993 (N_20993,N_19763,N_19971);
xnor U20994 (N_20994,N_19244,N_19280);
and U20995 (N_20995,N_19085,N_19408);
nand U20996 (N_20996,N_19207,N_19066);
or U20997 (N_20997,N_19499,N_19044);
and U20998 (N_20998,N_19982,N_19081);
or U20999 (N_20999,N_19418,N_19518);
and U21000 (N_21000,N_20995,N_20024);
xor U21001 (N_21001,N_20095,N_20101);
nor U21002 (N_21002,N_20984,N_20944);
nand U21003 (N_21003,N_20505,N_20950);
and U21004 (N_21004,N_20406,N_20844);
xor U21005 (N_21005,N_20362,N_20068);
xor U21006 (N_21006,N_20412,N_20263);
xnor U21007 (N_21007,N_20926,N_20635);
or U21008 (N_21008,N_20139,N_20616);
nor U21009 (N_21009,N_20979,N_20887);
xor U21010 (N_21010,N_20792,N_20879);
nand U21011 (N_21011,N_20389,N_20876);
nand U21012 (N_21012,N_20873,N_20728);
and U21013 (N_21013,N_20367,N_20173);
nand U21014 (N_21014,N_20503,N_20532);
or U21015 (N_21015,N_20742,N_20575);
and U21016 (N_21016,N_20752,N_20289);
xor U21017 (N_21017,N_20819,N_20768);
nand U21018 (N_21018,N_20494,N_20699);
nor U21019 (N_21019,N_20499,N_20996);
or U21020 (N_21020,N_20674,N_20772);
or U21021 (N_21021,N_20708,N_20871);
and U21022 (N_21022,N_20609,N_20080);
xor U21023 (N_21023,N_20200,N_20901);
and U21024 (N_21024,N_20211,N_20798);
nor U21025 (N_21025,N_20345,N_20631);
xnor U21026 (N_21026,N_20031,N_20084);
xnor U21027 (N_21027,N_20540,N_20223);
nor U21028 (N_21028,N_20981,N_20037);
xor U21029 (N_21029,N_20148,N_20859);
xnor U21030 (N_21030,N_20727,N_20565);
or U21031 (N_21031,N_20733,N_20191);
nor U21032 (N_21032,N_20543,N_20629);
and U21033 (N_21033,N_20707,N_20066);
and U21034 (N_21034,N_20920,N_20709);
and U21035 (N_21035,N_20022,N_20212);
or U21036 (N_21036,N_20482,N_20620);
nor U21037 (N_21037,N_20777,N_20647);
nand U21038 (N_21038,N_20663,N_20884);
and U21039 (N_21039,N_20098,N_20292);
nor U21040 (N_21040,N_20423,N_20824);
or U21041 (N_21041,N_20590,N_20257);
and U21042 (N_21042,N_20308,N_20176);
xnor U21043 (N_21043,N_20868,N_20195);
and U21044 (N_21044,N_20679,N_20854);
nor U21045 (N_21045,N_20045,N_20097);
or U21046 (N_21046,N_20099,N_20630);
and U21047 (N_21047,N_20608,N_20856);
nand U21048 (N_21048,N_20254,N_20365);
nor U21049 (N_21049,N_20640,N_20120);
xnor U21050 (N_21050,N_20786,N_20973);
and U21051 (N_21051,N_20426,N_20430);
and U21052 (N_21052,N_20581,N_20658);
nor U21053 (N_21053,N_20071,N_20875);
or U21054 (N_21054,N_20256,N_20619);
or U21055 (N_21055,N_20463,N_20048);
xnor U21056 (N_21056,N_20160,N_20753);
nor U21057 (N_21057,N_20162,N_20906);
xor U21058 (N_21058,N_20260,N_20056);
xnor U21059 (N_21059,N_20034,N_20246);
and U21060 (N_21060,N_20409,N_20520);
xnor U21061 (N_21061,N_20783,N_20407);
or U21062 (N_21062,N_20054,N_20703);
xor U21063 (N_21063,N_20963,N_20821);
nor U21064 (N_21064,N_20478,N_20541);
and U21065 (N_21065,N_20285,N_20327);
xor U21066 (N_21066,N_20044,N_20381);
nor U21067 (N_21067,N_20485,N_20416);
nor U21068 (N_21068,N_20003,N_20736);
nand U21069 (N_21069,N_20392,N_20317);
xor U21070 (N_21070,N_20228,N_20053);
or U21071 (N_21071,N_20323,N_20118);
xnor U21072 (N_21072,N_20998,N_20002);
xor U21073 (N_21073,N_20686,N_20559);
xor U21074 (N_21074,N_20291,N_20437);
and U21075 (N_21075,N_20239,N_20539);
or U21076 (N_21076,N_20304,N_20060);
nor U21077 (N_21077,N_20483,N_20496);
xor U21078 (N_21078,N_20976,N_20756);
xor U21079 (N_21079,N_20431,N_20073);
and U21080 (N_21080,N_20508,N_20602);
or U21081 (N_21081,N_20556,N_20125);
nand U21082 (N_21082,N_20848,N_20069);
nand U21083 (N_21083,N_20150,N_20174);
or U21084 (N_21084,N_20070,N_20550);
xor U21085 (N_21085,N_20332,N_20372);
nor U21086 (N_21086,N_20899,N_20420);
or U21087 (N_21087,N_20701,N_20645);
nor U21088 (N_21088,N_20447,N_20954);
nand U21089 (N_21089,N_20529,N_20270);
or U21090 (N_21090,N_20385,N_20921);
or U21091 (N_21091,N_20010,N_20877);
nor U21092 (N_21092,N_20583,N_20846);
and U21093 (N_21093,N_20769,N_20524);
nand U21094 (N_21094,N_20839,N_20997);
and U21095 (N_21095,N_20103,N_20595);
or U21096 (N_21096,N_20900,N_20810);
nand U21097 (N_21097,N_20438,N_20458);
nand U21098 (N_21098,N_20672,N_20049);
nand U21099 (N_21099,N_20725,N_20428);
or U21100 (N_21100,N_20591,N_20775);
nor U21101 (N_21101,N_20123,N_20082);
or U21102 (N_21102,N_20453,N_20171);
nor U21103 (N_21103,N_20641,N_20449);
and U21104 (N_21104,N_20882,N_20700);
nand U21105 (N_21105,N_20692,N_20273);
xnor U21106 (N_21106,N_20513,N_20491);
nor U21107 (N_21107,N_20925,N_20305);
or U21108 (N_21108,N_20587,N_20660);
and U21109 (N_21109,N_20360,N_20787);
and U21110 (N_21110,N_20857,N_20489);
or U21111 (N_21111,N_20353,N_20811);
nand U21112 (N_21112,N_20419,N_20612);
xnor U21113 (N_21113,N_20497,N_20653);
and U21114 (N_21114,N_20924,N_20953);
xnor U21115 (N_21115,N_20432,N_20959);
or U21116 (N_21116,N_20578,N_20555);
xor U21117 (N_21117,N_20898,N_20495);
nand U21118 (N_21118,N_20795,N_20737);
nor U21119 (N_21119,N_20347,N_20939);
or U21120 (N_21120,N_20274,N_20521);
nor U21121 (N_21121,N_20828,N_20001);
and U21122 (N_21122,N_20455,N_20450);
nor U21123 (N_21123,N_20134,N_20492);
nor U21124 (N_21124,N_20376,N_20033);
xnor U21125 (N_21125,N_20655,N_20067);
nor U21126 (N_21126,N_20029,N_20570);
nand U21127 (N_21127,N_20751,N_20517);
and U21128 (N_21128,N_20904,N_20040);
nand U21129 (N_21129,N_20009,N_20624);
xor U21130 (N_21130,N_20262,N_20222);
and U21131 (N_21131,N_20356,N_20185);
or U21132 (N_21132,N_20688,N_20301);
xnor U21133 (N_21133,N_20276,N_20471);
and U21134 (N_21134,N_20454,N_20863);
xor U21135 (N_21135,N_20827,N_20712);
xor U21136 (N_21136,N_20955,N_20664);
and U21137 (N_21137,N_20476,N_20579);
xnor U21138 (N_21138,N_20902,N_20149);
nand U21139 (N_21139,N_20395,N_20116);
xor U21140 (N_21140,N_20794,N_20272);
xnor U21141 (N_21141,N_20018,N_20357);
or U21142 (N_21142,N_20364,N_20597);
or U21143 (N_21143,N_20142,N_20962);
nor U21144 (N_21144,N_20853,N_20271);
or U21145 (N_21145,N_20467,N_20219);
nand U21146 (N_21146,N_20187,N_20415);
and U21147 (N_21147,N_20448,N_20157);
and U21148 (N_21148,N_20322,N_20724);
or U21149 (N_21149,N_20596,N_20178);
nor U21150 (N_21150,N_20404,N_20094);
xnor U21151 (N_21151,N_20108,N_20295);
nand U21152 (N_21152,N_20141,N_20030);
or U21153 (N_21153,N_20580,N_20417);
xnor U21154 (N_21154,N_20917,N_20860);
and U21155 (N_21155,N_20527,N_20711);
and U21156 (N_21156,N_20506,N_20636);
nand U21157 (N_21157,N_20368,N_20915);
and U21158 (N_21158,N_20177,N_20610);
or U21159 (N_21159,N_20230,N_20340);
nand U21160 (N_21160,N_20991,N_20622);
nand U21161 (N_21161,N_20850,N_20032);
xnor U21162 (N_21162,N_20716,N_20577);
and U21163 (N_21163,N_20440,N_20883);
nand U21164 (N_21164,N_20460,N_20279);
nor U21165 (N_21165,N_20302,N_20243);
nand U21166 (N_21166,N_20960,N_20153);
nor U21167 (N_21167,N_20748,N_20969);
nor U21168 (N_21168,N_20800,N_20321);
nor U21169 (N_21169,N_20885,N_20965);
nand U21170 (N_21170,N_20199,N_20628);
xor U21171 (N_21171,N_20210,N_20808);
or U21172 (N_21172,N_20779,N_20994);
xnor U21173 (N_21173,N_20764,N_20568);
nor U21174 (N_21174,N_20516,N_20375);
and U21175 (N_21175,N_20715,N_20490);
and U21176 (N_21176,N_20832,N_20281);
or U21177 (N_21177,N_20966,N_20078);
or U21178 (N_21178,N_20649,N_20967);
and U21179 (N_21179,N_20909,N_20232);
nand U21180 (N_21180,N_20740,N_20008);
and U21181 (N_21181,N_20350,N_20484);
nand U21182 (N_21182,N_20685,N_20754);
nand U21183 (N_21183,N_20651,N_20296);
nand U21184 (N_21184,N_20086,N_20538);
and U21185 (N_21185,N_20788,N_20470);
nand U21186 (N_21186,N_20830,N_20181);
nand U21187 (N_21187,N_20689,N_20734);
xor U21188 (N_21188,N_20702,N_20136);
or U21189 (N_21189,N_20836,N_20923);
nor U21190 (N_21190,N_20359,N_20479);
nand U21191 (N_21191,N_20698,N_20179);
nand U21192 (N_21192,N_20598,N_20789);
xor U21193 (N_21193,N_20571,N_20462);
nor U21194 (N_21194,N_20897,N_20207);
nand U21195 (N_21195,N_20025,N_20773);
or U21196 (N_21196,N_20722,N_20079);
xnor U21197 (N_21197,N_20584,N_20235);
and U21198 (N_21198,N_20093,N_20393);
nand U21199 (N_21199,N_20718,N_20983);
nor U21200 (N_21200,N_20601,N_20849);
nor U21201 (N_21201,N_20215,N_20766);
nand U21202 (N_21202,N_20000,N_20820);
or U21203 (N_21203,N_20390,N_20554);
and U21204 (N_21204,N_20047,N_20076);
or U21205 (N_21205,N_20300,N_20697);
xor U21206 (N_21206,N_20803,N_20158);
xor U21207 (N_21207,N_20444,N_20064);
nand U21208 (N_21208,N_20822,N_20439);
or U21209 (N_21209,N_20843,N_20189);
nor U21210 (N_21210,N_20102,N_20170);
nand U21211 (N_21211,N_20977,N_20972);
or U21212 (N_21212,N_20642,N_20361);
nand U21213 (N_21213,N_20293,N_20714);
nor U21214 (N_21214,N_20442,N_20964);
nor U21215 (N_21215,N_20472,N_20613);
nand U21216 (N_21216,N_20233,N_20269);
or U21217 (N_21217,N_20133,N_20004);
xor U21218 (N_21218,N_20312,N_20840);
or U21219 (N_21219,N_20077,N_20156);
or U21220 (N_21220,N_20227,N_20203);
nand U21221 (N_21221,N_20441,N_20760);
nor U21222 (N_21222,N_20366,N_20804);
and U21223 (N_21223,N_20988,N_20937);
and U21224 (N_21224,N_20932,N_20880);
xor U21225 (N_21225,N_20121,N_20085);
and U21226 (N_21226,N_20414,N_20287);
nor U21227 (N_21227,N_20138,N_20011);
or U21228 (N_21228,N_20041,N_20913);
xor U21229 (N_21229,N_20140,N_20346);
or U21230 (N_21230,N_20425,N_20706);
nor U21231 (N_21231,N_20949,N_20561);
nor U21232 (N_21232,N_20255,N_20643);
or U21233 (N_21233,N_20072,N_20695);
nor U21234 (N_21234,N_20750,N_20947);
nand U21235 (N_21235,N_20528,N_20413);
xnor U21236 (N_21236,N_20738,N_20801);
or U21237 (N_21237,N_20050,N_20562);
nor U21238 (N_21238,N_20500,N_20113);
and U21239 (N_21239,N_20745,N_20147);
nor U21240 (N_21240,N_20268,N_20433);
nand U21241 (N_21241,N_20758,N_20992);
and U21242 (N_21242,N_20242,N_20874);
nor U21243 (N_21243,N_20684,N_20411);
or U21244 (N_21244,N_20693,N_20192);
nand U21245 (N_21245,N_20184,N_20265);
or U21246 (N_21246,N_20014,N_20945);
xnor U21247 (N_21247,N_20280,N_20878);
xor U21248 (N_21248,N_20644,N_20240);
or U21249 (N_21249,N_20530,N_20143);
xnor U21250 (N_21250,N_20946,N_20297);
or U21251 (N_21251,N_20968,N_20107);
nand U21252 (N_21252,N_20343,N_20020);
nor U21253 (N_21253,N_20809,N_20126);
xor U21254 (N_21254,N_20152,N_20015);
nor U21255 (N_21255,N_20905,N_20858);
xnor U21256 (N_21256,N_20586,N_20594);
and U21257 (N_21257,N_20687,N_20721);
nor U21258 (N_21258,N_20719,N_20933);
xor U21259 (N_21259,N_20615,N_20109);
nor U21260 (N_21260,N_20936,N_20007);
nor U21261 (N_21261,N_20388,N_20816);
nand U21262 (N_21262,N_20951,N_20511);
and U21263 (N_21263,N_20535,N_20665);
and U21264 (N_21264,N_20916,N_20910);
nand U21265 (N_21265,N_20006,N_20564);
nand U21266 (N_21266,N_20614,N_20035);
nor U21267 (N_21267,N_20993,N_20646);
and U21268 (N_21268,N_20891,N_20852);
nand U21269 (N_21269,N_20893,N_20104);
nor U21270 (N_21270,N_20275,N_20331);
and U21271 (N_21271,N_20851,N_20551);
xnor U21272 (N_21272,N_20167,N_20611);
or U21273 (N_21273,N_20755,N_20978);
nor U21274 (N_21274,N_20743,N_20894);
and U21275 (N_21275,N_20791,N_20386);
nor U21276 (N_21276,N_20668,N_20400);
nor U21277 (N_21277,N_20514,N_20299);
nand U21278 (N_21278,N_20650,N_20785);
and U21279 (N_21279,N_20197,N_20046);
nor U21280 (N_21280,N_20573,N_20833);
nand U21281 (N_21281,N_20328,N_20481);
or U21282 (N_21282,N_20501,N_20717);
nor U21283 (N_21283,N_20021,N_20401);
or U21284 (N_21284,N_20464,N_20398);
xnor U21285 (N_21285,N_20468,N_20825);
xnor U21286 (N_21286,N_20831,N_20166);
nor U21287 (N_21287,N_20106,N_20216);
nand U21288 (N_21288,N_20911,N_20339);
nand U21289 (N_21289,N_20341,N_20731);
nand U21290 (N_21290,N_20866,N_20294);
nand U21291 (N_21291,N_20213,N_20761);
or U21292 (N_21292,N_20480,N_20934);
and U21293 (N_21293,N_20155,N_20576);
nand U21294 (N_21294,N_20572,N_20253);
nand U21295 (N_21295,N_20566,N_20971);
xor U21296 (N_21296,N_20394,N_20247);
nor U21297 (N_21297,N_20436,N_20445);
nand U21298 (N_21298,N_20100,N_20582);
and U21299 (N_21299,N_20473,N_20016);
xnor U21300 (N_21300,N_20313,N_20888);
or U21301 (N_21301,N_20694,N_20889);
and U21302 (N_21302,N_20316,N_20829);
or U21303 (N_21303,N_20338,N_20418);
and U21304 (N_21304,N_20678,N_20310);
nand U21305 (N_21305,N_20762,N_20986);
and U21306 (N_21306,N_20110,N_20378);
and U21307 (N_21307,N_20261,N_20793);
or U21308 (N_21308,N_20704,N_20330);
xor U21309 (N_21309,N_20111,N_20606);
nor U21310 (N_21310,N_20026,N_20796);
nand U21311 (N_21311,N_20845,N_20051);
and U21312 (N_21312,N_20600,N_20373);
xnor U21313 (N_21313,N_20574,N_20329);
or U21314 (N_21314,N_20286,N_20324);
nor U21315 (N_21315,N_20690,N_20318);
nor U21316 (N_21316,N_20661,N_20380);
nor U21317 (N_21317,N_20282,N_20402);
xor U21318 (N_21318,N_20774,N_20488);
xnor U21319 (N_21319,N_20465,N_20927);
and U21320 (N_21320,N_20446,N_20487);
or U21321 (N_21321,N_20940,N_20999);
xnor U21322 (N_21322,N_20930,N_20818);
or U21323 (N_21323,N_20421,N_20918);
xnor U21324 (N_21324,N_20218,N_20258);
or U21325 (N_21325,N_20352,N_20019);
and U21326 (N_21326,N_20982,N_20855);
and U21327 (N_21327,N_20870,N_20370);
and U21328 (N_21328,N_20985,N_20790);
xnor U21329 (N_21329,N_20941,N_20558);
or U21330 (N_21330,N_20677,N_20135);
nand U21331 (N_21331,N_20283,N_20563);
or U21332 (N_21332,N_20165,N_20974);
or U21333 (N_21333,N_20422,N_20290);
nand U21334 (N_21334,N_20128,N_20542);
nor U21335 (N_21335,N_20089,N_20334);
nand U21336 (N_21336,N_20059,N_20039);
and U21337 (N_21337,N_20063,N_20427);
nand U21338 (N_21338,N_20956,N_20259);
nor U21339 (N_21339,N_20990,N_20342);
nand U21340 (N_21340,N_20815,N_20112);
nand U21341 (N_21341,N_20593,N_20604);
xor U21342 (N_21342,N_20209,N_20236);
and U21343 (N_21343,N_20675,N_20132);
nand U21344 (N_21344,N_20137,N_20383);
and U21345 (N_21345,N_20131,N_20919);
and U21346 (N_21346,N_20410,N_20735);
nand U21347 (N_21347,N_20780,N_20812);
nor U21348 (N_21348,N_20266,N_20961);
nand U21349 (N_21349,N_20943,N_20518);
xor U21350 (N_21350,N_20314,N_20226);
or U21351 (N_21351,N_20869,N_20249);
xor U21352 (N_21352,N_20841,N_20217);
xnor U21353 (N_21353,N_20348,N_20129);
nor U21354 (N_21354,N_20623,N_20127);
or U21355 (N_21355,N_20847,N_20895);
and U21356 (N_21356,N_20507,N_20544);
nor U21357 (N_21357,N_20303,N_20408);
or U21358 (N_21358,N_20214,N_20119);
nor U21359 (N_21359,N_20377,N_20807);
xor U21360 (N_21360,N_20028,N_20669);
nand U21361 (N_21361,N_20928,N_20512);
xor U21362 (N_21362,N_20241,N_20929);
xor U21363 (N_21363,N_20767,N_20146);
nor U21364 (N_21364,N_20519,N_20813);
nor U21365 (N_21365,N_20403,N_20405);
xnor U21366 (N_21366,N_20567,N_20667);
nand U21367 (N_21367,N_20553,N_20835);
nor U21368 (N_21368,N_20662,N_20161);
or U21369 (N_21369,N_20429,N_20522);
nor U21370 (N_21370,N_20585,N_20552);
nand U21371 (N_21371,N_20201,N_20509);
nor U21372 (N_21372,N_20639,N_20309);
nor U21373 (N_21373,N_20526,N_20091);
and U21374 (N_21374,N_20952,N_20164);
nor U21375 (N_21375,N_20806,N_20837);
nor U21376 (N_21376,N_20151,N_20369);
and U21377 (N_21377,N_20115,N_20194);
and U21378 (N_21378,N_20523,N_20204);
or U21379 (N_21379,N_20681,N_20797);
nand U21380 (N_21380,N_20475,N_20379);
and U21381 (N_21381,N_20670,N_20435);
or U21382 (N_21382,N_20802,N_20560);
xor U21383 (N_21383,N_20907,N_20117);
xor U21384 (N_21384,N_20391,N_20676);
xor U21385 (N_21385,N_20912,N_20358);
and U21386 (N_21386,N_20778,N_20278);
xor U21387 (N_21387,N_20671,N_20648);
or U21388 (N_21388,N_20654,N_20055);
nand U21389 (N_21389,N_20746,N_20443);
nand U21390 (N_21390,N_20163,N_20335);
xor U21391 (N_21391,N_20105,N_20466);
nand U21392 (N_21392,N_20531,N_20186);
or U21393 (N_21393,N_20224,N_20231);
nor U21394 (N_21394,N_20970,N_20618);
xor U21395 (N_21395,N_20144,N_20680);
xnor U21396 (N_21396,N_20548,N_20225);
nand U21397 (N_21397,N_20975,N_20159);
xnor U21398 (N_21398,N_20720,N_20605);
or U21399 (N_21399,N_20634,N_20154);
nand U21400 (N_21400,N_20682,N_20145);
nand U21401 (N_21401,N_20267,N_20625);
nor U21402 (N_21402,N_20938,N_20457);
xor U21403 (N_21403,N_20190,N_20862);
nor U21404 (N_21404,N_20890,N_20931);
nand U21405 (N_21405,N_20763,N_20599);
or U21406 (N_21406,N_20245,N_20881);
or U21407 (N_21407,N_20914,N_20626);
nor U21408 (N_21408,N_20896,N_20087);
nor U21409 (N_21409,N_20486,N_20182);
and U21410 (N_21410,N_20399,N_20012);
xor U21411 (N_21411,N_20298,N_20248);
or U21412 (N_21412,N_20549,N_20451);
xnor U21413 (N_21413,N_20065,N_20452);
xnor U21414 (N_21414,N_20234,N_20765);
nor U21415 (N_21415,N_20168,N_20739);
nor U21416 (N_21416,N_20705,N_20657);
nor U21417 (N_21417,N_20384,N_20935);
and U21418 (N_21418,N_20730,N_20319);
nand U21419 (N_21419,N_20244,N_20320);
xor U21420 (N_21420,N_20942,N_20823);
or U21421 (N_21421,N_20536,N_20683);
or U21422 (N_21422,N_20922,N_20502);
nor U21423 (N_21423,N_20723,N_20202);
xor U21424 (N_21424,N_20220,N_20781);
nor U21425 (N_21425,N_20336,N_20696);
nand U21426 (N_21426,N_20534,N_20776);
xor U21427 (N_21427,N_20504,N_20043);
xnor U21428 (N_21428,N_20396,N_20096);
xor U21429 (N_21429,N_20784,N_20987);
or U21430 (N_21430,N_20948,N_20886);
nand U21431 (N_21431,N_20017,N_20172);
and U21432 (N_21432,N_20713,N_20757);
or U21433 (N_21433,N_20122,N_20958);
and U21434 (N_21434,N_20741,N_20169);
nand U21435 (N_21435,N_20656,N_20759);
nand U21436 (N_21436,N_20074,N_20498);
and U21437 (N_21437,N_20817,N_20980);
nand U21438 (N_21438,N_20387,N_20229);
and U21439 (N_21439,N_20867,N_20782);
and U21440 (N_21440,N_20805,N_20838);
nand U21441 (N_21441,N_20371,N_20545);
or U21442 (N_21442,N_20592,N_20252);
nand U21443 (N_21443,N_20251,N_20627);
nor U21444 (N_21444,N_20603,N_20525);
and U21445 (N_21445,N_20354,N_20013);
or U21446 (N_21446,N_20193,N_20374);
and U21447 (N_21447,N_20659,N_20311);
and U21448 (N_21448,N_20363,N_20284);
xor U21449 (N_21449,N_20510,N_20732);
xnor U21450 (N_21450,N_20461,N_20351);
or U21451 (N_21451,N_20673,N_20196);
nor U21452 (N_21452,N_20264,N_20617);
nand U21453 (N_21453,N_20206,N_20005);
xor U21454 (N_21454,N_20075,N_20770);
or U21455 (N_21455,N_20198,N_20277);
and U21456 (N_21456,N_20057,N_20569);
or U21457 (N_21457,N_20175,N_20337);
and U21458 (N_21458,N_20188,N_20546);
or U21459 (N_21459,N_20092,N_20892);
nor U21460 (N_21460,N_20183,N_20633);
nand U21461 (N_21461,N_20771,N_20090);
or U21462 (N_21462,N_20749,N_20474);
xnor U21463 (N_21463,N_20691,N_20062);
or U21464 (N_21464,N_20180,N_20083);
nor U21465 (N_21465,N_20872,N_20250);
nand U21466 (N_21466,N_20221,N_20355);
xnor U21467 (N_21467,N_20038,N_20477);
or U21468 (N_21468,N_20747,N_20469);
nand U21469 (N_21469,N_20865,N_20088);
nor U21470 (N_21470,N_20842,N_20908);
and U21471 (N_21471,N_20114,N_20333);
or U21472 (N_21472,N_20632,N_20397);
nand U21473 (N_21473,N_20861,N_20058);
nor U21474 (N_21474,N_20382,N_20557);
xnor U21475 (N_21475,N_20238,N_20052);
xor U21476 (N_21476,N_20061,N_20124);
or U21477 (N_21477,N_20814,N_20607);
xor U21478 (N_21478,N_20710,N_20989);
xor U21479 (N_21479,N_20456,N_20864);
nand U21480 (N_21480,N_20027,N_20957);
nor U21481 (N_21481,N_20826,N_20325);
or U21482 (N_21482,N_20459,N_20515);
nand U21483 (N_21483,N_20547,N_20799);
and U21484 (N_21484,N_20493,N_20537);
and U21485 (N_21485,N_20023,N_20666);
nor U21486 (N_21486,N_20652,N_20729);
nor U21487 (N_21487,N_20638,N_20637);
xor U21488 (N_21488,N_20349,N_20288);
or U21489 (N_21489,N_20315,N_20726);
nor U21490 (N_21490,N_20208,N_20424);
nor U21491 (N_21491,N_20434,N_20130);
nor U21492 (N_21492,N_20205,N_20533);
nor U21493 (N_21493,N_20621,N_20081);
and U21494 (N_21494,N_20306,N_20903);
xnor U21495 (N_21495,N_20344,N_20307);
nor U21496 (N_21496,N_20588,N_20326);
nor U21497 (N_21497,N_20834,N_20036);
nand U21498 (N_21498,N_20237,N_20042);
xnor U21499 (N_21499,N_20744,N_20589);
and U21500 (N_21500,N_20864,N_20618);
nand U21501 (N_21501,N_20680,N_20879);
nand U21502 (N_21502,N_20507,N_20370);
or U21503 (N_21503,N_20058,N_20857);
or U21504 (N_21504,N_20085,N_20399);
xnor U21505 (N_21505,N_20207,N_20543);
nand U21506 (N_21506,N_20311,N_20463);
or U21507 (N_21507,N_20069,N_20335);
xor U21508 (N_21508,N_20114,N_20025);
nand U21509 (N_21509,N_20313,N_20155);
and U21510 (N_21510,N_20638,N_20254);
nor U21511 (N_21511,N_20873,N_20301);
xnor U21512 (N_21512,N_20800,N_20500);
and U21513 (N_21513,N_20284,N_20156);
or U21514 (N_21514,N_20720,N_20553);
xnor U21515 (N_21515,N_20747,N_20367);
and U21516 (N_21516,N_20001,N_20339);
nand U21517 (N_21517,N_20226,N_20138);
or U21518 (N_21518,N_20070,N_20508);
or U21519 (N_21519,N_20479,N_20643);
xor U21520 (N_21520,N_20897,N_20821);
xnor U21521 (N_21521,N_20294,N_20029);
or U21522 (N_21522,N_20025,N_20615);
xnor U21523 (N_21523,N_20612,N_20518);
nand U21524 (N_21524,N_20748,N_20688);
and U21525 (N_21525,N_20861,N_20834);
xnor U21526 (N_21526,N_20264,N_20911);
nand U21527 (N_21527,N_20264,N_20460);
and U21528 (N_21528,N_20638,N_20603);
nor U21529 (N_21529,N_20977,N_20005);
xnor U21530 (N_21530,N_20760,N_20353);
nand U21531 (N_21531,N_20160,N_20969);
nand U21532 (N_21532,N_20429,N_20312);
or U21533 (N_21533,N_20323,N_20442);
or U21534 (N_21534,N_20660,N_20154);
and U21535 (N_21535,N_20585,N_20615);
and U21536 (N_21536,N_20315,N_20140);
nand U21537 (N_21537,N_20611,N_20347);
xnor U21538 (N_21538,N_20476,N_20346);
xor U21539 (N_21539,N_20432,N_20648);
xor U21540 (N_21540,N_20679,N_20079);
or U21541 (N_21541,N_20480,N_20247);
and U21542 (N_21542,N_20033,N_20618);
xnor U21543 (N_21543,N_20806,N_20702);
nand U21544 (N_21544,N_20617,N_20835);
or U21545 (N_21545,N_20870,N_20584);
xor U21546 (N_21546,N_20960,N_20882);
or U21547 (N_21547,N_20222,N_20888);
xnor U21548 (N_21548,N_20893,N_20585);
or U21549 (N_21549,N_20304,N_20196);
and U21550 (N_21550,N_20714,N_20604);
xnor U21551 (N_21551,N_20670,N_20459);
and U21552 (N_21552,N_20106,N_20496);
nand U21553 (N_21553,N_20434,N_20323);
and U21554 (N_21554,N_20051,N_20486);
and U21555 (N_21555,N_20153,N_20416);
and U21556 (N_21556,N_20428,N_20377);
nor U21557 (N_21557,N_20253,N_20806);
or U21558 (N_21558,N_20530,N_20236);
and U21559 (N_21559,N_20371,N_20324);
nand U21560 (N_21560,N_20454,N_20413);
xor U21561 (N_21561,N_20014,N_20808);
or U21562 (N_21562,N_20440,N_20042);
or U21563 (N_21563,N_20139,N_20809);
xnor U21564 (N_21564,N_20142,N_20197);
or U21565 (N_21565,N_20717,N_20661);
or U21566 (N_21566,N_20766,N_20820);
and U21567 (N_21567,N_20075,N_20305);
xnor U21568 (N_21568,N_20533,N_20195);
nand U21569 (N_21569,N_20192,N_20748);
nand U21570 (N_21570,N_20838,N_20831);
nor U21571 (N_21571,N_20562,N_20479);
or U21572 (N_21572,N_20921,N_20043);
nand U21573 (N_21573,N_20430,N_20432);
xor U21574 (N_21574,N_20053,N_20409);
nor U21575 (N_21575,N_20181,N_20649);
nand U21576 (N_21576,N_20126,N_20204);
xnor U21577 (N_21577,N_20841,N_20078);
nand U21578 (N_21578,N_20202,N_20328);
xnor U21579 (N_21579,N_20361,N_20098);
and U21580 (N_21580,N_20086,N_20466);
nor U21581 (N_21581,N_20768,N_20581);
nor U21582 (N_21582,N_20450,N_20393);
xor U21583 (N_21583,N_20457,N_20631);
or U21584 (N_21584,N_20333,N_20573);
or U21585 (N_21585,N_20394,N_20180);
nor U21586 (N_21586,N_20418,N_20738);
xnor U21587 (N_21587,N_20566,N_20885);
or U21588 (N_21588,N_20203,N_20242);
and U21589 (N_21589,N_20268,N_20989);
xor U21590 (N_21590,N_20489,N_20542);
nand U21591 (N_21591,N_20367,N_20795);
xor U21592 (N_21592,N_20509,N_20177);
xor U21593 (N_21593,N_20829,N_20067);
and U21594 (N_21594,N_20176,N_20516);
nand U21595 (N_21595,N_20244,N_20832);
and U21596 (N_21596,N_20341,N_20351);
nand U21597 (N_21597,N_20371,N_20014);
and U21598 (N_21598,N_20826,N_20783);
nor U21599 (N_21599,N_20956,N_20188);
or U21600 (N_21600,N_20006,N_20461);
nand U21601 (N_21601,N_20204,N_20210);
or U21602 (N_21602,N_20733,N_20715);
nor U21603 (N_21603,N_20672,N_20860);
nand U21604 (N_21604,N_20188,N_20373);
nor U21605 (N_21605,N_20857,N_20720);
and U21606 (N_21606,N_20501,N_20213);
and U21607 (N_21607,N_20827,N_20442);
nand U21608 (N_21608,N_20340,N_20433);
nor U21609 (N_21609,N_20422,N_20485);
or U21610 (N_21610,N_20757,N_20377);
xnor U21611 (N_21611,N_20171,N_20865);
xnor U21612 (N_21612,N_20929,N_20693);
xnor U21613 (N_21613,N_20843,N_20003);
or U21614 (N_21614,N_20285,N_20775);
nor U21615 (N_21615,N_20216,N_20336);
or U21616 (N_21616,N_20843,N_20432);
nand U21617 (N_21617,N_20429,N_20159);
xnor U21618 (N_21618,N_20323,N_20212);
or U21619 (N_21619,N_20212,N_20151);
xnor U21620 (N_21620,N_20386,N_20086);
nand U21621 (N_21621,N_20319,N_20831);
nor U21622 (N_21622,N_20320,N_20720);
and U21623 (N_21623,N_20692,N_20701);
or U21624 (N_21624,N_20417,N_20837);
nand U21625 (N_21625,N_20253,N_20160);
and U21626 (N_21626,N_20958,N_20618);
xnor U21627 (N_21627,N_20511,N_20172);
xnor U21628 (N_21628,N_20732,N_20719);
nor U21629 (N_21629,N_20232,N_20162);
or U21630 (N_21630,N_20077,N_20099);
xnor U21631 (N_21631,N_20387,N_20409);
or U21632 (N_21632,N_20456,N_20785);
nand U21633 (N_21633,N_20228,N_20525);
and U21634 (N_21634,N_20488,N_20807);
xnor U21635 (N_21635,N_20035,N_20536);
or U21636 (N_21636,N_20553,N_20817);
xor U21637 (N_21637,N_20728,N_20570);
xnor U21638 (N_21638,N_20826,N_20229);
nand U21639 (N_21639,N_20316,N_20673);
nor U21640 (N_21640,N_20209,N_20041);
or U21641 (N_21641,N_20854,N_20924);
xor U21642 (N_21642,N_20278,N_20224);
or U21643 (N_21643,N_20740,N_20339);
nand U21644 (N_21644,N_20347,N_20043);
or U21645 (N_21645,N_20369,N_20152);
nand U21646 (N_21646,N_20011,N_20748);
nand U21647 (N_21647,N_20882,N_20859);
and U21648 (N_21648,N_20214,N_20088);
nor U21649 (N_21649,N_20447,N_20519);
xor U21650 (N_21650,N_20461,N_20592);
and U21651 (N_21651,N_20501,N_20479);
or U21652 (N_21652,N_20333,N_20555);
nand U21653 (N_21653,N_20652,N_20871);
xor U21654 (N_21654,N_20986,N_20696);
and U21655 (N_21655,N_20755,N_20294);
xor U21656 (N_21656,N_20347,N_20060);
and U21657 (N_21657,N_20602,N_20351);
or U21658 (N_21658,N_20718,N_20159);
or U21659 (N_21659,N_20406,N_20412);
xnor U21660 (N_21660,N_20346,N_20991);
or U21661 (N_21661,N_20109,N_20948);
nor U21662 (N_21662,N_20192,N_20670);
xnor U21663 (N_21663,N_20200,N_20438);
xnor U21664 (N_21664,N_20658,N_20671);
or U21665 (N_21665,N_20184,N_20244);
xor U21666 (N_21666,N_20322,N_20830);
and U21667 (N_21667,N_20411,N_20147);
nand U21668 (N_21668,N_20396,N_20873);
nand U21669 (N_21669,N_20195,N_20042);
nand U21670 (N_21670,N_20839,N_20122);
or U21671 (N_21671,N_20600,N_20205);
nor U21672 (N_21672,N_20361,N_20953);
nor U21673 (N_21673,N_20491,N_20028);
and U21674 (N_21674,N_20389,N_20668);
and U21675 (N_21675,N_20505,N_20893);
nor U21676 (N_21676,N_20755,N_20810);
xnor U21677 (N_21677,N_20333,N_20932);
and U21678 (N_21678,N_20311,N_20635);
nand U21679 (N_21679,N_20073,N_20307);
xor U21680 (N_21680,N_20681,N_20180);
xor U21681 (N_21681,N_20194,N_20129);
and U21682 (N_21682,N_20151,N_20408);
or U21683 (N_21683,N_20015,N_20329);
nor U21684 (N_21684,N_20125,N_20346);
and U21685 (N_21685,N_20113,N_20912);
or U21686 (N_21686,N_20728,N_20938);
nor U21687 (N_21687,N_20154,N_20569);
xnor U21688 (N_21688,N_20582,N_20588);
nor U21689 (N_21689,N_20249,N_20709);
nor U21690 (N_21690,N_20689,N_20640);
and U21691 (N_21691,N_20876,N_20303);
nand U21692 (N_21692,N_20558,N_20503);
or U21693 (N_21693,N_20753,N_20885);
or U21694 (N_21694,N_20899,N_20990);
nor U21695 (N_21695,N_20685,N_20957);
and U21696 (N_21696,N_20010,N_20048);
and U21697 (N_21697,N_20149,N_20531);
xnor U21698 (N_21698,N_20922,N_20058);
xnor U21699 (N_21699,N_20312,N_20697);
nor U21700 (N_21700,N_20284,N_20913);
or U21701 (N_21701,N_20021,N_20615);
nand U21702 (N_21702,N_20081,N_20933);
or U21703 (N_21703,N_20774,N_20771);
or U21704 (N_21704,N_20077,N_20758);
nand U21705 (N_21705,N_20095,N_20479);
or U21706 (N_21706,N_20373,N_20650);
nor U21707 (N_21707,N_20568,N_20298);
nand U21708 (N_21708,N_20117,N_20951);
xor U21709 (N_21709,N_20162,N_20001);
xor U21710 (N_21710,N_20803,N_20665);
and U21711 (N_21711,N_20337,N_20769);
nand U21712 (N_21712,N_20967,N_20287);
and U21713 (N_21713,N_20876,N_20884);
and U21714 (N_21714,N_20142,N_20277);
and U21715 (N_21715,N_20004,N_20718);
or U21716 (N_21716,N_20251,N_20139);
nor U21717 (N_21717,N_20565,N_20511);
nand U21718 (N_21718,N_20578,N_20325);
nand U21719 (N_21719,N_20718,N_20471);
and U21720 (N_21720,N_20352,N_20689);
or U21721 (N_21721,N_20960,N_20372);
nor U21722 (N_21722,N_20739,N_20927);
nand U21723 (N_21723,N_20959,N_20374);
nand U21724 (N_21724,N_20091,N_20834);
nand U21725 (N_21725,N_20438,N_20593);
or U21726 (N_21726,N_20781,N_20900);
nand U21727 (N_21727,N_20287,N_20401);
nor U21728 (N_21728,N_20679,N_20117);
nor U21729 (N_21729,N_20378,N_20876);
and U21730 (N_21730,N_20770,N_20949);
or U21731 (N_21731,N_20230,N_20634);
or U21732 (N_21732,N_20990,N_20618);
and U21733 (N_21733,N_20617,N_20282);
nor U21734 (N_21734,N_20097,N_20479);
and U21735 (N_21735,N_20174,N_20026);
xor U21736 (N_21736,N_20359,N_20881);
nor U21737 (N_21737,N_20051,N_20369);
or U21738 (N_21738,N_20267,N_20836);
and U21739 (N_21739,N_20100,N_20414);
and U21740 (N_21740,N_20926,N_20651);
xor U21741 (N_21741,N_20176,N_20485);
nand U21742 (N_21742,N_20851,N_20559);
or U21743 (N_21743,N_20972,N_20234);
nor U21744 (N_21744,N_20380,N_20466);
nor U21745 (N_21745,N_20717,N_20294);
xor U21746 (N_21746,N_20275,N_20004);
xor U21747 (N_21747,N_20369,N_20304);
xnor U21748 (N_21748,N_20935,N_20603);
nand U21749 (N_21749,N_20834,N_20592);
nand U21750 (N_21750,N_20041,N_20525);
and U21751 (N_21751,N_20219,N_20159);
nor U21752 (N_21752,N_20913,N_20461);
nand U21753 (N_21753,N_20110,N_20255);
and U21754 (N_21754,N_20109,N_20681);
nand U21755 (N_21755,N_20951,N_20103);
nand U21756 (N_21756,N_20222,N_20461);
nor U21757 (N_21757,N_20401,N_20701);
nor U21758 (N_21758,N_20732,N_20702);
xor U21759 (N_21759,N_20308,N_20373);
or U21760 (N_21760,N_20171,N_20808);
or U21761 (N_21761,N_20544,N_20382);
nor U21762 (N_21762,N_20617,N_20926);
nand U21763 (N_21763,N_20066,N_20607);
xor U21764 (N_21764,N_20219,N_20532);
nor U21765 (N_21765,N_20607,N_20286);
nand U21766 (N_21766,N_20124,N_20912);
or U21767 (N_21767,N_20762,N_20135);
xnor U21768 (N_21768,N_20664,N_20074);
xor U21769 (N_21769,N_20282,N_20620);
nand U21770 (N_21770,N_20548,N_20493);
nor U21771 (N_21771,N_20806,N_20747);
and U21772 (N_21772,N_20771,N_20188);
xor U21773 (N_21773,N_20746,N_20452);
xnor U21774 (N_21774,N_20167,N_20096);
nand U21775 (N_21775,N_20406,N_20050);
nand U21776 (N_21776,N_20425,N_20182);
nor U21777 (N_21777,N_20299,N_20210);
xnor U21778 (N_21778,N_20632,N_20183);
nor U21779 (N_21779,N_20465,N_20847);
xnor U21780 (N_21780,N_20266,N_20199);
or U21781 (N_21781,N_20373,N_20048);
and U21782 (N_21782,N_20219,N_20338);
nand U21783 (N_21783,N_20260,N_20163);
nor U21784 (N_21784,N_20362,N_20618);
or U21785 (N_21785,N_20626,N_20423);
nand U21786 (N_21786,N_20993,N_20512);
xor U21787 (N_21787,N_20656,N_20082);
nand U21788 (N_21788,N_20987,N_20344);
and U21789 (N_21789,N_20143,N_20715);
or U21790 (N_21790,N_20899,N_20649);
xor U21791 (N_21791,N_20058,N_20102);
nand U21792 (N_21792,N_20155,N_20872);
or U21793 (N_21793,N_20317,N_20223);
nor U21794 (N_21794,N_20885,N_20404);
xnor U21795 (N_21795,N_20625,N_20293);
nor U21796 (N_21796,N_20756,N_20123);
or U21797 (N_21797,N_20435,N_20002);
nand U21798 (N_21798,N_20058,N_20996);
nand U21799 (N_21799,N_20417,N_20328);
nor U21800 (N_21800,N_20895,N_20892);
or U21801 (N_21801,N_20022,N_20943);
xnor U21802 (N_21802,N_20602,N_20160);
or U21803 (N_21803,N_20455,N_20213);
and U21804 (N_21804,N_20737,N_20965);
nor U21805 (N_21805,N_20330,N_20207);
xnor U21806 (N_21806,N_20422,N_20302);
or U21807 (N_21807,N_20163,N_20853);
or U21808 (N_21808,N_20282,N_20036);
and U21809 (N_21809,N_20976,N_20554);
nor U21810 (N_21810,N_20519,N_20085);
nand U21811 (N_21811,N_20951,N_20880);
and U21812 (N_21812,N_20974,N_20291);
or U21813 (N_21813,N_20954,N_20105);
nand U21814 (N_21814,N_20151,N_20094);
or U21815 (N_21815,N_20292,N_20170);
nor U21816 (N_21816,N_20857,N_20179);
and U21817 (N_21817,N_20086,N_20308);
and U21818 (N_21818,N_20686,N_20266);
nand U21819 (N_21819,N_20487,N_20340);
xor U21820 (N_21820,N_20669,N_20007);
xnor U21821 (N_21821,N_20564,N_20230);
nor U21822 (N_21822,N_20565,N_20233);
and U21823 (N_21823,N_20079,N_20041);
or U21824 (N_21824,N_20479,N_20341);
nand U21825 (N_21825,N_20895,N_20996);
nor U21826 (N_21826,N_20456,N_20566);
xnor U21827 (N_21827,N_20362,N_20972);
and U21828 (N_21828,N_20614,N_20513);
and U21829 (N_21829,N_20003,N_20386);
and U21830 (N_21830,N_20350,N_20984);
xnor U21831 (N_21831,N_20627,N_20741);
or U21832 (N_21832,N_20946,N_20090);
nand U21833 (N_21833,N_20699,N_20577);
nor U21834 (N_21834,N_20315,N_20080);
or U21835 (N_21835,N_20072,N_20029);
and U21836 (N_21836,N_20546,N_20952);
or U21837 (N_21837,N_20758,N_20115);
or U21838 (N_21838,N_20641,N_20026);
nand U21839 (N_21839,N_20819,N_20679);
nand U21840 (N_21840,N_20275,N_20964);
and U21841 (N_21841,N_20055,N_20958);
nor U21842 (N_21842,N_20694,N_20152);
xor U21843 (N_21843,N_20607,N_20054);
nor U21844 (N_21844,N_20858,N_20316);
and U21845 (N_21845,N_20979,N_20281);
xnor U21846 (N_21846,N_20472,N_20154);
nor U21847 (N_21847,N_20257,N_20830);
or U21848 (N_21848,N_20561,N_20849);
xnor U21849 (N_21849,N_20587,N_20528);
nand U21850 (N_21850,N_20852,N_20614);
and U21851 (N_21851,N_20121,N_20391);
or U21852 (N_21852,N_20577,N_20516);
or U21853 (N_21853,N_20594,N_20233);
nor U21854 (N_21854,N_20570,N_20342);
or U21855 (N_21855,N_20678,N_20515);
or U21856 (N_21856,N_20982,N_20680);
and U21857 (N_21857,N_20866,N_20336);
xnor U21858 (N_21858,N_20950,N_20027);
and U21859 (N_21859,N_20385,N_20712);
and U21860 (N_21860,N_20417,N_20433);
nor U21861 (N_21861,N_20796,N_20525);
or U21862 (N_21862,N_20164,N_20404);
or U21863 (N_21863,N_20741,N_20556);
nand U21864 (N_21864,N_20706,N_20104);
xnor U21865 (N_21865,N_20305,N_20280);
or U21866 (N_21866,N_20088,N_20881);
and U21867 (N_21867,N_20911,N_20005);
nand U21868 (N_21868,N_20764,N_20943);
nor U21869 (N_21869,N_20641,N_20068);
xnor U21870 (N_21870,N_20447,N_20279);
nor U21871 (N_21871,N_20311,N_20327);
and U21872 (N_21872,N_20241,N_20947);
nand U21873 (N_21873,N_20081,N_20330);
and U21874 (N_21874,N_20573,N_20262);
nor U21875 (N_21875,N_20929,N_20893);
and U21876 (N_21876,N_20718,N_20678);
nor U21877 (N_21877,N_20138,N_20549);
nand U21878 (N_21878,N_20930,N_20424);
xor U21879 (N_21879,N_20206,N_20790);
xor U21880 (N_21880,N_20185,N_20766);
nand U21881 (N_21881,N_20395,N_20133);
or U21882 (N_21882,N_20250,N_20145);
nor U21883 (N_21883,N_20773,N_20109);
xnor U21884 (N_21884,N_20506,N_20051);
or U21885 (N_21885,N_20904,N_20583);
nand U21886 (N_21886,N_20911,N_20590);
nor U21887 (N_21887,N_20529,N_20056);
nor U21888 (N_21888,N_20899,N_20091);
nor U21889 (N_21889,N_20968,N_20824);
nor U21890 (N_21890,N_20303,N_20218);
or U21891 (N_21891,N_20754,N_20689);
or U21892 (N_21892,N_20740,N_20075);
nor U21893 (N_21893,N_20466,N_20617);
and U21894 (N_21894,N_20223,N_20221);
nand U21895 (N_21895,N_20572,N_20030);
nor U21896 (N_21896,N_20269,N_20365);
xnor U21897 (N_21897,N_20262,N_20620);
or U21898 (N_21898,N_20666,N_20965);
and U21899 (N_21899,N_20623,N_20695);
nor U21900 (N_21900,N_20229,N_20450);
or U21901 (N_21901,N_20459,N_20088);
nor U21902 (N_21902,N_20558,N_20686);
or U21903 (N_21903,N_20618,N_20529);
nor U21904 (N_21904,N_20357,N_20824);
nor U21905 (N_21905,N_20873,N_20774);
xor U21906 (N_21906,N_20850,N_20388);
xor U21907 (N_21907,N_20075,N_20303);
nor U21908 (N_21908,N_20863,N_20487);
xnor U21909 (N_21909,N_20729,N_20478);
and U21910 (N_21910,N_20009,N_20407);
nor U21911 (N_21911,N_20337,N_20333);
or U21912 (N_21912,N_20137,N_20165);
nand U21913 (N_21913,N_20422,N_20609);
and U21914 (N_21914,N_20417,N_20149);
nand U21915 (N_21915,N_20556,N_20219);
nor U21916 (N_21916,N_20430,N_20647);
nor U21917 (N_21917,N_20323,N_20746);
nand U21918 (N_21918,N_20824,N_20847);
xor U21919 (N_21919,N_20470,N_20533);
and U21920 (N_21920,N_20031,N_20833);
or U21921 (N_21921,N_20967,N_20565);
xor U21922 (N_21922,N_20528,N_20150);
nor U21923 (N_21923,N_20990,N_20559);
xnor U21924 (N_21924,N_20715,N_20250);
nor U21925 (N_21925,N_20923,N_20458);
and U21926 (N_21926,N_20940,N_20511);
xor U21927 (N_21927,N_20450,N_20698);
nor U21928 (N_21928,N_20768,N_20500);
nor U21929 (N_21929,N_20780,N_20356);
nor U21930 (N_21930,N_20671,N_20071);
xor U21931 (N_21931,N_20458,N_20411);
nor U21932 (N_21932,N_20172,N_20932);
xor U21933 (N_21933,N_20510,N_20288);
nor U21934 (N_21934,N_20273,N_20808);
nor U21935 (N_21935,N_20035,N_20495);
xor U21936 (N_21936,N_20308,N_20644);
nor U21937 (N_21937,N_20663,N_20483);
or U21938 (N_21938,N_20976,N_20343);
nand U21939 (N_21939,N_20024,N_20385);
nand U21940 (N_21940,N_20727,N_20051);
and U21941 (N_21941,N_20705,N_20693);
nand U21942 (N_21942,N_20685,N_20046);
and U21943 (N_21943,N_20894,N_20811);
xnor U21944 (N_21944,N_20057,N_20200);
xor U21945 (N_21945,N_20629,N_20899);
xor U21946 (N_21946,N_20649,N_20242);
nor U21947 (N_21947,N_20249,N_20925);
and U21948 (N_21948,N_20462,N_20362);
xnor U21949 (N_21949,N_20197,N_20718);
or U21950 (N_21950,N_20933,N_20712);
nand U21951 (N_21951,N_20457,N_20881);
and U21952 (N_21952,N_20841,N_20045);
xor U21953 (N_21953,N_20148,N_20033);
nand U21954 (N_21954,N_20624,N_20905);
nand U21955 (N_21955,N_20811,N_20924);
xnor U21956 (N_21956,N_20310,N_20976);
xor U21957 (N_21957,N_20415,N_20071);
nand U21958 (N_21958,N_20231,N_20267);
nand U21959 (N_21959,N_20780,N_20118);
or U21960 (N_21960,N_20201,N_20751);
or U21961 (N_21961,N_20523,N_20480);
nand U21962 (N_21962,N_20327,N_20841);
nand U21963 (N_21963,N_20591,N_20657);
or U21964 (N_21964,N_20531,N_20495);
nand U21965 (N_21965,N_20930,N_20585);
nand U21966 (N_21966,N_20582,N_20542);
or U21967 (N_21967,N_20910,N_20824);
nor U21968 (N_21968,N_20309,N_20247);
and U21969 (N_21969,N_20934,N_20203);
nand U21970 (N_21970,N_20680,N_20851);
and U21971 (N_21971,N_20614,N_20422);
and U21972 (N_21972,N_20936,N_20300);
nand U21973 (N_21973,N_20018,N_20060);
xnor U21974 (N_21974,N_20231,N_20470);
nand U21975 (N_21975,N_20570,N_20719);
nor U21976 (N_21976,N_20239,N_20513);
xor U21977 (N_21977,N_20257,N_20531);
or U21978 (N_21978,N_20212,N_20088);
nand U21979 (N_21979,N_20865,N_20397);
and U21980 (N_21980,N_20781,N_20778);
and U21981 (N_21981,N_20777,N_20464);
nor U21982 (N_21982,N_20190,N_20336);
nor U21983 (N_21983,N_20491,N_20894);
xnor U21984 (N_21984,N_20056,N_20066);
xor U21985 (N_21985,N_20480,N_20935);
xor U21986 (N_21986,N_20128,N_20264);
and U21987 (N_21987,N_20080,N_20260);
nand U21988 (N_21988,N_20386,N_20772);
and U21989 (N_21989,N_20104,N_20627);
nor U21990 (N_21990,N_20269,N_20398);
nor U21991 (N_21991,N_20355,N_20080);
nor U21992 (N_21992,N_20015,N_20495);
nor U21993 (N_21993,N_20846,N_20599);
xor U21994 (N_21994,N_20635,N_20193);
and U21995 (N_21995,N_20162,N_20769);
nand U21996 (N_21996,N_20633,N_20045);
nand U21997 (N_21997,N_20409,N_20411);
and U21998 (N_21998,N_20705,N_20675);
and U21999 (N_21999,N_20813,N_20748);
nand U22000 (N_22000,N_21712,N_21682);
nor U22001 (N_22001,N_21605,N_21063);
xnor U22002 (N_22002,N_21872,N_21991);
and U22003 (N_22003,N_21793,N_21962);
nand U22004 (N_22004,N_21936,N_21649);
and U22005 (N_22005,N_21466,N_21791);
nor U22006 (N_22006,N_21027,N_21358);
xnor U22007 (N_22007,N_21173,N_21538);
and U22008 (N_22008,N_21365,N_21454);
or U22009 (N_22009,N_21688,N_21164);
nor U22010 (N_22010,N_21390,N_21951);
or U22011 (N_22011,N_21505,N_21205);
nor U22012 (N_22012,N_21092,N_21362);
xnor U22013 (N_22013,N_21786,N_21488);
and U22014 (N_22014,N_21705,N_21609);
xnor U22015 (N_22015,N_21217,N_21414);
nor U22016 (N_22016,N_21213,N_21635);
nand U22017 (N_22017,N_21133,N_21338);
or U22018 (N_22018,N_21896,N_21781);
and U22019 (N_22019,N_21687,N_21168);
nor U22020 (N_22020,N_21070,N_21835);
xor U22021 (N_22021,N_21306,N_21648);
and U22022 (N_22022,N_21859,N_21785);
nand U22023 (N_22023,N_21273,N_21129);
or U22024 (N_22024,N_21940,N_21715);
and U22025 (N_22025,N_21579,N_21776);
nand U22026 (N_22026,N_21446,N_21097);
or U22027 (N_22027,N_21714,N_21483);
xnor U22028 (N_22028,N_21572,N_21091);
and U22029 (N_22029,N_21053,N_21911);
nand U22030 (N_22030,N_21815,N_21704);
or U22031 (N_22031,N_21248,N_21669);
and U22032 (N_22032,N_21713,N_21980);
xor U22033 (N_22033,N_21462,N_21800);
xor U22034 (N_22034,N_21693,N_21310);
nand U22035 (N_22035,N_21566,N_21726);
and U22036 (N_22036,N_21549,N_21986);
nand U22037 (N_22037,N_21371,N_21025);
or U22038 (N_22038,N_21661,N_21313);
nand U22039 (N_22039,N_21254,N_21607);
or U22040 (N_22040,N_21860,N_21795);
nor U22041 (N_22041,N_21169,N_21207);
and U22042 (N_22042,N_21455,N_21469);
nor U22043 (N_22043,N_21270,N_21196);
nor U22044 (N_22044,N_21198,N_21342);
nor U22045 (N_22045,N_21385,N_21087);
nor U22046 (N_22046,N_21271,N_21482);
nor U22047 (N_22047,N_21354,N_21801);
or U22048 (N_22048,N_21743,N_21100);
xor U22049 (N_22049,N_21560,N_21664);
and U22050 (N_22050,N_21161,N_21770);
nor U22051 (N_22051,N_21866,N_21914);
nor U22052 (N_22052,N_21305,N_21151);
nand U22053 (N_22053,N_21002,N_21812);
and U22054 (N_22054,N_21646,N_21039);
nand U22055 (N_22055,N_21178,N_21094);
xnor U22056 (N_22056,N_21283,N_21355);
or U22057 (N_22057,N_21910,N_21622);
nand U22058 (N_22058,N_21465,N_21842);
xor U22059 (N_22059,N_21852,N_21337);
xor U22060 (N_22060,N_21948,N_21124);
and U22061 (N_22061,N_21890,N_21259);
nand U22062 (N_22062,N_21246,N_21925);
or U22063 (N_22063,N_21819,N_21432);
xor U22064 (N_22064,N_21437,N_21757);
and U22065 (N_22065,N_21279,N_21807);
and U22066 (N_22066,N_21899,N_21231);
nand U22067 (N_22067,N_21093,N_21453);
and U22068 (N_22068,N_21824,N_21000);
nor U22069 (N_22069,N_21944,N_21753);
xnor U22070 (N_22070,N_21473,N_21869);
or U22071 (N_22071,N_21536,N_21191);
nand U22072 (N_22072,N_21802,N_21810);
nor U22073 (N_22073,N_21877,N_21929);
nor U22074 (N_22074,N_21644,N_21406);
or U22075 (N_22075,N_21627,N_21838);
nand U22076 (N_22076,N_21917,N_21463);
nand U22077 (N_22077,N_21489,N_21061);
xnor U22078 (N_22078,N_21357,N_21546);
xnor U22079 (N_22079,N_21998,N_21398);
or U22080 (N_22080,N_21269,N_21327);
or U22081 (N_22081,N_21799,N_21486);
xor U22082 (N_22082,N_21267,N_21081);
xor U22083 (N_22083,N_21862,N_21253);
nor U22084 (N_22084,N_21435,N_21439);
and U22085 (N_22085,N_21710,N_21485);
xnor U22086 (N_22086,N_21449,N_21378);
xnor U22087 (N_22087,N_21677,N_21806);
or U22088 (N_22088,N_21245,N_21452);
or U22089 (N_22089,N_21729,N_21018);
nand U22090 (N_22090,N_21540,N_21008);
xnor U22091 (N_22091,N_21364,N_21846);
or U22092 (N_22092,N_21528,N_21578);
nand U22093 (N_22093,N_21317,N_21922);
or U22094 (N_22094,N_21755,N_21592);
or U22095 (N_22095,N_21159,N_21185);
or U22096 (N_22096,N_21663,N_21968);
xor U22097 (N_22097,N_21882,N_21274);
nand U22098 (N_22098,N_21915,N_21585);
and U22099 (N_22099,N_21695,N_21656);
nand U22100 (N_22100,N_21352,N_21156);
xnor U22101 (N_22101,N_21707,N_21557);
nand U22102 (N_22102,N_21766,N_21360);
and U22103 (N_22103,N_21029,N_21567);
nor U22104 (N_22104,N_21044,N_21670);
nor U22105 (N_22105,N_21484,N_21889);
xnor U22106 (N_22106,N_21820,N_21004);
nor U22107 (N_22107,N_21181,N_21665);
xor U22108 (N_22108,N_21510,N_21777);
nor U22109 (N_22109,N_21771,N_21376);
nor U22110 (N_22110,N_21830,N_21224);
nor U22111 (N_22111,N_21285,N_21192);
nor U22112 (N_22112,N_21532,N_21533);
and U22113 (N_22113,N_21932,N_21021);
nor U22114 (N_22114,N_21689,N_21772);
xnor U22115 (N_22115,N_21901,N_21085);
or U22116 (N_22116,N_21539,N_21754);
xor U22117 (N_22117,N_21904,N_21288);
or U22118 (N_22118,N_21878,N_21593);
xnor U22119 (N_22119,N_21808,N_21928);
xor U22120 (N_22120,N_21924,N_21997);
or U22121 (N_22121,N_21500,N_21424);
xor U22122 (N_22122,N_21598,N_21227);
and U22123 (N_22123,N_21933,N_21006);
nor U22124 (N_22124,N_21938,N_21076);
or U22125 (N_22125,N_21783,N_21407);
nand U22126 (N_22126,N_21410,N_21652);
nor U22127 (N_22127,N_21268,N_21903);
or U22128 (N_22128,N_21067,N_21126);
and U22129 (N_22129,N_21611,N_21134);
or U22130 (N_22130,N_21131,N_21303);
nand U22131 (N_22131,N_21017,N_21412);
and U22132 (N_22132,N_21975,N_21573);
and U22133 (N_22133,N_21887,N_21601);
or U22134 (N_22134,N_21291,N_21056);
xor U22135 (N_22135,N_21511,N_21966);
and U22136 (N_22136,N_21865,N_21767);
and U22137 (N_22137,N_21850,N_21803);
and U22138 (N_22138,N_21708,N_21316);
and U22139 (N_22139,N_21535,N_21956);
nand U22140 (N_22140,N_21604,N_21618);
or U22141 (N_22141,N_21072,N_21491);
nor U22142 (N_22142,N_21492,N_21993);
nor U22143 (N_22143,N_21702,N_21599);
nor U22144 (N_22144,N_21065,N_21554);
xnor U22145 (N_22145,N_21570,N_21828);
xnor U22146 (N_22146,N_21111,N_21400);
and U22147 (N_22147,N_21434,N_21871);
nor U22148 (N_22148,N_21375,N_21034);
or U22149 (N_22149,N_21955,N_21003);
or U22150 (N_22150,N_21633,N_21001);
or U22151 (N_22151,N_21608,N_21836);
and U22152 (N_22152,N_21071,N_21653);
or U22153 (N_22153,N_21613,N_21046);
or U22154 (N_22154,N_21210,N_21329);
xnor U22155 (N_22155,N_21894,N_21720);
or U22156 (N_22156,N_21119,N_21761);
nor U22157 (N_22157,N_21450,N_21768);
nor U22158 (N_22158,N_21615,N_21089);
nor U22159 (N_22159,N_21888,N_21361);
nand U22160 (N_22160,N_21632,N_21383);
or U22161 (N_22161,N_21293,N_21861);
nor U22162 (N_22162,N_21068,N_21983);
and U22163 (N_22163,N_21392,N_21393);
nor U22164 (N_22164,N_21154,N_21506);
nand U22165 (N_22165,N_21032,N_21879);
nand U22166 (N_22166,N_21988,N_21099);
nor U22167 (N_22167,N_21077,N_21654);
nor U22168 (N_22168,N_21897,N_21569);
and U22169 (N_22169,N_21222,N_21183);
nand U22170 (N_22170,N_21885,N_21884);
xor U22171 (N_22171,N_21722,N_21629);
nor U22172 (N_22172,N_21301,N_21199);
xnor U22173 (N_22173,N_21923,N_21582);
or U22174 (N_22174,N_21200,N_21149);
or U22175 (N_22175,N_21413,N_21110);
nand U22176 (N_22176,N_21289,N_21647);
nor U22177 (N_22177,N_21255,N_21165);
xor U22178 (N_22178,N_21543,N_21788);
nor U22179 (N_22179,N_21794,N_21234);
nand U22180 (N_22180,N_21942,N_21745);
and U22181 (N_22181,N_21645,N_21394);
and U22182 (N_22182,N_21396,N_21735);
or U22183 (N_22183,N_21740,N_21343);
or U22184 (N_22184,N_21128,N_21438);
and U22185 (N_22185,N_21937,N_21236);
xnor U22186 (N_22186,N_21934,N_21969);
xnor U22187 (N_22187,N_21155,N_21832);
nor U22188 (N_22188,N_21218,N_21818);
or U22189 (N_22189,N_21326,N_21822);
xor U22190 (N_22190,N_21177,N_21042);
or U22191 (N_22191,N_21706,N_21811);
nor U22192 (N_22192,N_21504,N_21575);
nand U22193 (N_22193,N_21606,N_21011);
and U22194 (N_22194,N_21130,N_21900);
xnor U22195 (N_22195,N_21941,N_21826);
xnor U22196 (N_22196,N_21694,N_21521);
xor U22197 (N_22197,N_21190,N_21610);
or U22198 (N_22198,N_21697,N_21717);
nor U22199 (N_22199,N_21841,N_21905);
or U22200 (N_22200,N_21858,N_21848);
nand U22201 (N_22201,N_21302,N_21215);
and U22202 (N_22202,N_21675,N_21122);
xor U22203 (N_22203,N_21105,N_21120);
xor U22204 (N_22204,N_21892,N_21079);
or U22205 (N_22205,N_21967,N_21958);
or U22206 (N_22206,N_21086,N_21686);
nor U22207 (N_22207,N_21395,N_21102);
or U22208 (N_22208,N_21143,N_21214);
and U22209 (N_22209,N_21014,N_21240);
xnor U22210 (N_22210,N_21223,N_21805);
or U22211 (N_22211,N_21363,N_21221);
nand U22212 (N_22212,N_21499,N_21749);
xnor U22213 (N_22213,N_21916,N_21278);
xor U22214 (N_22214,N_21103,N_21493);
nor U22215 (N_22215,N_21671,N_21262);
nor U22216 (N_22216,N_21368,N_21082);
or U22217 (N_22217,N_21583,N_21333);
nand U22218 (N_22218,N_21281,N_21049);
nand U22219 (N_22219,N_21537,N_21595);
nor U22220 (N_22220,N_21477,N_21977);
xnor U22221 (N_22221,N_21758,N_21837);
xnor U22222 (N_22222,N_21459,N_21487);
nor U22223 (N_22223,N_21060,N_21339);
nor U22224 (N_22224,N_21444,N_21284);
nand U22225 (N_22225,N_21429,N_21033);
nand U22226 (N_22226,N_21386,N_21321);
nor U22227 (N_22227,N_21296,N_21870);
nand U22228 (N_22228,N_21666,N_21351);
nand U22229 (N_22229,N_21926,N_21292);
and U22230 (N_22230,N_21513,N_21195);
and U22231 (N_22231,N_21346,N_21431);
nor U22232 (N_22232,N_21864,N_21171);
and U22233 (N_22233,N_21401,N_21447);
or U22234 (N_22234,N_21331,N_21445);
and U22235 (N_22235,N_21380,N_21636);
xnor U22236 (N_22236,N_21323,N_21348);
nor U22237 (N_22237,N_21732,N_21738);
nand U22238 (N_22238,N_21062,N_21733);
nor U22239 (N_22239,N_21990,N_21083);
nand U22240 (N_22240,N_21475,N_21055);
and U22241 (N_22241,N_21945,N_21849);
nand U22242 (N_22242,N_21409,N_21683);
and U22243 (N_22243,N_21202,N_21972);
and U22244 (N_22244,N_21280,N_21397);
nand U22245 (N_22245,N_21141,N_21565);
xnor U22246 (N_22246,N_21855,N_21495);
nor U22247 (N_22247,N_21624,N_21147);
xnor U22248 (N_22248,N_21287,N_21891);
nor U22249 (N_22249,N_21651,N_21035);
or U22250 (N_22250,N_21419,N_21229);
xor U22251 (N_22251,N_21698,N_21350);
or U22252 (N_22252,N_21947,N_21716);
xor U22253 (N_22253,N_21421,N_21881);
and U22254 (N_22254,N_21332,N_21209);
or U22255 (N_22255,N_21699,N_21369);
or U22256 (N_22256,N_21711,N_21760);
or U22257 (N_22257,N_21232,N_21544);
nand U22258 (N_22258,N_21529,N_21007);
and U22259 (N_22259,N_21531,N_21763);
or U22260 (N_22260,N_21256,N_21668);
and U22261 (N_22261,N_21643,N_21249);
or U22262 (N_22262,N_21561,N_21157);
and U22263 (N_22263,N_21679,N_21225);
and U22264 (N_22264,N_21964,N_21261);
or U22265 (N_22265,N_21718,N_21978);
nand U22266 (N_22266,N_21193,N_21797);
nor U22267 (N_22267,N_21873,N_21981);
and U22268 (N_22268,N_21789,N_21479);
nor U22269 (N_22269,N_21497,N_21108);
and U22270 (N_22270,N_21748,N_21244);
nor U22271 (N_22271,N_21010,N_21909);
and U22272 (N_22272,N_21286,N_21739);
nor U22273 (N_22273,N_21736,N_21809);
xnor U22274 (N_22274,N_21886,N_21744);
or U22275 (N_22275,N_21580,N_21825);
nor U22276 (N_22276,N_21050,N_21640);
or U22277 (N_22277,N_21659,N_21551);
nand U22278 (N_22278,N_21420,N_21160);
or U22279 (N_22279,N_21950,N_21023);
xor U22280 (N_22280,N_21180,N_21370);
nor U22281 (N_22281,N_21311,N_21912);
xor U22282 (N_22282,N_21075,N_21581);
or U22283 (N_22283,N_21005,N_21525);
xor U22284 (N_22284,N_21696,N_21919);
and U22285 (N_22285,N_21965,N_21073);
nor U22286 (N_22286,N_21300,N_21796);
xnor U22287 (N_22287,N_21047,N_21142);
or U22288 (N_22288,N_21031,N_21428);
xor U22289 (N_22289,N_21457,N_21979);
and U22290 (N_22290,N_21206,N_21069);
or U22291 (N_22291,N_21517,N_21555);
and U22292 (N_22292,N_21571,N_21960);
and U22293 (N_22293,N_21391,N_21084);
or U22294 (N_22294,N_21252,N_21526);
nor U22295 (N_22295,N_21631,N_21382);
and U22296 (N_22296,N_21752,N_21187);
xor U22297 (N_22297,N_21415,N_21762);
nand U22298 (N_22298,N_21472,N_21587);
xor U22299 (N_22299,N_21775,N_21325);
xnor U22300 (N_22300,N_21908,N_21136);
nand U22301 (N_22301,N_21625,N_21101);
and U22302 (N_22302,N_21064,N_21476);
nand U22303 (N_22303,N_21827,N_21448);
nor U22304 (N_22304,N_21700,N_21295);
nor U22305 (N_22305,N_21520,N_21863);
or U22306 (N_22306,N_21490,N_21427);
and U22307 (N_22307,N_21779,N_21931);
or U22308 (N_22308,N_21373,N_21436);
and U22309 (N_22309,N_21464,N_21139);
or U22310 (N_22310,N_21784,N_21541);
xor U22311 (N_22311,N_21674,N_21020);
xor U22312 (N_22312,N_21920,N_21603);
nand U22313 (N_22313,N_21260,N_21597);
xnor U22314 (N_22314,N_21530,N_21845);
nand U22315 (N_22315,N_21186,N_21829);
nand U22316 (N_22316,N_21673,N_21170);
xor U22317 (N_22317,N_21208,N_21389);
and U22318 (N_22318,N_21612,N_21773);
xor U22319 (N_22319,N_21843,N_21684);
and U22320 (N_22320,N_21742,N_21058);
xnor U22321 (N_22321,N_21523,N_21443);
nor U22322 (N_22322,N_21680,N_21201);
nor U22323 (N_22323,N_21408,N_21074);
nand U22324 (N_22324,N_21179,N_21125);
nand U22325 (N_22325,N_21913,N_21816);
and U22326 (N_22326,N_21096,N_21184);
or U22327 (N_22327,N_21411,N_21780);
or U22328 (N_22328,N_21322,N_21918);
and U22329 (N_22329,N_21764,N_21728);
or U22330 (N_22330,N_21774,N_21616);
nor U22331 (N_22331,N_21496,N_21038);
nand U22332 (N_22332,N_21344,N_21952);
xor U22333 (N_22333,N_21494,N_21468);
nand U22334 (N_22334,N_21949,N_21518);
nand U22335 (N_22335,N_21379,N_21556);
nor U22336 (N_22336,N_21216,N_21238);
nor U22337 (N_22337,N_21467,N_21297);
and U22338 (N_22338,N_21422,N_21782);
nor U22339 (N_22339,N_21558,N_21588);
and U22340 (N_22340,N_21174,N_21194);
nand U22341 (N_22341,N_21204,N_21778);
nand U22342 (N_22342,N_21703,N_21823);
nand U22343 (N_22343,N_21630,N_21115);
or U22344 (N_22344,N_21146,N_21586);
nand U22345 (N_22345,N_21349,N_21638);
nand U22346 (N_22346,N_21662,N_21921);
xnor U22347 (N_22347,N_21628,N_21876);
and U22348 (N_22348,N_21117,N_21963);
xor U22349 (N_22349,N_21522,N_21175);
xnor U22350 (N_22350,N_21095,N_21765);
nor U22351 (N_22351,N_21982,N_21377);
xnor U22352 (N_22352,N_21691,N_21241);
xor U22353 (N_22353,N_21999,N_21197);
or U22354 (N_22354,N_21239,N_21642);
nor U22355 (N_22355,N_21501,N_21471);
nand U22356 (N_22356,N_21048,N_21626);
nor U22357 (N_22357,N_21576,N_21856);
nor U22358 (N_22358,N_21264,N_21309);
nor U22359 (N_22359,N_21150,N_21430);
or U22360 (N_22360,N_21559,N_21813);
nand U22361 (N_22361,N_21009,N_21138);
or U22362 (N_22362,N_21750,N_21140);
or U22363 (N_22363,N_21080,N_21851);
xnor U22364 (N_22364,N_21243,N_21335);
nand U22365 (N_22365,N_21619,N_21515);
and U22366 (N_22366,N_21833,N_21875);
nand U22367 (N_22367,N_21634,N_21116);
or U22368 (N_22368,N_21868,N_21985);
nor U22369 (N_22369,N_21943,N_21040);
or U22370 (N_22370,N_21045,N_21534);
xnor U22371 (N_22371,N_21220,N_21498);
and U22372 (N_22372,N_21840,N_21078);
and U22373 (N_22373,N_21737,N_21387);
nor U22374 (N_22374,N_21562,N_21036);
xor U22375 (N_22375,N_21113,N_21992);
xor U22376 (N_22376,N_21163,N_21996);
nand U22377 (N_22377,N_21844,N_21328);
xor U22378 (N_22378,N_21366,N_21158);
and U22379 (N_22379,N_21481,N_21372);
xnor U22380 (N_22380,N_21509,N_21470);
and U22381 (N_22381,N_21347,N_21987);
nand U22382 (N_22382,N_21516,N_21106);
nand U22383 (N_22383,N_21416,N_21121);
and U22384 (N_22384,N_21594,N_21725);
nand U22385 (N_22385,N_21989,N_21502);
xnor U22386 (N_22386,N_21013,N_21650);
or U22387 (N_22387,N_21312,N_21553);
nor U22388 (N_22388,N_21660,N_21144);
and U22389 (N_22389,N_21568,N_21847);
xor U22390 (N_22390,N_21524,N_21584);
nor U22391 (N_22391,N_21821,N_21970);
xnor U22392 (N_22392,N_21589,N_21724);
xor U22393 (N_22393,N_21381,N_21266);
nor U22394 (N_22394,N_21162,N_21527);
nor U22395 (N_22395,N_21759,N_21374);
xnor U22396 (N_22396,N_21367,N_21623);
or U22397 (N_22397,N_21426,N_21247);
nor U22398 (N_22398,N_21016,N_21423);
nor U22399 (N_22399,N_21098,N_21024);
or U22400 (N_22400,N_21404,N_21188);
and U22401 (N_22401,N_21563,N_21104);
or U22402 (N_22402,N_21596,N_21456);
nand U22403 (N_22403,N_21953,N_21324);
xor U22404 (N_22404,N_21883,N_21230);
nor U22405 (N_22405,N_21730,N_21620);
nor U22406 (N_22406,N_21614,N_21514);
xnor U22407 (N_22407,N_21417,N_21641);
and U22408 (N_22408,N_21741,N_21550);
or U22409 (N_22409,N_21203,N_21734);
nand U22410 (N_22410,N_21577,N_21402);
nor U22411 (N_22411,N_21242,N_21330);
xnor U22412 (N_22412,N_21474,N_21685);
nor U22413 (N_22413,N_21314,N_21458);
and U22414 (N_22414,N_21817,N_21984);
nand U22415 (N_22415,N_21542,N_21057);
and U22416 (N_22416,N_21235,N_21405);
nor U22417 (N_22417,N_21356,N_21902);
xor U22418 (N_22418,N_21547,N_21480);
xor U22419 (N_22419,N_21804,N_21275);
xor U22420 (N_22420,N_21548,N_21219);
nor U22421 (N_22421,N_21359,N_21148);
or U22422 (N_22422,N_21552,N_21388);
xor U22423 (N_22423,N_21228,N_21692);
nor U22424 (N_22424,N_21441,N_21709);
nor U22425 (N_22425,N_21451,N_21345);
nor U22426 (N_22426,N_21746,N_21022);
nor U22427 (N_22427,N_21976,N_21336);
and U22428 (N_22428,N_21282,N_21090);
nand U22429 (N_22429,N_21907,N_21690);
and U22430 (N_22430,N_21959,N_21308);
nor U22431 (N_22431,N_21834,N_21545);
xnor U22432 (N_22432,N_21132,N_21166);
xnor U22433 (N_22433,N_21127,N_21798);
nor U22434 (N_22434,N_21418,N_21118);
xor U22435 (N_22435,N_21226,N_21257);
nor U22436 (N_22436,N_21026,N_21015);
or U22437 (N_22437,N_21874,N_21994);
nor U22438 (N_22438,N_21957,N_21425);
and U22439 (N_22439,N_21172,N_21137);
and U22440 (N_22440,N_21277,N_21676);
or U22441 (N_22441,N_21051,N_21112);
or U22442 (N_22442,N_21399,N_21028);
nand U22443 (N_22443,N_21440,N_21590);
xnor U22444 (N_22444,N_21574,N_21831);
and U22445 (N_22445,N_21319,N_21935);
or U22446 (N_22446,N_21756,N_21265);
and U22447 (N_22447,N_21353,N_21751);
nor U22448 (N_22448,N_21059,N_21176);
and U22449 (N_22449,N_21304,N_21681);
xnor U22450 (N_22450,N_21442,N_21995);
nand U22451 (N_22451,N_21189,N_21667);
xor U22452 (N_22452,N_21037,N_21971);
or U22453 (N_22453,N_21263,N_21299);
or U22454 (N_22454,N_21731,N_21946);
nor U22455 (N_22455,N_21012,N_21507);
or U22456 (N_22456,N_21600,N_21315);
xnor U22457 (N_22457,N_21272,N_21721);
nand U22458 (N_22458,N_21787,N_21839);
or U22459 (N_22459,N_21318,N_21602);
nand U22460 (N_22460,N_21639,N_21867);
and U22461 (N_22461,N_21320,N_21657);
nand U22462 (N_22462,N_21152,N_21294);
or U22463 (N_22463,N_21403,N_21961);
xor U22464 (N_22464,N_21727,N_21340);
xor U22465 (N_22465,N_21384,N_21719);
or U22466 (N_22466,N_21658,N_21052);
nand U22467 (N_22467,N_21433,N_21043);
nand U22468 (N_22468,N_21930,N_21123);
and U22469 (N_22469,N_21857,N_21814);
nor U22470 (N_22470,N_21107,N_21790);
nand U22471 (N_22471,N_21939,N_21334);
and U22472 (N_22472,N_21461,N_21853);
nand U22473 (N_22473,N_21250,N_21298);
or U22474 (N_22474,N_21898,N_21233);
xor U22475 (N_22475,N_21066,N_21030);
or U22476 (N_22476,N_21621,N_21769);
nand U22477 (N_22477,N_21276,N_21307);
nand U22478 (N_22478,N_21088,N_21927);
nor U22479 (N_22479,N_21974,N_21182);
and U22480 (N_22480,N_21564,N_21954);
and U22481 (N_22481,N_21251,N_21478);
or U22482 (N_22482,N_21019,N_21508);
nand U22483 (N_22483,N_21973,N_21591);
and U22484 (N_22484,N_21145,N_21895);
nor U22485 (N_22485,N_21792,N_21512);
and U22486 (N_22486,N_21237,N_21135);
xnor U22487 (N_22487,N_21211,N_21258);
xor U22488 (N_22488,N_21906,N_21460);
nor U22489 (N_22489,N_21880,N_21153);
nand U22490 (N_22490,N_21655,N_21637);
nand U22491 (N_22491,N_21054,N_21672);
xnor U22492 (N_22492,N_21167,N_21503);
or U22493 (N_22493,N_21723,N_21893);
nand U22494 (N_22494,N_21854,N_21041);
nor U22495 (N_22495,N_21212,N_21114);
nor U22496 (N_22496,N_21747,N_21617);
or U22497 (N_22497,N_21519,N_21678);
xor U22498 (N_22498,N_21290,N_21701);
or U22499 (N_22499,N_21341,N_21109);
xnor U22500 (N_22500,N_21499,N_21052);
and U22501 (N_22501,N_21616,N_21490);
xor U22502 (N_22502,N_21344,N_21129);
or U22503 (N_22503,N_21291,N_21816);
nand U22504 (N_22504,N_21930,N_21448);
xor U22505 (N_22505,N_21635,N_21363);
or U22506 (N_22506,N_21375,N_21706);
nand U22507 (N_22507,N_21236,N_21718);
nor U22508 (N_22508,N_21628,N_21688);
nor U22509 (N_22509,N_21195,N_21113);
nor U22510 (N_22510,N_21628,N_21591);
and U22511 (N_22511,N_21244,N_21228);
and U22512 (N_22512,N_21207,N_21448);
xnor U22513 (N_22513,N_21409,N_21951);
nor U22514 (N_22514,N_21884,N_21234);
nor U22515 (N_22515,N_21257,N_21115);
xor U22516 (N_22516,N_21572,N_21984);
nand U22517 (N_22517,N_21004,N_21167);
nand U22518 (N_22518,N_21565,N_21093);
xor U22519 (N_22519,N_21820,N_21723);
and U22520 (N_22520,N_21788,N_21565);
xnor U22521 (N_22521,N_21801,N_21316);
nor U22522 (N_22522,N_21362,N_21309);
and U22523 (N_22523,N_21722,N_21757);
and U22524 (N_22524,N_21053,N_21527);
nand U22525 (N_22525,N_21192,N_21775);
and U22526 (N_22526,N_21418,N_21478);
or U22527 (N_22527,N_21243,N_21675);
or U22528 (N_22528,N_21264,N_21780);
nand U22529 (N_22529,N_21805,N_21385);
or U22530 (N_22530,N_21311,N_21997);
and U22531 (N_22531,N_21790,N_21699);
xor U22532 (N_22532,N_21980,N_21859);
nand U22533 (N_22533,N_21283,N_21929);
nor U22534 (N_22534,N_21067,N_21737);
xnor U22535 (N_22535,N_21889,N_21129);
or U22536 (N_22536,N_21336,N_21775);
nor U22537 (N_22537,N_21681,N_21317);
and U22538 (N_22538,N_21187,N_21686);
xnor U22539 (N_22539,N_21068,N_21008);
nor U22540 (N_22540,N_21856,N_21273);
xor U22541 (N_22541,N_21764,N_21422);
nand U22542 (N_22542,N_21647,N_21518);
nor U22543 (N_22543,N_21069,N_21748);
or U22544 (N_22544,N_21530,N_21705);
xnor U22545 (N_22545,N_21654,N_21283);
or U22546 (N_22546,N_21440,N_21213);
and U22547 (N_22547,N_21258,N_21000);
or U22548 (N_22548,N_21501,N_21351);
xnor U22549 (N_22549,N_21462,N_21661);
nor U22550 (N_22550,N_21123,N_21486);
nor U22551 (N_22551,N_21113,N_21409);
or U22552 (N_22552,N_21966,N_21039);
and U22553 (N_22553,N_21823,N_21923);
or U22554 (N_22554,N_21424,N_21051);
and U22555 (N_22555,N_21836,N_21510);
nand U22556 (N_22556,N_21858,N_21535);
and U22557 (N_22557,N_21736,N_21084);
nor U22558 (N_22558,N_21768,N_21906);
xnor U22559 (N_22559,N_21330,N_21282);
nor U22560 (N_22560,N_21748,N_21571);
nand U22561 (N_22561,N_21213,N_21130);
nand U22562 (N_22562,N_21071,N_21472);
or U22563 (N_22563,N_21922,N_21563);
nand U22564 (N_22564,N_21328,N_21526);
xor U22565 (N_22565,N_21002,N_21125);
xnor U22566 (N_22566,N_21269,N_21690);
or U22567 (N_22567,N_21959,N_21817);
and U22568 (N_22568,N_21686,N_21263);
nand U22569 (N_22569,N_21783,N_21676);
xnor U22570 (N_22570,N_21707,N_21744);
and U22571 (N_22571,N_21471,N_21905);
xor U22572 (N_22572,N_21717,N_21522);
nand U22573 (N_22573,N_21771,N_21126);
nand U22574 (N_22574,N_21361,N_21351);
nand U22575 (N_22575,N_21995,N_21050);
and U22576 (N_22576,N_21620,N_21606);
nor U22577 (N_22577,N_21993,N_21313);
and U22578 (N_22578,N_21300,N_21454);
xor U22579 (N_22579,N_21482,N_21783);
and U22580 (N_22580,N_21173,N_21379);
nor U22581 (N_22581,N_21886,N_21806);
and U22582 (N_22582,N_21624,N_21580);
nand U22583 (N_22583,N_21919,N_21327);
or U22584 (N_22584,N_21751,N_21721);
xnor U22585 (N_22585,N_21228,N_21993);
nand U22586 (N_22586,N_21199,N_21175);
or U22587 (N_22587,N_21146,N_21561);
and U22588 (N_22588,N_21073,N_21791);
and U22589 (N_22589,N_21463,N_21540);
and U22590 (N_22590,N_21230,N_21556);
xnor U22591 (N_22591,N_21400,N_21153);
nand U22592 (N_22592,N_21667,N_21248);
xor U22593 (N_22593,N_21512,N_21148);
nand U22594 (N_22594,N_21638,N_21275);
xnor U22595 (N_22595,N_21606,N_21951);
nor U22596 (N_22596,N_21459,N_21290);
or U22597 (N_22597,N_21269,N_21202);
and U22598 (N_22598,N_21644,N_21480);
xnor U22599 (N_22599,N_21981,N_21528);
xnor U22600 (N_22600,N_21873,N_21946);
and U22601 (N_22601,N_21653,N_21462);
nand U22602 (N_22602,N_21160,N_21808);
or U22603 (N_22603,N_21028,N_21043);
xnor U22604 (N_22604,N_21732,N_21479);
xnor U22605 (N_22605,N_21068,N_21020);
and U22606 (N_22606,N_21080,N_21128);
xnor U22607 (N_22607,N_21237,N_21769);
and U22608 (N_22608,N_21736,N_21062);
and U22609 (N_22609,N_21918,N_21971);
xor U22610 (N_22610,N_21216,N_21625);
nor U22611 (N_22611,N_21114,N_21780);
and U22612 (N_22612,N_21519,N_21135);
or U22613 (N_22613,N_21986,N_21791);
or U22614 (N_22614,N_21151,N_21837);
or U22615 (N_22615,N_21003,N_21054);
nand U22616 (N_22616,N_21394,N_21678);
or U22617 (N_22617,N_21854,N_21919);
and U22618 (N_22618,N_21195,N_21262);
xnor U22619 (N_22619,N_21592,N_21911);
nor U22620 (N_22620,N_21642,N_21178);
xnor U22621 (N_22621,N_21214,N_21612);
nand U22622 (N_22622,N_21899,N_21447);
xnor U22623 (N_22623,N_21422,N_21502);
nor U22624 (N_22624,N_21380,N_21221);
or U22625 (N_22625,N_21138,N_21586);
nor U22626 (N_22626,N_21377,N_21223);
nand U22627 (N_22627,N_21988,N_21805);
nor U22628 (N_22628,N_21981,N_21375);
and U22629 (N_22629,N_21703,N_21716);
xor U22630 (N_22630,N_21422,N_21665);
nand U22631 (N_22631,N_21222,N_21798);
xor U22632 (N_22632,N_21962,N_21560);
xor U22633 (N_22633,N_21693,N_21889);
xor U22634 (N_22634,N_21847,N_21644);
or U22635 (N_22635,N_21044,N_21812);
nand U22636 (N_22636,N_21194,N_21014);
or U22637 (N_22637,N_21815,N_21205);
and U22638 (N_22638,N_21165,N_21147);
or U22639 (N_22639,N_21395,N_21707);
xor U22640 (N_22640,N_21336,N_21678);
nor U22641 (N_22641,N_21642,N_21573);
nor U22642 (N_22642,N_21824,N_21548);
and U22643 (N_22643,N_21940,N_21370);
xnor U22644 (N_22644,N_21940,N_21580);
nand U22645 (N_22645,N_21372,N_21834);
and U22646 (N_22646,N_21191,N_21635);
xor U22647 (N_22647,N_21442,N_21567);
xor U22648 (N_22648,N_21304,N_21348);
and U22649 (N_22649,N_21781,N_21716);
and U22650 (N_22650,N_21660,N_21860);
xnor U22651 (N_22651,N_21784,N_21033);
xnor U22652 (N_22652,N_21600,N_21720);
xor U22653 (N_22653,N_21600,N_21764);
nor U22654 (N_22654,N_21652,N_21667);
and U22655 (N_22655,N_21393,N_21701);
nand U22656 (N_22656,N_21540,N_21971);
or U22657 (N_22657,N_21176,N_21340);
and U22658 (N_22658,N_21355,N_21556);
or U22659 (N_22659,N_21589,N_21614);
nand U22660 (N_22660,N_21438,N_21442);
or U22661 (N_22661,N_21830,N_21723);
xor U22662 (N_22662,N_21725,N_21701);
nor U22663 (N_22663,N_21336,N_21401);
nand U22664 (N_22664,N_21075,N_21122);
xnor U22665 (N_22665,N_21232,N_21508);
and U22666 (N_22666,N_21353,N_21832);
nor U22667 (N_22667,N_21355,N_21605);
nand U22668 (N_22668,N_21863,N_21862);
nand U22669 (N_22669,N_21694,N_21878);
or U22670 (N_22670,N_21207,N_21642);
nand U22671 (N_22671,N_21498,N_21855);
and U22672 (N_22672,N_21896,N_21917);
nor U22673 (N_22673,N_21836,N_21978);
or U22674 (N_22674,N_21750,N_21396);
nand U22675 (N_22675,N_21003,N_21173);
or U22676 (N_22676,N_21367,N_21746);
nand U22677 (N_22677,N_21833,N_21634);
nor U22678 (N_22678,N_21828,N_21816);
xnor U22679 (N_22679,N_21961,N_21265);
xnor U22680 (N_22680,N_21924,N_21996);
or U22681 (N_22681,N_21159,N_21927);
nand U22682 (N_22682,N_21025,N_21310);
and U22683 (N_22683,N_21498,N_21784);
or U22684 (N_22684,N_21745,N_21054);
nand U22685 (N_22685,N_21130,N_21956);
or U22686 (N_22686,N_21269,N_21991);
nor U22687 (N_22687,N_21579,N_21913);
nand U22688 (N_22688,N_21990,N_21404);
xnor U22689 (N_22689,N_21853,N_21280);
nor U22690 (N_22690,N_21692,N_21927);
or U22691 (N_22691,N_21154,N_21756);
nor U22692 (N_22692,N_21065,N_21920);
nor U22693 (N_22693,N_21765,N_21695);
nand U22694 (N_22694,N_21883,N_21211);
or U22695 (N_22695,N_21855,N_21021);
nand U22696 (N_22696,N_21296,N_21867);
xnor U22697 (N_22697,N_21745,N_21998);
and U22698 (N_22698,N_21718,N_21128);
and U22699 (N_22699,N_21330,N_21933);
and U22700 (N_22700,N_21847,N_21451);
nand U22701 (N_22701,N_21023,N_21622);
nor U22702 (N_22702,N_21371,N_21960);
xor U22703 (N_22703,N_21317,N_21619);
or U22704 (N_22704,N_21781,N_21046);
nor U22705 (N_22705,N_21803,N_21134);
xnor U22706 (N_22706,N_21260,N_21397);
nand U22707 (N_22707,N_21033,N_21178);
nor U22708 (N_22708,N_21264,N_21844);
or U22709 (N_22709,N_21099,N_21404);
or U22710 (N_22710,N_21953,N_21899);
nand U22711 (N_22711,N_21786,N_21661);
xor U22712 (N_22712,N_21840,N_21439);
nand U22713 (N_22713,N_21810,N_21768);
xnor U22714 (N_22714,N_21362,N_21767);
or U22715 (N_22715,N_21764,N_21257);
nand U22716 (N_22716,N_21295,N_21020);
and U22717 (N_22717,N_21557,N_21714);
and U22718 (N_22718,N_21071,N_21413);
nand U22719 (N_22719,N_21880,N_21375);
xor U22720 (N_22720,N_21885,N_21878);
nor U22721 (N_22721,N_21097,N_21515);
and U22722 (N_22722,N_21455,N_21884);
or U22723 (N_22723,N_21163,N_21268);
nor U22724 (N_22724,N_21889,N_21078);
xnor U22725 (N_22725,N_21820,N_21270);
xor U22726 (N_22726,N_21204,N_21018);
and U22727 (N_22727,N_21713,N_21867);
and U22728 (N_22728,N_21184,N_21544);
nand U22729 (N_22729,N_21587,N_21521);
xor U22730 (N_22730,N_21651,N_21178);
xnor U22731 (N_22731,N_21027,N_21144);
and U22732 (N_22732,N_21200,N_21651);
xor U22733 (N_22733,N_21103,N_21710);
nand U22734 (N_22734,N_21666,N_21573);
xor U22735 (N_22735,N_21065,N_21734);
nand U22736 (N_22736,N_21817,N_21394);
nand U22737 (N_22737,N_21442,N_21713);
and U22738 (N_22738,N_21537,N_21208);
nand U22739 (N_22739,N_21106,N_21153);
xor U22740 (N_22740,N_21440,N_21651);
nand U22741 (N_22741,N_21901,N_21657);
nand U22742 (N_22742,N_21552,N_21429);
nor U22743 (N_22743,N_21580,N_21115);
nor U22744 (N_22744,N_21838,N_21328);
nor U22745 (N_22745,N_21704,N_21338);
nand U22746 (N_22746,N_21122,N_21209);
nor U22747 (N_22747,N_21740,N_21138);
xnor U22748 (N_22748,N_21835,N_21768);
nor U22749 (N_22749,N_21214,N_21557);
and U22750 (N_22750,N_21311,N_21415);
nor U22751 (N_22751,N_21557,N_21158);
and U22752 (N_22752,N_21705,N_21207);
nor U22753 (N_22753,N_21480,N_21502);
and U22754 (N_22754,N_21681,N_21313);
xor U22755 (N_22755,N_21514,N_21151);
nor U22756 (N_22756,N_21039,N_21999);
nor U22757 (N_22757,N_21980,N_21752);
and U22758 (N_22758,N_21549,N_21470);
and U22759 (N_22759,N_21079,N_21183);
xnor U22760 (N_22760,N_21287,N_21950);
nand U22761 (N_22761,N_21559,N_21035);
nor U22762 (N_22762,N_21034,N_21155);
nand U22763 (N_22763,N_21050,N_21192);
xor U22764 (N_22764,N_21134,N_21524);
xnor U22765 (N_22765,N_21166,N_21776);
nor U22766 (N_22766,N_21346,N_21463);
and U22767 (N_22767,N_21506,N_21805);
and U22768 (N_22768,N_21259,N_21750);
and U22769 (N_22769,N_21791,N_21655);
nor U22770 (N_22770,N_21799,N_21542);
xnor U22771 (N_22771,N_21030,N_21832);
xor U22772 (N_22772,N_21574,N_21612);
or U22773 (N_22773,N_21701,N_21812);
xor U22774 (N_22774,N_21967,N_21410);
or U22775 (N_22775,N_21198,N_21048);
and U22776 (N_22776,N_21927,N_21466);
nor U22777 (N_22777,N_21886,N_21683);
nor U22778 (N_22778,N_21844,N_21815);
or U22779 (N_22779,N_21186,N_21139);
nor U22780 (N_22780,N_21383,N_21619);
xnor U22781 (N_22781,N_21508,N_21820);
nand U22782 (N_22782,N_21339,N_21434);
or U22783 (N_22783,N_21757,N_21343);
xor U22784 (N_22784,N_21905,N_21444);
nor U22785 (N_22785,N_21794,N_21119);
nand U22786 (N_22786,N_21460,N_21772);
nor U22787 (N_22787,N_21057,N_21448);
or U22788 (N_22788,N_21576,N_21043);
and U22789 (N_22789,N_21564,N_21238);
and U22790 (N_22790,N_21167,N_21245);
xnor U22791 (N_22791,N_21416,N_21027);
nor U22792 (N_22792,N_21190,N_21120);
nand U22793 (N_22793,N_21437,N_21125);
or U22794 (N_22794,N_21440,N_21602);
nor U22795 (N_22795,N_21508,N_21304);
xor U22796 (N_22796,N_21940,N_21176);
xor U22797 (N_22797,N_21353,N_21849);
xnor U22798 (N_22798,N_21850,N_21367);
and U22799 (N_22799,N_21233,N_21900);
nor U22800 (N_22800,N_21045,N_21336);
nor U22801 (N_22801,N_21114,N_21708);
nor U22802 (N_22802,N_21281,N_21605);
or U22803 (N_22803,N_21830,N_21050);
nand U22804 (N_22804,N_21722,N_21184);
nor U22805 (N_22805,N_21403,N_21011);
nand U22806 (N_22806,N_21654,N_21134);
or U22807 (N_22807,N_21144,N_21498);
and U22808 (N_22808,N_21569,N_21391);
or U22809 (N_22809,N_21872,N_21037);
and U22810 (N_22810,N_21877,N_21411);
and U22811 (N_22811,N_21946,N_21862);
xor U22812 (N_22812,N_21979,N_21711);
xor U22813 (N_22813,N_21304,N_21091);
xnor U22814 (N_22814,N_21442,N_21147);
or U22815 (N_22815,N_21860,N_21643);
nand U22816 (N_22816,N_21055,N_21123);
and U22817 (N_22817,N_21960,N_21841);
xor U22818 (N_22818,N_21680,N_21212);
nand U22819 (N_22819,N_21758,N_21144);
nor U22820 (N_22820,N_21562,N_21147);
nor U22821 (N_22821,N_21246,N_21855);
xor U22822 (N_22822,N_21063,N_21612);
or U22823 (N_22823,N_21032,N_21471);
nand U22824 (N_22824,N_21033,N_21552);
nand U22825 (N_22825,N_21020,N_21198);
and U22826 (N_22826,N_21691,N_21726);
nand U22827 (N_22827,N_21119,N_21932);
and U22828 (N_22828,N_21644,N_21013);
or U22829 (N_22829,N_21445,N_21930);
and U22830 (N_22830,N_21252,N_21949);
or U22831 (N_22831,N_21223,N_21010);
and U22832 (N_22832,N_21089,N_21686);
or U22833 (N_22833,N_21077,N_21702);
xnor U22834 (N_22834,N_21111,N_21566);
nor U22835 (N_22835,N_21265,N_21866);
nand U22836 (N_22836,N_21533,N_21626);
nor U22837 (N_22837,N_21141,N_21335);
and U22838 (N_22838,N_21397,N_21023);
nor U22839 (N_22839,N_21586,N_21036);
xor U22840 (N_22840,N_21391,N_21396);
nand U22841 (N_22841,N_21072,N_21564);
or U22842 (N_22842,N_21981,N_21163);
xnor U22843 (N_22843,N_21755,N_21275);
xor U22844 (N_22844,N_21595,N_21919);
nand U22845 (N_22845,N_21719,N_21292);
xor U22846 (N_22846,N_21085,N_21385);
or U22847 (N_22847,N_21834,N_21522);
or U22848 (N_22848,N_21873,N_21935);
xnor U22849 (N_22849,N_21316,N_21983);
and U22850 (N_22850,N_21575,N_21199);
nor U22851 (N_22851,N_21816,N_21621);
nand U22852 (N_22852,N_21580,N_21076);
nor U22853 (N_22853,N_21982,N_21485);
and U22854 (N_22854,N_21041,N_21129);
nor U22855 (N_22855,N_21130,N_21449);
or U22856 (N_22856,N_21326,N_21386);
and U22857 (N_22857,N_21767,N_21819);
and U22858 (N_22858,N_21008,N_21729);
and U22859 (N_22859,N_21324,N_21318);
or U22860 (N_22860,N_21533,N_21035);
nor U22861 (N_22861,N_21468,N_21311);
and U22862 (N_22862,N_21951,N_21097);
or U22863 (N_22863,N_21819,N_21800);
nand U22864 (N_22864,N_21391,N_21394);
xnor U22865 (N_22865,N_21394,N_21182);
nor U22866 (N_22866,N_21637,N_21947);
xor U22867 (N_22867,N_21183,N_21077);
and U22868 (N_22868,N_21958,N_21608);
or U22869 (N_22869,N_21665,N_21246);
xor U22870 (N_22870,N_21474,N_21580);
nor U22871 (N_22871,N_21270,N_21953);
nand U22872 (N_22872,N_21974,N_21986);
nor U22873 (N_22873,N_21328,N_21377);
nand U22874 (N_22874,N_21116,N_21856);
nand U22875 (N_22875,N_21518,N_21941);
xor U22876 (N_22876,N_21834,N_21810);
nand U22877 (N_22877,N_21504,N_21929);
and U22878 (N_22878,N_21032,N_21505);
or U22879 (N_22879,N_21014,N_21407);
and U22880 (N_22880,N_21880,N_21175);
xor U22881 (N_22881,N_21618,N_21505);
nand U22882 (N_22882,N_21163,N_21707);
xor U22883 (N_22883,N_21541,N_21124);
and U22884 (N_22884,N_21602,N_21172);
nand U22885 (N_22885,N_21079,N_21615);
and U22886 (N_22886,N_21744,N_21328);
nor U22887 (N_22887,N_21037,N_21811);
nand U22888 (N_22888,N_21991,N_21304);
and U22889 (N_22889,N_21749,N_21141);
or U22890 (N_22890,N_21689,N_21516);
or U22891 (N_22891,N_21891,N_21210);
or U22892 (N_22892,N_21587,N_21081);
or U22893 (N_22893,N_21910,N_21785);
nor U22894 (N_22894,N_21422,N_21609);
xnor U22895 (N_22895,N_21039,N_21033);
and U22896 (N_22896,N_21780,N_21875);
nand U22897 (N_22897,N_21985,N_21301);
nor U22898 (N_22898,N_21098,N_21235);
xor U22899 (N_22899,N_21371,N_21743);
xor U22900 (N_22900,N_21016,N_21973);
nor U22901 (N_22901,N_21644,N_21869);
and U22902 (N_22902,N_21700,N_21456);
nor U22903 (N_22903,N_21487,N_21342);
nand U22904 (N_22904,N_21022,N_21708);
nor U22905 (N_22905,N_21619,N_21446);
or U22906 (N_22906,N_21961,N_21484);
xor U22907 (N_22907,N_21442,N_21253);
xnor U22908 (N_22908,N_21278,N_21392);
or U22909 (N_22909,N_21073,N_21747);
nand U22910 (N_22910,N_21774,N_21090);
nand U22911 (N_22911,N_21101,N_21936);
nor U22912 (N_22912,N_21005,N_21597);
xnor U22913 (N_22913,N_21240,N_21104);
nand U22914 (N_22914,N_21526,N_21225);
nor U22915 (N_22915,N_21287,N_21007);
nand U22916 (N_22916,N_21357,N_21472);
nor U22917 (N_22917,N_21332,N_21138);
or U22918 (N_22918,N_21645,N_21509);
nor U22919 (N_22919,N_21746,N_21193);
xnor U22920 (N_22920,N_21532,N_21018);
xnor U22921 (N_22921,N_21270,N_21825);
or U22922 (N_22922,N_21425,N_21261);
nor U22923 (N_22923,N_21322,N_21965);
nor U22924 (N_22924,N_21626,N_21231);
xor U22925 (N_22925,N_21186,N_21009);
xor U22926 (N_22926,N_21942,N_21711);
nor U22927 (N_22927,N_21806,N_21523);
and U22928 (N_22928,N_21838,N_21312);
nor U22929 (N_22929,N_21848,N_21592);
nand U22930 (N_22930,N_21653,N_21293);
and U22931 (N_22931,N_21539,N_21280);
nand U22932 (N_22932,N_21834,N_21644);
nand U22933 (N_22933,N_21760,N_21791);
and U22934 (N_22934,N_21878,N_21019);
nand U22935 (N_22935,N_21823,N_21970);
nor U22936 (N_22936,N_21356,N_21999);
nor U22937 (N_22937,N_21605,N_21854);
xnor U22938 (N_22938,N_21715,N_21634);
or U22939 (N_22939,N_21883,N_21395);
nor U22940 (N_22940,N_21541,N_21356);
nand U22941 (N_22941,N_21654,N_21053);
nor U22942 (N_22942,N_21563,N_21731);
xnor U22943 (N_22943,N_21887,N_21667);
xnor U22944 (N_22944,N_21138,N_21300);
nand U22945 (N_22945,N_21074,N_21480);
or U22946 (N_22946,N_21555,N_21299);
or U22947 (N_22947,N_21947,N_21000);
nor U22948 (N_22948,N_21762,N_21270);
and U22949 (N_22949,N_21142,N_21489);
nor U22950 (N_22950,N_21262,N_21823);
or U22951 (N_22951,N_21874,N_21771);
or U22952 (N_22952,N_21836,N_21388);
and U22953 (N_22953,N_21232,N_21616);
or U22954 (N_22954,N_21284,N_21422);
xor U22955 (N_22955,N_21571,N_21562);
nor U22956 (N_22956,N_21217,N_21458);
nor U22957 (N_22957,N_21899,N_21426);
or U22958 (N_22958,N_21674,N_21848);
xor U22959 (N_22959,N_21707,N_21907);
or U22960 (N_22960,N_21523,N_21092);
xnor U22961 (N_22961,N_21714,N_21146);
xor U22962 (N_22962,N_21102,N_21352);
xor U22963 (N_22963,N_21960,N_21204);
nor U22964 (N_22964,N_21618,N_21609);
xnor U22965 (N_22965,N_21541,N_21293);
and U22966 (N_22966,N_21385,N_21549);
and U22967 (N_22967,N_21477,N_21653);
and U22968 (N_22968,N_21101,N_21843);
or U22969 (N_22969,N_21112,N_21425);
nand U22970 (N_22970,N_21265,N_21433);
nand U22971 (N_22971,N_21552,N_21549);
or U22972 (N_22972,N_21630,N_21506);
nor U22973 (N_22973,N_21090,N_21534);
nand U22974 (N_22974,N_21297,N_21170);
xnor U22975 (N_22975,N_21972,N_21281);
or U22976 (N_22976,N_21516,N_21903);
nor U22977 (N_22977,N_21303,N_21826);
or U22978 (N_22978,N_21608,N_21164);
nand U22979 (N_22979,N_21828,N_21325);
or U22980 (N_22980,N_21167,N_21439);
or U22981 (N_22981,N_21652,N_21152);
or U22982 (N_22982,N_21850,N_21600);
nand U22983 (N_22983,N_21831,N_21688);
and U22984 (N_22984,N_21850,N_21585);
or U22985 (N_22985,N_21797,N_21702);
nor U22986 (N_22986,N_21671,N_21259);
or U22987 (N_22987,N_21363,N_21711);
xnor U22988 (N_22988,N_21415,N_21510);
xor U22989 (N_22989,N_21079,N_21407);
and U22990 (N_22990,N_21414,N_21005);
nand U22991 (N_22991,N_21382,N_21344);
nand U22992 (N_22992,N_21046,N_21622);
nor U22993 (N_22993,N_21522,N_21876);
nand U22994 (N_22994,N_21590,N_21690);
and U22995 (N_22995,N_21442,N_21069);
nand U22996 (N_22996,N_21867,N_21657);
and U22997 (N_22997,N_21311,N_21668);
or U22998 (N_22998,N_21656,N_21155);
nand U22999 (N_22999,N_21235,N_21295);
nor U23000 (N_23000,N_22737,N_22193);
nand U23001 (N_23001,N_22087,N_22186);
or U23002 (N_23002,N_22105,N_22360);
nand U23003 (N_23003,N_22464,N_22147);
xnor U23004 (N_23004,N_22916,N_22381);
and U23005 (N_23005,N_22316,N_22576);
nand U23006 (N_23006,N_22937,N_22945);
or U23007 (N_23007,N_22942,N_22514);
or U23008 (N_23008,N_22382,N_22770);
nor U23009 (N_23009,N_22660,N_22048);
xor U23010 (N_23010,N_22260,N_22228);
xor U23011 (N_23011,N_22149,N_22855);
nor U23012 (N_23012,N_22818,N_22593);
and U23013 (N_23013,N_22842,N_22136);
xnor U23014 (N_23014,N_22627,N_22182);
and U23015 (N_23015,N_22983,N_22556);
or U23016 (N_23016,N_22056,N_22095);
xor U23017 (N_23017,N_22534,N_22812);
nand U23018 (N_23018,N_22040,N_22807);
nand U23019 (N_23019,N_22749,N_22046);
or U23020 (N_23020,N_22229,N_22938);
xor U23021 (N_23021,N_22718,N_22947);
xnor U23022 (N_23022,N_22396,N_22751);
and U23023 (N_23023,N_22490,N_22117);
nand U23024 (N_23024,N_22765,N_22376);
and U23025 (N_23025,N_22476,N_22816);
and U23026 (N_23026,N_22634,N_22240);
and U23027 (N_23027,N_22791,N_22680);
xor U23028 (N_23028,N_22391,N_22478);
nor U23029 (N_23029,N_22120,N_22851);
or U23030 (N_23030,N_22298,N_22010);
or U23031 (N_23031,N_22601,N_22743);
xnor U23032 (N_23032,N_22652,N_22832);
or U23033 (N_23033,N_22263,N_22439);
nor U23034 (N_23034,N_22764,N_22038);
nand U23035 (N_23035,N_22503,N_22753);
and U23036 (N_23036,N_22370,N_22379);
or U23037 (N_23037,N_22787,N_22954);
nand U23038 (N_23038,N_22472,N_22362);
and U23039 (N_23039,N_22355,N_22258);
nand U23040 (N_23040,N_22070,N_22953);
nand U23041 (N_23041,N_22910,N_22375);
nor U23042 (N_23042,N_22421,N_22869);
xnor U23043 (N_23043,N_22694,N_22768);
nor U23044 (N_23044,N_22326,N_22191);
xor U23045 (N_23045,N_22663,N_22343);
or U23046 (N_23046,N_22825,N_22259);
or U23047 (N_23047,N_22469,N_22517);
and U23048 (N_23048,N_22371,N_22051);
xor U23049 (N_23049,N_22313,N_22559);
or U23050 (N_23050,N_22779,N_22889);
or U23051 (N_23051,N_22044,N_22146);
nor U23052 (N_23052,N_22011,N_22133);
nand U23053 (N_23053,N_22958,N_22032);
nand U23054 (N_23054,N_22819,N_22976);
nand U23055 (N_23055,N_22359,N_22446);
and U23056 (N_23056,N_22303,N_22811);
or U23057 (N_23057,N_22346,N_22693);
nor U23058 (N_23058,N_22001,N_22425);
nand U23059 (N_23059,N_22773,N_22473);
and U23060 (N_23060,N_22860,N_22985);
nand U23061 (N_23061,N_22158,N_22813);
nand U23062 (N_23062,N_22932,N_22555);
and U23063 (N_23063,N_22873,N_22658);
or U23064 (N_23064,N_22533,N_22792);
nand U23065 (N_23065,N_22602,N_22466);
or U23066 (N_23066,N_22447,N_22703);
nor U23067 (N_23067,N_22069,N_22404);
xnor U23068 (N_23068,N_22318,N_22744);
and U23069 (N_23069,N_22453,N_22670);
xnor U23070 (N_23070,N_22605,N_22285);
nor U23071 (N_23071,N_22296,N_22076);
xor U23072 (N_23072,N_22500,N_22969);
nor U23073 (N_23073,N_22831,N_22590);
nor U23074 (N_23074,N_22524,N_22757);
xnor U23075 (N_23075,N_22748,N_22308);
nor U23076 (N_23076,N_22383,N_22736);
nor U23077 (N_23077,N_22868,N_22102);
and U23078 (N_23078,N_22767,N_22913);
xor U23079 (N_23079,N_22920,N_22642);
nand U23080 (N_23080,N_22618,N_22635);
nand U23081 (N_23081,N_22717,N_22426);
or U23082 (N_23082,N_22054,N_22962);
xnor U23083 (N_23083,N_22554,N_22215);
xor U23084 (N_23084,N_22975,N_22072);
or U23085 (N_23085,N_22012,N_22934);
xor U23086 (N_23086,N_22584,N_22281);
xnor U23087 (N_23087,N_22894,N_22861);
xor U23088 (N_23088,N_22689,N_22110);
nor U23089 (N_23089,N_22544,N_22665);
nand U23090 (N_23090,N_22678,N_22294);
nor U23091 (N_23091,N_22314,N_22759);
nand U23092 (N_23092,N_22543,N_22883);
or U23093 (N_23093,N_22875,N_22045);
nor U23094 (N_23094,N_22836,N_22804);
and U23095 (N_23095,N_22239,N_22331);
nand U23096 (N_23096,N_22594,N_22939);
nand U23097 (N_23097,N_22327,N_22397);
and U23098 (N_23098,N_22495,N_22135);
and U23099 (N_23099,N_22457,N_22998);
and U23100 (N_23100,N_22290,N_22906);
and U23101 (N_23101,N_22852,N_22725);
nand U23102 (N_23102,N_22488,N_22848);
or U23103 (N_23103,N_22882,N_22980);
nand U23104 (N_23104,N_22282,N_22427);
nand U23105 (N_23105,N_22334,N_22774);
and U23106 (N_23106,N_22574,N_22650);
or U23107 (N_23107,N_22866,N_22399);
and U23108 (N_23108,N_22406,N_22292);
or U23109 (N_23109,N_22510,N_22518);
nand U23110 (N_23110,N_22793,N_22025);
or U23111 (N_23111,N_22946,N_22442);
xor U23112 (N_23112,N_22093,N_22429);
nor U23113 (N_23113,N_22086,N_22890);
or U23114 (N_23114,N_22777,N_22622);
or U23115 (N_23115,N_22254,N_22164);
xnor U23116 (N_23116,N_22050,N_22460);
xnor U23117 (N_23117,N_22161,N_22651);
nand U23118 (N_23118,N_22731,N_22413);
nor U23119 (N_23119,N_22871,N_22287);
and U23120 (N_23120,N_22888,N_22328);
or U23121 (N_23121,N_22487,N_22052);
or U23122 (N_23122,N_22530,N_22219);
nor U23123 (N_23123,N_22116,N_22322);
nand U23124 (N_23124,N_22702,N_22896);
and U23125 (N_23125,N_22539,N_22711);
nand U23126 (N_23126,N_22841,N_22157);
and U23127 (N_23127,N_22676,N_22756);
and U23128 (N_23128,N_22177,N_22121);
xor U23129 (N_23129,N_22267,N_22585);
nor U23130 (N_23130,N_22168,N_22310);
nor U23131 (N_23131,N_22837,N_22029);
and U23132 (N_23132,N_22206,N_22919);
nor U23133 (N_23133,N_22423,N_22808);
nand U23134 (N_23134,N_22424,N_22190);
nor U23135 (N_23135,N_22870,N_22451);
and U23136 (N_23136,N_22188,N_22907);
or U23137 (N_23137,N_22448,N_22276);
nand U23138 (N_23138,N_22918,N_22643);
or U23139 (N_23139,N_22794,N_22948);
nand U23140 (N_23140,N_22609,N_22293);
nand U23141 (N_23141,N_22220,N_22972);
or U23142 (N_23142,N_22659,N_22769);
and U23143 (N_23143,N_22151,N_22390);
or U23144 (N_23144,N_22686,N_22562);
nand U23145 (N_23145,N_22492,N_22245);
and U23146 (N_23146,N_22874,N_22925);
nor U23147 (N_23147,N_22705,N_22535);
nor U23148 (N_23148,N_22115,N_22415);
nand U23149 (N_23149,N_22595,N_22986);
xor U23150 (N_23150,N_22741,N_22823);
xnor U23151 (N_23151,N_22187,N_22824);
and U23152 (N_23152,N_22776,N_22089);
and U23153 (N_23153,N_22529,N_22775);
nor U23154 (N_23154,N_22781,N_22030);
and U23155 (N_23155,N_22257,N_22822);
and U23156 (N_23156,N_22859,N_22019);
nand U23157 (N_23157,N_22083,N_22144);
nor U23158 (N_23158,N_22600,N_22134);
nand U23159 (N_23159,N_22638,N_22927);
nor U23160 (N_23160,N_22653,N_22657);
xor U23161 (N_23161,N_22885,N_22410);
or U23162 (N_23162,N_22210,N_22007);
and U23163 (N_23163,N_22003,N_22984);
xnor U23164 (N_23164,N_22691,N_22536);
nor U23165 (N_23165,N_22389,N_22977);
or U23166 (N_23166,N_22491,N_22905);
and U23167 (N_23167,N_22204,N_22604);
nand U23168 (N_23168,N_22628,N_22027);
nand U23169 (N_23169,N_22037,N_22450);
nand U23170 (N_23170,N_22968,N_22912);
nor U23171 (N_23171,N_22815,N_22286);
nand U23172 (N_23172,N_22955,N_22911);
and U23173 (N_23173,N_22251,N_22277);
or U23174 (N_23174,N_22881,N_22671);
xor U23175 (N_23175,N_22988,N_22364);
xor U23176 (N_23176,N_22935,N_22053);
nor U23177 (N_23177,N_22057,N_22026);
xnor U23178 (N_23178,N_22903,N_22828);
nor U23179 (N_23179,N_22138,N_22728);
nor U23180 (N_23180,N_22648,N_22356);
and U23181 (N_23181,N_22299,N_22512);
or U23182 (N_23182,N_22632,N_22253);
xor U23183 (N_23183,N_22598,N_22797);
or U23184 (N_23184,N_22821,N_22546);
nor U23185 (N_23185,N_22696,N_22682);
nand U23186 (N_23186,N_22091,N_22724);
nor U23187 (N_23187,N_22944,N_22493);
nand U23188 (N_23188,N_22256,N_22952);
and U23189 (N_23189,N_22727,N_22617);
nor U23190 (N_23190,N_22119,N_22931);
nand U23191 (N_23191,N_22713,N_22437);
nand U23192 (N_23192,N_22471,N_22235);
nor U23193 (N_23193,N_22319,N_22175);
or U23194 (N_23194,N_22847,N_22137);
xnor U23195 (N_23195,N_22372,N_22486);
nor U23196 (N_23196,N_22675,N_22461);
xnor U23197 (N_23197,N_22683,N_22084);
nor U23198 (N_23198,N_22607,N_22378);
and U23199 (N_23199,N_22479,N_22009);
nor U23200 (N_23200,N_22068,N_22035);
nand U23201 (N_23201,N_22320,N_22170);
or U23202 (N_23202,N_22538,N_22747);
nor U23203 (N_23203,N_22152,N_22506);
nor U23204 (N_23204,N_22475,N_22306);
or U23205 (N_23205,N_22892,N_22042);
and U23206 (N_23206,N_22090,N_22879);
and U23207 (N_23207,N_22407,N_22330);
nand U23208 (N_23208,N_22982,N_22189);
xor U23209 (N_23209,N_22459,N_22649);
nor U23210 (N_23210,N_22402,N_22950);
and U23211 (N_23211,N_22470,N_22197);
or U23212 (N_23212,N_22557,N_22365);
xnor U23213 (N_23213,N_22722,N_22750);
xnor U23214 (N_23214,N_22698,N_22181);
nand U23215 (N_23215,N_22688,N_22405);
xor U23216 (N_23216,N_22560,N_22814);
nor U23217 (N_23217,N_22126,N_22021);
nor U23218 (N_23218,N_22926,N_22092);
and U23219 (N_23219,N_22000,N_22625);
nand U23220 (N_23220,N_22047,N_22978);
and U23221 (N_23221,N_22224,N_22008);
nor U23222 (N_23222,N_22681,N_22291);
nand U23223 (N_23223,N_22194,N_22071);
nor U23224 (N_23224,N_22352,N_22344);
or U23225 (N_23225,N_22013,N_22833);
xnor U23226 (N_23226,N_22278,N_22930);
nor U23227 (N_23227,N_22107,N_22522);
or U23228 (N_23228,N_22246,N_22261);
and U23229 (N_23229,N_22845,N_22513);
nor U23230 (N_23230,N_22033,N_22249);
nor U23231 (N_23231,N_22416,N_22179);
nor U23232 (N_23232,N_22097,N_22521);
xnor U23233 (N_23233,N_22531,N_22943);
xor U23234 (N_23234,N_22567,N_22353);
xnor U23235 (N_23235,N_22564,N_22184);
nor U23236 (N_23236,N_22264,N_22205);
or U23237 (N_23237,N_22225,N_22826);
nor U23238 (N_23238,N_22166,N_22760);
nor U23239 (N_23239,N_22865,N_22898);
xor U23240 (N_23240,N_22283,N_22080);
or U23241 (N_23241,N_22430,N_22171);
or U23242 (N_23242,N_22202,N_22803);
nand U23243 (N_23243,N_22398,N_22250);
nor U23244 (N_23244,N_22165,N_22839);
and U23245 (N_23245,N_22374,N_22991);
and U23246 (N_23246,N_22242,N_22348);
and U23247 (N_23247,N_22351,N_22150);
and U23248 (N_23248,N_22637,N_22148);
or U23249 (N_23249,N_22055,N_22674);
or U23250 (N_23250,N_22667,N_22746);
or U23251 (N_23251,N_22238,N_22685);
xnor U23252 (N_23252,N_22163,N_22965);
and U23253 (N_23253,N_22417,N_22963);
xor U23254 (N_23254,N_22730,N_22212);
and U23255 (N_23255,N_22369,N_22106);
nand U23256 (N_23256,N_22458,N_22311);
nor U23257 (N_23257,N_22065,N_22124);
or U23258 (N_23258,N_22856,N_22248);
and U23259 (N_23259,N_22199,N_22961);
nand U23260 (N_23260,N_22656,N_22272);
or U23261 (N_23261,N_22715,N_22673);
xor U23262 (N_23262,N_22237,N_22266);
nand U23263 (N_23263,N_22307,N_22908);
xnor U23264 (N_23264,N_22411,N_22432);
nor U23265 (N_23265,N_22599,N_22373);
or U23266 (N_23266,N_22668,N_22462);
nor U23267 (N_23267,N_22393,N_22226);
nand U23268 (N_23268,N_22018,N_22886);
nor U23269 (N_23269,N_22695,N_22716);
nor U23270 (N_23270,N_22332,N_22922);
or U23271 (N_23271,N_22213,N_22017);
or U23272 (N_23272,N_22572,N_22143);
and U23273 (N_23273,N_22154,N_22796);
xor U23274 (N_23274,N_22735,N_22173);
or U23275 (N_23275,N_22209,N_22569);
or U23276 (N_23276,N_22496,N_22850);
nand U23277 (N_23277,N_22477,N_22853);
nor U23278 (N_23278,N_22484,N_22341);
nand U23279 (N_23279,N_22094,N_22336);
or U23280 (N_23280,N_22960,N_22999);
xnor U23281 (N_23281,N_22720,N_22145);
xor U23282 (N_23282,N_22004,N_22100);
or U23283 (N_23283,N_22880,N_22200);
or U23284 (N_23284,N_22337,N_22243);
or U23285 (N_23285,N_22854,N_22591);
nand U23286 (N_23286,N_22541,N_22645);
and U23287 (N_23287,N_22707,N_22626);
or U23288 (N_23288,N_22615,N_22766);
xor U23289 (N_23289,N_22483,N_22553);
xor U23290 (N_23290,N_22414,N_22772);
nor U23291 (N_23291,N_22849,N_22444);
or U23292 (N_23292,N_22697,N_22449);
or U23293 (N_23293,N_22024,N_22131);
or U23294 (N_23294,N_22981,N_22552);
and U23295 (N_23295,N_22159,N_22515);
or U23296 (N_23296,N_22914,N_22629);
xor U23297 (N_23297,N_22621,N_22754);
xnor U23298 (N_23298,N_22509,N_22827);
or U23299 (N_23299,N_22494,N_22997);
nand U23300 (N_23300,N_22167,N_22203);
or U23301 (N_23301,N_22074,N_22269);
or U23302 (N_23302,N_22734,N_22661);
xor U23303 (N_23303,N_22059,N_22109);
or U23304 (N_23304,N_22993,N_22139);
nor U23305 (N_23305,N_22505,N_22403);
nand U23306 (N_23306,N_22511,N_22581);
and U23307 (N_23307,N_22122,N_22185);
nand U23308 (N_23308,N_22992,N_22247);
nand U23309 (N_23309,N_22474,N_22214);
xnor U23310 (N_23310,N_22422,N_22577);
nand U23311 (N_23311,N_22377,N_22786);
or U23312 (N_23312,N_22540,N_22028);
and U23313 (N_23313,N_22596,N_22840);
xor U23314 (N_23314,N_22669,N_22664);
nor U23315 (N_23315,N_22198,N_22394);
and U23316 (N_23316,N_22778,N_22006);
xnor U23317 (N_23317,N_22350,N_22140);
nand U23318 (N_23318,N_22295,N_22358);
nand U23319 (N_23319,N_22289,N_22435);
and U23320 (N_23320,N_22366,N_22844);
and U23321 (N_23321,N_22740,N_22232);
xnor U23322 (N_23322,N_22526,N_22989);
or U23323 (N_23323,N_22049,N_22565);
xor U23324 (N_23324,N_22739,N_22408);
nand U23325 (N_23325,N_22582,N_22901);
xnor U23326 (N_23326,N_22113,N_22606);
xnor U23327 (N_23327,N_22709,N_22915);
nor U23328 (N_23328,N_22798,N_22957);
nand U23329 (N_23329,N_22275,N_22592);
xor U23330 (N_23330,N_22789,N_22465);
or U23331 (N_23331,N_22301,N_22317);
and U23332 (N_23332,N_22802,N_22959);
nor U23333 (N_23333,N_22523,N_22867);
or U23334 (N_23334,N_22795,N_22633);
nand U23335 (N_23335,N_22485,N_22636);
nor U23336 (N_23336,N_22620,N_22088);
xnor U23337 (N_23337,N_22380,N_22118);
xor U23338 (N_23338,N_22532,N_22129);
and U23339 (N_23339,N_22994,N_22838);
nand U23340 (N_23340,N_22979,N_22647);
xnor U23341 (N_23341,N_22271,N_22112);
nor U23342 (N_23342,N_22297,N_22501);
xor U23343 (N_23343,N_22079,N_22733);
and U23344 (N_23344,N_22395,N_22917);
nand U23345 (N_23345,N_22103,N_22800);
nand U23346 (N_23346,N_22436,N_22611);
or U23347 (N_23347,N_22265,N_22085);
nand U23348 (N_23348,N_22412,N_22846);
and U23349 (N_23349,N_22909,N_22160);
nand U23350 (N_23350,N_22893,N_22304);
xnor U23351 (N_23351,N_22973,N_22454);
nand U23352 (N_23352,N_22809,N_22520);
and U23353 (N_23353,N_22216,N_22153);
xnor U23354 (N_23354,N_22690,N_22801);
and U23355 (N_23355,N_22762,N_22575);
or U23356 (N_23356,N_22700,N_22387);
or U23357 (N_23357,N_22340,N_22923);
xor U23358 (N_23358,N_22099,N_22921);
xnor U23359 (N_23359,N_22573,N_22843);
or U23360 (N_23360,N_22252,N_22699);
and U23361 (N_23361,N_22111,N_22612);
nand U23362 (N_23362,N_22002,N_22714);
or U23363 (N_23363,N_22418,N_22878);
xor U23364 (N_23364,N_22640,N_22234);
and U23365 (N_23365,N_22624,N_22964);
nor U23366 (N_23366,N_22672,N_22654);
and U23367 (N_23367,N_22876,N_22467);
nor U23368 (N_23368,N_22528,N_22587);
nand U23369 (N_23369,N_22400,N_22335);
and U23370 (N_23370,N_22174,N_22745);
or U23371 (N_23371,N_22858,N_22208);
or U23372 (N_23372,N_22178,N_22349);
xor U23373 (N_23373,N_22077,N_22971);
nand U23374 (N_23374,N_22223,N_22211);
or U23375 (N_23375,N_22949,N_22504);
or U23376 (N_23376,N_22244,N_22455);
nand U23377 (N_23377,N_22201,N_22098);
nor U23378 (N_23378,N_22262,N_22877);
xnor U23379 (N_23379,N_22101,N_22790);
nor U23380 (N_23380,N_22928,N_22639);
or U23381 (N_23381,N_22578,N_22233);
or U23382 (N_23382,N_22062,N_22619);
xor U23383 (N_23383,N_22031,N_22005);
nor U23384 (N_23384,N_22280,N_22441);
xor U23385 (N_23385,N_22338,N_22970);
xnor U23386 (N_23386,N_22561,N_22900);
or U23387 (N_23387,N_22563,N_22060);
or U23388 (N_23388,N_22217,N_22367);
and U23389 (N_23389,N_22630,N_22064);
nor U23390 (N_23390,N_22603,N_22176);
and U23391 (N_23391,N_22545,N_22662);
xor U23392 (N_23392,N_22114,N_22579);
nand U23393 (N_23393,N_22571,N_22712);
or U23394 (N_23394,N_22388,N_22684);
nor U23395 (N_23395,N_22058,N_22502);
xnor U23396 (N_23396,N_22785,N_22066);
xnor U23397 (N_23397,N_22566,N_22274);
and U23398 (N_23398,N_22279,N_22752);
or U23399 (N_23399,N_22073,N_22468);
nor U23400 (N_23400,N_22361,N_22897);
nor U23401 (N_23401,N_22255,N_22169);
nor U23402 (N_23402,N_22723,N_22996);
and U23403 (N_23403,N_22445,N_22610);
xor U23404 (N_23404,N_22456,N_22863);
nand U23405 (N_23405,N_22570,N_22721);
nor U23406 (N_23406,N_22550,N_22156);
xnor U23407 (N_23407,N_22940,N_22273);
or U23408 (N_23408,N_22872,N_22616);
nor U23409 (N_23409,N_22132,N_22096);
or U23410 (N_23410,N_22480,N_22321);
nand U23411 (N_23411,N_22155,N_22799);
nor U23412 (N_23412,N_22784,N_22589);
nor U23413 (N_23413,N_22368,N_22829);
nor U23414 (N_23414,N_22222,N_22288);
nor U23415 (N_23415,N_22312,N_22710);
nand U23416 (N_23416,N_22221,N_22130);
or U23417 (N_23417,N_22580,N_22241);
or U23418 (N_23418,N_22036,N_22782);
or U23419 (N_23419,N_22284,N_22041);
nand U23420 (N_23420,N_22558,N_22666);
nand U23421 (N_23421,N_22420,N_22864);
xor U23422 (N_23422,N_22428,N_22196);
or U23423 (N_23423,N_22519,N_22974);
and U23424 (N_23424,N_22392,N_22172);
nand U23425 (N_23425,N_22990,N_22904);
or U23426 (N_23426,N_22527,N_22995);
nor U23427 (N_23427,N_22758,N_22409);
or U23428 (N_23428,N_22588,N_22891);
and U23429 (N_23429,N_22401,N_22127);
xor U23430 (N_23430,N_22902,N_22333);
xnor U23431 (N_23431,N_22315,N_22951);
xor U23432 (N_23432,N_22679,N_22499);
nand U23433 (N_23433,N_22386,N_22763);
or U23434 (N_23434,N_22452,N_22780);
or U23435 (N_23435,N_22329,N_22507);
or U23436 (N_23436,N_22440,N_22726);
and U23437 (N_23437,N_22967,N_22419);
nand U23438 (N_23438,N_22236,N_22497);
and U23439 (N_23439,N_22270,N_22817);
nand U23440 (N_23440,N_22738,N_22956);
nand U23441 (N_23441,N_22623,N_22887);
nor U23442 (N_23442,N_22641,N_22342);
xnor U23443 (N_23443,N_22783,N_22933);
and U23444 (N_23444,N_22463,N_22613);
xor U23445 (N_23445,N_22324,N_22755);
or U23446 (N_23446,N_22104,N_22646);
xor U23447 (N_23447,N_22325,N_22692);
xor U23448 (N_23448,N_22732,N_22309);
or U23449 (N_23449,N_22719,N_22551);
or U23450 (N_23450,N_22482,N_22183);
nor U23451 (N_23451,N_22128,N_22195);
nor U23452 (N_23452,N_22583,N_22300);
nand U23453 (N_23453,N_22061,N_22742);
and U23454 (N_23454,N_22125,N_22548);
or U23455 (N_23455,N_22302,N_22227);
and U23456 (N_23456,N_22108,N_22078);
nand U23457 (N_23457,N_22385,N_22677);
and U23458 (N_23458,N_22941,N_22363);
nand U23459 (N_23459,N_22162,N_22537);
nor U23460 (N_23460,N_22433,N_22434);
and U23461 (N_23461,N_22016,N_22857);
or U23462 (N_23462,N_22542,N_22644);
or U23463 (N_23463,N_22384,N_22023);
and U23464 (N_23464,N_22708,N_22525);
nand U23465 (N_23465,N_22067,N_22608);
or U23466 (N_23466,N_22192,N_22015);
or U23467 (N_23467,N_22489,N_22020);
or U23468 (N_23468,N_22729,N_22508);
xnor U23469 (N_23469,N_22347,N_22022);
or U23470 (N_23470,N_22357,N_22323);
or U23471 (N_23471,N_22516,N_22034);
xor U23472 (N_23472,N_22345,N_22788);
nor U23473 (N_23473,N_22354,N_22230);
xor U23474 (N_23474,N_22043,N_22568);
nor U23475 (N_23475,N_22431,N_22014);
nor U23476 (N_23476,N_22180,N_22597);
nand U23477 (N_23477,N_22834,N_22929);
xnor U23478 (N_23478,N_22899,N_22081);
xor U23479 (N_23479,N_22631,N_22862);
xnor U23480 (N_23480,N_22655,N_22806);
or U23481 (N_23481,N_22498,N_22936);
and U23482 (N_23482,N_22123,N_22231);
and U23483 (N_23483,N_22987,N_22805);
nand U23484 (N_23484,N_22549,N_22339);
and U23485 (N_23485,N_22835,N_22830);
nor U23486 (N_23486,N_22966,N_22810);
and U23487 (N_23487,N_22141,N_22924);
nor U23488 (N_23488,N_22218,N_22687);
nor U23489 (N_23489,N_22614,N_22481);
or U23490 (N_23490,N_22761,N_22884);
or U23491 (N_23491,N_22771,N_22207);
nand U23492 (N_23492,N_22820,N_22586);
nand U23493 (N_23493,N_22039,N_22704);
and U23494 (N_23494,N_22063,N_22268);
nand U23495 (N_23495,N_22142,N_22082);
and U23496 (N_23496,N_22075,N_22706);
and U23497 (N_23497,N_22438,N_22305);
nand U23498 (N_23498,N_22547,N_22443);
and U23499 (N_23499,N_22701,N_22895);
xor U23500 (N_23500,N_22514,N_22661);
nand U23501 (N_23501,N_22263,N_22046);
nand U23502 (N_23502,N_22871,N_22316);
and U23503 (N_23503,N_22706,N_22975);
nor U23504 (N_23504,N_22133,N_22634);
nand U23505 (N_23505,N_22293,N_22538);
or U23506 (N_23506,N_22195,N_22936);
or U23507 (N_23507,N_22749,N_22457);
xnor U23508 (N_23508,N_22870,N_22397);
nand U23509 (N_23509,N_22136,N_22856);
xor U23510 (N_23510,N_22080,N_22126);
and U23511 (N_23511,N_22083,N_22018);
xor U23512 (N_23512,N_22344,N_22920);
nand U23513 (N_23513,N_22270,N_22108);
nand U23514 (N_23514,N_22121,N_22216);
and U23515 (N_23515,N_22291,N_22887);
and U23516 (N_23516,N_22502,N_22445);
and U23517 (N_23517,N_22111,N_22658);
nor U23518 (N_23518,N_22652,N_22572);
and U23519 (N_23519,N_22949,N_22525);
nor U23520 (N_23520,N_22632,N_22296);
and U23521 (N_23521,N_22147,N_22934);
xnor U23522 (N_23522,N_22904,N_22934);
or U23523 (N_23523,N_22410,N_22193);
nor U23524 (N_23524,N_22839,N_22430);
and U23525 (N_23525,N_22738,N_22860);
or U23526 (N_23526,N_22168,N_22550);
nand U23527 (N_23527,N_22027,N_22455);
xnor U23528 (N_23528,N_22908,N_22718);
nand U23529 (N_23529,N_22925,N_22027);
nor U23530 (N_23530,N_22198,N_22192);
and U23531 (N_23531,N_22928,N_22499);
and U23532 (N_23532,N_22504,N_22818);
and U23533 (N_23533,N_22633,N_22499);
nand U23534 (N_23534,N_22969,N_22545);
and U23535 (N_23535,N_22901,N_22330);
or U23536 (N_23536,N_22005,N_22034);
and U23537 (N_23537,N_22975,N_22999);
nor U23538 (N_23538,N_22378,N_22195);
nand U23539 (N_23539,N_22886,N_22331);
or U23540 (N_23540,N_22893,N_22514);
xor U23541 (N_23541,N_22085,N_22951);
xnor U23542 (N_23542,N_22916,N_22028);
xor U23543 (N_23543,N_22787,N_22761);
and U23544 (N_23544,N_22864,N_22304);
or U23545 (N_23545,N_22567,N_22111);
or U23546 (N_23546,N_22687,N_22446);
nor U23547 (N_23547,N_22329,N_22166);
and U23548 (N_23548,N_22633,N_22662);
and U23549 (N_23549,N_22438,N_22170);
nand U23550 (N_23550,N_22530,N_22749);
and U23551 (N_23551,N_22246,N_22404);
nand U23552 (N_23552,N_22144,N_22122);
or U23553 (N_23553,N_22188,N_22606);
xnor U23554 (N_23554,N_22211,N_22320);
nor U23555 (N_23555,N_22617,N_22691);
nor U23556 (N_23556,N_22452,N_22041);
and U23557 (N_23557,N_22787,N_22876);
and U23558 (N_23558,N_22877,N_22590);
nor U23559 (N_23559,N_22150,N_22108);
or U23560 (N_23560,N_22007,N_22623);
and U23561 (N_23561,N_22531,N_22016);
and U23562 (N_23562,N_22325,N_22370);
xor U23563 (N_23563,N_22186,N_22223);
or U23564 (N_23564,N_22782,N_22375);
or U23565 (N_23565,N_22689,N_22860);
nand U23566 (N_23566,N_22315,N_22249);
and U23567 (N_23567,N_22570,N_22231);
or U23568 (N_23568,N_22375,N_22382);
or U23569 (N_23569,N_22214,N_22028);
or U23570 (N_23570,N_22356,N_22093);
and U23571 (N_23571,N_22474,N_22534);
nor U23572 (N_23572,N_22117,N_22002);
and U23573 (N_23573,N_22824,N_22954);
xor U23574 (N_23574,N_22391,N_22038);
and U23575 (N_23575,N_22230,N_22176);
or U23576 (N_23576,N_22652,N_22317);
nand U23577 (N_23577,N_22726,N_22183);
or U23578 (N_23578,N_22607,N_22765);
or U23579 (N_23579,N_22864,N_22611);
or U23580 (N_23580,N_22090,N_22772);
or U23581 (N_23581,N_22816,N_22957);
nand U23582 (N_23582,N_22375,N_22937);
nor U23583 (N_23583,N_22189,N_22037);
nand U23584 (N_23584,N_22408,N_22309);
nor U23585 (N_23585,N_22571,N_22285);
and U23586 (N_23586,N_22914,N_22510);
or U23587 (N_23587,N_22356,N_22015);
and U23588 (N_23588,N_22363,N_22335);
nor U23589 (N_23589,N_22557,N_22675);
xnor U23590 (N_23590,N_22862,N_22876);
nor U23591 (N_23591,N_22037,N_22749);
nor U23592 (N_23592,N_22830,N_22754);
nand U23593 (N_23593,N_22507,N_22686);
nand U23594 (N_23594,N_22536,N_22593);
or U23595 (N_23595,N_22936,N_22636);
and U23596 (N_23596,N_22612,N_22039);
or U23597 (N_23597,N_22748,N_22631);
or U23598 (N_23598,N_22660,N_22793);
and U23599 (N_23599,N_22545,N_22835);
nand U23600 (N_23600,N_22102,N_22770);
nor U23601 (N_23601,N_22619,N_22483);
or U23602 (N_23602,N_22196,N_22590);
xnor U23603 (N_23603,N_22132,N_22038);
xnor U23604 (N_23604,N_22376,N_22144);
and U23605 (N_23605,N_22124,N_22748);
nand U23606 (N_23606,N_22398,N_22382);
nor U23607 (N_23607,N_22310,N_22471);
and U23608 (N_23608,N_22759,N_22922);
or U23609 (N_23609,N_22966,N_22245);
nand U23610 (N_23610,N_22256,N_22414);
nor U23611 (N_23611,N_22583,N_22030);
nor U23612 (N_23612,N_22172,N_22081);
nand U23613 (N_23613,N_22048,N_22486);
nand U23614 (N_23614,N_22703,N_22141);
and U23615 (N_23615,N_22531,N_22292);
nor U23616 (N_23616,N_22385,N_22591);
and U23617 (N_23617,N_22973,N_22157);
or U23618 (N_23618,N_22914,N_22152);
nand U23619 (N_23619,N_22328,N_22990);
nand U23620 (N_23620,N_22411,N_22870);
xor U23621 (N_23621,N_22121,N_22946);
nor U23622 (N_23622,N_22180,N_22799);
xor U23623 (N_23623,N_22013,N_22777);
nor U23624 (N_23624,N_22877,N_22920);
or U23625 (N_23625,N_22443,N_22245);
xnor U23626 (N_23626,N_22041,N_22179);
and U23627 (N_23627,N_22809,N_22194);
or U23628 (N_23628,N_22469,N_22707);
and U23629 (N_23629,N_22755,N_22923);
and U23630 (N_23630,N_22847,N_22002);
nand U23631 (N_23631,N_22319,N_22974);
nor U23632 (N_23632,N_22445,N_22243);
nor U23633 (N_23633,N_22084,N_22043);
xor U23634 (N_23634,N_22590,N_22585);
and U23635 (N_23635,N_22732,N_22118);
xor U23636 (N_23636,N_22404,N_22852);
nand U23637 (N_23637,N_22135,N_22313);
or U23638 (N_23638,N_22631,N_22440);
xor U23639 (N_23639,N_22039,N_22047);
or U23640 (N_23640,N_22897,N_22220);
nor U23641 (N_23641,N_22543,N_22776);
or U23642 (N_23642,N_22346,N_22077);
or U23643 (N_23643,N_22361,N_22418);
nor U23644 (N_23644,N_22523,N_22150);
xor U23645 (N_23645,N_22856,N_22603);
or U23646 (N_23646,N_22380,N_22787);
nor U23647 (N_23647,N_22608,N_22986);
nand U23648 (N_23648,N_22217,N_22973);
nor U23649 (N_23649,N_22884,N_22824);
and U23650 (N_23650,N_22225,N_22758);
nand U23651 (N_23651,N_22219,N_22068);
nand U23652 (N_23652,N_22098,N_22255);
nor U23653 (N_23653,N_22546,N_22731);
nor U23654 (N_23654,N_22457,N_22401);
nand U23655 (N_23655,N_22435,N_22615);
and U23656 (N_23656,N_22037,N_22718);
xnor U23657 (N_23657,N_22601,N_22517);
nand U23658 (N_23658,N_22991,N_22457);
nand U23659 (N_23659,N_22239,N_22329);
nand U23660 (N_23660,N_22641,N_22801);
nor U23661 (N_23661,N_22419,N_22313);
xnor U23662 (N_23662,N_22828,N_22572);
xor U23663 (N_23663,N_22588,N_22106);
or U23664 (N_23664,N_22731,N_22137);
or U23665 (N_23665,N_22976,N_22326);
nand U23666 (N_23666,N_22889,N_22593);
nor U23667 (N_23667,N_22171,N_22647);
nand U23668 (N_23668,N_22529,N_22829);
or U23669 (N_23669,N_22963,N_22709);
nor U23670 (N_23670,N_22672,N_22950);
nand U23671 (N_23671,N_22992,N_22420);
nand U23672 (N_23672,N_22735,N_22573);
or U23673 (N_23673,N_22210,N_22992);
nand U23674 (N_23674,N_22142,N_22525);
nor U23675 (N_23675,N_22669,N_22959);
nor U23676 (N_23676,N_22009,N_22583);
nand U23677 (N_23677,N_22867,N_22337);
xor U23678 (N_23678,N_22319,N_22839);
xnor U23679 (N_23679,N_22256,N_22163);
nand U23680 (N_23680,N_22787,N_22644);
or U23681 (N_23681,N_22048,N_22598);
or U23682 (N_23682,N_22547,N_22403);
or U23683 (N_23683,N_22442,N_22907);
xor U23684 (N_23684,N_22056,N_22237);
nand U23685 (N_23685,N_22738,N_22480);
and U23686 (N_23686,N_22420,N_22226);
nor U23687 (N_23687,N_22257,N_22436);
and U23688 (N_23688,N_22362,N_22569);
xor U23689 (N_23689,N_22138,N_22931);
nor U23690 (N_23690,N_22081,N_22231);
and U23691 (N_23691,N_22639,N_22519);
or U23692 (N_23692,N_22317,N_22489);
nand U23693 (N_23693,N_22603,N_22635);
xnor U23694 (N_23694,N_22227,N_22382);
xor U23695 (N_23695,N_22606,N_22105);
xnor U23696 (N_23696,N_22456,N_22962);
nand U23697 (N_23697,N_22200,N_22881);
or U23698 (N_23698,N_22976,N_22772);
xor U23699 (N_23699,N_22954,N_22664);
nand U23700 (N_23700,N_22791,N_22625);
nand U23701 (N_23701,N_22027,N_22704);
and U23702 (N_23702,N_22891,N_22556);
nor U23703 (N_23703,N_22228,N_22392);
and U23704 (N_23704,N_22635,N_22165);
nor U23705 (N_23705,N_22557,N_22396);
nor U23706 (N_23706,N_22782,N_22554);
nor U23707 (N_23707,N_22677,N_22654);
nor U23708 (N_23708,N_22797,N_22013);
xnor U23709 (N_23709,N_22274,N_22589);
or U23710 (N_23710,N_22037,N_22026);
nand U23711 (N_23711,N_22935,N_22936);
xor U23712 (N_23712,N_22804,N_22550);
xor U23713 (N_23713,N_22201,N_22874);
and U23714 (N_23714,N_22670,N_22553);
and U23715 (N_23715,N_22425,N_22404);
nor U23716 (N_23716,N_22852,N_22525);
xor U23717 (N_23717,N_22602,N_22628);
or U23718 (N_23718,N_22140,N_22847);
and U23719 (N_23719,N_22195,N_22851);
nand U23720 (N_23720,N_22905,N_22096);
nor U23721 (N_23721,N_22077,N_22990);
nand U23722 (N_23722,N_22557,N_22540);
nand U23723 (N_23723,N_22955,N_22616);
and U23724 (N_23724,N_22429,N_22605);
or U23725 (N_23725,N_22365,N_22546);
and U23726 (N_23726,N_22235,N_22650);
and U23727 (N_23727,N_22805,N_22495);
nand U23728 (N_23728,N_22067,N_22360);
nor U23729 (N_23729,N_22290,N_22082);
and U23730 (N_23730,N_22159,N_22466);
or U23731 (N_23731,N_22479,N_22095);
and U23732 (N_23732,N_22075,N_22377);
xnor U23733 (N_23733,N_22182,N_22364);
xnor U23734 (N_23734,N_22458,N_22296);
xnor U23735 (N_23735,N_22503,N_22647);
or U23736 (N_23736,N_22281,N_22669);
nor U23737 (N_23737,N_22850,N_22780);
xor U23738 (N_23738,N_22706,N_22280);
and U23739 (N_23739,N_22573,N_22217);
nand U23740 (N_23740,N_22757,N_22217);
xnor U23741 (N_23741,N_22668,N_22108);
and U23742 (N_23742,N_22117,N_22295);
nor U23743 (N_23743,N_22692,N_22375);
nor U23744 (N_23744,N_22813,N_22034);
nand U23745 (N_23745,N_22091,N_22482);
xor U23746 (N_23746,N_22955,N_22239);
nand U23747 (N_23747,N_22188,N_22171);
or U23748 (N_23748,N_22065,N_22419);
nor U23749 (N_23749,N_22136,N_22562);
or U23750 (N_23750,N_22332,N_22074);
or U23751 (N_23751,N_22534,N_22856);
xor U23752 (N_23752,N_22928,N_22159);
and U23753 (N_23753,N_22403,N_22134);
nor U23754 (N_23754,N_22589,N_22915);
nand U23755 (N_23755,N_22647,N_22328);
and U23756 (N_23756,N_22253,N_22091);
or U23757 (N_23757,N_22337,N_22151);
xnor U23758 (N_23758,N_22050,N_22292);
xor U23759 (N_23759,N_22075,N_22931);
and U23760 (N_23760,N_22850,N_22342);
xor U23761 (N_23761,N_22271,N_22721);
and U23762 (N_23762,N_22757,N_22103);
xor U23763 (N_23763,N_22823,N_22114);
nor U23764 (N_23764,N_22251,N_22987);
or U23765 (N_23765,N_22672,N_22942);
or U23766 (N_23766,N_22484,N_22707);
xor U23767 (N_23767,N_22631,N_22778);
and U23768 (N_23768,N_22502,N_22138);
nand U23769 (N_23769,N_22801,N_22896);
nor U23770 (N_23770,N_22132,N_22819);
xnor U23771 (N_23771,N_22342,N_22160);
nor U23772 (N_23772,N_22091,N_22989);
xnor U23773 (N_23773,N_22860,N_22492);
xor U23774 (N_23774,N_22631,N_22211);
or U23775 (N_23775,N_22772,N_22021);
xor U23776 (N_23776,N_22741,N_22802);
or U23777 (N_23777,N_22687,N_22125);
or U23778 (N_23778,N_22582,N_22738);
and U23779 (N_23779,N_22569,N_22841);
and U23780 (N_23780,N_22133,N_22078);
nor U23781 (N_23781,N_22718,N_22416);
nand U23782 (N_23782,N_22105,N_22980);
and U23783 (N_23783,N_22895,N_22355);
xnor U23784 (N_23784,N_22516,N_22907);
and U23785 (N_23785,N_22468,N_22954);
xor U23786 (N_23786,N_22960,N_22130);
and U23787 (N_23787,N_22341,N_22937);
nand U23788 (N_23788,N_22390,N_22934);
nor U23789 (N_23789,N_22700,N_22995);
nand U23790 (N_23790,N_22505,N_22108);
nand U23791 (N_23791,N_22024,N_22747);
nand U23792 (N_23792,N_22624,N_22019);
or U23793 (N_23793,N_22584,N_22930);
or U23794 (N_23794,N_22462,N_22909);
nand U23795 (N_23795,N_22078,N_22498);
nand U23796 (N_23796,N_22604,N_22857);
xor U23797 (N_23797,N_22424,N_22594);
nor U23798 (N_23798,N_22322,N_22931);
nand U23799 (N_23799,N_22054,N_22438);
nand U23800 (N_23800,N_22088,N_22722);
nand U23801 (N_23801,N_22240,N_22495);
or U23802 (N_23802,N_22033,N_22270);
nand U23803 (N_23803,N_22833,N_22601);
or U23804 (N_23804,N_22612,N_22190);
and U23805 (N_23805,N_22904,N_22785);
xor U23806 (N_23806,N_22947,N_22003);
and U23807 (N_23807,N_22052,N_22437);
and U23808 (N_23808,N_22162,N_22654);
nor U23809 (N_23809,N_22149,N_22089);
xnor U23810 (N_23810,N_22480,N_22213);
nor U23811 (N_23811,N_22231,N_22374);
nand U23812 (N_23812,N_22150,N_22310);
xor U23813 (N_23813,N_22688,N_22618);
xor U23814 (N_23814,N_22752,N_22711);
nor U23815 (N_23815,N_22729,N_22245);
nand U23816 (N_23816,N_22163,N_22694);
and U23817 (N_23817,N_22628,N_22089);
nand U23818 (N_23818,N_22624,N_22601);
nand U23819 (N_23819,N_22283,N_22931);
or U23820 (N_23820,N_22944,N_22908);
and U23821 (N_23821,N_22069,N_22105);
or U23822 (N_23822,N_22355,N_22255);
and U23823 (N_23823,N_22533,N_22513);
or U23824 (N_23824,N_22419,N_22969);
and U23825 (N_23825,N_22180,N_22694);
nand U23826 (N_23826,N_22877,N_22433);
and U23827 (N_23827,N_22494,N_22562);
nor U23828 (N_23828,N_22163,N_22899);
or U23829 (N_23829,N_22630,N_22976);
nand U23830 (N_23830,N_22018,N_22098);
xnor U23831 (N_23831,N_22507,N_22203);
nor U23832 (N_23832,N_22337,N_22368);
nor U23833 (N_23833,N_22915,N_22356);
or U23834 (N_23834,N_22760,N_22866);
xnor U23835 (N_23835,N_22602,N_22614);
nor U23836 (N_23836,N_22882,N_22782);
or U23837 (N_23837,N_22078,N_22464);
or U23838 (N_23838,N_22815,N_22602);
nand U23839 (N_23839,N_22226,N_22365);
and U23840 (N_23840,N_22352,N_22622);
or U23841 (N_23841,N_22944,N_22846);
and U23842 (N_23842,N_22395,N_22064);
nor U23843 (N_23843,N_22563,N_22611);
nand U23844 (N_23844,N_22764,N_22689);
nand U23845 (N_23845,N_22319,N_22006);
and U23846 (N_23846,N_22454,N_22509);
or U23847 (N_23847,N_22287,N_22596);
nand U23848 (N_23848,N_22454,N_22304);
nor U23849 (N_23849,N_22310,N_22485);
nand U23850 (N_23850,N_22984,N_22063);
and U23851 (N_23851,N_22243,N_22536);
xnor U23852 (N_23852,N_22515,N_22488);
xnor U23853 (N_23853,N_22948,N_22501);
xor U23854 (N_23854,N_22038,N_22905);
and U23855 (N_23855,N_22469,N_22876);
and U23856 (N_23856,N_22822,N_22810);
or U23857 (N_23857,N_22366,N_22712);
nor U23858 (N_23858,N_22388,N_22741);
or U23859 (N_23859,N_22477,N_22721);
and U23860 (N_23860,N_22358,N_22724);
and U23861 (N_23861,N_22341,N_22171);
nor U23862 (N_23862,N_22666,N_22588);
nor U23863 (N_23863,N_22806,N_22555);
or U23864 (N_23864,N_22266,N_22852);
xor U23865 (N_23865,N_22780,N_22413);
or U23866 (N_23866,N_22439,N_22845);
xnor U23867 (N_23867,N_22597,N_22369);
xnor U23868 (N_23868,N_22338,N_22129);
xor U23869 (N_23869,N_22068,N_22893);
and U23870 (N_23870,N_22321,N_22633);
xnor U23871 (N_23871,N_22453,N_22363);
xor U23872 (N_23872,N_22074,N_22091);
and U23873 (N_23873,N_22086,N_22782);
nor U23874 (N_23874,N_22809,N_22645);
nand U23875 (N_23875,N_22119,N_22448);
nand U23876 (N_23876,N_22622,N_22599);
nand U23877 (N_23877,N_22741,N_22863);
nand U23878 (N_23878,N_22316,N_22099);
nand U23879 (N_23879,N_22487,N_22315);
nand U23880 (N_23880,N_22514,N_22588);
and U23881 (N_23881,N_22333,N_22785);
xor U23882 (N_23882,N_22168,N_22099);
or U23883 (N_23883,N_22466,N_22487);
xor U23884 (N_23884,N_22070,N_22305);
xor U23885 (N_23885,N_22192,N_22597);
nand U23886 (N_23886,N_22572,N_22862);
nor U23887 (N_23887,N_22680,N_22983);
nand U23888 (N_23888,N_22905,N_22036);
xor U23889 (N_23889,N_22908,N_22688);
or U23890 (N_23890,N_22389,N_22771);
nand U23891 (N_23891,N_22771,N_22363);
and U23892 (N_23892,N_22780,N_22758);
nor U23893 (N_23893,N_22662,N_22123);
or U23894 (N_23894,N_22833,N_22175);
or U23895 (N_23895,N_22004,N_22260);
or U23896 (N_23896,N_22832,N_22582);
nor U23897 (N_23897,N_22157,N_22173);
or U23898 (N_23898,N_22514,N_22177);
nor U23899 (N_23899,N_22942,N_22136);
or U23900 (N_23900,N_22769,N_22058);
nand U23901 (N_23901,N_22860,N_22786);
or U23902 (N_23902,N_22778,N_22677);
or U23903 (N_23903,N_22101,N_22944);
and U23904 (N_23904,N_22370,N_22523);
nor U23905 (N_23905,N_22102,N_22522);
xor U23906 (N_23906,N_22744,N_22242);
xnor U23907 (N_23907,N_22880,N_22906);
or U23908 (N_23908,N_22348,N_22168);
nor U23909 (N_23909,N_22338,N_22085);
nand U23910 (N_23910,N_22196,N_22437);
or U23911 (N_23911,N_22755,N_22160);
and U23912 (N_23912,N_22231,N_22149);
or U23913 (N_23913,N_22723,N_22068);
nand U23914 (N_23914,N_22676,N_22177);
and U23915 (N_23915,N_22016,N_22305);
or U23916 (N_23916,N_22957,N_22633);
xnor U23917 (N_23917,N_22792,N_22565);
nor U23918 (N_23918,N_22719,N_22520);
or U23919 (N_23919,N_22644,N_22708);
nand U23920 (N_23920,N_22164,N_22096);
nand U23921 (N_23921,N_22501,N_22919);
or U23922 (N_23922,N_22489,N_22949);
and U23923 (N_23923,N_22350,N_22077);
or U23924 (N_23924,N_22801,N_22436);
and U23925 (N_23925,N_22609,N_22038);
nand U23926 (N_23926,N_22256,N_22036);
and U23927 (N_23927,N_22109,N_22891);
or U23928 (N_23928,N_22605,N_22124);
and U23929 (N_23929,N_22892,N_22218);
nand U23930 (N_23930,N_22972,N_22543);
nand U23931 (N_23931,N_22381,N_22554);
xor U23932 (N_23932,N_22093,N_22948);
nor U23933 (N_23933,N_22924,N_22227);
nor U23934 (N_23934,N_22046,N_22659);
or U23935 (N_23935,N_22114,N_22095);
and U23936 (N_23936,N_22511,N_22203);
or U23937 (N_23937,N_22161,N_22831);
nand U23938 (N_23938,N_22052,N_22929);
or U23939 (N_23939,N_22047,N_22854);
nor U23940 (N_23940,N_22491,N_22402);
nor U23941 (N_23941,N_22950,N_22411);
nand U23942 (N_23942,N_22388,N_22495);
nor U23943 (N_23943,N_22232,N_22922);
nor U23944 (N_23944,N_22274,N_22942);
and U23945 (N_23945,N_22859,N_22276);
xnor U23946 (N_23946,N_22817,N_22006);
or U23947 (N_23947,N_22294,N_22045);
or U23948 (N_23948,N_22155,N_22163);
nor U23949 (N_23949,N_22142,N_22465);
nand U23950 (N_23950,N_22623,N_22176);
and U23951 (N_23951,N_22180,N_22552);
xnor U23952 (N_23952,N_22314,N_22982);
nor U23953 (N_23953,N_22524,N_22808);
nor U23954 (N_23954,N_22329,N_22846);
nand U23955 (N_23955,N_22252,N_22563);
nor U23956 (N_23956,N_22336,N_22021);
and U23957 (N_23957,N_22921,N_22048);
nand U23958 (N_23958,N_22922,N_22227);
and U23959 (N_23959,N_22403,N_22926);
nand U23960 (N_23960,N_22467,N_22815);
or U23961 (N_23961,N_22896,N_22503);
nand U23962 (N_23962,N_22940,N_22888);
nand U23963 (N_23963,N_22402,N_22768);
xnor U23964 (N_23964,N_22859,N_22901);
nor U23965 (N_23965,N_22183,N_22285);
nand U23966 (N_23966,N_22783,N_22954);
nor U23967 (N_23967,N_22880,N_22718);
nor U23968 (N_23968,N_22238,N_22472);
nand U23969 (N_23969,N_22837,N_22308);
and U23970 (N_23970,N_22497,N_22098);
or U23971 (N_23971,N_22966,N_22273);
nand U23972 (N_23972,N_22814,N_22349);
and U23973 (N_23973,N_22233,N_22652);
and U23974 (N_23974,N_22401,N_22358);
nand U23975 (N_23975,N_22806,N_22291);
xnor U23976 (N_23976,N_22992,N_22199);
or U23977 (N_23977,N_22951,N_22402);
nand U23978 (N_23978,N_22319,N_22044);
nand U23979 (N_23979,N_22022,N_22956);
xor U23980 (N_23980,N_22870,N_22818);
or U23981 (N_23981,N_22033,N_22636);
nor U23982 (N_23982,N_22714,N_22648);
nand U23983 (N_23983,N_22391,N_22275);
nor U23984 (N_23984,N_22042,N_22340);
xnor U23985 (N_23985,N_22779,N_22956);
nand U23986 (N_23986,N_22058,N_22491);
and U23987 (N_23987,N_22788,N_22593);
nor U23988 (N_23988,N_22249,N_22969);
nor U23989 (N_23989,N_22337,N_22522);
nor U23990 (N_23990,N_22800,N_22442);
nor U23991 (N_23991,N_22255,N_22527);
nor U23992 (N_23992,N_22018,N_22705);
and U23993 (N_23993,N_22738,N_22844);
nand U23994 (N_23994,N_22062,N_22528);
nand U23995 (N_23995,N_22986,N_22528);
xor U23996 (N_23996,N_22918,N_22882);
nand U23997 (N_23997,N_22832,N_22950);
xnor U23998 (N_23998,N_22953,N_22449);
nor U23999 (N_23999,N_22446,N_22004);
xnor U24000 (N_24000,N_23157,N_23313);
or U24001 (N_24001,N_23019,N_23223);
nand U24002 (N_24002,N_23394,N_23284);
nor U24003 (N_24003,N_23675,N_23132);
and U24004 (N_24004,N_23321,N_23882);
nor U24005 (N_24005,N_23089,N_23240);
and U24006 (N_24006,N_23806,N_23176);
and U24007 (N_24007,N_23362,N_23414);
xor U24008 (N_24008,N_23274,N_23514);
or U24009 (N_24009,N_23179,N_23737);
or U24010 (N_24010,N_23359,N_23231);
or U24011 (N_24011,N_23234,N_23689);
or U24012 (N_24012,N_23183,N_23189);
xnor U24013 (N_24013,N_23392,N_23738);
or U24014 (N_24014,N_23066,N_23372);
or U24015 (N_24015,N_23273,N_23379);
nand U24016 (N_24016,N_23615,N_23923);
xnor U24017 (N_24017,N_23518,N_23925);
xor U24018 (N_24018,N_23540,N_23431);
xnor U24019 (N_24019,N_23896,N_23852);
nand U24020 (N_24020,N_23343,N_23100);
nor U24021 (N_24021,N_23690,N_23058);
and U24022 (N_24022,N_23940,N_23279);
or U24023 (N_24023,N_23190,N_23053);
nor U24024 (N_24024,N_23855,N_23853);
nor U24025 (N_24025,N_23626,N_23479);
nor U24026 (N_24026,N_23427,N_23520);
or U24027 (N_24027,N_23135,N_23011);
nand U24028 (N_24028,N_23287,N_23426);
or U24029 (N_24029,N_23204,N_23947);
nand U24030 (N_24030,N_23466,N_23785);
or U24031 (N_24031,N_23085,N_23091);
nor U24032 (N_24032,N_23782,N_23904);
nor U24033 (N_24033,N_23986,N_23922);
nand U24034 (N_24034,N_23030,N_23528);
nand U24035 (N_24035,N_23124,N_23798);
nor U24036 (N_24036,N_23692,N_23031);
nor U24037 (N_24037,N_23046,N_23230);
or U24038 (N_24038,N_23902,N_23489);
and U24039 (N_24039,N_23824,N_23086);
xnor U24040 (N_24040,N_23028,N_23914);
and U24041 (N_24041,N_23792,N_23472);
nand U24042 (N_24042,N_23254,N_23498);
nand U24043 (N_24043,N_23764,N_23718);
or U24044 (N_24044,N_23319,N_23935);
and U24045 (N_24045,N_23396,N_23171);
nand U24046 (N_24046,N_23126,N_23530);
xor U24047 (N_24047,N_23945,N_23791);
nor U24048 (N_24048,N_23004,N_23339);
and U24049 (N_24049,N_23468,N_23859);
nand U24050 (N_24050,N_23278,N_23251);
nand U24051 (N_24051,N_23756,N_23716);
xnor U24052 (N_24052,N_23741,N_23860);
xnor U24053 (N_24053,N_23570,N_23233);
or U24054 (N_24054,N_23780,N_23430);
nor U24055 (N_24055,N_23971,N_23163);
and U24056 (N_24056,N_23629,N_23476);
nand U24057 (N_24057,N_23025,N_23981);
or U24058 (N_24058,N_23774,N_23326);
nand U24059 (N_24059,N_23589,N_23699);
xnor U24060 (N_24060,N_23497,N_23338);
or U24061 (N_24061,N_23933,N_23453);
or U24062 (N_24062,N_23803,N_23207);
or U24063 (N_24063,N_23436,N_23827);
nor U24064 (N_24064,N_23460,N_23728);
nor U24065 (N_24065,N_23016,N_23351);
xor U24066 (N_24066,N_23143,N_23063);
nand U24067 (N_24067,N_23041,N_23921);
or U24068 (N_24068,N_23618,N_23154);
and U24069 (N_24069,N_23366,N_23247);
nor U24070 (N_24070,N_23382,N_23762);
xnor U24071 (N_24071,N_23691,N_23934);
and U24072 (N_24072,N_23329,N_23671);
xnor U24073 (N_24073,N_23161,N_23742);
nand U24074 (N_24074,N_23751,N_23409);
xor U24075 (N_24075,N_23378,N_23515);
nor U24076 (N_24076,N_23021,N_23113);
nor U24077 (N_24077,N_23197,N_23502);
nor U24078 (N_24078,N_23897,N_23425);
xnor U24079 (N_24079,N_23908,N_23758);
xnor U24080 (N_24080,N_23001,N_23121);
xnor U24081 (N_24081,N_23057,N_23309);
or U24082 (N_24082,N_23545,N_23707);
nand U24083 (N_24083,N_23282,N_23301);
or U24084 (N_24084,N_23964,N_23395);
nand U24085 (N_24085,N_23672,N_23535);
and U24086 (N_24086,N_23353,N_23187);
xor U24087 (N_24087,N_23790,N_23663);
and U24088 (N_24088,N_23628,N_23735);
or U24089 (N_24089,N_23843,N_23277);
nor U24090 (N_24090,N_23719,N_23302);
nor U24091 (N_24091,N_23448,N_23506);
xnor U24092 (N_24092,N_23052,N_23049);
nor U24093 (N_24093,N_23311,N_23314);
nand U24094 (N_24094,N_23641,N_23295);
and U24095 (N_24095,N_23386,N_23661);
or U24096 (N_24096,N_23345,N_23428);
nand U24097 (N_24097,N_23607,N_23634);
nor U24098 (N_24098,N_23038,N_23836);
or U24099 (N_24099,N_23920,N_23370);
nor U24100 (N_24100,N_23733,N_23048);
nand U24101 (N_24101,N_23300,N_23821);
nor U24102 (N_24102,N_23265,N_23554);
xnor U24103 (N_24103,N_23494,N_23673);
xor U24104 (N_24104,N_23638,N_23283);
xor U24105 (N_24105,N_23648,N_23595);
nor U24106 (N_24106,N_23109,N_23260);
or U24107 (N_24107,N_23772,N_23055);
or U24108 (N_24108,N_23172,N_23071);
and U24109 (N_24109,N_23341,N_23419);
and U24110 (N_24110,N_23894,N_23499);
or U24111 (N_24111,N_23434,N_23481);
nand U24112 (N_24112,N_23397,N_23169);
or U24113 (N_24113,N_23891,N_23591);
nor U24114 (N_24114,N_23929,N_23544);
xnor U24115 (N_24115,N_23484,N_23232);
and U24116 (N_24116,N_23994,N_23146);
nand U24117 (N_24117,N_23318,N_23660);
nand U24118 (N_24118,N_23070,N_23624);
and U24119 (N_24119,N_23639,N_23166);
nor U24120 (N_24120,N_23931,N_23103);
and U24121 (N_24121,N_23965,N_23950);
xnor U24122 (N_24122,N_23152,N_23145);
and U24123 (N_24123,N_23708,N_23608);
nand U24124 (N_24124,N_23308,N_23093);
nor U24125 (N_24125,N_23483,N_23203);
nor U24126 (N_24126,N_23839,N_23846);
or U24127 (N_24127,N_23125,N_23208);
nor U24128 (N_24128,N_23695,N_23294);
and U24129 (N_24129,N_23275,N_23034);
xor U24130 (N_24130,N_23850,N_23400);
nor U24131 (N_24131,N_23709,N_23477);
nand U24132 (N_24132,N_23867,N_23014);
nand U24133 (N_24133,N_23838,N_23482);
xor U24134 (N_24134,N_23401,N_23606);
nand U24135 (N_24135,N_23130,N_23969);
nor U24136 (N_24136,N_23511,N_23635);
xor U24137 (N_24137,N_23598,N_23706);
nand U24138 (N_24138,N_23927,N_23067);
and U24139 (N_24139,N_23559,N_23155);
and U24140 (N_24140,N_23555,N_23422);
or U24141 (N_24141,N_23061,N_23280);
xor U24142 (N_24142,N_23703,N_23438);
xor U24143 (N_24143,N_23315,N_23563);
or U24144 (N_24144,N_23101,N_23445);
or U24145 (N_24145,N_23771,N_23237);
and U24146 (N_24146,N_23220,N_23322);
and U24147 (N_24147,N_23465,N_23227);
nand U24148 (N_24148,N_23375,N_23115);
nor U24149 (N_24149,N_23120,N_23997);
nand U24150 (N_24150,N_23787,N_23610);
xor U24151 (N_24151,N_23022,N_23813);
nand U24152 (N_24152,N_23727,N_23676);
or U24153 (N_24153,N_23668,N_23987);
or U24154 (N_24154,N_23566,N_23948);
nor U24155 (N_24155,N_23887,N_23127);
xor U24156 (N_24156,N_23088,N_23087);
or U24157 (N_24157,N_23469,N_23677);
or U24158 (N_24158,N_23202,N_23435);
xor U24159 (N_24159,N_23236,N_23377);
and U24160 (N_24160,N_23212,N_23732);
xor U24161 (N_24161,N_23096,N_23794);
and U24162 (N_24162,N_23259,N_23939);
nor U24163 (N_24163,N_23678,N_23715);
or U24164 (N_24164,N_23873,N_23833);
and U24165 (N_24165,N_23527,N_23193);
xnor U24166 (N_24166,N_23334,N_23439);
and U24167 (N_24167,N_23398,N_23487);
and U24168 (N_24168,N_23105,N_23082);
nand U24169 (N_24169,N_23619,N_23862);
nor U24170 (N_24170,N_23131,N_23252);
and U24171 (N_24171,N_23578,N_23214);
xnor U24172 (N_24172,N_23122,N_23636);
or U24173 (N_24173,N_23463,N_23700);
xnor U24174 (N_24174,N_23449,N_23336);
nand U24175 (N_24175,N_23029,N_23106);
xnor U24176 (N_24176,N_23167,N_23516);
or U24177 (N_24177,N_23271,N_23561);
xnor U24178 (N_24178,N_23184,N_23342);
or U24179 (N_24179,N_23285,N_23770);
or U24180 (N_24180,N_23918,N_23363);
nor U24181 (N_24181,N_23305,N_23385);
xor U24182 (N_24182,N_23188,N_23826);
xnor U24183 (N_24183,N_23865,N_23954);
and U24184 (N_24184,N_23898,N_23474);
nor U24185 (N_24185,N_23462,N_23364);
nand U24186 (N_24186,N_23156,N_23452);
and U24187 (N_24187,N_23773,N_23538);
nand U24188 (N_24188,N_23604,N_23108);
nand U24189 (N_24189,N_23590,N_23075);
nand U24190 (N_24190,N_23289,N_23178);
nor U24191 (N_24191,N_23281,N_23213);
nand U24192 (N_24192,N_23560,N_23654);
nand U24193 (N_24193,N_23553,N_23745);
nand U24194 (N_24194,N_23493,N_23455);
and U24195 (N_24195,N_23817,N_23942);
nor U24196 (N_24196,N_23246,N_23084);
and U24197 (N_24197,N_23107,N_23829);
and U24198 (N_24198,N_23150,N_23786);
and U24199 (N_24199,N_23953,N_23993);
xnor U24200 (N_24200,N_23748,N_23759);
and U24201 (N_24201,N_23097,N_23702);
xor U24202 (N_24202,N_23244,N_23437);
and U24203 (N_24203,N_23858,N_23381);
nor U24204 (N_24204,N_23991,N_23704);
and U24205 (N_24205,N_23267,N_23946);
nor U24206 (N_24206,N_23222,N_23899);
or U24207 (N_24207,N_23424,N_23524);
xnor U24208 (N_24208,N_23870,N_23988);
nand U24209 (N_24209,N_23814,N_23693);
nand U24210 (N_24210,N_23446,N_23117);
xor U24211 (N_24211,N_23170,N_23492);
nor U24212 (N_24212,N_23299,N_23094);
nor U24213 (N_24213,N_23531,N_23831);
xnor U24214 (N_24214,N_23550,N_23651);
xnor U24215 (N_24215,N_23949,N_23136);
xnor U24216 (N_24216,N_23682,N_23881);
xor U24217 (N_24217,N_23627,N_23005);
xnor U24218 (N_24218,N_23142,N_23241);
nor U24219 (N_24219,N_23664,N_23513);
or U24220 (N_24220,N_23757,N_23797);
or U24221 (N_24221,N_23886,N_23072);
nand U24222 (N_24222,N_23637,N_23263);
or U24223 (N_24223,N_23253,N_23358);
nand U24224 (N_24224,N_23959,N_23781);
nand U24225 (N_24225,N_23532,N_23517);
xnor U24226 (N_24226,N_23478,N_23470);
nor U24227 (N_24227,N_23062,N_23543);
nor U24228 (N_24228,N_23646,N_23711);
nor U24229 (N_24229,N_23984,N_23841);
xnor U24230 (N_24230,N_23665,N_23760);
xnor U24231 (N_24231,N_23847,N_23480);
or U24232 (N_24232,N_23504,N_23198);
xor U24233 (N_24233,N_23743,N_23501);
nand U24234 (N_24234,N_23879,N_23625);
nor U24235 (N_24235,N_23851,N_23734);
nand U24236 (N_24236,N_23195,N_23412);
nor U24237 (N_24237,N_23020,N_23576);
and U24238 (N_24238,N_23266,N_23602);
nor U24239 (N_24239,N_23450,N_23832);
xnor U24240 (N_24240,N_23509,N_23201);
nor U24241 (N_24241,N_23164,N_23903);
nor U24242 (N_24242,N_23588,N_23215);
or U24243 (N_24243,N_23402,N_23390);
or U24244 (N_24244,N_23938,N_23652);
xor U24245 (N_24245,N_23649,N_23168);
nand U24246 (N_24246,N_23441,N_23573);
nand U24247 (N_24247,N_23816,N_23032);
or U24248 (N_24248,N_23036,N_23647);
or U24249 (N_24249,N_23650,N_23739);
nand U24250 (N_24250,N_23730,N_23679);
and U24251 (N_24251,N_23613,N_23906);
nor U24252 (N_24252,N_23023,N_23842);
xnor U24253 (N_24253,N_23328,N_23503);
or U24254 (N_24254,N_23864,N_23801);
nand U24255 (N_24255,N_23344,N_23944);
nor U24256 (N_24256,N_23490,N_23645);
or U24257 (N_24257,N_23261,N_23211);
nand U24258 (N_24258,N_23901,N_23874);
or U24259 (N_24259,N_23128,N_23407);
xor U24260 (N_24260,N_23955,N_23970);
and U24261 (N_24261,N_23026,N_23017);
nand U24262 (N_24262,N_23777,N_23916);
nor U24263 (N_24263,N_23205,N_23539);
or U24264 (N_24264,N_23888,N_23221);
or U24265 (N_24265,N_23697,N_23835);
nor U24266 (N_24266,N_23753,N_23985);
nand U24267 (N_24267,N_23060,N_23040);
xor U24268 (N_24268,N_23614,N_23064);
and U24269 (N_24269,N_23325,N_23235);
nor U24270 (N_24270,N_23868,N_23698);
nor U24271 (N_24271,N_23505,N_23225);
or U24272 (N_24272,N_23622,N_23391);
xor U24273 (N_24273,N_23616,N_23335);
nand U24274 (N_24274,N_23521,N_23642);
nor U24275 (N_24275,N_23767,N_23669);
and U24276 (N_24276,N_23393,N_23990);
xor U24277 (N_24277,N_23585,N_23983);
nor U24278 (N_24278,N_23877,N_23655);
nand U24279 (N_24279,N_23912,N_23769);
or U24280 (N_24280,N_23475,N_23837);
and U24281 (N_24281,N_23962,N_23805);
xnor U24282 (N_24282,N_23148,N_23793);
nor U24283 (N_24283,N_23209,N_23258);
nand U24284 (N_24284,N_23365,N_23444);
nand U24285 (N_24285,N_23541,N_23008);
or U24286 (N_24286,N_23349,N_23910);
nand U24287 (N_24287,N_23975,N_23963);
nor U24288 (N_24288,N_23069,N_23173);
and U24289 (N_24289,N_23324,N_23369);
and U24290 (N_24290,N_23750,N_23968);
or U24291 (N_24291,N_23423,N_23268);
or U24292 (N_24292,N_23245,N_23533);
nor U24293 (N_24293,N_23185,N_23534);
and U24294 (N_24294,N_23286,N_23112);
nand U24295 (N_24295,N_23226,N_23500);
nor U24296 (N_24296,N_23443,N_23788);
or U24297 (N_24297,N_23705,N_23726);
and U24298 (N_24298,N_23599,N_23141);
and U24299 (N_24299,N_23356,N_23825);
nor U24300 (N_24300,N_23844,N_23582);
nand U24301 (N_24301,N_23413,N_23957);
and U24302 (N_24302,N_23454,N_23909);
nand U24303 (N_24303,N_23416,N_23255);
nor U24304 (N_24304,N_23779,N_23768);
or U24305 (N_24305,N_23420,N_23383);
nand U24306 (N_24306,N_23384,N_23006);
and U24307 (N_24307,N_23134,N_23352);
nor U24308 (N_24308,N_23003,N_23355);
xnor U24309 (N_24309,N_23681,N_23159);
xor U24310 (N_24310,N_23035,N_23775);
nor U24311 (N_24311,N_23059,N_23556);
nand U24312 (N_24312,N_23111,N_23565);
nor U24313 (N_24313,N_23596,N_23256);
nor U24314 (N_24314,N_23696,N_23740);
xor U24315 (N_24315,N_23417,N_23812);
nor U24316 (N_24316,N_23546,N_23079);
or U24317 (N_24317,N_23736,N_23507);
xnor U24318 (N_24318,N_23978,N_23307);
nor U24319 (N_24319,N_23068,N_23194);
nand U24320 (N_24320,N_23744,N_23123);
or U24321 (N_24321,N_23755,N_23243);
xor U24322 (N_24322,N_23710,N_23009);
and U24323 (N_24323,N_23337,N_23292);
xor U24324 (N_24324,N_23415,N_23593);
nor U24325 (N_24325,N_23807,N_23206);
and U24326 (N_24326,N_23995,N_23713);
nand U24327 (N_24327,N_23139,N_23118);
xor U24328 (N_24328,N_23433,N_23104);
or U24329 (N_24329,N_23276,N_23992);
and U24330 (N_24330,N_23361,N_23459);
nand U24331 (N_24331,N_23442,N_23915);
xor U24332 (N_24332,N_23219,N_23941);
and U24333 (N_24333,N_23162,N_23044);
nand U24334 (N_24334,N_23848,N_23147);
or U24335 (N_24335,N_23373,N_23000);
or U24336 (N_24336,N_23815,N_23911);
nand U24337 (N_24337,N_23290,N_23819);
xnor U24338 (N_24338,N_23721,N_23092);
nand U24339 (N_24339,N_23175,N_23461);
and U24340 (N_24340,N_23239,N_23943);
nand U24341 (N_24341,N_23073,N_23789);
nor U24342 (N_24342,N_23577,N_23296);
nand U24343 (N_24343,N_23687,N_23784);
nor U24344 (N_24344,N_23180,N_23976);
nor U24345 (N_24345,N_23191,N_23429);
or U24346 (N_24346,N_23580,N_23572);
nand U24347 (N_24347,N_23849,N_23722);
nand U24348 (N_24348,N_23958,N_23542);
xor U24349 (N_24349,N_23996,N_23587);
nor U24350 (N_24350,N_23871,N_23323);
xnor U24351 (N_24351,N_23200,N_23007);
and U24352 (N_24352,N_23522,N_23458);
and U24353 (N_24353,N_23967,N_23659);
and U24354 (N_24354,N_23811,N_23583);
or U24355 (N_24355,N_23272,N_23042);
nand U24356 (N_24356,N_23304,N_23670);
xnor U24357 (N_24357,N_23937,N_23701);
and U24358 (N_24358,N_23269,N_23039);
nand U24359 (N_24359,N_23297,N_23488);
or U24360 (N_24360,N_23389,N_23242);
nand U24361 (N_24361,N_23980,N_23880);
or U24362 (N_24362,N_23876,N_23575);
nor U24363 (N_24363,N_23601,N_23796);
and U24364 (N_24364,N_23182,N_23250);
or U24365 (N_24365,N_23405,N_23037);
xor U24366 (N_24366,N_23317,N_23508);
and U24367 (N_24367,N_23081,N_23440);
nand U24368 (N_24368,N_23761,N_23347);
nor U24369 (N_24369,N_23486,N_23558);
and U24370 (N_24370,N_23350,N_23348);
and U24371 (N_24371,N_23605,N_23388);
and U24372 (N_24372,N_23262,N_23603);
or U24373 (N_24373,N_23644,N_23218);
xnor U24374 (N_24374,N_23804,N_23054);
xnor U24375 (N_24375,N_23529,N_23597);
nand U24376 (N_24376,N_23238,N_23810);
xnor U24377 (N_24377,N_23421,N_23018);
and U24378 (N_24378,N_23640,N_23116);
xnor U24379 (N_24379,N_23077,N_23763);
nor U24380 (N_24380,N_23594,N_23845);
and U24381 (N_24381,N_23766,N_23783);
and U24382 (N_24382,N_23432,N_23151);
nand U24383 (N_24383,N_23568,N_23892);
and U24384 (N_24384,N_23611,N_23919);
or U24385 (N_24385,N_23998,N_23800);
nor U24386 (N_24386,N_23694,N_23861);
nor U24387 (N_24387,N_23653,N_23633);
or U24388 (N_24388,N_23656,N_23537);
or U24389 (N_24389,N_23688,N_23288);
nand U24390 (N_24390,N_23808,N_23367);
xnor U24391 (N_24391,N_23306,N_23802);
xor U24392 (N_24392,N_23491,N_23620);
nor U24393 (N_24393,N_23410,N_23828);
nor U24394 (N_24394,N_23327,N_23133);
nand U24395 (N_24395,N_23926,N_23557);
nand U24396 (N_24396,N_23181,N_23579);
xor U24397 (N_24397,N_23680,N_23249);
nand U24398 (N_24398,N_23495,N_23229);
nor U24399 (N_24399,N_23406,N_23548);
or U24400 (N_24400,N_23936,N_23714);
nor U24401 (N_24401,N_23754,N_23002);
and U24402 (N_24402,N_23724,N_23749);
or U24403 (N_24403,N_23863,N_23643);
nor U24404 (N_24404,N_23884,N_23684);
and U24405 (N_24405,N_23569,N_23823);
and U24406 (N_24406,N_23723,N_23564);
and U24407 (N_24407,N_23371,N_23310);
and U24408 (N_24408,N_23331,N_23368);
nor U24409 (N_24409,N_23387,N_23818);
xnor U24410 (N_24410,N_23186,N_23144);
nand U24411 (N_24411,N_23224,N_23047);
and U24412 (N_24412,N_23717,N_23248);
and U24413 (N_24413,N_23900,N_23913);
and U24414 (N_24414,N_23137,N_23174);
or U24415 (N_24415,N_23210,N_23158);
nand U24416 (N_24416,N_23080,N_23519);
or U24417 (N_24417,N_23799,N_23746);
xnor U24418 (N_24418,N_23883,N_23999);
xor U24419 (N_24419,N_23076,N_23952);
and U24420 (N_24420,N_23765,N_23747);
nand U24421 (N_24421,N_23630,N_23257);
nand U24422 (N_24422,N_23729,N_23114);
and U24423 (N_24423,N_23216,N_23961);
nand U24424 (N_24424,N_23270,N_23612);
or U24425 (N_24425,N_23045,N_23333);
nand U24426 (N_24426,N_23403,N_23102);
xor U24427 (N_24427,N_23830,N_23192);
nand U24428 (N_24428,N_23623,N_23165);
xor U24429 (N_24429,N_23110,N_23464);
nor U24430 (N_24430,N_23418,N_23411);
or U24431 (N_24431,N_23907,N_23795);
xor U24432 (N_24432,N_23662,N_23512);
nand U24433 (N_24433,N_23683,N_23316);
and U24434 (N_24434,N_23293,N_23869);
nand U24435 (N_24435,N_23725,N_23467);
nor U24436 (N_24436,N_23354,N_23979);
nor U24437 (N_24437,N_23951,N_23917);
and U24438 (N_24438,N_23866,N_23840);
xor U24439 (N_24439,N_23010,N_23332);
nand U24440 (N_24440,N_23153,N_23330);
or U24441 (N_24441,N_23820,N_23834);
nor U24442 (N_24442,N_23551,N_23012);
or U24443 (N_24443,N_23857,N_23140);
nor U24444 (N_24444,N_23932,N_23346);
nor U24445 (N_24445,N_23631,N_23380);
nand U24446 (N_24446,N_23686,N_23974);
or U24447 (N_24447,N_23889,N_23024);
or U24448 (N_24448,N_23547,N_23228);
and U24449 (N_24449,N_23885,N_23720);
or U24450 (N_24450,N_23574,N_23050);
and U24451 (N_24451,N_23586,N_23562);
nand U24452 (N_24452,N_23473,N_23956);
xnor U24453 (N_24453,N_23138,N_23083);
nand U24454 (N_24454,N_23129,N_23878);
or U24455 (N_24455,N_23972,N_23581);
xnor U24456 (N_24456,N_23177,N_23320);
nand U24457 (N_24457,N_23982,N_23357);
nor U24458 (N_24458,N_23298,N_23099);
or U24459 (N_24459,N_23567,N_23658);
nor U24460 (N_24460,N_23621,N_23609);
and U24461 (N_24461,N_23264,N_23160);
nor U24462 (N_24462,N_23600,N_23526);
nor U24463 (N_24463,N_23875,N_23778);
or U24464 (N_24464,N_23056,N_23989);
nand U24465 (N_24465,N_23051,N_23065);
xnor U24466 (N_24466,N_23471,N_23895);
nor U24467 (N_24467,N_23033,N_23027);
and U24468 (N_24468,N_23924,N_23674);
or U24469 (N_24469,N_23095,N_23552);
or U24470 (N_24470,N_23374,N_23015);
or U24471 (N_24471,N_23013,N_23617);
nand U24472 (N_24472,N_23822,N_23457);
or U24473 (N_24473,N_23098,N_23312);
nand U24474 (N_24474,N_23856,N_23043);
nor U24475 (N_24475,N_23303,N_23456);
and U24476 (N_24476,N_23399,N_23149);
and U24477 (N_24477,N_23090,N_23657);
and U24478 (N_24478,N_23571,N_23666);
and U24479 (N_24479,N_23404,N_23632);
xor U24480 (N_24480,N_23977,N_23712);
or U24481 (N_24481,N_23928,N_23809);
xnor U24482 (N_24482,N_23199,N_23966);
or U24483 (N_24483,N_23854,N_23485);
xor U24484 (N_24484,N_23973,N_23930);
nand U24485 (N_24485,N_23525,N_23291);
nand U24486 (N_24486,N_23523,N_23340);
nand U24487 (N_24487,N_23196,N_23074);
nand U24488 (N_24488,N_23549,N_23496);
nand U24489 (N_24489,N_23685,N_23872);
nor U24490 (N_24490,N_23752,N_23510);
nor U24491 (N_24491,N_23776,N_23536);
xor U24492 (N_24492,N_23731,N_23447);
and U24493 (N_24493,N_23119,N_23667);
and U24494 (N_24494,N_23451,N_23905);
and U24495 (N_24495,N_23078,N_23592);
nor U24496 (N_24496,N_23360,N_23217);
xor U24497 (N_24497,N_23960,N_23584);
xor U24498 (N_24498,N_23893,N_23408);
nor U24499 (N_24499,N_23890,N_23376);
nand U24500 (N_24500,N_23690,N_23074);
xor U24501 (N_24501,N_23237,N_23021);
nor U24502 (N_24502,N_23170,N_23894);
nor U24503 (N_24503,N_23750,N_23296);
or U24504 (N_24504,N_23876,N_23738);
nor U24505 (N_24505,N_23507,N_23000);
nand U24506 (N_24506,N_23663,N_23560);
nor U24507 (N_24507,N_23728,N_23832);
xor U24508 (N_24508,N_23477,N_23212);
and U24509 (N_24509,N_23157,N_23471);
nor U24510 (N_24510,N_23979,N_23723);
nand U24511 (N_24511,N_23114,N_23671);
or U24512 (N_24512,N_23590,N_23620);
nor U24513 (N_24513,N_23835,N_23260);
and U24514 (N_24514,N_23922,N_23968);
xor U24515 (N_24515,N_23545,N_23654);
xnor U24516 (N_24516,N_23877,N_23042);
nand U24517 (N_24517,N_23675,N_23823);
nand U24518 (N_24518,N_23521,N_23166);
nor U24519 (N_24519,N_23678,N_23340);
and U24520 (N_24520,N_23035,N_23347);
nor U24521 (N_24521,N_23606,N_23730);
nand U24522 (N_24522,N_23891,N_23255);
nor U24523 (N_24523,N_23744,N_23361);
xnor U24524 (N_24524,N_23818,N_23661);
or U24525 (N_24525,N_23308,N_23533);
and U24526 (N_24526,N_23561,N_23055);
or U24527 (N_24527,N_23419,N_23605);
and U24528 (N_24528,N_23239,N_23830);
nor U24529 (N_24529,N_23620,N_23514);
nor U24530 (N_24530,N_23469,N_23987);
or U24531 (N_24531,N_23119,N_23219);
nand U24532 (N_24532,N_23353,N_23151);
and U24533 (N_24533,N_23337,N_23892);
nor U24534 (N_24534,N_23224,N_23508);
nand U24535 (N_24535,N_23854,N_23221);
or U24536 (N_24536,N_23594,N_23144);
xnor U24537 (N_24537,N_23981,N_23239);
nor U24538 (N_24538,N_23383,N_23337);
xor U24539 (N_24539,N_23458,N_23687);
nand U24540 (N_24540,N_23855,N_23748);
or U24541 (N_24541,N_23291,N_23479);
or U24542 (N_24542,N_23298,N_23950);
nor U24543 (N_24543,N_23260,N_23591);
nor U24544 (N_24544,N_23800,N_23825);
xnor U24545 (N_24545,N_23515,N_23335);
nor U24546 (N_24546,N_23122,N_23070);
nor U24547 (N_24547,N_23387,N_23472);
or U24548 (N_24548,N_23424,N_23490);
nor U24549 (N_24549,N_23499,N_23178);
nor U24550 (N_24550,N_23958,N_23409);
or U24551 (N_24551,N_23397,N_23960);
nand U24552 (N_24552,N_23693,N_23436);
nand U24553 (N_24553,N_23978,N_23178);
nand U24554 (N_24554,N_23056,N_23892);
nor U24555 (N_24555,N_23868,N_23796);
and U24556 (N_24556,N_23745,N_23274);
or U24557 (N_24557,N_23740,N_23891);
xnor U24558 (N_24558,N_23198,N_23727);
nor U24559 (N_24559,N_23256,N_23772);
xnor U24560 (N_24560,N_23208,N_23568);
nand U24561 (N_24561,N_23533,N_23573);
xor U24562 (N_24562,N_23100,N_23633);
nand U24563 (N_24563,N_23833,N_23292);
or U24564 (N_24564,N_23117,N_23316);
nor U24565 (N_24565,N_23034,N_23179);
nand U24566 (N_24566,N_23494,N_23330);
nand U24567 (N_24567,N_23482,N_23560);
xnor U24568 (N_24568,N_23670,N_23779);
and U24569 (N_24569,N_23016,N_23774);
xor U24570 (N_24570,N_23247,N_23936);
xnor U24571 (N_24571,N_23572,N_23033);
xor U24572 (N_24572,N_23391,N_23170);
xor U24573 (N_24573,N_23725,N_23938);
nand U24574 (N_24574,N_23191,N_23610);
nor U24575 (N_24575,N_23952,N_23612);
xnor U24576 (N_24576,N_23008,N_23236);
xor U24577 (N_24577,N_23233,N_23707);
nor U24578 (N_24578,N_23444,N_23564);
xnor U24579 (N_24579,N_23110,N_23770);
or U24580 (N_24580,N_23330,N_23438);
nor U24581 (N_24581,N_23085,N_23469);
nand U24582 (N_24582,N_23717,N_23772);
nor U24583 (N_24583,N_23807,N_23047);
nand U24584 (N_24584,N_23419,N_23893);
nor U24585 (N_24585,N_23071,N_23315);
nand U24586 (N_24586,N_23826,N_23246);
or U24587 (N_24587,N_23895,N_23279);
nand U24588 (N_24588,N_23252,N_23267);
and U24589 (N_24589,N_23908,N_23731);
nor U24590 (N_24590,N_23949,N_23055);
nand U24591 (N_24591,N_23801,N_23982);
and U24592 (N_24592,N_23225,N_23080);
nor U24593 (N_24593,N_23338,N_23104);
xor U24594 (N_24594,N_23625,N_23802);
xnor U24595 (N_24595,N_23923,N_23806);
xor U24596 (N_24596,N_23682,N_23482);
and U24597 (N_24597,N_23004,N_23332);
and U24598 (N_24598,N_23657,N_23774);
and U24599 (N_24599,N_23664,N_23848);
nor U24600 (N_24600,N_23932,N_23651);
nand U24601 (N_24601,N_23317,N_23890);
nand U24602 (N_24602,N_23360,N_23420);
nor U24603 (N_24603,N_23885,N_23537);
or U24604 (N_24604,N_23437,N_23295);
nand U24605 (N_24605,N_23615,N_23249);
nor U24606 (N_24606,N_23700,N_23984);
xnor U24607 (N_24607,N_23365,N_23268);
or U24608 (N_24608,N_23998,N_23997);
nand U24609 (N_24609,N_23447,N_23349);
nor U24610 (N_24610,N_23722,N_23848);
and U24611 (N_24611,N_23829,N_23497);
nand U24612 (N_24612,N_23189,N_23937);
or U24613 (N_24613,N_23684,N_23716);
xnor U24614 (N_24614,N_23990,N_23028);
nand U24615 (N_24615,N_23901,N_23286);
and U24616 (N_24616,N_23129,N_23836);
and U24617 (N_24617,N_23606,N_23651);
xor U24618 (N_24618,N_23742,N_23873);
or U24619 (N_24619,N_23581,N_23843);
and U24620 (N_24620,N_23247,N_23114);
or U24621 (N_24621,N_23699,N_23158);
or U24622 (N_24622,N_23277,N_23180);
or U24623 (N_24623,N_23863,N_23171);
nand U24624 (N_24624,N_23413,N_23603);
xnor U24625 (N_24625,N_23375,N_23549);
nor U24626 (N_24626,N_23346,N_23709);
nor U24627 (N_24627,N_23929,N_23113);
nand U24628 (N_24628,N_23114,N_23897);
nand U24629 (N_24629,N_23138,N_23115);
and U24630 (N_24630,N_23021,N_23803);
and U24631 (N_24631,N_23701,N_23588);
nand U24632 (N_24632,N_23883,N_23149);
xor U24633 (N_24633,N_23839,N_23864);
nor U24634 (N_24634,N_23415,N_23809);
nand U24635 (N_24635,N_23639,N_23991);
xor U24636 (N_24636,N_23052,N_23748);
nand U24637 (N_24637,N_23189,N_23076);
or U24638 (N_24638,N_23536,N_23664);
nand U24639 (N_24639,N_23404,N_23618);
and U24640 (N_24640,N_23207,N_23797);
and U24641 (N_24641,N_23192,N_23897);
xor U24642 (N_24642,N_23993,N_23778);
nand U24643 (N_24643,N_23750,N_23978);
nor U24644 (N_24644,N_23334,N_23551);
or U24645 (N_24645,N_23867,N_23825);
or U24646 (N_24646,N_23936,N_23925);
nor U24647 (N_24647,N_23856,N_23341);
or U24648 (N_24648,N_23806,N_23576);
xor U24649 (N_24649,N_23978,N_23239);
and U24650 (N_24650,N_23947,N_23816);
or U24651 (N_24651,N_23916,N_23867);
and U24652 (N_24652,N_23338,N_23178);
and U24653 (N_24653,N_23775,N_23387);
or U24654 (N_24654,N_23755,N_23735);
or U24655 (N_24655,N_23953,N_23606);
nor U24656 (N_24656,N_23955,N_23108);
and U24657 (N_24657,N_23224,N_23792);
nor U24658 (N_24658,N_23099,N_23847);
or U24659 (N_24659,N_23406,N_23502);
nand U24660 (N_24660,N_23254,N_23146);
nor U24661 (N_24661,N_23749,N_23593);
xnor U24662 (N_24662,N_23650,N_23790);
and U24663 (N_24663,N_23320,N_23863);
and U24664 (N_24664,N_23548,N_23329);
nand U24665 (N_24665,N_23584,N_23355);
nand U24666 (N_24666,N_23853,N_23005);
nor U24667 (N_24667,N_23634,N_23404);
xor U24668 (N_24668,N_23870,N_23781);
xor U24669 (N_24669,N_23160,N_23406);
or U24670 (N_24670,N_23360,N_23369);
nand U24671 (N_24671,N_23595,N_23643);
nor U24672 (N_24672,N_23596,N_23329);
and U24673 (N_24673,N_23761,N_23542);
or U24674 (N_24674,N_23757,N_23664);
or U24675 (N_24675,N_23042,N_23534);
nand U24676 (N_24676,N_23102,N_23475);
or U24677 (N_24677,N_23600,N_23991);
nor U24678 (N_24678,N_23217,N_23595);
nor U24679 (N_24679,N_23199,N_23054);
and U24680 (N_24680,N_23904,N_23136);
or U24681 (N_24681,N_23532,N_23161);
nand U24682 (N_24682,N_23869,N_23172);
and U24683 (N_24683,N_23979,N_23660);
xor U24684 (N_24684,N_23263,N_23895);
nor U24685 (N_24685,N_23858,N_23825);
nor U24686 (N_24686,N_23615,N_23245);
nand U24687 (N_24687,N_23421,N_23191);
nor U24688 (N_24688,N_23954,N_23249);
and U24689 (N_24689,N_23023,N_23715);
nor U24690 (N_24690,N_23555,N_23791);
nor U24691 (N_24691,N_23929,N_23014);
xor U24692 (N_24692,N_23548,N_23560);
or U24693 (N_24693,N_23329,N_23317);
or U24694 (N_24694,N_23319,N_23355);
nor U24695 (N_24695,N_23140,N_23684);
or U24696 (N_24696,N_23290,N_23921);
and U24697 (N_24697,N_23401,N_23024);
nand U24698 (N_24698,N_23100,N_23340);
xor U24699 (N_24699,N_23459,N_23681);
and U24700 (N_24700,N_23074,N_23305);
or U24701 (N_24701,N_23472,N_23004);
xor U24702 (N_24702,N_23866,N_23914);
xor U24703 (N_24703,N_23591,N_23835);
xor U24704 (N_24704,N_23481,N_23895);
and U24705 (N_24705,N_23944,N_23834);
nand U24706 (N_24706,N_23033,N_23258);
nor U24707 (N_24707,N_23898,N_23531);
nor U24708 (N_24708,N_23655,N_23085);
nand U24709 (N_24709,N_23497,N_23847);
nor U24710 (N_24710,N_23676,N_23975);
nand U24711 (N_24711,N_23476,N_23160);
nor U24712 (N_24712,N_23928,N_23331);
or U24713 (N_24713,N_23910,N_23273);
nand U24714 (N_24714,N_23609,N_23197);
nor U24715 (N_24715,N_23540,N_23231);
nor U24716 (N_24716,N_23376,N_23132);
nand U24717 (N_24717,N_23063,N_23961);
xnor U24718 (N_24718,N_23521,N_23563);
and U24719 (N_24719,N_23657,N_23174);
nor U24720 (N_24720,N_23896,N_23816);
and U24721 (N_24721,N_23646,N_23666);
and U24722 (N_24722,N_23358,N_23698);
and U24723 (N_24723,N_23488,N_23977);
xnor U24724 (N_24724,N_23156,N_23139);
and U24725 (N_24725,N_23863,N_23027);
nor U24726 (N_24726,N_23278,N_23317);
xor U24727 (N_24727,N_23226,N_23169);
and U24728 (N_24728,N_23355,N_23486);
nand U24729 (N_24729,N_23570,N_23323);
nor U24730 (N_24730,N_23158,N_23162);
or U24731 (N_24731,N_23810,N_23606);
xor U24732 (N_24732,N_23014,N_23432);
nand U24733 (N_24733,N_23491,N_23062);
xor U24734 (N_24734,N_23609,N_23433);
nand U24735 (N_24735,N_23495,N_23460);
xor U24736 (N_24736,N_23849,N_23065);
or U24737 (N_24737,N_23837,N_23737);
or U24738 (N_24738,N_23856,N_23193);
or U24739 (N_24739,N_23076,N_23298);
nor U24740 (N_24740,N_23729,N_23477);
nand U24741 (N_24741,N_23402,N_23235);
or U24742 (N_24742,N_23993,N_23939);
nand U24743 (N_24743,N_23076,N_23718);
and U24744 (N_24744,N_23901,N_23873);
xnor U24745 (N_24745,N_23167,N_23777);
or U24746 (N_24746,N_23347,N_23008);
or U24747 (N_24747,N_23203,N_23919);
nor U24748 (N_24748,N_23972,N_23311);
and U24749 (N_24749,N_23157,N_23601);
nand U24750 (N_24750,N_23960,N_23607);
and U24751 (N_24751,N_23380,N_23547);
or U24752 (N_24752,N_23870,N_23314);
xor U24753 (N_24753,N_23810,N_23128);
nand U24754 (N_24754,N_23137,N_23055);
xnor U24755 (N_24755,N_23984,N_23166);
and U24756 (N_24756,N_23401,N_23082);
and U24757 (N_24757,N_23156,N_23113);
and U24758 (N_24758,N_23331,N_23934);
xnor U24759 (N_24759,N_23561,N_23740);
nand U24760 (N_24760,N_23024,N_23400);
and U24761 (N_24761,N_23006,N_23113);
nand U24762 (N_24762,N_23347,N_23514);
and U24763 (N_24763,N_23667,N_23463);
or U24764 (N_24764,N_23326,N_23922);
nor U24765 (N_24765,N_23961,N_23899);
nand U24766 (N_24766,N_23172,N_23612);
nand U24767 (N_24767,N_23910,N_23209);
or U24768 (N_24768,N_23342,N_23424);
and U24769 (N_24769,N_23542,N_23063);
and U24770 (N_24770,N_23025,N_23279);
and U24771 (N_24771,N_23422,N_23644);
or U24772 (N_24772,N_23336,N_23746);
nor U24773 (N_24773,N_23134,N_23819);
nor U24774 (N_24774,N_23423,N_23547);
nand U24775 (N_24775,N_23559,N_23050);
or U24776 (N_24776,N_23337,N_23617);
and U24777 (N_24777,N_23174,N_23352);
nor U24778 (N_24778,N_23563,N_23152);
nand U24779 (N_24779,N_23420,N_23255);
and U24780 (N_24780,N_23838,N_23056);
nand U24781 (N_24781,N_23308,N_23367);
and U24782 (N_24782,N_23774,N_23797);
nand U24783 (N_24783,N_23255,N_23498);
xor U24784 (N_24784,N_23777,N_23604);
and U24785 (N_24785,N_23261,N_23567);
nor U24786 (N_24786,N_23071,N_23642);
nand U24787 (N_24787,N_23501,N_23920);
nand U24788 (N_24788,N_23345,N_23171);
nand U24789 (N_24789,N_23788,N_23636);
nor U24790 (N_24790,N_23210,N_23004);
nand U24791 (N_24791,N_23712,N_23082);
nand U24792 (N_24792,N_23789,N_23571);
and U24793 (N_24793,N_23330,N_23527);
and U24794 (N_24794,N_23246,N_23919);
and U24795 (N_24795,N_23993,N_23592);
or U24796 (N_24796,N_23036,N_23801);
nor U24797 (N_24797,N_23015,N_23433);
or U24798 (N_24798,N_23376,N_23383);
and U24799 (N_24799,N_23841,N_23721);
xnor U24800 (N_24800,N_23887,N_23902);
or U24801 (N_24801,N_23723,N_23353);
nor U24802 (N_24802,N_23288,N_23765);
nor U24803 (N_24803,N_23900,N_23470);
and U24804 (N_24804,N_23918,N_23869);
or U24805 (N_24805,N_23036,N_23234);
nand U24806 (N_24806,N_23958,N_23200);
nor U24807 (N_24807,N_23368,N_23283);
or U24808 (N_24808,N_23766,N_23389);
nor U24809 (N_24809,N_23114,N_23270);
xor U24810 (N_24810,N_23977,N_23238);
xor U24811 (N_24811,N_23116,N_23988);
nand U24812 (N_24812,N_23389,N_23977);
xnor U24813 (N_24813,N_23072,N_23190);
and U24814 (N_24814,N_23016,N_23435);
xnor U24815 (N_24815,N_23626,N_23324);
nand U24816 (N_24816,N_23679,N_23148);
or U24817 (N_24817,N_23828,N_23137);
or U24818 (N_24818,N_23781,N_23844);
and U24819 (N_24819,N_23141,N_23449);
nand U24820 (N_24820,N_23135,N_23834);
and U24821 (N_24821,N_23026,N_23469);
xor U24822 (N_24822,N_23193,N_23454);
or U24823 (N_24823,N_23873,N_23262);
nor U24824 (N_24824,N_23404,N_23976);
or U24825 (N_24825,N_23529,N_23287);
and U24826 (N_24826,N_23834,N_23411);
nand U24827 (N_24827,N_23216,N_23077);
nor U24828 (N_24828,N_23934,N_23737);
nor U24829 (N_24829,N_23532,N_23365);
nand U24830 (N_24830,N_23140,N_23707);
or U24831 (N_24831,N_23156,N_23501);
and U24832 (N_24832,N_23177,N_23810);
nand U24833 (N_24833,N_23286,N_23356);
and U24834 (N_24834,N_23190,N_23657);
nor U24835 (N_24835,N_23784,N_23146);
and U24836 (N_24836,N_23283,N_23657);
nor U24837 (N_24837,N_23141,N_23180);
xor U24838 (N_24838,N_23350,N_23380);
or U24839 (N_24839,N_23336,N_23228);
and U24840 (N_24840,N_23684,N_23248);
and U24841 (N_24841,N_23953,N_23828);
nand U24842 (N_24842,N_23498,N_23615);
or U24843 (N_24843,N_23971,N_23602);
nor U24844 (N_24844,N_23705,N_23054);
nand U24845 (N_24845,N_23925,N_23389);
or U24846 (N_24846,N_23586,N_23324);
nor U24847 (N_24847,N_23327,N_23111);
xnor U24848 (N_24848,N_23645,N_23159);
xor U24849 (N_24849,N_23085,N_23343);
nand U24850 (N_24850,N_23843,N_23265);
xnor U24851 (N_24851,N_23078,N_23340);
nand U24852 (N_24852,N_23850,N_23598);
nor U24853 (N_24853,N_23360,N_23039);
xor U24854 (N_24854,N_23576,N_23663);
nand U24855 (N_24855,N_23557,N_23157);
xnor U24856 (N_24856,N_23477,N_23076);
nand U24857 (N_24857,N_23712,N_23435);
and U24858 (N_24858,N_23632,N_23852);
or U24859 (N_24859,N_23866,N_23126);
or U24860 (N_24860,N_23044,N_23670);
or U24861 (N_24861,N_23020,N_23350);
xor U24862 (N_24862,N_23708,N_23213);
nor U24863 (N_24863,N_23496,N_23024);
nand U24864 (N_24864,N_23563,N_23690);
and U24865 (N_24865,N_23031,N_23456);
nand U24866 (N_24866,N_23225,N_23079);
nor U24867 (N_24867,N_23358,N_23162);
nand U24868 (N_24868,N_23039,N_23333);
xnor U24869 (N_24869,N_23637,N_23305);
nand U24870 (N_24870,N_23372,N_23393);
xnor U24871 (N_24871,N_23309,N_23118);
xor U24872 (N_24872,N_23851,N_23486);
and U24873 (N_24873,N_23262,N_23342);
nor U24874 (N_24874,N_23970,N_23370);
nor U24875 (N_24875,N_23182,N_23343);
nor U24876 (N_24876,N_23989,N_23526);
or U24877 (N_24877,N_23800,N_23771);
nor U24878 (N_24878,N_23616,N_23196);
and U24879 (N_24879,N_23913,N_23564);
nand U24880 (N_24880,N_23085,N_23948);
nor U24881 (N_24881,N_23587,N_23240);
nor U24882 (N_24882,N_23424,N_23649);
and U24883 (N_24883,N_23554,N_23257);
nor U24884 (N_24884,N_23592,N_23458);
nand U24885 (N_24885,N_23000,N_23138);
nand U24886 (N_24886,N_23595,N_23111);
or U24887 (N_24887,N_23769,N_23175);
or U24888 (N_24888,N_23264,N_23817);
xnor U24889 (N_24889,N_23761,N_23775);
and U24890 (N_24890,N_23969,N_23262);
and U24891 (N_24891,N_23609,N_23987);
or U24892 (N_24892,N_23114,N_23750);
nand U24893 (N_24893,N_23799,N_23673);
nand U24894 (N_24894,N_23620,N_23109);
nor U24895 (N_24895,N_23592,N_23051);
nand U24896 (N_24896,N_23204,N_23051);
or U24897 (N_24897,N_23341,N_23871);
and U24898 (N_24898,N_23709,N_23600);
and U24899 (N_24899,N_23537,N_23696);
nor U24900 (N_24900,N_23055,N_23242);
and U24901 (N_24901,N_23215,N_23451);
nor U24902 (N_24902,N_23506,N_23438);
nor U24903 (N_24903,N_23062,N_23327);
nor U24904 (N_24904,N_23592,N_23144);
nand U24905 (N_24905,N_23981,N_23249);
or U24906 (N_24906,N_23580,N_23810);
or U24907 (N_24907,N_23010,N_23485);
nand U24908 (N_24908,N_23864,N_23437);
or U24909 (N_24909,N_23757,N_23402);
and U24910 (N_24910,N_23643,N_23868);
nand U24911 (N_24911,N_23377,N_23023);
and U24912 (N_24912,N_23805,N_23019);
nand U24913 (N_24913,N_23830,N_23079);
and U24914 (N_24914,N_23108,N_23666);
xnor U24915 (N_24915,N_23557,N_23901);
or U24916 (N_24916,N_23297,N_23761);
xor U24917 (N_24917,N_23166,N_23203);
nor U24918 (N_24918,N_23763,N_23904);
xor U24919 (N_24919,N_23201,N_23200);
or U24920 (N_24920,N_23481,N_23052);
or U24921 (N_24921,N_23790,N_23142);
nand U24922 (N_24922,N_23406,N_23526);
xor U24923 (N_24923,N_23430,N_23124);
or U24924 (N_24924,N_23625,N_23478);
nor U24925 (N_24925,N_23319,N_23933);
xor U24926 (N_24926,N_23399,N_23030);
and U24927 (N_24927,N_23908,N_23019);
or U24928 (N_24928,N_23371,N_23540);
and U24929 (N_24929,N_23881,N_23781);
xor U24930 (N_24930,N_23807,N_23592);
and U24931 (N_24931,N_23446,N_23005);
xor U24932 (N_24932,N_23659,N_23436);
nand U24933 (N_24933,N_23878,N_23791);
or U24934 (N_24934,N_23826,N_23904);
or U24935 (N_24935,N_23424,N_23358);
nor U24936 (N_24936,N_23440,N_23579);
and U24937 (N_24937,N_23027,N_23543);
xor U24938 (N_24938,N_23753,N_23465);
or U24939 (N_24939,N_23096,N_23828);
nand U24940 (N_24940,N_23562,N_23542);
nand U24941 (N_24941,N_23647,N_23906);
and U24942 (N_24942,N_23375,N_23825);
and U24943 (N_24943,N_23652,N_23819);
nor U24944 (N_24944,N_23913,N_23217);
nor U24945 (N_24945,N_23410,N_23318);
nand U24946 (N_24946,N_23319,N_23070);
and U24947 (N_24947,N_23384,N_23675);
and U24948 (N_24948,N_23106,N_23327);
nor U24949 (N_24949,N_23321,N_23738);
or U24950 (N_24950,N_23823,N_23081);
nand U24951 (N_24951,N_23051,N_23290);
or U24952 (N_24952,N_23659,N_23744);
nand U24953 (N_24953,N_23499,N_23957);
nor U24954 (N_24954,N_23099,N_23286);
and U24955 (N_24955,N_23117,N_23865);
nor U24956 (N_24956,N_23293,N_23785);
xnor U24957 (N_24957,N_23848,N_23081);
and U24958 (N_24958,N_23536,N_23043);
xnor U24959 (N_24959,N_23499,N_23192);
nor U24960 (N_24960,N_23081,N_23362);
nand U24961 (N_24961,N_23511,N_23050);
or U24962 (N_24962,N_23460,N_23731);
or U24963 (N_24963,N_23709,N_23474);
nand U24964 (N_24964,N_23180,N_23338);
or U24965 (N_24965,N_23183,N_23499);
xnor U24966 (N_24966,N_23479,N_23831);
or U24967 (N_24967,N_23262,N_23396);
nor U24968 (N_24968,N_23438,N_23600);
or U24969 (N_24969,N_23735,N_23326);
or U24970 (N_24970,N_23396,N_23878);
or U24971 (N_24971,N_23352,N_23682);
or U24972 (N_24972,N_23033,N_23452);
and U24973 (N_24973,N_23038,N_23333);
and U24974 (N_24974,N_23877,N_23359);
nor U24975 (N_24975,N_23381,N_23794);
and U24976 (N_24976,N_23112,N_23619);
nand U24977 (N_24977,N_23588,N_23731);
and U24978 (N_24978,N_23309,N_23173);
or U24979 (N_24979,N_23614,N_23113);
nor U24980 (N_24980,N_23086,N_23912);
xnor U24981 (N_24981,N_23777,N_23482);
nand U24982 (N_24982,N_23564,N_23360);
nand U24983 (N_24983,N_23443,N_23281);
nor U24984 (N_24984,N_23342,N_23548);
and U24985 (N_24985,N_23668,N_23626);
nand U24986 (N_24986,N_23669,N_23640);
nor U24987 (N_24987,N_23208,N_23513);
or U24988 (N_24988,N_23501,N_23328);
nor U24989 (N_24989,N_23569,N_23842);
or U24990 (N_24990,N_23134,N_23644);
xnor U24991 (N_24991,N_23805,N_23954);
xor U24992 (N_24992,N_23628,N_23741);
xnor U24993 (N_24993,N_23192,N_23814);
nor U24994 (N_24994,N_23047,N_23694);
nor U24995 (N_24995,N_23977,N_23241);
and U24996 (N_24996,N_23560,N_23817);
or U24997 (N_24997,N_23208,N_23312);
xor U24998 (N_24998,N_23780,N_23026);
nand U24999 (N_24999,N_23698,N_23822);
xor UO_0 (O_0,N_24340,N_24897);
or UO_1 (O_1,N_24813,N_24935);
xnor UO_2 (O_2,N_24635,N_24148);
xor UO_3 (O_3,N_24481,N_24200);
xor UO_4 (O_4,N_24176,N_24109);
and UO_5 (O_5,N_24375,N_24927);
nand UO_6 (O_6,N_24325,N_24485);
and UO_7 (O_7,N_24968,N_24855);
nor UO_8 (O_8,N_24564,N_24226);
nand UO_9 (O_9,N_24419,N_24005);
nor UO_10 (O_10,N_24085,N_24364);
xnor UO_11 (O_11,N_24346,N_24812);
nand UO_12 (O_12,N_24929,N_24628);
nor UO_13 (O_13,N_24688,N_24700);
nand UO_14 (O_14,N_24772,N_24184);
and UO_15 (O_15,N_24951,N_24382);
nand UO_16 (O_16,N_24166,N_24095);
nand UO_17 (O_17,N_24482,N_24472);
and UO_18 (O_18,N_24724,N_24396);
nand UO_19 (O_19,N_24796,N_24163);
nor UO_20 (O_20,N_24222,N_24048);
nor UO_21 (O_21,N_24317,N_24742);
xor UO_22 (O_22,N_24969,N_24685);
xnor UO_23 (O_23,N_24411,N_24713);
and UO_24 (O_24,N_24064,N_24767);
xnor UO_25 (O_25,N_24517,N_24494);
xor UO_26 (O_26,N_24406,N_24634);
or UO_27 (O_27,N_24321,N_24050);
xor UO_28 (O_28,N_24535,N_24227);
and UO_29 (O_29,N_24750,N_24906);
xnor UO_30 (O_30,N_24316,N_24285);
xor UO_31 (O_31,N_24056,N_24502);
or UO_32 (O_32,N_24119,N_24255);
nor UO_33 (O_33,N_24695,N_24279);
and UO_34 (O_34,N_24033,N_24426);
nand UO_35 (O_35,N_24353,N_24577);
nor UO_36 (O_36,N_24116,N_24570);
nand UO_37 (O_37,N_24617,N_24299);
and UO_38 (O_38,N_24079,N_24246);
nand UO_39 (O_39,N_24687,N_24682);
xnor UO_40 (O_40,N_24066,N_24212);
nor UO_41 (O_41,N_24598,N_24548);
xor UO_42 (O_42,N_24083,N_24488);
or UO_43 (O_43,N_24618,N_24558);
xnor UO_44 (O_44,N_24276,N_24918);
and UO_45 (O_45,N_24169,N_24515);
and UO_46 (O_46,N_24017,N_24420);
nor UO_47 (O_47,N_24841,N_24689);
and UO_48 (O_48,N_24096,N_24057);
nand UO_49 (O_49,N_24547,N_24881);
nand UO_50 (O_50,N_24605,N_24757);
nor UO_51 (O_51,N_24082,N_24160);
and UO_52 (O_52,N_24916,N_24231);
or UO_53 (O_53,N_24985,N_24904);
xnor UO_54 (O_54,N_24320,N_24527);
or UO_55 (O_55,N_24500,N_24010);
nand UO_56 (O_56,N_24754,N_24770);
or UO_57 (O_57,N_24251,N_24891);
xnor UO_58 (O_58,N_24681,N_24671);
nor UO_59 (O_59,N_24940,N_24778);
xnor UO_60 (O_60,N_24442,N_24138);
nand UO_61 (O_61,N_24936,N_24505);
nand UO_62 (O_62,N_24704,N_24009);
xor UO_63 (O_63,N_24518,N_24070);
or UO_64 (O_64,N_24541,N_24567);
nand UO_65 (O_65,N_24125,N_24779);
xor UO_66 (O_66,N_24699,N_24270);
nor UO_67 (O_67,N_24571,N_24478);
nand UO_68 (O_68,N_24021,N_24871);
or UO_69 (O_69,N_24181,N_24859);
xor UO_70 (O_70,N_24984,N_24954);
xnor UO_71 (O_71,N_24911,N_24961);
or UO_72 (O_72,N_24344,N_24917);
nand UO_73 (O_73,N_24880,N_24072);
nor UO_74 (O_74,N_24458,N_24452);
or UO_75 (O_75,N_24361,N_24828);
and UO_76 (O_76,N_24823,N_24804);
xnor UO_77 (O_77,N_24188,N_24877);
xnor UO_78 (O_78,N_24496,N_24373);
and UO_79 (O_79,N_24701,N_24493);
nor UO_80 (O_80,N_24013,N_24221);
and UO_81 (O_81,N_24920,N_24797);
nor UO_82 (O_82,N_24622,N_24878);
and UO_83 (O_83,N_24947,N_24908);
xnor UO_84 (O_84,N_24683,N_24922);
xor UO_85 (O_85,N_24150,N_24736);
and UO_86 (O_86,N_24168,N_24213);
and UO_87 (O_87,N_24211,N_24606);
nor UO_88 (O_88,N_24412,N_24410);
nor UO_89 (O_89,N_24233,N_24789);
xnor UO_90 (O_90,N_24781,N_24768);
xnor UO_91 (O_91,N_24840,N_24582);
or UO_92 (O_92,N_24962,N_24029);
and UO_93 (O_93,N_24665,N_24381);
nand UO_94 (O_94,N_24413,N_24275);
nor UO_95 (O_95,N_24308,N_24332);
or UO_96 (O_96,N_24826,N_24012);
or UO_97 (O_97,N_24650,N_24195);
nand UO_98 (O_98,N_24845,N_24731);
nand UO_99 (O_99,N_24497,N_24347);
nand UO_100 (O_100,N_24937,N_24358);
and UO_101 (O_101,N_24106,N_24800);
nor UO_102 (O_102,N_24297,N_24436);
xnor UO_103 (O_103,N_24484,N_24374);
nand UO_104 (O_104,N_24851,N_24139);
or UO_105 (O_105,N_24171,N_24508);
or UO_106 (O_106,N_24730,N_24258);
nand UO_107 (O_107,N_24591,N_24283);
xnor UO_108 (O_108,N_24892,N_24210);
nor UO_109 (O_109,N_24471,N_24235);
xor UO_110 (O_110,N_24080,N_24763);
nand UO_111 (O_111,N_24025,N_24323);
nor UO_112 (O_112,N_24640,N_24630);
or UO_113 (O_113,N_24854,N_24870);
and UO_114 (O_114,N_24957,N_24161);
or UO_115 (O_115,N_24203,N_24749);
nor UO_116 (O_116,N_24745,N_24241);
and UO_117 (O_117,N_24561,N_24165);
and UO_118 (O_118,N_24128,N_24666);
and UO_119 (O_119,N_24130,N_24093);
and UO_120 (O_120,N_24696,N_24007);
and UO_121 (O_121,N_24026,N_24707);
or UO_122 (O_122,N_24926,N_24274);
or UO_123 (O_123,N_24456,N_24248);
nor UO_124 (O_124,N_24247,N_24782);
xor UO_125 (O_125,N_24549,N_24811);
xnor UO_126 (O_126,N_24566,N_24073);
or UO_127 (O_127,N_24022,N_24403);
or UO_128 (O_128,N_24584,N_24737);
and UO_129 (O_129,N_24291,N_24748);
xnor UO_130 (O_130,N_24014,N_24301);
or UO_131 (O_131,N_24495,N_24455);
and UO_132 (O_132,N_24016,N_24405);
xnor UO_133 (O_133,N_24239,N_24893);
xor UO_134 (O_134,N_24512,N_24821);
or UO_135 (O_135,N_24451,N_24977);
xnor UO_136 (O_136,N_24232,N_24620);
xor UO_137 (O_137,N_24397,N_24679);
and UO_138 (O_138,N_24199,N_24292);
xnor UO_139 (O_139,N_24694,N_24846);
nor UO_140 (O_140,N_24857,N_24611);
nand UO_141 (O_141,N_24525,N_24592);
nand UO_142 (O_142,N_24424,N_24417);
xor UO_143 (O_143,N_24914,N_24179);
or UO_144 (O_144,N_24253,N_24267);
or UO_145 (O_145,N_24649,N_24629);
and UO_146 (O_146,N_24595,N_24103);
nand UO_147 (O_147,N_24089,N_24147);
and UO_148 (O_148,N_24244,N_24579);
nand UO_149 (O_149,N_24313,N_24815);
xor UO_150 (O_150,N_24142,N_24980);
xnor UO_151 (O_151,N_24051,N_24581);
and UO_152 (O_152,N_24747,N_24967);
and UO_153 (O_153,N_24145,N_24334);
and UO_154 (O_154,N_24639,N_24047);
nor UO_155 (O_155,N_24479,N_24858);
nor UO_156 (O_156,N_24492,N_24583);
xnor UO_157 (O_157,N_24428,N_24949);
nand UO_158 (O_158,N_24834,N_24349);
or UO_159 (O_159,N_24438,N_24798);
and UO_160 (O_160,N_24625,N_24609);
nand UO_161 (O_161,N_24658,N_24467);
nand UO_162 (O_162,N_24603,N_24589);
and UO_163 (O_163,N_24551,N_24860);
or UO_164 (O_164,N_24766,N_24003);
and UO_165 (O_165,N_24069,N_24955);
nor UO_166 (O_166,N_24993,N_24769);
xnor UO_167 (O_167,N_24209,N_24764);
nor UO_168 (O_168,N_24623,N_24554);
nor UO_169 (O_169,N_24758,N_24557);
and UO_170 (O_170,N_24060,N_24787);
nor UO_171 (O_171,N_24612,N_24314);
and UO_172 (O_172,N_24296,N_24019);
xnor UO_173 (O_173,N_24336,N_24593);
or UO_174 (O_174,N_24569,N_24457);
xnor UO_175 (O_175,N_24979,N_24018);
and UO_176 (O_176,N_24883,N_24751);
nor UO_177 (O_177,N_24928,N_24616);
nor UO_178 (O_178,N_24943,N_24814);
nand UO_179 (O_179,N_24850,N_24229);
xor UO_180 (O_180,N_24157,N_24654);
or UO_181 (O_181,N_24712,N_24099);
nand UO_182 (O_182,N_24559,N_24646);
and UO_183 (O_183,N_24372,N_24365);
nand UO_184 (O_184,N_24453,N_24652);
xnor UO_185 (O_185,N_24727,N_24890);
nand UO_186 (O_186,N_24975,N_24674);
and UO_187 (O_187,N_24444,N_24068);
or UO_188 (O_188,N_24193,N_24636);
and UO_189 (O_189,N_24122,N_24035);
and UO_190 (O_190,N_24172,N_24454);
nand UO_191 (O_191,N_24034,N_24404);
and UO_192 (O_192,N_24348,N_24054);
nor UO_193 (O_193,N_24944,N_24948);
nand UO_194 (O_194,N_24820,N_24264);
and UO_195 (O_195,N_24809,N_24065);
and UO_196 (O_196,N_24486,N_24534);
and UO_197 (O_197,N_24038,N_24819);
or UO_198 (O_198,N_24434,N_24208);
nand UO_199 (O_199,N_24825,N_24450);
or UO_200 (O_200,N_24596,N_24907);
xor UO_201 (O_201,N_24847,N_24988);
nand UO_202 (O_202,N_24587,N_24714);
nor UO_203 (O_203,N_24164,N_24449);
nor UO_204 (O_204,N_24071,N_24115);
or UO_205 (O_205,N_24888,N_24670);
or UO_206 (O_206,N_24362,N_24537);
and UO_207 (O_207,N_24392,N_24565);
and UO_208 (O_208,N_24919,N_24990);
nand UO_209 (O_209,N_24705,N_24322);
nor UO_210 (O_210,N_24597,N_24153);
nand UO_211 (O_211,N_24894,N_24972);
nand UO_212 (O_212,N_24245,N_24111);
and UO_213 (O_213,N_24509,N_24205);
xor UO_214 (O_214,N_24389,N_24697);
nor UO_215 (O_215,N_24266,N_24744);
nor UO_216 (O_216,N_24844,N_24530);
or UO_217 (O_217,N_24271,N_24607);
nor UO_218 (O_218,N_24669,N_24873);
nor UO_219 (O_219,N_24415,N_24189);
or UO_220 (O_220,N_24831,N_24131);
and UO_221 (O_221,N_24884,N_24357);
and UO_222 (O_222,N_24086,N_24499);
nand UO_223 (O_223,N_24773,N_24159);
and UO_224 (O_224,N_24049,N_24141);
and UO_225 (O_225,N_24960,N_24715);
nand UO_226 (O_226,N_24576,N_24252);
or UO_227 (O_227,N_24204,N_24218);
xnor UO_228 (O_228,N_24108,N_24262);
or UO_229 (O_229,N_24522,N_24838);
and UO_230 (O_230,N_24761,N_24608);
nand UO_231 (O_231,N_24872,N_24938);
nand UO_232 (O_232,N_24808,N_24342);
nor UO_233 (O_233,N_24995,N_24638);
or UO_234 (O_234,N_24234,N_24501);
and UO_235 (O_235,N_24889,N_24986);
nor UO_236 (O_236,N_24028,N_24690);
nor UO_237 (O_237,N_24552,N_24945);
nand UO_238 (O_238,N_24536,N_24573);
nor UO_239 (O_239,N_24011,N_24864);
xor UO_240 (O_240,N_24799,N_24777);
and UO_241 (O_241,N_24925,N_24786);
and UO_242 (O_242,N_24818,N_24981);
or UO_243 (O_243,N_24709,N_24384);
or UO_244 (O_244,N_24101,N_24895);
and UO_245 (O_245,N_24100,N_24407);
nor UO_246 (O_246,N_24088,N_24989);
and UO_247 (O_247,N_24046,N_24642);
and UO_248 (O_248,N_24775,N_24243);
xnor UO_249 (O_249,N_24824,N_24513);
and UO_250 (O_250,N_24655,N_24331);
xnor UO_251 (O_251,N_24723,N_24600);
or UO_252 (O_252,N_24152,N_24575);
nor UO_253 (O_253,N_24958,N_24260);
nand UO_254 (O_254,N_24963,N_24946);
or UO_255 (O_255,N_24081,N_24303);
nor UO_256 (O_256,N_24335,N_24836);
xor UO_257 (O_257,N_24966,N_24752);
nor UO_258 (O_258,N_24601,N_24829);
nand UO_259 (O_259,N_24684,N_24563);
nand UO_260 (O_260,N_24237,N_24146);
xor UO_261 (O_261,N_24330,N_24341);
and UO_262 (O_262,N_24110,N_24753);
or UO_263 (O_263,N_24368,N_24439);
and UO_264 (O_264,N_24310,N_24923);
nand UO_265 (O_265,N_24273,N_24462);
and UO_266 (O_266,N_24466,N_24662);
or UO_267 (O_267,N_24098,N_24090);
nand UO_268 (O_268,N_24711,N_24776);
nor UO_269 (O_269,N_24540,N_24132);
or UO_270 (O_270,N_24097,N_24004);
nand UO_271 (O_271,N_24249,N_24350);
and UO_272 (O_272,N_24913,N_24343);
nand UO_273 (O_273,N_24491,N_24939);
and UO_274 (O_274,N_24293,N_24887);
nand UO_275 (O_275,N_24398,N_24610);
nand UO_276 (O_276,N_24852,N_24602);
xor UO_277 (O_277,N_24653,N_24528);
xor UO_278 (O_278,N_24214,N_24000);
nand UO_279 (O_279,N_24490,N_24498);
nor UO_280 (O_280,N_24514,N_24151);
or UO_281 (O_281,N_24521,N_24519);
and UO_282 (O_282,N_24127,N_24615);
and UO_283 (O_283,N_24287,N_24733);
nor UO_284 (O_284,N_24660,N_24738);
and UO_285 (O_285,N_24732,N_24366);
xnor UO_286 (O_286,N_24771,N_24399);
or UO_287 (O_287,N_24686,N_24394);
or UO_288 (O_288,N_24158,N_24312);
nand UO_289 (O_289,N_24459,N_24790);
and UO_290 (O_290,N_24942,N_24667);
and UO_291 (O_291,N_24144,N_24680);
nor UO_292 (O_292,N_24269,N_24043);
nand UO_293 (O_293,N_24041,N_24216);
nand UO_294 (O_294,N_24402,N_24386);
or UO_295 (O_295,N_24553,N_24959);
xnor UO_296 (O_296,N_24031,N_24794);
and UO_297 (O_297,N_24673,N_24126);
or UO_298 (O_298,N_24520,N_24228);
xnor UO_299 (O_299,N_24656,N_24862);
and UO_300 (O_300,N_24186,N_24061);
xor UO_301 (O_301,N_24734,N_24604);
nor UO_302 (O_302,N_24201,N_24102);
xor UO_303 (O_303,N_24867,N_24133);
and UO_304 (O_304,N_24706,N_24032);
nand UO_305 (O_305,N_24174,N_24370);
xor UO_306 (O_306,N_24698,N_24503);
and UO_307 (O_307,N_24924,N_24318);
and UO_308 (O_308,N_24915,N_24746);
nor UO_309 (O_309,N_24333,N_24268);
nor UO_310 (O_310,N_24037,N_24903);
or UO_311 (O_311,N_24676,N_24578);
nor UO_312 (O_312,N_24261,N_24044);
xor UO_313 (O_313,N_24632,N_24027);
xor UO_314 (O_314,N_24118,N_24105);
nor UO_315 (O_315,N_24934,N_24114);
nor UO_316 (O_316,N_24791,N_24162);
or UO_317 (O_317,N_24822,N_24516);
and UO_318 (O_318,N_24440,N_24997);
or UO_319 (O_319,N_24645,N_24780);
xor UO_320 (O_320,N_24816,N_24352);
xnor UO_321 (O_321,N_24277,N_24827);
nand UO_322 (O_322,N_24590,N_24124);
or UO_323 (O_323,N_24236,N_24477);
or UO_324 (O_324,N_24154,N_24801);
xnor UO_325 (O_325,N_24058,N_24288);
nor UO_326 (O_326,N_24902,N_24053);
nand UO_327 (O_327,N_24865,N_24351);
nor UO_328 (O_328,N_24722,N_24793);
nand UO_329 (O_329,N_24976,N_24401);
nand UO_330 (O_330,N_24941,N_24830);
or UO_331 (O_331,N_24329,N_24555);
nor UO_332 (O_332,N_24839,N_24950);
xnor UO_333 (O_333,N_24123,N_24356);
xor UO_334 (O_334,N_24194,N_24429);
nor UO_335 (O_335,N_24633,N_24192);
or UO_336 (O_336,N_24533,N_24691);
nand UO_337 (O_337,N_24886,N_24994);
and UO_338 (O_338,N_24476,N_24726);
and UO_339 (O_339,N_24281,N_24468);
nand UO_340 (O_340,N_24987,N_24933);
or UO_341 (O_341,N_24294,N_24339);
nor UO_342 (O_342,N_24983,N_24874);
nor UO_343 (O_343,N_24002,N_24075);
or UO_344 (O_344,N_24544,N_24999);
xor UO_345 (O_345,N_24015,N_24421);
nor UO_346 (O_346,N_24784,N_24084);
nor UO_347 (O_347,N_24143,N_24637);
xnor UO_348 (O_348,N_24447,N_24720);
and UO_349 (O_349,N_24416,N_24901);
and UO_350 (O_350,N_24956,N_24759);
nor UO_351 (O_351,N_24363,N_24112);
or UO_352 (O_352,N_24197,N_24526);
and UO_353 (O_353,N_24448,N_24059);
nor UO_354 (O_354,N_24572,N_24074);
nor UO_355 (O_355,N_24223,N_24998);
nor UO_356 (O_356,N_24921,N_24562);
xnor UO_357 (O_357,N_24295,N_24324);
nor UO_358 (O_358,N_24121,N_24896);
nor UO_359 (O_359,N_24849,N_24621);
nor UO_360 (O_360,N_24067,N_24393);
xor UO_361 (O_361,N_24580,N_24242);
and UO_362 (O_362,N_24414,N_24149);
or UO_363 (O_363,N_24077,N_24030);
nand UO_364 (O_364,N_24302,N_24326);
or UO_365 (O_365,N_24224,N_24190);
and UO_366 (O_366,N_24735,N_24390);
xor UO_367 (O_367,N_24328,N_24259);
or UO_368 (O_368,N_24788,N_24107);
nor UO_369 (O_369,N_24473,N_24225);
nor UO_370 (O_370,N_24008,N_24431);
xnor UO_371 (O_371,N_24187,N_24129);
nand UO_372 (O_372,N_24055,N_24045);
nor UO_373 (O_373,N_24869,N_24991);
nor UO_374 (O_374,N_24092,N_24932);
xnor UO_375 (O_375,N_24659,N_24483);
nand UO_376 (O_376,N_24379,N_24641);
or UO_377 (O_377,N_24408,N_24418);
and UO_378 (O_378,N_24369,N_24523);
xnor UO_379 (O_379,N_24023,N_24177);
and UO_380 (O_380,N_24693,N_24740);
or UO_381 (O_381,N_24524,N_24219);
and UO_382 (O_382,N_24719,N_24973);
and UO_383 (O_383,N_24644,N_24378);
nand UO_384 (O_384,N_24464,N_24042);
nand UO_385 (O_385,N_24367,N_24465);
nand UO_386 (O_386,N_24510,N_24354);
nand UO_387 (O_387,N_24539,N_24175);
xnor UO_388 (O_388,N_24140,N_24432);
nand UO_389 (O_389,N_24729,N_24309);
xnor UO_390 (O_390,N_24657,N_24574);
or UO_391 (O_391,N_24556,N_24721);
or UO_392 (O_392,N_24377,N_24040);
nor UO_393 (O_393,N_24952,N_24215);
or UO_394 (O_394,N_24446,N_24463);
nand UO_395 (O_395,N_24137,N_24376);
and UO_396 (O_396,N_24155,N_24807);
nor UO_397 (O_397,N_24550,N_24487);
nand UO_398 (O_398,N_24774,N_24507);
and UO_399 (O_399,N_24832,N_24395);
and UO_400 (O_400,N_24594,N_24511);
nor UO_401 (O_401,N_24094,N_24588);
xor UO_402 (O_402,N_24238,N_24538);
nor UO_403 (O_403,N_24992,N_24543);
or UO_404 (O_404,N_24619,N_24387);
xnor UO_405 (O_405,N_24185,N_24052);
or UO_406 (O_406,N_24792,N_24202);
and UO_407 (O_407,N_24806,N_24435);
or UO_408 (O_408,N_24024,N_24586);
nor UO_409 (O_409,N_24360,N_24180);
nor UO_410 (O_410,N_24206,N_24461);
nand UO_411 (O_411,N_24783,N_24805);
nor UO_412 (O_412,N_24425,N_24718);
nor UO_413 (O_413,N_24337,N_24388);
xnor UO_414 (O_414,N_24422,N_24626);
nor UO_415 (O_415,N_24624,N_24167);
xnor UO_416 (O_416,N_24437,N_24087);
xnor UO_417 (O_417,N_24359,N_24879);
and UO_418 (O_418,N_24643,N_24964);
nand UO_419 (O_419,N_24848,N_24755);
nor UO_420 (O_420,N_24982,N_24866);
or UO_421 (O_421,N_24263,N_24863);
nor UO_422 (O_422,N_24545,N_24423);
xor UO_423 (O_423,N_24278,N_24971);
or UO_424 (O_424,N_24480,N_24409);
and UO_425 (O_425,N_24882,N_24311);
or UO_426 (O_426,N_24802,N_24675);
nor UO_427 (O_427,N_24739,N_24661);
or UO_428 (O_428,N_24298,N_24648);
nand UO_429 (O_429,N_24965,N_24756);
and UO_430 (O_430,N_24355,N_24930);
or UO_431 (O_431,N_24702,N_24391);
nand UO_432 (O_432,N_24529,N_24230);
and UO_433 (O_433,N_24542,N_24716);
nor UO_434 (O_434,N_24795,N_24198);
or UO_435 (O_435,N_24256,N_24445);
xor UO_436 (O_436,N_24304,N_24020);
nor UO_437 (O_437,N_24474,N_24282);
or UO_438 (O_438,N_24909,N_24760);
xnor UO_439 (O_439,N_24953,N_24315);
nor UO_440 (O_440,N_24978,N_24156);
and UO_441 (O_441,N_24837,N_24651);
nand UO_442 (O_442,N_24672,N_24817);
and UO_443 (O_443,N_24380,N_24250);
or UO_444 (O_444,N_24183,N_24400);
nand UO_445 (O_445,N_24931,N_24170);
nor UO_446 (O_446,N_24280,N_24531);
xor UO_447 (O_447,N_24076,N_24868);
or UO_448 (O_448,N_24178,N_24861);
nor UO_449 (O_449,N_24475,N_24614);
nand UO_450 (O_450,N_24289,N_24272);
nand UO_451 (O_451,N_24546,N_24063);
nor UO_452 (O_452,N_24506,N_24599);
nor UO_453 (O_453,N_24785,N_24762);
nor UO_454 (O_454,N_24443,N_24876);
and UO_455 (O_455,N_24504,N_24678);
nand UO_456 (O_456,N_24006,N_24240);
nor UO_457 (O_457,N_24196,N_24703);
nor UO_458 (O_458,N_24104,N_24290);
nor UO_459 (O_459,N_24217,N_24307);
nand UO_460 (O_460,N_24433,N_24568);
xnor UO_461 (O_461,N_24327,N_24338);
or UO_462 (O_462,N_24717,N_24134);
xor UO_463 (O_463,N_24036,N_24460);
and UO_464 (O_464,N_24173,N_24427);
nand UO_465 (O_465,N_24842,N_24113);
nor UO_466 (O_466,N_24254,N_24469);
nor UO_467 (O_467,N_24001,N_24710);
nand UO_468 (O_468,N_24853,N_24585);
nand UO_469 (O_469,N_24725,N_24843);
or UO_470 (O_470,N_24974,N_24532);
or UO_471 (O_471,N_24692,N_24743);
nand UO_472 (O_472,N_24306,N_24300);
or UO_473 (O_473,N_24383,N_24885);
nand UO_474 (O_474,N_24385,N_24708);
nand UO_475 (O_475,N_24286,N_24120);
xnor UO_476 (O_476,N_24265,N_24613);
xnor UO_477 (O_477,N_24078,N_24284);
xnor UO_478 (O_478,N_24135,N_24430);
nor UO_479 (O_479,N_24856,N_24039);
and UO_480 (O_480,N_24900,N_24117);
and UO_481 (O_481,N_24627,N_24996);
nand UO_482 (O_482,N_24631,N_24305);
nor UO_483 (O_483,N_24875,N_24905);
and UO_484 (O_484,N_24371,N_24489);
or UO_485 (O_485,N_24898,N_24560);
xor UO_486 (O_486,N_24663,N_24803);
or UO_487 (O_487,N_24441,N_24899);
or UO_488 (O_488,N_24677,N_24207);
or UO_489 (O_489,N_24345,N_24191);
nor UO_490 (O_490,N_24668,N_24062);
and UO_491 (O_491,N_24810,N_24182);
nor UO_492 (O_492,N_24833,N_24647);
nand UO_493 (O_493,N_24728,N_24220);
or UO_494 (O_494,N_24765,N_24835);
nor UO_495 (O_495,N_24257,N_24741);
and UO_496 (O_496,N_24136,N_24970);
and UO_497 (O_497,N_24470,N_24912);
and UO_498 (O_498,N_24319,N_24091);
or UO_499 (O_499,N_24910,N_24664);
nand UO_500 (O_500,N_24241,N_24480);
nor UO_501 (O_501,N_24380,N_24727);
xor UO_502 (O_502,N_24543,N_24370);
xor UO_503 (O_503,N_24196,N_24700);
and UO_504 (O_504,N_24254,N_24219);
nor UO_505 (O_505,N_24052,N_24044);
nor UO_506 (O_506,N_24244,N_24437);
nand UO_507 (O_507,N_24720,N_24138);
xor UO_508 (O_508,N_24454,N_24050);
xnor UO_509 (O_509,N_24968,N_24810);
or UO_510 (O_510,N_24973,N_24801);
nor UO_511 (O_511,N_24959,N_24303);
nor UO_512 (O_512,N_24807,N_24343);
xor UO_513 (O_513,N_24611,N_24493);
xor UO_514 (O_514,N_24351,N_24282);
xnor UO_515 (O_515,N_24201,N_24918);
nor UO_516 (O_516,N_24197,N_24439);
or UO_517 (O_517,N_24382,N_24717);
xor UO_518 (O_518,N_24597,N_24527);
or UO_519 (O_519,N_24082,N_24652);
xnor UO_520 (O_520,N_24232,N_24035);
xor UO_521 (O_521,N_24841,N_24701);
nand UO_522 (O_522,N_24593,N_24730);
and UO_523 (O_523,N_24686,N_24591);
or UO_524 (O_524,N_24785,N_24433);
nand UO_525 (O_525,N_24892,N_24355);
nor UO_526 (O_526,N_24636,N_24932);
nor UO_527 (O_527,N_24458,N_24209);
xor UO_528 (O_528,N_24015,N_24848);
or UO_529 (O_529,N_24059,N_24510);
or UO_530 (O_530,N_24536,N_24750);
nand UO_531 (O_531,N_24086,N_24753);
or UO_532 (O_532,N_24804,N_24127);
xor UO_533 (O_533,N_24239,N_24505);
and UO_534 (O_534,N_24706,N_24271);
or UO_535 (O_535,N_24153,N_24771);
and UO_536 (O_536,N_24695,N_24564);
nor UO_537 (O_537,N_24415,N_24201);
or UO_538 (O_538,N_24371,N_24234);
nand UO_539 (O_539,N_24611,N_24303);
or UO_540 (O_540,N_24587,N_24071);
and UO_541 (O_541,N_24908,N_24716);
and UO_542 (O_542,N_24803,N_24033);
nand UO_543 (O_543,N_24082,N_24767);
and UO_544 (O_544,N_24321,N_24926);
nand UO_545 (O_545,N_24158,N_24555);
xnor UO_546 (O_546,N_24774,N_24375);
nor UO_547 (O_547,N_24560,N_24267);
xnor UO_548 (O_548,N_24156,N_24953);
and UO_549 (O_549,N_24988,N_24460);
nand UO_550 (O_550,N_24017,N_24395);
nor UO_551 (O_551,N_24287,N_24603);
nand UO_552 (O_552,N_24083,N_24102);
xor UO_553 (O_553,N_24761,N_24142);
nand UO_554 (O_554,N_24607,N_24116);
nand UO_555 (O_555,N_24747,N_24767);
nand UO_556 (O_556,N_24762,N_24478);
nand UO_557 (O_557,N_24367,N_24146);
nor UO_558 (O_558,N_24565,N_24662);
xnor UO_559 (O_559,N_24913,N_24566);
or UO_560 (O_560,N_24337,N_24561);
nor UO_561 (O_561,N_24594,N_24053);
and UO_562 (O_562,N_24897,N_24876);
nand UO_563 (O_563,N_24571,N_24165);
and UO_564 (O_564,N_24053,N_24152);
or UO_565 (O_565,N_24060,N_24848);
or UO_566 (O_566,N_24065,N_24235);
nand UO_567 (O_567,N_24836,N_24827);
xnor UO_568 (O_568,N_24299,N_24821);
or UO_569 (O_569,N_24004,N_24510);
or UO_570 (O_570,N_24029,N_24206);
or UO_571 (O_571,N_24133,N_24077);
nor UO_572 (O_572,N_24854,N_24558);
and UO_573 (O_573,N_24137,N_24289);
xnor UO_574 (O_574,N_24359,N_24161);
nand UO_575 (O_575,N_24660,N_24955);
and UO_576 (O_576,N_24813,N_24770);
nor UO_577 (O_577,N_24902,N_24386);
nand UO_578 (O_578,N_24504,N_24390);
and UO_579 (O_579,N_24114,N_24578);
xor UO_580 (O_580,N_24090,N_24919);
nor UO_581 (O_581,N_24953,N_24641);
nor UO_582 (O_582,N_24394,N_24048);
xnor UO_583 (O_583,N_24582,N_24950);
and UO_584 (O_584,N_24393,N_24983);
and UO_585 (O_585,N_24220,N_24405);
and UO_586 (O_586,N_24361,N_24880);
nand UO_587 (O_587,N_24339,N_24675);
or UO_588 (O_588,N_24050,N_24064);
xnor UO_589 (O_589,N_24396,N_24391);
and UO_590 (O_590,N_24931,N_24658);
nand UO_591 (O_591,N_24746,N_24070);
xnor UO_592 (O_592,N_24332,N_24963);
nor UO_593 (O_593,N_24585,N_24126);
and UO_594 (O_594,N_24024,N_24949);
nor UO_595 (O_595,N_24472,N_24667);
nor UO_596 (O_596,N_24380,N_24513);
and UO_597 (O_597,N_24933,N_24504);
or UO_598 (O_598,N_24596,N_24487);
nand UO_599 (O_599,N_24095,N_24600);
or UO_600 (O_600,N_24671,N_24371);
nor UO_601 (O_601,N_24007,N_24226);
nand UO_602 (O_602,N_24140,N_24521);
nand UO_603 (O_603,N_24983,N_24859);
and UO_604 (O_604,N_24774,N_24455);
or UO_605 (O_605,N_24271,N_24854);
nand UO_606 (O_606,N_24295,N_24518);
nand UO_607 (O_607,N_24924,N_24294);
and UO_608 (O_608,N_24706,N_24164);
or UO_609 (O_609,N_24878,N_24458);
nor UO_610 (O_610,N_24687,N_24556);
or UO_611 (O_611,N_24993,N_24592);
or UO_612 (O_612,N_24378,N_24980);
xnor UO_613 (O_613,N_24309,N_24261);
nand UO_614 (O_614,N_24048,N_24796);
and UO_615 (O_615,N_24594,N_24020);
nand UO_616 (O_616,N_24798,N_24027);
or UO_617 (O_617,N_24974,N_24990);
xor UO_618 (O_618,N_24000,N_24520);
nor UO_619 (O_619,N_24875,N_24756);
and UO_620 (O_620,N_24532,N_24838);
nand UO_621 (O_621,N_24984,N_24480);
nor UO_622 (O_622,N_24945,N_24343);
xor UO_623 (O_623,N_24167,N_24646);
or UO_624 (O_624,N_24220,N_24342);
xnor UO_625 (O_625,N_24684,N_24522);
or UO_626 (O_626,N_24961,N_24868);
xnor UO_627 (O_627,N_24751,N_24499);
or UO_628 (O_628,N_24457,N_24964);
and UO_629 (O_629,N_24107,N_24553);
xor UO_630 (O_630,N_24463,N_24933);
nor UO_631 (O_631,N_24993,N_24187);
xor UO_632 (O_632,N_24639,N_24479);
xor UO_633 (O_633,N_24107,N_24137);
or UO_634 (O_634,N_24335,N_24024);
and UO_635 (O_635,N_24799,N_24989);
and UO_636 (O_636,N_24211,N_24119);
or UO_637 (O_637,N_24961,N_24164);
and UO_638 (O_638,N_24383,N_24911);
and UO_639 (O_639,N_24988,N_24372);
nand UO_640 (O_640,N_24298,N_24931);
or UO_641 (O_641,N_24812,N_24971);
nor UO_642 (O_642,N_24533,N_24101);
nand UO_643 (O_643,N_24231,N_24932);
xnor UO_644 (O_644,N_24109,N_24755);
xnor UO_645 (O_645,N_24216,N_24672);
or UO_646 (O_646,N_24206,N_24421);
nand UO_647 (O_647,N_24960,N_24050);
or UO_648 (O_648,N_24999,N_24985);
or UO_649 (O_649,N_24359,N_24933);
nor UO_650 (O_650,N_24004,N_24469);
or UO_651 (O_651,N_24734,N_24946);
or UO_652 (O_652,N_24856,N_24102);
xor UO_653 (O_653,N_24307,N_24403);
and UO_654 (O_654,N_24111,N_24455);
nor UO_655 (O_655,N_24054,N_24676);
or UO_656 (O_656,N_24128,N_24374);
and UO_657 (O_657,N_24136,N_24816);
xnor UO_658 (O_658,N_24028,N_24181);
nand UO_659 (O_659,N_24594,N_24750);
nor UO_660 (O_660,N_24952,N_24856);
nor UO_661 (O_661,N_24468,N_24148);
and UO_662 (O_662,N_24177,N_24545);
nand UO_663 (O_663,N_24862,N_24531);
nor UO_664 (O_664,N_24815,N_24604);
xor UO_665 (O_665,N_24122,N_24808);
xnor UO_666 (O_666,N_24833,N_24038);
nor UO_667 (O_667,N_24750,N_24277);
nand UO_668 (O_668,N_24927,N_24717);
xor UO_669 (O_669,N_24451,N_24351);
and UO_670 (O_670,N_24706,N_24212);
and UO_671 (O_671,N_24908,N_24408);
xor UO_672 (O_672,N_24455,N_24105);
nor UO_673 (O_673,N_24246,N_24024);
or UO_674 (O_674,N_24674,N_24938);
nand UO_675 (O_675,N_24852,N_24678);
or UO_676 (O_676,N_24199,N_24290);
nand UO_677 (O_677,N_24343,N_24197);
and UO_678 (O_678,N_24292,N_24124);
xnor UO_679 (O_679,N_24147,N_24985);
nand UO_680 (O_680,N_24470,N_24940);
or UO_681 (O_681,N_24243,N_24208);
and UO_682 (O_682,N_24496,N_24116);
or UO_683 (O_683,N_24556,N_24366);
or UO_684 (O_684,N_24769,N_24408);
nor UO_685 (O_685,N_24157,N_24387);
xor UO_686 (O_686,N_24811,N_24259);
and UO_687 (O_687,N_24168,N_24104);
nor UO_688 (O_688,N_24480,N_24955);
xnor UO_689 (O_689,N_24326,N_24709);
or UO_690 (O_690,N_24197,N_24732);
and UO_691 (O_691,N_24358,N_24031);
and UO_692 (O_692,N_24768,N_24715);
and UO_693 (O_693,N_24712,N_24274);
or UO_694 (O_694,N_24777,N_24251);
and UO_695 (O_695,N_24087,N_24458);
and UO_696 (O_696,N_24917,N_24029);
nand UO_697 (O_697,N_24953,N_24884);
nand UO_698 (O_698,N_24336,N_24041);
and UO_699 (O_699,N_24618,N_24664);
nor UO_700 (O_700,N_24554,N_24408);
and UO_701 (O_701,N_24287,N_24516);
xnor UO_702 (O_702,N_24746,N_24157);
nor UO_703 (O_703,N_24815,N_24829);
xnor UO_704 (O_704,N_24978,N_24212);
xnor UO_705 (O_705,N_24025,N_24664);
nand UO_706 (O_706,N_24925,N_24226);
xor UO_707 (O_707,N_24110,N_24819);
xor UO_708 (O_708,N_24354,N_24390);
nand UO_709 (O_709,N_24776,N_24144);
and UO_710 (O_710,N_24697,N_24578);
xor UO_711 (O_711,N_24930,N_24868);
xnor UO_712 (O_712,N_24922,N_24213);
and UO_713 (O_713,N_24557,N_24147);
nand UO_714 (O_714,N_24183,N_24303);
xnor UO_715 (O_715,N_24603,N_24884);
or UO_716 (O_716,N_24298,N_24437);
nand UO_717 (O_717,N_24095,N_24233);
nor UO_718 (O_718,N_24932,N_24326);
and UO_719 (O_719,N_24561,N_24822);
and UO_720 (O_720,N_24840,N_24617);
or UO_721 (O_721,N_24468,N_24055);
and UO_722 (O_722,N_24372,N_24164);
and UO_723 (O_723,N_24478,N_24243);
xnor UO_724 (O_724,N_24026,N_24954);
nand UO_725 (O_725,N_24464,N_24545);
or UO_726 (O_726,N_24406,N_24871);
or UO_727 (O_727,N_24573,N_24520);
xor UO_728 (O_728,N_24733,N_24324);
nand UO_729 (O_729,N_24986,N_24760);
or UO_730 (O_730,N_24198,N_24678);
nand UO_731 (O_731,N_24539,N_24183);
nor UO_732 (O_732,N_24118,N_24543);
or UO_733 (O_733,N_24127,N_24071);
nor UO_734 (O_734,N_24134,N_24642);
xor UO_735 (O_735,N_24448,N_24333);
nand UO_736 (O_736,N_24135,N_24296);
nor UO_737 (O_737,N_24505,N_24620);
xnor UO_738 (O_738,N_24684,N_24636);
nor UO_739 (O_739,N_24170,N_24229);
nand UO_740 (O_740,N_24831,N_24298);
xnor UO_741 (O_741,N_24596,N_24523);
xnor UO_742 (O_742,N_24779,N_24927);
xnor UO_743 (O_743,N_24631,N_24257);
or UO_744 (O_744,N_24760,N_24375);
and UO_745 (O_745,N_24622,N_24335);
and UO_746 (O_746,N_24123,N_24331);
or UO_747 (O_747,N_24088,N_24147);
nor UO_748 (O_748,N_24468,N_24470);
nand UO_749 (O_749,N_24323,N_24860);
nor UO_750 (O_750,N_24398,N_24901);
nor UO_751 (O_751,N_24132,N_24522);
nor UO_752 (O_752,N_24159,N_24092);
and UO_753 (O_753,N_24797,N_24271);
xnor UO_754 (O_754,N_24035,N_24460);
nand UO_755 (O_755,N_24619,N_24599);
nand UO_756 (O_756,N_24108,N_24475);
nand UO_757 (O_757,N_24289,N_24325);
and UO_758 (O_758,N_24854,N_24676);
nand UO_759 (O_759,N_24058,N_24037);
nor UO_760 (O_760,N_24988,N_24355);
nand UO_761 (O_761,N_24542,N_24934);
xor UO_762 (O_762,N_24596,N_24425);
nand UO_763 (O_763,N_24515,N_24829);
xor UO_764 (O_764,N_24450,N_24500);
nand UO_765 (O_765,N_24672,N_24785);
xor UO_766 (O_766,N_24962,N_24920);
and UO_767 (O_767,N_24262,N_24966);
or UO_768 (O_768,N_24249,N_24900);
xnor UO_769 (O_769,N_24432,N_24113);
xnor UO_770 (O_770,N_24492,N_24434);
xnor UO_771 (O_771,N_24438,N_24240);
xor UO_772 (O_772,N_24185,N_24098);
nor UO_773 (O_773,N_24385,N_24002);
nor UO_774 (O_774,N_24093,N_24399);
or UO_775 (O_775,N_24555,N_24060);
xor UO_776 (O_776,N_24210,N_24482);
nor UO_777 (O_777,N_24938,N_24350);
or UO_778 (O_778,N_24535,N_24763);
nand UO_779 (O_779,N_24980,N_24222);
or UO_780 (O_780,N_24042,N_24815);
nor UO_781 (O_781,N_24062,N_24565);
nor UO_782 (O_782,N_24337,N_24830);
xnor UO_783 (O_783,N_24649,N_24955);
xor UO_784 (O_784,N_24755,N_24918);
and UO_785 (O_785,N_24630,N_24433);
or UO_786 (O_786,N_24728,N_24797);
nand UO_787 (O_787,N_24431,N_24361);
xnor UO_788 (O_788,N_24817,N_24646);
and UO_789 (O_789,N_24479,N_24921);
and UO_790 (O_790,N_24437,N_24477);
nor UO_791 (O_791,N_24114,N_24935);
xnor UO_792 (O_792,N_24035,N_24435);
nor UO_793 (O_793,N_24405,N_24496);
xor UO_794 (O_794,N_24521,N_24736);
nor UO_795 (O_795,N_24793,N_24381);
nand UO_796 (O_796,N_24234,N_24167);
and UO_797 (O_797,N_24834,N_24269);
nand UO_798 (O_798,N_24522,N_24577);
xor UO_799 (O_799,N_24993,N_24148);
or UO_800 (O_800,N_24292,N_24557);
xnor UO_801 (O_801,N_24794,N_24996);
nor UO_802 (O_802,N_24974,N_24635);
nand UO_803 (O_803,N_24740,N_24033);
xnor UO_804 (O_804,N_24087,N_24834);
nor UO_805 (O_805,N_24463,N_24795);
xor UO_806 (O_806,N_24973,N_24198);
xnor UO_807 (O_807,N_24926,N_24695);
nand UO_808 (O_808,N_24145,N_24484);
nor UO_809 (O_809,N_24832,N_24207);
xor UO_810 (O_810,N_24202,N_24847);
xnor UO_811 (O_811,N_24404,N_24638);
nand UO_812 (O_812,N_24220,N_24754);
nor UO_813 (O_813,N_24450,N_24378);
xnor UO_814 (O_814,N_24468,N_24636);
and UO_815 (O_815,N_24873,N_24228);
and UO_816 (O_816,N_24012,N_24190);
and UO_817 (O_817,N_24938,N_24328);
nand UO_818 (O_818,N_24881,N_24213);
or UO_819 (O_819,N_24624,N_24094);
and UO_820 (O_820,N_24764,N_24225);
xor UO_821 (O_821,N_24476,N_24371);
and UO_822 (O_822,N_24952,N_24554);
nand UO_823 (O_823,N_24403,N_24933);
nor UO_824 (O_824,N_24649,N_24676);
xor UO_825 (O_825,N_24415,N_24656);
and UO_826 (O_826,N_24288,N_24048);
nor UO_827 (O_827,N_24355,N_24557);
nor UO_828 (O_828,N_24841,N_24263);
or UO_829 (O_829,N_24735,N_24486);
and UO_830 (O_830,N_24130,N_24016);
nand UO_831 (O_831,N_24244,N_24334);
or UO_832 (O_832,N_24604,N_24899);
and UO_833 (O_833,N_24188,N_24816);
nand UO_834 (O_834,N_24414,N_24692);
xnor UO_835 (O_835,N_24031,N_24548);
and UO_836 (O_836,N_24595,N_24107);
nor UO_837 (O_837,N_24002,N_24277);
and UO_838 (O_838,N_24545,N_24695);
or UO_839 (O_839,N_24571,N_24534);
or UO_840 (O_840,N_24988,N_24528);
nand UO_841 (O_841,N_24876,N_24874);
and UO_842 (O_842,N_24063,N_24118);
nor UO_843 (O_843,N_24303,N_24828);
nor UO_844 (O_844,N_24412,N_24371);
and UO_845 (O_845,N_24327,N_24927);
and UO_846 (O_846,N_24490,N_24933);
and UO_847 (O_847,N_24811,N_24863);
or UO_848 (O_848,N_24944,N_24834);
and UO_849 (O_849,N_24758,N_24581);
nand UO_850 (O_850,N_24234,N_24687);
xnor UO_851 (O_851,N_24106,N_24699);
xnor UO_852 (O_852,N_24784,N_24286);
or UO_853 (O_853,N_24248,N_24541);
and UO_854 (O_854,N_24483,N_24536);
and UO_855 (O_855,N_24704,N_24556);
nor UO_856 (O_856,N_24882,N_24336);
xor UO_857 (O_857,N_24364,N_24768);
xor UO_858 (O_858,N_24252,N_24963);
and UO_859 (O_859,N_24409,N_24672);
nand UO_860 (O_860,N_24164,N_24538);
or UO_861 (O_861,N_24728,N_24822);
nand UO_862 (O_862,N_24998,N_24295);
nor UO_863 (O_863,N_24362,N_24938);
nand UO_864 (O_864,N_24618,N_24727);
and UO_865 (O_865,N_24176,N_24000);
xnor UO_866 (O_866,N_24709,N_24562);
and UO_867 (O_867,N_24645,N_24891);
nand UO_868 (O_868,N_24724,N_24033);
xnor UO_869 (O_869,N_24663,N_24677);
nor UO_870 (O_870,N_24928,N_24145);
nand UO_871 (O_871,N_24503,N_24127);
and UO_872 (O_872,N_24291,N_24036);
and UO_873 (O_873,N_24250,N_24309);
nand UO_874 (O_874,N_24822,N_24798);
and UO_875 (O_875,N_24772,N_24866);
and UO_876 (O_876,N_24302,N_24197);
xor UO_877 (O_877,N_24278,N_24915);
xnor UO_878 (O_878,N_24501,N_24082);
nor UO_879 (O_879,N_24891,N_24527);
and UO_880 (O_880,N_24627,N_24249);
and UO_881 (O_881,N_24672,N_24797);
nand UO_882 (O_882,N_24136,N_24112);
nand UO_883 (O_883,N_24799,N_24418);
and UO_884 (O_884,N_24593,N_24744);
or UO_885 (O_885,N_24504,N_24461);
or UO_886 (O_886,N_24999,N_24680);
nand UO_887 (O_887,N_24019,N_24794);
nor UO_888 (O_888,N_24001,N_24017);
and UO_889 (O_889,N_24864,N_24133);
xor UO_890 (O_890,N_24655,N_24952);
nor UO_891 (O_891,N_24081,N_24604);
xnor UO_892 (O_892,N_24006,N_24205);
and UO_893 (O_893,N_24985,N_24699);
and UO_894 (O_894,N_24076,N_24399);
or UO_895 (O_895,N_24217,N_24477);
or UO_896 (O_896,N_24625,N_24578);
nor UO_897 (O_897,N_24328,N_24601);
nand UO_898 (O_898,N_24151,N_24898);
nor UO_899 (O_899,N_24494,N_24020);
or UO_900 (O_900,N_24331,N_24959);
nand UO_901 (O_901,N_24998,N_24373);
nor UO_902 (O_902,N_24849,N_24664);
or UO_903 (O_903,N_24000,N_24086);
and UO_904 (O_904,N_24995,N_24005);
xor UO_905 (O_905,N_24340,N_24064);
xnor UO_906 (O_906,N_24358,N_24649);
xor UO_907 (O_907,N_24720,N_24702);
nor UO_908 (O_908,N_24070,N_24606);
and UO_909 (O_909,N_24632,N_24615);
or UO_910 (O_910,N_24359,N_24325);
xnor UO_911 (O_911,N_24889,N_24944);
nand UO_912 (O_912,N_24702,N_24876);
nor UO_913 (O_913,N_24692,N_24735);
and UO_914 (O_914,N_24641,N_24593);
nor UO_915 (O_915,N_24349,N_24529);
or UO_916 (O_916,N_24682,N_24914);
xnor UO_917 (O_917,N_24504,N_24748);
nand UO_918 (O_918,N_24035,N_24701);
or UO_919 (O_919,N_24971,N_24221);
xor UO_920 (O_920,N_24085,N_24820);
nand UO_921 (O_921,N_24882,N_24557);
or UO_922 (O_922,N_24636,N_24966);
xor UO_923 (O_923,N_24837,N_24340);
nand UO_924 (O_924,N_24180,N_24599);
and UO_925 (O_925,N_24720,N_24766);
nor UO_926 (O_926,N_24011,N_24599);
xnor UO_927 (O_927,N_24393,N_24113);
and UO_928 (O_928,N_24042,N_24296);
nand UO_929 (O_929,N_24549,N_24666);
nor UO_930 (O_930,N_24029,N_24447);
nand UO_931 (O_931,N_24046,N_24934);
xnor UO_932 (O_932,N_24561,N_24944);
and UO_933 (O_933,N_24349,N_24662);
nor UO_934 (O_934,N_24008,N_24690);
nand UO_935 (O_935,N_24974,N_24551);
or UO_936 (O_936,N_24622,N_24883);
xor UO_937 (O_937,N_24666,N_24828);
nor UO_938 (O_938,N_24429,N_24410);
xor UO_939 (O_939,N_24256,N_24423);
and UO_940 (O_940,N_24376,N_24348);
and UO_941 (O_941,N_24296,N_24532);
or UO_942 (O_942,N_24441,N_24343);
or UO_943 (O_943,N_24024,N_24589);
and UO_944 (O_944,N_24885,N_24339);
nor UO_945 (O_945,N_24104,N_24436);
nor UO_946 (O_946,N_24869,N_24864);
and UO_947 (O_947,N_24877,N_24217);
xnor UO_948 (O_948,N_24363,N_24454);
nor UO_949 (O_949,N_24692,N_24589);
xnor UO_950 (O_950,N_24097,N_24125);
and UO_951 (O_951,N_24560,N_24687);
nor UO_952 (O_952,N_24495,N_24651);
nand UO_953 (O_953,N_24064,N_24266);
and UO_954 (O_954,N_24584,N_24681);
and UO_955 (O_955,N_24240,N_24544);
or UO_956 (O_956,N_24698,N_24522);
xor UO_957 (O_957,N_24772,N_24286);
or UO_958 (O_958,N_24456,N_24383);
and UO_959 (O_959,N_24935,N_24106);
nor UO_960 (O_960,N_24790,N_24556);
or UO_961 (O_961,N_24027,N_24934);
nand UO_962 (O_962,N_24934,N_24904);
nor UO_963 (O_963,N_24724,N_24140);
nand UO_964 (O_964,N_24469,N_24050);
nor UO_965 (O_965,N_24957,N_24728);
or UO_966 (O_966,N_24339,N_24352);
nand UO_967 (O_967,N_24075,N_24228);
and UO_968 (O_968,N_24593,N_24857);
or UO_969 (O_969,N_24801,N_24830);
and UO_970 (O_970,N_24366,N_24112);
nand UO_971 (O_971,N_24403,N_24073);
and UO_972 (O_972,N_24662,N_24055);
xor UO_973 (O_973,N_24691,N_24267);
nand UO_974 (O_974,N_24592,N_24225);
xnor UO_975 (O_975,N_24779,N_24652);
or UO_976 (O_976,N_24762,N_24034);
and UO_977 (O_977,N_24563,N_24269);
nor UO_978 (O_978,N_24227,N_24450);
or UO_979 (O_979,N_24612,N_24934);
xnor UO_980 (O_980,N_24627,N_24323);
nand UO_981 (O_981,N_24103,N_24713);
xnor UO_982 (O_982,N_24944,N_24958);
and UO_983 (O_983,N_24883,N_24491);
or UO_984 (O_984,N_24215,N_24341);
or UO_985 (O_985,N_24828,N_24595);
nor UO_986 (O_986,N_24333,N_24485);
xor UO_987 (O_987,N_24880,N_24109);
nand UO_988 (O_988,N_24253,N_24164);
and UO_989 (O_989,N_24602,N_24509);
nand UO_990 (O_990,N_24369,N_24822);
or UO_991 (O_991,N_24623,N_24074);
xor UO_992 (O_992,N_24711,N_24798);
or UO_993 (O_993,N_24211,N_24547);
xor UO_994 (O_994,N_24274,N_24040);
or UO_995 (O_995,N_24844,N_24103);
nand UO_996 (O_996,N_24492,N_24897);
or UO_997 (O_997,N_24902,N_24724);
nor UO_998 (O_998,N_24226,N_24911);
nand UO_999 (O_999,N_24563,N_24089);
xnor UO_1000 (O_1000,N_24523,N_24461);
or UO_1001 (O_1001,N_24669,N_24928);
or UO_1002 (O_1002,N_24854,N_24362);
or UO_1003 (O_1003,N_24419,N_24682);
nand UO_1004 (O_1004,N_24002,N_24530);
xnor UO_1005 (O_1005,N_24141,N_24400);
nand UO_1006 (O_1006,N_24281,N_24330);
xor UO_1007 (O_1007,N_24646,N_24945);
nor UO_1008 (O_1008,N_24124,N_24153);
nor UO_1009 (O_1009,N_24966,N_24574);
or UO_1010 (O_1010,N_24172,N_24168);
nand UO_1011 (O_1011,N_24560,N_24699);
and UO_1012 (O_1012,N_24882,N_24424);
xnor UO_1013 (O_1013,N_24535,N_24826);
or UO_1014 (O_1014,N_24949,N_24732);
or UO_1015 (O_1015,N_24551,N_24253);
or UO_1016 (O_1016,N_24461,N_24979);
xnor UO_1017 (O_1017,N_24164,N_24689);
nand UO_1018 (O_1018,N_24926,N_24292);
xor UO_1019 (O_1019,N_24043,N_24803);
or UO_1020 (O_1020,N_24038,N_24333);
nor UO_1021 (O_1021,N_24480,N_24269);
nor UO_1022 (O_1022,N_24337,N_24748);
and UO_1023 (O_1023,N_24581,N_24989);
xnor UO_1024 (O_1024,N_24841,N_24231);
xor UO_1025 (O_1025,N_24097,N_24910);
nand UO_1026 (O_1026,N_24149,N_24447);
xnor UO_1027 (O_1027,N_24118,N_24301);
nor UO_1028 (O_1028,N_24352,N_24231);
and UO_1029 (O_1029,N_24894,N_24942);
and UO_1030 (O_1030,N_24620,N_24309);
and UO_1031 (O_1031,N_24557,N_24992);
nor UO_1032 (O_1032,N_24235,N_24227);
and UO_1033 (O_1033,N_24956,N_24197);
nand UO_1034 (O_1034,N_24586,N_24272);
nand UO_1035 (O_1035,N_24115,N_24699);
nand UO_1036 (O_1036,N_24170,N_24643);
and UO_1037 (O_1037,N_24529,N_24745);
and UO_1038 (O_1038,N_24048,N_24461);
xnor UO_1039 (O_1039,N_24457,N_24421);
or UO_1040 (O_1040,N_24701,N_24597);
or UO_1041 (O_1041,N_24963,N_24664);
xor UO_1042 (O_1042,N_24620,N_24094);
or UO_1043 (O_1043,N_24733,N_24542);
xor UO_1044 (O_1044,N_24432,N_24256);
and UO_1045 (O_1045,N_24446,N_24379);
xor UO_1046 (O_1046,N_24861,N_24209);
and UO_1047 (O_1047,N_24577,N_24856);
and UO_1048 (O_1048,N_24402,N_24181);
nor UO_1049 (O_1049,N_24008,N_24853);
xnor UO_1050 (O_1050,N_24998,N_24702);
and UO_1051 (O_1051,N_24516,N_24418);
nor UO_1052 (O_1052,N_24951,N_24268);
and UO_1053 (O_1053,N_24108,N_24441);
nand UO_1054 (O_1054,N_24632,N_24298);
and UO_1055 (O_1055,N_24789,N_24229);
and UO_1056 (O_1056,N_24466,N_24100);
xnor UO_1057 (O_1057,N_24086,N_24270);
or UO_1058 (O_1058,N_24522,N_24360);
and UO_1059 (O_1059,N_24363,N_24092);
or UO_1060 (O_1060,N_24031,N_24870);
xor UO_1061 (O_1061,N_24238,N_24534);
nand UO_1062 (O_1062,N_24163,N_24922);
nor UO_1063 (O_1063,N_24595,N_24148);
or UO_1064 (O_1064,N_24586,N_24799);
nor UO_1065 (O_1065,N_24959,N_24734);
and UO_1066 (O_1066,N_24699,N_24557);
nand UO_1067 (O_1067,N_24358,N_24408);
and UO_1068 (O_1068,N_24585,N_24777);
or UO_1069 (O_1069,N_24650,N_24698);
and UO_1070 (O_1070,N_24336,N_24447);
or UO_1071 (O_1071,N_24220,N_24881);
xnor UO_1072 (O_1072,N_24534,N_24857);
nand UO_1073 (O_1073,N_24896,N_24612);
nand UO_1074 (O_1074,N_24412,N_24544);
or UO_1075 (O_1075,N_24784,N_24869);
and UO_1076 (O_1076,N_24209,N_24130);
nor UO_1077 (O_1077,N_24494,N_24863);
xnor UO_1078 (O_1078,N_24506,N_24840);
nand UO_1079 (O_1079,N_24400,N_24356);
xnor UO_1080 (O_1080,N_24675,N_24732);
xor UO_1081 (O_1081,N_24958,N_24762);
or UO_1082 (O_1082,N_24539,N_24268);
nor UO_1083 (O_1083,N_24371,N_24646);
and UO_1084 (O_1084,N_24006,N_24152);
nor UO_1085 (O_1085,N_24111,N_24200);
or UO_1086 (O_1086,N_24355,N_24422);
or UO_1087 (O_1087,N_24795,N_24840);
or UO_1088 (O_1088,N_24308,N_24962);
nand UO_1089 (O_1089,N_24366,N_24871);
xor UO_1090 (O_1090,N_24948,N_24984);
nor UO_1091 (O_1091,N_24682,N_24868);
and UO_1092 (O_1092,N_24646,N_24470);
and UO_1093 (O_1093,N_24875,N_24715);
nor UO_1094 (O_1094,N_24489,N_24206);
and UO_1095 (O_1095,N_24992,N_24963);
xor UO_1096 (O_1096,N_24802,N_24940);
and UO_1097 (O_1097,N_24549,N_24608);
and UO_1098 (O_1098,N_24577,N_24058);
xnor UO_1099 (O_1099,N_24041,N_24547);
nor UO_1100 (O_1100,N_24978,N_24487);
or UO_1101 (O_1101,N_24898,N_24134);
nand UO_1102 (O_1102,N_24331,N_24521);
nand UO_1103 (O_1103,N_24906,N_24496);
nand UO_1104 (O_1104,N_24267,N_24967);
and UO_1105 (O_1105,N_24438,N_24276);
or UO_1106 (O_1106,N_24143,N_24384);
nor UO_1107 (O_1107,N_24593,N_24459);
nand UO_1108 (O_1108,N_24008,N_24597);
xnor UO_1109 (O_1109,N_24967,N_24618);
xor UO_1110 (O_1110,N_24889,N_24322);
and UO_1111 (O_1111,N_24719,N_24912);
nor UO_1112 (O_1112,N_24077,N_24756);
or UO_1113 (O_1113,N_24024,N_24596);
nand UO_1114 (O_1114,N_24476,N_24246);
and UO_1115 (O_1115,N_24821,N_24889);
and UO_1116 (O_1116,N_24376,N_24600);
nand UO_1117 (O_1117,N_24809,N_24710);
nand UO_1118 (O_1118,N_24505,N_24459);
or UO_1119 (O_1119,N_24048,N_24664);
nor UO_1120 (O_1120,N_24300,N_24304);
or UO_1121 (O_1121,N_24700,N_24399);
nand UO_1122 (O_1122,N_24881,N_24103);
or UO_1123 (O_1123,N_24008,N_24280);
xor UO_1124 (O_1124,N_24152,N_24871);
and UO_1125 (O_1125,N_24507,N_24148);
or UO_1126 (O_1126,N_24733,N_24860);
xnor UO_1127 (O_1127,N_24072,N_24296);
nor UO_1128 (O_1128,N_24344,N_24795);
xnor UO_1129 (O_1129,N_24740,N_24085);
nor UO_1130 (O_1130,N_24736,N_24629);
nand UO_1131 (O_1131,N_24992,N_24060);
nand UO_1132 (O_1132,N_24401,N_24289);
xor UO_1133 (O_1133,N_24889,N_24842);
and UO_1134 (O_1134,N_24868,N_24846);
or UO_1135 (O_1135,N_24086,N_24416);
nor UO_1136 (O_1136,N_24431,N_24948);
nor UO_1137 (O_1137,N_24907,N_24176);
nand UO_1138 (O_1138,N_24711,N_24763);
xnor UO_1139 (O_1139,N_24005,N_24277);
or UO_1140 (O_1140,N_24034,N_24390);
xor UO_1141 (O_1141,N_24640,N_24241);
nand UO_1142 (O_1142,N_24880,N_24794);
and UO_1143 (O_1143,N_24446,N_24047);
nor UO_1144 (O_1144,N_24969,N_24845);
or UO_1145 (O_1145,N_24892,N_24524);
and UO_1146 (O_1146,N_24641,N_24037);
nor UO_1147 (O_1147,N_24101,N_24740);
and UO_1148 (O_1148,N_24141,N_24672);
nand UO_1149 (O_1149,N_24318,N_24615);
nor UO_1150 (O_1150,N_24336,N_24754);
or UO_1151 (O_1151,N_24260,N_24275);
xor UO_1152 (O_1152,N_24568,N_24598);
nand UO_1153 (O_1153,N_24794,N_24249);
xnor UO_1154 (O_1154,N_24847,N_24734);
nor UO_1155 (O_1155,N_24507,N_24483);
and UO_1156 (O_1156,N_24228,N_24106);
xor UO_1157 (O_1157,N_24405,N_24383);
nor UO_1158 (O_1158,N_24642,N_24896);
xnor UO_1159 (O_1159,N_24915,N_24517);
and UO_1160 (O_1160,N_24457,N_24973);
or UO_1161 (O_1161,N_24458,N_24212);
or UO_1162 (O_1162,N_24191,N_24947);
nor UO_1163 (O_1163,N_24161,N_24225);
nand UO_1164 (O_1164,N_24290,N_24629);
nand UO_1165 (O_1165,N_24271,N_24700);
nor UO_1166 (O_1166,N_24200,N_24985);
xnor UO_1167 (O_1167,N_24331,N_24186);
xnor UO_1168 (O_1168,N_24390,N_24208);
and UO_1169 (O_1169,N_24954,N_24839);
xor UO_1170 (O_1170,N_24756,N_24603);
or UO_1171 (O_1171,N_24526,N_24579);
nand UO_1172 (O_1172,N_24308,N_24533);
and UO_1173 (O_1173,N_24233,N_24799);
nor UO_1174 (O_1174,N_24677,N_24812);
nor UO_1175 (O_1175,N_24583,N_24643);
xor UO_1176 (O_1176,N_24821,N_24274);
nand UO_1177 (O_1177,N_24571,N_24946);
or UO_1178 (O_1178,N_24124,N_24079);
and UO_1179 (O_1179,N_24236,N_24424);
nand UO_1180 (O_1180,N_24181,N_24780);
xnor UO_1181 (O_1181,N_24070,N_24286);
xor UO_1182 (O_1182,N_24996,N_24273);
or UO_1183 (O_1183,N_24841,N_24183);
nor UO_1184 (O_1184,N_24672,N_24037);
and UO_1185 (O_1185,N_24205,N_24445);
nor UO_1186 (O_1186,N_24865,N_24535);
xnor UO_1187 (O_1187,N_24447,N_24931);
or UO_1188 (O_1188,N_24384,N_24153);
nand UO_1189 (O_1189,N_24335,N_24267);
nor UO_1190 (O_1190,N_24600,N_24136);
or UO_1191 (O_1191,N_24657,N_24649);
or UO_1192 (O_1192,N_24870,N_24829);
nand UO_1193 (O_1193,N_24206,N_24524);
and UO_1194 (O_1194,N_24567,N_24867);
and UO_1195 (O_1195,N_24233,N_24947);
nor UO_1196 (O_1196,N_24516,N_24787);
and UO_1197 (O_1197,N_24303,N_24614);
and UO_1198 (O_1198,N_24205,N_24998);
nor UO_1199 (O_1199,N_24051,N_24177);
nand UO_1200 (O_1200,N_24405,N_24655);
and UO_1201 (O_1201,N_24388,N_24021);
nor UO_1202 (O_1202,N_24417,N_24758);
nor UO_1203 (O_1203,N_24188,N_24889);
and UO_1204 (O_1204,N_24224,N_24697);
and UO_1205 (O_1205,N_24013,N_24791);
or UO_1206 (O_1206,N_24696,N_24635);
nand UO_1207 (O_1207,N_24858,N_24608);
xnor UO_1208 (O_1208,N_24202,N_24811);
nand UO_1209 (O_1209,N_24957,N_24494);
and UO_1210 (O_1210,N_24777,N_24527);
nor UO_1211 (O_1211,N_24067,N_24340);
nor UO_1212 (O_1212,N_24613,N_24490);
or UO_1213 (O_1213,N_24257,N_24286);
xor UO_1214 (O_1214,N_24482,N_24227);
nor UO_1215 (O_1215,N_24275,N_24618);
nor UO_1216 (O_1216,N_24755,N_24053);
nand UO_1217 (O_1217,N_24839,N_24022);
or UO_1218 (O_1218,N_24279,N_24857);
nor UO_1219 (O_1219,N_24093,N_24910);
nand UO_1220 (O_1220,N_24036,N_24578);
or UO_1221 (O_1221,N_24948,N_24316);
nor UO_1222 (O_1222,N_24068,N_24500);
or UO_1223 (O_1223,N_24037,N_24586);
and UO_1224 (O_1224,N_24870,N_24051);
and UO_1225 (O_1225,N_24656,N_24482);
nor UO_1226 (O_1226,N_24926,N_24015);
and UO_1227 (O_1227,N_24333,N_24824);
and UO_1228 (O_1228,N_24584,N_24538);
nand UO_1229 (O_1229,N_24572,N_24950);
or UO_1230 (O_1230,N_24828,N_24699);
and UO_1231 (O_1231,N_24836,N_24138);
xnor UO_1232 (O_1232,N_24292,N_24608);
and UO_1233 (O_1233,N_24882,N_24255);
nand UO_1234 (O_1234,N_24445,N_24532);
xnor UO_1235 (O_1235,N_24356,N_24060);
xor UO_1236 (O_1236,N_24885,N_24572);
xor UO_1237 (O_1237,N_24222,N_24448);
nor UO_1238 (O_1238,N_24408,N_24192);
xor UO_1239 (O_1239,N_24187,N_24199);
nor UO_1240 (O_1240,N_24880,N_24594);
and UO_1241 (O_1241,N_24349,N_24763);
nand UO_1242 (O_1242,N_24724,N_24712);
and UO_1243 (O_1243,N_24919,N_24602);
nor UO_1244 (O_1244,N_24767,N_24157);
and UO_1245 (O_1245,N_24388,N_24042);
nor UO_1246 (O_1246,N_24409,N_24335);
xor UO_1247 (O_1247,N_24653,N_24792);
or UO_1248 (O_1248,N_24490,N_24617);
xnor UO_1249 (O_1249,N_24170,N_24221);
xor UO_1250 (O_1250,N_24958,N_24721);
nor UO_1251 (O_1251,N_24770,N_24167);
xnor UO_1252 (O_1252,N_24845,N_24555);
nand UO_1253 (O_1253,N_24834,N_24004);
nand UO_1254 (O_1254,N_24644,N_24669);
nor UO_1255 (O_1255,N_24206,N_24370);
xnor UO_1256 (O_1256,N_24204,N_24997);
or UO_1257 (O_1257,N_24264,N_24068);
nand UO_1258 (O_1258,N_24686,N_24636);
xor UO_1259 (O_1259,N_24292,N_24365);
xnor UO_1260 (O_1260,N_24782,N_24231);
or UO_1261 (O_1261,N_24336,N_24545);
nand UO_1262 (O_1262,N_24572,N_24638);
nor UO_1263 (O_1263,N_24054,N_24025);
nand UO_1264 (O_1264,N_24068,N_24063);
and UO_1265 (O_1265,N_24240,N_24648);
xnor UO_1266 (O_1266,N_24604,N_24447);
nor UO_1267 (O_1267,N_24233,N_24864);
and UO_1268 (O_1268,N_24375,N_24377);
nand UO_1269 (O_1269,N_24410,N_24219);
and UO_1270 (O_1270,N_24051,N_24376);
or UO_1271 (O_1271,N_24471,N_24750);
or UO_1272 (O_1272,N_24331,N_24818);
nand UO_1273 (O_1273,N_24550,N_24066);
and UO_1274 (O_1274,N_24216,N_24853);
or UO_1275 (O_1275,N_24906,N_24993);
xnor UO_1276 (O_1276,N_24049,N_24503);
nand UO_1277 (O_1277,N_24123,N_24329);
nand UO_1278 (O_1278,N_24695,N_24960);
nor UO_1279 (O_1279,N_24514,N_24838);
and UO_1280 (O_1280,N_24624,N_24353);
xor UO_1281 (O_1281,N_24971,N_24580);
and UO_1282 (O_1282,N_24388,N_24093);
nand UO_1283 (O_1283,N_24619,N_24310);
or UO_1284 (O_1284,N_24444,N_24220);
or UO_1285 (O_1285,N_24602,N_24929);
or UO_1286 (O_1286,N_24239,N_24119);
or UO_1287 (O_1287,N_24669,N_24850);
and UO_1288 (O_1288,N_24377,N_24810);
and UO_1289 (O_1289,N_24341,N_24565);
nand UO_1290 (O_1290,N_24126,N_24410);
and UO_1291 (O_1291,N_24018,N_24699);
xor UO_1292 (O_1292,N_24701,N_24944);
nor UO_1293 (O_1293,N_24288,N_24147);
and UO_1294 (O_1294,N_24969,N_24384);
nand UO_1295 (O_1295,N_24976,N_24404);
nand UO_1296 (O_1296,N_24980,N_24202);
nand UO_1297 (O_1297,N_24766,N_24019);
nor UO_1298 (O_1298,N_24775,N_24875);
xnor UO_1299 (O_1299,N_24366,N_24133);
or UO_1300 (O_1300,N_24048,N_24771);
and UO_1301 (O_1301,N_24624,N_24753);
xnor UO_1302 (O_1302,N_24914,N_24442);
xor UO_1303 (O_1303,N_24287,N_24487);
nor UO_1304 (O_1304,N_24945,N_24892);
xnor UO_1305 (O_1305,N_24122,N_24158);
or UO_1306 (O_1306,N_24243,N_24839);
xor UO_1307 (O_1307,N_24529,N_24181);
and UO_1308 (O_1308,N_24699,N_24566);
or UO_1309 (O_1309,N_24203,N_24450);
nand UO_1310 (O_1310,N_24696,N_24753);
nand UO_1311 (O_1311,N_24310,N_24902);
and UO_1312 (O_1312,N_24703,N_24788);
nand UO_1313 (O_1313,N_24740,N_24804);
nor UO_1314 (O_1314,N_24449,N_24652);
nand UO_1315 (O_1315,N_24015,N_24279);
nor UO_1316 (O_1316,N_24537,N_24665);
xnor UO_1317 (O_1317,N_24786,N_24818);
xnor UO_1318 (O_1318,N_24843,N_24779);
or UO_1319 (O_1319,N_24667,N_24910);
and UO_1320 (O_1320,N_24493,N_24235);
nand UO_1321 (O_1321,N_24708,N_24667);
nand UO_1322 (O_1322,N_24032,N_24276);
and UO_1323 (O_1323,N_24146,N_24266);
and UO_1324 (O_1324,N_24672,N_24378);
xnor UO_1325 (O_1325,N_24171,N_24273);
or UO_1326 (O_1326,N_24191,N_24943);
and UO_1327 (O_1327,N_24618,N_24249);
nor UO_1328 (O_1328,N_24085,N_24564);
nand UO_1329 (O_1329,N_24872,N_24526);
nand UO_1330 (O_1330,N_24497,N_24929);
xor UO_1331 (O_1331,N_24034,N_24773);
and UO_1332 (O_1332,N_24046,N_24388);
nor UO_1333 (O_1333,N_24667,N_24229);
nor UO_1334 (O_1334,N_24731,N_24892);
nand UO_1335 (O_1335,N_24696,N_24639);
and UO_1336 (O_1336,N_24480,N_24818);
xor UO_1337 (O_1337,N_24776,N_24529);
or UO_1338 (O_1338,N_24528,N_24371);
xnor UO_1339 (O_1339,N_24732,N_24044);
or UO_1340 (O_1340,N_24515,N_24854);
or UO_1341 (O_1341,N_24073,N_24785);
nor UO_1342 (O_1342,N_24460,N_24367);
or UO_1343 (O_1343,N_24978,N_24536);
xor UO_1344 (O_1344,N_24437,N_24248);
nor UO_1345 (O_1345,N_24664,N_24136);
nand UO_1346 (O_1346,N_24421,N_24638);
xnor UO_1347 (O_1347,N_24424,N_24804);
and UO_1348 (O_1348,N_24123,N_24224);
nand UO_1349 (O_1349,N_24474,N_24233);
xor UO_1350 (O_1350,N_24666,N_24605);
nor UO_1351 (O_1351,N_24954,N_24043);
xnor UO_1352 (O_1352,N_24124,N_24636);
or UO_1353 (O_1353,N_24945,N_24198);
nor UO_1354 (O_1354,N_24991,N_24530);
nor UO_1355 (O_1355,N_24864,N_24295);
nor UO_1356 (O_1356,N_24052,N_24360);
nand UO_1357 (O_1357,N_24201,N_24535);
nand UO_1358 (O_1358,N_24174,N_24077);
nor UO_1359 (O_1359,N_24193,N_24642);
and UO_1360 (O_1360,N_24986,N_24611);
xor UO_1361 (O_1361,N_24961,N_24784);
nand UO_1362 (O_1362,N_24995,N_24304);
and UO_1363 (O_1363,N_24636,N_24207);
or UO_1364 (O_1364,N_24840,N_24859);
or UO_1365 (O_1365,N_24431,N_24413);
nor UO_1366 (O_1366,N_24371,N_24029);
nor UO_1367 (O_1367,N_24613,N_24059);
and UO_1368 (O_1368,N_24402,N_24326);
nand UO_1369 (O_1369,N_24075,N_24226);
and UO_1370 (O_1370,N_24902,N_24409);
and UO_1371 (O_1371,N_24091,N_24360);
and UO_1372 (O_1372,N_24462,N_24193);
or UO_1373 (O_1373,N_24864,N_24451);
and UO_1374 (O_1374,N_24710,N_24950);
xor UO_1375 (O_1375,N_24097,N_24268);
nand UO_1376 (O_1376,N_24327,N_24305);
nand UO_1377 (O_1377,N_24065,N_24817);
xor UO_1378 (O_1378,N_24422,N_24404);
nor UO_1379 (O_1379,N_24624,N_24360);
xor UO_1380 (O_1380,N_24652,N_24471);
nor UO_1381 (O_1381,N_24246,N_24133);
nand UO_1382 (O_1382,N_24952,N_24642);
and UO_1383 (O_1383,N_24217,N_24910);
and UO_1384 (O_1384,N_24403,N_24077);
or UO_1385 (O_1385,N_24760,N_24786);
xnor UO_1386 (O_1386,N_24535,N_24169);
or UO_1387 (O_1387,N_24143,N_24523);
or UO_1388 (O_1388,N_24726,N_24283);
nor UO_1389 (O_1389,N_24160,N_24862);
nor UO_1390 (O_1390,N_24712,N_24651);
nand UO_1391 (O_1391,N_24901,N_24926);
nand UO_1392 (O_1392,N_24892,N_24051);
and UO_1393 (O_1393,N_24934,N_24565);
or UO_1394 (O_1394,N_24007,N_24329);
and UO_1395 (O_1395,N_24953,N_24120);
or UO_1396 (O_1396,N_24032,N_24320);
xor UO_1397 (O_1397,N_24251,N_24443);
nand UO_1398 (O_1398,N_24006,N_24815);
nor UO_1399 (O_1399,N_24022,N_24550);
nand UO_1400 (O_1400,N_24911,N_24646);
and UO_1401 (O_1401,N_24133,N_24706);
nand UO_1402 (O_1402,N_24277,N_24157);
xnor UO_1403 (O_1403,N_24828,N_24759);
nand UO_1404 (O_1404,N_24288,N_24567);
xor UO_1405 (O_1405,N_24929,N_24226);
or UO_1406 (O_1406,N_24691,N_24997);
and UO_1407 (O_1407,N_24541,N_24901);
nand UO_1408 (O_1408,N_24731,N_24620);
xnor UO_1409 (O_1409,N_24915,N_24636);
nor UO_1410 (O_1410,N_24480,N_24474);
xnor UO_1411 (O_1411,N_24821,N_24666);
and UO_1412 (O_1412,N_24574,N_24244);
nor UO_1413 (O_1413,N_24729,N_24706);
xor UO_1414 (O_1414,N_24608,N_24677);
and UO_1415 (O_1415,N_24834,N_24307);
nor UO_1416 (O_1416,N_24808,N_24270);
xnor UO_1417 (O_1417,N_24888,N_24313);
or UO_1418 (O_1418,N_24443,N_24942);
and UO_1419 (O_1419,N_24810,N_24244);
and UO_1420 (O_1420,N_24258,N_24526);
nand UO_1421 (O_1421,N_24746,N_24736);
nand UO_1422 (O_1422,N_24572,N_24205);
or UO_1423 (O_1423,N_24575,N_24580);
nor UO_1424 (O_1424,N_24820,N_24817);
and UO_1425 (O_1425,N_24390,N_24211);
and UO_1426 (O_1426,N_24574,N_24973);
or UO_1427 (O_1427,N_24422,N_24641);
xnor UO_1428 (O_1428,N_24229,N_24321);
xnor UO_1429 (O_1429,N_24172,N_24048);
nand UO_1430 (O_1430,N_24041,N_24323);
and UO_1431 (O_1431,N_24753,N_24229);
nor UO_1432 (O_1432,N_24726,N_24423);
xor UO_1433 (O_1433,N_24912,N_24413);
xor UO_1434 (O_1434,N_24590,N_24336);
nor UO_1435 (O_1435,N_24664,N_24103);
nand UO_1436 (O_1436,N_24569,N_24515);
xnor UO_1437 (O_1437,N_24367,N_24703);
nand UO_1438 (O_1438,N_24632,N_24012);
nand UO_1439 (O_1439,N_24820,N_24789);
nand UO_1440 (O_1440,N_24179,N_24430);
nand UO_1441 (O_1441,N_24373,N_24814);
xnor UO_1442 (O_1442,N_24552,N_24046);
xnor UO_1443 (O_1443,N_24401,N_24915);
xnor UO_1444 (O_1444,N_24257,N_24438);
and UO_1445 (O_1445,N_24055,N_24675);
nand UO_1446 (O_1446,N_24382,N_24294);
or UO_1447 (O_1447,N_24962,N_24998);
xor UO_1448 (O_1448,N_24402,N_24723);
or UO_1449 (O_1449,N_24397,N_24534);
nor UO_1450 (O_1450,N_24568,N_24888);
nand UO_1451 (O_1451,N_24578,N_24639);
or UO_1452 (O_1452,N_24906,N_24428);
and UO_1453 (O_1453,N_24213,N_24380);
nand UO_1454 (O_1454,N_24647,N_24605);
nand UO_1455 (O_1455,N_24780,N_24163);
nand UO_1456 (O_1456,N_24668,N_24737);
nand UO_1457 (O_1457,N_24965,N_24258);
nor UO_1458 (O_1458,N_24072,N_24684);
nand UO_1459 (O_1459,N_24219,N_24465);
nor UO_1460 (O_1460,N_24649,N_24250);
xor UO_1461 (O_1461,N_24943,N_24542);
nor UO_1462 (O_1462,N_24995,N_24361);
nand UO_1463 (O_1463,N_24258,N_24524);
or UO_1464 (O_1464,N_24572,N_24481);
nand UO_1465 (O_1465,N_24353,N_24847);
or UO_1466 (O_1466,N_24676,N_24711);
xnor UO_1467 (O_1467,N_24373,N_24675);
and UO_1468 (O_1468,N_24695,N_24313);
or UO_1469 (O_1469,N_24568,N_24227);
or UO_1470 (O_1470,N_24085,N_24952);
or UO_1471 (O_1471,N_24297,N_24464);
xnor UO_1472 (O_1472,N_24667,N_24958);
or UO_1473 (O_1473,N_24807,N_24639);
or UO_1474 (O_1474,N_24519,N_24153);
xor UO_1475 (O_1475,N_24799,N_24802);
and UO_1476 (O_1476,N_24206,N_24694);
and UO_1477 (O_1477,N_24560,N_24926);
nor UO_1478 (O_1478,N_24248,N_24289);
or UO_1479 (O_1479,N_24307,N_24596);
and UO_1480 (O_1480,N_24399,N_24172);
or UO_1481 (O_1481,N_24978,N_24550);
nor UO_1482 (O_1482,N_24562,N_24649);
xnor UO_1483 (O_1483,N_24559,N_24894);
nand UO_1484 (O_1484,N_24013,N_24094);
xnor UO_1485 (O_1485,N_24440,N_24002);
xor UO_1486 (O_1486,N_24784,N_24696);
and UO_1487 (O_1487,N_24787,N_24500);
xor UO_1488 (O_1488,N_24706,N_24642);
nand UO_1489 (O_1489,N_24715,N_24144);
or UO_1490 (O_1490,N_24378,N_24998);
or UO_1491 (O_1491,N_24487,N_24855);
nor UO_1492 (O_1492,N_24085,N_24589);
and UO_1493 (O_1493,N_24214,N_24918);
nand UO_1494 (O_1494,N_24980,N_24972);
nand UO_1495 (O_1495,N_24209,N_24396);
xnor UO_1496 (O_1496,N_24890,N_24566);
nor UO_1497 (O_1497,N_24687,N_24700);
xnor UO_1498 (O_1498,N_24773,N_24916);
nand UO_1499 (O_1499,N_24711,N_24846);
xnor UO_1500 (O_1500,N_24536,N_24422);
xor UO_1501 (O_1501,N_24452,N_24655);
nand UO_1502 (O_1502,N_24642,N_24859);
and UO_1503 (O_1503,N_24164,N_24400);
or UO_1504 (O_1504,N_24798,N_24416);
nor UO_1505 (O_1505,N_24587,N_24088);
nor UO_1506 (O_1506,N_24734,N_24134);
nand UO_1507 (O_1507,N_24850,N_24196);
xnor UO_1508 (O_1508,N_24370,N_24060);
nor UO_1509 (O_1509,N_24664,N_24482);
nand UO_1510 (O_1510,N_24192,N_24801);
and UO_1511 (O_1511,N_24683,N_24227);
and UO_1512 (O_1512,N_24942,N_24082);
nor UO_1513 (O_1513,N_24986,N_24638);
nand UO_1514 (O_1514,N_24626,N_24565);
nor UO_1515 (O_1515,N_24095,N_24230);
nor UO_1516 (O_1516,N_24994,N_24178);
nor UO_1517 (O_1517,N_24530,N_24963);
nor UO_1518 (O_1518,N_24997,N_24007);
or UO_1519 (O_1519,N_24189,N_24915);
or UO_1520 (O_1520,N_24062,N_24841);
xnor UO_1521 (O_1521,N_24164,N_24853);
nand UO_1522 (O_1522,N_24317,N_24670);
xor UO_1523 (O_1523,N_24963,N_24630);
xnor UO_1524 (O_1524,N_24376,N_24428);
or UO_1525 (O_1525,N_24446,N_24696);
nand UO_1526 (O_1526,N_24023,N_24620);
and UO_1527 (O_1527,N_24669,N_24832);
or UO_1528 (O_1528,N_24596,N_24609);
nor UO_1529 (O_1529,N_24661,N_24465);
and UO_1530 (O_1530,N_24562,N_24696);
and UO_1531 (O_1531,N_24344,N_24866);
or UO_1532 (O_1532,N_24349,N_24389);
nor UO_1533 (O_1533,N_24146,N_24806);
xnor UO_1534 (O_1534,N_24670,N_24032);
or UO_1535 (O_1535,N_24199,N_24894);
or UO_1536 (O_1536,N_24323,N_24357);
or UO_1537 (O_1537,N_24352,N_24604);
or UO_1538 (O_1538,N_24869,N_24032);
xnor UO_1539 (O_1539,N_24212,N_24170);
xnor UO_1540 (O_1540,N_24398,N_24324);
xnor UO_1541 (O_1541,N_24385,N_24834);
and UO_1542 (O_1542,N_24919,N_24281);
or UO_1543 (O_1543,N_24361,N_24669);
or UO_1544 (O_1544,N_24258,N_24795);
xor UO_1545 (O_1545,N_24425,N_24118);
nand UO_1546 (O_1546,N_24995,N_24138);
or UO_1547 (O_1547,N_24930,N_24290);
xor UO_1548 (O_1548,N_24619,N_24412);
nand UO_1549 (O_1549,N_24697,N_24462);
xor UO_1550 (O_1550,N_24034,N_24806);
and UO_1551 (O_1551,N_24248,N_24152);
nor UO_1552 (O_1552,N_24297,N_24891);
xnor UO_1553 (O_1553,N_24472,N_24528);
nor UO_1554 (O_1554,N_24096,N_24755);
nor UO_1555 (O_1555,N_24298,N_24795);
and UO_1556 (O_1556,N_24557,N_24038);
and UO_1557 (O_1557,N_24669,N_24497);
or UO_1558 (O_1558,N_24463,N_24532);
and UO_1559 (O_1559,N_24381,N_24596);
xor UO_1560 (O_1560,N_24680,N_24440);
nand UO_1561 (O_1561,N_24646,N_24753);
xor UO_1562 (O_1562,N_24161,N_24340);
or UO_1563 (O_1563,N_24754,N_24649);
nor UO_1564 (O_1564,N_24809,N_24573);
xnor UO_1565 (O_1565,N_24482,N_24438);
nand UO_1566 (O_1566,N_24653,N_24320);
or UO_1567 (O_1567,N_24842,N_24147);
xor UO_1568 (O_1568,N_24948,N_24083);
or UO_1569 (O_1569,N_24602,N_24208);
or UO_1570 (O_1570,N_24251,N_24878);
nand UO_1571 (O_1571,N_24860,N_24505);
and UO_1572 (O_1572,N_24141,N_24702);
and UO_1573 (O_1573,N_24323,N_24308);
nand UO_1574 (O_1574,N_24424,N_24063);
nand UO_1575 (O_1575,N_24284,N_24755);
xnor UO_1576 (O_1576,N_24311,N_24198);
nor UO_1577 (O_1577,N_24731,N_24867);
xnor UO_1578 (O_1578,N_24076,N_24059);
or UO_1579 (O_1579,N_24744,N_24453);
and UO_1580 (O_1580,N_24447,N_24463);
nor UO_1581 (O_1581,N_24232,N_24149);
nand UO_1582 (O_1582,N_24374,N_24323);
nor UO_1583 (O_1583,N_24935,N_24646);
xnor UO_1584 (O_1584,N_24034,N_24341);
or UO_1585 (O_1585,N_24125,N_24709);
nand UO_1586 (O_1586,N_24905,N_24515);
nor UO_1587 (O_1587,N_24338,N_24244);
nor UO_1588 (O_1588,N_24352,N_24923);
or UO_1589 (O_1589,N_24479,N_24196);
xnor UO_1590 (O_1590,N_24488,N_24929);
nand UO_1591 (O_1591,N_24552,N_24032);
nor UO_1592 (O_1592,N_24444,N_24426);
and UO_1593 (O_1593,N_24440,N_24833);
nor UO_1594 (O_1594,N_24770,N_24488);
or UO_1595 (O_1595,N_24636,N_24213);
and UO_1596 (O_1596,N_24802,N_24195);
nor UO_1597 (O_1597,N_24892,N_24088);
or UO_1598 (O_1598,N_24760,N_24516);
xor UO_1599 (O_1599,N_24158,N_24718);
nand UO_1600 (O_1600,N_24154,N_24048);
nor UO_1601 (O_1601,N_24469,N_24067);
or UO_1602 (O_1602,N_24400,N_24241);
or UO_1603 (O_1603,N_24258,N_24112);
and UO_1604 (O_1604,N_24442,N_24248);
or UO_1605 (O_1605,N_24450,N_24576);
nand UO_1606 (O_1606,N_24221,N_24871);
nand UO_1607 (O_1607,N_24296,N_24696);
and UO_1608 (O_1608,N_24620,N_24704);
xor UO_1609 (O_1609,N_24031,N_24994);
and UO_1610 (O_1610,N_24478,N_24183);
or UO_1611 (O_1611,N_24894,N_24461);
nand UO_1612 (O_1612,N_24288,N_24763);
xor UO_1613 (O_1613,N_24167,N_24249);
nand UO_1614 (O_1614,N_24466,N_24091);
or UO_1615 (O_1615,N_24001,N_24503);
nand UO_1616 (O_1616,N_24388,N_24280);
and UO_1617 (O_1617,N_24923,N_24019);
nand UO_1618 (O_1618,N_24462,N_24952);
xnor UO_1619 (O_1619,N_24360,N_24890);
and UO_1620 (O_1620,N_24244,N_24333);
xor UO_1621 (O_1621,N_24398,N_24695);
nor UO_1622 (O_1622,N_24045,N_24248);
or UO_1623 (O_1623,N_24900,N_24520);
and UO_1624 (O_1624,N_24212,N_24721);
nand UO_1625 (O_1625,N_24358,N_24629);
nand UO_1626 (O_1626,N_24214,N_24669);
and UO_1627 (O_1627,N_24947,N_24417);
and UO_1628 (O_1628,N_24916,N_24775);
nand UO_1629 (O_1629,N_24107,N_24194);
nand UO_1630 (O_1630,N_24091,N_24130);
and UO_1631 (O_1631,N_24640,N_24104);
and UO_1632 (O_1632,N_24608,N_24937);
and UO_1633 (O_1633,N_24562,N_24745);
nor UO_1634 (O_1634,N_24922,N_24110);
and UO_1635 (O_1635,N_24618,N_24903);
and UO_1636 (O_1636,N_24175,N_24907);
xnor UO_1637 (O_1637,N_24584,N_24050);
or UO_1638 (O_1638,N_24669,N_24539);
or UO_1639 (O_1639,N_24240,N_24626);
or UO_1640 (O_1640,N_24731,N_24053);
nand UO_1641 (O_1641,N_24731,N_24415);
and UO_1642 (O_1642,N_24108,N_24621);
or UO_1643 (O_1643,N_24124,N_24449);
and UO_1644 (O_1644,N_24747,N_24880);
or UO_1645 (O_1645,N_24651,N_24307);
or UO_1646 (O_1646,N_24093,N_24977);
xor UO_1647 (O_1647,N_24771,N_24524);
nor UO_1648 (O_1648,N_24862,N_24506);
xor UO_1649 (O_1649,N_24896,N_24201);
and UO_1650 (O_1650,N_24931,N_24755);
and UO_1651 (O_1651,N_24858,N_24167);
or UO_1652 (O_1652,N_24090,N_24461);
nor UO_1653 (O_1653,N_24881,N_24681);
nand UO_1654 (O_1654,N_24060,N_24349);
nand UO_1655 (O_1655,N_24444,N_24755);
xnor UO_1656 (O_1656,N_24078,N_24803);
and UO_1657 (O_1657,N_24552,N_24726);
nor UO_1658 (O_1658,N_24798,N_24819);
xnor UO_1659 (O_1659,N_24438,N_24602);
xor UO_1660 (O_1660,N_24721,N_24014);
xor UO_1661 (O_1661,N_24587,N_24322);
xor UO_1662 (O_1662,N_24971,N_24486);
or UO_1663 (O_1663,N_24007,N_24265);
nand UO_1664 (O_1664,N_24164,N_24263);
nor UO_1665 (O_1665,N_24346,N_24736);
and UO_1666 (O_1666,N_24227,N_24349);
and UO_1667 (O_1667,N_24998,N_24909);
xnor UO_1668 (O_1668,N_24020,N_24292);
and UO_1669 (O_1669,N_24935,N_24860);
and UO_1670 (O_1670,N_24491,N_24403);
xor UO_1671 (O_1671,N_24272,N_24401);
nor UO_1672 (O_1672,N_24982,N_24038);
nand UO_1673 (O_1673,N_24825,N_24833);
xor UO_1674 (O_1674,N_24093,N_24334);
nand UO_1675 (O_1675,N_24041,N_24908);
xor UO_1676 (O_1676,N_24936,N_24506);
or UO_1677 (O_1677,N_24273,N_24773);
or UO_1678 (O_1678,N_24201,N_24871);
nand UO_1679 (O_1679,N_24286,N_24002);
nor UO_1680 (O_1680,N_24259,N_24775);
and UO_1681 (O_1681,N_24183,N_24669);
nor UO_1682 (O_1682,N_24207,N_24327);
or UO_1683 (O_1683,N_24014,N_24108);
nand UO_1684 (O_1684,N_24506,N_24637);
nand UO_1685 (O_1685,N_24162,N_24359);
xor UO_1686 (O_1686,N_24701,N_24542);
and UO_1687 (O_1687,N_24054,N_24296);
xor UO_1688 (O_1688,N_24497,N_24491);
nor UO_1689 (O_1689,N_24926,N_24161);
xnor UO_1690 (O_1690,N_24760,N_24521);
xnor UO_1691 (O_1691,N_24233,N_24097);
nand UO_1692 (O_1692,N_24766,N_24101);
xor UO_1693 (O_1693,N_24369,N_24735);
nor UO_1694 (O_1694,N_24715,N_24361);
or UO_1695 (O_1695,N_24428,N_24081);
xnor UO_1696 (O_1696,N_24382,N_24160);
or UO_1697 (O_1697,N_24620,N_24604);
nand UO_1698 (O_1698,N_24973,N_24915);
nor UO_1699 (O_1699,N_24098,N_24538);
xor UO_1700 (O_1700,N_24654,N_24955);
nand UO_1701 (O_1701,N_24485,N_24773);
or UO_1702 (O_1702,N_24782,N_24847);
or UO_1703 (O_1703,N_24430,N_24851);
nand UO_1704 (O_1704,N_24662,N_24248);
and UO_1705 (O_1705,N_24671,N_24824);
xnor UO_1706 (O_1706,N_24667,N_24394);
nor UO_1707 (O_1707,N_24278,N_24083);
or UO_1708 (O_1708,N_24747,N_24335);
and UO_1709 (O_1709,N_24377,N_24657);
or UO_1710 (O_1710,N_24068,N_24341);
xor UO_1711 (O_1711,N_24077,N_24122);
xor UO_1712 (O_1712,N_24936,N_24474);
and UO_1713 (O_1713,N_24239,N_24168);
nor UO_1714 (O_1714,N_24366,N_24030);
and UO_1715 (O_1715,N_24437,N_24042);
or UO_1716 (O_1716,N_24510,N_24174);
and UO_1717 (O_1717,N_24628,N_24707);
or UO_1718 (O_1718,N_24475,N_24329);
nor UO_1719 (O_1719,N_24572,N_24606);
or UO_1720 (O_1720,N_24437,N_24376);
xnor UO_1721 (O_1721,N_24266,N_24613);
or UO_1722 (O_1722,N_24006,N_24749);
and UO_1723 (O_1723,N_24789,N_24573);
nor UO_1724 (O_1724,N_24311,N_24728);
nand UO_1725 (O_1725,N_24483,N_24975);
and UO_1726 (O_1726,N_24583,N_24574);
nand UO_1727 (O_1727,N_24306,N_24089);
or UO_1728 (O_1728,N_24791,N_24700);
xnor UO_1729 (O_1729,N_24372,N_24143);
and UO_1730 (O_1730,N_24118,N_24657);
xor UO_1731 (O_1731,N_24475,N_24625);
and UO_1732 (O_1732,N_24016,N_24415);
nor UO_1733 (O_1733,N_24915,N_24709);
and UO_1734 (O_1734,N_24652,N_24075);
and UO_1735 (O_1735,N_24302,N_24716);
xnor UO_1736 (O_1736,N_24300,N_24998);
nor UO_1737 (O_1737,N_24966,N_24692);
or UO_1738 (O_1738,N_24705,N_24080);
nand UO_1739 (O_1739,N_24578,N_24137);
nand UO_1740 (O_1740,N_24858,N_24541);
or UO_1741 (O_1741,N_24361,N_24190);
nor UO_1742 (O_1742,N_24650,N_24536);
xor UO_1743 (O_1743,N_24585,N_24041);
xor UO_1744 (O_1744,N_24497,N_24108);
nor UO_1745 (O_1745,N_24911,N_24034);
xor UO_1746 (O_1746,N_24816,N_24487);
xnor UO_1747 (O_1747,N_24559,N_24051);
nand UO_1748 (O_1748,N_24167,N_24963);
or UO_1749 (O_1749,N_24251,N_24302);
nand UO_1750 (O_1750,N_24274,N_24941);
nand UO_1751 (O_1751,N_24796,N_24051);
and UO_1752 (O_1752,N_24359,N_24986);
or UO_1753 (O_1753,N_24859,N_24400);
or UO_1754 (O_1754,N_24367,N_24167);
and UO_1755 (O_1755,N_24034,N_24351);
nand UO_1756 (O_1756,N_24470,N_24221);
nand UO_1757 (O_1757,N_24229,N_24736);
xor UO_1758 (O_1758,N_24211,N_24069);
xor UO_1759 (O_1759,N_24067,N_24125);
or UO_1760 (O_1760,N_24147,N_24119);
nand UO_1761 (O_1761,N_24009,N_24722);
xor UO_1762 (O_1762,N_24738,N_24836);
nor UO_1763 (O_1763,N_24228,N_24978);
xor UO_1764 (O_1764,N_24792,N_24442);
xor UO_1765 (O_1765,N_24274,N_24641);
nor UO_1766 (O_1766,N_24931,N_24783);
and UO_1767 (O_1767,N_24834,N_24929);
and UO_1768 (O_1768,N_24231,N_24273);
and UO_1769 (O_1769,N_24416,N_24408);
nand UO_1770 (O_1770,N_24544,N_24722);
or UO_1771 (O_1771,N_24872,N_24016);
nor UO_1772 (O_1772,N_24003,N_24241);
and UO_1773 (O_1773,N_24093,N_24353);
or UO_1774 (O_1774,N_24406,N_24109);
or UO_1775 (O_1775,N_24687,N_24528);
nor UO_1776 (O_1776,N_24698,N_24514);
xnor UO_1777 (O_1777,N_24225,N_24777);
nor UO_1778 (O_1778,N_24000,N_24027);
nor UO_1779 (O_1779,N_24118,N_24907);
and UO_1780 (O_1780,N_24589,N_24954);
and UO_1781 (O_1781,N_24128,N_24356);
and UO_1782 (O_1782,N_24270,N_24957);
nor UO_1783 (O_1783,N_24802,N_24397);
nor UO_1784 (O_1784,N_24446,N_24205);
or UO_1785 (O_1785,N_24218,N_24449);
nor UO_1786 (O_1786,N_24092,N_24673);
or UO_1787 (O_1787,N_24500,N_24931);
nor UO_1788 (O_1788,N_24707,N_24885);
nand UO_1789 (O_1789,N_24186,N_24571);
xor UO_1790 (O_1790,N_24827,N_24725);
and UO_1791 (O_1791,N_24188,N_24080);
and UO_1792 (O_1792,N_24087,N_24890);
and UO_1793 (O_1793,N_24897,N_24111);
nand UO_1794 (O_1794,N_24453,N_24198);
and UO_1795 (O_1795,N_24395,N_24867);
and UO_1796 (O_1796,N_24333,N_24921);
xor UO_1797 (O_1797,N_24594,N_24673);
and UO_1798 (O_1798,N_24325,N_24884);
and UO_1799 (O_1799,N_24111,N_24390);
nor UO_1800 (O_1800,N_24953,N_24430);
and UO_1801 (O_1801,N_24234,N_24654);
and UO_1802 (O_1802,N_24016,N_24592);
or UO_1803 (O_1803,N_24130,N_24397);
xor UO_1804 (O_1804,N_24726,N_24652);
xor UO_1805 (O_1805,N_24600,N_24324);
nand UO_1806 (O_1806,N_24584,N_24984);
nor UO_1807 (O_1807,N_24763,N_24303);
or UO_1808 (O_1808,N_24910,N_24543);
or UO_1809 (O_1809,N_24249,N_24475);
nand UO_1810 (O_1810,N_24288,N_24947);
nand UO_1811 (O_1811,N_24812,N_24098);
nand UO_1812 (O_1812,N_24563,N_24494);
or UO_1813 (O_1813,N_24162,N_24806);
nand UO_1814 (O_1814,N_24709,N_24910);
xor UO_1815 (O_1815,N_24014,N_24442);
nand UO_1816 (O_1816,N_24112,N_24726);
xnor UO_1817 (O_1817,N_24501,N_24026);
xnor UO_1818 (O_1818,N_24374,N_24219);
xnor UO_1819 (O_1819,N_24471,N_24499);
xor UO_1820 (O_1820,N_24529,N_24454);
and UO_1821 (O_1821,N_24764,N_24415);
nand UO_1822 (O_1822,N_24451,N_24076);
nand UO_1823 (O_1823,N_24124,N_24880);
or UO_1824 (O_1824,N_24293,N_24768);
nand UO_1825 (O_1825,N_24244,N_24603);
xnor UO_1826 (O_1826,N_24367,N_24613);
nor UO_1827 (O_1827,N_24218,N_24338);
and UO_1828 (O_1828,N_24776,N_24180);
nor UO_1829 (O_1829,N_24659,N_24687);
nor UO_1830 (O_1830,N_24700,N_24899);
and UO_1831 (O_1831,N_24110,N_24267);
and UO_1832 (O_1832,N_24283,N_24543);
nand UO_1833 (O_1833,N_24839,N_24828);
nor UO_1834 (O_1834,N_24448,N_24390);
nor UO_1835 (O_1835,N_24270,N_24082);
nand UO_1836 (O_1836,N_24335,N_24316);
nor UO_1837 (O_1837,N_24467,N_24710);
and UO_1838 (O_1838,N_24406,N_24865);
and UO_1839 (O_1839,N_24868,N_24038);
and UO_1840 (O_1840,N_24066,N_24334);
and UO_1841 (O_1841,N_24967,N_24431);
or UO_1842 (O_1842,N_24311,N_24168);
nand UO_1843 (O_1843,N_24734,N_24455);
nand UO_1844 (O_1844,N_24220,N_24446);
and UO_1845 (O_1845,N_24462,N_24457);
nand UO_1846 (O_1846,N_24241,N_24201);
xnor UO_1847 (O_1847,N_24702,N_24774);
nand UO_1848 (O_1848,N_24798,N_24157);
or UO_1849 (O_1849,N_24605,N_24221);
nor UO_1850 (O_1850,N_24942,N_24722);
and UO_1851 (O_1851,N_24184,N_24176);
xor UO_1852 (O_1852,N_24886,N_24745);
and UO_1853 (O_1853,N_24051,N_24447);
or UO_1854 (O_1854,N_24293,N_24395);
nand UO_1855 (O_1855,N_24374,N_24422);
and UO_1856 (O_1856,N_24354,N_24163);
xor UO_1857 (O_1857,N_24398,N_24248);
nand UO_1858 (O_1858,N_24952,N_24901);
nor UO_1859 (O_1859,N_24211,N_24712);
or UO_1860 (O_1860,N_24063,N_24435);
or UO_1861 (O_1861,N_24373,N_24642);
and UO_1862 (O_1862,N_24007,N_24127);
nor UO_1863 (O_1863,N_24355,N_24883);
xnor UO_1864 (O_1864,N_24860,N_24697);
or UO_1865 (O_1865,N_24335,N_24158);
nand UO_1866 (O_1866,N_24502,N_24826);
xor UO_1867 (O_1867,N_24004,N_24380);
and UO_1868 (O_1868,N_24625,N_24765);
and UO_1869 (O_1869,N_24599,N_24832);
or UO_1870 (O_1870,N_24863,N_24197);
xor UO_1871 (O_1871,N_24371,N_24864);
nor UO_1872 (O_1872,N_24938,N_24874);
xor UO_1873 (O_1873,N_24038,N_24345);
xor UO_1874 (O_1874,N_24676,N_24864);
and UO_1875 (O_1875,N_24480,N_24896);
nor UO_1876 (O_1876,N_24332,N_24198);
or UO_1877 (O_1877,N_24908,N_24963);
and UO_1878 (O_1878,N_24393,N_24638);
xnor UO_1879 (O_1879,N_24702,N_24509);
nor UO_1880 (O_1880,N_24390,N_24050);
or UO_1881 (O_1881,N_24250,N_24232);
and UO_1882 (O_1882,N_24711,N_24243);
or UO_1883 (O_1883,N_24130,N_24782);
xnor UO_1884 (O_1884,N_24523,N_24894);
nor UO_1885 (O_1885,N_24227,N_24489);
and UO_1886 (O_1886,N_24257,N_24895);
xor UO_1887 (O_1887,N_24025,N_24081);
nand UO_1888 (O_1888,N_24191,N_24531);
or UO_1889 (O_1889,N_24968,N_24476);
and UO_1890 (O_1890,N_24134,N_24678);
xor UO_1891 (O_1891,N_24069,N_24885);
nor UO_1892 (O_1892,N_24289,N_24609);
and UO_1893 (O_1893,N_24583,N_24695);
and UO_1894 (O_1894,N_24126,N_24456);
or UO_1895 (O_1895,N_24840,N_24526);
nand UO_1896 (O_1896,N_24171,N_24476);
and UO_1897 (O_1897,N_24496,N_24079);
and UO_1898 (O_1898,N_24549,N_24314);
xor UO_1899 (O_1899,N_24397,N_24492);
xor UO_1900 (O_1900,N_24002,N_24314);
xor UO_1901 (O_1901,N_24988,N_24357);
nor UO_1902 (O_1902,N_24660,N_24860);
xnor UO_1903 (O_1903,N_24542,N_24307);
nand UO_1904 (O_1904,N_24373,N_24755);
nand UO_1905 (O_1905,N_24860,N_24279);
xnor UO_1906 (O_1906,N_24312,N_24292);
and UO_1907 (O_1907,N_24239,N_24078);
nand UO_1908 (O_1908,N_24527,N_24899);
nor UO_1909 (O_1909,N_24781,N_24119);
or UO_1910 (O_1910,N_24190,N_24112);
nor UO_1911 (O_1911,N_24338,N_24362);
xnor UO_1912 (O_1912,N_24265,N_24149);
or UO_1913 (O_1913,N_24247,N_24929);
nand UO_1914 (O_1914,N_24708,N_24946);
nor UO_1915 (O_1915,N_24062,N_24228);
nor UO_1916 (O_1916,N_24538,N_24070);
xor UO_1917 (O_1917,N_24204,N_24987);
nand UO_1918 (O_1918,N_24898,N_24067);
nand UO_1919 (O_1919,N_24064,N_24227);
nor UO_1920 (O_1920,N_24201,N_24376);
and UO_1921 (O_1921,N_24556,N_24794);
and UO_1922 (O_1922,N_24413,N_24242);
nand UO_1923 (O_1923,N_24203,N_24806);
xnor UO_1924 (O_1924,N_24562,N_24980);
and UO_1925 (O_1925,N_24389,N_24340);
and UO_1926 (O_1926,N_24306,N_24636);
or UO_1927 (O_1927,N_24108,N_24527);
nand UO_1928 (O_1928,N_24579,N_24788);
nand UO_1929 (O_1929,N_24861,N_24092);
nand UO_1930 (O_1930,N_24876,N_24297);
nand UO_1931 (O_1931,N_24924,N_24424);
or UO_1932 (O_1932,N_24744,N_24447);
xor UO_1933 (O_1933,N_24168,N_24918);
and UO_1934 (O_1934,N_24052,N_24993);
xor UO_1935 (O_1935,N_24599,N_24750);
and UO_1936 (O_1936,N_24385,N_24066);
nor UO_1937 (O_1937,N_24792,N_24242);
or UO_1938 (O_1938,N_24445,N_24515);
or UO_1939 (O_1939,N_24048,N_24029);
nand UO_1940 (O_1940,N_24685,N_24096);
nand UO_1941 (O_1941,N_24306,N_24339);
or UO_1942 (O_1942,N_24413,N_24758);
xor UO_1943 (O_1943,N_24985,N_24878);
xor UO_1944 (O_1944,N_24731,N_24133);
and UO_1945 (O_1945,N_24343,N_24917);
xnor UO_1946 (O_1946,N_24396,N_24997);
or UO_1947 (O_1947,N_24937,N_24602);
nand UO_1948 (O_1948,N_24315,N_24454);
or UO_1949 (O_1949,N_24646,N_24181);
and UO_1950 (O_1950,N_24506,N_24799);
xor UO_1951 (O_1951,N_24295,N_24651);
nor UO_1952 (O_1952,N_24085,N_24871);
or UO_1953 (O_1953,N_24277,N_24131);
xor UO_1954 (O_1954,N_24741,N_24209);
nand UO_1955 (O_1955,N_24028,N_24033);
and UO_1956 (O_1956,N_24208,N_24921);
or UO_1957 (O_1957,N_24565,N_24643);
xor UO_1958 (O_1958,N_24655,N_24650);
and UO_1959 (O_1959,N_24868,N_24651);
nand UO_1960 (O_1960,N_24807,N_24953);
nand UO_1961 (O_1961,N_24341,N_24612);
and UO_1962 (O_1962,N_24579,N_24896);
nand UO_1963 (O_1963,N_24662,N_24071);
or UO_1964 (O_1964,N_24345,N_24377);
nor UO_1965 (O_1965,N_24633,N_24513);
xor UO_1966 (O_1966,N_24398,N_24170);
and UO_1967 (O_1967,N_24471,N_24730);
xor UO_1968 (O_1968,N_24374,N_24056);
xnor UO_1969 (O_1969,N_24038,N_24569);
xor UO_1970 (O_1970,N_24963,N_24917);
nor UO_1971 (O_1971,N_24871,N_24164);
nand UO_1972 (O_1972,N_24177,N_24519);
nor UO_1973 (O_1973,N_24487,N_24333);
or UO_1974 (O_1974,N_24372,N_24339);
nor UO_1975 (O_1975,N_24268,N_24304);
xnor UO_1976 (O_1976,N_24926,N_24476);
or UO_1977 (O_1977,N_24507,N_24760);
xnor UO_1978 (O_1978,N_24697,N_24685);
and UO_1979 (O_1979,N_24417,N_24703);
nor UO_1980 (O_1980,N_24736,N_24490);
and UO_1981 (O_1981,N_24993,N_24165);
nand UO_1982 (O_1982,N_24104,N_24718);
nor UO_1983 (O_1983,N_24430,N_24233);
xor UO_1984 (O_1984,N_24632,N_24715);
nor UO_1985 (O_1985,N_24050,N_24870);
nand UO_1986 (O_1986,N_24981,N_24291);
nor UO_1987 (O_1987,N_24681,N_24497);
and UO_1988 (O_1988,N_24226,N_24424);
or UO_1989 (O_1989,N_24688,N_24860);
xor UO_1990 (O_1990,N_24031,N_24491);
nand UO_1991 (O_1991,N_24866,N_24417);
or UO_1992 (O_1992,N_24300,N_24411);
and UO_1993 (O_1993,N_24051,N_24803);
and UO_1994 (O_1994,N_24924,N_24714);
xnor UO_1995 (O_1995,N_24976,N_24683);
nor UO_1996 (O_1996,N_24319,N_24434);
nand UO_1997 (O_1997,N_24165,N_24971);
nand UO_1998 (O_1998,N_24891,N_24684);
xor UO_1999 (O_1999,N_24544,N_24341);
nor UO_2000 (O_2000,N_24813,N_24599);
nor UO_2001 (O_2001,N_24696,N_24416);
and UO_2002 (O_2002,N_24947,N_24146);
and UO_2003 (O_2003,N_24231,N_24946);
or UO_2004 (O_2004,N_24801,N_24945);
or UO_2005 (O_2005,N_24199,N_24651);
nor UO_2006 (O_2006,N_24403,N_24632);
xor UO_2007 (O_2007,N_24998,N_24231);
xor UO_2008 (O_2008,N_24574,N_24041);
or UO_2009 (O_2009,N_24433,N_24233);
or UO_2010 (O_2010,N_24021,N_24596);
nand UO_2011 (O_2011,N_24955,N_24948);
or UO_2012 (O_2012,N_24398,N_24295);
nor UO_2013 (O_2013,N_24761,N_24940);
or UO_2014 (O_2014,N_24995,N_24422);
and UO_2015 (O_2015,N_24859,N_24942);
or UO_2016 (O_2016,N_24170,N_24489);
xnor UO_2017 (O_2017,N_24101,N_24434);
nor UO_2018 (O_2018,N_24241,N_24796);
nor UO_2019 (O_2019,N_24388,N_24820);
nand UO_2020 (O_2020,N_24649,N_24927);
nor UO_2021 (O_2021,N_24038,N_24948);
or UO_2022 (O_2022,N_24851,N_24295);
xnor UO_2023 (O_2023,N_24474,N_24217);
or UO_2024 (O_2024,N_24981,N_24310);
nor UO_2025 (O_2025,N_24531,N_24362);
or UO_2026 (O_2026,N_24675,N_24735);
and UO_2027 (O_2027,N_24832,N_24051);
xor UO_2028 (O_2028,N_24686,N_24963);
or UO_2029 (O_2029,N_24482,N_24441);
nor UO_2030 (O_2030,N_24388,N_24947);
nor UO_2031 (O_2031,N_24582,N_24071);
nor UO_2032 (O_2032,N_24674,N_24203);
nand UO_2033 (O_2033,N_24042,N_24932);
xor UO_2034 (O_2034,N_24415,N_24998);
xor UO_2035 (O_2035,N_24510,N_24531);
nand UO_2036 (O_2036,N_24762,N_24468);
or UO_2037 (O_2037,N_24992,N_24604);
nand UO_2038 (O_2038,N_24884,N_24886);
or UO_2039 (O_2039,N_24153,N_24060);
and UO_2040 (O_2040,N_24709,N_24001);
or UO_2041 (O_2041,N_24560,N_24724);
and UO_2042 (O_2042,N_24350,N_24358);
nand UO_2043 (O_2043,N_24238,N_24152);
nor UO_2044 (O_2044,N_24204,N_24687);
and UO_2045 (O_2045,N_24415,N_24350);
xnor UO_2046 (O_2046,N_24220,N_24752);
xor UO_2047 (O_2047,N_24026,N_24220);
and UO_2048 (O_2048,N_24268,N_24804);
or UO_2049 (O_2049,N_24952,N_24970);
nand UO_2050 (O_2050,N_24729,N_24014);
nand UO_2051 (O_2051,N_24274,N_24989);
nand UO_2052 (O_2052,N_24088,N_24775);
and UO_2053 (O_2053,N_24823,N_24128);
and UO_2054 (O_2054,N_24239,N_24648);
nand UO_2055 (O_2055,N_24339,N_24253);
nand UO_2056 (O_2056,N_24003,N_24870);
xnor UO_2057 (O_2057,N_24221,N_24224);
or UO_2058 (O_2058,N_24294,N_24155);
xor UO_2059 (O_2059,N_24342,N_24394);
or UO_2060 (O_2060,N_24856,N_24376);
xor UO_2061 (O_2061,N_24497,N_24896);
nor UO_2062 (O_2062,N_24242,N_24751);
and UO_2063 (O_2063,N_24050,N_24809);
nand UO_2064 (O_2064,N_24156,N_24836);
or UO_2065 (O_2065,N_24390,N_24138);
and UO_2066 (O_2066,N_24550,N_24969);
or UO_2067 (O_2067,N_24293,N_24897);
nand UO_2068 (O_2068,N_24608,N_24520);
nor UO_2069 (O_2069,N_24353,N_24087);
or UO_2070 (O_2070,N_24906,N_24053);
nand UO_2071 (O_2071,N_24853,N_24609);
and UO_2072 (O_2072,N_24613,N_24786);
or UO_2073 (O_2073,N_24606,N_24746);
or UO_2074 (O_2074,N_24342,N_24694);
and UO_2075 (O_2075,N_24552,N_24043);
and UO_2076 (O_2076,N_24106,N_24167);
or UO_2077 (O_2077,N_24703,N_24186);
nor UO_2078 (O_2078,N_24960,N_24799);
nand UO_2079 (O_2079,N_24698,N_24226);
and UO_2080 (O_2080,N_24278,N_24731);
nor UO_2081 (O_2081,N_24988,N_24188);
nor UO_2082 (O_2082,N_24847,N_24180);
xnor UO_2083 (O_2083,N_24750,N_24948);
nor UO_2084 (O_2084,N_24059,N_24142);
nor UO_2085 (O_2085,N_24722,N_24756);
xor UO_2086 (O_2086,N_24113,N_24180);
xor UO_2087 (O_2087,N_24905,N_24128);
xor UO_2088 (O_2088,N_24865,N_24185);
nand UO_2089 (O_2089,N_24693,N_24754);
and UO_2090 (O_2090,N_24564,N_24014);
and UO_2091 (O_2091,N_24147,N_24349);
nand UO_2092 (O_2092,N_24307,N_24455);
and UO_2093 (O_2093,N_24438,N_24982);
or UO_2094 (O_2094,N_24372,N_24412);
xor UO_2095 (O_2095,N_24773,N_24260);
xor UO_2096 (O_2096,N_24904,N_24134);
and UO_2097 (O_2097,N_24918,N_24726);
nand UO_2098 (O_2098,N_24342,N_24476);
or UO_2099 (O_2099,N_24575,N_24873);
or UO_2100 (O_2100,N_24119,N_24149);
nand UO_2101 (O_2101,N_24207,N_24339);
xor UO_2102 (O_2102,N_24842,N_24585);
xnor UO_2103 (O_2103,N_24920,N_24915);
xor UO_2104 (O_2104,N_24700,N_24921);
or UO_2105 (O_2105,N_24783,N_24895);
or UO_2106 (O_2106,N_24422,N_24395);
and UO_2107 (O_2107,N_24128,N_24507);
nand UO_2108 (O_2108,N_24529,N_24431);
nand UO_2109 (O_2109,N_24045,N_24864);
or UO_2110 (O_2110,N_24491,N_24922);
or UO_2111 (O_2111,N_24347,N_24784);
nor UO_2112 (O_2112,N_24331,N_24291);
xnor UO_2113 (O_2113,N_24298,N_24212);
or UO_2114 (O_2114,N_24143,N_24120);
or UO_2115 (O_2115,N_24523,N_24011);
and UO_2116 (O_2116,N_24169,N_24116);
or UO_2117 (O_2117,N_24211,N_24958);
nor UO_2118 (O_2118,N_24628,N_24351);
or UO_2119 (O_2119,N_24610,N_24236);
or UO_2120 (O_2120,N_24324,N_24319);
and UO_2121 (O_2121,N_24114,N_24684);
nand UO_2122 (O_2122,N_24674,N_24309);
nand UO_2123 (O_2123,N_24714,N_24347);
nor UO_2124 (O_2124,N_24474,N_24184);
xor UO_2125 (O_2125,N_24086,N_24623);
nand UO_2126 (O_2126,N_24905,N_24014);
and UO_2127 (O_2127,N_24682,N_24573);
and UO_2128 (O_2128,N_24899,N_24659);
nor UO_2129 (O_2129,N_24188,N_24861);
and UO_2130 (O_2130,N_24795,N_24655);
xnor UO_2131 (O_2131,N_24391,N_24012);
xnor UO_2132 (O_2132,N_24651,N_24072);
or UO_2133 (O_2133,N_24899,N_24553);
or UO_2134 (O_2134,N_24424,N_24504);
nor UO_2135 (O_2135,N_24132,N_24842);
or UO_2136 (O_2136,N_24509,N_24270);
or UO_2137 (O_2137,N_24040,N_24670);
xor UO_2138 (O_2138,N_24272,N_24724);
or UO_2139 (O_2139,N_24790,N_24779);
xnor UO_2140 (O_2140,N_24334,N_24816);
xor UO_2141 (O_2141,N_24528,N_24262);
nor UO_2142 (O_2142,N_24417,N_24526);
xnor UO_2143 (O_2143,N_24269,N_24020);
or UO_2144 (O_2144,N_24158,N_24869);
and UO_2145 (O_2145,N_24663,N_24428);
xor UO_2146 (O_2146,N_24454,N_24055);
or UO_2147 (O_2147,N_24775,N_24593);
nand UO_2148 (O_2148,N_24364,N_24543);
nor UO_2149 (O_2149,N_24531,N_24352);
nor UO_2150 (O_2150,N_24801,N_24606);
or UO_2151 (O_2151,N_24624,N_24898);
xor UO_2152 (O_2152,N_24323,N_24825);
xor UO_2153 (O_2153,N_24408,N_24249);
and UO_2154 (O_2154,N_24283,N_24568);
nand UO_2155 (O_2155,N_24600,N_24765);
or UO_2156 (O_2156,N_24898,N_24095);
xor UO_2157 (O_2157,N_24987,N_24447);
or UO_2158 (O_2158,N_24695,N_24520);
or UO_2159 (O_2159,N_24291,N_24522);
and UO_2160 (O_2160,N_24543,N_24111);
or UO_2161 (O_2161,N_24697,N_24885);
nor UO_2162 (O_2162,N_24717,N_24257);
xor UO_2163 (O_2163,N_24904,N_24587);
and UO_2164 (O_2164,N_24276,N_24027);
or UO_2165 (O_2165,N_24159,N_24973);
or UO_2166 (O_2166,N_24214,N_24129);
xor UO_2167 (O_2167,N_24615,N_24218);
and UO_2168 (O_2168,N_24962,N_24605);
or UO_2169 (O_2169,N_24084,N_24990);
or UO_2170 (O_2170,N_24580,N_24087);
or UO_2171 (O_2171,N_24134,N_24049);
nor UO_2172 (O_2172,N_24455,N_24374);
nor UO_2173 (O_2173,N_24102,N_24249);
xnor UO_2174 (O_2174,N_24628,N_24372);
or UO_2175 (O_2175,N_24209,N_24617);
nand UO_2176 (O_2176,N_24139,N_24035);
or UO_2177 (O_2177,N_24167,N_24706);
nor UO_2178 (O_2178,N_24964,N_24305);
nor UO_2179 (O_2179,N_24152,N_24251);
or UO_2180 (O_2180,N_24276,N_24653);
nor UO_2181 (O_2181,N_24788,N_24189);
xnor UO_2182 (O_2182,N_24222,N_24735);
nor UO_2183 (O_2183,N_24155,N_24914);
or UO_2184 (O_2184,N_24147,N_24069);
and UO_2185 (O_2185,N_24267,N_24456);
nor UO_2186 (O_2186,N_24033,N_24763);
or UO_2187 (O_2187,N_24349,N_24667);
nand UO_2188 (O_2188,N_24521,N_24864);
xnor UO_2189 (O_2189,N_24832,N_24596);
nand UO_2190 (O_2190,N_24255,N_24957);
nand UO_2191 (O_2191,N_24219,N_24986);
or UO_2192 (O_2192,N_24520,N_24255);
xor UO_2193 (O_2193,N_24926,N_24486);
xor UO_2194 (O_2194,N_24249,N_24824);
and UO_2195 (O_2195,N_24656,N_24716);
nand UO_2196 (O_2196,N_24871,N_24826);
nor UO_2197 (O_2197,N_24814,N_24992);
and UO_2198 (O_2198,N_24803,N_24285);
nand UO_2199 (O_2199,N_24331,N_24449);
nor UO_2200 (O_2200,N_24419,N_24694);
nor UO_2201 (O_2201,N_24298,N_24928);
and UO_2202 (O_2202,N_24213,N_24758);
or UO_2203 (O_2203,N_24484,N_24159);
xor UO_2204 (O_2204,N_24718,N_24232);
or UO_2205 (O_2205,N_24533,N_24689);
nand UO_2206 (O_2206,N_24204,N_24214);
and UO_2207 (O_2207,N_24543,N_24403);
nor UO_2208 (O_2208,N_24373,N_24950);
or UO_2209 (O_2209,N_24944,N_24984);
or UO_2210 (O_2210,N_24862,N_24972);
nor UO_2211 (O_2211,N_24490,N_24006);
xor UO_2212 (O_2212,N_24838,N_24742);
xnor UO_2213 (O_2213,N_24780,N_24790);
or UO_2214 (O_2214,N_24364,N_24704);
nor UO_2215 (O_2215,N_24774,N_24668);
nor UO_2216 (O_2216,N_24271,N_24490);
or UO_2217 (O_2217,N_24266,N_24088);
or UO_2218 (O_2218,N_24683,N_24481);
xnor UO_2219 (O_2219,N_24359,N_24228);
and UO_2220 (O_2220,N_24931,N_24496);
nor UO_2221 (O_2221,N_24862,N_24189);
or UO_2222 (O_2222,N_24251,N_24580);
or UO_2223 (O_2223,N_24670,N_24606);
xor UO_2224 (O_2224,N_24452,N_24233);
and UO_2225 (O_2225,N_24388,N_24624);
or UO_2226 (O_2226,N_24914,N_24799);
nand UO_2227 (O_2227,N_24879,N_24901);
and UO_2228 (O_2228,N_24626,N_24038);
nor UO_2229 (O_2229,N_24386,N_24983);
nand UO_2230 (O_2230,N_24189,N_24314);
and UO_2231 (O_2231,N_24590,N_24008);
or UO_2232 (O_2232,N_24598,N_24037);
xnor UO_2233 (O_2233,N_24325,N_24879);
or UO_2234 (O_2234,N_24715,N_24254);
and UO_2235 (O_2235,N_24444,N_24892);
or UO_2236 (O_2236,N_24780,N_24252);
nor UO_2237 (O_2237,N_24703,N_24150);
and UO_2238 (O_2238,N_24499,N_24791);
nor UO_2239 (O_2239,N_24249,N_24272);
nand UO_2240 (O_2240,N_24560,N_24630);
xnor UO_2241 (O_2241,N_24718,N_24527);
nand UO_2242 (O_2242,N_24679,N_24693);
nor UO_2243 (O_2243,N_24457,N_24379);
xor UO_2244 (O_2244,N_24450,N_24444);
nand UO_2245 (O_2245,N_24854,N_24282);
nand UO_2246 (O_2246,N_24253,N_24620);
nand UO_2247 (O_2247,N_24964,N_24697);
or UO_2248 (O_2248,N_24889,N_24430);
and UO_2249 (O_2249,N_24748,N_24940);
and UO_2250 (O_2250,N_24483,N_24352);
and UO_2251 (O_2251,N_24615,N_24171);
nand UO_2252 (O_2252,N_24369,N_24268);
nor UO_2253 (O_2253,N_24853,N_24759);
nor UO_2254 (O_2254,N_24819,N_24210);
and UO_2255 (O_2255,N_24709,N_24242);
nand UO_2256 (O_2256,N_24738,N_24650);
and UO_2257 (O_2257,N_24251,N_24517);
xor UO_2258 (O_2258,N_24462,N_24797);
xor UO_2259 (O_2259,N_24247,N_24028);
and UO_2260 (O_2260,N_24559,N_24724);
nand UO_2261 (O_2261,N_24357,N_24246);
and UO_2262 (O_2262,N_24325,N_24392);
nor UO_2263 (O_2263,N_24678,N_24373);
and UO_2264 (O_2264,N_24548,N_24392);
nand UO_2265 (O_2265,N_24222,N_24418);
xnor UO_2266 (O_2266,N_24060,N_24403);
xor UO_2267 (O_2267,N_24474,N_24977);
or UO_2268 (O_2268,N_24224,N_24351);
or UO_2269 (O_2269,N_24586,N_24727);
xor UO_2270 (O_2270,N_24268,N_24742);
xnor UO_2271 (O_2271,N_24970,N_24133);
and UO_2272 (O_2272,N_24336,N_24330);
xor UO_2273 (O_2273,N_24406,N_24459);
nand UO_2274 (O_2274,N_24587,N_24790);
nor UO_2275 (O_2275,N_24748,N_24902);
nor UO_2276 (O_2276,N_24616,N_24941);
or UO_2277 (O_2277,N_24128,N_24317);
or UO_2278 (O_2278,N_24331,N_24661);
nand UO_2279 (O_2279,N_24901,N_24186);
and UO_2280 (O_2280,N_24594,N_24658);
nand UO_2281 (O_2281,N_24189,N_24841);
nand UO_2282 (O_2282,N_24966,N_24156);
nand UO_2283 (O_2283,N_24167,N_24659);
xnor UO_2284 (O_2284,N_24179,N_24438);
nor UO_2285 (O_2285,N_24846,N_24141);
nor UO_2286 (O_2286,N_24709,N_24315);
and UO_2287 (O_2287,N_24671,N_24617);
xor UO_2288 (O_2288,N_24678,N_24618);
and UO_2289 (O_2289,N_24978,N_24626);
nand UO_2290 (O_2290,N_24978,N_24508);
nand UO_2291 (O_2291,N_24662,N_24383);
nand UO_2292 (O_2292,N_24789,N_24853);
xnor UO_2293 (O_2293,N_24845,N_24754);
or UO_2294 (O_2294,N_24099,N_24524);
xnor UO_2295 (O_2295,N_24089,N_24830);
and UO_2296 (O_2296,N_24848,N_24909);
nor UO_2297 (O_2297,N_24610,N_24314);
xor UO_2298 (O_2298,N_24414,N_24521);
or UO_2299 (O_2299,N_24365,N_24799);
xnor UO_2300 (O_2300,N_24431,N_24227);
or UO_2301 (O_2301,N_24764,N_24382);
and UO_2302 (O_2302,N_24462,N_24863);
or UO_2303 (O_2303,N_24357,N_24927);
xor UO_2304 (O_2304,N_24810,N_24598);
xor UO_2305 (O_2305,N_24438,N_24543);
and UO_2306 (O_2306,N_24102,N_24168);
nor UO_2307 (O_2307,N_24060,N_24430);
nand UO_2308 (O_2308,N_24858,N_24209);
nand UO_2309 (O_2309,N_24342,N_24175);
xor UO_2310 (O_2310,N_24008,N_24329);
or UO_2311 (O_2311,N_24506,N_24479);
nand UO_2312 (O_2312,N_24671,N_24670);
xor UO_2313 (O_2313,N_24587,N_24768);
xnor UO_2314 (O_2314,N_24929,N_24552);
and UO_2315 (O_2315,N_24862,N_24113);
nor UO_2316 (O_2316,N_24678,N_24328);
nand UO_2317 (O_2317,N_24097,N_24814);
xor UO_2318 (O_2318,N_24067,N_24901);
or UO_2319 (O_2319,N_24513,N_24312);
nand UO_2320 (O_2320,N_24192,N_24802);
or UO_2321 (O_2321,N_24281,N_24266);
nand UO_2322 (O_2322,N_24519,N_24973);
xor UO_2323 (O_2323,N_24814,N_24613);
xor UO_2324 (O_2324,N_24401,N_24802);
and UO_2325 (O_2325,N_24492,N_24931);
and UO_2326 (O_2326,N_24695,N_24245);
nor UO_2327 (O_2327,N_24482,N_24856);
xor UO_2328 (O_2328,N_24552,N_24760);
xnor UO_2329 (O_2329,N_24012,N_24568);
nor UO_2330 (O_2330,N_24551,N_24927);
xnor UO_2331 (O_2331,N_24288,N_24702);
nand UO_2332 (O_2332,N_24787,N_24488);
or UO_2333 (O_2333,N_24574,N_24937);
nor UO_2334 (O_2334,N_24840,N_24698);
xor UO_2335 (O_2335,N_24038,N_24149);
nor UO_2336 (O_2336,N_24660,N_24776);
xor UO_2337 (O_2337,N_24532,N_24478);
and UO_2338 (O_2338,N_24261,N_24598);
and UO_2339 (O_2339,N_24479,N_24117);
nor UO_2340 (O_2340,N_24687,N_24767);
nor UO_2341 (O_2341,N_24669,N_24589);
nor UO_2342 (O_2342,N_24468,N_24310);
or UO_2343 (O_2343,N_24307,N_24923);
nor UO_2344 (O_2344,N_24857,N_24397);
or UO_2345 (O_2345,N_24894,N_24867);
or UO_2346 (O_2346,N_24299,N_24865);
and UO_2347 (O_2347,N_24526,N_24887);
nand UO_2348 (O_2348,N_24009,N_24333);
or UO_2349 (O_2349,N_24400,N_24461);
xnor UO_2350 (O_2350,N_24406,N_24154);
xor UO_2351 (O_2351,N_24470,N_24945);
nand UO_2352 (O_2352,N_24665,N_24581);
nand UO_2353 (O_2353,N_24938,N_24845);
nor UO_2354 (O_2354,N_24670,N_24124);
nor UO_2355 (O_2355,N_24067,N_24468);
nor UO_2356 (O_2356,N_24048,N_24033);
xnor UO_2357 (O_2357,N_24756,N_24171);
and UO_2358 (O_2358,N_24384,N_24174);
and UO_2359 (O_2359,N_24596,N_24321);
nor UO_2360 (O_2360,N_24699,N_24633);
nor UO_2361 (O_2361,N_24204,N_24613);
or UO_2362 (O_2362,N_24153,N_24672);
and UO_2363 (O_2363,N_24903,N_24097);
and UO_2364 (O_2364,N_24923,N_24527);
or UO_2365 (O_2365,N_24368,N_24456);
nor UO_2366 (O_2366,N_24104,N_24951);
nand UO_2367 (O_2367,N_24847,N_24444);
xor UO_2368 (O_2368,N_24894,N_24086);
or UO_2369 (O_2369,N_24321,N_24815);
xnor UO_2370 (O_2370,N_24101,N_24522);
xor UO_2371 (O_2371,N_24013,N_24685);
or UO_2372 (O_2372,N_24858,N_24304);
xor UO_2373 (O_2373,N_24809,N_24667);
xor UO_2374 (O_2374,N_24305,N_24726);
nor UO_2375 (O_2375,N_24501,N_24302);
or UO_2376 (O_2376,N_24642,N_24286);
or UO_2377 (O_2377,N_24612,N_24669);
and UO_2378 (O_2378,N_24764,N_24743);
nand UO_2379 (O_2379,N_24207,N_24309);
or UO_2380 (O_2380,N_24720,N_24986);
or UO_2381 (O_2381,N_24160,N_24813);
or UO_2382 (O_2382,N_24361,N_24676);
nor UO_2383 (O_2383,N_24990,N_24511);
and UO_2384 (O_2384,N_24439,N_24490);
and UO_2385 (O_2385,N_24403,N_24757);
xnor UO_2386 (O_2386,N_24808,N_24983);
nor UO_2387 (O_2387,N_24257,N_24523);
or UO_2388 (O_2388,N_24136,N_24750);
xor UO_2389 (O_2389,N_24792,N_24158);
nand UO_2390 (O_2390,N_24814,N_24188);
and UO_2391 (O_2391,N_24451,N_24718);
and UO_2392 (O_2392,N_24637,N_24059);
nand UO_2393 (O_2393,N_24066,N_24089);
and UO_2394 (O_2394,N_24513,N_24829);
and UO_2395 (O_2395,N_24838,N_24324);
xor UO_2396 (O_2396,N_24252,N_24535);
xnor UO_2397 (O_2397,N_24382,N_24141);
xor UO_2398 (O_2398,N_24658,N_24473);
xor UO_2399 (O_2399,N_24682,N_24426);
xnor UO_2400 (O_2400,N_24565,N_24107);
nor UO_2401 (O_2401,N_24399,N_24450);
and UO_2402 (O_2402,N_24413,N_24691);
or UO_2403 (O_2403,N_24118,N_24647);
xnor UO_2404 (O_2404,N_24720,N_24601);
or UO_2405 (O_2405,N_24302,N_24872);
xnor UO_2406 (O_2406,N_24292,N_24153);
or UO_2407 (O_2407,N_24342,N_24664);
or UO_2408 (O_2408,N_24763,N_24463);
nor UO_2409 (O_2409,N_24331,N_24780);
xor UO_2410 (O_2410,N_24957,N_24109);
and UO_2411 (O_2411,N_24327,N_24146);
nor UO_2412 (O_2412,N_24171,N_24914);
and UO_2413 (O_2413,N_24616,N_24191);
or UO_2414 (O_2414,N_24228,N_24789);
or UO_2415 (O_2415,N_24761,N_24496);
nand UO_2416 (O_2416,N_24175,N_24430);
and UO_2417 (O_2417,N_24166,N_24637);
nand UO_2418 (O_2418,N_24742,N_24847);
nor UO_2419 (O_2419,N_24350,N_24411);
nand UO_2420 (O_2420,N_24503,N_24665);
nor UO_2421 (O_2421,N_24324,N_24014);
or UO_2422 (O_2422,N_24525,N_24407);
xnor UO_2423 (O_2423,N_24958,N_24994);
nor UO_2424 (O_2424,N_24729,N_24454);
nand UO_2425 (O_2425,N_24035,N_24573);
nor UO_2426 (O_2426,N_24229,N_24027);
and UO_2427 (O_2427,N_24574,N_24675);
and UO_2428 (O_2428,N_24184,N_24698);
nand UO_2429 (O_2429,N_24856,N_24617);
nand UO_2430 (O_2430,N_24969,N_24436);
and UO_2431 (O_2431,N_24045,N_24156);
nor UO_2432 (O_2432,N_24112,N_24044);
xnor UO_2433 (O_2433,N_24581,N_24633);
nand UO_2434 (O_2434,N_24356,N_24697);
and UO_2435 (O_2435,N_24808,N_24393);
or UO_2436 (O_2436,N_24668,N_24475);
nor UO_2437 (O_2437,N_24517,N_24666);
nor UO_2438 (O_2438,N_24088,N_24953);
nor UO_2439 (O_2439,N_24345,N_24331);
or UO_2440 (O_2440,N_24559,N_24117);
xnor UO_2441 (O_2441,N_24117,N_24464);
xor UO_2442 (O_2442,N_24489,N_24909);
nor UO_2443 (O_2443,N_24830,N_24665);
nor UO_2444 (O_2444,N_24218,N_24702);
or UO_2445 (O_2445,N_24197,N_24800);
nor UO_2446 (O_2446,N_24488,N_24241);
and UO_2447 (O_2447,N_24783,N_24616);
or UO_2448 (O_2448,N_24575,N_24339);
xnor UO_2449 (O_2449,N_24272,N_24545);
or UO_2450 (O_2450,N_24833,N_24667);
xor UO_2451 (O_2451,N_24734,N_24807);
nor UO_2452 (O_2452,N_24562,N_24152);
xor UO_2453 (O_2453,N_24952,N_24448);
nand UO_2454 (O_2454,N_24389,N_24140);
or UO_2455 (O_2455,N_24703,N_24012);
and UO_2456 (O_2456,N_24484,N_24619);
nand UO_2457 (O_2457,N_24197,N_24581);
nor UO_2458 (O_2458,N_24834,N_24500);
and UO_2459 (O_2459,N_24282,N_24707);
xnor UO_2460 (O_2460,N_24330,N_24215);
or UO_2461 (O_2461,N_24599,N_24937);
or UO_2462 (O_2462,N_24771,N_24927);
and UO_2463 (O_2463,N_24179,N_24196);
nor UO_2464 (O_2464,N_24265,N_24776);
nor UO_2465 (O_2465,N_24038,N_24061);
nand UO_2466 (O_2466,N_24200,N_24806);
or UO_2467 (O_2467,N_24077,N_24321);
xnor UO_2468 (O_2468,N_24031,N_24569);
nor UO_2469 (O_2469,N_24387,N_24333);
nand UO_2470 (O_2470,N_24292,N_24272);
and UO_2471 (O_2471,N_24861,N_24418);
nor UO_2472 (O_2472,N_24370,N_24369);
and UO_2473 (O_2473,N_24394,N_24176);
nor UO_2474 (O_2474,N_24692,N_24313);
xor UO_2475 (O_2475,N_24142,N_24737);
nand UO_2476 (O_2476,N_24627,N_24363);
nor UO_2477 (O_2477,N_24092,N_24061);
nor UO_2478 (O_2478,N_24744,N_24201);
xor UO_2479 (O_2479,N_24440,N_24018);
or UO_2480 (O_2480,N_24700,N_24015);
nand UO_2481 (O_2481,N_24727,N_24755);
nand UO_2482 (O_2482,N_24866,N_24199);
and UO_2483 (O_2483,N_24710,N_24982);
and UO_2484 (O_2484,N_24702,N_24464);
nor UO_2485 (O_2485,N_24392,N_24365);
xnor UO_2486 (O_2486,N_24570,N_24567);
and UO_2487 (O_2487,N_24720,N_24052);
and UO_2488 (O_2488,N_24358,N_24409);
xor UO_2489 (O_2489,N_24941,N_24598);
xor UO_2490 (O_2490,N_24980,N_24696);
nand UO_2491 (O_2491,N_24452,N_24221);
nand UO_2492 (O_2492,N_24418,N_24608);
nor UO_2493 (O_2493,N_24051,N_24174);
and UO_2494 (O_2494,N_24087,N_24564);
nand UO_2495 (O_2495,N_24103,N_24916);
and UO_2496 (O_2496,N_24159,N_24988);
xor UO_2497 (O_2497,N_24604,N_24787);
and UO_2498 (O_2498,N_24899,N_24651);
and UO_2499 (O_2499,N_24509,N_24285);
nor UO_2500 (O_2500,N_24633,N_24784);
nor UO_2501 (O_2501,N_24201,N_24144);
nand UO_2502 (O_2502,N_24950,N_24687);
or UO_2503 (O_2503,N_24698,N_24492);
and UO_2504 (O_2504,N_24045,N_24240);
xor UO_2505 (O_2505,N_24617,N_24817);
nor UO_2506 (O_2506,N_24187,N_24521);
or UO_2507 (O_2507,N_24322,N_24121);
nand UO_2508 (O_2508,N_24471,N_24057);
or UO_2509 (O_2509,N_24147,N_24960);
and UO_2510 (O_2510,N_24680,N_24455);
nor UO_2511 (O_2511,N_24564,N_24318);
and UO_2512 (O_2512,N_24504,N_24147);
nor UO_2513 (O_2513,N_24605,N_24507);
xnor UO_2514 (O_2514,N_24216,N_24840);
xor UO_2515 (O_2515,N_24989,N_24251);
nand UO_2516 (O_2516,N_24233,N_24519);
nand UO_2517 (O_2517,N_24187,N_24235);
or UO_2518 (O_2518,N_24338,N_24276);
or UO_2519 (O_2519,N_24943,N_24453);
or UO_2520 (O_2520,N_24286,N_24731);
or UO_2521 (O_2521,N_24794,N_24426);
or UO_2522 (O_2522,N_24385,N_24484);
nor UO_2523 (O_2523,N_24326,N_24470);
nor UO_2524 (O_2524,N_24010,N_24659);
and UO_2525 (O_2525,N_24362,N_24991);
xnor UO_2526 (O_2526,N_24722,N_24733);
nor UO_2527 (O_2527,N_24127,N_24742);
xnor UO_2528 (O_2528,N_24143,N_24655);
or UO_2529 (O_2529,N_24850,N_24949);
or UO_2530 (O_2530,N_24200,N_24534);
nor UO_2531 (O_2531,N_24408,N_24255);
or UO_2532 (O_2532,N_24938,N_24747);
xor UO_2533 (O_2533,N_24427,N_24069);
nor UO_2534 (O_2534,N_24335,N_24829);
nor UO_2535 (O_2535,N_24482,N_24233);
nand UO_2536 (O_2536,N_24869,N_24663);
nand UO_2537 (O_2537,N_24131,N_24355);
nand UO_2538 (O_2538,N_24080,N_24904);
nand UO_2539 (O_2539,N_24650,N_24505);
and UO_2540 (O_2540,N_24985,N_24584);
nor UO_2541 (O_2541,N_24377,N_24491);
xnor UO_2542 (O_2542,N_24537,N_24717);
and UO_2543 (O_2543,N_24034,N_24576);
and UO_2544 (O_2544,N_24260,N_24051);
nor UO_2545 (O_2545,N_24794,N_24513);
nand UO_2546 (O_2546,N_24975,N_24080);
nand UO_2547 (O_2547,N_24148,N_24050);
nor UO_2548 (O_2548,N_24719,N_24763);
nor UO_2549 (O_2549,N_24073,N_24580);
xnor UO_2550 (O_2550,N_24776,N_24731);
or UO_2551 (O_2551,N_24019,N_24607);
nand UO_2552 (O_2552,N_24563,N_24026);
xor UO_2553 (O_2553,N_24893,N_24890);
or UO_2554 (O_2554,N_24764,N_24379);
nand UO_2555 (O_2555,N_24489,N_24215);
nor UO_2556 (O_2556,N_24621,N_24306);
or UO_2557 (O_2557,N_24710,N_24649);
xor UO_2558 (O_2558,N_24011,N_24178);
or UO_2559 (O_2559,N_24858,N_24519);
xor UO_2560 (O_2560,N_24270,N_24027);
nand UO_2561 (O_2561,N_24231,N_24424);
nor UO_2562 (O_2562,N_24926,N_24739);
and UO_2563 (O_2563,N_24518,N_24130);
and UO_2564 (O_2564,N_24833,N_24478);
xnor UO_2565 (O_2565,N_24822,N_24439);
or UO_2566 (O_2566,N_24448,N_24718);
xor UO_2567 (O_2567,N_24164,N_24808);
nor UO_2568 (O_2568,N_24357,N_24844);
nand UO_2569 (O_2569,N_24483,N_24562);
nand UO_2570 (O_2570,N_24003,N_24908);
or UO_2571 (O_2571,N_24616,N_24093);
xnor UO_2572 (O_2572,N_24615,N_24629);
nor UO_2573 (O_2573,N_24295,N_24687);
or UO_2574 (O_2574,N_24650,N_24495);
xnor UO_2575 (O_2575,N_24907,N_24145);
nor UO_2576 (O_2576,N_24486,N_24804);
and UO_2577 (O_2577,N_24971,N_24086);
or UO_2578 (O_2578,N_24210,N_24447);
xnor UO_2579 (O_2579,N_24541,N_24610);
nor UO_2580 (O_2580,N_24900,N_24176);
and UO_2581 (O_2581,N_24178,N_24330);
nor UO_2582 (O_2582,N_24773,N_24793);
nand UO_2583 (O_2583,N_24135,N_24171);
xor UO_2584 (O_2584,N_24263,N_24482);
nor UO_2585 (O_2585,N_24353,N_24685);
nand UO_2586 (O_2586,N_24590,N_24554);
and UO_2587 (O_2587,N_24345,N_24880);
nor UO_2588 (O_2588,N_24647,N_24826);
or UO_2589 (O_2589,N_24437,N_24418);
and UO_2590 (O_2590,N_24737,N_24424);
nand UO_2591 (O_2591,N_24825,N_24436);
xnor UO_2592 (O_2592,N_24810,N_24924);
nor UO_2593 (O_2593,N_24770,N_24221);
nand UO_2594 (O_2594,N_24910,N_24547);
nor UO_2595 (O_2595,N_24149,N_24267);
nor UO_2596 (O_2596,N_24918,N_24666);
nor UO_2597 (O_2597,N_24919,N_24350);
xor UO_2598 (O_2598,N_24883,N_24326);
and UO_2599 (O_2599,N_24228,N_24824);
xor UO_2600 (O_2600,N_24785,N_24714);
or UO_2601 (O_2601,N_24835,N_24183);
or UO_2602 (O_2602,N_24864,N_24944);
or UO_2603 (O_2603,N_24750,N_24240);
or UO_2604 (O_2604,N_24915,N_24782);
and UO_2605 (O_2605,N_24428,N_24297);
nand UO_2606 (O_2606,N_24882,N_24252);
or UO_2607 (O_2607,N_24505,N_24598);
nand UO_2608 (O_2608,N_24274,N_24714);
xor UO_2609 (O_2609,N_24533,N_24537);
or UO_2610 (O_2610,N_24152,N_24107);
and UO_2611 (O_2611,N_24585,N_24352);
and UO_2612 (O_2612,N_24873,N_24188);
nor UO_2613 (O_2613,N_24672,N_24864);
nand UO_2614 (O_2614,N_24919,N_24238);
nand UO_2615 (O_2615,N_24851,N_24536);
nand UO_2616 (O_2616,N_24603,N_24203);
nand UO_2617 (O_2617,N_24062,N_24886);
or UO_2618 (O_2618,N_24804,N_24015);
nor UO_2619 (O_2619,N_24920,N_24583);
nor UO_2620 (O_2620,N_24941,N_24470);
xnor UO_2621 (O_2621,N_24131,N_24115);
or UO_2622 (O_2622,N_24302,N_24062);
nor UO_2623 (O_2623,N_24685,N_24875);
xnor UO_2624 (O_2624,N_24791,N_24521);
xnor UO_2625 (O_2625,N_24649,N_24376);
or UO_2626 (O_2626,N_24844,N_24354);
or UO_2627 (O_2627,N_24217,N_24762);
and UO_2628 (O_2628,N_24889,N_24687);
nand UO_2629 (O_2629,N_24331,N_24380);
and UO_2630 (O_2630,N_24005,N_24077);
nand UO_2631 (O_2631,N_24770,N_24866);
and UO_2632 (O_2632,N_24572,N_24436);
or UO_2633 (O_2633,N_24119,N_24784);
and UO_2634 (O_2634,N_24084,N_24241);
nand UO_2635 (O_2635,N_24021,N_24097);
and UO_2636 (O_2636,N_24657,N_24606);
and UO_2637 (O_2637,N_24083,N_24026);
nand UO_2638 (O_2638,N_24005,N_24183);
xor UO_2639 (O_2639,N_24963,N_24753);
nand UO_2640 (O_2640,N_24763,N_24263);
nor UO_2641 (O_2641,N_24783,N_24096);
and UO_2642 (O_2642,N_24911,N_24715);
nor UO_2643 (O_2643,N_24955,N_24413);
and UO_2644 (O_2644,N_24907,N_24874);
xor UO_2645 (O_2645,N_24832,N_24358);
xor UO_2646 (O_2646,N_24260,N_24603);
and UO_2647 (O_2647,N_24427,N_24060);
or UO_2648 (O_2648,N_24942,N_24957);
nor UO_2649 (O_2649,N_24690,N_24659);
xnor UO_2650 (O_2650,N_24185,N_24631);
nand UO_2651 (O_2651,N_24797,N_24770);
and UO_2652 (O_2652,N_24472,N_24835);
nor UO_2653 (O_2653,N_24943,N_24948);
nand UO_2654 (O_2654,N_24139,N_24656);
or UO_2655 (O_2655,N_24018,N_24690);
or UO_2656 (O_2656,N_24904,N_24314);
xnor UO_2657 (O_2657,N_24399,N_24575);
xor UO_2658 (O_2658,N_24936,N_24444);
xor UO_2659 (O_2659,N_24878,N_24200);
nand UO_2660 (O_2660,N_24111,N_24260);
or UO_2661 (O_2661,N_24326,N_24142);
and UO_2662 (O_2662,N_24261,N_24877);
nor UO_2663 (O_2663,N_24094,N_24486);
or UO_2664 (O_2664,N_24866,N_24235);
nor UO_2665 (O_2665,N_24325,N_24447);
and UO_2666 (O_2666,N_24576,N_24613);
or UO_2667 (O_2667,N_24440,N_24311);
and UO_2668 (O_2668,N_24763,N_24156);
nor UO_2669 (O_2669,N_24999,N_24783);
or UO_2670 (O_2670,N_24648,N_24604);
xor UO_2671 (O_2671,N_24695,N_24319);
xnor UO_2672 (O_2672,N_24176,N_24072);
and UO_2673 (O_2673,N_24194,N_24006);
nor UO_2674 (O_2674,N_24750,N_24841);
nor UO_2675 (O_2675,N_24251,N_24312);
xnor UO_2676 (O_2676,N_24567,N_24988);
nand UO_2677 (O_2677,N_24196,N_24697);
nand UO_2678 (O_2678,N_24151,N_24387);
xnor UO_2679 (O_2679,N_24698,N_24543);
nand UO_2680 (O_2680,N_24944,N_24950);
and UO_2681 (O_2681,N_24620,N_24076);
nand UO_2682 (O_2682,N_24672,N_24148);
nand UO_2683 (O_2683,N_24631,N_24512);
nand UO_2684 (O_2684,N_24887,N_24934);
nor UO_2685 (O_2685,N_24517,N_24646);
nand UO_2686 (O_2686,N_24003,N_24578);
nor UO_2687 (O_2687,N_24624,N_24317);
and UO_2688 (O_2688,N_24979,N_24315);
nand UO_2689 (O_2689,N_24388,N_24434);
nor UO_2690 (O_2690,N_24791,N_24836);
xor UO_2691 (O_2691,N_24295,N_24633);
nand UO_2692 (O_2692,N_24049,N_24990);
xnor UO_2693 (O_2693,N_24588,N_24539);
nor UO_2694 (O_2694,N_24182,N_24461);
nor UO_2695 (O_2695,N_24225,N_24125);
nand UO_2696 (O_2696,N_24245,N_24041);
xnor UO_2697 (O_2697,N_24815,N_24149);
or UO_2698 (O_2698,N_24984,N_24305);
xnor UO_2699 (O_2699,N_24770,N_24485);
and UO_2700 (O_2700,N_24723,N_24902);
nor UO_2701 (O_2701,N_24316,N_24015);
and UO_2702 (O_2702,N_24705,N_24861);
or UO_2703 (O_2703,N_24186,N_24884);
and UO_2704 (O_2704,N_24257,N_24800);
xnor UO_2705 (O_2705,N_24255,N_24063);
nor UO_2706 (O_2706,N_24603,N_24966);
xor UO_2707 (O_2707,N_24644,N_24788);
and UO_2708 (O_2708,N_24114,N_24650);
xnor UO_2709 (O_2709,N_24867,N_24804);
and UO_2710 (O_2710,N_24908,N_24989);
or UO_2711 (O_2711,N_24488,N_24999);
nand UO_2712 (O_2712,N_24474,N_24279);
xor UO_2713 (O_2713,N_24110,N_24030);
xnor UO_2714 (O_2714,N_24450,N_24436);
and UO_2715 (O_2715,N_24076,N_24401);
xor UO_2716 (O_2716,N_24614,N_24837);
nand UO_2717 (O_2717,N_24808,N_24444);
nor UO_2718 (O_2718,N_24607,N_24519);
nor UO_2719 (O_2719,N_24019,N_24470);
or UO_2720 (O_2720,N_24850,N_24769);
xnor UO_2721 (O_2721,N_24245,N_24276);
nand UO_2722 (O_2722,N_24997,N_24534);
nor UO_2723 (O_2723,N_24665,N_24002);
nand UO_2724 (O_2724,N_24519,N_24461);
and UO_2725 (O_2725,N_24965,N_24940);
nand UO_2726 (O_2726,N_24388,N_24464);
nor UO_2727 (O_2727,N_24792,N_24349);
and UO_2728 (O_2728,N_24971,N_24873);
and UO_2729 (O_2729,N_24429,N_24981);
and UO_2730 (O_2730,N_24429,N_24421);
nand UO_2731 (O_2731,N_24554,N_24476);
or UO_2732 (O_2732,N_24944,N_24849);
or UO_2733 (O_2733,N_24531,N_24989);
or UO_2734 (O_2734,N_24845,N_24212);
xnor UO_2735 (O_2735,N_24861,N_24507);
and UO_2736 (O_2736,N_24723,N_24796);
nand UO_2737 (O_2737,N_24823,N_24626);
or UO_2738 (O_2738,N_24351,N_24391);
xor UO_2739 (O_2739,N_24955,N_24501);
and UO_2740 (O_2740,N_24349,N_24178);
or UO_2741 (O_2741,N_24645,N_24382);
nor UO_2742 (O_2742,N_24944,N_24946);
nand UO_2743 (O_2743,N_24751,N_24722);
nor UO_2744 (O_2744,N_24913,N_24536);
nor UO_2745 (O_2745,N_24482,N_24497);
nand UO_2746 (O_2746,N_24873,N_24913);
nand UO_2747 (O_2747,N_24337,N_24457);
or UO_2748 (O_2748,N_24519,N_24065);
nor UO_2749 (O_2749,N_24152,N_24278);
nor UO_2750 (O_2750,N_24549,N_24564);
xnor UO_2751 (O_2751,N_24280,N_24624);
and UO_2752 (O_2752,N_24179,N_24167);
nor UO_2753 (O_2753,N_24015,N_24666);
nand UO_2754 (O_2754,N_24845,N_24521);
xnor UO_2755 (O_2755,N_24254,N_24980);
and UO_2756 (O_2756,N_24655,N_24134);
nand UO_2757 (O_2757,N_24110,N_24243);
nor UO_2758 (O_2758,N_24004,N_24161);
nor UO_2759 (O_2759,N_24012,N_24369);
nand UO_2760 (O_2760,N_24334,N_24305);
nor UO_2761 (O_2761,N_24565,N_24628);
xor UO_2762 (O_2762,N_24844,N_24748);
xnor UO_2763 (O_2763,N_24083,N_24596);
nor UO_2764 (O_2764,N_24767,N_24656);
nand UO_2765 (O_2765,N_24556,N_24919);
nor UO_2766 (O_2766,N_24996,N_24092);
xor UO_2767 (O_2767,N_24351,N_24839);
and UO_2768 (O_2768,N_24410,N_24482);
and UO_2769 (O_2769,N_24846,N_24697);
and UO_2770 (O_2770,N_24125,N_24697);
nand UO_2771 (O_2771,N_24009,N_24125);
or UO_2772 (O_2772,N_24801,N_24007);
and UO_2773 (O_2773,N_24353,N_24843);
and UO_2774 (O_2774,N_24892,N_24107);
or UO_2775 (O_2775,N_24322,N_24077);
or UO_2776 (O_2776,N_24469,N_24082);
xor UO_2777 (O_2777,N_24060,N_24747);
nor UO_2778 (O_2778,N_24130,N_24697);
and UO_2779 (O_2779,N_24375,N_24843);
nand UO_2780 (O_2780,N_24762,N_24903);
nor UO_2781 (O_2781,N_24911,N_24382);
xor UO_2782 (O_2782,N_24210,N_24493);
and UO_2783 (O_2783,N_24533,N_24984);
and UO_2784 (O_2784,N_24362,N_24881);
or UO_2785 (O_2785,N_24043,N_24799);
xnor UO_2786 (O_2786,N_24204,N_24928);
and UO_2787 (O_2787,N_24892,N_24640);
nor UO_2788 (O_2788,N_24409,N_24362);
xnor UO_2789 (O_2789,N_24814,N_24236);
nand UO_2790 (O_2790,N_24712,N_24008);
and UO_2791 (O_2791,N_24035,N_24001);
or UO_2792 (O_2792,N_24693,N_24563);
xnor UO_2793 (O_2793,N_24516,N_24081);
nand UO_2794 (O_2794,N_24339,N_24139);
nor UO_2795 (O_2795,N_24708,N_24380);
xnor UO_2796 (O_2796,N_24735,N_24553);
or UO_2797 (O_2797,N_24309,N_24139);
or UO_2798 (O_2798,N_24839,N_24284);
or UO_2799 (O_2799,N_24046,N_24669);
xnor UO_2800 (O_2800,N_24113,N_24615);
nand UO_2801 (O_2801,N_24956,N_24725);
xor UO_2802 (O_2802,N_24655,N_24345);
or UO_2803 (O_2803,N_24250,N_24813);
xnor UO_2804 (O_2804,N_24227,N_24148);
and UO_2805 (O_2805,N_24533,N_24581);
nand UO_2806 (O_2806,N_24539,N_24039);
and UO_2807 (O_2807,N_24044,N_24007);
and UO_2808 (O_2808,N_24550,N_24408);
xnor UO_2809 (O_2809,N_24791,N_24607);
nand UO_2810 (O_2810,N_24124,N_24501);
nor UO_2811 (O_2811,N_24097,N_24430);
nor UO_2812 (O_2812,N_24693,N_24171);
and UO_2813 (O_2813,N_24971,N_24203);
nor UO_2814 (O_2814,N_24545,N_24691);
and UO_2815 (O_2815,N_24947,N_24345);
nand UO_2816 (O_2816,N_24403,N_24180);
and UO_2817 (O_2817,N_24683,N_24499);
or UO_2818 (O_2818,N_24538,N_24373);
or UO_2819 (O_2819,N_24498,N_24927);
or UO_2820 (O_2820,N_24029,N_24564);
nand UO_2821 (O_2821,N_24291,N_24129);
nand UO_2822 (O_2822,N_24731,N_24239);
or UO_2823 (O_2823,N_24792,N_24673);
or UO_2824 (O_2824,N_24560,N_24845);
nand UO_2825 (O_2825,N_24129,N_24830);
xor UO_2826 (O_2826,N_24326,N_24340);
or UO_2827 (O_2827,N_24517,N_24047);
nand UO_2828 (O_2828,N_24774,N_24607);
nand UO_2829 (O_2829,N_24786,N_24035);
or UO_2830 (O_2830,N_24829,N_24292);
or UO_2831 (O_2831,N_24276,N_24655);
xnor UO_2832 (O_2832,N_24955,N_24475);
xor UO_2833 (O_2833,N_24025,N_24727);
or UO_2834 (O_2834,N_24113,N_24548);
nand UO_2835 (O_2835,N_24717,N_24728);
xor UO_2836 (O_2836,N_24689,N_24517);
and UO_2837 (O_2837,N_24909,N_24986);
or UO_2838 (O_2838,N_24531,N_24078);
or UO_2839 (O_2839,N_24598,N_24838);
xor UO_2840 (O_2840,N_24387,N_24602);
and UO_2841 (O_2841,N_24327,N_24116);
or UO_2842 (O_2842,N_24954,N_24155);
and UO_2843 (O_2843,N_24337,N_24625);
nand UO_2844 (O_2844,N_24926,N_24929);
or UO_2845 (O_2845,N_24805,N_24024);
or UO_2846 (O_2846,N_24653,N_24103);
nand UO_2847 (O_2847,N_24908,N_24863);
and UO_2848 (O_2848,N_24240,N_24945);
nor UO_2849 (O_2849,N_24617,N_24943);
xnor UO_2850 (O_2850,N_24798,N_24231);
xnor UO_2851 (O_2851,N_24649,N_24762);
nor UO_2852 (O_2852,N_24997,N_24586);
nand UO_2853 (O_2853,N_24626,N_24519);
or UO_2854 (O_2854,N_24489,N_24737);
nor UO_2855 (O_2855,N_24410,N_24849);
nor UO_2856 (O_2856,N_24183,N_24011);
or UO_2857 (O_2857,N_24890,N_24179);
and UO_2858 (O_2858,N_24551,N_24155);
nor UO_2859 (O_2859,N_24165,N_24146);
nor UO_2860 (O_2860,N_24583,N_24283);
nor UO_2861 (O_2861,N_24998,N_24567);
and UO_2862 (O_2862,N_24870,N_24573);
and UO_2863 (O_2863,N_24040,N_24624);
or UO_2864 (O_2864,N_24533,N_24075);
and UO_2865 (O_2865,N_24971,N_24102);
and UO_2866 (O_2866,N_24605,N_24242);
nor UO_2867 (O_2867,N_24841,N_24917);
xnor UO_2868 (O_2868,N_24193,N_24387);
or UO_2869 (O_2869,N_24597,N_24575);
nand UO_2870 (O_2870,N_24380,N_24263);
nor UO_2871 (O_2871,N_24749,N_24573);
xor UO_2872 (O_2872,N_24323,N_24652);
nand UO_2873 (O_2873,N_24459,N_24088);
nor UO_2874 (O_2874,N_24774,N_24718);
nor UO_2875 (O_2875,N_24791,N_24265);
xnor UO_2876 (O_2876,N_24828,N_24263);
nand UO_2877 (O_2877,N_24105,N_24457);
nor UO_2878 (O_2878,N_24336,N_24603);
nor UO_2879 (O_2879,N_24347,N_24979);
or UO_2880 (O_2880,N_24437,N_24262);
and UO_2881 (O_2881,N_24855,N_24050);
nor UO_2882 (O_2882,N_24054,N_24176);
nand UO_2883 (O_2883,N_24169,N_24042);
or UO_2884 (O_2884,N_24206,N_24483);
and UO_2885 (O_2885,N_24458,N_24367);
nor UO_2886 (O_2886,N_24236,N_24191);
nor UO_2887 (O_2887,N_24960,N_24585);
xor UO_2888 (O_2888,N_24379,N_24439);
nor UO_2889 (O_2889,N_24979,N_24912);
or UO_2890 (O_2890,N_24531,N_24456);
and UO_2891 (O_2891,N_24145,N_24916);
xnor UO_2892 (O_2892,N_24214,N_24610);
nor UO_2893 (O_2893,N_24795,N_24728);
nand UO_2894 (O_2894,N_24396,N_24230);
xnor UO_2895 (O_2895,N_24618,N_24210);
nand UO_2896 (O_2896,N_24047,N_24367);
nor UO_2897 (O_2897,N_24134,N_24814);
nand UO_2898 (O_2898,N_24472,N_24248);
xor UO_2899 (O_2899,N_24406,N_24471);
nor UO_2900 (O_2900,N_24666,N_24228);
xor UO_2901 (O_2901,N_24993,N_24345);
or UO_2902 (O_2902,N_24830,N_24800);
or UO_2903 (O_2903,N_24560,N_24051);
nor UO_2904 (O_2904,N_24467,N_24242);
and UO_2905 (O_2905,N_24555,N_24373);
xnor UO_2906 (O_2906,N_24534,N_24332);
nor UO_2907 (O_2907,N_24477,N_24023);
nand UO_2908 (O_2908,N_24626,N_24052);
xor UO_2909 (O_2909,N_24919,N_24217);
xor UO_2910 (O_2910,N_24082,N_24974);
or UO_2911 (O_2911,N_24285,N_24236);
nand UO_2912 (O_2912,N_24497,N_24646);
nand UO_2913 (O_2913,N_24135,N_24366);
nor UO_2914 (O_2914,N_24724,N_24820);
nand UO_2915 (O_2915,N_24175,N_24665);
and UO_2916 (O_2916,N_24176,N_24500);
nor UO_2917 (O_2917,N_24015,N_24907);
nand UO_2918 (O_2918,N_24399,N_24191);
or UO_2919 (O_2919,N_24875,N_24212);
nand UO_2920 (O_2920,N_24224,N_24350);
or UO_2921 (O_2921,N_24553,N_24097);
or UO_2922 (O_2922,N_24565,N_24347);
and UO_2923 (O_2923,N_24084,N_24119);
or UO_2924 (O_2924,N_24067,N_24341);
nor UO_2925 (O_2925,N_24227,N_24903);
or UO_2926 (O_2926,N_24205,N_24462);
or UO_2927 (O_2927,N_24512,N_24302);
nand UO_2928 (O_2928,N_24542,N_24623);
nor UO_2929 (O_2929,N_24275,N_24764);
xnor UO_2930 (O_2930,N_24006,N_24546);
or UO_2931 (O_2931,N_24163,N_24232);
nor UO_2932 (O_2932,N_24597,N_24594);
nor UO_2933 (O_2933,N_24118,N_24411);
xor UO_2934 (O_2934,N_24568,N_24120);
or UO_2935 (O_2935,N_24597,N_24631);
and UO_2936 (O_2936,N_24130,N_24620);
nor UO_2937 (O_2937,N_24708,N_24974);
nand UO_2938 (O_2938,N_24053,N_24108);
or UO_2939 (O_2939,N_24080,N_24323);
or UO_2940 (O_2940,N_24979,N_24580);
or UO_2941 (O_2941,N_24069,N_24065);
nor UO_2942 (O_2942,N_24424,N_24408);
xor UO_2943 (O_2943,N_24155,N_24962);
nand UO_2944 (O_2944,N_24854,N_24525);
and UO_2945 (O_2945,N_24934,N_24762);
and UO_2946 (O_2946,N_24063,N_24475);
or UO_2947 (O_2947,N_24534,N_24478);
and UO_2948 (O_2948,N_24360,N_24685);
xnor UO_2949 (O_2949,N_24759,N_24690);
or UO_2950 (O_2950,N_24595,N_24026);
or UO_2951 (O_2951,N_24047,N_24522);
nor UO_2952 (O_2952,N_24348,N_24574);
xnor UO_2953 (O_2953,N_24775,N_24430);
nor UO_2954 (O_2954,N_24400,N_24365);
and UO_2955 (O_2955,N_24187,N_24436);
or UO_2956 (O_2956,N_24893,N_24492);
nand UO_2957 (O_2957,N_24424,N_24227);
nand UO_2958 (O_2958,N_24455,N_24494);
xor UO_2959 (O_2959,N_24973,N_24349);
or UO_2960 (O_2960,N_24633,N_24987);
or UO_2961 (O_2961,N_24029,N_24669);
and UO_2962 (O_2962,N_24992,N_24969);
nor UO_2963 (O_2963,N_24854,N_24240);
nor UO_2964 (O_2964,N_24959,N_24453);
nor UO_2965 (O_2965,N_24409,N_24792);
nor UO_2966 (O_2966,N_24372,N_24750);
xor UO_2967 (O_2967,N_24696,N_24928);
and UO_2968 (O_2968,N_24307,N_24499);
nor UO_2969 (O_2969,N_24155,N_24576);
xnor UO_2970 (O_2970,N_24225,N_24720);
nand UO_2971 (O_2971,N_24004,N_24579);
or UO_2972 (O_2972,N_24574,N_24913);
and UO_2973 (O_2973,N_24398,N_24223);
or UO_2974 (O_2974,N_24283,N_24192);
nor UO_2975 (O_2975,N_24252,N_24843);
and UO_2976 (O_2976,N_24305,N_24992);
xnor UO_2977 (O_2977,N_24714,N_24691);
xor UO_2978 (O_2978,N_24817,N_24454);
nand UO_2979 (O_2979,N_24961,N_24262);
nor UO_2980 (O_2980,N_24633,N_24504);
nand UO_2981 (O_2981,N_24486,N_24158);
nor UO_2982 (O_2982,N_24723,N_24909);
and UO_2983 (O_2983,N_24431,N_24280);
xor UO_2984 (O_2984,N_24586,N_24248);
or UO_2985 (O_2985,N_24222,N_24757);
nor UO_2986 (O_2986,N_24249,N_24068);
xor UO_2987 (O_2987,N_24242,N_24655);
and UO_2988 (O_2988,N_24051,N_24133);
nand UO_2989 (O_2989,N_24670,N_24035);
and UO_2990 (O_2990,N_24063,N_24709);
xor UO_2991 (O_2991,N_24668,N_24938);
nand UO_2992 (O_2992,N_24277,N_24655);
nand UO_2993 (O_2993,N_24892,N_24290);
nand UO_2994 (O_2994,N_24567,N_24409);
and UO_2995 (O_2995,N_24581,N_24028);
xor UO_2996 (O_2996,N_24648,N_24224);
and UO_2997 (O_2997,N_24148,N_24119);
xnor UO_2998 (O_2998,N_24427,N_24557);
nand UO_2999 (O_2999,N_24943,N_24937);
endmodule