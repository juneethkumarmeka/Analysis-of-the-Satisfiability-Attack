module basic_500_3000_500_60_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_65,In_379);
and U1 (N_1,In_204,In_498);
or U2 (N_2,In_131,In_290);
and U3 (N_3,In_4,In_159);
and U4 (N_4,In_428,In_2);
nor U5 (N_5,In_45,In_161);
and U6 (N_6,In_56,In_43);
and U7 (N_7,In_110,In_256);
or U8 (N_8,In_404,In_480);
or U9 (N_9,In_3,In_75);
or U10 (N_10,In_13,In_128);
and U11 (N_11,In_400,In_457);
or U12 (N_12,In_318,In_314);
and U13 (N_13,In_153,In_89);
and U14 (N_14,In_430,In_420);
nand U15 (N_15,In_36,In_281);
or U16 (N_16,In_349,In_450);
nor U17 (N_17,In_439,In_178);
or U18 (N_18,In_257,In_491);
nor U19 (N_19,In_344,In_162);
nand U20 (N_20,In_396,In_390);
or U21 (N_21,In_367,In_332);
nand U22 (N_22,In_405,In_463);
or U23 (N_23,In_120,In_435);
or U24 (N_24,In_326,In_499);
nand U25 (N_25,In_299,In_252);
or U26 (N_26,In_490,In_248);
nor U27 (N_27,In_223,In_164);
and U28 (N_28,In_66,In_460);
nor U29 (N_29,In_239,In_98);
or U30 (N_30,In_482,In_412);
nand U31 (N_31,In_35,In_316);
nand U32 (N_32,In_456,In_339);
or U33 (N_33,In_145,In_81);
and U34 (N_34,In_144,In_214);
or U35 (N_35,In_307,In_308);
and U36 (N_36,In_88,In_293);
and U37 (N_37,In_364,In_429);
nand U38 (N_38,In_215,In_15);
nand U39 (N_39,In_250,In_315);
nor U40 (N_40,In_287,In_298);
nor U41 (N_41,In_224,In_355);
or U42 (N_42,In_21,In_126);
nor U43 (N_43,In_485,In_113);
nand U44 (N_44,In_286,In_166);
nor U45 (N_45,In_475,In_20);
nand U46 (N_46,In_442,In_233);
nor U47 (N_47,In_279,In_397);
or U48 (N_48,In_52,In_30);
nor U49 (N_49,In_322,In_212);
and U50 (N_50,In_380,In_391);
and U51 (N_51,In_271,In_92);
or U52 (N_52,N_45,In_320);
nand U53 (N_53,In_359,In_372);
and U54 (N_54,In_181,In_80);
nand U55 (N_55,In_48,In_292);
nand U56 (N_56,In_234,In_109);
nor U57 (N_57,In_445,In_115);
nor U58 (N_58,In_305,In_259);
and U59 (N_59,In_276,In_329);
nand U60 (N_60,N_44,In_353);
nor U61 (N_61,In_246,In_73);
and U62 (N_62,In_107,In_9);
nor U63 (N_63,In_179,In_229);
and U64 (N_64,N_29,N_25);
and U65 (N_65,In_97,In_177);
and U66 (N_66,In_94,In_365);
or U67 (N_67,In_330,In_347);
or U68 (N_68,In_213,In_392);
and U69 (N_69,In_394,In_206);
or U70 (N_70,In_407,In_225);
and U71 (N_71,In_174,In_302);
nand U72 (N_72,In_373,In_395);
nor U73 (N_73,In_284,In_23);
xor U74 (N_74,In_325,In_471);
or U75 (N_75,In_467,In_348);
nand U76 (N_76,N_4,In_44);
and U77 (N_77,In_415,N_41);
and U78 (N_78,In_64,In_87);
or U79 (N_79,In_388,In_247);
nand U80 (N_80,In_103,In_492);
nor U81 (N_81,In_438,In_300);
nand U82 (N_82,In_282,In_139);
and U83 (N_83,In_78,In_7);
nor U84 (N_84,In_67,In_436);
nor U85 (N_85,In_389,N_35);
and U86 (N_86,In_195,In_142);
nor U87 (N_87,N_9,In_297);
nor U88 (N_88,In_207,In_453);
and U89 (N_89,N_33,N_34);
and U90 (N_90,In_51,In_25);
and U91 (N_91,In_474,In_49);
or U92 (N_92,In_346,N_48);
nand U93 (N_93,In_190,N_0);
nor U94 (N_94,In_419,In_459);
nor U95 (N_95,In_193,In_335);
nand U96 (N_96,In_187,In_61);
or U97 (N_97,In_345,In_40);
or U98 (N_98,In_0,In_433);
and U99 (N_99,In_155,In_116);
and U100 (N_100,In_150,In_50);
nor U101 (N_101,N_72,In_356);
and U102 (N_102,In_102,In_211);
nand U103 (N_103,In_461,In_173);
and U104 (N_104,N_68,In_185);
and U105 (N_105,N_50,In_28);
or U106 (N_106,In_220,N_89);
or U107 (N_107,In_93,In_125);
or U108 (N_108,N_60,In_437);
and U109 (N_109,In_427,N_15);
or U110 (N_110,In_141,In_446);
and U111 (N_111,In_455,In_494);
and U112 (N_112,In_452,In_197);
nand U113 (N_113,In_312,In_238);
or U114 (N_114,In_321,In_301);
xnor U115 (N_115,In_260,In_488);
nand U116 (N_116,In_63,In_383);
and U117 (N_117,N_1,In_263);
or U118 (N_118,In_447,In_68);
nand U119 (N_119,In_358,N_3);
xnor U120 (N_120,N_51,In_294);
nor U121 (N_121,In_458,In_351);
nand U122 (N_122,In_289,N_36);
nor U123 (N_123,In_38,In_117);
nor U124 (N_124,N_54,In_273);
nor U125 (N_125,In_118,In_241);
and U126 (N_126,In_283,In_146);
nor U127 (N_127,In_47,In_418);
or U128 (N_128,N_85,In_194);
nand U129 (N_129,In_310,In_403);
nand U130 (N_130,In_341,In_129);
nand U131 (N_131,In_242,In_483);
or U132 (N_132,In_333,In_134);
or U133 (N_133,N_18,In_19);
nand U134 (N_134,In_278,N_8);
or U135 (N_135,In_11,In_100);
nand U136 (N_136,In_170,In_199);
and U137 (N_137,In_338,N_39);
and U138 (N_138,In_83,N_97);
or U139 (N_139,In_148,In_72);
or U140 (N_140,In_236,In_484);
nand U141 (N_141,In_169,In_105);
nand U142 (N_142,In_154,N_76);
and U143 (N_143,N_99,In_465);
or U144 (N_144,In_431,In_147);
and U145 (N_145,N_77,In_217);
nand U146 (N_146,N_37,N_43);
nor U147 (N_147,N_92,In_473);
nor U148 (N_148,N_5,In_386);
and U149 (N_149,N_13,In_265);
nand U150 (N_150,In_269,In_138);
nor U151 (N_151,In_253,N_73);
and U152 (N_152,In_493,N_106);
or U153 (N_153,N_132,In_37);
and U154 (N_154,In_327,N_2);
and U155 (N_155,In_149,In_272);
nor U156 (N_156,N_87,In_10);
nor U157 (N_157,N_47,N_22);
and U158 (N_158,In_410,In_244);
nand U159 (N_159,N_137,In_409);
and U160 (N_160,N_17,N_30);
nor U161 (N_161,N_108,In_165);
nor U162 (N_162,In_231,N_28);
and U163 (N_163,In_34,N_123);
nand U164 (N_164,In_479,In_378);
nor U165 (N_165,N_90,N_124);
or U166 (N_166,In_156,In_16);
and U167 (N_167,In_441,In_313);
or U168 (N_168,In_375,In_132);
nor U169 (N_169,In_137,In_425);
and U170 (N_170,In_340,N_91);
or U171 (N_171,In_168,In_95);
or U172 (N_172,N_143,In_189);
nand U173 (N_173,N_31,In_472);
and U174 (N_174,N_125,In_426);
nand U175 (N_175,In_200,In_368);
xor U176 (N_176,In_449,In_411);
or U177 (N_177,N_59,In_57);
and U178 (N_178,N_114,In_91);
or U179 (N_179,In_258,In_466);
and U180 (N_180,N_78,In_74);
nand U181 (N_181,In_124,In_434);
nor U182 (N_182,N_110,In_121);
nand U183 (N_183,In_454,In_86);
nand U184 (N_184,In_443,N_71);
and U185 (N_185,N_84,In_470);
or U186 (N_186,N_12,N_81);
nand U187 (N_187,N_116,In_387);
nand U188 (N_188,In_221,In_432);
or U189 (N_189,In_85,In_202);
nand U190 (N_190,In_481,In_377);
nand U191 (N_191,N_140,In_270);
or U192 (N_192,In_423,In_317);
nand U193 (N_193,N_120,In_254);
and U194 (N_194,In_402,In_366);
or U195 (N_195,In_328,In_143);
nor U196 (N_196,In_324,In_267);
nand U197 (N_197,N_112,In_255);
or U198 (N_198,N_95,N_146);
and U199 (N_199,In_136,In_209);
and U200 (N_200,N_178,N_180);
and U201 (N_201,In_381,N_138);
and U202 (N_202,In_401,In_69);
nand U203 (N_203,N_52,N_161);
nand U204 (N_204,In_235,In_249);
or U205 (N_205,N_171,In_22);
and U206 (N_206,N_109,In_352);
nor U207 (N_207,In_203,In_183);
and U208 (N_208,In_261,In_476);
nand U209 (N_209,In_274,In_323);
and U210 (N_210,In_106,N_93);
nand U211 (N_211,N_142,In_188);
nand U212 (N_212,N_62,In_8);
nor U213 (N_213,N_186,In_489);
and U214 (N_214,In_151,In_354);
nor U215 (N_215,In_487,N_57);
and U216 (N_216,N_154,N_75);
and U217 (N_217,In_350,N_128);
or U218 (N_218,N_152,N_46);
nand U219 (N_219,In_264,In_33);
or U220 (N_220,N_198,In_62);
or U221 (N_221,N_61,N_173);
nor U222 (N_222,N_7,N_86);
nand U223 (N_223,In_230,In_167);
nor U224 (N_224,In_160,N_14);
nor U225 (N_225,N_150,In_14);
nand U226 (N_226,In_266,In_198);
nand U227 (N_227,N_115,N_118);
or U228 (N_228,In_127,In_76);
and U229 (N_229,In_382,In_413);
xnor U230 (N_230,In_1,N_183);
nand U231 (N_231,N_167,In_495);
and U232 (N_232,N_181,In_296);
nand U233 (N_233,In_398,In_245);
or U234 (N_234,N_107,N_156);
nor U235 (N_235,In_357,In_304);
and U236 (N_236,In_384,N_122);
nor U237 (N_237,N_105,N_74);
or U238 (N_238,In_370,In_451);
nand U239 (N_239,In_54,N_197);
nor U240 (N_240,N_182,In_222);
or U241 (N_241,N_53,N_6);
and U242 (N_242,In_112,In_414);
and U243 (N_243,In_227,In_104);
or U244 (N_244,N_96,In_361);
or U245 (N_245,In_24,N_80);
nand U246 (N_246,In_306,In_122);
nor U247 (N_247,In_440,N_193);
nand U248 (N_248,In_478,In_275);
nand U249 (N_249,In_180,N_83);
or U250 (N_250,In_277,In_295);
or U251 (N_251,N_119,N_165);
xor U252 (N_252,N_194,N_103);
or U253 (N_253,In_99,In_399);
nand U254 (N_254,N_247,In_343);
nand U255 (N_255,N_222,N_100);
or U256 (N_256,In_42,In_39);
nor U257 (N_257,N_175,In_191);
nand U258 (N_258,In_416,N_63);
nand U259 (N_259,N_139,N_230);
and U260 (N_260,In_108,In_422);
nor U261 (N_261,N_188,N_214);
nor U262 (N_262,N_179,N_241);
and U263 (N_263,N_160,N_20);
nor U264 (N_264,N_243,N_70);
nand U265 (N_265,N_206,N_169);
or U266 (N_266,In_251,N_233);
or U267 (N_267,N_205,N_136);
and U268 (N_268,N_134,In_336);
nand U269 (N_269,N_189,N_218);
nand U270 (N_270,In_309,N_219);
nor U271 (N_271,In_291,N_144);
nand U272 (N_272,In_114,N_133);
nor U273 (N_273,N_19,N_121);
nand U274 (N_274,In_468,N_201);
nand U275 (N_275,In_311,In_196);
nand U276 (N_276,N_69,In_496);
and U277 (N_277,N_234,In_374);
or U278 (N_278,N_58,N_40);
nor U279 (N_279,In_280,N_141);
nand U280 (N_280,N_215,N_248);
nand U281 (N_281,N_237,N_153);
nand U282 (N_282,N_212,N_10);
nor U283 (N_283,In_158,N_225);
and U284 (N_284,N_204,In_163);
and U285 (N_285,N_209,In_424);
and U286 (N_286,In_17,N_113);
nand U287 (N_287,N_168,N_155);
nand U288 (N_288,In_130,In_417);
nor U289 (N_289,N_226,In_218);
and U290 (N_290,In_101,In_176);
and U291 (N_291,N_27,N_221);
or U292 (N_292,N_232,In_133);
nor U293 (N_293,In_171,N_249);
and U294 (N_294,In_243,N_242);
or U295 (N_295,N_42,N_162);
or U296 (N_296,N_238,In_201);
and U297 (N_297,In_462,N_130);
and U298 (N_298,N_104,N_224);
or U299 (N_299,In_369,In_228);
and U300 (N_300,N_294,N_276);
and U301 (N_301,N_111,N_261);
nand U302 (N_302,N_172,N_163);
and U303 (N_303,N_217,In_53);
or U304 (N_304,N_292,In_175);
nor U305 (N_305,N_56,N_257);
nand U306 (N_306,In_182,N_259);
or U307 (N_307,N_157,N_166);
nand U308 (N_308,In_58,In_27);
or U309 (N_309,In_186,In_18);
or U310 (N_310,N_255,N_228);
or U311 (N_311,N_23,N_126);
or U312 (N_312,In_157,N_266);
and U313 (N_313,In_363,N_199);
nor U314 (N_314,N_82,N_252);
or U315 (N_315,In_84,In_337);
or U316 (N_316,N_271,In_29);
or U317 (N_317,N_11,N_273);
nand U318 (N_318,In_172,N_246);
and U319 (N_319,In_448,N_94);
or U320 (N_320,In_342,N_170);
and U321 (N_321,In_111,N_102);
nand U322 (N_322,In_226,N_177);
or U323 (N_323,N_147,In_70);
nand U324 (N_324,N_275,In_152);
nand U325 (N_325,N_216,N_245);
or U326 (N_326,N_210,N_256);
nor U327 (N_327,In_6,In_334);
xnor U328 (N_328,In_123,N_277);
or U329 (N_329,N_287,N_101);
and U330 (N_330,N_270,N_289);
nand U331 (N_331,N_98,N_158);
or U332 (N_332,N_135,In_393);
nor U333 (N_333,N_159,N_293);
or U334 (N_334,N_66,N_202);
nand U335 (N_335,N_24,N_286);
and U336 (N_336,N_283,N_200);
nor U337 (N_337,N_262,In_385);
and U338 (N_338,In_303,N_272);
nor U339 (N_339,N_88,N_298);
and U340 (N_340,In_421,In_371);
or U341 (N_341,N_21,N_67);
and U342 (N_342,N_264,N_213);
nand U343 (N_343,In_240,In_444);
or U344 (N_344,In_331,N_145);
or U345 (N_345,N_290,N_295);
nor U346 (N_346,In_12,N_16);
nand U347 (N_347,In_135,In_31);
nor U348 (N_348,In_192,In_32);
nor U349 (N_349,N_253,N_274);
nor U350 (N_350,N_236,N_55);
nor U351 (N_351,N_339,In_210);
nand U352 (N_352,N_269,N_347);
or U353 (N_353,N_337,N_320);
and U354 (N_354,In_406,N_227);
and U355 (N_355,N_129,N_174);
nand U356 (N_356,N_240,N_250);
nand U357 (N_357,N_307,In_268);
nor U358 (N_358,N_302,N_296);
nor U359 (N_359,N_325,N_260);
and U360 (N_360,In_82,N_319);
nor U361 (N_361,N_329,In_469);
nor U362 (N_362,N_326,N_191);
nor U363 (N_363,N_151,In_237);
nor U364 (N_364,In_71,N_207);
nor U365 (N_365,In_96,N_348);
nor U366 (N_366,In_77,N_345);
nor U367 (N_367,N_279,N_117);
nand U368 (N_368,N_211,N_32);
nand U369 (N_369,N_323,N_333);
or U370 (N_370,N_223,In_41);
nor U371 (N_371,N_278,N_79);
xnor U372 (N_372,In_319,In_486);
nand U373 (N_373,N_334,N_304);
nand U374 (N_374,N_299,In_184);
nor U375 (N_375,N_331,N_321);
nand U376 (N_376,N_324,In_5);
and U377 (N_377,N_127,N_330);
and U378 (N_378,N_305,N_340);
nor U379 (N_379,In_477,In_262);
nand U380 (N_380,In_90,N_309);
and U381 (N_381,N_318,N_315);
nor U382 (N_382,N_332,N_195);
nand U383 (N_383,N_65,N_297);
nand U384 (N_384,N_220,N_190);
or U385 (N_385,N_346,N_322);
nand U386 (N_386,N_282,N_244);
nor U387 (N_387,N_288,N_26);
nor U388 (N_388,N_267,N_149);
and U389 (N_389,N_303,N_196);
nand U390 (N_390,N_312,In_497);
nand U391 (N_391,N_310,N_281);
nand U392 (N_392,N_265,In_360);
nor U393 (N_393,In_408,In_205);
and U394 (N_394,In_59,N_314);
and U395 (N_395,N_328,N_284);
or U396 (N_396,In_26,N_317);
and U397 (N_397,N_229,N_306);
nand U398 (N_398,N_349,N_185);
and U399 (N_399,N_342,In_219);
nand U400 (N_400,N_285,N_338);
nand U401 (N_401,In_119,N_358);
and U402 (N_402,N_254,N_387);
or U403 (N_403,N_396,N_368);
nor U404 (N_404,N_389,N_374);
and U405 (N_405,N_388,N_176);
and U406 (N_406,N_291,N_393);
or U407 (N_407,In_216,N_352);
nand U408 (N_408,N_384,In_46);
and U409 (N_409,In_362,N_148);
nand U410 (N_410,N_357,N_385);
and U411 (N_411,N_316,In_55);
nand U412 (N_412,In_79,N_64);
or U413 (N_413,N_377,N_353);
nor U414 (N_414,N_38,N_187);
and U415 (N_415,N_370,N_373);
or U416 (N_416,In_60,N_351);
and U417 (N_417,N_362,N_371);
nor U418 (N_418,N_382,N_268);
or U419 (N_419,In_208,N_364);
and U420 (N_420,N_327,N_300);
nand U421 (N_421,N_231,N_394);
nand U422 (N_422,N_251,N_208);
nand U423 (N_423,N_397,N_344);
nand U424 (N_424,N_376,N_378);
nor U425 (N_425,N_184,N_239);
nand U426 (N_426,N_380,N_263);
nor U427 (N_427,N_383,In_140);
nand U428 (N_428,N_369,N_359);
and U429 (N_429,N_192,N_235);
or U430 (N_430,N_49,In_288);
nor U431 (N_431,N_392,N_301);
or U432 (N_432,N_381,N_308);
nor U433 (N_433,N_350,N_356);
or U434 (N_434,N_372,N_355);
and U435 (N_435,N_258,N_399);
and U436 (N_436,In_232,N_313);
nand U437 (N_437,N_354,N_365);
nand U438 (N_438,N_164,N_395);
nor U439 (N_439,N_311,N_390);
or U440 (N_440,N_336,N_363);
and U441 (N_441,In_285,In_464);
or U442 (N_442,N_375,N_341);
and U443 (N_443,In_376,N_379);
or U444 (N_444,N_335,N_280);
and U445 (N_445,N_361,N_398);
nor U446 (N_446,N_360,N_366);
or U447 (N_447,N_343,N_203);
and U448 (N_448,N_386,N_391);
xnor U449 (N_449,N_131,N_367);
nor U450 (N_450,N_444,N_400);
and U451 (N_451,N_447,N_420);
and U452 (N_452,N_405,N_422);
and U453 (N_453,N_421,N_416);
and U454 (N_454,N_441,N_406);
or U455 (N_455,N_418,N_438);
nand U456 (N_456,N_413,N_401);
nor U457 (N_457,N_428,N_424);
nand U458 (N_458,N_404,N_410);
nor U459 (N_459,N_429,N_408);
or U460 (N_460,N_417,N_435);
or U461 (N_461,N_432,N_411);
or U462 (N_462,N_433,N_440);
or U463 (N_463,N_439,N_412);
nor U464 (N_464,N_437,N_434);
nand U465 (N_465,N_415,N_448);
and U466 (N_466,N_423,N_442);
nor U467 (N_467,N_446,N_407);
nor U468 (N_468,N_449,N_403);
nor U469 (N_469,N_427,N_443);
nand U470 (N_470,N_426,N_409);
and U471 (N_471,N_425,N_431);
or U472 (N_472,N_419,N_414);
and U473 (N_473,N_402,N_436);
nor U474 (N_474,N_445,N_430);
or U475 (N_475,N_404,N_435);
or U476 (N_476,N_433,N_446);
nor U477 (N_477,N_425,N_424);
and U478 (N_478,N_431,N_442);
and U479 (N_479,N_403,N_442);
and U480 (N_480,N_404,N_417);
and U481 (N_481,N_428,N_437);
nand U482 (N_482,N_446,N_435);
nand U483 (N_483,N_408,N_420);
and U484 (N_484,N_444,N_428);
or U485 (N_485,N_439,N_442);
nor U486 (N_486,N_420,N_402);
or U487 (N_487,N_441,N_447);
or U488 (N_488,N_443,N_410);
or U489 (N_489,N_436,N_419);
nand U490 (N_490,N_412,N_416);
or U491 (N_491,N_441,N_411);
nor U492 (N_492,N_438,N_449);
and U493 (N_493,N_432,N_400);
nand U494 (N_494,N_411,N_405);
nand U495 (N_495,N_417,N_432);
and U496 (N_496,N_403,N_400);
nand U497 (N_497,N_435,N_419);
and U498 (N_498,N_444,N_442);
nor U499 (N_499,N_407,N_406);
xor U500 (N_500,N_453,N_498);
or U501 (N_501,N_472,N_484);
and U502 (N_502,N_471,N_479);
nor U503 (N_503,N_475,N_494);
and U504 (N_504,N_450,N_473);
and U505 (N_505,N_490,N_469);
and U506 (N_506,N_499,N_462);
nand U507 (N_507,N_460,N_464);
and U508 (N_508,N_474,N_456);
nand U509 (N_509,N_495,N_488);
nor U510 (N_510,N_487,N_455);
nand U511 (N_511,N_457,N_465);
and U512 (N_512,N_458,N_493);
nor U513 (N_513,N_467,N_477);
nand U514 (N_514,N_451,N_480);
nor U515 (N_515,N_492,N_454);
and U516 (N_516,N_463,N_452);
nand U517 (N_517,N_466,N_491);
nor U518 (N_518,N_470,N_496);
nor U519 (N_519,N_468,N_483);
nor U520 (N_520,N_461,N_497);
nor U521 (N_521,N_481,N_486);
nand U522 (N_522,N_476,N_482);
nand U523 (N_523,N_489,N_485);
nor U524 (N_524,N_459,N_478);
and U525 (N_525,N_470,N_462);
or U526 (N_526,N_476,N_495);
or U527 (N_527,N_491,N_468);
nand U528 (N_528,N_484,N_488);
and U529 (N_529,N_462,N_468);
and U530 (N_530,N_452,N_467);
nor U531 (N_531,N_491,N_498);
nand U532 (N_532,N_499,N_450);
and U533 (N_533,N_484,N_475);
nand U534 (N_534,N_451,N_470);
nand U535 (N_535,N_476,N_464);
nor U536 (N_536,N_466,N_469);
and U537 (N_537,N_491,N_472);
and U538 (N_538,N_479,N_475);
or U539 (N_539,N_496,N_467);
nand U540 (N_540,N_462,N_480);
or U541 (N_541,N_484,N_480);
nor U542 (N_542,N_464,N_455);
xor U543 (N_543,N_464,N_452);
or U544 (N_544,N_461,N_495);
or U545 (N_545,N_480,N_464);
and U546 (N_546,N_497,N_488);
nand U547 (N_547,N_453,N_450);
or U548 (N_548,N_465,N_476);
and U549 (N_549,N_459,N_465);
or U550 (N_550,N_537,N_532);
nand U551 (N_551,N_500,N_538);
nand U552 (N_552,N_547,N_530);
nand U553 (N_553,N_527,N_501);
xor U554 (N_554,N_515,N_526);
nand U555 (N_555,N_509,N_543);
nand U556 (N_556,N_540,N_523);
and U557 (N_557,N_514,N_521);
nand U558 (N_558,N_528,N_545);
nand U559 (N_559,N_502,N_516);
or U560 (N_560,N_535,N_512);
and U561 (N_561,N_508,N_529);
nor U562 (N_562,N_504,N_546);
nand U563 (N_563,N_519,N_536);
nand U564 (N_564,N_510,N_506);
and U565 (N_565,N_533,N_541);
nand U566 (N_566,N_548,N_505);
nand U567 (N_567,N_534,N_517);
and U568 (N_568,N_525,N_544);
and U569 (N_569,N_503,N_524);
and U570 (N_570,N_518,N_520);
nor U571 (N_571,N_511,N_507);
or U572 (N_572,N_539,N_542);
nor U573 (N_573,N_513,N_549);
nor U574 (N_574,N_531,N_522);
and U575 (N_575,N_506,N_517);
and U576 (N_576,N_520,N_544);
nor U577 (N_577,N_531,N_538);
or U578 (N_578,N_538,N_520);
nand U579 (N_579,N_532,N_531);
nor U580 (N_580,N_504,N_501);
nor U581 (N_581,N_520,N_527);
nor U582 (N_582,N_503,N_506);
and U583 (N_583,N_500,N_517);
and U584 (N_584,N_534,N_533);
nand U585 (N_585,N_518,N_504);
nor U586 (N_586,N_532,N_534);
and U587 (N_587,N_501,N_525);
nand U588 (N_588,N_528,N_525);
or U589 (N_589,N_545,N_540);
nand U590 (N_590,N_542,N_513);
and U591 (N_591,N_522,N_502);
and U592 (N_592,N_526,N_519);
nand U593 (N_593,N_510,N_519);
nand U594 (N_594,N_520,N_512);
xor U595 (N_595,N_504,N_508);
or U596 (N_596,N_531,N_527);
nor U597 (N_597,N_512,N_513);
nand U598 (N_598,N_546,N_514);
nand U599 (N_599,N_546,N_500);
or U600 (N_600,N_583,N_582);
nor U601 (N_601,N_594,N_562);
nand U602 (N_602,N_561,N_567);
and U603 (N_603,N_556,N_566);
or U604 (N_604,N_585,N_555);
xor U605 (N_605,N_568,N_589);
nor U606 (N_606,N_553,N_573);
or U607 (N_607,N_554,N_564);
nand U608 (N_608,N_563,N_591);
nor U609 (N_609,N_576,N_596);
nor U610 (N_610,N_597,N_558);
or U611 (N_611,N_592,N_577);
nor U612 (N_612,N_557,N_551);
nor U613 (N_613,N_572,N_550);
xnor U614 (N_614,N_570,N_559);
nor U615 (N_615,N_593,N_599);
and U616 (N_616,N_584,N_588);
nor U617 (N_617,N_552,N_595);
nand U618 (N_618,N_569,N_575);
or U619 (N_619,N_579,N_580);
xor U620 (N_620,N_586,N_581);
nor U621 (N_621,N_571,N_598);
or U622 (N_622,N_587,N_574);
nor U623 (N_623,N_578,N_590);
or U624 (N_624,N_565,N_560);
nor U625 (N_625,N_578,N_555);
nor U626 (N_626,N_558,N_577);
nor U627 (N_627,N_582,N_588);
or U628 (N_628,N_591,N_587);
or U629 (N_629,N_576,N_595);
nor U630 (N_630,N_591,N_552);
and U631 (N_631,N_552,N_593);
or U632 (N_632,N_569,N_568);
or U633 (N_633,N_580,N_556);
and U634 (N_634,N_579,N_585);
and U635 (N_635,N_573,N_593);
nand U636 (N_636,N_587,N_575);
nand U637 (N_637,N_565,N_571);
and U638 (N_638,N_567,N_590);
nand U639 (N_639,N_591,N_550);
nor U640 (N_640,N_598,N_568);
nand U641 (N_641,N_562,N_575);
and U642 (N_642,N_579,N_584);
nand U643 (N_643,N_598,N_563);
nor U644 (N_644,N_552,N_587);
or U645 (N_645,N_568,N_561);
nor U646 (N_646,N_566,N_591);
nor U647 (N_647,N_552,N_596);
and U648 (N_648,N_563,N_550);
nor U649 (N_649,N_555,N_590);
nand U650 (N_650,N_637,N_623);
and U651 (N_651,N_646,N_639);
or U652 (N_652,N_633,N_600);
or U653 (N_653,N_649,N_631);
nor U654 (N_654,N_647,N_628);
and U655 (N_655,N_627,N_626);
and U656 (N_656,N_617,N_644);
nor U657 (N_657,N_645,N_611);
or U658 (N_658,N_629,N_640);
and U659 (N_659,N_630,N_615);
nor U660 (N_660,N_648,N_643);
nor U661 (N_661,N_620,N_619);
and U662 (N_662,N_618,N_613);
nor U663 (N_663,N_634,N_612);
nand U664 (N_664,N_614,N_642);
nand U665 (N_665,N_632,N_607);
or U666 (N_666,N_606,N_638);
or U667 (N_667,N_625,N_616);
or U668 (N_668,N_602,N_609);
nand U669 (N_669,N_601,N_608);
nand U670 (N_670,N_624,N_641);
or U671 (N_671,N_622,N_610);
and U672 (N_672,N_603,N_605);
or U673 (N_673,N_604,N_621);
nand U674 (N_674,N_636,N_635);
nor U675 (N_675,N_628,N_613);
and U676 (N_676,N_639,N_644);
and U677 (N_677,N_608,N_628);
and U678 (N_678,N_638,N_614);
nand U679 (N_679,N_632,N_616);
and U680 (N_680,N_623,N_624);
and U681 (N_681,N_628,N_627);
nand U682 (N_682,N_622,N_619);
nand U683 (N_683,N_622,N_612);
nor U684 (N_684,N_643,N_640);
and U685 (N_685,N_627,N_630);
nor U686 (N_686,N_618,N_634);
and U687 (N_687,N_634,N_630);
and U688 (N_688,N_637,N_601);
or U689 (N_689,N_647,N_646);
nand U690 (N_690,N_612,N_645);
nand U691 (N_691,N_626,N_611);
or U692 (N_692,N_640,N_605);
nor U693 (N_693,N_621,N_638);
nand U694 (N_694,N_628,N_642);
and U695 (N_695,N_632,N_611);
or U696 (N_696,N_623,N_618);
nand U697 (N_697,N_626,N_607);
or U698 (N_698,N_641,N_611);
and U699 (N_699,N_606,N_611);
nor U700 (N_700,N_666,N_683);
or U701 (N_701,N_665,N_671);
nor U702 (N_702,N_680,N_678);
or U703 (N_703,N_676,N_697);
and U704 (N_704,N_696,N_687);
nor U705 (N_705,N_651,N_681);
nor U706 (N_706,N_667,N_669);
and U707 (N_707,N_698,N_662);
and U708 (N_708,N_679,N_685);
and U709 (N_709,N_694,N_688);
or U710 (N_710,N_664,N_693);
nand U711 (N_711,N_653,N_660);
or U712 (N_712,N_668,N_656);
nand U713 (N_713,N_674,N_657);
or U714 (N_714,N_689,N_692);
nor U715 (N_715,N_652,N_677);
nor U716 (N_716,N_695,N_659);
and U717 (N_717,N_684,N_691);
nand U718 (N_718,N_682,N_650);
nor U719 (N_719,N_663,N_690);
nor U720 (N_720,N_654,N_670);
nand U721 (N_721,N_658,N_672);
xor U722 (N_722,N_686,N_699);
nor U723 (N_723,N_675,N_661);
nand U724 (N_724,N_673,N_655);
and U725 (N_725,N_652,N_699);
nand U726 (N_726,N_699,N_654);
nor U727 (N_727,N_654,N_678);
or U728 (N_728,N_664,N_691);
nand U729 (N_729,N_689,N_655);
and U730 (N_730,N_679,N_699);
nand U731 (N_731,N_650,N_692);
and U732 (N_732,N_661,N_699);
nor U733 (N_733,N_651,N_694);
and U734 (N_734,N_671,N_698);
nor U735 (N_735,N_667,N_697);
nor U736 (N_736,N_690,N_656);
nor U737 (N_737,N_672,N_692);
or U738 (N_738,N_687,N_665);
or U739 (N_739,N_672,N_679);
and U740 (N_740,N_657,N_686);
nand U741 (N_741,N_665,N_699);
and U742 (N_742,N_656,N_688);
nor U743 (N_743,N_679,N_665);
nor U744 (N_744,N_674,N_675);
and U745 (N_745,N_653,N_688);
or U746 (N_746,N_682,N_686);
and U747 (N_747,N_652,N_685);
nor U748 (N_748,N_661,N_671);
and U749 (N_749,N_654,N_688);
and U750 (N_750,N_730,N_706);
nor U751 (N_751,N_711,N_713);
nand U752 (N_752,N_701,N_700);
nand U753 (N_753,N_709,N_714);
and U754 (N_754,N_745,N_728);
and U755 (N_755,N_723,N_704);
nand U756 (N_756,N_720,N_719);
nor U757 (N_757,N_712,N_739);
nand U758 (N_758,N_717,N_705);
nor U759 (N_759,N_727,N_716);
and U760 (N_760,N_748,N_725);
nor U761 (N_761,N_715,N_743);
and U762 (N_762,N_735,N_703);
and U763 (N_763,N_724,N_736);
and U764 (N_764,N_741,N_738);
nand U765 (N_765,N_710,N_734);
nand U766 (N_766,N_742,N_726);
or U767 (N_767,N_737,N_749);
nand U768 (N_768,N_731,N_740);
nor U769 (N_769,N_721,N_718);
or U770 (N_770,N_708,N_702);
nor U771 (N_771,N_722,N_733);
nand U772 (N_772,N_747,N_707);
or U773 (N_773,N_732,N_729);
nor U774 (N_774,N_746,N_744);
nand U775 (N_775,N_723,N_736);
and U776 (N_776,N_714,N_700);
and U777 (N_777,N_740,N_748);
nand U778 (N_778,N_743,N_724);
or U779 (N_779,N_730,N_731);
or U780 (N_780,N_748,N_729);
and U781 (N_781,N_706,N_724);
nand U782 (N_782,N_721,N_708);
nand U783 (N_783,N_705,N_715);
nor U784 (N_784,N_740,N_746);
and U785 (N_785,N_717,N_744);
or U786 (N_786,N_715,N_734);
or U787 (N_787,N_717,N_732);
and U788 (N_788,N_745,N_742);
or U789 (N_789,N_734,N_720);
nor U790 (N_790,N_737,N_720);
nor U791 (N_791,N_734,N_748);
or U792 (N_792,N_738,N_742);
and U793 (N_793,N_749,N_720);
nor U794 (N_794,N_732,N_747);
nand U795 (N_795,N_746,N_728);
nor U796 (N_796,N_741,N_740);
and U797 (N_797,N_724,N_716);
and U798 (N_798,N_726,N_715);
and U799 (N_799,N_742,N_729);
nand U800 (N_800,N_750,N_778);
nand U801 (N_801,N_755,N_773);
nor U802 (N_802,N_775,N_764);
and U803 (N_803,N_758,N_753);
or U804 (N_804,N_788,N_782);
or U805 (N_805,N_767,N_791);
and U806 (N_806,N_766,N_781);
and U807 (N_807,N_754,N_769);
or U808 (N_808,N_784,N_787);
or U809 (N_809,N_771,N_797);
nand U810 (N_810,N_779,N_770);
and U811 (N_811,N_776,N_763);
or U812 (N_812,N_757,N_794);
or U813 (N_813,N_792,N_789);
nor U814 (N_814,N_756,N_772);
or U815 (N_815,N_777,N_761);
and U816 (N_816,N_793,N_759);
nor U817 (N_817,N_751,N_799);
and U818 (N_818,N_786,N_752);
nand U819 (N_819,N_796,N_762);
or U820 (N_820,N_785,N_765);
or U821 (N_821,N_795,N_790);
nor U822 (N_822,N_774,N_780);
and U823 (N_823,N_768,N_798);
nor U824 (N_824,N_783,N_760);
nor U825 (N_825,N_759,N_756);
nor U826 (N_826,N_793,N_790);
or U827 (N_827,N_789,N_777);
and U828 (N_828,N_764,N_752);
and U829 (N_829,N_789,N_760);
and U830 (N_830,N_759,N_753);
nor U831 (N_831,N_785,N_774);
nand U832 (N_832,N_761,N_793);
nor U833 (N_833,N_758,N_789);
or U834 (N_834,N_764,N_788);
nand U835 (N_835,N_781,N_750);
nand U836 (N_836,N_755,N_790);
nand U837 (N_837,N_799,N_784);
nor U838 (N_838,N_772,N_788);
or U839 (N_839,N_753,N_797);
or U840 (N_840,N_797,N_799);
and U841 (N_841,N_783,N_768);
and U842 (N_842,N_756,N_779);
nor U843 (N_843,N_762,N_779);
nor U844 (N_844,N_783,N_797);
nor U845 (N_845,N_795,N_760);
or U846 (N_846,N_768,N_782);
xor U847 (N_847,N_768,N_769);
and U848 (N_848,N_754,N_777);
and U849 (N_849,N_777,N_763);
nor U850 (N_850,N_812,N_834);
nand U851 (N_851,N_802,N_805);
and U852 (N_852,N_818,N_800);
and U853 (N_853,N_836,N_822);
nor U854 (N_854,N_811,N_821);
nand U855 (N_855,N_801,N_823);
nand U856 (N_856,N_826,N_815);
and U857 (N_857,N_843,N_808);
and U858 (N_858,N_831,N_806);
xnor U859 (N_859,N_814,N_829);
and U860 (N_860,N_824,N_841);
and U861 (N_861,N_832,N_827);
or U862 (N_862,N_848,N_849);
nand U863 (N_863,N_816,N_830);
or U864 (N_864,N_819,N_845);
nand U865 (N_865,N_813,N_820);
and U866 (N_866,N_803,N_844);
nor U867 (N_867,N_809,N_817);
and U868 (N_868,N_847,N_810);
or U869 (N_869,N_840,N_825);
xnor U870 (N_870,N_807,N_838);
nand U871 (N_871,N_828,N_839);
and U872 (N_872,N_835,N_833);
or U873 (N_873,N_846,N_842);
nor U874 (N_874,N_837,N_804);
nor U875 (N_875,N_823,N_835);
or U876 (N_876,N_817,N_807);
or U877 (N_877,N_839,N_826);
xnor U878 (N_878,N_844,N_832);
nand U879 (N_879,N_830,N_807);
or U880 (N_880,N_844,N_828);
nor U881 (N_881,N_839,N_848);
nor U882 (N_882,N_848,N_822);
xor U883 (N_883,N_811,N_826);
or U884 (N_884,N_841,N_835);
nand U885 (N_885,N_843,N_831);
and U886 (N_886,N_816,N_833);
and U887 (N_887,N_804,N_807);
nand U888 (N_888,N_821,N_845);
nor U889 (N_889,N_848,N_802);
and U890 (N_890,N_817,N_801);
nor U891 (N_891,N_847,N_817);
nor U892 (N_892,N_816,N_811);
and U893 (N_893,N_823,N_840);
and U894 (N_894,N_804,N_841);
or U895 (N_895,N_837,N_836);
and U896 (N_896,N_839,N_801);
nand U897 (N_897,N_830,N_822);
nor U898 (N_898,N_812,N_811);
or U899 (N_899,N_848,N_816);
or U900 (N_900,N_875,N_887);
nand U901 (N_901,N_895,N_854);
nand U902 (N_902,N_859,N_876);
or U903 (N_903,N_860,N_871);
and U904 (N_904,N_889,N_851);
or U905 (N_905,N_862,N_890);
nand U906 (N_906,N_899,N_884);
or U907 (N_907,N_865,N_852);
nand U908 (N_908,N_885,N_866);
nor U909 (N_909,N_867,N_864);
nor U910 (N_910,N_880,N_869);
nor U911 (N_911,N_898,N_870);
xor U912 (N_912,N_856,N_874);
nor U913 (N_913,N_897,N_893);
or U914 (N_914,N_888,N_873);
nor U915 (N_915,N_853,N_892);
and U916 (N_916,N_879,N_850);
and U917 (N_917,N_878,N_877);
nor U918 (N_918,N_894,N_868);
and U919 (N_919,N_896,N_857);
and U920 (N_920,N_855,N_858);
nor U921 (N_921,N_886,N_882);
nand U922 (N_922,N_881,N_863);
nand U923 (N_923,N_883,N_861);
and U924 (N_924,N_872,N_891);
nor U925 (N_925,N_896,N_875);
nor U926 (N_926,N_877,N_890);
nand U927 (N_927,N_880,N_867);
or U928 (N_928,N_851,N_883);
nor U929 (N_929,N_860,N_875);
nor U930 (N_930,N_857,N_864);
nor U931 (N_931,N_897,N_877);
or U932 (N_932,N_887,N_872);
nand U933 (N_933,N_870,N_852);
nand U934 (N_934,N_862,N_865);
or U935 (N_935,N_875,N_851);
and U936 (N_936,N_891,N_871);
nor U937 (N_937,N_851,N_888);
and U938 (N_938,N_898,N_895);
or U939 (N_939,N_874,N_881);
or U940 (N_940,N_855,N_896);
and U941 (N_941,N_860,N_883);
or U942 (N_942,N_854,N_885);
nand U943 (N_943,N_899,N_878);
nand U944 (N_944,N_864,N_856);
nor U945 (N_945,N_851,N_873);
and U946 (N_946,N_886,N_862);
and U947 (N_947,N_875,N_856);
nor U948 (N_948,N_861,N_877);
nor U949 (N_949,N_851,N_876);
xnor U950 (N_950,N_918,N_946);
or U951 (N_951,N_942,N_944);
and U952 (N_952,N_904,N_912);
nor U953 (N_953,N_949,N_929);
nor U954 (N_954,N_938,N_931);
nor U955 (N_955,N_941,N_907);
or U956 (N_956,N_935,N_937);
nor U957 (N_957,N_922,N_925);
nor U958 (N_958,N_908,N_936);
and U959 (N_959,N_926,N_923);
or U960 (N_960,N_909,N_916);
nor U961 (N_961,N_948,N_947);
and U962 (N_962,N_945,N_921);
or U963 (N_963,N_920,N_911);
nand U964 (N_964,N_905,N_934);
nor U965 (N_965,N_900,N_940);
nand U966 (N_966,N_927,N_902);
and U967 (N_967,N_903,N_939);
nand U968 (N_968,N_913,N_915);
nand U969 (N_969,N_914,N_932);
or U970 (N_970,N_917,N_901);
nand U971 (N_971,N_906,N_943);
nor U972 (N_972,N_928,N_910);
nor U973 (N_973,N_930,N_933);
nand U974 (N_974,N_919,N_924);
nor U975 (N_975,N_924,N_947);
nor U976 (N_976,N_904,N_901);
nor U977 (N_977,N_919,N_906);
and U978 (N_978,N_929,N_911);
and U979 (N_979,N_925,N_900);
nor U980 (N_980,N_925,N_924);
nor U981 (N_981,N_912,N_929);
nand U982 (N_982,N_932,N_941);
nor U983 (N_983,N_931,N_906);
or U984 (N_984,N_942,N_902);
and U985 (N_985,N_925,N_944);
and U986 (N_986,N_916,N_905);
nor U987 (N_987,N_916,N_938);
nand U988 (N_988,N_904,N_939);
xnor U989 (N_989,N_913,N_940);
and U990 (N_990,N_909,N_914);
nor U991 (N_991,N_933,N_935);
nand U992 (N_992,N_942,N_910);
or U993 (N_993,N_934,N_924);
and U994 (N_994,N_942,N_940);
or U995 (N_995,N_949,N_941);
or U996 (N_996,N_932,N_905);
nor U997 (N_997,N_907,N_918);
nand U998 (N_998,N_945,N_925);
and U999 (N_999,N_942,N_922);
nor U1000 (N_1000,N_964,N_973);
nor U1001 (N_1001,N_988,N_978);
or U1002 (N_1002,N_965,N_957);
nand U1003 (N_1003,N_980,N_974);
nand U1004 (N_1004,N_958,N_977);
and U1005 (N_1005,N_963,N_966);
nand U1006 (N_1006,N_979,N_975);
nor U1007 (N_1007,N_999,N_993);
nor U1008 (N_1008,N_962,N_959);
and U1009 (N_1009,N_997,N_960);
and U1010 (N_1010,N_972,N_967);
nor U1011 (N_1011,N_970,N_994);
nand U1012 (N_1012,N_990,N_991);
nor U1013 (N_1013,N_996,N_952);
nor U1014 (N_1014,N_976,N_998);
or U1015 (N_1015,N_955,N_985);
and U1016 (N_1016,N_981,N_968);
and U1017 (N_1017,N_953,N_995);
nor U1018 (N_1018,N_954,N_969);
nand U1019 (N_1019,N_951,N_984);
and U1020 (N_1020,N_989,N_986);
nor U1021 (N_1021,N_987,N_982);
and U1022 (N_1022,N_971,N_992);
nand U1023 (N_1023,N_950,N_983);
nor U1024 (N_1024,N_961,N_956);
or U1025 (N_1025,N_979,N_969);
or U1026 (N_1026,N_961,N_971);
and U1027 (N_1027,N_985,N_970);
or U1028 (N_1028,N_976,N_959);
nor U1029 (N_1029,N_958,N_990);
or U1030 (N_1030,N_978,N_995);
or U1031 (N_1031,N_952,N_962);
or U1032 (N_1032,N_954,N_960);
or U1033 (N_1033,N_990,N_962);
and U1034 (N_1034,N_990,N_959);
or U1035 (N_1035,N_970,N_968);
nand U1036 (N_1036,N_997,N_989);
or U1037 (N_1037,N_995,N_966);
or U1038 (N_1038,N_996,N_956);
and U1039 (N_1039,N_975,N_978);
nand U1040 (N_1040,N_989,N_955);
or U1041 (N_1041,N_956,N_951);
nor U1042 (N_1042,N_971,N_957);
and U1043 (N_1043,N_970,N_952);
or U1044 (N_1044,N_981,N_969);
nand U1045 (N_1045,N_960,N_956);
nand U1046 (N_1046,N_981,N_985);
or U1047 (N_1047,N_985,N_996);
nor U1048 (N_1048,N_988,N_951);
or U1049 (N_1049,N_972,N_993);
nor U1050 (N_1050,N_1026,N_1019);
and U1051 (N_1051,N_1044,N_1007);
and U1052 (N_1052,N_1040,N_1035);
xor U1053 (N_1053,N_1025,N_1039);
or U1054 (N_1054,N_1015,N_1016);
or U1055 (N_1055,N_1048,N_1038);
and U1056 (N_1056,N_1029,N_1023);
nor U1057 (N_1057,N_1033,N_1042);
nand U1058 (N_1058,N_1028,N_1014);
nor U1059 (N_1059,N_1034,N_1013);
and U1060 (N_1060,N_1006,N_1022);
and U1061 (N_1061,N_1004,N_1020);
nor U1062 (N_1062,N_1009,N_1046);
nor U1063 (N_1063,N_1008,N_1031);
nor U1064 (N_1064,N_1018,N_1036);
nand U1065 (N_1065,N_1030,N_1012);
and U1066 (N_1066,N_1027,N_1032);
nor U1067 (N_1067,N_1041,N_1002);
or U1068 (N_1068,N_1024,N_1045);
nand U1069 (N_1069,N_1037,N_1005);
nor U1070 (N_1070,N_1011,N_1003);
or U1071 (N_1071,N_1001,N_1021);
and U1072 (N_1072,N_1049,N_1017);
nand U1073 (N_1073,N_1000,N_1010);
nor U1074 (N_1074,N_1043,N_1047);
nand U1075 (N_1075,N_1016,N_1035);
nand U1076 (N_1076,N_1045,N_1018);
nor U1077 (N_1077,N_1038,N_1005);
nand U1078 (N_1078,N_1006,N_1034);
and U1079 (N_1079,N_1027,N_1033);
nand U1080 (N_1080,N_1026,N_1015);
nand U1081 (N_1081,N_1032,N_1020);
nor U1082 (N_1082,N_1019,N_1001);
nor U1083 (N_1083,N_1024,N_1028);
nor U1084 (N_1084,N_1013,N_1016);
and U1085 (N_1085,N_1000,N_1025);
nand U1086 (N_1086,N_1040,N_1017);
xnor U1087 (N_1087,N_1045,N_1037);
and U1088 (N_1088,N_1016,N_1028);
nand U1089 (N_1089,N_1023,N_1022);
nor U1090 (N_1090,N_1020,N_1044);
and U1091 (N_1091,N_1022,N_1040);
and U1092 (N_1092,N_1001,N_1002);
or U1093 (N_1093,N_1007,N_1018);
and U1094 (N_1094,N_1007,N_1009);
nand U1095 (N_1095,N_1013,N_1049);
and U1096 (N_1096,N_1046,N_1022);
and U1097 (N_1097,N_1028,N_1029);
and U1098 (N_1098,N_1028,N_1018);
nor U1099 (N_1099,N_1022,N_1014);
nor U1100 (N_1100,N_1056,N_1095);
nor U1101 (N_1101,N_1062,N_1064);
or U1102 (N_1102,N_1075,N_1067);
nor U1103 (N_1103,N_1052,N_1058);
and U1104 (N_1104,N_1097,N_1055);
or U1105 (N_1105,N_1087,N_1094);
nor U1106 (N_1106,N_1061,N_1099);
nand U1107 (N_1107,N_1057,N_1081);
nor U1108 (N_1108,N_1059,N_1069);
nor U1109 (N_1109,N_1060,N_1090);
nor U1110 (N_1110,N_1093,N_1096);
and U1111 (N_1111,N_1065,N_1054);
nor U1112 (N_1112,N_1080,N_1070);
nand U1113 (N_1113,N_1071,N_1091);
or U1114 (N_1114,N_1053,N_1051);
and U1115 (N_1115,N_1079,N_1089);
and U1116 (N_1116,N_1074,N_1072);
nand U1117 (N_1117,N_1092,N_1084);
nor U1118 (N_1118,N_1066,N_1082);
or U1119 (N_1119,N_1063,N_1098);
and U1120 (N_1120,N_1083,N_1050);
nand U1121 (N_1121,N_1076,N_1086);
nor U1122 (N_1122,N_1068,N_1085);
nor U1123 (N_1123,N_1073,N_1078);
nor U1124 (N_1124,N_1077,N_1088);
nor U1125 (N_1125,N_1072,N_1063);
nor U1126 (N_1126,N_1061,N_1082);
nand U1127 (N_1127,N_1086,N_1077);
nand U1128 (N_1128,N_1079,N_1070);
nor U1129 (N_1129,N_1059,N_1066);
nand U1130 (N_1130,N_1078,N_1065);
xnor U1131 (N_1131,N_1053,N_1071);
nand U1132 (N_1132,N_1081,N_1071);
and U1133 (N_1133,N_1090,N_1061);
nand U1134 (N_1134,N_1070,N_1093);
and U1135 (N_1135,N_1062,N_1060);
and U1136 (N_1136,N_1075,N_1088);
or U1137 (N_1137,N_1089,N_1085);
or U1138 (N_1138,N_1067,N_1052);
and U1139 (N_1139,N_1081,N_1070);
nor U1140 (N_1140,N_1084,N_1087);
and U1141 (N_1141,N_1088,N_1096);
and U1142 (N_1142,N_1096,N_1055);
nor U1143 (N_1143,N_1079,N_1081);
or U1144 (N_1144,N_1061,N_1050);
nand U1145 (N_1145,N_1070,N_1053);
nor U1146 (N_1146,N_1070,N_1086);
nand U1147 (N_1147,N_1094,N_1095);
xnor U1148 (N_1148,N_1084,N_1098);
or U1149 (N_1149,N_1088,N_1074);
and U1150 (N_1150,N_1113,N_1119);
and U1151 (N_1151,N_1103,N_1104);
or U1152 (N_1152,N_1137,N_1115);
and U1153 (N_1153,N_1139,N_1147);
nand U1154 (N_1154,N_1126,N_1123);
and U1155 (N_1155,N_1111,N_1142);
nor U1156 (N_1156,N_1117,N_1144);
nor U1157 (N_1157,N_1118,N_1129);
nand U1158 (N_1158,N_1140,N_1125);
nor U1159 (N_1159,N_1130,N_1132);
nand U1160 (N_1160,N_1112,N_1101);
and U1161 (N_1161,N_1135,N_1100);
nor U1162 (N_1162,N_1149,N_1109);
nand U1163 (N_1163,N_1105,N_1131);
nand U1164 (N_1164,N_1127,N_1138);
nor U1165 (N_1165,N_1145,N_1146);
nor U1166 (N_1166,N_1141,N_1122);
nand U1167 (N_1167,N_1133,N_1120);
and U1168 (N_1168,N_1136,N_1143);
and U1169 (N_1169,N_1124,N_1134);
nand U1170 (N_1170,N_1116,N_1108);
and U1171 (N_1171,N_1110,N_1148);
nand U1172 (N_1172,N_1107,N_1102);
nor U1173 (N_1173,N_1121,N_1128);
or U1174 (N_1174,N_1114,N_1106);
or U1175 (N_1175,N_1112,N_1124);
nor U1176 (N_1176,N_1131,N_1113);
nor U1177 (N_1177,N_1118,N_1142);
nand U1178 (N_1178,N_1131,N_1112);
nor U1179 (N_1179,N_1109,N_1105);
or U1180 (N_1180,N_1125,N_1134);
nand U1181 (N_1181,N_1146,N_1108);
nand U1182 (N_1182,N_1126,N_1142);
or U1183 (N_1183,N_1125,N_1108);
and U1184 (N_1184,N_1118,N_1149);
or U1185 (N_1185,N_1125,N_1148);
and U1186 (N_1186,N_1106,N_1112);
nor U1187 (N_1187,N_1145,N_1102);
nand U1188 (N_1188,N_1123,N_1144);
and U1189 (N_1189,N_1147,N_1109);
nor U1190 (N_1190,N_1134,N_1145);
or U1191 (N_1191,N_1109,N_1100);
and U1192 (N_1192,N_1137,N_1116);
or U1193 (N_1193,N_1125,N_1136);
and U1194 (N_1194,N_1146,N_1116);
or U1195 (N_1195,N_1149,N_1102);
nor U1196 (N_1196,N_1132,N_1131);
nand U1197 (N_1197,N_1128,N_1126);
and U1198 (N_1198,N_1131,N_1147);
and U1199 (N_1199,N_1100,N_1146);
or U1200 (N_1200,N_1191,N_1189);
nand U1201 (N_1201,N_1161,N_1150);
nor U1202 (N_1202,N_1184,N_1156);
or U1203 (N_1203,N_1195,N_1179);
nor U1204 (N_1204,N_1171,N_1199);
nor U1205 (N_1205,N_1153,N_1196);
or U1206 (N_1206,N_1154,N_1152);
and U1207 (N_1207,N_1158,N_1185);
nor U1208 (N_1208,N_1151,N_1167);
or U1209 (N_1209,N_1198,N_1178);
or U1210 (N_1210,N_1160,N_1174);
nor U1211 (N_1211,N_1172,N_1162);
and U1212 (N_1212,N_1182,N_1176);
nor U1213 (N_1213,N_1170,N_1197);
and U1214 (N_1214,N_1177,N_1186);
and U1215 (N_1215,N_1192,N_1164);
nand U1216 (N_1216,N_1163,N_1183);
and U1217 (N_1217,N_1173,N_1159);
or U1218 (N_1218,N_1181,N_1175);
nand U1219 (N_1219,N_1194,N_1188);
nor U1220 (N_1220,N_1157,N_1193);
or U1221 (N_1221,N_1165,N_1166);
nand U1222 (N_1222,N_1187,N_1180);
nand U1223 (N_1223,N_1169,N_1155);
nand U1224 (N_1224,N_1190,N_1168);
or U1225 (N_1225,N_1184,N_1161);
or U1226 (N_1226,N_1174,N_1183);
or U1227 (N_1227,N_1168,N_1189);
xnor U1228 (N_1228,N_1198,N_1150);
nand U1229 (N_1229,N_1160,N_1170);
or U1230 (N_1230,N_1183,N_1166);
nand U1231 (N_1231,N_1194,N_1174);
nand U1232 (N_1232,N_1166,N_1169);
and U1233 (N_1233,N_1191,N_1183);
nor U1234 (N_1234,N_1193,N_1174);
nor U1235 (N_1235,N_1192,N_1154);
or U1236 (N_1236,N_1179,N_1191);
and U1237 (N_1237,N_1185,N_1166);
nand U1238 (N_1238,N_1183,N_1167);
and U1239 (N_1239,N_1182,N_1164);
nor U1240 (N_1240,N_1178,N_1169);
nand U1241 (N_1241,N_1196,N_1187);
nand U1242 (N_1242,N_1157,N_1150);
nor U1243 (N_1243,N_1167,N_1150);
and U1244 (N_1244,N_1171,N_1192);
or U1245 (N_1245,N_1154,N_1191);
nor U1246 (N_1246,N_1164,N_1184);
nor U1247 (N_1247,N_1168,N_1194);
xor U1248 (N_1248,N_1165,N_1161);
nand U1249 (N_1249,N_1164,N_1198);
and U1250 (N_1250,N_1248,N_1222);
and U1251 (N_1251,N_1244,N_1206);
or U1252 (N_1252,N_1215,N_1228);
nor U1253 (N_1253,N_1243,N_1239);
or U1254 (N_1254,N_1209,N_1210);
nand U1255 (N_1255,N_1218,N_1249);
nand U1256 (N_1256,N_1231,N_1203);
and U1257 (N_1257,N_1235,N_1225);
nand U1258 (N_1258,N_1245,N_1241);
nand U1259 (N_1259,N_1240,N_1212);
nor U1260 (N_1260,N_1204,N_1227);
nand U1261 (N_1261,N_1238,N_1200);
nor U1262 (N_1262,N_1202,N_1208);
nor U1263 (N_1263,N_1205,N_1223);
and U1264 (N_1264,N_1224,N_1219);
and U1265 (N_1265,N_1230,N_1236);
or U1266 (N_1266,N_1201,N_1211);
or U1267 (N_1267,N_1221,N_1246);
nor U1268 (N_1268,N_1216,N_1207);
nor U1269 (N_1269,N_1220,N_1233);
or U1270 (N_1270,N_1229,N_1237);
and U1271 (N_1271,N_1213,N_1234);
nand U1272 (N_1272,N_1242,N_1226);
nand U1273 (N_1273,N_1247,N_1214);
nand U1274 (N_1274,N_1217,N_1232);
nand U1275 (N_1275,N_1237,N_1230);
nand U1276 (N_1276,N_1233,N_1216);
or U1277 (N_1277,N_1221,N_1240);
or U1278 (N_1278,N_1214,N_1233);
nand U1279 (N_1279,N_1213,N_1229);
and U1280 (N_1280,N_1214,N_1220);
nor U1281 (N_1281,N_1237,N_1239);
and U1282 (N_1282,N_1232,N_1227);
or U1283 (N_1283,N_1241,N_1227);
nor U1284 (N_1284,N_1202,N_1206);
or U1285 (N_1285,N_1247,N_1210);
and U1286 (N_1286,N_1228,N_1235);
nor U1287 (N_1287,N_1236,N_1211);
and U1288 (N_1288,N_1246,N_1204);
xor U1289 (N_1289,N_1244,N_1213);
nor U1290 (N_1290,N_1219,N_1209);
or U1291 (N_1291,N_1222,N_1237);
and U1292 (N_1292,N_1206,N_1236);
and U1293 (N_1293,N_1234,N_1245);
or U1294 (N_1294,N_1249,N_1239);
and U1295 (N_1295,N_1212,N_1227);
nand U1296 (N_1296,N_1244,N_1243);
or U1297 (N_1297,N_1212,N_1221);
and U1298 (N_1298,N_1243,N_1217);
and U1299 (N_1299,N_1218,N_1208);
nand U1300 (N_1300,N_1293,N_1281);
nor U1301 (N_1301,N_1253,N_1290);
or U1302 (N_1302,N_1271,N_1251);
or U1303 (N_1303,N_1282,N_1297);
and U1304 (N_1304,N_1285,N_1259);
nor U1305 (N_1305,N_1257,N_1267);
and U1306 (N_1306,N_1280,N_1256);
and U1307 (N_1307,N_1250,N_1286);
nand U1308 (N_1308,N_1295,N_1255);
or U1309 (N_1309,N_1277,N_1269);
nor U1310 (N_1310,N_1276,N_1262);
nor U1311 (N_1311,N_1268,N_1266);
nand U1312 (N_1312,N_1299,N_1261);
nor U1313 (N_1313,N_1289,N_1263);
and U1314 (N_1314,N_1254,N_1258);
nor U1315 (N_1315,N_1265,N_1272);
nor U1316 (N_1316,N_1298,N_1291);
and U1317 (N_1317,N_1260,N_1288);
nand U1318 (N_1318,N_1274,N_1275);
nor U1319 (N_1319,N_1284,N_1287);
nor U1320 (N_1320,N_1283,N_1273);
or U1321 (N_1321,N_1270,N_1294);
and U1322 (N_1322,N_1296,N_1264);
or U1323 (N_1323,N_1252,N_1279);
nor U1324 (N_1324,N_1278,N_1292);
or U1325 (N_1325,N_1289,N_1294);
nand U1326 (N_1326,N_1260,N_1254);
and U1327 (N_1327,N_1280,N_1271);
nand U1328 (N_1328,N_1290,N_1298);
or U1329 (N_1329,N_1257,N_1281);
and U1330 (N_1330,N_1291,N_1259);
and U1331 (N_1331,N_1280,N_1285);
and U1332 (N_1332,N_1298,N_1273);
nand U1333 (N_1333,N_1289,N_1251);
or U1334 (N_1334,N_1252,N_1270);
nand U1335 (N_1335,N_1262,N_1274);
nand U1336 (N_1336,N_1256,N_1253);
or U1337 (N_1337,N_1281,N_1256);
nor U1338 (N_1338,N_1271,N_1270);
and U1339 (N_1339,N_1279,N_1272);
and U1340 (N_1340,N_1270,N_1298);
nor U1341 (N_1341,N_1278,N_1299);
or U1342 (N_1342,N_1288,N_1290);
nand U1343 (N_1343,N_1295,N_1297);
nor U1344 (N_1344,N_1269,N_1294);
nor U1345 (N_1345,N_1254,N_1291);
nand U1346 (N_1346,N_1299,N_1274);
and U1347 (N_1347,N_1253,N_1294);
and U1348 (N_1348,N_1271,N_1253);
nor U1349 (N_1349,N_1293,N_1250);
and U1350 (N_1350,N_1314,N_1347);
and U1351 (N_1351,N_1305,N_1310);
nor U1352 (N_1352,N_1315,N_1338);
and U1353 (N_1353,N_1345,N_1318);
or U1354 (N_1354,N_1321,N_1330);
or U1355 (N_1355,N_1324,N_1307);
and U1356 (N_1356,N_1302,N_1322);
and U1357 (N_1357,N_1316,N_1328);
and U1358 (N_1358,N_1313,N_1326);
or U1359 (N_1359,N_1342,N_1343);
or U1360 (N_1360,N_1300,N_1337);
or U1361 (N_1361,N_1306,N_1320);
nand U1362 (N_1362,N_1341,N_1303);
nor U1363 (N_1363,N_1344,N_1339);
nand U1364 (N_1364,N_1346,N_1340);
and U1365 (N_1365,N_1308,N_1325);
nor U1366 (N_1366,N_1312,N_1349);
and U1367 (N_1367,N_1301,N_1334);
nor U1368 (N_1368,N_1335,N_1309);
nand U1369 (N_1369,N_1332,N_1348);
nor U1370 (N_1370,N_1317,N_1327);
or U1371 (N_1371,N_1333,N_1311);
or U1372 (N_1372,N_1319,N_1323);
nor U1373 (N_1373,N_1336,N_1304);
and U1374 (N_1374,N_1331,N_1329);
and U1375 (N_1375,N_1301,N_1307);
or U1376 (N_1376,N_1321,N_1340);
nand U1377 (N_1377,N_1304,N_1321);
and U1378 (N_1378,N_1332,N_1303);
and U1379 (N_1379,N_1301,N_1339);
nor U1380 (N_1380,N_1342,N_1306);
or U1381 (N_1381,N_1316,N_1348);
and U1382 (N_1382,N_1340,N_1313);
or U1383 (N_1383,N_1338,N_1329);
nand U1384 (N_1384,N_1345,N_1306);
nor U1385 (N_1385,N_1339,N_1324);
and U1386 (N_1386,N_1323,N_1312);
and U1387 (N_1387,N_1332,N_1310);
nand U1388 (N_1388,N_1324,N_1308);
and U1389 (N_1389,N_1309,N_1315);
and U1390 (N_1390,N_1317,N_1346);
and U1391 (N_1391,N_1320,N_1330);
nor U1392 (N_1392,N_1341,N_1346);
nor U1393 (N_1393,N_1343,N_1307);
nor U1394 (N_1394,N_1300,N_1312);
or U1395 (N_1395,N_1328,N_1330);
nor U1396 (N_1396,N_1313,N_1342);
or U1397 (N_1397,N_1327,N_1337);
nand U1398 (N_1398,N_1345,N_1325);
or U1399 (N_1399,N_1342,N_1341);
or U1400 (N_1400,N_1366,N_1378);
nor U1401 (N_1401,N_1367,N_1386);
or U1402 (N_1402,N_1389,N_1374);
nor U1403 (N_1403,N_1369,N_1365);
nor U1404 (N_1404,N_1351,N_1379);
and U1405 (N_1405,N_1382,N_1354);
or U1406 (N_1406,N_1371,N_1355);
or U1407 (N_1407,N_1377,N_1391);
or U1408 (N_1408,N_1364,N_1363);
and U1409 (N_1409,N_1398,N_1380);
and U1410 (N_1410,N_1353,N_1390);
and U1411 (N_1411,N_1392,N_1357);
nand U1412 (N_1412,N_1394,N_1393);
or U1413 (N_1413,N_1387,N_1396);
or U1414 (N_1414,N_1397,N_1362);
or U1415 (N_1415,N_1399,N_1385);
and U1416 (N_1416,N_1356,N_1384);
nor U1417 (N_1417,N_1360,N_1368);
or U1418 (N_1418,N_1358,N_1359);
and U1419 (N_1419,N_1350,N_1372);
nor U1420 (N_1420,N_1381,N_1395);
nor U1421 (N_1421,N_1388,N_1383);
and U1422 (N_1422,N_1376,N_1370);
nand U1423 (N_1423,N_1352,N_1361);
nand U1424 (N_1424,N_1375,N_1373);
and U1425 (N_1425,N_1375,N_1357);
and U1426 (N_1426,N_1387,N_1379);
or U1427 (N_1427,N_1364,N_1350);
or U1428 (N_1428,N_1363,N_1357);
nor U1429 (N_1429,N_1361,N_1370);
nor U1430 (N_1430,N_1373,N_1382);
or U1431 (N_1431,N_1356,N_1392);
and U1432 (N_1432,N_1385,N_1377);
nand U1433 (N_1433,N_1378,N_1358);
nand U1434 (N_1434,N_1398,N_1354);
or U1435 (N_1435,N_1380,N_1366);
and U1436 (N_1436,N_1358,N_1366);
and U1437 (N_1437,N_1398,N_1367);
or U1438 (N_1438,N_1390,N_1374);
nand U1439 (N_1439,N_1399,N_1372);
or U1440 (N_1440,N_1398,N_1373);
nand U1441 (N_1441,N_1371,N_1383);
or U1442 (N_1442,N_1365,N_1364);
nand U1443 (N_1443,N_1383,N_1367);
or U1444 (N_1444,N_1375,N_1361);
nand U1445 (N_1445,N_1350,N_1395);
and U1446 (N_1446,N_1370,N_1363);
nor U1447 (N_1447,N_1399,N_1384);
and U1448 (N_1448,N_1382,N_1374);
or U1449 (N_1449,N_1381,N_1383);
or U1450 (N_1450,N_1417,N_1444);
or U1451 (N_1451,N_1448,N_1416);
nor U1452 (N_1452,N_1415,N_1423);
nor U1453 (N_1453,N_1428,N_1429);
or U1454 (N_1454,N_1432,N_1421);
and U1455 (N_1455,N_1441,N_1438);
and U1456 (N_1456,N_1445,N_1447);
and U1457 (N_1457,N_1401,N_1430);
nand U1458 (N_1458,N_1412,N_1400);
and U1459 (N_1459,N_1408,N_1424);
or U1460 (N_1460,N_1419,N_1405);
nor U1461 (N_1461,N_1435,N_1403);
or U1462 (N_1462,N_1411,N_1427);
or U1463 (N_1463,N_1404,N_1407);
xor U1464 (N_1464,N_1418,N_1413);
or U1465 (N_1465,N_1439,N_1437);
or U1466 (N_1466,N_1414,N_1409);
nand U1467 (N_1467,N_1431,N_1446);
or U1468 (N_1468,N_1449,N_1420);
nor U1469 (N_1469,N_1433,N_1434);
nand U1470 (N_1470,N_1422,N_1406);
and U1471 (N_1471,N_1440,N_1426);
nand U1472 (N_1472,N_1436,N_1443);
and U1473 (N_1473,N_1410,N_1402);
nand U1474 (N_1474,N_1442,N_1425);
or U1475 (N_1475,N_1401,N_1420);
nand U1476 (N_1476,N_1407,N_1439);
xnor U1477 (N_1477,N_1412,N_1420);
and U1478 (N_1478,N_1447,N_1402);
nand U1479 (N_1479,N_1430,N_1409);
or U1480 (N_1480,N_1411,N_1438);
nand U1481 (N_1481,N_1445,N_1422);
nand U1482 (N_1482,N_1413,N_1404);
nor U1483 (N_1483,N_1416,N_1400);
nand U1484 (N_1484,N_1446,N_1427);
nand U1485 (N_1485,N_1415,N_1448);
nand U1486 (N_1486,N_1422,N_1446);
nor U1487 (N_1487,N_1408,N_1409);
or U1488 (N_1488,N_1415,N_1416);
nand U1489 (N_1489,N_1447,N_1420);
or U1490 (N_1490,N_1407,N_1427);
and U1491 (N_1491,N_1423,N_1435);
nand U1492 (N_1492,N_1410,N_1426);
nor U1493 (N_1493,N_1411,N_1446);
and U1494 (N_1494,N_1442,N_1427);
nor U1495 (N_1495,N_1429,N_1400);
nor U1496 (N_1496,N_1408,N_1447);
or U1497 (N_1497,N_1447,N_1404);
nor U1498 (N_1498,N_1401,N_1425);
or U1499 (N_1499,N_1401,N_1424);
and U1500 (N_1500,N_1470,N_1489);
nand U1501 (N_1501,N_1461,N_1487);
nand U1502 (N_1502,N_1485,N_1466);
nor U1503 (N_1503,N_1491,N_1468);
or U1504 (N_1504,N_1467,N_1475);
nand U1505 (N_1505,N_1452,N_1450);
and U1506 (N_1506,N_1497,N_1492);
and U1507 (N_1507,N_1472,N_1499);
or U1508 (N_1508,N_1481,N_1458);
and U1509 (N_1509,N_1465,N_1496);
nand U1510 (N_1510,N_1488,N_1484);
nor U1511 (N_1511,N_1456,N_1495);
or U1512 (N_1512,N_1476,N_1483);
nor U1513 (N_1513,N_1474,N_1459);
nor U1514 (N_1514,N_1473,N_1460);
nor U1515 (N_1515,N_1453,N_1469);
and U1516 (N_1516,N_1480,N_1479);
nand U1517 (N_1517,N_1478,N_1454);
nand U1518 (N_1518,N_1451,N_1490);
or U1519 (N_1519,N_1494,N_1493);
nor U1520 (N_1520,N_1462,N_1477);
nor U1521 (N_1521,N_1486,N_1498);
nor U1522 (N_1522,N_1463,N_1471);
or U1523 (N_1523,N_1457,N_1464);
and U1524 (N_1524,N_1455,N_1482);
nand U1525 (N_1525,N_1462,N_1480);
nor U1526 (N_1526,N_1456,N_1499);
or U1527 (N_1527,N_1476,N_1467);
or U1528 (N_1528,N_1486,N_1469);
nand U1529 (N_1529,N_1476,N_1494);
and U1530 (N_1530,N_1451,N_1494);
or U1531 (N_1531,N_1459,N_1497);
or U1532 (N_1532,N_1497,N_1487);
and U1533 (N_1533,N_1453,N_1455);
and U1534 (N_1534,N_1471,N_1481);
and U1535 (N_1535,N_1493,N_1498);
nand U1536 (N_1536,N_1492,N_1475);
and U1537 (N_1537,N_1450,N_1460);
nand U1538 (N_1538,N_1467,N_1451);
nor U1539 (N_1539,N_1496,N_1495);
and U1540 (N_1540,N_1479,N_1459);
nor U1541 (N_1541,N_1471,N_1496);
or U1542 (N_1542,N_1472,N_1489);
nand U1543 (N_1543,N_1487,N_1459);
and U1544 (N_1544,N_1486,N_1489);
and U1545 (N_1545,N_1452,N_1458);
nand U1546 (N_1546,N_1479,N_1458);
or U1547 (N_1547,N_1456,N_1472);
or U1548 (N_1548,N_1484,N_1483);
nor U1549 (N_1549,N_1455,N_1460);
and U1550 (N_1550,N_1533,N_1542);
xnor U1551 (N_1551,N_1518,N_1543);
and U1552 (N_1552,N_1536,N_1537);
nor U1553 (N_1553,N_1547,N_1548);
nor U1554 (N_1554,N_1511,N_1549);
nor U1555 (N_1555,N_1535,N_1546);
nand U1556 (N_1556,N_1508,N_1509);
nor U1557 (N_1557,N_1514,N_1503);
nand U1558 (N_1558,N_1510,N_1522);
nor U1559 (N_1559,N_1527,N_1529);
nor U1560 (N_1560,N_1519,N_1525);
nand U1561 (N_1561,N_1501,N_1526);
or U1562 (N_1562,N_1539,N_1515);
nand U1563 (N_1563,N_1524,N_1506);
nor U1564 (N_1564,N_1534,N_1544);
nand U1565 (N_1565,N_1512,N_1520);
nand U1566 (N_1566,N_1523,N_1532);
nand U1567 (N_1567,N_1530,N_1504);
or U1568 (N_1568,N_1540,N_1507);
or U1569 (N_1569,N_1531,N_1541);
nand U1570 (N_1570,N_1505,N_1517);
nand U1571 (N_1571,N_1502,N_1545);
nand U1572 (N_1572,N_1500,N_1513);
nand U1573 (N_1573,N_1528,N_1516);
nor U1574 (N_1574,N_1538,N_1521);
nor U1575 (N_1575,N_1509,N_1500);
nand U1576 (N_1576,N_1522,N_1506);
nor U1577 (N_1577,N_1532,N_1513);
and U1578 (N_1578,N_1541,N_1525);
or U1579 (N_1579,N_1544,N_1516);
nor U1580 (N_1580,N_1512,N_1505);
nand U1581 (N_1581,N_1527,N_1512);
nor U1582 (N_1582,N_1545,N_1542);
and U1583 (N_1583,N_1507,N_1536);
or U1584 (N_1584,N_1544,N_1519);
nor U1585 (N_1585,N_1526,N_1545);
and U1586 (N_1586,N_1535,N_1518);
or U1587 (N_1587,N_1523,N_1540);
or U1588 (N_1588,N_1505,N_1540);
nand U1589 (N_1589,N_1503,N_1518);
nor U1590 (N_1590,N_1545,N_1524);
or U1591 (N_1591,N_1502,N_1504);
nand U1592 (N_1592,N_1516,N_1521);
nand U1593 (N_1593,N_1521,N_1522);
and U1594 (N_1594,N_1541,N_1545);
nor U1595 (N_1595,N_1527,N_1510);
and U1596 (N_1596,N_1522,N_1513);
nor U1597 (N_1597,N_1517,N_1501);
nor U1598 (N_1598,N_1504,N_1532);
nand U1599 (N_1599,N_1549,N_1522);
nor U1600 (N_1600,N_1583,N_1588);
and U1601 (N_1601,N_1594,N_1565);
and U1602 (N_1602,N_1597,N_1560);
and U1603 (N_1603,N_1592,N_1571);
nand U1604 (N_1604,N_1558,N_1575);
or U1605 (N_1605,N_1564,N_1585);
nand U1606 (N_1606,N_1595,N_1578);
nand U1607 (N_1607,N_1557,N_1580);
nor U1608 (N_1608,N_1599,N_1589);
nand U1609 (N_1609,N_1573,N_1551);
nand U1610 (N_1610,N_1587,N_1581);
nand U1611 (N_1611,N_1591,N_1563);
nand U1612 (N_1612,N_1568,N_1596);
nor U1613 (N_1613,N_1598,N_1554);
nand U1614 (N_1614,N_1590,N_1561);
and U1615 (N_1615,N_1593,N_1566);
or U1616 (N_1616,N_1550,N_1586);
or U1617 (N_1617,N_1579,N_1572);
and U1618 (N_1618,N_1556,N_1555);
or U1619 (N_1619,N_1552,N_1574);
nand U1620 (N_1620,N_1569,N_1567);
nand U1621 (N_1621,N_1553,N_1584);
or U1622 (N_1622,N_1582,N_1577);
or U1623 (N_1623,N_1576,N_1570);
and U1624 (N_1624,N_1559,N_1562);
nand U1625 (N_1625,N_1554,N_1571);
nor U1626 (N_1626,N_1569,N_1555);
nand U1627 (N_1627,N_1566,N_1550);
nand U1628 (N_1628,N_1557,N_1559);
nor U1629 (N_1629,N_1583,N_1591);
nor U1630 (N_1630,N_1560,N_1582);
nand U1631 (N_1631,N_1591,N_1593);
or U1632 (N_1632,N_1550,N_1556);
nor U1633 (N_1633,N_1564,N_1570);
nor U1634 (N_1634,N_1577,N_1563);
and U1635 (N_1635,N_1589,N_1579);
or U1636 (N_1636,N_1591,N_1598);
or U1637 (N_1637,N_1578,N_1591);
nor U1638 (N_1638,N_1584,N_1574);
nand U1639 (N_1639,N_1592,N_1552);
and U1640 (N_1640,N_1578,N_1580);
nand U1641 (N_1641,N_1572,N_1565);
nand U1642 (N_1642,N_1556,N_1553);
nand U1643 (N_1643,N_1576,N_1569);
nand U1644 (N_1644,N_1566,N_1570);
or U1645 (N_1645,N_1562,N_1596);
and U1646 (N_1646,N_1562,N_1558);
or U1647 (N_1647,N_1554,N_1595);
and U1648 (N_1648,N_1561,N_1567);
or U1649 (N_1649,N_1556,N_1594);
and U1650 (N_1650,N_1635,N_1606);
nor U1651 (N_1651,N_1633,N_1637);
nor U1652 (N_1652,N_1639,N_1632);
and U1653 (N_1653,N_1646,N_1630);
and U1654 (N_1654,N_1626,N_1631);
and U1655 (N_1655,N_1634,N_1625);
nor U1656 (N_1656,N_1618,N_1605);
or U1657 (N_1657,N_1645,N_1607);
nor U1658 (N_1658,N_1610,N_1624);
nor U1659 (N_1659,N_1615,N_1614);
and U1660 (N_1660,N_1629,N_1622);
nor U1661 (N_1661,N_1636,N_1600);
nor U1662 (N_1662,N_1613,N_1619);
nand U1663 (N_1663,N_1612,N_1621);
or U1664 (N_1664,N_1647,N_1604);
and U1665 (N_1665,N_1623,N_1609);
and U1666 (N_1666,N_1648,N_1641);
nand U1667 (N_1667,N_1628,N_1644);
nor U1668 (N_1668,N_1601,N_1611);
and U1669 (N_1669,N_1640,N_1617);
or U1670 (N_1670,N_1642,N_1649);
and U1671 (N_1671,N_1616,N_1643);
or U1672 (N_1672,N_1603,N_1608);
nand U1673 (N_1673,N_1638,N_1602);
nand U1674 (N_1674,N_1620,N_1627);
and U1675 (N_1675,N_1610,N_1632);
or U1676 (N_1676,N_1630,N_1609);
and U1677 (N_1677,N_1620,N_1606);
nor U1678 (N_1678,N_1643,N_1605);
nand U1679 (N_1679,N_1600,N_1644);
nand U1680 (N_1680,N_1618,N_1640);
and U1681 (N_1681,N_1644,N_1639);
nand U1682 (N_1682,N_1619,N_1611);
nand U1683 (N_1683,N_1607,N_1628);
nor U1684 (N_1684,N_1627,N_1640);
nand U1685 (N_1685,N_1625,N_1644);
or U1686 (N_1686,N_1606,N_1625);
nor U1687 (N_1687,N_1630,N_1611);
nor U1688 (N_1688,N_1631,N_1639);
nor U1689 (N_1689,N_1624,N_1628);
or U1690 (N_1690,N_1620,N_1638);
nand U1691 (N_1691,N_1604,N_1613);
or U1692 (N_1692,N_1603,N_1604);
nand U1693 (N_1693,N_1604,N_1630);
nand U1694 (N_1694,N_1626,N_1643);
or U1695 (N_1695,N_1616,N_1621);
or U1696 (N_1696,N_1619,N_1601);
and U1697 (N_1697,N_1632,N_1647);
nand U1698 (N_1698,N_1603,N_1617);
and U1699 (N_1699,N_1628,N_1618);
nand U1700 (N_1700,N_1698,N_1675);
and U1701 (N_1701,N_1650,N_1697);
or U1702 (N_1702,N_1687,N_1685);
and U1703 (N_1703,N_1654,N_1663);
nor U1704 (N_1704,N_1695,N_1691);
nor U1705 (N_1705,N_1688,N_1673);
xor U1706 (N_1706,N_1668,N_1669);
nand U1707 (N_1707,N_1689,N_1682);
or U1708 (N_1708,N_1660,N_1656);
nor U1709 (N_1709,N_1670,N_1690);
or U1710 (N_1710,N_1665,N_1684);
nand U1711 (N_1711,N_1672,N_1651);
nand U1712 (N_1712,N_1699,N_1658);
nand U1713 (N_1713,N_1676,N_1666);
and U1714 (N_1714,N_1678,N_1674);
and U1715 (N_1715,N_1693,N_1680);
or U1716 (N_1716,N_1694,N_1664);
nand U1717 (N_1717,N_1661,N_1657);
nor U1718 (N_1718,N_1692,N_1653);
and U1719 (N_1719,N_1686,N_1679);
nand U1720 (N_1720,N_1662,N_1681);
or U1721 (N_1721,N_1683,N_1667);
nor U1722 (N_1722,N_1659,N_1677);
xor U1723 (N_1723,N_1652,N_1696);
or U1724 (N_1724,N_1655,N_1671);
and U1725 (N_1725,N_1670,N_1668);
or U1726 (N_1726,N_1654,N_1689);
nor U1727 (N_1727,N_1698,N_1669);
nor U1728 (N_1728,N_1679,N_1666);
nor U1729 (N_1729,N_1691,N_1699);
and U1730 (N_1730,N_1698,N_1666);
nor U1731 (N_1731,N_1669,N_1688);
or U1732 (N_1732,N_1674,N_1676);
and U1733 (N_1733,N_1689,N_1681);
nand U1734 (N_1734,N_1663,N_1684);
nand U1735 (N_1735,N_1686,N_1660);
nand U1736 (N_1736,N_1681,N_1670);
and U1737 (N_1737,N_1653,N_1677);
or U1738 (N_1738,N_1694,N_1665);
nand U1739 (N_1739,N_1670,N_1666);
and U1740 (N_1740,N_1663,N_1681);
and U1741 (N_1741,N_1668,N_1689);
nor U1742 (N_1742,N_1692,N_1655);
or U1743 (N_1743,N_1670,N_1688);
or U1744 (N_1744,N_1673,N_1658);
nand U1745 (N_1745,N_1662,N_1690);
and U1746 (N_1746,N_1693,N_1679);
or U1747 (N_1747,N_1687,N_1659);
nor U1748 (N_1748,N_1686,N_1685);
and U1749 (N_1749,N_1673,N_1698);
xor U1750 (N_1750,N_1734,N_1736);
and U1751 (N_1751,N_1701,N_1740);
nor U1752 (N_1752,N_1712,N_1721);
nand U1753 (N_1753,N_1724,N_1749);
or U1754 (N_1754,N_1716,N_1703);
or U1755 (N_1755,N_1746,N_1726);
and U1756 (N_1756,N_1748,N_1717);
and U1757 (N_1757,N_1743,N_1727);
and U1758 (N_1758,N_1733,N_1729);
or U1759 (N_1759,N_1745,N_1728);
nand U1760 (N_1760,N_1718,N_1702);
and U1761 (N_1761,N_1720,N_1742);
and U1762 (N_1762,N_1708,N_1738);
nand U1763 (N_1763,N_1710,N_1700);
nor U1764 (N_1764,N_1719,N_1705);
xnor U1765 (N_1765,N_1709,N_1713);
and U1766 (N_1766,N_1741,N_1731);
nand U1767 (N_1767,N_1730,N_1737);
nor U1768 (N_1768,N_1706,N_1722);
nand U1769 (N_1769,N_1735,N_1715);
and U1770 (N_1770,N_1732,N_1714);
or U1771 (N_1771,N_1707,N_1704);
nor U1772 (N_1772,N_1711,N_1747);
nor U1773 (N_1773,N_1723,N_1725);
nand U1774 (N_1774,N_1744,N_1739);
nand U1775 (N_1775,N_1747,N_1707);
nor U1776 (N_1776,N_1710,N_1732);
or U1777 (N_1777,N_1730,N_1746);
nand U1778 (N_1778,N_1724,N_1714);
nand U1779 (N_1779,N_1708,N_1748);
nor U1780 (N_1780,N_1700,N_1724);
and U1781 (N_1781,N_1715,N_1744);
nor U1782 (N_1782,N_1732,N_1702);
nand U1783 (N_1783,N_1749,N_1747);
nand U1784 (N_1784,N_1734,N_1707);
nor U1785 (N_1785,N_1743,N_1742);
or U1786 (N_1786,N_1723,N_1747);
nand U1787 (N_1787,N_1742,N_1725);
nand U1788 (N_1788,N_1725,N_1709);
and U1789 (N_1789,N_1724,N_1740);
nor U1790 (N_1790,N_1711,N_1740);
and U1791 (N_1791,N_1713,N_1747);
or U1792 (N_1792,N_1707,N_1737);
nand U1793 (N_1793,N_1735,N_1746);
or U1794 (N_1794,N_1739,N_1741);
and U1795 (N_1795,N_1729,N_1749);
nor U1796 (N_1796,N_1707,N_1744);
or U1797 (N_1797,N_1721,N_1737);
nor U1798 (N_1798,N_1744,N_1735);
nand U1799 (N_1799,N_1724,N_1717);
and U1800 (N_1800,N_1773,N_1777);
and U1801 (N_1801,N_1757,N_1750);
or U1802 (N_1802,N_1778,N_1755);
nand U1803 (N_1803,N_1752,N_1761);
and U1804 (N_1804,N_1771,N_1791);
or U1805 (N_1805,N_1786,N_1758);
nor U1806 (N_1806,N_1782,N_1764);
and U1807 (N_1807,N_1790,N_1769);
xnor U1808 (N_1808,N_1793,N_1797);
nand U1809 (N_1809,N_1774,N_1775);
nor U1810 (N_1810,N_1770,N_1785);
and U1811 (N_1811,N_1766,N_1763);
nor U1812 (N_1812,N_1772,N_1779);
nor U1813 (N_1813,N_1780,N_1796);
nor U1814 (N_1814,N_1783,N_1754);
nor U1815 (N_1815,N_1781,N_1756);
nand U1816 (N_1816,N_1776,N_1789);
and U1817 (N_1817,N_1788,N_1798);
and U1818 (N_1818,N_1768,N_1759);
and U1819 (N_1819,N_1762,N_1760);
or U1820 (N_1820,N_1792,N_1794);
nor U1821 (N_1821,N_1795,N_1765);
nor U1822 (N_1822,N_1751,N_1799);
nand U1823 (N_1823,N_1767,N_1784);
and U1824 (N_1824,N_1787,N_1753);
nor U1825 (N_1825,N_1767,N_1769);
or U1826 (N_1826,N_1774,N_1755);
xnor U1827 (N_1827,N_1780,N_1776);
and U1828 (N_1828,N_1779,N_1773);
or U1829 (N_1829,N_1762,N_1761);
nand U1830 (N_1830,N_1762,N_1768);
or U1831 (N_1831,N_1780,N_1763);
or U1832 (N_1832,N_1762,N_1763);
nor U1833 (N_1833,N_1767,N_1779);
nand U1834 (N_1834,N_1790,N_1773);
nor U1835 (N_1835,N_1774,N_1780);
nor U1836 (N_1836,N_1796,N_1787);
nor U1837 (N_1837,N_1756,N_1778);
or U1838 (N_1838,N_1791,N_1759);
nor U1839 (N_1839,N_1794,N_1760);
nor U1840 (N_1840,N_1759,N_1750);
nand U1841 (N_1841,N_1770,N_1784);
nor U1842 (N_1842,N_1750,N_1764);
nor U1843 (N_1843,N_1756,N_1761);
nor U1844 (N_1844,N_1784,N_1797);
xnor U1845 (N_1845,N_1773,N_1758);
nand U1846 (N_1846,N_1758,N_1765);
nor U1847 (N_1847,N_1757,N_1796);
and U1848 (N_1848,N_1769,N_1758);
nor U1849 (N_1849,N_1776,N_1795);
or U1850 (N_1850,N_1802,N_1845);
nand U1851 (N_1851,N_1829,N_1849);
nand U1852 (N_1852,N_1832,N_1839);
or U1853 (N_1853,N_1840,N_1814);
nor U1854 (N_1854,N_1827,N_1844);
and U1855 (N_1855,N_1841,N_1825);
nand U1856 (N_1856,N_1817,N_1836);
and U1857 (N_1857,N_1822,N_1815);
nand U1858 (N_1858,N_1820,N_1821);
nor U1859 (N_1859,N_1810,N_1800);
nand U1860 (N_1860,N_1842,N_1805);
and U1861 (N_1861,N_1834,N_1813);
nand U1862 (N_1862,N_1835,N_1809);
nand U1863 (N_1863,N_1848,N_1804);
nand U1864 (N_1864,N_1837,N_1846);
and U1865 (N_1865,N_1816,N_1843);
and U1866 (N_1866,N_1818,N_1812);
or U1867 (N_1867,N_1823,N_1847);
nand U1868 (N_1868,N_1830,N_1808);
and U1869 (N_1869,N_1819,N_1801);
and U1870 (N_1870,N_1838,N_1833);
nor U1871 (N_1871,N_1826,N_1806);
nor U1872 (N_1872,N_1811,N_1824);
and U1873 (N_1873,N_1807,N_1803);
nor U1874 (N_1874,N_1828,N_1831);
or U1875 (N_1875,N_1849,N_1811);
nor U1876 (N_1876,N_1835,N_1840);
nand U1877 (N_1877,N_1838,N_1819);
or U1878 (N_1878,N_1821,N_1847);
and U1879 (N_1879,N_1826,N_1814);
or U1880 (N_1880,N_1810,N_1841);
or U1881 (N_1881,N_1846,N_1814);
and U1882 (N_1882,N_1827,N_1840);
nand U1883 (N_1883,N_1819,N_1837);
or U1884 (N_1884,N_1811,N_1833);
or U1885 (N_1885,N_1829,N_1815);
or U1886 (N_1886,N_1847,N_1846);
nor U1887 (N_1887,N_1800,N_1846);
nor U1888 (N_1888,N_1807,N_1815);
nand U1889 (N_1889,N_1832,N_1819);
and U1890 (N_1890,N_1805,N_1823);
nor U1891 (N_1891,N_1808,N_1840);
or U1892 (N_1892,N_1836,N_1804);
and U1893 (N_1893,N_1829,N_1802);
or U1894 (N_1894,N_1834,N_1824);
and U1895 (N_1895,N_1800,N_1811);
nor U1896 (N_1896,N_1845,N_1833);
nand U1897 (N_1897,N_1841,N_1823);
and U1898 (N_1898,N_1817,N_1818);
or U1899 (N_1899,N_1847,N_1814);
nor U1900 (N_1900,N_1863,N_1873);
or U1901 (N_1901,N_1884,N_1874);
nand U1902 (N_1902,N_1867,N_1885);
and U1903 (N_1903,N_1864,N_1889);
and U1904 (N_1904,N_1877,N_1865);
nor U1905 (N_1905,N_1876,N_1859);
and U1906 (N_1906,N_1897,N_1891);
nor U1907 (N_1907,N_1853,N_1866);
nand U1908 (N_1908,N_1881,N_1898);
nand U1909 (N_1909,N_1890,N_1883);
nand U1910 (N_1910,N_1882,N_1869);
nor U1911 (N_1911,N_1879,N_1851);
and U1912 (N_1912,N_1862,N_1895);
nor U1913 (N_1913,N_1896,N_1892);
nor U1914 (N_1914,N_1857,N_1886);
and U1915 (N_1915,N_1852,N_1887);
and U1916 (N_1916,N_1875,N_1868);
and U1917 (N_1917,N_1888,N_1854);
or U1918 (N_1918,N_1850,N_1894);
or U1919 (N_1919,N_1871,N_1878);
or U1920 (N_1920,N_1855,N_1860);
or U1921 (N_1921,N_1870,N_1899);
or U1922 (N_1922,N_1893,N_1872);
or U1923 (N_1923,N_1856,N_1858);
and U1924 (N_1924,N_1880,N_1861);
or U1925 (N_1925,N_1893,N_1856);
and U1926 (N_1926,N_1850,N_1870);
and U1927 (N_1927,N_1866,N_1875);
and U1928 (N_1928,N_1872,N_1896);
nor U1929 (N_1929,N_1895,N_1897);
nor U1930 (N_1930,N_1883,N_1884);
nor U1931 (N_1931,N_1884,N_1886);
nand U1932 (N_1932,N_1861,N_1860);
or U1933 (N_1933,N_1860,N_1882);
or U1934 (N_1934,N_1895,N_1892);
and U1935 (N_1935,N_1856,N_1851);
and U1936 (N_1936,N_1866,N_1890);
and U1937 (N_1937,N_1862,N_1855);
or U1938 (N_1938,N_1853,N_1877);
nor U1939 (N_1939,N_1892,N_1851);
nor U1940 (N_1940,N_1897,N_1885);
nand U1941 (N_1941,N_1883,N_1895);
and U1942 (N_1942,N_1888,N_1859);
and U1943 (N_1943,N_1868,N_1883);
nand U1944 (N_1944,N_1868,N_1881);
or U1945 (N_1945,N_1894,N_1861);
and U1946 (N_1946,N_1884,N_1862);
nor U1947 (N_1947,N_1862,N_1859);
nor U1948 (N_1948,N_1869,N_1898);
nand U1949 (N_1949,N_1893,N_1864);
and U1950 (N_1950,N_1930,N_1925);
nand U1951 (N_1951,N_1913,N_1928);
or U1952 (N_1952,N_1910,N_1918);
and U1953 (N_1953,N_1922,N_1932);
nand U1954 (N_1954,N_1916,N_1940);
nand U1955 (N_1955,N_1946,N_1908);
and U1956 (N_1956,N_1909,N_1921);
nor U1957 (N_1957,N_1920,N_1907);
nand U1958 (N_1958,N_1919,N_1942);
and U1959 (N_1959,N_1929,N_1914);
or U1960 (N_1960,N_1933,N_1900);
nor U1961 (N_1961,N_1931,N_1915);
nor U1962 (N_1962,N_1905,N_1901);
or U1963 (N_1963,N_1923,N_1936);
nor U1964 (N_1964,N_1911,N_1906);
nor U1965 (N_1965,N_1902,N_1944);
nor U1966 (N_1966,N_1941,N_1917);
nand U1967 (N_1967,N_1935,N_1924);
or U1968 (N_1968,N_1945,N_1904);
nor U1969 (N_1969,N_1903,N_1937);
nor U1970 (N_1970,N_1927,N_1947);
or U1971 (N_1971,N_1926,N_1934);
and U1972 (N_1972,N_1912,N_1938);
or U1973 (N_1973,N_1948,N_1939);
nand U1974 (N_1974,N_1949,N_1943);
or U1975 (N_1975,N_1922,N_1931);
or U1976 (N_1976,N_1904,N_1938);
nand U1977 (N_1977,N_1929,N_1904);
or U1978 (N_1978,N_1914,N_1927);
or U1979 (N_1979,N_1917,N_1929);
or U1980 (N_1980,N_1945,N_1902);
or U1981 (N_1981,N_1914,N_1946);
nor U1982 (N_1982,N_1943,N_1901);
or U1983 (N_1983,N_1914,N_1939);
xor U1984 (N_1984,N_1948,N_1902);
or U1985 (N_1985,N_1915,N_1925);
nor U1986 (N_1986,N_1923,N_1919);
and U1987 (N_1987,N_1931,N_1944);
nor U1988 (N_1988,N_1908,N_1941);
and U1989 (N_1989,N_1905,N_1949);
nor U1990 (N_1990,N_1918,N_1949);
and U1991 (N_1991,N_1934,N_1932);
nor U1992 (N_1992,N_1911,N_1927);
nor U1993 (N_1993,N_1926,N_1909);
and U1994 (N_1994,N_1943,N_1929);
nand U1995 (N_1995,N_1919,N_1905);
nand U1996 (N_1996,N_1932,N_1943);
nand U1997 (N_1997,N_1943,N_1939);
nand U1998 (N_1998,N_1918,N_1937);
nor U1999 (N_1999,N_1914,N_1912);
or U2000 (N_2000,N_1996,N_1976);
nand U2001 (N_2001,N_1983,N_1991);
and U2002 (N_2002,N_1960,N_1978);
nand U2003 (N_2003,N_1987,N_1956);
xnor U2004 (N_2004,N_1950,N_1966);
and U2005 (N_2005,N_1999,N_1992);
nand U2006 (N_2006,N_1995,N_1997);
and U2007 (N_2007,N_1969,N_1988);
nand U2008 (N_2008,N_1975,N_1968);
and U2009 (N_2009,N_1954,N_1952);
nor U2010 (N_2010,N_1994,N_1989);
and U2011 (N_2011,N_1990,N_1951);
and U2012 (N_2012,N_1971,N_1986);
nand U2013 (N_2013,N_1973,N_1981);
nor U2014 (N_2014,N_1974,N_1980);
and U2015 (N_2015,N_1964,N_1984);
nand U2016 (N_2016,N_1970,N_1965);
nand U2017 (N_2017,N_1957,N_1958);
nor U2018 (N_2018,N_1962,N_1977);
or U2019 (N_2019,N_1959,N_1967);
nand U2020 (N_2020,N_1955,N_1998);
or U2021 (N_2021,N_1972,N_1985);
nand U2022 (N_2022,N_1961,N_1979);
nand U2023 (N_2023,N_1993,N_1953);
and U2024 (N_2024,N_1982,N_1963);
nor U2025 (N_2025,N_1983,N_1976);
and U2026 (N_2026,N_1990,N_1965);
nand U2027 (N_2027,N_1951,N_1993);
or U2028 (N_2028,N_1998,N_1973);
and U2029 (N_2029,N_1988,N_1950);
nand U2030 (N_2030,N_1956,N_1975);
and U2031 (N_2031,N_1967,N_1979);
and U2032 (N_2032,N_1959,N_1990);
and U2033 (N_2033,N_1975,N_1990);
nand U2034 (N_2034,N_1983,N_1978);
nor U2035 (N_2035,N_1961,N_1989);
nor U2036 (N_2036,N_1967,N_1968);
and U2037 (N_2037,N_1958,N_1977);
or U2038 (N_2038,N_1959,N_1962);
nand U2039 (N_2039,N_1963,N_1989);
and U2040 (N_2040,N_1986,N_1993);
or U2041 (N_2041,N_1976,N_1950);
or U2042 (N_2042,N_1989,N_1960);
and U2043 (N_2043,N_1953,N_1964);
nor U2044 (N_2044,N_1993,N_1974);
xor U2045 (N_2045,N_1977,N_1951);
nand U2046 (N_2046,N_1973,N_1964);
nand U2047 (N_2047,N_1960,N_1973);
nor U2048 (N_2048,N_1973,N_1963);
or U2049 (N_2049,N_1956,N_1969);
and U2050 (N_2050,N_2015,N_2007);
nand U2051 (N_2051,N_2019,N_2011);
nand U2052 (N_2052,N_2010,N_2043);
xor U2053 (N_2053,N_2022,N_2038);
nor U2054 (N_2054,N_2001,N_2023);
nor U2055 (N_2055,N_2032,N_2004);
or U2056 (N_2056,N_2045,N_2000);
and U2057 (N_2057,N_2005,N_2035);
nor U2058 (N_2058,N_2037,N_2033);
and U2059 (N_2059,N_2030,N_2002);
xnor U2060 (N_2060,N_2003,N_2042);
nand U2061 (N_2061,N_2034,N_2016);
nand U2062 (N_2062,N_2029,N_2012);
or U2063 (N_2063,N_2041,N_2039);
and U2064 (N_2064,N_2040,N_2025);
nand U2065 (N_2065,N_2008,N_2046);
nand U2066 (N_2066,N_2013,N_2014);
nor U2067 (N_2067,N_2028,N_2027);
nand U2068 (N_2068,N_2006,N_2031);
or U2069 (N_2069,N_2048,N_2024);
nor U2070 (N_2070,N_2049,N_2018);
and U2071 (N_2071,N_2021,N_2036);
or U2072 (N_2072,N_2017,N_2009);
nand U2073 (N_2073,N_2047,N_2026);
and U2074 (N_2074,N_2044,N_2020);
nor U2075 (N_2075,N_2008,N_2036);
nor U2076 (N_2076,N_2044,N_2048);
nor U2077 (N_2077,N_2021,N_2034);
nand U2078 (N_2078,N_2033,N_2042);
or U2079 (N_2079,N_2035,N_2041);
and U2080 (N_2080,N_2000,N_2008);
nor U2081 (N_2081,N_2027,N_2031);
or U2082 (N_2082,N_2005,N_2012);
and U2083 (N_2083,N_2008,N_2044);
nand U2084 (N_2084,N_2037,N_2018);
nand U2085 (N_2085,N_2035,N_2047);
or U2086 (N_2086,N_2006,N_2042);
or U2087 (N_2087,N_2027,N_2030);
nand U2088 (N_2088,N_2000,N_2010);
nand U2089 (N_2089,N_2025,N_2030);
nand U2090 (N_2090,N_2010,N_2005);
or U2091 (N_2091,N_2012,N_2039);
and U2092 (N_2092,N_2042,N_2038);
and U2093 (N_2093,N_2014,N_2007);
nor U2094 (N_2094,N_2016,N_2020);
nor U2095 (N_2095,N_2014,N_2032);
and U2096 (N_2096,N_2006,N_2011);
nand U2097 (N_2097,N_2034,N_2042);
and U2098 (N_2098,N_2000,N_2024);
or U2099 (N_2099,N_2010,N_2029);
nand U2100 (N_2100,N_2084,N_2078);
or U2101 (N_2101,N_2054,N_2091);
or U2102 (N_2102,N_2074,N_2070);
nor U2103 (N_2103,N_2092,N_2093);
nand U2104 (N_2104,N_2073,N_2077);
nor U2105 (N_2105,N_2088,N_2089);
nor U2106 (N_2106,N_2059,N_2081);
or U2107 (N_2107,N_2096,N_2061);
or U2108 (N_2108,N_2094,N_2083);
nand U2109 (N_2109,N_2071,N_2080);
nand U2110 (N_2110,N_2072,N_2085);
nand U2111 (N_2111,N_2064,N_2075);
nor U2112 (N_2112,N_2056,N_2050);
and U2113 (N_2113,N_2086,N_2063);
and U2114 (N_2114,N_2060,N_2057);
xor U2115 (N_2115,N_2067,N_2058);
or U2116 (N_2116,N_2068,N_2099);
nand U2117 (N_2117,N_2065,N_2090);
nand U2118 (N_2118,N_2079,N_2053);
or U2119 (N_2119,N_2062,N_2095);
nor U2120 (N_2120,N_2055,N_2069);
nor U2121 (N_2121,N_2097,N_2082);
nand U2122 (N_2122,N_2066,N_2051);
nand U2123 (N_2123,N_2087,N_2052);
nor U2124 (N_2124,N_2076,N_2098);
or U2125 (N_2125,N_2087,N_2065);
nor U2126 (N_2126,N_2059,N_2067);
or U2127 (N_2127,N_2074,N_2053);
nor U2128 (N_2128,N_2089,N_2078);
and U2129 (N_2129,N_2089,N_2062);
or U2130 (N_2130,N_2094,N_2067);
nor U2131 (N_2131,N_2052,N_2064);
nor U2132 (N_2132,N_2079,N_2087);
nor U2133 (N_2133,N_2079,N_2056);
and U2134 (N_2134,N_2094,N_2077);
nor U2135 (N_2135,N_2080,N_2097);
nand U2136 (N_2136,N_2051,N_2085);
or U2137 (N_2137,N_2062,N_2087);
nor U2138 (N_2138,N_2097,N_2055);
nor U2139 (N_2139,N_2060,N_2089);
and U2140 (N_2140,N_2079,N_2078);
and U2141 (N_2141,N_2072,N_2082);
nand U2142 (N_2142,N_2056,N_2076);
and U2143 (N_2143,N_2051,N_2054);
and U2144 (N_2144,N_2060,N_2061);
nor U2145 (N_2145,N_2071,N_2085);
nand U2146 (N_2146,N_2068,N_2075);
and U2147 (N_2147,N_2082,N_2090);
or U2148 (N_2148,N_2095,N_2072);
nand U2149 (N_2149,N_2051,N_2075);
nor U2150 (N_2150,N_2114,N_2116);
nor U2151 (N_2151,N_2108,N_2133);
and U2152 (N_2152,N_2142,N_2141);
nor U2153 (N_2153,N_2126,N_2136);
and U2154 (N_2154,N_2132,N_2130);
nand U2155 (N_2155,N_2118,N_2106);
and U2156 (N_2156,N_2138,N_2134);
nand U2157 (N_2157,N_2135,N_2103);
nor U2158 (N_2158,N_2120,N_2122);
nand U2159 (N_2159,N_2124,N_2112);
nand U2160 (N_2160,N_2147,N_2101);
or U2161 (N_2161,N_2105,N_2119);
nor U2162 (N_2162,N_2115,N_2111);
nand U2163 (N_2163,N_2128,N_2148);
and U2164 (N_2164,N_2146,N_2107);
nand U2165 (N_2165,N_2123,N_2145);
or U2166 (N_2166,N_2127,N_2131);
nor U2167 (N_2167,N_2117,N_2129);
and U2168 (N_2168,N_2125,N_2100);
or U2169 (N_2169,N_2137,N_2140);
and U2170 (N_2170,N_2139,N_2113);
or U2171 (N_2171,N_2121,N_2104);
and U2172 (N_2172,N_2144,N_2143);
nor U2173 (N_2173,N_2149,N_2102);
nor U2174 (N_2174,N_2110,N_2109);
and U2175 (N_2175,N_2145,N_2119);
or U2176 (N_2176,N_2111,N_2145);
nor U2177 (N_2177,N_2131,N_2145);
nand U2178 (N_2178,N_2102,N_2116);
or U2179 (N_2179,N_2131,N_2121);
or U2180 (N_2180,N_2149,N_2103);
or U2181 (N_2181,N_2113,N_2136);
nor U2182 (N_2182,N_2145,N_2142);
or U2183 (N_2183,N_2107,N_2130);
or U2184 (N_2184,N_2129,N_2105);
and U2185 (N_2185,N_2108,N_2103);
nor U2186 (N_2186,N_2126,N_2147);
nor U2187 (N_2187,N_2127,N_2145);
or U2188 (N_2188,N_2112,N_2146);
nand U2189 (N_2189,N_2147,N_2136);
nor U2190 (N_2190,N_2113,N_2106);
and U2191 (N_2191,N_2119,N_2110);
or U2192 (N_2192,N_2132,N_2105);
or U2193 (N_2193,N_2143,N_2111);
and U2194 (N_2194,N_2129,N_2145);
and U2195 (N_2195,N_2107,N_2142);
and U2196 (N_2196,N_2133,N_2143);
and U2197 (N_2197,N_2107,N_2131);
and U2198 (N_2198,N_2108,N_2136);
nor U2199 (N_2199,N_2127,N_2114);
or U2200 (N_2200,N_2157,N_2184);
nand U2201 (N_2201,N_2178,N_2163);
nor U2202 (N_2202,N_2187,N_2169);
or U2203 (N_2203,N_2155,N_2185);
or U2204 (N_2204,N_2195,N_2188);
and U2205 (N_2205,N_2153,N_2173);
or U2206 (N_2206,N_2164,N_2152);
or U2207 (N_2207,N_2151,N_2183);
nand U2208 (N_2208,N_2177,N_2193);
and U2209 (N_2209,N_2171,N_2191);
nand U2210 (N_2210,N_2172,N_2167);
nor U2211 (N_2211,N_2186,N_2168);
or U2212 (N_2212,N_2189,N_2179);
or U2213 (N_2213,N_2181,N_2199);
or U2214 (N_2214,N_2175,N_2158);
and U2215 (N_2215,N_2192,N_2160);
nor U2216 (N_2216,N_2165,N_2198);
and U2217 (N_2217,N_2196,N_2190);
or U2218 (N_2218,N_2180,N_2154);
and U2219 (N_2219,N_2159,N_2174);
nor U2220 (N_2220,N_2197,N_2166);
nor U2221 (N_2221,N_2161,N_2194);
nand U2222 (N_2222,N_2176,N_2156);
nand U2223 (N_2223,N_2162,N_2170);
or U2224 (N_2224,N_2150,N_2182);
or U2225 (N_2225,N_2156,N_2157);
and U2226 (N_2226,N_2182,N_2152);
nand U2227 (N_2227,N_2179,N_2194);
nand U2228 (N_2228,N_2191,N_2161);
nor U2229 (N_2229,N_2160,N_2196);
nor U2230 (N_2230,N_2155,N_2154);
or U2231 (N_2231,N_2185,N_2159);
nor U2232 (N_2232,N_2181,N_2182);
and U2233 (N_2233,N_2183,N_2181);
and U2234 (N_2234,N_2192,N_2198);
and U2235 (N_2235,N_2164,N_2189);
nor U2236 (N_2236,N_2160,N_2194);
nor U2237 (N_2237,N_2151,N_2154);
or U2238 (N_2238,N_2189,N_2180);
and U2239 (N_2239,N_2181,N_2160);
nand U2240 (N_2240,N_2182,N_2169);
and U2241 (N_2241,N_2184,N_2179);
nor U2242 (N_2242,N_2179,N_2185);
nand U2243 (N_2243,N_2187,N_2184);
nor U2244 (N_2244,N_2156,N_2182);
nor U2245 (N_2245,N_2172,N_2189);
and U2246 (N_2246,N_2158,N_2160);
xnor U2247 (N_2247,N_2179,N_2167);
nand U2248 (N_2248,N_2166,N_2183);
and U2249 (N_2249,N_2180,N_2166);
and U2250 (N_2250,N_2227,N_2217);
and U2251 (N_2251,N_2218,N_2220);
and U2252 (N_2252,N_2237,N_2249);
nand U2253 (N_2253,N_2219,N_2246);
and U2254 (N_2254,N_2207,N_2205);
nand U2255 (N_2255,N_2206,N_2239);
nor U2256 (N_2256,N_2221,N_2215);
nand U2257 (N_2257,N_2232,N_2209);
and U2258 (N_2258,N_2226,N_2212);
nand U2259 (N_2259,N_2236,N_2244);
and U2260 (N_2260,N_2230,N_2201);
nor U2261 (N_2261,N_2247,N_2235);
and U2262 (N_2262,N_2225,N_2211);
and U2263 (N_2263,N_2234,N_2202);
or U2264 (N_2264,N_2233,N_2214);
or U2265 (N_2265,N_2222,N_2228);
nor U2266 (N_2266,N_2241,N_2213);
or U2267 (N_2267,N_2242,N_2224);
and U2268 (N_2268,N_2231,N_2208);
or U2269 (N_2269,N_2245,N_2248);
and U2270 (N_2270,N_2223,N_2216);
nor U2271 (N_2271,N_2240,N_2210);
nor U2272 (N_2272,N_2203,N_2204);
nor U2273 (N_2273,N_2229,N_2243);
nor U2274 (N_2274,N_2200,N_2238);
nor U2275 (N_2275,N_2241,N_2212);
and U2276 (N_2276,N_2235,N_2221);
nand U2277 (N_2277,N_2238,N_2233);
and U2278 (N_2278,N_2201,N_2227);
nand U2279 (N_2279,N_2220,N_2247);
nand U2280 (N_2280,N_2213,N_2206);
nand U2281 (N_2281,N_2212,N_2215);
nor U2282 (N_2282,N_2225,N_2206);
or U2283 (N_2283,N_2206,N_2214);
or U2284 (N_2284,N_2218,N_2244);
xor U2285 (N_2285,N_2245,N_2226);
and U2286 (N_2286,N_2245,N_2202);
or U2287 (N_2287,N_2231,N_2213);
and U2288 (N_2288,N_2234,N_2228);
or U2289 (N_2289,N_2214,N_2200);
or U2290 (N_2290,N_2241,N_2204);
and U2291 (N_2291,N_2225,N_2205);
nor U2292 (N_2292,N_2209,N_2227);
and U2293 (N_2293,N_2202,N_2239);
or U2294 (N_2294,N_2239,N_2237);
or U2295 (N_2295,N_2233,N_2226);
nand U2296 (N_2296,N_2242,N_2247);
nor U2297 (N_2297,N_2246,N_2247);
and U2298 (N_2298,N_2227,N_2216);
nand U2299 (N_2299,N_2200,N_2213);
nand U2300 (N_2300,N_2279,N_2276);
nand U2301 (N_2301,N_2291,N_2281);
nand U2302 (N_2302,N_2295,N_2288);
nor U2303 (N_2303,N_2273,N_2250);
or U2304 (N_2304,N_2289,N_2297);
and U2305 (N_2305,N_2278,N_2256);
nor U2306 (N_2306,N_2284,N_2254);
and U2307 (N_2307,N_2265,N_2270);
nand U2308 (N_2308,N_2277,N_2285);
nor U2309 (N_2309,N_2268,N_2298);
and U2310 (N_2310,N_2251,N_2290);
or U2311 (N_2311,N_2253,N_2272);
and U2312 (N_2312,N_2252,N_2258);
or U2313 (N_2313,N_2283,N_2263);
nand U2314 (N_2314,N_2282,N_2274);
and U2315 (N_2315,N_2255,N_2262);
nor U2316 (N_2316,N_2286,N_2264);
or U2317 (N_2317,N_2267,N_2287);
and U2318 (N_2318,N_2294,N_2259);
nand U2319 (N_2319,N_2261,N_2260);
or U2320 (N_2320,N_2271,N_2299);
and U2321 (N_2321,N_2275,N_2269);
and U2322 (N_2322,N_2280,N_2293);
nor U2323 (N_2323,N_2266,N_2296);
nor U2324 (N_2324,N_2292,N_2257);
and U2325 (N_2325,N_2290,N_2269);
and U2326 (N_2326,N_2293,N_2254);
and U2327 (N_2327,N_2272,N_2267);
or U2328 (N_2328,N_2273,N_2266);
nor U2329 (N_2329,N_2251,N_2285);
nand U2330 (N_2330,N_2259,N_2257);
or U2331 (N_2331,N_2272,N_2252);
or U2332 (N_2332,N_2296,N_2288);
and U2333 (N_2333,N_2256,N_2263);
nor U2334 (N_2334,N_2291,N_2257);
nor U2335 (N_2335,N_2287,N_2259);
nor U2336 (N_2336,N_2263,N_2260);
nand U2337 (N_2337,N_2262,N_2278);
and U2338 (N_2338,N_2296,N_2274);
nand U2339 (N_2339,N_2295,N_2273);
nor U2340 (N_2340,N_2290,N_2266);
or U2341 (N_2341,N_2272,N_2290);
and U2342 (N_2342,N_2298,N_2254);
and U2343 (N_2343,N_2252,N_2271);
nand U2344 (N_2344,N_2264,N_2268);
and U2345 (N_2345,N_2278,N_2285);
and U2346 (N_2346,N_2254,N_2271);
and U2347 (N_2347,N_2266,N_2250);
nand U2348 (N_2348,N_2257,N_2298);
nor U2349 (N_2349,N_2289,N_2250);
nand U2350 (N_2350,N_2302,N_2313);
nor U2351 (N_2351,N_2336,N_2330);
nand U2352 (N_2352,N_2307,N_2340);
nor U2353 (N_2353,N_2308,N_2335);
nand U2354 (N_2354,N_2347,N_2329);
and U2355 (N_2355,N_2322,N_2333);
nand U2356 (N_2356,N_2314,N_2331);
or U2357 (N_2357,N_2339,N_2312);
and U2358 (N_2358,N_2319,N_2326);
or U2359 (N_2359,N_2309,N_2343);
and U2360 (N_2360,N_2327,N_2344);
nand U2361 (N_2361,N_2315,N_2348);
and U2362 (N_2362,N_2301,N_2341);
or U2363 (N_2363,N_2337,N_2320);
nand U2364 (N_2364,N_2345,N_2321);
and U2365 (N_2365,N_2349,N_2328);
nor U2366 (N_2366,N_2317,N_2305);
or U2367 (N_2367,N_2323,N_2325);
or U2368 (N_2368,N_2334,N_2324);
nor U2369 (N_2369,N_2304,N_2316);
and U2370 (N_2370,N_2306,N_2346);
and U2371 (N_2371,N_2300,N_2338);
and U2372 (N_2372,N_2310,N_2342);
nor U2373 (N_2373,N_2332,N_2311);
nand U2374 (N_2374,N_2303,N_2318);
or U2375 (N_2375,N_2306,N_2315);
nand U2376 (N_2376,N_2308,N_2344);
nor U2377 (N_2377,N_2311,N_2345);
nand U2378 (N_2378,N_2337,N_2340);
nor U2379 (N_2379,N_2301,N_2317);
and U2380 (N_2380,N_2323,N_2309);
nand U2381 (N_2381,N_2318,N_2312);
and U2382 (N_2382,N_2326,N_2348);
nor U2383 (N_2383,N_2346,N_2332);
and U2384 (N_2384,N_2336,N_2335);
or U2385 (N_2385,N_2344,N_2346);
or U2386 (N_2386,N_2346,N_2330);
nor U2387 (N_2387,N_2347,N_2311);
nand U2388 (N_2388,N_2347,N_2338);
nor U2389 (N_2389,N_2319,N_2327);
nand U2390 (N_2390,N_2332,N_2308);
and U2391 (N_2391,N_2306,N_2304);
nand U2392 (N_2392,N_2320,N_2321);
and U2393 (N_2393,N_2335,N_2322);
nor U2394 (N_2394,N_2324,N_2344);
or U2395 (N_2395,N_2310,N_2306);
or U2396 (N_2396,N_2326,N_2302);
nor U2397 (N_2397,N_2322,N_2345);
or U2398 (N_2398,N_2308,N_2320);
nor U2399 (N_2399,N_2317,N_2349);
or U2400 (N_2400,N_2371,N_2364);
nand U2401 (N_2401,N_2393,N_2365);
nand U2402 (N_2402,N_2377,N_2399);
nand U2403 (N_2403,N_2355,N_2387);
or U2404 (N_2404,N_2353,N_2388);
nor U2405 (N_2405,N_2369,N_2375);
nand U2406 (N_2406,N_2374,N_2356);
and U2407 (N_2407,N_2395,N_2358);
nor U2408 (N_2408,N_2384,N_2390);
and U2409 (N_2409,N_2385,N_2396);
nor U2410 (N_2410,N_2354,N_2379);
or U2411 (N_2411,N_2372,N_2359);
nor U2412 (N_2412,N_2391,N_2383);
and U2413 (N_2413,N_2373,N_2368);
nand U2414 (N_2414,N_2378,N_2361);
and U2415 (N_2415,N_2386,N_2363);
and U2416 (N_2416,N_2382,N_2397);
nor U2417 (N_2417,N_2357,N_2367);
nand U2418 (N_2418,N_2362,N_2380);
nand U2419 (N_2419,N_2351,N_2392);
or U2420 (N_2420,N_2366,N_2352);
nor U2421 (N_2421,N_2381,N_2350);
nor U2422 (N_2422,N_2370,N_2398);
and U2423 (N_2423,N_2360,N_2389);
nand U2424 (N_2424,N_2394,N_2376);
nand U2425 (N_2425,N_2391,N_2390);
nand U2426 (N_2426,N_2379,N_2370);
and U2427 (N_2427,N_2380,N_2351);
nor U2428 (N_2428,N_2377,N_2370);
or U2429 (N_2429,N_2386,N_2397);
nand U2430 (N_2430,N_2356,N_2386);
nand U2431 (N_2431,N_2372,N_2351);
or U2432 (N_2432,N_2394,N_2368);
or U2433 (N_2433,N_2389,N_2382);
and U2434 (N_2434,N_2383,N_2363);
or U2435 (N_2435,N_2357,N_2364);
nand U2436 (N_2436,N_2374,N_2368);
and U2437 (N_2437,N_2350,N_2389);
and U2438 (N_2438,N_2367,N_2352);
nand U2439 (N_2439,N_2360,N_2386);
and U2440 (N_2440,N_2394,N_2387);
and U2441 (N_2441,N_2356,N_2377);
nor U2442 (N_2442,N_2375,N_2395);
or U2443 (N_2443,N_2378,N_2389);
and U2444 (N_2444,N_2371,N_2377);
or U2445 (N_2445,N_2390,N_2357);
nor U2446 (N_2446,N_2368,N_2358);
or U2447 (N_2447,N_2362,N_2386);
nor U2448 (N_2448,N_2382,N_2398);
nand U2449 (N_2449,N_2396,N_2380);
nand U2450 (N_2450,N_2418,N_2425);
nor U2451 (N_2451,N_2429,N_2428);
nor U2452 (N_2452,N_2431,N_2404);
or U2453 (N_2453,N_2419,N_2443);
and U2454 (N_2454,N_2438,N_2407);
nor U2455 (N_2455,N_2445,N_2414);
nor U2456 (N_2456,N_2415,N_2437);
nand U2457 (N_2457,N_2422,N_2402);
and U2458 (N_2458,N_2433,N_2435);
nand U2459 (N_2459,N_2406,N_2446);
or U2460 (N_2460,N_2448,N_2436);
nor U2461 (N_2461,N_2440,N_2447);
nor U2462 (N_2462,N_2432,N_2401);
and U2463 (N_2463,N_2424,N_2442);
nand U2464 (N_2464,N_2417,N_2427);
nand U2465 (N_2465,N_2421,N_2403);
nand U2466 (N_2466,N_2416,N_2434);
or U2467 (N_2467,N_2449,N_2409);
and U2468 (N_2468,N_2420,N_2426);
or U2469 (N_2469,N_2410,N_2439);
and U2470 (N_2470,N_2423,N_2430);
and U2471 (N_2471,N_2408,N_2411);
or U2472 (N_2472,N_2444,N_2441);
nand U2473 (N_2473,N_2412,N_2400);
and U2474 (N_2474,N_2405,N_2413);
and U2475 (N_2475,N_2435,N_2400);
and U2476 (N_2476,N_2445,N_2431);
or U2477 (N_2477,N_2411,N_2418);
nand U2478 (N_2478,N_2420,N_2413);
and U2479 (N_2479,N_2409,N_2408);
or U2480 (N_2480,N_2435,N_2412);
nor U2481 (N_2481,N_2400,N_2448);
nor U2482 (N_2482,N_2411,N_2430);
and U2483 (N_2483,N_2410,N_2426);
or U2484 (N_2484,N_2415,N_2410);
and U2485 (N_2485,N_2433,N_2443);
or U2486 (N_2486,N_2417,N_2448);
or U2487 (N_2487,N_2404,N_2445);
nor U2488 (N_2488,N_2424,N_2420);
nor U2489 (N_2489,N_2413,N_2429);
nand U2490 (N_2490,N_2433,N_2407);
nand U2491 (N_2491,N_2411,N_2415);
or U2492 (N_2492,N_2446,N_2408);
and U2493 (N_2493,N_2421,N_2423);
nand U2494 (N_2494,N_2432,N_2427);
and U2495 (N_2495,N_2422,N_2401);
xor U2496 (N_2496,N_2405,N_2424);
and U2497 (N_2497,N_2408,N_2412);
nor U2498 (N_2498,N_2421,N_2430);
and U2499 (N_2499,N_2421,N_2411);
nand U2500 (N_2500,N_2475,N_2496);
nand U2501 (N_2501,N_2495,N_2493);
nor U2502 (N_2502,N_2467,N_2484);
nand U2503 (N_2503,N_2469,N_2480);
nand U2504 (N_2504,N_2492,N_2471);
and U2505 (N_2505,N_2486,N_2450);
or U2506 (N_2506,N_2464,N_2490);
nand U2507 (N_2507,N_2466,N_2487);
or U2508 (N_2508,N_2463,N_2455);
nor U2509 (N_2509,N_2494,N_2452);
or U2510 (N_2510,N_2457,N_2454);
or U2511 (N_2511,N_2474,N_2499);
and U2512 (N_2512,N_2456,N_2489);
or U2513 (N_2513,N_2485,N_2481);
nand U2514 (N_2514,N_2451,N_2482);
nor U2515 (N_2515,N_2472,N_2470);
or U2516 (N_2516,N_2498,N_2461);
or U2517 (N_2517,N_2476,N_2478);
or U2518 (N_2518,N_2453,N_2483);
or U2519 (N_2519,N_2458,N_2497);
and U2520 (N_2520,N_2479,N_2460);
nor U2521 (N_2521,N_2462,N_2465);
nand U2522 (N_2522,N_2477,N_2491);
nor U2523 (N_2523,N_2473,N_2459);
nor U2524 (N_2524,N_2468,N_2488);
and U2525 (N_2525,N_2488,N_2480);
nand U2526 (N_2526,N_2480,N_2459);
nand U2527 (N_2527,N_2470,N_2460);
nand U2528 (N_2528,N_2459,N_2482);
nor U2529 (N_2529,N_2461,N_2456);
nor U2530 (N_2530,N_2462,N_2466);
and U2531 (N_2531,N_2460,N_2458);
nand U2532 (N_2532,N_2484,N_2462);
nand U2533 (N_2533,N_2465,N_2456);
and U2534 (N_2534,N_2467,N_2490);
or U2535 (N_2535,N_2450,N_2490);
nand U2536 (N_2536,N_2475,N_2474);
nor U2537 (N_2537,N_2474,N_2488);
and U2538 (N_2538,N_2480,N_2454);
and U2539 (N_2539,N_2479,N_2493);
nand U2540 (N_2540,N_2458,N_2456);
or U2541 (N_2541,N_2458,N_2465);
and U2542 (N_2542,N_2495,N_2475);
and U2543 (N_2543,N_2491,N_2458);
and U2544 (N_2544,N_2466,N_2461);
and U2545 (N_2545,N_2461,N_2460);
nand U2546 (N_2546,N_2480,N_2455);
and U2547 (N_2547,N_2477,N_2495);
and U2548 (N_2548,N_2462,N_2481);
nor U2549 (N_2549,N_2476,N_2453);
and U2550 (N_2550,N_2525,N_2547);
xor U2551 (N_2551,N_2521,N_2503);
or U2552 (N_2552,N_2544,N_2537);
nor U2553 (N_2553,N_2505,N_2526);
or U2554 (N_2554,N_2531,N_2539);
nand U2555 (N_2555,N_2512,N_2523);
or U2556 (N_2556,N_2532,N_2507);
nor U2557 (N_2557,N_2549,N_2501);
and U2558 (N_2558,N_2504,N_2510);
xor U2559 (N_2559,N_2528,N_2516);
nor U2560 (N_2560,N_2522,N_2533);
nand U2561 (N_2561,N_2514,N_2519);
and U2562 (N_2562,N_2524,N_2536);
nor U2563 (N_2563,N_2500,N_2527);
nor U2564 (N_2564,N_2546,N_2511);
nor U2565 (N_2565,N_2517,N_2548);
nand U2566 (N_2566,N_2506,N_2509);
nand U2567 (N_2567,N_2530,N_2520);
and U2568 (N_2568,N_2538,N_2543);
nand U2569 (N_2569,N_2502,N_2541);
nand U2570 (N_2570,N_2518,N_2535);
nor U2571 (N_2571,N_2542,N_2513);
nor U2572 (N_2572,N_2540,N_2545);
and U2573 (N_2573,N_2515,N_2508);
or U2574 (N_2574,N_2529,N_2534);
or U2575 (N_2575,N_2521,N_2541);
or U2576 (N_2576,N_2536,N_2519);
nand U2577 (N_2577,N_2521,N_2515);
nand U2578 (N_2578,N_2522,N_2506);
and U2579 (N_2579,N_2525,N_2516);
nand U2580 (N_2580,N_2510,N_2530);
nand U2581 (N_2581,N_2549,N_2543);
or U2582 (N_2582,N_2521,N_2523);
and U2583 (N_2583,N_2521,N_2500);
or U2584 (N_2584,N_2542,N_2504);
or U2585 (N_2585,N_2529,N_2513);
or U2586 (N_2586,N_2506,N_2516);
and U2587 (N_2587,N_2501,N_2548);
nor U2588 (N_2588,N_2524,N_2549);
and U2589 (N_2589,N_2530,N_2504);
nor U2590 (N_2590,N_2517,N_2507);
and U2591 (N_2591,N_2505,N_2530);
or U2592 (N_2592,N_2549,N_2532);
nor U2593 (N_2593,N_2505,N_2536);
nor U2594 (N_2594,N_2534,N_2517);
and U2595 (N_2595,N_2536,N_2506);
nor U2596 (N_2596,N_2517,N_2518);
or U2597 (N_2597,N_2528,N_2524);
xor U2598 (N_2598,N_2521,N_2536);
nand U2599 (N_2599,N_2504,N_2522);
nand U2600 (N_2600,N_2561,N_2570);
or U2601 (N_2601,N_2556,N_2569);
nand U2602 (N_2602,N_2571,N_2580);
nor U2603 (N_2603,N_2560,N_2585);
and U2604 (N_2604,N_2550,N_2558);
or U2605 (N_2605,N_2573,N_2552);
nand U2606 (N_2606,N_2572,N_2592);
and U2607 (N_2607,N_2586,N_2597);
and U2608 (N_2608,N_2576,N_2581);
and U2609 (N_2609,N_2564,N_2577);
or U2610 (N_2610,N_2554,N_2578);
or U2611 (N_2611,N_2575,N_2563);
nand U2612 (N_2612,N_2596,N_2583);
nand U2613 (N_2613,N_2594,N_2599);
nor U2614 (N_2614,N_2567,N_2579);
nor U2615 (N_2615,N_2587,N_2559);
nand U2616 (N_2616,N_2591,N_2595);
nand U2617 (N_2617,N_2562,N_2582);
and U2618 (N_2618,N_2589,N_2588);
nand U2619 (N_2619,N_2557,N_2584);
and U2620 (N_2620,N_2551,N_2555);
and U2621 (N_2621,N_2590,N_2565);
nor U2622 (N_2622,N_2598,N_2574);
or U2623 (N_2623,N_2553,N_2568);
or U2624 (N_2624,N_2593,N_2566);
and U2625 (N_2625,N_2595,N_2580);
and U2626 (N_2626,N_2581,N_2572);
and U2627 (N_2627,N_2578,N_2558);
and U2628 (N_2628,N_2594,N_2570);
and U2629 (N_2629,N_2574,N_2599);
and U2630 (N_2630,N_2583,N_2555);
and U2631 (N_2631,N_2586,N_2590);
and U2632 (N_2632,N_2597,N_2577);
or U2633 (N_2633,N_2553,N_2587);
nand U2634 (N_2634,N_2555,N_2594);
nand U2635 (N_2635,N_2566,N_2556);
or U2636 (N_2636,N_2576,N_2586);
nor U2637 (N_2637,N_2586,N_2550);
or U2638 (N_2638,N_2581,N_2566);
nand U2639 (N_2639,N_2557,N_2588);
or U2640 (N_2640,N_2560,N_2570);
nor U2641 (N_2641,N_2553,N_2562);
nor U2642 (N_2642,N_2554,N_2589);
or U2643 (N_2643,N_2557,N_2553);
nand U2644 (N_2644,N_2581,N_2553);
and U2645 (N_2645,N_2572,N_2566);
nand U2646 (N_2646,N_2570,N_2596);
or U2647 (N_2647,N_2554,N_2579);
and U2648 (N_2648,N_2573,N_2597);
or U2649 (N_2649,N_2571,N_2560);
and U2650 (N_2650,N_2634,N_2611);
nand U2651 (N_2651,N_2614,N_2635);
and U2652 (N_2652,N_2616,N_2608);
or U2653 (N_2653,N_2640,N_2624);
nand U2654 (N_2654,N_2623,N_2646);
nand U2655 (N_2655,N_2630,N_2643);
and U2656 (N_2656,N_2647,N_2648);
or U2657 (N_2657,N_2613,N_2602);
or U2658 (N_2658,N_2600,N_2607);
and U2659 (N_2659,N_2637,N_2632);
or U2660 (N_2660,N_2609,N_2605);
or U2661 (N_2661,N_2601,N_2628);
and U2662 (N_2662,N_2644,N_2612);
nand U2663 (N_2663,N_2645,N_2631);
nand U2664 (N_2664,N_2638,N_2603);
or U2665 (N_2665,N_2639,N_2618);
or U2666 (N_2666,N_2626,N_2649);
nand U2667 (N_2667,N_2622,N_2627);
or U2668 (N_2668,N_2606,N_2625);
and U2669 (N_2669,N_2642,N_2615);
nand U2670 (N_2670,N_2617,N_2621);
or U2671 (N_2671,N_2629,N_2604);
and U2672 (N_2672,N_2620,N_2633);
and U2673 (N_2673,N_2641,N_2636);
and U2674 (N_2674,N_2610,N_2619);
nor U2675 (N_2675,N_2617,N_2608);
nor U2676 (N_2676,N_2623,N_2632);
and U2677 (N_2677,N_2636,N_2630);
nor U2678 (N_2678,N_2604,N_2619);
or U2679 (N_2679,N_2642,N_2631);
or U2680 (N_2680,N_2646,N_2624);
and U2681 (N_2681,N_2640,N_2620);
nor U2682 (N_2682,N_2646,N_2622);
nand U2683 (N_2683,N_2609,N_2631);
and U2684 (N_2684,N_2646,N_2642);
and U2685 (N_2685,N_2633,N_2618);
nand U2686 (N_2686,N_2630,N_2642);
and U2687 (N_2687,N_2649,N_2642);
or U2688 (N_2688,N_2609,N_2617);
and U2689 (N_2689,N_2648,N_2613);
or U2690 (N_2690,N_2617,N_2618);
nor U2691 (N_2691,N_2635,N_2622);
nor U2692 (N_2692,N_2649,N_2635);
nand U2693 (N_2693,N_2603,N_2643);
and U2694 (N_2694,N_2647,N_2634);
or U2695 (N_2695,N_2624,N_2608);
nor U2696 (N_2696,N_2627,N_2616);
or U2697 (N_2697,N_2633,N_2622);
nor U2698 (N_2698,N_2604,N_2630);
or U2699 (N_2699,N_2644,N_2616);
or U2700 (N_2700,N_2683,N_2654);
nor U2701 (N_2701,N_2688,N_2698);
or U2702 (N_2702,N_2689,N_2663);
nand U2703 (N_2703,N_2686,N_2657);
and U2704 (N_2704,N_2687,N_2694);
nand U2705 (N_2705,N_2660,N_2651);
nand U2706 (N_2706,N_2659,N_2656);
and U2707 (N_2707,N_2685,N_2668);
nand U2708 (N_2708,N_2682,N_2692);
or U2709 (N_2709,N_2696,N_2672);
or U2710 (N_2710,N_2665,N_2684);
and U2711 (N_2711,N_2669,N_2690);
nor U2712 (N_2712,N_2695,N_2679);
and U2713 (N_2713,N_2650,N_2681);
nor U2714 (N_2714,N_2658,N_2670);
or U2715 (N_2715,N_2678,N_2676);
nor U2716 (N_2716,N_2693,N_2666);
nor U2717 (N_2717,N_2661,N_2662);
nand U2718 (N_2718,N_2652,N_2673);
or U2719 (N_2719,N_2664,N_2671);
or U2720 (N_2720,N_2674,N_2675);
or U2721 (N_2721,N_2691,N_2653);
or U2722 (N_2722,N_2697,N_2699);
nand U2723 (N_2723,N_2677,N_2655);
or U2724 (N_2724,N_2667,N_2680);
nand U2725 (N_2725,N_2681,N_2684);
and U2726 (N_2726,N_2684,N_2659);
nor U2727 (N_2727,N_2664,N_2651);
nand U2728 (N_2728,N_2651,N_2670);
or U2729 (N_2729,N_2673,N_2697);
or U2730 (N_2730,N_2686,N_2666);
or U2731 (N_2731,N_2690,N_2686);
nor U2732 (N_2732,N_2689,N_2664);
and U2733 (N_2733,N_2678,N_2663);
or U2734 (N_2734,N_2698,N_2695);
nand U2735 (N_2735,N_2673,N_2684);
xnor U2736 (N_2736,N_2681,N_2672);
or U2737 (N_2737,N_2658,N_2673);
or U2738 (N_2738,N_2696,N_2651);
or U2739 (N_2739,N_2665,N_2688);
nand U2740 (N_2740,N_2669,N_2657);
or U2741 (N_2741,N_2677,N_2673);
and U2742 (N_2742,N_2654,N_2681);
nor U2743 (N_2743,N_2675,N_2650);
nand U2744 (N_2744,N_2692,N_2678);
xnor U2745 (N_2745,N_2668,N_2653);
nor U2746 (N_2746,N_2699,N_2668);
nor U2747 (N_2747,N_2668,N_2659);
or U2748 (N_2748,N_2699,N_2692);
or U2749 (N_2749,N_2689,N_2661);
nand U2750 (N_2750,N_2733,N_2725);
or U2751 (N_2751,N_2703,N_2726);
or U2752 (N_2752,N_2714,N_2746);
nor U2753 (N_2753,N_2706,N_2721);
nor U2754 (N_2754,N_2722,N_2720);
nor U2755 (N_2755,N_2710,N_2736);
nor U2756 (N_2756,N_2729,N_2712);
nor U2757 (N_2757,N_2705,N_2700);
or U2758 (N_2758,N_2739,N_2724);
or U2759 (N_2759,N_2732,N_2701);
and U2760 (N_2760,N_2749,N_2731);
or U2761 (N_2761,N_2713,N_2704);
and U2762 (N_2762,N_2723,N_2718);
nand U2763 (N_2763,N_2707,N_2730);
nor U2764 (N_2764,N_2748,N_2737);
xor U2765 (N_2765,N_2738,N_2741);
and U2766 (N_2766,N_2709,N_2735);
and U2767 (N_2767,N_2747,N_2702);
and U2768 (N_2768,N_2715,N_2743);
and U2769 (N_2769,N_2740,N_2716);
nand U2770 (N_2770,N_2708,N_2734);
nand U2771 (N_2771,N_2728,N_2745);
nor U2772 (N_2772,N_2711,N_2719);
nor U2773 (N_2773,N_2744,N_2727);
and U2774 (N_2774,N_2742,N_2717);
and U2775 (N_2775,N_2734,N_2737);
or U2776 (N_2776,N_2705,N_2710);
or U2777 (N_2777,N_2733,N_2724);
nand U2778 (N_2778,N_2711,N_2740);
nor U2779 (N_2779,N_2703,N_2705);
xor U2780 (N_2780,N_2739,N_2748);
or U2781 (N_2781,N_2706,N_2737);
nand U2782 (N_2782,N_2719,N_2734);
and U2783 (N_2783,N_2700,N_2718);
or U2784 (N_2784,N_2748,N_2731);
and U2785 (N_2785,N_2736,N_2725);
nand U2786 (N_2786,N_2702,N_2719);
or U2787 (N_2787,N_2724,N_2701);
nand U2788 (N_2788,N_2748,N_2717);
nand U2789 (N_2789,N_2719,N_2706);
nand U2790 (N_2790,N_2736,N_2724);
and U2791 (N_2791,N_2746,N_2712);
xnor U2792 (N_2792,N_2727,N_2732);
nor U2793 (N_2793,N_2717,N_2718);
or U2794 (N_2794,N_2713,N_2737);
and U2795 (N_2795,N_2735,N_2716);
or U2796 (N_2796,N_2707,N_2727);
xnor U2797 (N_2797,N_2734,N_2740);
nor U2798 (N_2798,N_2703,N_2749);
nor U2799 (N_2799,N_2728,N_2740);
or U2800 (N_2800,N_2772,N_2798);
and U2801 (N_2801,N_2762,N_2751);
nor U2802 (N_2802,N_2797,N_2782);
or U2803 (N_2803,N_2754,N_2799);
or U2804 (N_2804,N_2756,N_2792);
nand U2805 (N_2805,N_2790,N_2753);
nor U2806 (N_2806,N_2773,N_2768);
nor U2807 (N_2807,N_2765,N_2781);
nand U2808 (N_2808,N_2796,N_2789);
or U2809 (N_2809,N_2775,N_2793);
or U2810 (N_2810,N_2776,N_2752);
and U2811 (N_2811,N_2778,N_2786);
or U2812 (N_2812,N_2770,N_2755);
nand U2813 (N_2813,N_2785,N_2759);
nand U2814 (N_2814,N_2780,N_2760);
nand U2815 (N_2815,N_2767,N_2757);
nand U2816 (N_2816,N_2783,N_2758);
nand U2817 (N_2817,N_2763,N_2771);
nand U2818 (N_2818,N_2769,N_2779);
nor U2819 (N_2819,N_2791,N_2777);
nor U2820 (N_2820,N_2795,N_2774);
nor U2821 (N_2821,N_2750,N_2766);
or U2822 (N_2822,N_2794,N_2787);
nor U2823 (N_2823,N_2788,N_2764);
nand U2824 (N_2824,N_2761,N_2784);
or U2825 (N_2825,N_2754,N_2777);
nand U2826 (N_2826,N_2761,N_2774);
nand U2827 (N_2827,N_2786,N_2797);
nor U2828 (N_2828,N_2762,N_2760);
and U2829 (N_2829,N_2791,N_2766);
and U2830 (N_2830,N_2790,N_2758);
nand U2831 (N_2831,N_2775,N_2754);
nand U2832 (N_2832,N_2758,N_2771);
or U2833 (N_2833,N_2758,N_2752);
nor U2834 (N_2834,N_2781,N_2788);
nor U2835 (N_2835,N_2798,N_2768);
or U2836 (N_2836,N_2784,N_2785);
nand U2837 (N_2837,N_2783,N_2799);
and U2838 (N_2838,N_2766,N_2775);
nor U2839 (N_2839,N_2750,N_2792);
nor U2840 (N_2840,N_2797,N_2751);
or U2841 (N_2841,N_2773,N_2780);
nor U2842 (N_2842,N_2770,N_2788);
nand U2843 (N_2843,N_2761,N_2779);
and U2844 (N_2844,N_2765,N_2769);
and U2845 (N_2845,N_2758,N_2767);
nand U2846 (N_2846,N_2784,N_2790);
and U2847 (N_2847,N_2792,N_2751);
or U2848 (N_2848,N_2776,N_2750);
nand U2849 (N_2849,N_2782,N_2766);
nand U2850 (N_2850,N_2805,N_2818);
or U2851 (N_2851,N_2804,N_2839);
or U2852 (N_2852,N_2811,N_2849);
or U2853 (N_2853,N_2822,N_2840);
nor U2854 (N_2854,N_2830,N_2803);
and U2855 (N_2855,N_2820,N_2843);
or U2856 (N_2856,N_2819,N_2825);
and U2857 (N_2857,N_2832,N_2814);
nor U2858 (N_2858,N_2801,N_2826);
and U2859 (N_2859,N_2824,N_2834);
and U2860 (N_2860,N_2812,N_2847);
nand U2861 (N_2861,N_2844,N_2848);
and U2862 (N_2862,N_2823,N_2836);
nand U2863 (N_2863,N_2800,N_2807);
and U2864 (N_2864,N_2845,N_2821);
and U2865 (N_2865,N_2810,N_2829);
and U2866 (N_2866,N_2831,N_2817);
or U2867 (N_2867,N_2816,N_2806);
and U2868 (N_2868,N_2841,N_2828);
and U2869 (N_2869,N_2835,N_2833);
or U2870 (N_2870,N_2815,N_2808);
nor U2871 (N_2871,N_2802,N_2827);
nor U2872 (N_2872,N_2813,N_2838);
nand U2873 (N_2873,N_2809,N_2842);
nand U2874 (N_2874,N_2837,N_2846);
nand U2875 (N_2875,N_2817,N_2821);
nand U2876 (N_2876,N_2808,N_2807);
or U2877 (N_2877,N_2834,N_2815);
or U2878 (N_2878,N_2811,N_2808);
nor U2879 (N_2879,N_2804,N_2837);
nor U2880 (N_2880,N_2802,N_2810);
or U2881 (N_2881,N_2829,N_2808);
nand U2882 (N_2882,N_2826,N_2811);
nor U2883 (N_2883,N_2830,N_2839);
nand U2884 (N_2884,N_2834,N_2822);
nand U2885 (N_2885,N_2848,N_2824);
or U2886 (N_2886,N_2813,N_2819);
or U2887 (N_2887,N_2841,N_2821);
and U2888 (N_2888,N_2832,N_2847);
or U2889 (N_2889,N_2841,N_2820);
nor U2890 (N_2890,N_2812,N_2828);
or U2891 (N_2891,N_2843,N_2849);
nor U2892 (N_2892,N_2823,N_2816);
and U2893 (N_2893,N_2808,N_2831);
or U2894 (N_2894,N_2811,N_2836);
and U2895 (N_2895,N_2844,N_2819);
nand U2896 (N_2896,N_2807,N_2837);
and U2897 (N_2897,N_2810,N_2811);
or U2898 (N_2898,N_2809,N_2838);
or U2899 (N_2899,N_2806,N_2837);
or U2900 (N_2900,N_2866,N_2857);
nand U2901 (N_2901,N_2853,N_2887);
or U2902 (N_2902,N_2873,N_2865);
nor U2903 (N_2903,N_2886,N_2893);
nor U2904 (N_2904,N_2871,N_2891);
and U2905 (N_2905,N_2882,N_2861);
nand U2906 (N_2906,N_2895,N_2898);
or U2907 (N_2907,N_2867,N_2868);
nor U2908 (N_2908,N_2883,N_2869);
nand U2909 (N_2909,N_2856,N_2894);
nor U2910 (N_2910,N_2880,N_2872);
nand U2911 (N_2911,N_2890,N_2881);
or U2912 (N_2912,N_2859,N_2899);
xnor U2913 (N_2913,N_2850,N_2889);
or U2914 (N_2914,N_2884,N_2879);
nor U2915 (N_2915,N_2854,N_2864);
or U2916 (N_2916,N_2892,N_2876);
nor U2917 (N_2917,N_2877,N_2896);
or U2918 (N_2918,N_2860,N_2863);
nor U2919 (N_2919,N_2855,N_2851);
nand U2920 (N_2920,N_2852,N_2870);
or U2921 (N_2921,N_2878,N_2897);
or U2922 (N_2922,N_2858,N_2875);
and U2923 (N_2923,N_2885,N_2874);
nand U2924 (N_2924,N_2862,N_2888);
nor U2925 (N_2925,N_2861,N_2894);
or U2926 (N_2926,N_2862,N_2850);
nor U2927 (N_2927,N_2856,N_2886);
nand U2928 (N_2928,N_2862,N_2851);
nor U2929 (N_2929,N_2866,N_2871);
and U2930 (N_2930,N_2853,N_2855);
nor U2931 (N_2931,N_2851,N_2899);
nor U2932 (N_2932,N_2888,N_2853);
nor U2933 (N_2933,N_2899,N_2897);
and U2934 (N_2934,N_2855,N_2888);
or U2935 (N_2935,N_2862,N_2899);
xnor U2936 (N_2936,N_2878,N_2883);
nor U2937 (N_2937,N_2881,N_2863);
nand U2938 (N_2938,N_2898,N_2854);
xor U2939 (N_2939,N_2862,N_2864);
or U2940 (N_2940,N_2881,N_2874);
nand U2941 (N_2941,N_2896,N_2880);
nor U2942 (N_2942,N_2855,N_2869);
nand U2943 (N_2943,N_2863,N_2882);
nand U2944 (N_2944,N_2879,N_2854);
nand U2945 (N_2945,N_2864,N_2889);
and U2946 (N_2946,N_2859,N_2876);
or U2947 (N_2947,N_2854,N_2878);
nand U2948 (N_2948,N_2857,N_2853);
and U2949 (N_2949,N_2884,N_2899);
nor U2950 (N_2950,N_2945,N_2926);
and U2951 (N_2951,N_2933,N_2938);
xor U2952 (N_2952,N_2923,N_2917);
and U2953 (N_2953,N_2921,N_2919);
nand U2954 (N_2954,N_2928,N_2924);
nand U2955 (N_2955,N_2925,N_2915);
and U2956 (N_2956,N_2922,N_2901);
and U2957 (N_2957,N_2912,N_2946);
nor U2958 (N_2958,N_2927,N_2935);
and U2959 (N_2959,N_2936,N_2939);
and U2960 (N_2960,N_2920,N_2907);
nor U2961 (N_2961,N_2934,N_2905);
nand U2962 (N_2962,N_2941,N_2944);
nand U2963 (N_2963,N_2949,N_2931);
and U2964 (N_2964,N_2932,N_2909);
or U2965 (N_2965,N_2904,N_2913);
or U2966 (N_2966,N_2911,N_2914);
nand U2967 (N_2967,N_2948,N_2916);
or U2968 (N_2968,N_2900,N_2903);
or U2969 (N_2969,N_2908,N_2942);
nand U2970 (N_2970,N_2930,N_2906);
and U2971 (N_2971,N_2929,N_2902);
and U2972 (N_2972,N_2937,N_2947);
nor U2973 (N_2973,N_2940,N_2943);
or U2974 (N_2974,N_2918,N_2910);
nor U2975 (N_2975,N_2933,N_2915);
nor U2976 (N_2976,N_2916,N_2903);
and U2977 (N_2977,N_2916,N_2900);
nor U2978 (N_2978,N_2920,N_2917);
nand U2979 (N_2979,N_2949,N_2905);
nand U2980 (N_2980,N_2927,N_2930);
nand U2981 (N_2981,N_2926,N_2944);
and U2982 (N_2982,N_2929,N_2907);
and U2983 (N_2983,N_2946,N_2922);
or U2984 (N_2984,N_2946,N_2909);
and U2985 (N_2985,N_2938,N_2903);
and U2986 (N_2986,N_2912,N_2945);
and U2987 (N_2987,N_2938,N_2900);
nand U2988 (N_2988,N_2943,N_2941);
nor U2989 (N_2989,N_2930,N_2945);
and U2990 (N_2990,N_2904,N_2919);
nand U2991 (N_2991,N_2925,N_2927);
nor U2992 (N_2992,N_2917,N_2902);
nand U2993 (N_2993,N_2936,N_2932);
nor U2994 (N_2994,N_2947,N_2912);
or U2995 (N_2995,N_2912,N_2916);
nand U2996 (N_2996,N_2930,N_2948);
or U2997 (N_2997,N_2922,N_2945);
nor U2998 (N_2998,N_2904,N_2940);
xnor U2999 (N_2999,N_2928,N_2906);
nor UO_0 (O_0,N_2974,N_2982);
nand UO_1 (O_1,N_2956,N_2970);
and UO_2 (O_2,N_2960,N_2988);
or UO_3 (O_3,N_2975,N_2992);
nor UO_4 (O_4,N_2971,N_2957);
or UO_5 (O_5,N_2991,N_2998);
or UO_6 (O_6,N_2973,N_2996);
or UO_7 (O_7,N_2961,N_2980);
and UO_8 (O_8,N_2997,N_2950);
nor UO_9 (O_9,N_2999,N_2954);
and UO_10 (O_10,N_2993,N_2994);
nand UO_11 (O_11,N_2990,N_2964);
and UO_12 (O_12,N_2977,N_2962);
and UO_13 (O_13,N_2995,N_2987);
or UO_14 (O_14,N_2958,N_2984);
nor UO_15 (O_15,N_2953,N_2981);
nand UO_16 (O_16,N_2985,N_2969);
nand UO_17 (O_17,N_2967,N_2965);
nand UO_18 (O_18,N_2959,N_2955);
or UO_19 (O_19,N_2983,N_2986);
nand UO_20 (O_20,N_2976,N_2963);
and UO_21 (O_21,N_2972,N_2979);
nor UO_22 (O_22,N_2989,N_2951);
or UO_23 (O_23,N_2968,N_2952);
and UO_24 (O_24,N_2978,N_2966);
or UO_25 (O_25,N_2972,N_2981);
nand UO_26 (O_26,N_2981,N_2988);
nand UO_27 (O_27,N_2984,N_2961);
and UO_28 (O_28,N_2969,N_2968);
nor UO_29 (O_29,N_2951,N_2961);
nor UO_30 (O_30,N_2994,N_2969);
and UO_31 (O_31,N_2966,N_2994);
and UO_32 (O_32,N_2986,N_2974);
or UO_33 (O_33,N_2984,N_2978);
or UO_34 (O_34,N_2959,N_2954);
nand UO_35 (O_35,N_2967,N_2955);
nand UO_36 (O_36,N_2979,N_2954);
and UO_37 (O_37,N_2983,N_2956);
nand UO_38 (O_38,N_2982,N_2966);
and UO_39 (O_39,N_2956,N_2954);
or UO_40 (O_40,N_2950,N_2973);
nand UO_41 (O_41,N_2997,N_2991);
nor UO_42 (O_42,N_2968,N_2999);
nand UO_43 (O_43,N_2997,N_2964);
nor UO_44 (O_44,N_2993,N_2957);
nand UO_45 (O_45,N_2965,N_2959);
nor UO_46 (O_46,N_2980,N_2970);
nor UO_47 (O_47,N_2979,N_2990);
nand UO_48 (O_48,N_2953,N_2972);
nor UO_49 (O_49,N_2970,N_2972);
and UO_50 (O_50,N_2981,N_2958);
nand UO_51 (O_51,N_2975,N_2980);
or UO_52 (O_52,N_2992,N_2981);
nor UO_53 (O_53,N_2986,N_2987);
nor UO_54 (O_54,N_2961,N_2965);
or UO_55 (O_55,N_2985,N_2980);
nor UO_56 (O_56,N_2969,N_2977);
or UO_57 (O_57,N_2986,N_2950);
nor UO_58 (O_58,N_2987,N_2966);
or UO_59 (O_59,N_2986,N_2953);
nand UO_60 (O_60,N_2974,N_2996);
or UO_61 (O_61,N_2990,N_2957);
and UO_62 (O_62,N_2952,N_2982);
or UO_63 (O_63,N_2966,N_2950);
and UO_64 (O_64,N_2991,N_2962);
nor UO_65 (O_65,N_2975,N_2968);
nor UO_66 (O_66,N_2956,N_2984);
nand UO_67 (O_67,N_2955,N_2972);
nor UO_68 (O_68,N_2973,N_2955);
nor UO_69 (O_69,N_2964,N_2976);
nor UO_70 (O_70,N_2986,N_2959);
and UO_71 (O_71,N_2984,N_2993);
nor UO_72 (O_72,N_2983,N_2989);
nor UO_73 (O_73,N_2961,N_2987);
nand UO_74 (O_74,N_2963,N_2954);
or UO_75 (O_75,N_2971,N_2987);
nand UO_76 (O_76,N_2993,N_2967);
nor UO_77 (O_77,N_2988,N_2978);
nand UO_78 (O_78,N_2978,N_2956);
xor UO_79 (O_79,N_2965,N_2987);
or UO_80 (O_80,N_2978,N_2990);
or UO_81 (O_81,N_2991,N_2950);
or UO_82 (O_82,N_2962,N_2986);
nand UO_83 (O_83,N_2988,N_2963);
nand UO_84 (O_84,N_2994,N_2982);
or UO_85 (O_85,N_2963,N_2972);
or UO_86 (O_86,N_2973,N_2969);
and UO_87 (O_87,N_2959,N_2973);
nand UO_88 (O_88,N_2957,N_2970);
nand UO_89 (O_89,N_2979,N_2956);
and UO_90 (O_90,N_2991,N_2988);
nor UO_91 (O_91,N_2978,N_2968);
nand UO_92 (O_92,N_2968,N_2987);
nand UO_93 (O_93,N_2971,N_2981);
nor UO_94 (O_94,N_2960,N_2982);
nand UO_95 (O_95,N_2980,N_2965);
nand UO_96 (O_96,N_2991,N_2956);
nor UO_97 (O_97,N_2966,N_2988);
nor UO_98 (O_98,N_2983,N_2954);
or UO_99 (O_99,N_2962,N_2988);
nand UO_100 (O_100,N_2982,N_2954);
nor UO_101 (O_101,N_2992,N_2976);
nand UO_102 (O_102,N_2998,N_2995);
or UO_103 (O_103,N_2991,N_2969);
nand UO_104 (O_104,N_2954,N_2995);
nor UO_105 (O_105,N_2953,N_2976);
or UO_106 (O_106,N_2972,N_2956);
nand UO_107 (O_107,N_2960,N_2961);
nand UO_108 (O_108,N_2967,N_2976);
nand UO_109 (O_109,N_2985,N_2961);
or UO_110 (O_110,N_2977,N_2963);
and UO_111 (O_111,N_2981,N_2961);
nor UO_112 (O_112,N_2950,N_2955);
nor UO_113 (O_113,N_2962,N_2984);
nor UO_114 (O_114,N_2974,N_2968);
nand UO_115 (O_115,N_2961,N_2955);
and UO_116 (O_116,N_2967,N_2986);
or UO_117 (O_117,N_2992,N_2984);
and UO_118 (O_118,N_2958,N_2971);
nor UO_119 (O_119,N_2974,N_2963);
and UO_120 (O_120,N_2995,N_2975);
nand UO_121 (O_121,N_2962,N_2978);
nand UO_122 (O_122,N_2956,N_2958);
nand UO_123 (O_123,N_2953,N_2995);
or UO_124 (O_124,N_2959,N_2989);
nand UO_125 (O_125,N_2976,N_2994);
nand UO_126 (O_126,N_2962,N_2994);
or UO_127 (O_127,N_2975,N_2971);
and UO_128 (O_128,N_2992,N_2964);
nand UO_129 (O_129,N_2954,N_2993);
or UO_130 (O_130,N_2988,N_2953);
nand UO_131 (O_131,N_2952,N_2954);
nand UO_132 (O_132,N_2962,N_2964);
and UO_133 (O_133,N_2964,N_2995);
nor UO_134 (O_134,N_2970,N_2981);
nand UO_135 (O_135,N_2965,N_2983);
and UO_136 (O_136,N_2968,N_2986);
and UO_137 (O_137,N_2976,N_2951);
and UO_138 (O_138,N_2975,N_2997);
nor UO_139 (O_139,N_2985,N_2991);
and UO_140 (O_140,N_2982,N_2978);
and UO_141 (O_141,N_2978,N_2972);
xor UO_142 (O_142,N_2982,N_2951);
and UO_143 (O_143,N_2972,N_2967);
nand UO_144 (O_144,N_2972,N_2986);
nor UO_145 (O_145,N_2988,N_2990);
and UO_146 (O_146,N_2959,N_2993);
nor UO_147 (O_147,N_2975,N_2979);
nor UO_148 (O_148,N_2960,N_2957);
and UO_149 (O_149,N_2955,N_2970);
and UO_150 (O_150,N_2980,N_2979);
xnor UO_151 (O_151,N_2998,N_2985);
nor UO_152 (O_152,N_2998,N_2952);
or UO_153 (O_153,N_2976,N_2950);
nor UO_154 (O_154,N_2954,N_2996);
nor UO_155 (O_155,N_2991,N_2975);
nand UO_156 (O_156,N_2968,N_2993);
or UO_157 (O_157,N_2992,N_2985);
nand UO_158 (O_158,N_2981,N_2994);
and UO_159 (O_159,N_2974,N_2987);
or UO_160 (O_160,N_2960,N_2970);
and UO_161 (O_161,N_2964,N_2960);
and UO_162 (O_162,N_2975,N_2950);
and UO_163 (O_163,N_2996,N_2953);
or UO_164 (O_164,N_2994,N_2992);
or UO_165 (O_165,N_2978,N_2963);
nor UO_166 (O_166,N_2969,N_2960);
or UO_167 (O_167,N_2954,N_2991);
nor UO_168 (O_168,N_2960,N_2986);
and UO_169 (O_169,N_2970,N_2998);
nand UO_170 (O_170,N_2978,N_2976);
nand UO_171 (O_171,N_2951,N_2999);
nor UO_172 (O_172,N_2970,N_2986);
nor UO_173 (O_173,N_2960,N_2991);
and UO_174 (O_174,N_2997,N_2984);
and UO_175 (O_175,N_2962,N_2952);
nor UO_176 (O_176,N_2984,N_2995);
or UO_177 (O_177,N_2986,N_2992);
or UO_178 (O_178,N_2962,N_2998);
and UO_179 (O_179,N_2951,N_2974);
nor UO_180 (O_180,N_2958,N_2991);
nand UO_181 (O_181,N_2952,N_2972);
or UO_182 (O_182,N_2982,N_2975);
nor UO_183 (O_183,N_2954,N_2984);
and UO_184 (O_184,N_2984,N_2964);
nand UO_185 (O_185,N_2995,N_2974);
and UO_186 (O_186,N_2978,N_2965);
or UO_187 (O_187,N_2996,N_2950);
nand UO_188 (O_188,N_2999,N_2992);
nor UO_189 (O_189,N_2983,N_2997);
or UO_190 (O_190,N_2955,N_2956);
nand UO_191 (O_191,N_2979,N_2968);
or UO_192 (O_192,N_2962,N_2967);
nor UO_193 (O_193,N_2969,N_2988);
nand UO_194 (O_194,N_2953,N_2980);
nor UO_195 (O_195,N_2971,N_2988);
or UO_196 (O_196,N_2971,N_2973);
nand UO_197 (O_197,N_2995,N_2979);
and UO_198 (O_198,N_2985,N_2983);
or UO_199 (O_199,N_2956,N_2990);
nand UO_200 (O_200,N_2999,N_2961);
nor UO_201 (O_201,N_2998,N_2969);
nor UO_202 (O_202,N_2953,N_2961);
nand UO_203 (O_203,N_2992,N_2954);
or UO_204 (O_204,N_2986,N_2969);
nor UO_205 (O_205,N_2956,N_2982);
or UO_206 (O_206,N_2998,N_2987);
or UO_207 (O_207,N_2965,N_2998);
nor UO_208 (O_208,N_2996,N_2981);
nand UO_209 (O_209,N_2958,N_2985);
nor UO_210 (O_210,N_2974,N_2977);
nand UO_211 (O_211,N_2958,N_2989);
nor UO_212 (O_212,N_2958,N_2962);
or UO_213 (O_213,N_2986,N_2985);
and UO_214 (O_214,N_2962,N_2976);
xnor UO_215 (O_215,N_2952,N_2958);
and UO_216 (O_216,N_2994,N_2963);
xor UO_217 (O_217,N_2969,N_2951);
nor UO_218 (O_218,N_2977,N_2989);
and UO_219 (O_219,N_2953,N_2963);
or UO_220 (O_220,N_2980,N_2959);
or UO_221 (O_221,N_2969,N_2980);
nand UO_222 (O_222,N_2963,N_2984);
nand UO_223 (O_223,N_2976,N_2955);
xor UO_224 (O_224,N_2956,N_2988);
and UO_225 (O_225,N_2988,N_2974);
nand UO_226 (O_226,N_2998,N_2976);
or UO_227 (O_227,N_2974,N_2994);
and UO_228 (O_228,N_2962,N_2971);
nor UO_229 (O_229,N_2955,N_2980);
and UO_230 (O_230,N_2963,N_2999);
nand UO_231 (O_231,N_2951,N_2964);
and UO_232 (O_232,N_2970,N_2971);
or UO_233 (O_233,N_2968,N_2957);
nand UO_234 (O_234,N_2981,N_2968);
nor UO_235 (O_235,N_2975,N_2962);
or UO_236 (O_236,N_2972,N_2950);
and UO_237 (O_237,N_2985,N_2995);
nand UO_238 (O_238,N_2989,N_2985);
nand UO_239 (O_239,N_2951,N_2960);
or UO_240 (O_240,N_2986,N_2958);
nor UO_241 (O_241,N_2988,N_2964);
nor UO_242 (O_242,N_2965,N_2990);
and UO_243 (O_243,N_2999,N_2990);
nand UO_244 (O_244,N_2970,N_2982);
nand UO_245 (O_245,N_2959,N_2990);
and UO_246 (O_246,N_2997,N_2988);
and UO_247 (O_247,N_2992,N_2983);
and UO_248 (O_248,N_2993,N_2955);
nand UO_249 (O_249,N_2972,N_2997);
or UO_250 (O_250,N_2966,N_2979);
nor UO_251 (O_251,N_2974,N_2969);
or UO_252 (O_252,N_2992,N_2991);
nor UO_253 (O_253,N_2984,N_2998);
nor UO_254 (O_254,N_2962,N_2979);
nand UO_255 (O_255,N_2968,N_2982);
nor UO_256 (O_256,N_2972,N_2991);
nor UO_257 (O_257,N_2990,N_2963);
nand UO_258 (O_258,N_2976,N_2958);
nor UO_259 (O_259,N_2981,N_2969);
nor UO_260 (O_260,N_2998,N_2988);
nor UO_261 (O_261,N_2978,N_2959);
nor UO_262 (O_262,N_2965,N_2952);
and UO_263 (O_263,N_2996,N_2956);
or UO_264 (O_264,N_2986,N_2998);
nand UO_265 (O_265,N_2962,N_2973);
nor UO_266 (O_266,N_2985,N_2975);
nor UO_267 (O_267,N_2961,N_2998);
nor UO_268 (O_268,N_2974,N_2954);
nor UO_269 (O_269,N_2970,N_2962);
or UO_270 (O_270,N_2983,N_2951);
or UO_271 (O_271,N_2989,N_2967);
nand UO_272 (O_272,N_2995,N_2956);
nand UO_273 (O_273,N_2958,N_2998);
nor UO_274 (O_274,N_2966,N_2981);
and UO_275 (O_275,N_2956,N_2998);
nor UO_276 (O_276,N_2974,N_2978);
or UO_277 (O_277,N_2954,N_2961);
or UO_278 (O_278,N_2979,N_2951);
and UO_279 (O_279,N_2974,N_2955);
and UO_280 (O_280,N_2968,N_2954);
nor UO_281 (O_281,N_2971,N_2954);
nor UO_282 (O_282,N_2993,N_2972);
nand UO_283 (O_283,N_2991,N_2996);
nand UO_284 (O_284,N_2991,N_2994);
or UO_285 (O_285,N_2987,N_2980);
nor UO_286 (O_286,N_2990,N_2993);
and UO_287 (O_287,N_2957,N_2964);
nor UO_288 (O_288,N_2986,N_2978);
and UO_289 (O_289,N_2996,N_2986);
and UO_290 (O_290,N_2962,N_2997);
and UO_291 (O_291,N_2959,N_2981);
and UO_292 (O_292,N_2952,N_2997);
and UO_293 (O_293,N_2997,N_2951);
or UO_294 (O_294,N_2990,N_2952);
and UO_295 (O_295,N_2977,N_2972);
nand UO_296 (O_296,N_2993,N_2989);
and UO_297 (O_297,N_2956,N_2973);
and UO_298 (O_298,N_2979,N_2976);
nor UO_299 (O_299,N_2996,N_2958);
nor UO_300 (O_300,N_2973,N_2974);
and UO_301 (O_301,N_2994,N_2967);
nor UO_302 (O_302,N_2964,N_2968);
or UO_303 (O_303,N_2960,N_2955);
nor UO_304 (O_304,N_2952,N_2993);
nand UO_305 (O_305,N_2971,N_2974);
xnor UO_306 (O_306,N_2961,N_2969);
nand UO_307 (O_307,N_2999,N_2971);
and UO_308 (O_308,N_2995,N_2997);
and UO_309 (O_309,N_2983,N_2979);
nor UO_310 (O_310,N_2967,N_2950);
nand UO_311 (O_311,N_2963,N_2980);
nand UO_312 (O_312,N_2992,N_2958);
and UO_313 (O_313,N_2995,N_2951);
or UO_314 (O_314,N_2952,N_2995);
or UO_315 (O_315,N_2999,N_2965);
or UO_316 (O_316,N_2979,N_2994);
nor UO_317 (O_317,N_2956,N_2968);
nand UO_318 (O_318,N_2962,N_2957);
and UO_319 (O_319,N_2950,N_2990);
and UO_320 (O_320,N_2950,N_2965);
nand UO_321 (O_321,N_2987,N_2994);
nand UO_322 (O_322,N_2959,N_2983);
and UO_323 (O_323,N_2980,N_2976);
and UO_324 (O_324,N_2977,N_2983);
nand UO_325 (O_325,N_2950,N_2989);
and UO_326 (O_326,N_2950,N_2992);
nand UO_327 (O_327,N_2964,N_2959);
or UO_328 (O_328,N_2970,N_2996);
nand UO_329 (O_329,N_2996,N_2971);
nand UO_330 (O_330,N_2990,N_2976);
nor UO_331 (O_331,N_2987,N_2984);
nand UO_332 (O_332,N_2966,N_2989);
or UO_333 (O_333,N_2958,N_2995);
or UO_334 (O_334,N_2991,N_2977);
and UO_335 (O_335,N_2999,N_2962);
or UO_336 (O_336,N_2952,N_2992);
nor UO_337 (O_337,N_2988,N_2992);
nand UO_338 (O_338,N_2989,N_2956);
or UO_339 (O_339,N_2977,N_2997);
nand UO_340 (O_340,N_2991,N_2964);
or UO_341 (O_341,N_2980,N_2967);
or UO_342 (O_342,N_2982,N_2987);
and UO_343 (O_343,N_2975,N_2978);
or UO_344 (O_344,N_2970,N_2994);
and UO_345 (O_345,N_2969,N_2971);
nor UO_346 (O_346,N_2970,N_2969);
nor UO_347 (O_347,N_2997,N_2993);
and UO_348 (O_348,N_2967,N_2992);
nor UO_349 (O_349,N_2968,N_2965);
and UO_350 (O_350,N_2999,N_2976);
or UO_351 (O_351,N_2981,N_2997);
and UO_352 (O_352,N_2987,N_2958);
and UO_353 (O_353,N_2990,N_2954);
nor UO_354 (O_354,N_2989,N_2976);
nand UO_355 (O_355,N_2972,N_2980);
nand UO_356 (O_356,N_2990,N_2977);
nand UO_357 (O_357,N_2953,N_2992);
or UO_358 (O_358,N_2963,N_2960);
or UO_359 (O_359,N_2988,N_2984);
or UO_360 (O_360,N_2995,N_2963);
and UO_361 (O_361,N_2998,N_2994);
and UO_362 (O_362,N_2960,N_2975);
and UO_363 (O_363,N_2991,N_2993);
nand UO_364 (O_364,N_2980,N_2958);
nand UO_365 (O_365,N_2974,N_2979);
nor UO_366 (O_366,N_2953,N_2965);
or UO_367 (O_367,N_2996,N_2952);
and UO_368 (O_368,N_2978,N_2979);
and UO_369 (O_369,N_2959,N_2977);
nand UO_370 (O_370,N_2983,N_2970);
and UO_371 (O_371,N_2974,N_2953);
or UO_372 (O_372,N_2975,N_2994);
and UO_373 (O_373,N_2962,N_2951);
nor UO_374 (O_374,N_2962,N_2980);
or UO_375 (O_375,N_2969,N_2983);
and UO_376 (O_376,N_2951,N_2959);
nor UO_377 (O_377,N_2962,N_2966);
and UO_378 (O_378,N_2963,N_2959);
nor UO_379 (O_379,N_2999,N_2986);
nand UO_380 (O_380,N_2973,N_2975);
nor UO_381 (O_381,N_2984,N_2955);
nand UO_382 (O_382,N_2965,N_2972);
and UO_383 (O_383,N_2964,N_2965);
or UO_384 (O_384,N_2955,N_2965);
and UO_385 (O_385,N_2981,N_2998);
nand UO_386 (O_386,N_2987,N_2954);
nand UO_387 (O_387,N_2955,N_2991);
or UO_388 (O_388,N_2959,N_2975);
nand UO_389 (O_389,N_2995,N_2993);
nand UO_390 (O_390,N_2998,N_2951);
nor UO_391 (O_391,N_2951,N_2996);
or UO_392 (O_392,N_2957,N_2985);
nand UO_393 (O_393,N_2969,N_2995);
nor UO_394 (O_394,N_2985,N_2966);
or UO_395 (O_395,N_2966,N_2969);
nor UO_396 (O_396,N_2973,N_2983);
and UO_397 (O_397,N_2988,N_2994);
nand UO_398 (O_398,N_2977,N_2982);
nor UO_399 (O_399,N_2991,N_2989);
or UO_400 (O_400,N_2969,N_2976);
nor UO_401 (O_401,N_2953,N_2956);
nand UO_402 (O_402,N_2992,N_2957);
nand UO_403 (O_403,N_2967,N_2978);
or UO_404 (O_404,N_2972,N_2975);
or UO_405 (O_405,N_2998,N_2955);
or UO_406 (O_406,N_2998,N_2983);
nand UO_407 (O_407,N_2998,N_2977);
or UO_408 (O_408,N_2988,N_2993);
and UO_409 (O_409,N_2967,N_2969);
and UO_410 (O_410,N_2963,N_2970);
and UO_411 (O_411,N_2999,N_2987);
or UO_412 (O_412,N_2972,N_2992);
nand UO_413 (O_413,N_2986,N_2993);
or UO_414 (O_414,N_2998,N_2974);
nor UO_415 (O_415,N_2994,N_2954);
or UO_416 (O_416,N_2951,N_2967);
and UO_417 (O_417,N_2977,N_2958);
nand UO_418 (O_418,N_2983,N_2981);
or UO_419 (O_419,N_2958,N_2973);
and UO_420 (O_420,N_2988,N_2976);
and UO_421 (O_421,N_2961,N_2952);
nor UO_422 (O_422,N_2983,N_2972);
nand UO_423 (O_423,N_2984,N_2969);
nor UO_424 (O_424,N_2979,N_2982);
nand UO_425 (O_425,N_2953,N_2957);
and UO_426 (O_426,N_2994,N_2984);
and UO_427 (O_427,N_2951,N_2994);
or UO_428 (O_428,N_2963,N_2986);
nand UO_429 (O_429,N_2990,N_2962);
nand UO_430 (O_430,N_2968,N_2972);
nand UO_431 (O_431,N_2999,N_2984);
or UO_432 (O_432,N_2978,N_2970);
nor UO_433 (O_433,N_2999,N_2955);
or UO_434 (O_434,N_2996,N_2972);
nor UO_435 (O_435,N_2974,N_2992);
and UO_436 (O_436,N_2964,N_2994);
nand UO_437 (O_437,N_2981,N_2952);
nor UO_438 (O_438,N_2967,N_2979);
or UO_439 (O_439,N_2990,N_2970);
nor UO_440 (O_440,N_2996,N_2969);
nor UO_441 (O_441,N_2955,N_2966);
and UO_442 (O_442,N_2959,N_2971);
or UO_443 (O_443,N_2968,N_2989);
or UO_444 (O_444,N_2976,N_2957);
nand UO_445 (O_445,N_2955,N_2982);
nor UO_446 (O_446,N_2993,N_2999);
nand UO_447 (O_447,N_2976,N_2995);
nand UO_448 (O_448,N_2980,N_2974);
or UO_449 (O_449,N_2981,N_2963);
and UO_450 (O_450,N_2965,N_2976);
and UO_451 (O_451,N_2971,N_2968);
xor UO_452 (O_452,N_2954,N_2977);
or UO_453 (O_453,N_2980,N_2952);
nand UO_454 (O_454,N_2996,N_2998);
and UO_455 (O_455,N_2970,N_2961);
and UO_456 (O_456,N_2955,N_2995);
nor UO_457 (O_457,N_2966,N_2963);
nand UO_458 (O_458,N_2972,N_2990);
and UO_459 (O_459,N_2992,N_2965);
or UO_460 (O_460,N_2972,N_2988);
nor UO_461 (O_461,N_2959,N_2957);
nor UO_462 (O_462,N_2971,N_2976);
or UO_463 (O_463,N_2975,N_2957);
nor UO_464 (O_464,N_2964,N_2979);
and UO_465 (O_465,N_2988,N_2952);
or UO_466 (O_466,N_2987,N_2962);
xor UO_467 (O_467,N_2955,N_2987);
nand UO_468 (O_468,N_2978,N_2997);
or UO_469 (O_469,N_2970,N_2991);
or UO_470 (O_470,N_2988,N_2965);
or UO_471 (O_471,N_2999,N_2981);
nor UO_472 (O_472,N_2954,N_2980);
or UO_473 (O_473,N_2989,N_2970);
and UO_474 (O_474,N_2990,N_2967);
and UO_475 (O_475,N_2990,N_2969);
nor UO_476 (O_476,N_2963,N_2983);
and UO_477 (O_477,N_2970,N_2992);
or UO_478 (O_478,N_2963,N_2965);
nand UO_479 (O_479,N_2968,N_2950);
nor UO_480 (O_480,N_2974,N_2997);
or UO_481 (O_481,N_2997,N_2954);
and UO_482 (O_482,N_2999,N_2956);
or UO_483 (O_483,N_2962,N_2995);
nor UO_484 (O_484,N_2989,N_2962);
nand UO_485 (O_485,N_2952,N_2977);
or UO_486 (O_486,N_2950,N_2971);
and UO_487 (O_487,N_2960,N_2959);
nor UO_488 (O_488,N_2983,N_2991);
or UO_489 (O_489,N_2997,N_2980);
or UO_490 (O_490,N_2997,N_2961);
nor UO_491 (O_491,N_2978,N_2995);
nor UO_492 (O_492,N_2960,N_2996);
or UO_493 (O_493,N_2966,N_2991);
or UO_494 (O_494,N_2973,N_2961);
nor UO_495 (O_495,N_2963,N_2964);
nand UO_496 (O_496,N_2970,N_2979);
nand UO_497 (O_497,N_2958,N_2990);
or UO_498 (O_498,N_2997,N_2970);
nor UO_499 (O_499,N_2958,N_2970);
endmodule