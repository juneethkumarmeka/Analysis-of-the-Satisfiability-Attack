module basic_500_3000_500_5_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_102,In_0);
nand U1 (N_1,In_202,In_146);
or U2 (N_2,In_217,In_397);
nand U3 (N_3,In_280,In_398);
or U4 (N_4,In_55,In_124);
or U5 (N_5,In_471,In_76);
nand U6 (N_6,In_433,In_100);
xnor U7 (N_7,In_497,In_449);
xor U8 (N_8,In_261,In_253);
or U9 (N_9,In_1,In_276);
xor U10 (N_10,In_307,In_298);
or U11 (N_11,In_467,In_244);
and U12 (N_12,In_126,In_204);
and U13 (N_13,In_74,In_336);
nor U14 (N_14,In_288,In_189);
and U15 (N_15,In_389,In_360);
nand U16 (N_16,In_291,In_211);
and U17 (N_17,In_195,In_314);
nor U18 (N_18,In_89,In_401);
nor U19 (N_19,In_194,In_64);
nor U20 (N_20,In_82,In_94);
and U21 (N_21,In_366,In_270);
nand U22 (N_22,In_429,In_395);
nor U23 (N_23,In_460,In_453);
xor U24 (N_24,In_410,In_255);
and U25 (N_25,In_425,In_435);
nand U26 (N_26,In_56,In_456);
nor U27 (N_27,In_328,In_411);
nand U28 (N_28,In_125,In_35);
nor U29 (N_29,In_295,In_152);
xnor U30 (N_30,In_220,In_313);
and U31 (N_31,In_231,In_134);
and U32 (N_32,In_485,In_234);
or U33 (N_33,In_308,In_71);
xor U34 (N_34,In_72,In_310);
xnor U35 (N_35,In_495,In_163);
and U36 (N_36,In_451,In_446);
nor U37 (N_37,In_484,In_299);
xnor U38 (N_38,In_454,In_476);
and U39 (N_39,In_116,In_239);
nand U40 (N_40,In_426,In_235);
or U41 (N_41,In_22,In_326);
or U42 (N_42,In_359,In_387);
or U43 (N_43,In_169,In_265);
or U44 (N_44,In_138,In_296);
nand U45 (N_45,In_30,In_370);
or U46 (N_46,In_373,In_148);
or U47 (N_47,In_461,In_334);
nor U48 (N_48,In_90,In_463);
nand U49 (N_49,In_69,In_442);
and U50 (N_50,In_482,In_98);
xor U51 (N_51,In_40,In_251);
xor U52 (N_52,In_242,In_477);
or U53 (N_53,In_187,In_23);
nand U54 (N_54,In_107,In_414);
and U55 (N_55,In_381,In_315);
or U56 (N_56,In_240,In_88);
and U57 (N_57,In_427,In_290);
xor U58 (N_58,In_31,In_147);
nand U59 (N_59,In_120,In_52);
or U60 (N_60,In_440,In_16);
xnor U61 (N_61,In_101,In_237);
nand U62 (N_62,In_306,In_252);
or U63 (N_63,In_149,In_362);
and U64 (N_64,In_340,In_434);
nor U65 (N_65,In_182,In_341);
xor U66 (N_66,In_418,In_208);
xnor U67 (N_67,In_218,In_378);
xor U68 (N_68,In_272,In_85);
nor U69 (N_69,In_26,In_29);
xor U70 (N_70,In_324,In_93);
xnor U71 (N_71,In_99,In_407);
xor U72 (N_72,In_221,In_273);
nor U73 (N_73,In_197,In_171);
and U74 (N_74,In_267,In_110);
xor U75 (N_75,In_376,In_266);
xor U76 (N_76,In_329,In_275);
and U77 (N_77,In_292,In_105);
nor U78 (N_78,In_419,In_281);
xnor U79 (N_79,In_65,In_203);
nor U80 (N_80,In_496,In_6);
and U81 (N_81,In_32,In_229);
or U82 (N_82,In_232,In_351);
xor U83 (N_83,In_175,In_210);
xor U84 (N_84,In_493,In_44);
and U85 (N_85,In_172,In_422);
and U86 (N_86,In_257,In_137);
nor U87 (N_87,In_445,In_75);
xnor U88 (N_88,In_303,In_478);
or U89 (N_89,In_36,In_127);
or U90 (N_90,In_345,In_14);
nand U91 (N_91,In_347,In_153);
or U92 (N_92,In_457,In_103);
and U93 (N_93,In_348,In_25);
or U94 (N_94,In_183,In_489);
and U95 (N_95,In_161,In_46);
or U96 (N_96,In_406,In_135);
nand U97 (N_97,In_186,In_423);
or U98 (N_98,In_198,In_15);
and U99 (N_99,In_11,In_420);
or U100 (N_100,In_188,In_41);
nor U101 (N_101,In_132,In_123);
or U102 (N_102,In_193,In_335);
or U103 (N_103,In_415,In_466);
or U104 (N_104,In_167,In_325);
and U105 (N_105,In_176,In_474);
and U106 (N_106,In_7,In_18);
xnor U107 (N_107,In_122,In_47);
nor U108 (N_108,In_177,In_191);
xor U109 (N_109,In_473,In_151);
nor U110 (N_110,In_439,In_164);
nor U111 (N_111,In_140,In_357);
nand U112 (N_112,In_367,In_54);
or U113 (N_113,In_256,In_154);
and U114 (N_114,In_45,In_58);
nor U115 (N_115,In_196,In_405);
nor U116 (N_116,In_342,In_375);
xnor U117 (N_117,In_27,In_430);
and U118 (N_118,In_213,In_91);
and U119 (N_119,In_403,In_42);
nand U120 (N_120,In_386,In_380);
or U121 (N_121,In_368,In_271);
and U122 (N_122,In_323,In_209);
nor U123 (N_123,In_77,In_67);
xnor U124 (N_124,In_60,In_216);
and U125 (N_125,In_86,In_322);
xor U126 (N_126,In_155,In_113);
nand U127 (N_127,In_309,In_481);
nor U128 (N_128,In_394,In_277);
and U129 (N_129,In_241,In_258);
xor U130 (N_130,In_352,In_417);
nor U131 (N_131,In_480,In_2);
or U132 (N_132,In_79,In_80);
xor U133 (N_133,In_206,In_37);
and U134 (N_134,In_133,In_184);
and U135 (N_135,In_185,In_450);
nor U136 (N_136,In_498,In_28);
nor U137 (N_137,In_259,In_353);
nor U138 (N_138,In_248,In_443);
nand U139 (N_139,In_301,In_374);
xor U140 (N_140,In_83,In_143);
and U141 (N_141,In_379,In_24);
nor U142 (N_142,In_119,In_179);
and U143 (N_143,In_207,In_114);
and U144 (N_144,In_247,In_444);
and U145 (N_145,In_59,In_441);
or U146 (N_146,In_377,In_431);
and U147 (N_147,In_312,In_199);
and U148 (N_148,In_274,In_371);
and U149 (N_149,In_284,In_402);
or U150 (N_150,In_283,In_409);
nor U151 (N_151,In_363,In_21);
or U152 (N_152,In_78,In_319);
nand U153 (N_153,In_10,In_84);
nand U154 (N_154,In_246,In_393);
or U155 (N_155,In_9,In_174);
or U156 (N_156,In_87,In_396);
or U157 (N_157,In_62,In_150);
nor U158 (N_158,In_404,In_160);
nor U159 (N_159,In_285,In_413);
and U160 (N_160,In_162,In_302);
or U161 (N_161,In_5,In_95);
xnor U162 (N_162,In_200,In_364);
and U163 (N_163,In_349,In_487);
xor U164 (N_164,In_63,In_8);
xnor U165 (N_165,In_390,In_156);
or U166 (N_166,In_236,In_282);
xnor U167 (N_167,In_178,In_447);
and U168 (N_168,In_233,In_212);
xor U169 (N_169,In_190,In_412);
xnor U170 (N_170,In_33,In_157);
nor U171 (N_171,In_320,In_262);
or U172 (N_172,In_278,In_486);
and U173 (N_173,In_499,In_392);
nand U174 (N_174,In_205,In_38);
or U175 (N_175,In_475,In_385);
or U176 (N_176,In_317,In_421);
nor U177 (N_177,In_3,In_223);
or U178 (N_178,In_269,In_399);
xor U179 (N_179,In_382,In_459);
nor U180 (N_180,In_142,In_224);
and U181 (N_181,In_343,In_346);
or U182 (N_182,In_372,In_383);
xnor U183 (N_183,In_462,In_51);
nor U184 (N_184,In_311,In_145);
nand U185 (N_185,In_245,In_327);
xor U186 (N_186,In_355,In_264);
xor U187 (N_187,In_168,In_130);
nand U188 (N_188,In_294,In_330);
xnor U189 (N_189,In_339,In_452);
xor U190 (N_190,In_365,In_333);
nand U191 (N_191,In_391,In_469);
and U192 (N_192,In_408,In_458);
nand U193 (N_193,In_289,In_19);
or U194 (N_194,In_260,In_238);
xor U195 (N_195,In_361,In_222);
or U196 (N_196,In_166,In_39);
nand U197 (N_197,In_356,In_226);
and U198 (N_198,In_432,In_490);
nor U199 (N_199,In_424,In_111);
xor U200 (N_200,In_73,In_455);
nor U201 (N_201,In_117,In_49);
or U202 (N_202,In_214,In_57);
and U203 (N_203,In_332,In_141);
nor U204 (N_204,In_465,In_437);
nor U205 (N_205,In_227,In_448);
nand U206 (N_206,In_13,In_263);
and U207 (N_207,In_136,In_472);
or U208 (N_208,In_344,In_384);
or U209 (N_209,In_97,In_304);
xor U210 (N_210,In_121,In_61);
and U211 (N_211,In_12,In_369);
or U212 (N_212,In_192,In_488);
nand U213 (N_213,In_66,In_300);
nor U214 (N_214,In_128,In_20);
nand U215 (N_215,In_109,In_331);
and U216 (N_216,In_165,In_43);
nand U217 (N_217,In_118,In_305);
or U218 (N_218,In_106,In_4);
and U219 (N_219,In_464,In_337);
xor U220 (N_220,In_358,In_388);
and U221 (N_221,In_92,In_159);
nand U222 (N_222,In_470,In_287);
nand U223 (N_223,In_173,In_293);
xnor U224 (N_224,In_479,In_492);
nor U225 (N_225,In_68,In_201);
xnor U226 (N_226,In_243,In_400);
nand U227 (N_227,In_34,In_338);
or U228 (N_228,In_50,In_250);
nor U229 (N_229,In_354,In_321);
or U230 (N_230,In_131,In_17);
and U231 (N_231,In_225,In_228);
xor U232 (N_232,In_104,In_268);
nor U233 (N_233,In_53,In_316);
and U234 (N_234,In_181,In_468);
and U235 (N_235,In_139,In_491);
xor U236 (N_236,In_108,In_254);
nand U237 (N_237,In_249,In_318);
xor U238 (N_238,In_350,In_219);
xor U239 (N_239,In_112,In_96);
xnor U240 (N_240,In_158,In_279);
nor U241 (N_241,In_436,In_180);
nand U242 (N_242,In_115,In_438);
nand U243 (N_243,In_129,In_48);
xor U244 (N_244,In_483,In_81);
xnor U245 (N_245,In_215,In_230);
and U246 (N_246,In_297,In_494);
and U247 (N_247,In_428,In_70);
xor U248 (N_248,In_416,In_286);
xor U249 (N_249,In_170,In_144);
or U250 (N_250,In_40,In_219);
nand U251 (N_251,In_323,In_441);
and U252 (N_252,In_361,In_413);
nand U253 (N_253,In_270,In_235);
nand U254 (N_254,In_379,In_233);
and U255 (N_255,In_22,In_213);
xnor U256 (N_256,In_458,In_405);
nand U257 (N_257,In_263,In_50);
nor U258 (N_258,In_307,In_143);
and U259 (N_259,In_279,In_447);
nor U260 (N_260,In_254,In_158);
nand U261 (N_261,In_383,In_90);
nand U262 (N_262,In_451,In_333);
nand U263 (N_263,In_63,In_419);
and U264 (N_264,In_409,In_62);
and U265 (N_265,In_146,In_176);
and U266 (N_266,In_333,In_354);
nor U267 (N_267,In_355,In_318);
or U268 (N_268,In_473,In_221);
and U269 (N_269,In_453,In_194);
nor U270 (N_270,In_270,In_230);
xor U271 (N_271,In_72,In_59);
nand U272 (N_272,In_232,In_294);
or U273 (N_273,In_247,In_213);
and U274 (N_274,In_400,In_389);
or U275 (N_275,In_233,In_15);
xnor U276 (N_276,In_281,In_139);
xor U277 (N_277,In_240,In_254);
nor U278 (N_278,In_232,In_248);
and U279 (N_279,In_182,In_36);
xnor U280 (N_280,In_139,In_259);
xnor U281 (N_281,In_295,In_402);
nor U282 (N_282,In_188,In_412);
or U283 (N_283,In_307,In_201);
or U284 (N_284,In_175,In_84);
xor U285 (N_285,In_200,In_412);
xor U286 (N_286,In_35,In_287);
nor U287 (N_287,In_254,In_426);
xor U288 (N_288,In_40,In_198);
or U289 (N_289,In_410,In_471);
xnor U290 (N_290,In_393,In_453);
or U291 (N_291,In_47,In_490);
or U292 (N_292,In_341,In_260);
and U293 (N_293,In_459,In_481);
and U294 (N_294,In_432,In_71);
nor U295 (N_295,In_451,In_422);
nand U296 (N_296,In_368,In_86);
and U297 (N_297,In_490,In_488);
or U298 (N_298,In_26,In_22);
and U299 (N_299,In_496,In_212);
nor U300 (N_300,In_114,In_293);
or U301 (N_301,In_446,In_366);
nor U302 (N_302,In_445,In_377);
or U303 (N_303,In_420,In_197);
or U304 (N_304,In_473,In_362);
or U305 (N_305,In_424,In_155);
or U306 (N_306,In_14,In_157);
xor U307 (N_307,In_399,In_297);
or U308 (N_308,In_285,In_243);
xnor U309 (N_309,In_380,In_59);
or U310 (N_310,In_0,In_399);
nor U311 (N_311,In_255,In_199);
and U312 (N_312,In_410,In_411);
xnor U313 (N_313,In_45,In_405);
nor U314 (N_314,In_426,In_300);
nand U315 (N_315,In_427,In_377);
nor U316 (N_316,In_235,In_85);
and U317 (N_317,In_212,In_476);
or U318 (N_318,In_65,In_456);
or U319 (N_319,In_444,In_68);
nand U320 (N_320,In_365,In_260);
nor U321 (N_321,In_294,In_46);
xnor U322 (N_322,In_234,In_182);
nand U323 (N_323,In_171,In_199);
and U324 (N_324,In_150,In_377);
xnor U325 (N_325,In_187,In_34);
nor U326 (N_326,In_124,In_232);
xnor U327 (N_327,In_62,In_380);
or U328 (N_328,In_124,In_81);
or U329 (N_329,In_324,In_159);
xnor U330 (N_330,In_389,In_296);
or U331 (N_331,In_423,In_122);
nor U332 (N_332,In_62,In_291);
nand U333 (N_333,In_319,In_430);
and U334 (N_334,In_187,In_396);
nand U335 (N_335,In_307,In_9);
and U336 (N_336,In_430,In_387);
or U337 (N_337,In_17,In_345);
or U338 (N_338,In_357,In_68);
nor U339 (N_339,In_444,In_201);
or U340 (N_340,In_4,In_44);
or U341 (N_341,In_258,In_89);
xor U342 (N_342,In_132,In_103);
nand U343 (N_343,In_56,In_375);
nand U344 (N_344,In_204,In_203);
nor U345 (N_345,In_202,In_232);
or U346 (N_346,In_280,In_379);
or U347 (N_347,In_22,In_66);
nand U348 (N_348,In_168,In_12);
nand U349 (N_349,In_381,In_278);
xor U350 (N_350,In_99,In_20);
and U351 (N_351,In_259,In_283);
or U352 (N_352,In_165,In_350);
xnor U353 (N_353,In_318,In_220);
nor U354 (N_354,In_254,In_395);
or U355 (N_355,In_224,In_430);
nand U356 (N_356,In_134,In_150);
and U357 (N_357,In_53,In_275);
nor U358 (N_358,In_191,In_249);
nor U359 (N_359,In_10,In_252);
nand U360 (N_360,In_262,In_377);
xnor U361 (N_361,In_45,In_118);
nand U362 (N_362,In_115,In_121);
or U363 (N_363,In_148,In_483);
nand U364 (N_364,In_436,In_375);
or U365 (N_365,In_15,In_288);
xor U366 (N_366,In_83,In_301);
nand U367 (N_367,In_493,In_62);
and U368 (N_368,In_328,In_82);
xnor U369 (N_369,In_317,In_34);
and U370 (N_370,In_158,In_261);
nor U371 (N_371,In_437,In_66);
or U372 (N_372,In_479,In_370);
or U373 (N_373,In_354,In_304);
xnor U374 (N_374,In_63,In_43);
xor U375 (N_375,In_444,In_439);
nand U376 (N_376,In_161,In_124);
or U377 (N_377,In_492,In_325);
nand U378 (N_378,In_55,In_297);
xor U379 (N_379,In_446,In_181);
and U380 (N_380,In_41,In_337);
or U381 (N_381,In_450,In_24);
and U382 (N_382,In_446,In_484);
and U383 (N_383,In_417,In_228);
nand U384 (N_384,In_304,In_221);
nor U385 (N_385,In_481,In_137);
or U386 (N_386,In_319,In_302);
nand U387 (N_387,In_149,In_352);
nand U388 (N_388,In_339,In_248);
xor U389 (N_389,In_303,In_175);
or U390 (N_390,In_21,In_454);
or U391 (N_391,In_159,In_242);
nand U392 (N_392,In_364,In_14);
or U393 (N_393,In_74,In_29);
nand U394 (N_394,In_245,In_469);
and U395 (N_395,In_478,In_489);
xor U396 (N_396,In_76,In_202);
and U397 (N_397,In_48,In_160);
xor U398 (N_398,In_376,In_355);
nand U399 (N_399,In_360,In_337);
nand U400 (N_400,In_161,In_255);
xnor U401 (N_401,In_118,In_32);
nor U402 (N_402,In_444,In_265);
nand U403 (N_403,In_354,In_254);
and U404 (N_404,In_438,In_191);
nor U405 (N_405,In_120,In_9);
nor U406 (N_406,In_452,In_186);
and U407 (N_407,In_476,In_386);
and U408 (N_408,In_68,In_6);
nor U409 (N_409,In_261,In_147);
and U410 (N_410,In_137,In_230);
xor U411 (N_411,In_186,In_266);
and U412 (N_412,In_305,In_480);
xor U413 (N_413,In_349,In_323);
nand U414 (N_414,In_449,In_433);
or U415 (N_415,In_29,In_233);
xnor U416 (N_416,In_459,In_6);
and U417 (N_417,In_328,In_231);
nor U418 (N_418,In_311,In_330);
or U419 (N_419,In_59,In_93);
xor U420 (N_420,In_169,In_412);
xor U421 (N_421,In_233,In_324);
xnor U422 (N_422,In_95,In_415);
or U423 (N_423,In_208,In_260);
nor U424 (N_424,In_124,In_248);
xor U425 (N_425,In_455,In_412);
xnor U426 (N_426,In_7,In_478);
xnor U427 (N_427,In_436,In_325);
nand U428 (N_428,In_252,In_125);
and U429 (N_429,In_39,In_278);
nor U430 (N_430,In_315,In_69);
nor U431 (N_431,In_194,In_401);
nand U432 (N_432,In_353,In_424);
nor U433 (N_433,In_411,In_66);
xor U434 (N_434,In_464,In_52);
and U435 (N_435,In_348,In_491);
nand U436 (N_436,In_232,In_42);
nor U437 (N_437,In_213,In_1);
or U438 (N_438,In_383,In_251);
xor U439 (N_439,In_274,In_426);
and U440 (N_440,In_186,In_215);
or U441 (N_441,In_123,In_475);
and U442 (N_442,In_405,In_259);
xnor U443 (N_443,In_387,In_457);
nand U444 (N_444,In_263,In_313);
nor U445 (N_445,In_154,In_376);
nand U446 (N_446,In_101,In_134);
nand U447 (N_447,In_465,In_348);
nor U448 (N_448,In_152,In_445);
xor U449 (N_449,In_248,In_256);
nor U450 (N_450,In_427,In_175);
and U451 (N_451,In_12,In_266);
xnor U452 (N_452,In_214,In_396);
nand U453 (N_453,In_452,In_157);
or U454 (N_454,In_381,In_110);
or U455 (N_455,In_128,In_146);
and U456 (N_456,In_293,In_116);
and U457 (N_457,In_242,In_216);
or U458 (N_458,In_106,In_408);
and U459 (N_459,In_142,In_495);
nand U460 (N_460,In_140,In_344);
nor U461 (N_461,In_104,In_328);
xnor U462 (N_462,In_325,In_119);
and U463 (N_463,In_418,In_57);
or U464 (N_464,In_362,In_435);
and U465 (N_465,In_449,In_254);
and U466 (N_466,In_199,In_33);
nor U467 (N_467,In_363,In_297);
nand U468 (N_468,In_72,In_22);
nor U469 (N_469,In_57,In_183);
xor U470 (N_470,In_185,In_103);
and U471 (N_471,In_89,In_374);
nor U472 (N_472,In_438,In_300);
nand U473 (N_473,In_257,In_388);
nor U474 (N_474,In_351,In_359);
nand U475 (N_475,In_424,In_178);
and U476 (N_476,In_380,In_433);
and U477 (N_477,In_174,In_181);
xnor U478 (N_478,In_115,In_246);
nor U479 (N_479,In_218,In_485);
and U480 (N_480,In_255,In_219);
and U481 (N_481,In_227,In_112);
or U482 (N_482,In_474,In_155);
nor U483 (N_483,In_49,In_375);
or U484 (N_484,In_193,In_409);
and U485 (N_485,In_453,In_312);
or U486 (N_486,In_305,In_44);
nor U487 (N_487,In_336,In_150);
nor U488 (N_488,In_213,In_240);
xor U489 (N_489,In_82,In_77);
and U490 (N_490,In_366,In_35);
nand U491 (N_491,In_75,In_467);
and U492 (N_492,In_263,In_210);
or U493 (N_493,In_98,In_70);
or U494 (N_494,In_413,In_129);
and U495 (N_495,In_322,In_30);
or U496 (N_496,In_312,In_385);
and U497 (N_497,In_202,In_251);
and U498 (N_498,In_358,In_492);
nor U499 (N_499,In_179,In_389);
nor U500 (N_500,In_164,In_138);
and U501 (N_501,In_475,In_274);
xor U502 (N_502,In_236,In_140);
or U503 (N_503,In_479,In_449);
nor U504 (N_504,In_85,In_65);
xor U505 (N_505,In_33,In_105);
and U506 (N_506,In_128,In_277);
or U507 (N_507,In_247,In_414);
and U508 (N_508,In_443,In_485);
or U509 (N_509,In_135,In_119);
nor U510 (N_510,In_197,In_376);
or U511 (N_511,In_246,In_39);
nand U512 (N_512,In_106,In_231);
nor U513 (N_513,In_114,In_202);
and U514 (N_514,In_49,In_204);
nand U515 (N_515,In_325,In_107);
nand U516 (N_516,In_89,In_464);
or U517 (N_517,In_102,In_342);
or U518 (N_518,In_377,In_157);
nor U519 (N_519,In_216,In_77);
or U520 (N_520,In_104,In_261);
nor U521 (N_521,In_326,In_66);
xor U522 (N_522,In_155,In_349);
xnor U523 (N_523,In_145,In_370);
nand U524 (N_524,In_173,In_287);
or U525 (N_525,In_228,In_316);
xnor U526 (N_526,In_363,In_420);
nand U527 (N_527,In_161,In_214);
xnor U528 (N_528,In_173,In_254);
nand U529 (N_529,In_311,In_300);
nor U530 (N_530,In_294,In_195);
xor U531 (N_531,In_103,In_4);
and U532 (N_532,In_23,In_419);
nor U533 (N_533,In_311,In_253);
xor U534 (N_534,In_397,In_301);
xnor U535 (N_535,In_387,In_375);
xor U536 (N_536,In_228,In_14);
or U537 (N_537,In_219,In_77);
nor U538 (N_538,In_237,In_494);
and U539 (N_539,In_261,In_77);
or U540 (N_540,In_108,In_286);
xor U541 (N_541,In_432,In_118);
nor U542 (N_542,In_118,In_249);
and U543 (N_543,In_291,In_258);
nand U544 (N_544,In_23,In_5);
and U545 (N_545,In_411,In_31);
or U546 (N_546,In_414,In_173);
or U547 (N_547,In_271,In_39);
xor U548 (N_548,In_78,In_49);
or U549 (N_549,In_115,In_137);
xor U550 (N_550,In_155,In_332);
nor U551 (N_551,In_425,In_412);
or U552 (N_552,In_460,In_496);
nor U553 (N_553,In_41,In_310);
or U554 (N_554,In_278,In_222);
xnor U555 (N_555,In_185,In_114);
xor U556 (N_556,In_56,In_75);
nand U557 (N_557,In_182,In_133);
xor U558 (N_558,In_443,In_461);
and U559 (N_559,In_280,In_265);
or U560 (N_560,In_32,In_6);
and U561 (N_561,In_285,In_439);
xor U562 (N_562,In_473,In_320);
or U563 (N_563,In_375,In_28);
or U564 (N_564,In_49,In_196);
xor U565 (N_565,In_444,In_448);
nor U566 (N_566,In_170,In_288);
and U567 (N_567,In_230,In_245);
xor U568 (N_568,In_387,In_272);
nand U569 (N_569,In_236,In_54);
or U570 (N_570,In_245,In_449);
nand U571 (N_571,In_474,In_16);
nand U572 (N_572,In_126,In_309);
xor U573 (N_573,In_230,In_5);
or U574 (N_574,In_77,In_140);
xnor U575 (N_575,In_203,In_444);
xnor U576 (N_576,In_470,In_48);
nor U577 (N_577,In_468,In_41);
nand U578 (N_578,In_284,In_270);
and U579 (N_579,In_472,In_195);
nor U580 (N_580,In_281,In_236);
xnor U581 (N_581,In_58,In_258);
or U582 (N_582,In_499,In_141);
xnor U583 (N_583,In_499,In_67);
or U584 (N_584,In_367,In_183);
xor U585 (N_585,In_157,In_333);
or U586 (N_586,In_477,In_245);
and U587 (N_587,In_192,In_305);
and U588 (N_588,In_77,In_456);
nor U589 (N_589,In_188,In_490);
xnor U590 (N_590,In_186,In_224);
and U591 (N_591,In_399,In_415);
xor U592 (N_592,In_266,In_455);
xor U593 (N_593,In_193,In_188);
nor U594 (N_594,In_73,In_215);
nand U595 (N_595,In_234,In_192);
xor U596 (N_596,In_94,In_93);
xor U597 (N_597,In_369,In_473);
nor U598 (N_598,In_32,In_464);
nand U599 (N_599,In_291,In_371);
nor U600 (N_600,N_73,N_408);
and U601 (N_601,N_483,N_264);
or U602 (N_602,N_143,N_506);
and U603 (N_603,N_135,N_293);
and U604 (N_604,N_580,N_520);
nor U605 (N_605,N_377,N_364);
and U606 (N_606,N_8,N_15);
nor U607 (N_607,N_297,N_204);
xnor U608 (N_608,N_479,N_272);
xnor U609 (N_609,N_395,N_549);
nand U610 (N_610,N_527,N_283);
nor U611 (N_611,N_249,N_501);
or U612 (N_612,N_474,N_446);
xor U613 (N_613,N_512,N_218);
and U614 (N_614,N_548,N_401);
nand U615 (N_615,N_90,N_213);
xnor U616 (N_616,N_544,N_211);
or U617 (N_617,N_255,N_39);
and U618 (N_618,N_329,N_299);
and U619 (N_619,N_107,N_323);
or U620 (N_620,N_239,N_170);
nand U621 (N_621,N_57,N_358);
xor U622 (N_622,N_43,N_71);
nor U623 (N_623,N_351,N_102);
xnor U624 (N_624,N_109,N_275);
nand U625 (N_625,N_509,N_360);
xor U626 (N_626,N_20,N_147);
nor U627 (N_627,N_366,N_407);
and U628 (N_628,N_159,N_592);
or U629 (N_629,N_497,N_139);
xnor U630 (N_630,N_310,N_251);
xnor U631 (N_631,N_182,N_457);
and U632 (N_632,N_270,N_405);
and U633 (N_633,N_210,N_511);
xnor U634 (N_634,N_594,N_243);
or U635 (N_635,N_104,N_30);
nand U636 (N_636,N_37,N_234);
xor U637 (N_637,N_153,N_48);
or U638 (N_638,N_78,N_375);
and U639 (N_639,N_216,N_228);
nor U640 (N_640,N_58,N_498);
xnor U641 (N_641,N_412,N_394);
nor U642 (N_642,N_451,N_562);
or U643 (N_643,N_224,N_36);
or U644 (N_644,N_301,N_522);
xor U645 (N_645,N_595,N_349);
xor U646 (N_646,N_438,N_25);
xnor U647 (N_647,N_123,N_185);
nand U648 (N_648,N_164,N_391);
and U649 (N_649,N_357,N_588);
xnor U650 (N_650,N_574,N_523);
and U651 (N_651,N_140,N_263);
and U652 (N_652,N_440,N_235);
nor U653 (N_653,N_284,N_385);
or U654 (N_654,N_546,N_266);
and U655 (N_655,N_324,N_347);
xor U656 (N_656,N_124,N_97);
nand U657 (N_657,N_274,N_525);
nor U658 (N_658,N_427,N_230);
nor U659 (N_659,N_116,N_47);
xor U660 (N_660,N_286,N_332);
nand U661 (N_661,N_417,N_89);
xnor U662 (N_662,N_543,N_486);
nand U663 (N_663,N_507,N_325);
nand U664 (N_664,N_128,N_484);
and U665 (N_665,N_447,N_376);
nand U666 (N_666,N_277,N_4);
and U667 (N_667,N_160,N_191);
or U668 (N_668,N_584,N_478);
xor U669 (N_669,N_433,N_241);
nor U670 (N_670,N_510,N_19);
xor U671 (N_671,N_261,N_348);
nand U672 (N_672,N_396,N_101);
nand U673 (N_673,N_365,N_133);
nand U674 (N_674,N_345,N_453);
or U675 (N_675,N_537,N_488);
xnor U676 (N_676,N_561,N_17);
or U677 (N_677,N_340,N_529);
nand U678 (N_678,N_473,N_10);
xor U679 (N_679,N_505,N_6);
nor U680 (N_680,N_285,N_398);
and U681 (N_681,N_56,N_445);
nor U682 (N_682,N_0,N_552);
or U683 (N_683,N_186,N_175);
and U684 (N_684,N_196,N_553);
nor U685 (N_685,N_485,N_183);
or U686 (N_686,N_536,N_29);
nand U687 (N_687,N_26,N_156);
xor U688 (N_688,N_125,N_289);
and U689 (N_689,N_384,N_9);
xnor U690 (N_690,N_12,N_45);
or U691 (N_691,N_545,N_226);
and U692 (N_692,N_268,N_113);
and U693 (N_693,N_87,N_23);
and U694 (N_694,N_526,N_62);
nor U695 (N_695,N_161,N_163);
xor U696 (N_696,N_237,N_132);
and U697 (N_697,N_111,N_359);
or U698 (N_698,N_259,N_54);
nor U699 (N_699,N_282,N_246);
and U700 (N_700,N_7,N_406);
nand U701 (N_701,N_343,N_114);
xnor U702 (N_702,N_229,N_491);
nand U703 (N_703,N_294,N_413);
or U704 (N_704,N_141,N_233);
and U705 (N_705,N_292,N_492);
xor U706 (N_706,N_112,N_317);
and U707 (N_707,N_75,N_419);
nand U708 (N_708,N_579,N_311);
nand U709 (N_709,N_55,N_572);
nor U710 (N_710,N_344,N_444);
or U711 (N_711,N_203,N_32);
nand U712 (N_712,N_247,N_475);
and U713 (N_713,N_571,N_421);
xor U714 (N_714,N_110,N_434);
or U715 (N_715,N_180,N_431);
nand U716 (N_716,N_515,N_363);
nand U717 (N_717,N_212,N_381);
nor U718 (N_718,N_157,N_201);
and U719 (N_719,N_312,N_207);
xor U720 (N_720,N_416,N_248);
and U721 (N_721,N_521,N_389);
nand U722 (N_722,N_300,N_287);
nand U723 (N_723,N_350,N_69);
xnor U724 (N_724,N_585,N_16);
nand U725 (N_725,N_296,N_593);
nand U726 (N_726,N_334,N_280);
nor U727 (N_727,N_555,N_302);
or U728 (N_728,N_392,N_319);
xnor U729 (N_729,N_24,N_439);
xnor U730 (N_730,N_198,N_77);
xnor U731 (N_731,N_469,N_72);
xor U732 (N_732,N_200,N_223);
and U733 (N_733,N_590,N_22);
xnor U734 (N_734,N_118,N_414);
nand U735 (N_735,N_468,N_137);
nand U736 (N_736,N_441,N_151);
nand U737 (N_737,N_108,N_91);
nand U738 (N_738,N_291,N_267);
and U739 (N_739,N_99,N_346);
nand U740 (N_740,N_424,N_119);
xnor U741 (N_741,N_60,N_192);
nor U742 (N_742,N_410,N_452);
nor U743 (N_743,N_361,N_217);
and U744 (N_744,N_369,N_477);
nor U745 (N_745,N_70,N_27);
xor U746 (N_746,N_244,N_276);
and U747 (N_747,N_535,N_539);
nand U748 (N_748,N_356,N_463);
nor U749 (N_749,N_74,N_262);
and U750 (N_750,N_298,N_121);
nand U751 (N_751,N_209,N_333);
xor U752 (N_752,N_500,N_155);
nor U753 (N_753,N_13,N_489);
and U754 (N_754,N_245,N_397);
or U755 (N_755,N_308,N_541);
nor U756 (N_756,N_158,N_558);
and U757 (N_757,N_126,N_331);
nand U758 (N_758,N_28,N_481);
or U759 (N_759,N_82,N_557);
nand U760 (N_760,N_464,N_232);
nor U761 (N_761,N_265,N_573);
xnor U762 (N_762,N_459,N_95);
nand U763 (N_763,N_31,N_254);
xnor U764 (N_764,N_465,N_378);
xnor U765 (N_765,N_214,N_250);
or U766 (N_766,N_355,N_220);
or U767 (N_767,N_518,N_21);
nor U768 (N_768,N_542,N_53);
nor U769 (N_769,N_472,N_260);
xor U770 (N_770,N_508,N_171);
nor U771 (N_771,N_50,N_130);
or U772 (N_772,N_46,N_400);
or U773 (N_773,N_456,N_68);
or U774 (N_774,N_448,N_513);
nand U775 (N_775,N_194,N_563);
nand U776 (N_776,N_197,N_168);
nor U777 (N_777,N_547,N_409);
or U778 (N_778,N_52,N_195);
xor U779 (N_779,N_339,N_370);
and U780 (N_780,N_295,N_278);
nand U781 (N_781,N_576,N_252);
nor U782 (N_782,N_63,N_51);
nand U783 (N_783,N_2,N_532);
or U784 (N_784,N_504,N_436);
and U785 (N_785,N_393,N_176);
xnor U786 (N_786,N_190,N_538);
and U787 (N_787,N_503,N_399);
or U788 (N_788,N_181,N_458);
nor U789 (N_789,N_86,N_496);
nand U790 (N_790,N_519,N_5);
and U791 (N_791,N_437,N_368);
or U792 (N_792,N_534,N_582);
nor U793 (N_793,N_142,N_411);
xor U794 (N_794,N_514,N_129);
xnor U795 (N_795,N_383,N_240);
nor U796 (N_796,N_455,N_403);
nand U797 (N_797,N_96,N_425);
or U798 (N_798,N_335,N_65);
and U799 (N_799,N_257,N_84);
and U800 (N_800,N_146,N_40);
or U801 (N_801,N_551,N_597);
or U802 (N_802,N_426,N_253);
nand U803 (N_803,N_460,N_236);
xnor U804 (N_804,N_386,N_388);
xnor U805 (N_805,N_154,N_583);
nand U806 (N_806,N_318,N_569);
nor U807 (N_807,N_428,N_288);
nor U808 (N_808,N_353,N_152);
nor U809 (N_809,N_258,N_178);
nand U810 (N_810,N_336,N_493);
nor U811 (N_811,N_415,N_326);
xnor U812 (N_812,N_305,N_327);
and U813 (N_813,N_367,N_94);
or U814 (N_814,N_131,N_304);
xnor U815 (N_815,N_581,N_322);
or U816 (N_816,N_35,N_379);
or U817 (N_817,N_144,N_120);
nand U818 (N_818,N_578,N_49);
nand U819 (N_819,N_14,N_188);
nor U820 (N_820,N_134,N_462);
nand U821 (N_821,N_315,N_502);
nor U822 (N_822,N_122,N_81);
nor U823 (N_823,N_169,N_174);
nor U824 (N_824,N_61,N_517);
and U825 (N_825,N_1,N_471);
nand U826 (N_826,N_41,N_342);
nand U827 (N_827,N_93,N_443);
nor U828 (N_828,N_575,N_495);
and U829 (N_829,N_256,N_85);
and U830 (N_830,N_150,N_466);
and U831 (N_831,N_172,N_387);
nor U832 (N_832,N_480,N_568);
xor U833 (N_833,N_487,N_442);
nor U834 (N_834,N_596,N_127);
or U835 (N_835,N_162,N_402);
or U836 (N_836,N_225,N_149);
nand U837 (N_837,N_148,N_103);
and U838 (N_838,N_313,N_167);
xnor U839 (N_839,N_117,N_570);
nor U840 (N_840,N_177,N_80);
xnor U841 (N_841,N_33,N_373);
nand U842 (N_842,N_187,N_587);
or U843 (N_843,N_238,N_166);
xor U844 (N_844,N_524,N_18);
nor U845 (N_845,N_11,N_420);
or U846 (N_846,N_106,N_321);
and U847 (N_847,N_461,N_309);
nor U848 (N_848,N_554,N_34);
nand U849 (N_849,N_273,N_222);
or U850 (N_850,N_76,N_432);
nor U851 (N_851,N_316,N_189);
nand U852 (N_852,N_599,N_42);
or U853 (N_853,N_567,N_138);
nor U854 (N_854,N_314,N_476);
xor U855 (N_855,N_550,N_560);
or U856 (N_856,N_450,N_242);
nand U857 (N_857,N_227,N_528);
nor U858 (N_858,N_577,N_430);
and U859 (N_859,N_372,N_184);
xor U860 (N_860,N_374,N_422);
xnor U861 (N_861,N_64,N_206);
or U862 (N_862,N_98,N_59);
xnor U863 (N_863,N_330,N_499);
or U864 (N_864,N_423,N_362);
and U865 (N_865,N_328,N_435);
and U866 (N_866,N_83,N_390);
nor U867 (N_867,N_67,N_165);
nor U868 (N_868,N_559,N_208);
and U869 (N_869,N_115,N_92);
nor U870 (N_870,N_490,N_586);
and U871 (N_871,N_199,N_467);
and U872 (N_872,N_589,N_290);
xor U873 (N_873,N_516,N_79);
or U874 (N_874,N_320,N_145);
nand U875 (N_875,N_556,N_337);
xnor U876 (N_876,N_231,N_281);
and U877 (N_877,N_38,N_566);
xor U878 (N_878,N_540,N_44);
or U879 (N_879,N_565,N_202);
xnor U880 (N_880,N_591,N_338);
xnor U881 (N_881,N_100,N_219);
and U882 (N_882,N_494,N_470);
and U883 (N_883,N_454,N_382);
or U884 (N_884,N_179,N_279);
nand U885 (N_885,N_307,N_341);
and U886 (N_886,N_531,N_105);
or U887 (N_887,N_271,N_371);
or U888 (N_888,N_380,N_66);
and U889 (N_889,N_193,N_418);
and U890 (N_890,N_598,N_3);
nor U891 (N_891,N_215,N_429);
xnor U892 (N_892,N_173,N_221);
nand U893 (N_893,N_269,N_136);
xnor U894 (N_894,N_564,N_404);
xnor U895 (N_895,N_530,N_533);
nor U896 (N_896,N_205,N_352);
and U897 (N_897,N_449,N_306);
nor U898 (N_898,N_354,N_303);
nand U899 (N_899,N_88,N_482);
or U900 (N_900,N_457,N_573);
nor U901 (N_901,N_343,N_146);
xor U902 (N_902,N_225,N_71);
or U903 (N_903,N_292,N_167);
nor U904 (N_904,N_56,N_160);
xnor U905 (N_905,N_281,N_22);
or U906 (N_906,N_150,N_101);
or U907 (N_907,N_252,N_245);
xor U908 (N_908,N_220,N_300);
nor U909 (N_909,N_456,N_493);
and U910 (N_910,N_78,N_562);
xor U911 (N_911,N_409,N_545);
nand U912 (N_912,N_407,N_412);
or U913 (N_913,N_383,N_297);
nor U914 (N_914,N_283,N_77);
or U915 (N_915,N_121,N_553);
nand U916 (N_916,N_406,N_260);
and U917 (N_917,N_486,N_36);
and U918 (N_918,N_154,N_13);
or U919 (N_919,N_254,N_246);
nor U920 (N_920,N_242,N_542);
nand U921 (N_921,N_206,N_544);
nor U922 (N_922,N_99,N_69);
nand U923 (N_923,N_234,N_130);
xnor U924 (N_924,N_518,N_11);
or U925 (N_925,N_311,N_114);
or U926 (N_926,N_225,N_445);
nand U927 (N_927,N_103,N_527);
nand U928 (N_928,N_295,N_89);
xor U929 (N_929,N_290,N_363);
nor U930 (N_930,N_37,N_136);
nand U931 (N_931,N_321,N_236);
nand U932 (N_932,N_484,N_163);
nor U933 (N_933,N_258,N_377);
xor U934 (N_934,N_264,N_571);
or U935 (N_935,N_342,N_246);
and U936 (N_936,N_546,N_421);
nor U937 (N_937,N_53,N_248);
xnor U938 (N_938,N_76,N_16);
xor U939 (N_939,N_562,N_208);
xor U940 (N_940,N_307,N_157);
nor U941 (N_941,N_442,N_494);
and U942 (N_942,N_126,N_278);
xnor U943 (N_943,N_330,N_452);
nor U944 (N_944,N_307,N_417);
nor U945 (N_945,N_46,N_516);
xnor U946 (N_946,N_530,N_85);
nand U947 (N_947,N_324,N_192);
or U948 (N_948,N_565,N_290);
xor U949 (N_949,N_539,N_281);
and U950 (N_950,N_375,N_261);
or U951 (N_951,N_175,N_9);
nand U952 (N_952,N_157,N_481);
or U953 (N_953,N_221,N_455);
or U954 (N_954,N_7,N_152);
and U955 (N_955,N_34,N_46);
and U956 (N_956,N_383,N_457);
or U957 (N_957,N_272,N_419);
or U958 (N_958,N_22,N_75);
nand U959 (N_959,N_365,N_89);
and U960 (N_960,N_127,N_504);
xor U961 (N_961,N_192,N_78);
xnor U962 (N_962,N_563,N_228);
and U963 (N_963,N_16,N_466);
nor U964 (N_964,N_106,N_564);
or U965 (N_965,N_241,N_278);
or U966 (N_966,N_268,N_422);
xor U967 (N_967,N_229,N_37);
or U968 (N_968,N_581,N_302);
and U969 (N_969,N_399,N_249);
and U970 (N_970,N_234,N_502);
nand U971 (N_971,N_372,N_128);
or U972 (N_972,N_282,N_196);
xor U973 (N_973,N_486,N_56);
and U974 (N_974,N_98,N_378);
nand U975 (N_975,N_449,N_573);
xor U976 (N_976,N_502,N_100);
xnor U977 (N_977,N_494,N_364);
nand U978 (N_978,N_552,N_461);
xor U979 (N_979,N_389,N_427);
and U980 (N_980,N_356,N_110);
or U981 (N_981,N_599,N_93);
nand U982 (N_982,N_449,N_478);
nor U983 (N_983,N_414,N_456);
or U984 (N_984,N_326,N_412);
and U985 (N_985,N_447,N_466);
and U986 (N_986,N_191,N_564);
nor U987 (N_987,N_2,N_147);
and U988 (N_988,N_146,N_440);
nand U989 (N_989,N_75,N_142);
xor U990 (N_990,N_98,N_56);
nor U991 (N_991,N_115,N_155);
nand U992 (N_992,N_406,N_275);
and U993 (N_993,N_368,N_565);
and U994 (N_994,N_542,N_336);
nand U995 (N_995,N_224,N_340);
nor U996 (N_996,N_536,N_169);
or U997 (N_997,N_44,N_273);
nor U998 (N_998,N_28,N_257);
nor U999 (N_999,N_62,N_165);
or U1000 (N_1000,N_10,N_87);
nand U1001 (N_1001,N_309,N_501);
or U1002 (N_1002,N_431,N_480);
or U1003 (N_1003,N_100,N_107);
nand U1004 (N_1004,N_597,N_390);
xor U1005 (N_1005,N_122,N_306);
and U1006 (N_1006,N_434,N_570);
or U1007 (N_1007,N_352,N_158);
and U1008 (N_1008,N_54,N_514);
nand U1009 (N_1009,N_258,N_200);
xor U1010 (N_1010,N_214,N_186);
nor U1011 (N_1011,N_212,N_203);
xnor U1012 (N_1012,N_211,N_339);
nor U1013 (N_1013,N_136,N_555);
nand U1014 (N_1014,N_50,N_271);
xnor U1015 (N_1015,N_457,N_461);
nor U1016 (N_1016,N_252,N_374);
nor U1017 (N_1017,N_474,N_331);
nand U1018 (N_1018,N_115,N_177);
nand U1019 (N_1019,N_467,N_543);
nand U1020 (N_1020,N_223,N_147);
or U1021 (N_1021,N_373,N_332);
xor U1022 (N_1022,N_376,N_243);
nor U1023 (N_1023,N_479,N_457);
nor U1024 (N_1024,N_110,N_438);
xnor U1025 (N_1025,N_20,N_285);
nand U1026 (N_1026,N_376,N_456);
or U1027 (N_1027,N_390,N_114);
or U1028 (N_1028,N_253,N_528);
and U1029 (N_1029,N_594,N_114);
nand U1030 (N_1030,N_132,N_69);
and U1031 (N_1031,N_184,N_191);
nand U1032 (N_1032,N_321,N_78);
xor U1033 (N_1033,N_33,N_79);
and U1034 (N_1034,N_495,N_278);
nand U1035 (N_1035,N_377,N_472);
nand U1036 (N_1036,N_156,N_309);
nand U1037 (N_1037,N_410,N_510);
nand U1038 (N_1038,N_228,N_101);
nand U1039 (N_1039,N_569,N_63);
nand U1040 (N_1040,N_116,N_551);
nor U1041 (N_1041,N_69,N_70);
xor U1042 (N_1042,N_321,N_45);
xnor U1043 (N_1043,N_442,N_260);
and U1044 (N_1044,N_208,N_46);
nand U1045 (N_1045,N_56,N_549);
nand U1046 (N_1046,N_284,N_371);
xnor U1047 (N_1047,N_312,N_389);
nor U1048 (N_1048,N_199,N_113);
xnor U1049 (N_1049,N_325,N_207);
or U1050 (N_1050,N_148,N_388);
or U1051 (N_1051,N_151,N_93);
and U1052 (N_1052,N_224,N_529);
nor U1053 (N_1053,N_96,N_474);
and U1054 (N_1054,N_521,N_355);
nand U1055 (N_1055,N_263,N_157);
nand U1056 (N_1056,N_465,N_130);
and U1057 (N_1057,N_121,N_388);
or U1058 (N_1058,N_336,N_199);
or U1059 (N_1059,N_139,N_323);
xor U1060 (N_1060,N_401,N_154);
nor U1061 (N_1061,N_290,N_480);
or U1062 (N_1062,N_348,N_293);
or U1063 (N_1063,N_183,N_467);
nand U1064 (N_1064,N_20,N_537);
xor U1065 (N_1065,N_233,N_343);
or U1066 (N_1066,N_495,N_421);
nor U1067 (N_1067,N_168,N_352);
or U1068 (N_1068,N_194,N_472);
xor U1069 (N_1069,N_85,N_583);
nand U1070 (N_1070,N_302,N_512);
nor U1071 (N_1071,N_151,N_34);
and U1072 (N_1072,N_518,N_335);
nand U1073 (N_1073,N_590,N_480);
xor U1074 (N_1074,N_508,N_135);
or U1075 (N_1075,N_184,N_404);
or U1076 (N_1076,N_407,N_496);
and U1077 (N_1077,N_270,N_493);
xnor U1078 (N_1078,N_583,N_500);
and U1079 (N_1079,N_180,N_566);
xnor U1080 (N_1080,N_41,N_184);
xnor U1081 (N_1081,N_440,N_295);
and U1082 (N_1082,N_443,N_55);
nand U1083 (N_1083,N_412,N_314);
and U1084 (N_1084,N_167,N_510);
nor U1085 (N_1085,N_162,N_289);
nor U1086 (N_1086,N_272,N_498);
xnor U1087 (N_1087,N_1,N_182);
nand U1088 (N_1088,N_211,N_529);
nand U1089 (N_1089,N_228,N_490);
and U1090 (N_1090,N_367,N_476);
nand U1091 (N_1091,N_218,N_157);
nand U1092 (N_1092,N_101,N_548);
and U1093 (N_1093,N_528,N_244);
or U1094 (N_1094,N_104,N_83);
xor U1095 (N_1095,N_448,N_311);
nor U1096 (N_1096,N_143,N_220);
or U1097 (N_1097,N_119,N_270);
nor U1098 (N_1098,N_335,N_467);
and U1099 (N_1099,N_292,N_488);
nand U1100 (N_1100,N_276,N_318);
nor U1101 (N_1101,N_323,N_374);
nand U1102 (N_1102,N_334,N_541);
nand U1103 (N_1103,N_439,N_37);
nor U1104 (N_1104,N_40,N_185);
nand U1105 (N_1105,N_7,N_19);
and U1106 (N_1106,N_596,N_149);
or U1107 (N_1107,N_333,N_266);
nor U1108 (N_1108,N_132,N_160);
and U1109 (N_1109,N_257,N_143);
nor U1110 (N_1110,N_591,N_363);
nand U1111 (N_1111,N_149,N_401);
and U1112 (N_1112,N_44,N_85);
or U1113 (N_1113,N_74,N_537);
nand U1114 (N_1114,N_59,N_439);
xor U1115 (N_1115,N_165,N_203);
and U1116 (N_1116,N_237,N_558);
nor U1117 (N_1117,N_546,N_149);
and U1118 (N_1118,N_505,N_532);
or U1119 (N_1119,N_75,N_27);
nand U1120 (N_1120,N_490,N_374);
nor U1121 (N_1121,N_418,N_0);
and U1122 (N_1122,N_118,N_406);
nand U1123 (N_1123,N_31,N_167);
nand U1124 (N_1124,N_510,N_457);
or U1125 (N_1125,N_308,N_12);
nand U1126 (N_1126,N_222,N_29);
nand U1127 (N_1127,N_450,N_141);
xnor U1128 (N_1128,N_517,N_541);
nor U1129 (N_1129,N_99,N_419);
or U1130 (N_1130,N_388,N_118);
nor U1131 (N_1131,N_163,N_487);
xor U1132 (N_1132,N_486,N_75);
and U1133 (N_1133,N_488,N_0);
nand U1134 (N_1134,N_17,N_441);
nor U1135 (N_1135,N_265,N_181);
and U1136 (N_1136,N_95,N_234);
or U1137 (N_1137,N_1,N_100);
and U1138 (N_1138,N_261,N_70);
nor U1139 (N_1139,N_54,N_440);
or U1140 (N_1140,N_385,N_501);
or U1141 (N_1141,N_241,N_402);
xor U1142 (N_1142,N_265,N_205);
xnor U1143 (N_1143,N_393,N_170);
and U1144 (N_1144,N_274,N_424);
xor U1145 (N_1145,N_373,N_591);
or U1146 (N_1146,N_381,N_565);
xor U1147 (N_1147,N_225,N_95);
nor U1148 (N_1148,N_413,N_42);
and U1149 (N_1149,N_285,N_88);
nor U1150 (N_1150,N_565,N_108);
nand U1151 (N_1151,N_316,N_472);
nor U1152 (N_1152,N_272,N_107);
or U1153 (N_1153,N_360,N_433);
xor U1154 (N_1154,N_157,N_488);
nor U1155 (N_1155,N_374,N_142);
nand U1156 (N_1156,N_13,N_531);
and U1157 (N_1157,N_356,N_163);
and U1158 (N_1158,N_594,N_284);
and U1159 (N_1159,N_177,N_433);
xnor U1160 (N_1160,N_378,N_388);
or U1161 (N_1161,N_491,N_487);
nand U1162 (N_1162,N_469,N_49);
nand U1163 (N_1163,N_416,N_112);
or U1164 (N_1164,N_452,N_351);
nand U1165 (N_1165,N_173,N_530);
and U1166 (N_1166,N_200,N_591);
nor U1167 (N_1167,N_164,N_131);
nor U1168 (N_1168,N_35,N_419);
and U1169 (N_1169,N_171,N_429);
xnor U1170 (N_1170,N_192,N_370);
xor U1171 (N_1171,N_263,N_595);
nor U1172 (N_1172,N_417,N_63);
or U1173 (N_1173,N_211,N_101);
nor U1174 (N_1174,N_435,N_599);
nand U1175 (N_1175,N_85,N_22);
xnor U1176 (N_1176,N_131,N_116);
nand U1177 (N_1177,N_399,N_376);
and U1178 (N_1178,N_199,N_100);
nand U1179 (N_1179,N_106,N_552);
xnor U1180 (N_1180,N_113,N_374);
and U1181 (N_1181,N_452,N_389);
or U1182 (N_1182,N_196,N_399);
nor U1183 (N_1183,N_175,N_329);
nand U1184 (N_1184,N_272,N_70);
nand U1185 (N_1185,N_464,N_577);
and U1186 (N_1186,N_40,N_246);
xor U1187 (N_1187,N_117,N_346);
xnor U1188 (N_1188,N_45,N_556);
or U1189 (N_1189,N_367,N_429);
nand U1190 (N_1190,N_497,N_381);
nor U1191 (N_1191,N_405,N_55);
or U1192 (N_1192,N_449,N_200);
nor U1193 (N_1193,N_99,N_487);
xor U1194 (N_1194,N_488,N_372);
or U1195 (N_1195,N_486,N_138);
and U1196 (N_1196,N_362,N_593);
xor U1197 (N_1197,N_482,N_396);
and U1198 (N_1198,N_77,N_573);
xor U1199 (N_1199,N_296,N_448);
nor U1200 (N_1200,N_1027,N_886);
and U1201 (N_1201,N_720,N_721);
nor U1202 (N_1202,N_961,N_842);
nand U1203 (N_1203,N_1129,N_1183);
or U1204 (N_1204,N_1008,N_667);
nor U1205 (N_1205,N_923,N_1022);
nor U1206 (N_1206,N_1017,N_710);
xnor U1207 (N_1207,N_871,N_782);
nand U1208 (N_1208,N_688,N_1081);
xor U1209 (N_1209,N_724,N_1077);
and U1210 (N_1210,N_1187,N_723);
and U1211 (N_1211,N_905,N_637);
nor U1212 (N_1212,N_821,N_1135);
nand U1213 (N_1213,N_1080,N_948);
or U1214 (N_1214,N_1001,N_830);
nand U1215 (N_1215,N_1009,N_1007);
or U1216 (N_1216,N_715,N_623);
or U1217 (N_1217,N_1145,N_808);
and U1218 (N_1218,N_658,N_1079);
nand U1219 (N_1219,N_747,N_832);
xnor U1220 (N_1220,N_736,N_616);
or U1221 (N_1221,N_659,N_802);
or U1222 (N_1222,N_962,N_1174);
nand U1223 (N_1223,N_761,N_997);
and U1224 (N_1224,N_823,N_986);
and U1225 (N_1225,N_1072,N_1115);
or U1226 (N_1226,N_712,N_977);
xor U1227 (N_1227,N_955,N_838);
nand U1228 (N_1228,N_1128,N_970);
nor U1229 (N_1229,N_1110,N_1157);
or U1230 (N_1230,N_1147,N_765);
nand U1231 (N_1231,N_1020,N_868);
nand U1232 (N_1232,N_1002,N_725);
xor U1233 (N_1233,N_1033,N_922);
nor U1234 (N_1234,N_915,N_770);
or U1235 (N_1235,N_863,N_991);
xor U1236 (N_1236,N_971,N_927);
nor U1237 (N_1237,N_984,N_1182);
and U1238 (N_1238,N_646,N_665);
or U1239 (N_1239,N_1066,N_1124);
nand U1240 (N_1240,N_914,N_1006);
or U1241 (N_1241,N_894,N_1053);
nor U1242 (N_1242,N_714,N_919);
xor U1243 (N_1243,N_632,N_979);
nor U1244 (N_1244,N_1090,N_648);
nand U1245 (N_1245,N_729,N_936);
nand U1246 (N_1246,N_1031,N_898);
xor U1247 (N_1247,N_615,N_760);
or U1248 (N_1248,N_814,N_1076);
and U1249 (N_1249,N_687,N_943);
or U1250 (N_1250,N_969,N_1156);
nand U1251 (N_1251,N_1107,N_1125);
xor U1252 (N_1252,N_899,N_636);
xnor U1253 (N_1253,N_829,N_811);
and U1254 (N_1254,N_656,N_705);
nor U1255 (N_1255,N_1134,N_738);
or U1256 (N_1256,N_1087,N_630);
nor U1257 (N_1257,N_956,N_1180);
or U1258 (N_1258,N_1127,N_836);
and U1259 (N_1259,N_966,N_912);
xor U1260 (N_1260,N_870,N_860);
or U1261 (N_1261,N_1165,N_1068);
nor U1262 (N_1262,N_768,N_1028);
nand U1263 (N_1263,N_673,N_624);
nand U1264 (N_1264,N_680,N_670);
xor U1265 (N_1265,N_1178,N_792);
nand U1266 (N_1266,N_1016,N_1138);
or U1267 (N_1267,N_799,N_764);
nor U1268 (N_1268,N_803,N_1162);
and U1269 (N_1269,N_989,N_1116);
or U1270 (N_1270,N_626,N_1024);
xnor U1271 (N_1271,N_1158,N_917);
nand U1272 (N_1272,N_990,N_866);
or U1273 (N_1273,N_1000,N_628);
nor U1274 (N_1274,N_635,N_884);
xnor U1275 (N_1275,N_1189,N_801);
or U1276 (N_1276,N_751,N_900);
or U1277 (N_1277,N_776,N_1188);
nor U1278 (N_1278,N_907,N_683);
and U1279 (N_1279,N_1169,N_749);
and U1280 (N_1280,N_1190,N_995);
nor U1281 (N_1281,N_1039,N_1060);
nor U1282 (N_1282,N_753,N_824);
nor U1283 (N_1283,N_1163,N_775);
xor U1284 (N_1284,N_817,N_819);
and U1285 (N_1285,N_652,N_1003);
xnor U1286 (N_1286,N_1114,N_735);
nand U1287 (N_1287,N_1166,N_748);
and U1288 (N_1288,N_1095,N_978);
or U1289 (N_1289,N_773,N_769);
nand U1290 (N_1290,N_1143,N_1063);
nand U1291 (N_1291,N_1177,N_812);
nor U1292 (N_1292,N_1025,N_852);
and U1293 (N_1293,N_1054,N_717);
xnor U1294 (N_1294,N_794,N_826);
nor U1295 (N_1295,N_825,N_650);
nand U1296 (N_1296,N_784,N_1148);
nor U1297 (N_1297,N_758,N_611);
and U1298 (N_1298,N_828,N_1052);
or U1299 (N_1299,N_861,N_1109);
nand U1300 (N_1300,N_653,N_762);
or U1301 (N_1301,N_859,N_633);
nor U1302 (N_1302,N_918,N_1161);
nand U1303 (N_1303,N_1103,N_1193);
and U1304 (N_1304,N_718,N_704);
or U1305 (N_1305,N_700,N_920);
or U1306 (N_1306,N_963,N_1062);
and U1307 (N_1307,N_879,N_1194);
or U1308 (N_1308,N_1048,N_675);
nor U1309 (N_1309,N_690,N_668);
and U1310 (N_1310,N_925,N_935);
and U1311 (N_1311,N_994,N_600);
nand U1312 (N_1312,N_677,N_851);
and U1313 (N_1313,N_981,N_1132);
nor U1314 (N_1314,N_1196,N_1082);
nor U1315 (N_1315,N_713,N_921);
xnor U1316 (N_1316,N_897,N_983);
xor U1317 (N_1317,N_1045,N_1184);
xnor U1318 (N_1318,N_875,N_754);
and U1319 (N_1319,N_1035,N_982);
and U1320 (N_1320,N_728,N_845);
and U1321 (N_1321,N_746,N_678);
and U1322 (N_1322,N_744,N_810);
or U1323 (N_1323,N_785,N_601);
nand U1324 (N_1324,N_904,N_662);
or U1325 (N_1325,N_1179,N_664);
nor U1326 (N_1326,N_992,N_644);
or U1327 (N_1327,N_1101,N_1086);
and U1328 (N_1328,N_681,N_787);
nor U1329 (N_1329,N_657,N_973);
or U1330 (N_1330,N_1153,N_934);
nor U1331 (N_1331,N_610,N_1120);
or U1332 (N_1332,N_1155,N_679);
xnor U1333 (N_1333,N_790,N_820);
nor U1334 (N_1334,N_649,N_783);
nand U1335 (N_1335,N_752,N_706);
xnor U1336 (N_1336,N_620,N_1105);
or U1337 (N_1337,N_1089,N_1119);
nand U1338 (N_1338,N_685,N_763);
nor U1339 (N_1339,N_913,N_987);
nor U1340 (N_1340,N_1170,N_822);
nand U1341 (N_1341,N_716,N_813);
nand U1342 (N_1342,N_1160,N_686);
and U1343 (N_1343,N_1099,N_1151);
nor U1344 (N_1344,N_631,N_745);
xor U1345 (N_1345,N_1102,N_1118);
and U1346 (N_1346,N_938,N_780);
xnor U1347 (N_1347,N_1198,N_931);
xnor U1348 (N_1348,N_873,N_800);
nor U1349 (N_1349,N_1093,N_797);
xnor U1350 (N_1350,N_696,N_909);
nand U1351 (N_1351,N_1019,N_639);
xor U1352 (N_1352,N_1186,N_654);
nand U1353 (N_1353,N_789,N_609);
xnor U1354 (N_1354,N_888,N_726);
or U1355 (N_1355,N_878,N_739);
xnor U1356 (N_1356,N_872,N_1171);
and U1357 (N_1357,N_818,N_841);
or U1358 (N_1358,N_734,N_876);
or U1359 (N_1359,N_1149,N_694);
or U1360 (N_1360,N_1175,N_887);
and U1361 (N_1361,N_1191,N_902);
and U1362 (N_1362,N_965,N_1041);
xnor U1363 (N_1363,N_689,N_711);
xor U1364 (N_1364,N_737,N_1071);
and U1365 (N_1365,N_730,N_1167);
and U1366 (N_1366,N_857,N_809);
or U1367 (N_1367,N_940,N_805);
and U1368 (N_1368,N_1070,N_853);
nor U1369 (N_1369,N_1168,N_750);
or U1370 (N_1370,N_771,N_608);
xor U1371 (N_1371,N_1075,N_950);
or U1372 (N_1372,N_933,N_953);
nand U1373 (N_1373,N_779,N_756);
or U1374 (N_1374,N_1146,N_699);
or U1375 (N_1375,N_960,N_869);
nand U1376 (N_1376,N_1021,N_1085);
nor U1377 (N_1377,N_1139,N_910);
nand U1378 (N_1378,N_602,N_669);
or U1379 (N_1379,N_1164,N_757);
or U1380 (N_1380,N_937,N_942);
or U1381 (N_1381,N_660,N_1043);
nand U1382 (N_1382,N_702,N_890);
nand U1383 (N_1383,N_618,N_759);
or U1384 (N_1384,N_945,N_831);
nor U1385 (N_1385,N_619,N_676);
and U1386 (N_1386,N_772,N_1195);
or U1387 (N_1387,N_740,N_613);
nand U1388 (N_1388,N_947,N_793);
nor U1389 (N_1389,N_889,N_815);
or U1390 (N_1390,N_949,N_642);
nand U1391 (N_1391,N_774,N_911);
or U1392 (N_1392,N_895,N_951);
or U1393 (N_1393,N_906,N_614);
and U1394 (N_1394,N_1047,N_980);
and U1395 (N_1395,N_858,N_1074);
and U1396 (N_1396,N_1140,N_959);
nor U1397 (N_1397,N_682,N_1131);
nor U1398 (N_1398,N_691,N_1049);
or U1399 (N_1399,N_892,N_1181);
nor U1400 (N_1400,N_622,N_671);
and U1401 (N_1401,N_972,N_1057);
or U1402 (N_1402,N_1098,N_1097);
nor U1403 (N_1403,N_621,N_1044);
nor U1404 (N_1404,N_946,N_964);
nor U1405 (N_1405,N_1192,N_1199);
xor U1406 (N_1406,N_1108,N_1011);
nand U1407 (N_1407,N_928,N_1111);
and U1408 (N_1408,N_638,N_645);
xnor U1409 (N_1409,N_985,N_1152);
xor U1410 (N_1410,N_835,N_847);
xor U1411 (N_1411,N_840,N_939);
nand U1412 (N_1412,N_1065,N_1150);
or U1413 (N_1413,N_743,N_786);
or U1414 (N_1414,N_874,N_1172);
xor U1415 (N_1415,N_778,N_796);
or U1416 (N_1416,N_975,N_1042);
nand U1417 (N_1417,N_1067,N_952);
xnor U1418 (N_1418,N_1010,N_719);
xnor U1419 (N_1419,N_1126,N_695);
or U1420 (N_1420,N_893,N_954);
nand U1421 (N_1421,N_1036,N_967);
xor U1422 (N_1422,N_607,N_701);
or U1423 (N_1423,N_854,N_976);
and U1424 (N_1424,N_647,N_1104);
nor U1425 (N_1425,N_1113,N_862);
nand U1426 (N_1426,N_1176,N_1197);
and U1427 (N_1427,N_697,N_1112);
xnor U1428 (N_1428,N_837,N_993);
xnor U1429 (N_1429,N_722,N_604);
xor U1430 (N_1430,N_1015,N_807);
nand U1431 (N_1431,N_629,N_741);
or U1432 (N_1432,N_767,N_968);
nand U1433 (N_1433,N_1029,N_1023);
or U1434 (N_1434,N_1030,N_833);
xnor U1435 (N_1435,N_1159,N_666);
or U1436 (N_1436,N_634,N_707);
nor U1437 (N_1437,N_1032,N_1055);
and U1438 (N_1438,N_1083,N_1046);
xnor U1439 (N_1439,N_856,N_742);
xor U1440 (N_1440,N_839,N_908);
and U1441 (N_1441,N_844,N_684);
nand U1442 (N_1442,N_777,N_672);
or U1443 (N_1443,N_1144,N_944);
nand U1444 (N_1444,N_731,N_843);
or U1445 (N_1445,N_880,N_885);
nand U1446 (N_1446,N_1094,N_1096);
nor U1447 (N_1447,N_846,N_727);
or U1448 (N_1448,N_891,N_1091);
nor U1449 (N_1449,N_903,N_1123);
xnor U1450 (N_1450,N_1121,N_1013);
nor U1451 (N_1451,N_999,N_998);
xor U1452 (N_1452,N_606,N_929);
xor U1453 (N_1453,N_1173,N_930);
or U1454 (N_1454,N_867,N_1088);
nand U1455 (N_1455,N_617,N_1012);
xnor U1456 (N_1456,N_625,N_651);
nor U1457 (N_1457,N_864,N_834);
nand U1458 (N_1458,N_1005,N_1137);
nor U1459 (N_1459,N_766,N_709);
xnor U1460 (N_1460,N_1014,N_804);
nand U1461 (N_1461,N_848,N_1026);
nand U1462 (N_1462,N_855,N_901);
or U1463 (N_1463,N_1142,N_1034);
nor U1464 (N_1464,N_1037,N_643);
or U1465 (N_1465,N_1106,N_941);
nor U1466 (N_1466,N_732,N_603);
or U1467 (N_1467,N_1051,N_1059);
or U1468 (N_1468,N_1004,N_816);
xnor U1469 (N_1469,N_932,N_1056);
nor U1470 (N_1470,N_877,N_1130);
xor U1471 (N_1471,N_663,N_1133);
or U1472 (N_1472,N_1064,N_674);
nand U1473 (N_1473,N_881,N_1073);
nand U1474 (N_1474,N_640,N_896);
xnor U1475 (N_1475,N_1141,N_641);
nor U1476 (N_1476,N_692,N_849);
and U1477 (N_1477,N_795,N_883);
nand U1478 (N_1478,N_882,N_788);
and U1479 (N_1479,N_1078,N_703);
xnor U1480 (N_1480,N_1100,N_850);
nor U1481 (N_1481,N_1092,N_1061);
nor U1482 (N_1482,N_926,N_605);
or U1483 (N_1483,N_865,N_1136);
and U1484 (N_1484,N_791,N_996);
nor U1485 (N_1485,N_798,N_781);
or U1486 (N_1486,N_698,N_733);
nand U1487 (N_1487,N_1084,N_957);
nor U1488 (N_1488,N_661,N_693);
and U1489 (N_1489,N_827,N_974);
nor U1490 (N_1490,N_1122,N_1058);
nor U1491 (N_1491,N_988,N_924);
nand U1492 (N_1492,N_958,N_1050);
and U1493 (N_1493,N_627,N_655);
nor U1494 (N_1494,N_612,N_755);
or U1495 (N_1495,N_806,N_1117);
nor U1496 (N_1496,N_1040,N_1185);
or U1497 (N_1497,N_1154,N_1038);
xnor U1498 (N_1498,N_1069,N_708);
nand U1499 (N_1499,N_916,N_1018);
xnor U1500 (N_1500,N_689,N_897);
nor U1501 (N_1501,N_1013,N_648);
and U1502 (N_1502,N_790,N_939);
or U1503 (N_1503,N_846,N_806);
xor U1504 (N_1504,N_1090,N_620);
xnor U1505 (N_1505,N_919,N_860);
xnor U1506 (N_1506,N_1111,N_998);
xnor U1507 (N_1507,N_895,N_1081);
xnor U1508 (N_1508,N_753,N_1093);
and U1509 (N_1509,N_869,N_635);
xor U1510 (N_1510,N_733,N_700);
and U1511 (N_1511,N_753,N_686);
nand U1512 (N_1512,N_1156,N_1185);
and U1513 (N_1513,N_1029,N_1078);
nor U1514 (N_1514,N_673,N_945);
or U1515 (N_1515,N_864,N_1154);
xnor U1516 (N_1516,N_804,N_661);
and U1517 (N_1517,N_856,N_1155);
or U1518 (N_1518,N_741,N_882);
nand U1519 (N_1519,N_901,N_871);
and U1520 (N_1520,N_649,N_924);
or U1521 (N_1521,N_1051,N_893);
nand U1522 (N_1522,N_834,N_1093);
nor U1523 (N_1523,N_1006,N_903);
and U1524 (N_1524,N_874,N_984);
and U1525 (N_1525,N_830,N_981);
and U1526 (N_1526,N_844,N_1132);
and U1527 (N_1527,N_862,N_628);
nor U1528 (N_1528,N_732,N_656);
nand U1529 (N_1529,N_1108,N_662);
xnor U1530 (N_1530,N_1022,N_628);
and U1531 (N_1531,N_1132,N_1138);
or U1532 (N_1532,N_620,N_694);
and U1533 (N_1533,N_1016,N_730);
nand U1534 (N_1534,N_1113,N_675);
nand U1535 (N_1535,N_1197,N_1007);
xor U1536 (N_1536,N_1042,N_1098);
xor U1537 (N_1537,N_1162,N_660);
nor U1538 (N_1538,N_620,N_1101);
nand U1539 (N_1539,N_807,N_624);
xor U1540 (N_1540,N_998,N_991);
or U1541 (N_1541,N_633,N_806);
and U1542 (N_1542,N_714,N_884);
xnor U1543 (N_1543,N_912,N_729);
and U1544 (N_1544,N_674,N_917);
and U1545 (N_1545,N_794,N_1086);
and U1546 (N_1546,N_903,N_698);
nor U1547 (N_1547,N_642,N_1052);
or U1548 (N_1548,N_1164,N_958);
and U1549 (N_1549,N_1026,N_851);
nor U1550 (N_1550,N_1059,N_602);
nor U1551 (N_1551,N_833,N_809);
nand U1552 (N_1552,N_869,N_926);
or U1553 (N_1553,N_745,N_915);
xor U1554 (N_1554,N_806,N_748);
or U1555 (N_1555,N_990,N_930);
xnor U1556 (N_1556,N_781,N_1053);
or U1557 (N_1557,N_1125,N_919);
and U1558 (N_1558,N_955,N_707);
nand U1559 (N_1559,N_776,N_1183);
or U1560 (N_1560,N_788,N_1143);
or U1561 (N_1561,N_602,N_1009);
nand U1562 (N_1562,N_967,N_1142);
nand U1563 (N_1563,N_836,N_609);
xor U1564 (N_1564,N_1000,N_870);
nor U1565 (N_1565,N_800,N_1085);
nor U1566 (N_1566,N_831,N_1192);
and U1567 (N_1567,N_1066,N_797);
nand U1568 (N_1568,N_1172,N_652);
nor U1569 (N_1569,N_733,N_1029);
nor U1570 (N_1570,N_873,N_1101);
or U1571 (N_1571,N_1151,N_1013);
nand U1572 (N_1572,N_692,N_942);
or U1573 (N_1573,N_1049,N_662);
or U1574 (N_1574,N_600,N_743);
and U1575 (N_1575,N_706,N_1026);
or U1576 (N_1576,N_733,N_734);
and U1577 (N_1577,N_1137,N_893);
and U1578 (N_1578,N_675,N_1099);
xor U1579 (N_1579,N_1099,N_828);
xor U1580 (N_1580,N_958,N_618);
xnor U1581 (N_1581,N_921,N_1003);
or U1582 (N_1582,N_625,N_724);
and U1583 (N_1583,N_822,N_715);
xor U1584 (N_1584,N_603,N_1049);
and U1585 (N_1585,N_737,N_1160);
xor U1586 (N_1586,N_633,N_978);
nand U1587 (N_1587,N_906,N_644);
xnor U1588 (N_1588,N_1106,N_871);
and U1589 (N_1589,N_731,N_1128);
nor U1590 (N_1590,N_1132,N_1021);
or U1591 (N_1591,N_842,N_1188);
nor U1592 (N_1592,N_631,N_1175);
nand U1593 (N_1593,N_804,N_900);
nor U1594 (N_1594,N_906,N_700);
nor U1595 (N_1595,N_902,N_1077);
or U1596 (N_1596,N_610,N_1088);
nand U1597 (N_1597,N_873,N_625);
xor U1598 (N_1598,N_1119,N_860);
nand U1599 (N_1599,N_995,N_1049);
nand U1600 (N_1600,N_1068,N_861);
or U1601 (N_1601,N_766,N_1096);
and U1602 (N_1602,N_891,N_1056);
xor U1603 (N_1603,N_1148,N_622);
or U1604 (N_1604,N_1046,N_690);
nand U1605 (N_1605,N_869,N_610);
nor U1606 (N_1606,N_810,N_944);
xor U1607 (N_1607,N_877,N_790);
or U1608 (N_1608,N_1170,N_1075);
and U1609 (N_1609,N_922,N_891);
nand U1610 (N_1610,N_868,N_823);
nor U1611 (N_1611,N_948,N_730);
nor U1612 (N_1612,N_905,N_1001);
nor U1613 (N_1613,N_921,N_934);
xnor U1614 (N_1614,N_1108,N_840);
or U1615 (N_1615,N_886,N_940);
and U1616 (N_1616,N_1117,N_847);
nor U1617 (N_1617,N_819,N_1105);
nand U1618 (N_1618,N_973,N_782);
nor U1619 (N_1619,N_1039,N_1028);
nor U1620 (N_1620,N_764,N_767);
nor U1621 (N_1621,N_881,N_817);
nor U1622 (N_1622,N_744,N_865);
nand U1623 (N_1623,N_962,N_1087);
and U1624 (N_1624,N_923,N_798);
and U1625 (N_1625,N_1002,N_920);
xnor U1626 (N_1626,N_657,N_672);
nand U1627 (N_1627,N_953,N_1019);
nor U1628 (N_1628,N_863,N_971);
and U1629 (N_1629,N_1144,N_840);
or U1630 (N_1630,N_907,N_998);
xnor U1631 (N_1631,N_945,N_800);
xor U1632 (N_1632,N_1092,N_1012);
or U1633 (N_1633,N_1183,N_790);
nor U1634 (N_1634,N_901,N_1120);
and U1635 (N_1635,N_815,N_1076);
nor U1636 (N_1636,N_730,N_663);
nand U1637 (N_1637,N_1172,N_962);
nor U1638 (N_1638,N_885,N_1119);
xnor U1639 (N_1639,N_771,N_795);
and U1640 (N_1640,N_910,N_1181);
and U1641 (N_1641,N_1185,N_1139);
or U1642 (N_1642,N_829,N_868);
nand U1643 (N_1643,N_624,N_797);
nand U1644 (N_1644,N_1081,N_765);
xor U1645 (N_1645,N_693,N_1192);
or U1646 (N_1646,N_988,N_1000);
or U1647 (N_1647,N_736,N_1054);
nand U1648 (N_1648,N_799,N_632);
and U1649 (N_1649,N_607,N_611);
xor U1650 (N_1650,N_723,N_671);
xnor U1651 (N_1651,N_1105,N_668);
xnor U1652 (N_1652,N_670,N_959);
and U1653 (N_1653,N_686,N_1183);
xnor U1654 (N_1654,N_1109,N_1035);
nor U1655 (N_1655,N_841,N_756);
or U1656 (N_1656,N_984,N_1150);
nand U1657 (N_1657,N_643,N_802);
xnor U1658 (N_1658,N_887,N_1167);
nand U1659 (N_1659,N_912,N_1028);
nand U1660 (N_1660,N_667,N_940);
nand U1661 (N_1661,N_613,N_656);
xnor U1662 (N_1662,N_747,N_986);
nor U1663 (N_1663,N_920,N_613);
nand U1664 (N_1664,N_923,N_1170);
or U1665 (N_1665,N_983,N_903);
xor U1666 (N_1666,N_1102,N_776);
nor U1667 (N_1667,N_1198,N_1149);
xor U1668 (N_1668,N_1198,N_770);
nand U1669 (N_1669,N_1009,N_800);
nand U1670 (N_1670,N_990,N_634);
nor U1671 (N_1671,N_1133,N_653);
or U1672 (N_1672,N_611,N_755);
xnor U1673 (N_1673,N_649,N_1058);
nor U1674 (N_1674,N_1103,N_1134);
or U1675 (N_1675,N_755,N_930);
nand U1676 (N_1676,N_808,N_1070);
nor U1677 (N_1677,N_825,N_774);
nor U1678 (N_1678,N_997,N_653);
or U1679 (N_1679,N_1170,N_893);
nand U1680 (N_1680,N_648,N_687);
and U1681 (N_1681,N_809,N_759);
nor U1682 (N_1682,N_1052,N_716);
nand U1683 (N_1683,N_1037,N_1153);
or U1684 (N_1684,N_616,N_1068);
nand U1685 (N_1685,N_630,N_1176);
nor U1686 (N_1686,N_954,N_1175);
or U1687 (N_1687,N_1006,N_626);
xor U1688 (N_1688,N_1048,N_1174);
or U1689 (N_1689,N_618,N_1081);
nand U1690 (N_1690,N_953,N_975);
or U1691 (N_1691,N_647,N_1035);
nor U1692 (N_1692,N_817,N_803);
and U1693 (N_1693,N_929,N_1050);
or U1694 (N_1694,N_977,N_723);
nor U1695 (N_1695,N_1162,N_827);
nor U1696 (N_1696,N_817,N_845);
nor U1697 (N_1697,N_682,N_1038);
nor U1698 (N_1698,N_1162,N_1112);
nand U1699 (N_1699,N_1035,N_873);
xnor U1700 (N_1700,N_935,N_747);
or U1701 (N_1701,N_615,N_605);
and U1702 (N_1702,N_713,N_619);
nand U1703 (N_1703,N_1024,N_1064);
nor U1704 (N_1704,N_810,N_1084);
xnor U1705 (N_1705,N_715,N_684);
nand U1706 (N_1706,N_1152,N_1114);
xor U1707 (N_1707,N_885,N_1120);
xor U1708 (N_1708,N_636,N_916);
nand U1709 (N_1709,N_1184,N_838);
nor U1710 (N_1710,N_1119,N_873);
nor U1711 (N_1711,N_1148,N_963);
nand U1712 (N_1712,N_965,N_1191);
xnor U1713 (N_1713,N_997,N_687);
or U1714 (N_1714,N_670,N_790);
nor U1715 (N_1715,N_1181,N_719);
and U1716 (N_1716,N_1068,N_1161);
and U1717 (N_1717,N_862,N_881);
xor U1718 (N_1718,N_866,N_1129);
or U1719 (N_1719,N_657,N_756);
and U1720 (N_1720,N_730,N_761);
xor U1721 (N_1721,N_1110,N_1179);
nand U1722 (N_1722,N_628,N_844);
and U1723 (N_1723,N_1105,N_755);
and U1724 (N_1724,N_769,N_705);
or U1725 (N_1725,N_686,N_837);
xor U1726 (N_1726,N_727,N_929);
nand U1727 (N_1727,N_747,N_821);
and U1728 (N_1728,N_977,N_918);
nand U1729 (N_1729,N_1099,N_1165);
nor U1730 (N_1730,N_777,N_1019);
or U1731 (N_1731,N_1112,N_771);
nand U1732 (N_1732,N_838,N_753);
nand U1733 (N_1733,N_1013,N_1100);
or U1734 (N_1734,N_982,N_609);
or U1735 (N_1735,N_1110,N_802);
and U1736 (N_1736,N_931,N_997);
nand U1737 (N_1737,N_1169,N_877);
xnor U1738 (N_1738,N_1173,N_924);
nand U1739 (N_1739,N_906,N_608);
and U1740 (N_1740,N_1037,N_859);
and U1741 (N_1741,N_1080,N_603);
and U1742 (N_1742,N_740,N_1198);
nor U1743 (N_1743,N_748,N_953);
or U1744 (N_1744,N_700,N_1196);
xnor U1745 (N_1745,N_908,N_707);
and U1746 (N_1746,N_600,N_702);
and U1747 (N_1747,N_1023,N_923);
xnor U1748 (N_1748,N_806,N_1158);
nand U1749 (N_1749,N_614,N_853);
xor U1750 (N_1750,N_1080,N_776);
xnor U1751 (N_1751,N_804,N_1195);
or U1752 (N_1752,N_668,N_1120);
nand U1753 (N_1753,N_996,N_798);
or U1754 (N_1754,N_600,N_644);
or U1755 (N_1755,N_1072,N_892);
xnor U1756 (N_1756,N_765,N_857);
and U1757 (N_1757,N_646,N_1038);
or U1758 (N_1758,N_735,N_965);
or U1759 (N_1759,N_791,N_999);
and U1760 (N_1760,N_849,N_896);
nand U1761 (N_1761,N_931,N_875);
nand U1762 (N_1762,N_859,N_882);
or U1763 (N_1763,N_1169,N_1083);
xnor U1764 (N_1764,N_1176,N_880);
xor U1765 (N_1765,N_949,N_1181);
nand U1766 (N_1766,N_1082,N_802);
or U1767 (N_1767,N_639,N_1030);
xnor U1768 (N_1768,N_728,N_615);
and U1769 (N_1769,N_688,N_610);
nand U1770 (N_1770,N_804,N_825);
or U1771 (N_1771,N_820,N_809);
xor U1772 (N_1772,N_795,N_692);
xnor U1773 (N_1773,N_1133,N_886);
or U1774 (N_1774,N_985,N_789);
or U1775 (N_1775,N_1187,N_908);
nand U1776 (N_1776,N_609,N_1166);
xor U1777 (N_1777,N_980,N_604);
xnor U1778 (N_1778,N_1064,N_872);
or U1779 (N_1779,N_889,N_602);
nand U1780 (N_1780,N_1041,N_1056);
nor U1781 (N_1781,N_929,N_1080);
nand U1782 (N_1782,N_910,N_867);
nand U1783 (N_1783,N_1128,N_1191);
nor U1784 (N_1784,N_725,N_1173);
nand U1785 (N_1785,N_960,N_601);
and U1786 (N_1786,N_929,N_1130);
and U1787 (N_1787,N_683,N_825);
nand U1788 (N_1788,N_653,N_1165);
nand U1789 (N_1789,N_850,N_891);
xnor U1790 (N_1790,N_887,N_986);
and U1791 (N_1791,N_1101,N_954);
xor U1792 (N_1792,N_987,N_771);
xor U1793 (N_1793,N_1072,N_969);
nand U1794 (N_1794,N_922,N_1051);
nor U1795 (N_1795,N_766,N_1187);
nor U1796 (N_1796,N_1104,N_651);
and U1797 (N_1797,N_684,N_618);
and U1798 (N_1798,N_683,N_1003);
nor U1799 (N_1799,N_1126,N_998);
xor U1800 (N_1800,N_1450,N_1745);
nor U1801 (N_1801,N_1509,N_1412);
and U1802 (N_1802,N_1624,N_1219);
nor U1803 (N_1803,N_1573,N_1478);
nand U1804 (N_1804,N_1685,N_1783);
nand U1805 (N_1805,N_1331,N_1421);
and U1806 (N_1806,N_1488,N_1440);
nor U1807 (N_1807,N_1787,N_1645);
and U1808 (N_1808,N_1530,N_1283);
nor U1809 (N_1809,N_1311,N_1607);
xor U1810 (N_1810,N_1553,N_1286);
nand U1811 (N_1811,N_1308,N_1524);
or U1812 (N_1812,N_1718,N_1425);
and U1813 (N_1813,N_1340,N_1677);
and U1814 (N_1814,N_1538,N_1738);
or U1815 (N_1815,N_1442,N_1373);
and U1816 (N_1816,N_1426,N_1504);
and U1817 (N_1817,N_1248,N_1265);
xor U1818 (N_1818,N_1556,N_1616);
or U1819 (N_1819,N_1471,N_1346);
or U1820 (N_1820,N_1764,N_1643);
nand U1821 (N_1821,N_1254,N_1510);
xnor U1822 (N_1822,N_1379,N_1497);
nor U1823 (N_1823,N_1227,N_1695);
nand U1824 (N_1824,N_1518,N_1558);
or U1825 (N_1825,N_1415,N_1662);
and U1826 (N_1826,N_1794,N_1336);
nand U1827 (N_1827,N_1690,N_1266);
nor U1828 (N_1828,N_1231,N_1585);
and U1829 (N_1829,N_1343,N_1441);
or U1830 (N_1830,N_1743,N_1703);
and U1831 (N_1831,N_1572,N_1768);
nor U1832 (N_1832,N_1213,N_1411);
nor U1833 (N_1833,N_1674,N_1692);
or U1834 (N_1834,N_1390,N_1201);
and U1835 (N_1835,N_1544,N_1322);
or U1836 (N_1836,N_1375,N_1431);
nand U1837 (N_1837,N_1527,N_1420);
xnor U1838 (N_1838,N_1280,N_1586);
or U1839 (N_1839,N_1461,N_1615);
xnor U1840 (N_1840,N_1403,N_1563);
nor U1841 (N_1841,N_1514,N_1584);
nor U1842 (N_1842,N_1617,N_1378);
or U1843 (N_1843,N_1759,N_1376);
or U1844 (N_1844,N_1779,N_1430);
nand U1845 (N_1845,N_1487,N_1224);
nand U1846 (N_1846,N_1797,N_1484);
or U1847 (N_1847,N_1316,N_1795);
nand U1848 (N_1848,N_1720,N_1257);
xnor U1849 (N_1849,N_1503,N_1305);
and U1850 (N_1850,N_1385,N_1742);
xnor U1851 (N_1851,N_1771,N_1543);
xor U1852 (N_1852,N_1292,N_1715);
xnor U1853 (N_1853,N_1750,N_1708);
nor U1854 (N_1854,N_1408,N_1449);
nor U1855 (N_1855,N_1472,N_1479);
nor U1856 (N_1856,N_1749,N_1329);
nor U1857 (N_1857,N_1782,N_1583);
or U1858 (N_1858,N_1606,N_1595);
nand U1859 (N_1859,N_1374,N_1770);
nor U1860 (N_1860,N_1744,N_1491);
or U1861 (N_1861,N_1414,N_1529);
nand U1862 (N_1862,N_1383,N_1476);
and U1863 (N_1863,N_1398,N_1466);
or U1864 (N_1864,N_1396,N_1650);
nand U1865 (N_1865,N_1661,N_1774);
nor U1866 (N_1866,N_1549,N_1330);
or U1867 (N_1867,N_1763,N_1263);
and U1868 (N_1868,N_1796,N_1542);
or U1869 (N_1869,N_1608,N_1345);
or U1870 (N_1870,N_1299,N_1678);
nor U1871 (N_1871,N_1247,N_1788);
nor U1872 (N_1872,N_1511,N_1729);
or U1873 (N_1873,N_1657,N_1255);
nor U1874 (N_1874,N_1591,N_1459);
xor U1875 (N_1875,N_1666,N_1681);
and U1876 (N_1876,N_1437,N_1658);
nand U1877 (N_1877,N_1653,N_1339);
nor U1878 (N_1878,N_1647,N_1306);
and U1879 (N_1879,N_1222,N_1627);
xor U1880 (N_1880,N_1550,N_1539);
nor U1881 (N_1881,N_1724,N_1712);
nand U1882 (N_1882,N_1716,N_1238);
nand U1883 (N_1883,N_1673,N_1601);
and U1884 (N_1884,N_1559,N_1684);
and U1885 (N_1885,N_1633,N_1520);
and U1886 (N_1886,N_1364,N_1436);
nand U1887 (N_1887,N_1334,N_1335);
nor U1888 (N_1888,N_1675,N_1215);
or U1889 (N_1889,N_1792,N_1646);
nand U1890 (N_1890,N_1748,N_1506);
or U1891 (N_1891,N_1752,N_1648);
nand U1892 (N_1892,N_1216,N_1735);
xnor U1893 (N_1893,N_1337,N_1282);
and U1894 (N_1894,N_1571,N_1602);
nand U1895 (N_1895,N_1482,N_1686);
and U1896 (N_1896,N_1251,N_1264);
nand U1897 (N_1897,N_1279,N_1532);
or U1898 (N_1898,N_1576,N_1272);
nand U1899 (N_1899,N_1784,N_1734);
nor U1900 (N_1900,N_1649,N_1598);
xnor U1901 (N_1901,N_1456,N_1728);
and U1902 (N_1902,N_1697,N_1400);
xor U1903 (N_1903,N_1664,N_1758);
nor U1904 (N_1904,N_1221,N_1276);
nor U1905 (N_1905,N_1551,N_1704);
xor U1906 (N_1906,N_1409,N_1365);
xor U1907 (N_1907,N_1355,N_1707);
xor U1908 (N_1908,N_1386,N_1367);
xor U1909 (N_1909,N_1567,N_1470);
xnor U1910 (N_1910,N_1212,N_1424);
or U1911 (N_1911,N_1432,N_1244);
nand U1912 (N_1912,N_1302,N_1326);
nand U1913 (N_1913,N_1290,N_1687);
xor U1914 (N_1914,N_1610,N_1512);
and U1915 (N_1915,N_1274,N_1361);
or U1916 (N_1916,N_1402,N_1565);
nand U1917 (N_1917,N_1469,N_1651);
nor U1918 (N_1918,N_1297,N_1620);
and U1919 (N_1919,N_1528,N_1790);
nand U1920 (N_1920,N_1405,N_1701);
xor U1921 (N_1921,N_1575,N_1592);
xnor U1922 (N_1922,N_1756,N_1419);
nand U1923 (N_1923,N_1632,N_1760);
or U1924 (N_1924,N_1508,N_1249);
nor U1925 (N_1925,N_1635,N_1229);
and U1926 (N_1926,N_1714,N_1676);
nor U1927 (N_1927,N_1751,N_1753);
nand U1928 (N_1928,N_1682,N_1581);
or U1929 (N_1929,N_1536,N_1291);
and U1930 (N_1930,N_1372,N_1641);
nand U1931 (N_1931,N_1269,N_1435);
nand U1932 (N_1932,N_1545,N_1516);
and U1933 (N_1933,N_1665,N_1477);
xnor U1934 (N_1934,N_1799,N_1663);
xor U1935 (N_1935,N_1596,N_1303);
xor U1936 (N_1936,N_1287,N_1636);
or U1937 (N_1937,N_1533,N_1500);
nor U1938 (N_1938,N_1446,N_1644);
nor U1939 (N_1939,N_1320,N_1775);
or U1940 (N_1940,N_1786,N_1496);
xnor U1941 (N_1941,N_1341,N_1347);
and U1942 (N_1942,N_1368,N_1732);
or U1943 (N_1943,N_1258,N_1207);
nor U1944 (N_1944,N_1670,N_1259);
nor U1945 (N_1945,N_1566,N_1296);
and U1946 (N_1946,N_1318,N_1239);
or U1947 (N_1947,N_1310,N_1580);
and U1948 (N_1948,N_1468,N_1522);
xor U1949 (N_1949,N_1631,N_1353);
xor U1950 (N_1950,N_1726,N_1240);
nand U1951 (N_1951,N_1394,N_1531);
or U1952 (N_1952,N_1540,N_1217);
xnor U1953 (N_1953,N_1698,N_1593);
and U1954 (N_1954,N_1439,N_1767);
nand U1955 (N_1955,N_1669,N_1315);
and U1956 (N_1956,N_1659,N_1218);
and U1957 (N_1957,N_1301,N_1391);
or U1958 (N_1958,N_1246,N_1349);
or U1959 (N_1959,N_1600,N_1730);
and U1960 (N_1960,N_1594,N_1313);
or U1961 (N_1961,N_1214,N_1458);
or U1962 (N_1962,N_1689,N_1423);
xnor U1963 (N_1963,N_1589,N_1380);
and U1964 (N_1964,N_1381,N_1754);
or U1965 (N_1965,N_1691,N_1605);
and U1966 (N_1966,N_1481,N_1725);
nor U1967 (N_1967,N_1284,N_1569);
nor U1968 (N_1968,N_1384,N_1358);
and U1969 (N_1969,N_1772,N_1210);
nor U1970 (N_1970,N_1505,N_1554);
nand U1971 (N_1971,N_1234,N_1789);
nand U1972 (N_1972,N_1702,N_1314);
nand U1973 (N_1973,N_1696,N_1778);
and U1974 (N_1974,N_1711,N_1465);
or U1975 (N_1975,N_1434,N_1612);
nor U1976 (N_1976,N_1525,N_1289);
or U1977 (N_1977,N_1526,N_1236);
nor U1978 (N_1978,N_1727,N_1328);
nor U1979 (N_1979,N_1502,N_1304);
and U1980 (N_1980,N_1668,N_1388);
nand U1981 (N_1981,N_1588,N_1679);
and U1982 (N_1982,N_1416,N_1209);
nor U1983 (N_1983,N_1392,N_1521);
nor U1984 (N_1984,N_1312,N_1233);
and U1985 (N_1985,N_1639,N_1253);
nor U1986 (N_1986,N_1332,N_1327);
nor U1987 (N_1987,N_1579,N_1319);
or U1988 (N_1988,N_1428,N_1309);
nand U1989 (N_1989,N_1321,N_1307);
or U1990 (N_1990,N_1324,N_1443);
xnor U1991 (N_1991,N_1293,N_1363);
and U1992 (N_1992,N_1317,N_1204);
and U1993 (N_1993,N_1235,N_1245);
or U1994 (N_1994,N_1473,N_1746);
or U1995 (N_1995,N_1709,N_1781);
or U1996 (N_1996,N_1377,N_1582);
xnor U1997 (N_1997,N_1205,N_1277);
nand U1998 (N_1998,N_1741,N_1467);
xnor U1999 (N_1999,N_1495,N_1577);
or U2000 (N_2000,N_1688,N_1492);
nor U2001 (N_2001,N_1776,N_1348);
and U2002 (N_2002,N_1357,N_1252);
nor U2003 (N_2003,N_1773,N_1241);
xnor U2004 (N_2004,N_1404,N_1629);
nor U2005 (N_2005,N_1621,N_1694);
nand U2006 (N_2006,N_1541,N_1693);
or U2007 (N_2007,N_1275,N_1228);
and U2008 (N_2008,N_1777,N_1791);
and U2009 (N_2009,N_1519,N_1613);
and U2010 (N_2010,N_1226,N_1230);
or U2011 (N_2011,N_1483,N_1660);
and U2012 (N_2012,N_1557,N_1700);
or U2013 (N_2013,N_1603,N_1202);
nand U2014 (N_2014,N_1705,N_1338);
and U2015 (N_2015,N_1418,N_1298);
and U2016 (N_2016,N_1498,N_1351);
and U2017 (N_2017,N_1389,N_1407);
and U2018 (N_2018,N_1268,N_1737);
nor U2019 (N_2019,N_1628,N_1342);
nand U2020 (N_2020,N_1453,N_1270);
or U2021 (N_2021,N_1208,N_1387);
and U2022 (N_2022,N_1300,N_1578);
nand U2023 (N_2023,N_1634,N_1288);
xor U2024 (N_2024,N_1537,N_1517);
nor U2025 (N_2025,N_1507,N_1356);
xnor U2026 (N_2026,N_1486,N_1755);
xor U2027 (N_2027,N_1574,N_1623);
nand U2028 (N_2028,N_1640,N_1652);
xnor U2029 (N_2029,N_1344,N_1740);
and U2030 (N_2030,N_1560,N_1766);
or U2031 (N_2031,N_1395,N_1490);
xor U2032 (N_2032,N_1294,N_1671);
nor U2033 (N_2033,N_1417,N_1371);
nand U2034 (N_2034,N_1609,N_1422);
nor U2035 (N_2035,N_1278,N_1410);
xor U2036 (N_2036,N_1444,N_1590);
nor U2037 (N_2037,N_1447,N_1350);
and U2038 (N_2038,N_1562,N_1587);
and U2039 (N_2039,N_1489,N_1736);
nand U2040 (N_2040,N_1499,N_1451);
or U2041 (N_2041,N_1535,N_1798);
nor U2042 (N_2042,N_1366,N_1262);
nand U2043 (N_2043,N_1256,N_1599);
xnor U2044 (N_2044,N_1785,N_1780);
or U2045 (N_2045,N_1485,N_1382);
nor U2046 (N_2046,N_1765,N_1354);
or U2047 (N_2047,N_1757,N_1733);
nor U2048 (N_2048,N_1237,N_1513);
nor U2049 (N_2049,N_1655,N_1200);
nor U2050 (N_2050,N_1457,N_1547);
nor U2051 (N_2051,N_1243,N_1656);
nand U2052 (N_2052,N_1555,N_1534);
and U2053 (N_2053,N_1413,N_1427);
nand U2054 (N_2054,N_1464,N_1455);
and U2055 (N_2055,N_1762,N_1261);
and U2056 (N_2056,N_1433,N_1438);
nand U2057 (N_2057,N_1722,N_1448);
xor U2058 (N_2058,N_1564,N_1552);
xnor U2059 (N_2059,N_1225,N_1501);
xnor U2060 (N_2060,N_1672,N_1680);
and U2061 (N_2061,N_1642,N_1618);
nor U2062 (N_2062,N_1271,N_1360);
xnor U2063 (N_2063,N_1323,N_1761);
xor U2064 (N_2064,N_1739,N_1769);
or U2065 (N_2065,N_1359,N_1295);
and U2066 (N_2066,N_1713,N_1597);
xnor U2067 (N_2067,N_1706,N_1452);
or U2068 (N_2068,N_1223,N_1475);
or U2069 (N_2069,N_1242,N_1285);
and U2070 (N_2070,N_1710,N_1220);
nand U2071 (N_2071,N_1570,N_1494);
and U2072 (N_2072,N_1625,N_1654);
and U2073 (N_2073,N_1699,N_1614);
or U2074 (N_2074,N_1445,N_1747);
or U2075 (N_2075,N_1211,N_1463);
and U2076 (N_2076,N_1474,N_1250);
xor U2077 (N_2077,N_1622,N_1619);
xor U2078 (N_2078,N_1397,N_1515);
xor U2079 (N_2079,N_1546,N_1638);
nor U2080 (N_2080,N_1406,N_1429);
and U2081 (N_2081,N_1454,N_1370);
or U2082 (N_2082,N_1723,N_1203);
and U2083 (N_2083,N_1717,N_1281);
or U2084 (N_2084,N_1206,N_1523);
or U2085 (N_2085,N_1325,N_1462);
and U2086 (N_2086,N_1493,N_1626);
nand U2087 (N_2087,N_1568,N_1401);
nand U2088 (N_2088,N_1460,N_1630);
or U2089 (N_2089,N_1604,N_1273);
or U2090 (N_2090,N_1719,N_1637);
nand U2091 (N_2091,N_1561,N_1362);
nor U2092 (N_2092,N_1352,N_1793);
nor U2093 (N_2093,N_1369,N_1731);
nor U2094 (N_2094,N_1333,N_1611);
and U2095 (N_2095,N_1267,N_1667);
and U2096 (N_2096,N_1232,N_1480);
xnor U2097 (N_2097,N_1721,N_1683);
and U2098 (N_2098,N_1399,N_1393);
xnor U2099 (N_2099,N_1548,N_1260);
nor U2100 (N_2100,N_1585,N_1219);
or U2101 (N_2101,N_1633,N_1324);
and U2102 (N_2102,N_1203,N_1527);
and U2103 (N_2103,N_1771,N_1614);
and U2104 (N_2104,N_1750,N_1771);
or U2105 (N_2105,N_1209,N_1431);
nor U2106 (N_2106,N_1684,N_1427);
or U2107 (N_2107,N_1453,N_1385);
and U2108 (N_2108,N_1761,N_1751);
nand U2109 (N_2109,N_1365,N_1485);
nor U2110 (N_2110,N_1621,N_1291);
nand U2111 (N_2111,N_1776,N_1255);
or U2112 (N_2112,N_1726,N_1513);
nor U2113 (N_2113,N_1497,N_1756);
xor U2114 (N_2114,N_1673,N_1311);
xnor U2115 (N_2115,N_1523,N_1625);
and U2116 (N_2116,N_1321,N_1618);
xor U2117 (N_2117,N_1719,N_1262);
and U2118 (N_2118,N_1693,N_1616);
nor U2119 (N_2119,N_1765,N_1788);
or U2120 (N_2120,N_1581,N_1264);
and U2121 (N_2121,N_1714,N_1650);
nor U2122 (N_2122,N_1526,N_1568);
nand U2123 (N_2123,N_1386,N_1311);
xor U2124 (N_2124,N_1551,N_1339);
xor U2125 (N_2125,N_1703,N_1453);
nor U2126 (N_2126,N_1320,N_1481);
and U2127 (N_2127,N_1311,N_1557);
nand U2128 (N_2128,N_1333,N_1310);
and U2129 (N_2129,N_1373,N_1590);
nand U2130 (N_2130,N_1301,N_1346);
or U2131 (N_2131,N_1340,N_1374);
nor U2132 (N_2132,N_1794,N_1225);
nand U2133 (N_2133,N_1347,N_1473);
xor U2134 (N_2134,N_1691,N_1250);
or U2135 (N_2135,N_1400,N_1690);
and U2136 (N_2136,N_1709,N_1430);
xnor U2137 (N_2137,N_1733,N_1403);
xor U2138 (N_2138,N_1556,N_1672);
or U2139 (N_2139,N_1311,N_1586);
xnor U2140 (N_2140,N_1639,N_1303);
xnor U2141 (N_2141,N_1386,N_1696);
xnor U2142 (N_2142,N_1702,N_1794);
nor U2143 (N_2143,N_1313,N_1623);
and U2144 (N_2144,N_1764,N_1258);
and U2145 (N_2145,N_1597,N_1380);
and U2146 (N_2146,N_1586,N_1568);
xor U2147 (N_2147,N_1771,N_1747);
nor U2148 (N_2148,N_1729,N_1292);
nand U2149 (N_2149,N_1734,N_1659);
or U2150 (N_2150,N_1480,N_1642);
or U2151 (N_2151,N_1780,N_1537);
and U2152 (N_2152,N_1355,N_1646);
and U2153 (N_2153,N_1479,N_1513);
or U2154 (N_2154,N_1582,N_1311);
xnor U2155 (N_2155,N_1675,N_1723);
and U2156 (N_2156,N_1734,N_1458);
or U2157 (N_2157,N_1731,N_1616);
nor U2158 (N_2158,N_1561,N_1201);
or U2159 (N_2159,N_1427,N_1432);
or U2160 (N_2160,N_1698,N_1497);
nand U2161 (N_2161,N_1460,N_1361);
nand U2162 (N_2162,N_1708,N_1683);
nand U2163 (N_2163,N_1604,N_1333);
nand U2164 (N_2164,N_1574,N_1737);
nand U2165 (N_2165,N_1595,N_1359);
nor U2166 (N_2166,N_1355,N_1746);
nor U2167 (N_2167,N_1298,N_1619);
xor U2168 (N_2168,N_1454,N_1544);
nor U2169 (N_2169,N_1442,N_1584);
xnor U2170 (N_2170,N_1763,N_1549);
xor U2171 (N_2171,N_1320,N_1273);
nor U2172 (N_2172,N_1496,N_1758);
and U2173 (N_2173,N_1538,N_1415);
xnor U2174 (N_2174,N_1242,N_1600);
xor U2175 (N_2175,N_1746,N_1269);
nand U2176 (N_2176,N_1545,N_1471);
nand U2177 (N_2177,N_1457,N_1743);
and U2178 (N_2178,N_1496,N_1469);
nor U2179 (N_2179,N_1551,N_1281);
nand U2180 (N_2180,N_1371,N_1588);
xor U2181 (N_2181,N_1366,N_1333);
nand U2182 (N_2182,N_1486,N_1670);
or U2183 (N_2183,N_1512,N_1478);
or U2184 (N_2184,N_1557,N_1329);
or U2185 (N_2185,N_1523,N_1585);
nand U2186 (N_2186,N_1383,N_1242);
nor U2187 (N_2187,N_1368,N_1602);
or U2188 (N_2188,N_1780,N_1297);
and U2189 (N_2189,N_1281,N_1683);
nand U2190 (N_2190,N_1347,N_1572);
and U2191 (N_2191,N_1535,N_1793);
nand U2192 (N_2192,N_1615,N_1387);
xnor U2193 (N_2193,N_1516,N_1469);
or U2194 (N_2194,N_1762,N_1223);
and U2195 (N_2195,N_1438,N_1663);
or U2196 (N_2196,N_1216,N_1205);
nand U2197 (N_2197,N_1517,N_1662);
xor U2198 (N_2198,N_1223,N_1673);
nor U2199 (N_2199,N_1329,N_1735);
and U2200 (N_2200,N_1222,N_1528);
xnor U2201 (N_2201,N_1627,N_1593);
nor U2202 (N_2202,N_1713,N_1285);
nor U2203 (N_2203,N_1485,N_1575);
nor U2204 (N_2204,N_1489,N_1608);
nor U2205 (N_2205,N_1222,N_1337);
xor U2206 (N_2206,N_1276,N_1376);
or U2207 (N_2207,N_1711,N_1738);
nor U2208 (N_2208,N_1327,N_1748);
and U2209 (N_2209,N_1492,N_1476);
nand U2210 (N_2210,N_1588,N_1203);
xor U2211 (N_2211,N_1322,N_1641);
or U2212 (N_2212,N_1428,N_1266);
nor U2213 (N_2213,N_1640,N_1307);
and U2214 (N_2214,N_1508,N_1328);
nand U2215 (N_2215,N_1202,N_1460);
and U2216 (N_2216,N_1311,N_1652);
xnor U2217 (N_2217,N_1431,N_1467);
nand U2218 (N_2218,N_1652,N_1235);
and U2219 (N_2219,N_1327,N_1530);
or U2220 (N_2220,N_1597,N_1391);
or U2221 (N_2221,N_1766,N_1263);
nor U2222 (N_2222,N_1486,N_1282);
xnor U2223 (N_2223,N_1314,N_1609);
or U2224 (N_2224,N_1210,N_1319);
and U2225 (N_2225,N_1262,N_1798);
or U2226 (N_2226,N_1359,N_1426);
nor U2227 (N_2227,N_1464,N_1202);
nor U2228 (N_2228,N_1352,N_1716);
or U2229 (N_2229,N_1291,N_1694);
or U2230 (N_2230,N_1689,N_1366);
and U2231 (N_2231,N_1306,N_1464);
and U2232 (N_2232,N_1260,N_1565);
nand U2233 (N_2233,N_1398,N_1750);
xor U2234 (N_2234,N_1345,N_1595);
or U2235 (N_2235,N_1296,N_1441);
or U2236 (N_2236,N_1218,N_1668);
nor U2237 (N_2237,N_1579,N_1292);
nand U2238 (N_2238,N_1684,N_1570);
and U2239 (N_2239,N_1523,N_1708);
and U2240 (N_2240,N_1655,N_1244);
nand U2241 (N_2241,N_1764,N_1742);
and U2242 (N_2242,N_1642,N_1399);
xnor U2243 (N_2243,N_1300,N_1773);
nor U2244 (N_2244,N_1276,N_1520);
or U2245 (N_2245,N_1661,N_1330);
xnor U2246 (N_2246,N_1618,N_1334);
or U2247 (N_2247,N_1726,N_1598);
nand U2248 (N_2248,N_1480,N_1707);
and U2249 (N_2249,N_1361,N_1202);
nand U2250 (N_2250,N_1750,N_1719);
xor U2251 (N_2251,N_1541,N_1456);
xnor U2252 (N_2252,N_1749,N_1508);
or U2253 (N_2253,N_1450,N_1430);
nand U2254 (N_2254,N_1324,N_1418);
or U2255 (N_2255,N_1262,N_1579);
xnor U2256 (N_2256,N_1306,N_1388);
and U2257 (N_2257,N_1711,N_1222);
or U2258 (N_2258,N_1552,N_1665);
xor U2259 (N_2259,N_1736,N_1591);
xnor U2260 (N_2260,N_1694,N_1778);
nand U2261 (N_2261,N_1502,N_1630);
nand U2262 (N_2262,N_1278,N_1220);
nor U2263 (N_2263,N_1325,N_1735);
nand U2264 (N_2264,N_1752,N_1345);
or U2265 (N_2265,N_1291,N_1440);
nor U2266 (N_2266,N_1495,N_1218);
and U2267 (N_2267,N_1603,N_1297);
nand U2268 (N_2268,N_1230,N_1583);
xnor U2269 (N_2269,N_1784,N_1571);
or U2270 (N_2270,N_1688,N_1392);
or U2271 (N_2271,N_1639,N_1418);
nor U2272 (N_2272,N_1780,N_1464);
or U2273 (N_2273,N_1759,N_1545);
nor U2274 (N_2274,N_1280,N_1438);
or U2275 (N_2275,N_1458,N_1276);
nor U2276 (N_2276,N_1726,N_1395);
xor U2277 (N_2277,N_1320,N_1497);
nand U2278 (N_2278,N_1557,N_1756);
nand U2279 (N_2279,N_1724,N_1497);
xor U2280 (N_2280,N_1773,N_1205);
and U2281 (N_2281,N_1614,N_1510);
and U2282 (N_2282,N_1437,N_1349);
xor U2283 (N_2283,N_1357,N_1479);
nor U2284 (N_2284,N_1471,N_1235);
xor U2285 (N_2285,N_1751,N_1460);
and U2286 (N_2286,N_1758,N_1349);
nor U2287 (N_2287,N_1771,N_1572);
and U2288 (N_2288,N_1520,N_1267);
nand U2289 (N_2289,N_1327,N_1745);
nand U2290 (N_2290,N_1724,N_1744);
or U2291 (N_2291,N_1310,N_1719);
nand U2292 (N_2292,N_1581,N_1665);
xor U2293 (N_2293,N_1536,N_1279);
xnor U2294 (N_2294,N_1212,N_1590);
or U2295 (N_2295,N_1731,N_1212);
and U2296 (N_2296,N_1560,N_1215);
nor U2297 (N_2297,N_1224,N_1514);
or U2298 (N_2298,N_1560,N_1613);
nand U2299 (N_2299,N_1423,N_1579);
nand U2300 (N_2300,N_1732,N_1620);
nand U2301 (N_2301,N_1780,N_1798);
nor U2302 (N_2302,N_1247,N_1745);
nor U2303 (N_2303,N_1598,N_1343);
nand U2304 (N_2304,N_1589,N_1214);
nand U2305 (N_2305,N_1441,N_1780);
nand U2306 (N_2306,N_1365,N_1270);
nand U2307 (N_2307,N_1277,N_1774);
nor U2308 (N_2308,N_1524,N_1372);
and U2309 (N_2309,N_1222,N_1629);
nand U2310 (N_2310,N_1518,N_1541);
and U2311 (N_2311,N_1781,N_1296);
nor U2312 (N_2312,N_1252,N_1290);
and U2313 (N_2313,N_1474,N_1204);
and U2314 (N_2314,N_1299,N_1358);
xnor U2315 (N_2315,N_1234,N_1467);
or U2316 (N_2316,N_1665,N_1213);
or U2317 (N_2317,N_1305,N_1720);
nand U2318 (N_2318,N_1269,N_1259);
xnor U2319 (N_2319,N_1746,N_1216);
nand U2320 (N_2320,N_1445,N_1268);
and U2321 (N_2321,N_1534,N_1208);
nand U2322 (N_2322,N_1532,N_1472);
or U2323 (N_2323,N_1551,N_1662);
nand U2324 (N_2324,N_1322,N_1333);
nand U2325 (N_2325,N_1246,N_1589);
xnor U2326 (N_2326,N_1213,N_1538);
nand U2327 (N_2327,N_1675,N_1745);
nor U2328 (N_2328,N_1457,N_1363);
xor U2329 (N_2329,N_1567,N_1541);
xor U2330 (N_2330,N_1496,N_1390);
nand U2331 (N_2331,N_1472,N_1585);
nand U2332 (N_2332,N_1621,N_1368);
or U2333 (N_2333,N_1211,N_1497);
nand U2334 (N_2334,N_1761,N_1677);
or U2335 (N_2335,N_1528,N_1741);
nor U2336 (N_2336,N_1435,N_1367);
or U2337 (N_2337,N_1711,N_1243);
and U2338 (N_2338,N_1411,N_1225);
xor U2339 (N_2339,N_1355,N_1798);
xnor U2340 (N_2340,N_1229,N_1724);
xnor U2341 (N_2341,N_1280,N_1454);
xnor U2342 (N_2342,N_1303,N_1755);
nand U2343 (N_2343,N_1466,N_1747);
or U2344 (N_2344,N_1246,N_1649);
and U2345 (N_2345,N_1473,N_1715);
nand U2346 (N_2346,N_1310,N_1709);
and U2347 (N_2347,N_1340,N_1604);
or U2348 (N_2348,N_1311,N_1203);
or U2349 (N_2349,N_1332,N_1275);
nand U2350 (N_2350,N_1392,N_1592);
or U2351 (N_2351,N_1734,N_1481);
and U2352 (N_2352,N_1726,N_1521);
or U2353 (N_2353,N_1346,N_1418);
and U2354 (N_2354,N_1580,N_1207);
or U2355 (N_2355,N_1318,N_1578);
nor U2356 (N_2356,N_1359,N_1208);
nand U2357 (N_2357,N_1555,N_1658);
nand U2358 (N_2358,N_1660,N_1340);
and U2359 (N_2359,N_1587,N_1393);
or U2360 (N_2360,N_1604,N_1352);
nand U2361 (N_2361,N_1469,N_1591);
or U2362 (N_2362,N_1561,N_1568);
nor U2363 (N_2363,N_1216,N_1245);
and U2364 (N_2364,N_1310,N_1200);
nor U2365 (N_2365,N_1602,N_1682);
or U2366 (N_2366,N_1558,N_1630);
or U2367 (N_2367,N_1290,N_1645);
nand U2368 (N_2368,N_1474,N_1559);
nor U2369 (N_2369,N_1322,N_1565);
and U2370 (N_2370,N_1311,N_1626);
nor U2371 (N_2371,N_1461,N_1632);
nand U2372 (N_2372,N_1454,N_1243);
nand U2373 (N_2373,N_1640,N_1231);
nor U2374 (N_2374,N_1627,N_1499);
xnor U2375 (N_2375,N_1735,N_1421);
and U2376 (N_2376,N_1560,N_1534);
xor U2377 (N_2377,N_1467,N_1643);
nand U2378 (N_2378,N_1475,N_1525);
or U2379 (N_2379,N_1683,N_1264);
nand U2380 (N_2380,N_1365,N_1323);
and U2381 (N_2381,N_1752,N_1456);
nor U2382 (N_2382,N_1504,N_1410);
nand U2383 (N_2383,N_1667,N_1290);
nor U2384 (N_2384,N_1707,N_1278);
xnor U2385 (N_2385,N_1373,N_1216);
xor U2386 (N_2386,N_1213,N_1544);
nor U2387 (N_2387,N_1385,N_1780);
nor U2388 (N_2388,N_1431,N_1756);
and U2389 (N_2389,N_1255,N_1466);
xor U2390 (N_2390,N_1539,N_1720);
nand U2391 (N_2391,N_1633,N_1524);
and U2392 (N_2392,N_1741,N_1322);
or U2393 (N_2393,N_1543,N_1706);
nor U2394 (N_2394,N_1666,N_1537);
nor U2395 (N_2395,N_1213,N_1777);
and U2396 (N_2396,N_1215,N_1616);
nor U2397 (N_2397,N_1515,N_1503);
xnor U2398 (N_2398,N_1680,N_1760);
xnor U2399 (N_2399,N_1366,N_1723);
xnor U2400 (N_2400,N_2039,N_2067);
xnor U2401 (N_2401,N_1976,N_2382);
or U2402 (N_2402,N_1963,N_1883);
xor U2403 (N_2403,N_2189,N_2178);
or U2404 (N_2404,N_2234,N_2045);
xor U2405 (N_2405,N_2001,N_1887);
or U2406 (N_2406,N_2163,N_2381);
nand U2407 (N_2407,N_1861,N_2250);
and U2408 (N_2408,N_1930,N_2175);
nor U2409 (N_2409,N_2048,N_2364);
nand U2410 (N_2410,N_1873,N_2092);
nand U2411 (N_2411,N_1928,N_1856);
xnor U2412 (N_2412,N_2065,N_1837);
nand U2413 (N_2413,N_1903,N_2113);
or U2414 (N_2414,N_1966,N_2357);
nor U2415 (N_2415,N_2077,N_1944);
and U2416 (N_2416,N_1961,N_1847);
and U2417 (N_2417,N_2371,N_2119);
nand U2418 (N_2418,N_2379,N_2015);
and U2419 (N_2419,N_2011,N_1989);
and U2420 (N_2420,N_1886,N_1901);
or U2421 (N_2421,N_2235,N_1945);
or U2422 (N_2422,N_2316,N_2262);
xnor U2423 (N_2423,N_1821,N_2298);
or U2424 (N_2424,N_2319,N_2172);
nor U2425 (N_2425,N_2056,N_2356);
or U2426 (N_2426,N_1958,N_2278);
or U2427 (N_2427,N_2004,N_2302);
nor U2428 (N_2428,N_2117,N_2006);
or U2429 (N_2429,N_2360,N_1932);
xnor U2430 (N_2430,N_2130,N_2259);
and U2431 (N_2431,N_2207,N_2080);
xnor U2432 (N_2432,N_2297,N_1996);
xnor U2433 (N_2433,N_1864,N_1857);
nor U2434 (N_2434,N_2229,N_1809);
or U2435 (N_2435,N_1891,N_2343);
nor U2436 (N_2436,N_1827,N_2396);
nor U2437 (N_2437,N_2210,N_2332);
nand U2438 (N_2438,N_2188,N_1898);
and U2439 (N_2439,N_2196,N_2224);
or U2440 (N_2440,N_1906,N_2191);
nand U2441 (N_2441,N_2152,N_2208);
nor U2442 (N_2442,N_2069,N_2078);
nand U2443 (N_2443,N_2283,N_2288);
or U2444 (N_2444,N_1855,N_2099);
nand U2445 (N_2445,N_2068,N_1853);
nand U2446 (N_2446,N_2009,N_2263);
nor U2447 (N_2447,N_1962,N_1943);
and U2448 (N_2448,N_2213,N_1851);
nor U2449 (N_2449,N_1889,N_2007);
and U2450 (N_2450,N_2076,N_2243);
nand U2451 (N_2451,N_1916,N_2249);
xor U2452 (N_2452,N_2087,N_2136);
nor U2453 (N_2453,N_2184,N_2135);
and U2454 (N_2454,N_1813,N_1979);
xor U2455 (N_2455,N_2383,N_2033);
or U2456 (N_2456,N_2399,N_2385);
nand U2457 (N_2457,N_1900,N_1994);
and U2458 (N_2458,N_2174,N_2304);
or U2459 (N_2459,N_1841,N_2389);
and U2460 (N_2460,N_2301,N_1879);
xnor U2461 (N_2461,N_1805,N_2269);
and U2462 (N_2462,N_2390,N_2395);
and U2463 (N_2463,N_2293,N_2139);
or U2464 (N_2464,N_2326,N_2226);
nor U2465 (N_2465,N_1806,N_2317);
and U2466 (N_2466,N_2374,N_1843);
nand U2467 (N_2467,N_1955,N_2367);
nor U2468 (N_2468,N_2232,N_1824);
xor U2469 (N_2469,N_2325,N_1890);
nand U2470 (N_2470,N_2378,N_2031);
nor U2471 (N_2471,N_2314,N_1967);
nor U2472 (N_2472,N_2377,N_2195);
nand U2473 (N_2473,N_2336,N_2159);
nand U2474 (N_2474,N_2217,N_2013);
xnor U2475 (N_2475,N_2372,N_2164);
xor U2476 (N_2476,N_2362,N_2233);
xnor U2477 (N_2477,N_2331,N_1876);
nand U2478 (N_2478,N_2018,N_2355);
xor U2479 (N_2479,N_1998,N_1836);
or U2480 (N_2480,N_1986,N_1811);
or U2481 (N_2481,N_1862,N_2179);
nor U2482 (N_2482,N_1965,N_2176);
xor U2483 (N_2483,N_2157,N_2248);
nor U2484 (N_2484,N_2185,N_2275);
and U2485 (N_2485,N_1865,N_1907);
or U2486 (N_2486,N_1812,N_2260);
nand U2487 (N_2487,N_2141,N_1984);
or U2488 (N_2488,N_2267,N_2097);
nor U2489 (N_2489,N_1867,N_2026);
xor U2490 (N_2490,N_1893,N_2061);
nor U2491 (N_2491,N_1973,N_2064);
nand U2492 (N_2492,N_2155,N_1803);
or U2493 (N_2493,N_2255,N_2323);
xnor U2494 (N_2494,N_2270,N_1840);
xor U2495 (N_2495,N_2041,N_2131);
or U2496 (N_2496,N_1937,N_2165);
nor U2497 (N_2497,N_1938,N_2287);
xor U2498 (N_2498,N_2016,N_2114);
and U2499 (N_2499,N_1957,N_2116);
nor U2500 (N_2500,N_1810,N_2388);
nand U2501 (N_2501,N_1991,N_2230);
and U2502 (N_2502,N_2201,N_2118);
nor U2503 (N_2503,N_1920,N_2149);
and U2504 (N_2504,N_2375,N_2036);
and U2505 (N_2505,N_2008,N_2303);
xnor U2506 (N_2506,N_2205,N_2052);
or U2507 (N_2507,N_2012,N_1845);
and U2508 (N_2508,N_1968,N_2063);
and U2509 (N_2509,N_2066,N_2245);
and U2510 (N_2510,N_1804,N_2140);
and U2511 (N_2511,N_2392,N_2327);
or U2512 (N_2512,N_2274,N_2158);
xor U2513 (N_2513,N_2346,N_2352);
xnor U2514 (N_2514,N_2111,N_2032);
or U2515 (N_2515,N_1871,N_2264);
nand U2516 (N_2516,N_1858,N_1995);
nand U2517 (N_2517,N_2014,N_2137);
nand U2518 (N_2518,N_2047,N_2095);
nand U2519 (N_2519,N_1972,N_2121);
xnor U2520 (N_2520,N_1970,N_2242);
and U2521 (N_2521,N_2342,N_2156);
or U2522 (N_2522,N_2206,N_2285);
or U2523 (N_2523,N_1919,N_2289);
nor U2524 (N_2524,N_1951,N_1825);
and U2525 (N_2525,N_1981,N_2177);
or U2526 (N_2526,N_1926,N_2348);
and U2527 (N_2527,N_2295,N_1915);
nand U2528 (N_2528,N_2101,N_1828);
and U2529 (N_2529,N_2394,N_2199);
and U2530 (N_2530,N_1917,N_1880);
or U2531 (N_2531,N_1854,N_2286);
xor U2532 (N_2532,N_2086,N_2102);
nor U2533 (N_2533,N_2082,N_2306);
or U2534 (N_2534,N_2161,N_2143);
or U2535 (N_2535,N_2202,N_2105);
and U2536 (N_2536,N_2349,N_2236);
and U2537 (N_2537,N_1829,N_1849);
nor U2538 (N_2538,N_1801,N_1808);
nand U2539 (N_2539,N_2110,N_2350);
nor U2540 (N_2540,N_2222,N_1800);
nor U2541 (N_2541,N_2180,N_2334);
or U2542 (N_2542,N_2329,N_2171);
nor U2543 (N_2543,N_2017,N_1936);
or U2544 (N_2544,N_2160,N_2313);
and U2545 (N_2545,N_1913,N_1911);
or U2546 (N_2546,N_2055,N_2219);
nor U2547 (N_2547,N_2088,N_2238);
and U2548 (N_2548,N_2376,N_2025);
or U2549 (N_2549,N_1934,N_2128);
or U2550 (N_2550,N_2221,N_2090);
or U2551 (N_2551,N_2062,N_2335);
or U2552 (N_2552,N_1977,N_2386);
nor U2553 (N_2553,N_2261,N_1933);
nand U2554 (N_2554,N_1842,N_1908);
nor U2555 (N_2555,N_2265,N_1838);
nand U2556 (N_2556,N_2005,N_2125);
and U2557 (N_2557,N_1969,N_2333);
or U2558 (N_2558,N_2028,N_2091);
nor U2559 (N_2559,N_1953,N_1910);
nand U2560 (N_2560,N_1868,N_2251);
nor U2561 (N_2561,N_1832,N_1863);
xor U2562 (N_2562,N_2257,N_1807);
nand U2563 (N_2563,N_2312,N_1954);
nand U2564 (N_2564,N_1940,N_2256);
and U2565 (N_2565,N_1814,N_1947);
nor U2566 (N_2566,N_2190,N_2145);
and U2567 (N_2567,N_1848,N_2059);
nand U2568 (N_2568,N_2182,N_2281);
and U2569 (N_2569,N_2366,N_1939);
nor U2570 (N_2570,N_2038,N_2134);
or U2571 (N_2571,N_2307,N_2123);
or U2572 (N_2572,N_1921,N_2387);
and U2573 (N_2573,N_2290,N_1831);
and U2574 (N_2574,N_2054,N_2299);
nand U2575 (N_2575,N_1833,N_2146);
nand U2576 (N_2576,N_2070,N_1844);
nor U2577 (N_2577,N_1822,N_2104);
or U2578 (N_2578,N_2339,N_2084);
xor U2579 (N_2579,N_1877,N_2049);
or U2580 (N_2580,N_1830,N_2169);
xnor U2581 (N_2581,N_1978,N_2183);
and U2582 (N_2582,N_1892,N_1860);
and U2583 (N_2583,N_2057,N_2079);
nor U2584 (N_2584,N_2073,N_2223);
nor U2585 (N_2585,N_2363,N_1941);
xnor U2586 (N_2586,N_2291,N_2050);
nor U2587 (N_2587,N_1881,N_2280);
nor U2588 (N_2588,N_2369,N_2240);
nand U2589 (N_2589,N_1895,N_2107);
and U2590 (N_2590,N_2397,N_2034);
nand U2591 (N_2591,N_1905,N_2225);
xnor U2592 (N_2592,N_2072,N_2126);
nand U2593 (N_2593,N_1950,N_1914);
nor U2594 (N_2594,N_2258,N_2344);
xnor U2595 (N_2595,N_1990,N_2368);
nor U2596 (N_2596,N_2096,N_2365);
nand U2597 (N_2597,N_2153,N_2268);
and U2598 (N_2598,N_2060,N_2138);
nand U2599 (N_2599,N_2109,N_2305);
nand U2600 (N_2600,N_2043,N_2115);
and U2601 (N_2601,N_1959,N_1818);
xnor U2602 (N_2602,N_2373,N_2051);
xor U2603 (N_2603,N_2168,N_2181);
nand U2604 (N_2604,N_2030,N_1997);
nor U2605 (N_2605,N_2003,N_1894);
nand U2606 (N_2606,N_2296,N_2231);
nor U2607 (N_2607,N_1902,N_2330);
or U2608 (N_2608,N_2020,N_1866);
nand U2609 (N_2609,N_1948,N_2227);
or U2610 (N_2610,N_2284,N_2186);
and U2611 (N_2611,N_2127,N_2380);
or U2612 (N_2612,N_2211,N_2276);
nor U2613 (N_2613,N_2112,N_2083);
nor U2614 (N_2614,N_1802,N_2204);
nor U2615 (N_2615,N_2273,N_1918);
and U2616 (N_2616,N_2228,N_1850);
or U2617 (N_2617,N_1852,N_1885);
and U2618 (N_2618,N_1999,N_2282);
or U2619 (N_2619,N_1909,N_2324);
xor U2620 (N_2620,N_2359,N_2279);
or U2621 (N_2621,N_2010,N_2272);
nand U2622 (N_2622,N_2021,N_1935);
and U2623 (N_2623,N_1927,N_2247);
nand U2624 (N_2624,N_1923,N_1992);
xnor U2625 (N_2625,N_1983,N_1875);
nand U2626 (N_2626,N_1980,N_2340);
xnor U2627 (N_2627,N_1859,N_2133);
xor U2628 (N_2628,N_2300,N_1987);
nand U2629 (N_2629,N_2192,N_2193);
or U2630 (N_2630,N_2085,N_1956);
nand U2631 (N_2631,N_1869,N_2214);
or U2632 (N_2632,N_1896,N_1819);
and U2633 (N_2633,N_1839,N_1912);
and U2634 (N_2634,N_1846,N_2308);
or U2635 (N_2635,N_2081,N_2022);
or U2636 (N_2636,N_2142,N_2321);
and U2637 (N_2637,N_2311,N_2074);
or U2638 (N_2638,N_2294,N_2198);
nand U2639 (N_2639,N_2029,N_2239);
nor U2640 (N_2640,N_2002,N_1929);
and U2641 (N_2641,N_2241,N_1975);
or U2642 (N_2642,N_2370,N_1971);
nand U2643 (N_2643,N_2212,N_2218);
nor U2644 (N_2644,N_2194,N_2393);
and U2645 (N_2645,N_2197,N_2108);
or U2646 (N_2646,N_1942,N_2132);
xnor U2647 (N_2647,N_2338,N_2252);
or U2648 (N_2648,N_1816,N_1931);
nand U2649 (N_2649,N_2266,N_1988);
xor U2650 (N_2650,N_2094,N_2322);
nand U2651 (N_2651,N_2147,N_2209);
and U2652 (N_2652,N_1897,N_2046);
xor U2653 (N_2653,N_1974,N_2220);
and U2654 (N_2654,N_2042,N_1826);
nor U2655 (N_2655,N_2358,N_2098);
nand U2656 (N_2656,N_2315,N_1964);
xor U2657 (N_2657,N_1960,N_2044);
and U2658 (N_2658,N_2309,N_2071);
xor U2659 (N_2659,N_2341,N_2122);
nand U2660 (N_2660,N_2148,N_2027);
or U2661 (N_2661,N_2246,N_1874);
xnor U2662 (N_2662,N_1835,N_2353);
nand U2663 (N_2663,N_2391,N_1882);
xnor U2664 (N_2664,N_2173,N_2024);
nand U2665 (N_2665,N_1823,N_1888);
or U2666 (N_2666,N_2384,N_1872);
and U2667 (N_2667,N_2253,N_2216);
nor U2668 (N_2668,N_1993,N_1952);
or U2669 (N_2669,N_1878,N_2347);
nor U2670 (N_2670,N_2129,N_2244);
nand U2671 (N_2671,N_2093,N_1834);
or U2672 (N_2672,N_2040,N_2058);
and U2673 (N_2673,N_2154,N_2167);
nor U2674 (N_2674,N_2328,N_2203);
and U2675 (N_2675,N_1946,N_2000);
nand U2676 (N_2676,N_2354,N_2053);
and U2677 (N_2677,N_2170,N_2124);
nor U2678 (N_2678,N_2277,N_2292);
nand U2679 (N_2679,N_1925,N_2037);
nor U2680 (N_2680,N_2351,N_2310);
and U2681 (N_2681,N_2023,N_2345);
or U2682 (N_2682,N_2151,N_2075);
or U2683 (N_2683,N_2120,N_2271);
and U2684 (N_2684,N_2200,N_1820);
xor U2685 (N_2685,N_2019,N_2144);
and U2686 (N_2686,N_1815,N_2398);
nor U2687 (N_2687,N_2150,N_1985);
and U2688 (N_2688,N_2337,N_2254);
nand U2689 (N_2689,N_1924,N_1904);
nor U2690 (N_2690,N_2166,N_2100);
and U2691 (N_2691,N_2187,N_1982);
nand U2692 (N_2692,N_1899,N_1817);
or U2693 (N_2693,N_2089,N_2320);
and U2694 (N_2694,N_2215,N_1922);
or U2695 (N_2695,N_2035,N_1884);
nor U2696 (N_2696,N_1949,N_2237);
and U2697 (N_2697,N_2162,N_2103);
nor U2698 (N_2698,N_2106,N_2318);
nand U2699 (N_2699,N_2361,N_1870);
nor U2700 (N_2700,N_2013,N_2282);
and U2701 (N_2701,N_1925,N_2318);
nand U2702 (N_2702,N_2330,N_2043);
nor U2703 (N_2703,N_2186,N_2058);
nand U2704 (N_2704,N_2305,N_2381);
or U2705 (N_2705,N_1985,N_1818);
or U2706 (N_2706,N_2068,N_2296);
nor U2707 (N_2707,N_1954,N_2273);
nand U2708 (N_2708,N_2325,N_2310);
or U2709 (N_2709,N_1935,N_1913);
nand U2710 (N_2710,N_2309,N_2101);
and U2711 (N_2711,N_2004,N_2122);
nor U2712 (N_2712,N_2194,N_2230);
nor U2713 (N_2713,N_2391,N_1859);
nor U2714 (N_2714,N_2026,N_2270);
or U2715 (N_2715,N_1894,N_2115);
nor U2716 (N_2716,N_1825,N_1905);
xnor U2717 (N_2717,N_2194,N_2337);
or U2718 (N_2718,N_2397,N_2292);
and U2719 (N_2719,N_2370,N_2335);
xor U2720 (N_2720,N_1931,N_2191);
nand U2721 (N_2721,N_1836,N_2346);
and U2722 (N_2722,N_2375,N_2091);
nor U2723 (N_2723,N_2073,N_2310);
and U2724 (N_2724,N_2144,N_1877);
xor U2725 (N_2725,N_2273,N_1907);
nand U2726 (N_2726,N_2080,N_1975);
nor U2727 (N_2727,N_1966,N_2013);
nor U2728 (N_2728,N_1916,N_2080);
xnor U2729 (N_2729,N_2383,N_1846);
and U2730 (N_2730,N_2111,N_2142);
nor U2731 (N_2731,N_1967,N_2041);
nor U2732 (N_2732,N_1858,N_1930);
nor U2733 (N_2733,N_1867,N_2105);
nor U2734 (N_2734,N_2387,N_2059);
xor U2735 (N_2735,N_2169,N_2229);
or U2736 (N_2736,N_2125,N_1981);
xnor U2737 (N_2737,N_2006,N_1846);
or U2738 (N_2738,N_1972,N_2103);
and U2739 (N_2739,N_2244,N_2006);
nand U2740 (N_2740,N_2337,N_1884);
xor U2741 (N_2741,N_2111,N_2267);
or U2742 (N_2742,N_2310,N_2033);
and U2743 (N_2743,N_1996,N_2128);
nand U2744 (N_2744,N_2173,N_2232);
nor U2745 (N_2745,N_1974,N_2071);
xor U2746 (N_2746,N_2380,N_1938);
or U2747 (N_2747,N_1906,N_2392);
nor U2748 (N_2748,N_1884,N_1833);
xnor U2749 (N_2749,N_2274,N_2348);
or U2750 (N_2750,N_2086,N_2045);
or U2751 (N_2751,N_2398,N_1883);
nand U2752 (N_2752,N_1881,N_2187);
and U2753 (N_2753,N_2157,N_2358);
and U2754 (N_2754,N_2151,N_2212);
nand U2755 (N_2755,N_1824,N_2393);
xnor U2756 (N_2756,N_2072,N_2191);
nand U2757 (N_2757,N_2237,N_2367);
or U2758 (N_2758,N_2399,N_2264);
nand U2759 (N_2759,N_2352,N_2355);
nand U2760 (N_2760,N_1885,N_1928);
nand U2761 (N_2761,N_2031,N_2222);
nand U2762 (N_2762,N_1974,N_1817);
and U2763 (N_2763,N_1945,N_1841);
and U2764 (N_2764,N_2034,N_2217);
and U2765 (N_2765,N_1936,N_2107);
xor U2766 (N_2766,N_2027,N_2292);
xor U2767 (N_2767,N_2351,N_2033);
or U2768 (N_2768,N_2138,N_2390);
nand U2769 (N_2769,N_1886,N_1872);
or U2770 (N_2770,N_2341,N_2010);
or U2771 (N_2771,N_2310,N_2335);
nor U2772 (N_2772,N_2108,N_2383);
or U2773 (N_2773,N_1852,N_2190);
xor U2774 (N_2774,N_2333,N_1893);
nor U2775 (N_2775,N_2321,N_2354);
or U2776 (N_2776,N_2220,N_2048);
and U2777 (N_2777,N_2128,N_2300);
nand U2778 (N_2778,N_2048,N_1873);
xnor U2779 (N_2779,N_1895,N_1891);
or U2780 (N_2780,N_2096,N_2017);
nor U2781 (N_2781,N_1826,N_2073);
and U2782 (N_2782,N_1950,N_2099);
or U2783 (N_2783,N_2222,N_1927);
or U2784 (N_2784,N_2113,N_2033);
nand U2785 (N_2785,N_2202,N_2072);
nand U2786 (N_2786,N_2057,N_1835);
xnor U2787 (N_2787,N_1901,N_1996);
nor U2788 (N_2788,N_2230,N_2008);
nor U2789 (N_2789,N_2356,N_2041);
or U2790 (N_2790,N_2230,N_2104);
and U2791 (N_2791,N_1920,N_2013);
and U2792 (N_2792,N_1822,N_2189);
nand U2793 (N_2793,N_1913,N_2292);
xor U2794 (N_2794,N_2145,N_2057);
and U2795 (N_2795,N_1919,N_2339);
nand U2796 (N_2796,N_2346,N_2359);
nor U2797 (N_2797,N_2393,N_2095);
or U2798 (N_2798,N_2077,N_1935);
or U2799 (N_2799,N_2230,N_2395);
xnor U2800 (N_2800,N_1889,N_2314);
nor U2801 (N_2801,N_1825,N_1999);
and U2802 (N_2802,N_2254,N_2342);
xnor U2803 (N_2803,N_2247,N_2220);
or U2804 (N_2804,N_1847,N_2271);
nand U2805 (N_2805,N_2177,N_1914);
xnor U2806 (N_2806,N_2173,N_1956);
or U2807 (N_2807,N_2029,N_1858);
nor U2808 (N_2808,N_2117,N_2211);
and U2809 (N_2809,N_1952,N_2390);
or U2810 (N_2810,N_2271,N_2280);
nand U2811 (N_2811,N_1835,N_1889);
or U2812 (N_2812,N_2104,N_2091);
xor U2813 (N_2813,N_2329,N_1845);
nor U2814 (N_2814,N_1954,N_1810);
and U2815 (N_2815,N_2064,N_2253);
and U2816 (N_2816,N_2048,N_1825);
xor U2817 (N_2817,N_2327,N_2345);
or U2818 (N_2818,N_2380,N_2025);
or U2819 (N_2819,N_2148,N_2025);
and U2820 (N_2820,N_1983,N_2339);
nand U2821 (N_2821,N_2261,N_1800);
and U2822 (N_2822,N_2005,N_2344);
xnor U2823 (N_2823,N_1951,N_2018);
xor U2824 (N_2824,N_1995,N_1804);
nor U2825 (N_2825,N_2196,N_2156);
or U2826 (N_2826,N_2306,N_1843);
xnor U2827 (N_2827,N_1932,N_1958);
or U2828 (N_2828,N_2061,N_1975);
nand U2829 (N_2829,N_2024,N_2074);
nand U2830 (N_2830,N_2185,N_1913);
nor U2831 (N_2831,N_2167,N_2149);
and U2832 (N_2832,N_1818,N_1920);
xor U2833 (N_2833,N_2332,N_2001);
and U2834 (N_2834,N_1899,N_2298);
and U2835 (N_2835,N_2186,N_2372);
nand U2836 (N_2836,N_2391,N_2172);
nand U2837 (N_2837,N_2384,N_2030);
or U2838 (N_2838,N_2354,N_2331);
and U2839 (N_2839,N_2319,N_2141);
and U2840 (N_2840,N_2185,N_2258);
nand U2841 (N_2841,N_2324,N_2010);
and U2842 (N_2842,N_2296,N_2236);
nor U2843 (N_2843,N_2277,N_1810);
nand U2844 (N_2844,N_2213,N_1971);
and U2845 (N_2845,N_1806,N_2281);
and U2846 (N_2846,N_1861,N_1911);
and U2847 (N_2847,N_2115,N_1878);
xor U2848 (N_2848,N_2382,N_2064);
nor U2849 (N_2849,N_1847,N_2362);
xor U2850 (N_2850,N_1832,N_1928);
or U2851 (N_2851,N_1938,N_1887);
nor U2852 (N_2852,N_2343,N_2213);
nand U2853 (N_2853,N_2101,N_2212);
and U2854 (N_2854,N_2117,N_2237);
nor U2855 (N_2855,N_2263,N_2223);
or U2856 (N_2856,N_1886,N_1957);
xnor U2857 (N_2857,N_1892,N_2055);
nor U2858 (N_2858,N_2325,N_2395);
or U2859 (N_2859,N_1933,N_2390);
or U2860 (N_2860,N_2332,N_2023);
or U2861 (N_2861,N_2221,N_1854);
and U2862 (N_2862,N_1907,N_1987);
or U2863 (N_2863,N_2037,N_2245);
and U2864 (N_2864,N_2025,N_2242);
xnor U2865 (N_2865,N_2034,N_1917);
nor U2866 (N_2866,N_2105,N_2267);
xor U2867 (N_2867,N_1860,N_2004);
nor U2868 (N_2868,N_1879,N_1967);
or U2869 (N_2869,N_2014,N_2034);
nand U2870 (N_2870,N_2266,N_2260);
nand U2871 (N_2871,N_1998,N_1960);
or U2872 (N_2872,N_1833,N_2326);
xor U2873 (N_2873,N_2156,N_2316);
and U2874 (N_2874,N_2076,N_2325);
nor U2875 (N_2875,N_2011,N_2015);
nand U2876 (N_2876,N_2097,N_2298);
and U2877 (N_2877,N_2060,N_2252);
xor U2878 (N_2878,N_2005,N_2095);
and U2879 (N_2879,N_2355,N_2327);
and U2880 (N_2880,N_2213,N_2250);
and U2881 (N_2881,N_2235,N_2102);
nor U2882 (N_2882,N_1836,N_2377);
xnor U2883 (N_2883,N_2336,N_2379);
xor U2884 (N_2884,N_2298,N_2062);
nor U2885 (N_2885,N_2270,N_1835);
nor U2886 (N_2886,N_1909,N_2109);
xor U2887 (N_2887,N_2077,N_1918);
and U2888 (N_2888,N_1859,N_2075);
or U2889 (N_2889,N_1956,N_2382);
and U2890 (N_2890,N_2111,N_1954);
or U2891 (N_2891,N_2308,N_2211);
xnor U2892 (N_2892,N_2374,N_2324);
or U2893 (N_2893,N_1905,N_2101);
and U2894 (N_2894,N_1948,N_2367);
or U2895 (N_2895,N_2385,N_1840);
or U2896 (N_2896,N_1900,N_2306);
and U2897 (N_2897,N_2387,N_2255);
nor U2898 (N_2898,N_2135,N_2310);
or U2899 (N_2899,N_2000,N_1978);
nand U2900 (N_2900,N_2291,N_2259);
nand U2901 (N_2901,N_2336,N_2267);
xnor U2902 (N_2902,N_2054,N_1959);
nor U2903 (N_2903,N_2397,N_1829);
nor U2904 (N_2904,N_1819,N_1978);
nor U2905 (N_2905,N_2388,N_2277);
and U2906 (N_2906,N_1992,N_1995);
or U2907 (N_2907,N_2108,N_1899);
and U2908 (N_2908,N_2227,N_2267);
xnor U2909 (N_2909,N_2336,N_2148);
and U2910 (N_2910,N_2004,N_1959);
xor U2911 (N_2911,N_2287,N_2248);
nand U2912 (N_2912,N_2049,N_1986);
nand U2913 (N_2913,N_2093,N_2318);
nor U2914 (N_2914,N_2300,N_2181);
xnor U2915 (N_2915,N_1827,N_1951);
nand U2916 (N_2916,N_1829,N_2166);
nor U2917 (N_2917,N_2116,N_2353);
nand U2918 (N_2918,N_2192,N_1941);
xnor U2919 (N_2919,N_1912,N_1814);
and U2920 (N_2920,N_2033,N_1854);
nand U2921 (N_2921,N_1833,N_2341);
or U2922 (N_2922,N_2380,N_2245);
or U2923 (N_2923,N_2238,N_2370);
or U2924 (N_2924,N_2135,N_1987);
nor U2925 (N_2925,N_1857,N_2274);
xnor U2926 (N_2926,N_2159,N_2187);
xor U2927 (N_2927,N_1983,N_2381);
xnor U2928 (N_2928,N_2266,N_2216);
nor U2929 (N_2929,N_2115,N_2250);
nor U2930 (N_2930,N_1985,N_2189);
nand U2931 (N_2931,N_1869,N_2038);
and U2932 (N_2932,N_2158,N_2102);
and U2933 (N_2933,N_2394,N_1831);
xnor U2934 (N_2934,N_2023,N_2014);
nand U2935 (N_2935,N_1840,N_1884);
nor U2936 (N_2936,N_2015,N_2308);
nor U2937 (N_2937,N_2290,N_1890);
xnor U2938 (N_2938,N_2216,N_2094);
or U2939 (N_2939,N_1987,N_1952);
nor U2940 (N_2940,N_2054,N_2292);
xnor U2941 (N_2941,N_1980,N_2054);
nand U2942 (N_2942,N_2370,N_2119);
nand U2943 (N_2943,N_1819,N_2070);
or U2944 (N_2944,N_2065,N_1802);
nor U2945 (N_2945,N_2336,N_1967);
nand U2946 (N_2946,N_2198,N_2344);
xor U2947 (N_2947,N_2068,N_2303);
or U2948 (N_2948,N_2069,N_2292);
and U2949 (N_2949,N_1907,N_1844);
xor U2950 (N_2950,N_2190,N_2308);
or U2951 (N_2951,N_2235,N_2390);
and U2952 (N_2952,N_2285,N_1872);
xnor U2953 (N_2953,N_1806,N_2002);
and U2954 (N_2954,N_2332,N_1806);
and U2955 (N_2955,N_2217,N_2128);
and U2956 (N_2956,N_2274,N_2157);
nand U2957 (N_2957,N_1972,N_2188);
nand U2958 (N_2958,N_1896,N_2266);
or U2959 (N_2959,N_2044,N_2240);
nor U2960 (N_2960,N_2365,N_1812);
nand U2961 (N_2961,N_1867,N_2094);
nor U2962 (N_2962,N_2204,N_2262);
nor U2963 (N_2963,N_2240,N_2138);
nor U2964 (N_2964,N_2147,N_2073);
nand U2965 (N_2965,N_1827,N_1958);
and U2966 (N_2966,N_2289,N_2112);
nand U2967 (N_2967,N_2284,N_1838);
xnor U2968 (N_2968,N_1933,N_1903);
xnor U2969 (N_2969,N_2009,N_2170);
nand U2970 (N_2970,N_1954,N_1964);
and U2971 (N_2971,N_1949,N_2029);
or U2972 (N_2972,N_2355,N_2287);
or U2973 (N_2973,N_2256,N_2055);
xnor U2974 (N_2974,N_2310,N_1850);
xor U2975 (N_2975,N_2261,N_2174);
and U2976 (N_2976,N_1996,N_2140);
and U2977 (N_2977,N_1975,N_1890);
or U2978 (N_2978,N_2087,N_1893);
and U2979 (N_2979,N_2117,N_2202);
and U2980 (N_2980,N_1918,N_2050);
and U2981 (N_2981,N_1945,N_2136);
or U2982 (N_2982,N_1861,N_1848);
nor U2983 (N_2983,N_2243,N_2148);
or U2984 (N_2984,N_1986,N_2130);
and U2985 (N_2985,N_1815,N_2346);
nand U2986 (N_2986,N_1962,N_2087);
and U2987 (N_2987,N_2334,N_2086);
xnor U2988 (N_2988,N_1841,N_2197);
xor U2989 (N_2989,N_2091,N_2382);
or U2990 (N_2990,N_2169,N_2289);
or U2991 (N_2991,N_2195,N_1915);
nor U2992 (N_2992,N_2278,N_1911);
nand U2993 (N_2993,N_2382,N_1850);
nor U2994 (N_2994,N_2234,N_1833);
xnor U2995 (N_2995,N_1826,N_2137);
or U2996 (N_2996,N_2237,N_1933);
or U2997 (N_2997,N_1856,N_1880);
xnor U2998 (N_2998,N_2067,N_1969);
and U2999 (N_2999,N_1957,N_2342);
or UO_0 (O_0,N_2604,N_2674);
nor UO_1 (O_1,N_2440,N_2574);
nand UO_2 (O_2,N_2417,N_2893);
nand UO_3 (O_3,N_2435,N_2805);
or UO_4 (O_4,N_2712,N_2739);
nand UO_5 (O_5,N_2447,N_2534);
nand UO_6 (O_6,N_2575,N_2837);
nand UO_7 (O_7,N_2754,N_2445);
and UO_8 (O_8,N_2949,N_2617);
or UO_9 (O_9,N_2791,N_2726);
nand UO_10 (O_10,N_2539,N_2661);
or UO_11 (O_11,N_2662,N_2564);
nand UO_12 (O_12,N_2875,N_2593);
or UO_13 (O_13,N_2678,N_2597);
or UO_14 (O_14,N_2522,N_2693);
and UO_15 (O_15,N_2563,N_2886);
and UO_16 (O_16,N_2671,N_2813);
or UO_17 (O_17,N_2732,N_2869);
nor UO_18 (O_18,N_2470,N_2959);
and UO_19 (O_19,N_2681,N_2498);
nor UO_20 (O_20,N_2481,N_2997);
or UO_21 (O_21,N_2737,N_2629);
nand UO_22 (O_22,N_2586,N_2816);
nand UO_23 (O_23,N_2588,N_2882);
and UO_24 (O_24,N_2938,N_2720);
nand UO_25 (O_25,N_2550,N_2967);
xnor UO_26 (O_26,N_2434,N_2957);
xnor UO_27 (O_27,N_2413,N_2790);
xnor UO_28 (O_28,N_2426,N_2632);
and UO_29 (O_29,N_2489,N_2424);
and UO_30 (O_30,N_2985,N_2702);
nor UO_31 (O_31,N_2803,N_2628);
or UO_32 (O_32,N_2659,N_2746);
nor UO_33 (O_33,N_2826,N_2404);
or UO_34 (O_34,N_2589,N_2897);
xnor UO_35 (O_35,N_2703,N_2598);
nand UO_36 (O_36,N_2821,N_2640);
xnor UO_37 (O_37,N_2443,N_2694);
or UO_38 (O_38,N_2902,N_2636);
and UO_39 (O_39,N_2735,N_2706);
xnor UO_40 (O_40,N_2545,N_2861);
nor UO_41 (O_41,N_2623,N_2918);
nand UO_42 (O_42,N_2559,N_2438);
nor UO_43 (O_43,N_2976,N_2465);
and UO_44 (O_44,N_2998,N_2543);
and UO_45 (O_45,N_2439,N_2412);
xnor UO_46 (O_46,N_2649,N_2848);
and UO_47 (O_47,N_2572,N_2827);
nor UO_48 (O_48,N_2457,N_2936);
xor UO_49 (O_49,N_2762,N_2890);
nand UO_50 (O_50,N_2418,N_2609);
and UO_51 (O_51,N_2981,N_2843);
or UO_52 (O_52,N_2740,N_2437);
and UO_53 (O_53,N_2458,N_2874);
xor UO_54 (O_54,N_2829,N_2601);
nand UO_55 (O_55,N_2819,N_2983);
nor UO_56 (O_56,N_2904,N_2809);
xnor UO_57 (O_57,N_2855,N_2556);
and UO_58 (O_58,N_2555,N_2419);
or UO_59 (O_59,N_2715,N_2579);
and UO_60 (O_60,N_2653,N_2991);
or UO_61 (O_61,N_2505,N_2774);
nor UO_62 (O_62,N_2898,N_2728);
nor UO_63 (O_63,N_2734,N_2517);
nor UO_64 (O_64,N_2776,N_2511);
or UO_65 (O_65,N_2951,N_2646);
or UO_66 (O_66,N_2449,N_2885);
or UO_67 (O_67,N_2525,N_2554);
nor UO_68 (O_68,N_2596,N_2789);
and UO_69 (O_69,N_2411,N_2941);
or UO_70 (O_70,N_2521,N_2558);
and UO_71 (O_71,N_2849,N_2704);
nor UO_72 (O_72,N_2839,N_2570);
nor UO_73 (O_73,N_2451,N_2838);
nand UO_74 (O_74,N_2479,N_2812);
and UO_75 (O_75,N_2752,N_2710);
nand UO_76 (O_76,N_2787,N_2456);
and UO_77 (O_77,N_2663,N_2937);
and UO_78 (O_78,N_2782,N_2468);
and UO_79 (O_79,N_2568,N_2698);
nor UO_80 (O_80,N_2431,N_2648);
xor UO_81 (O_81,N_2892,N_2778);
or UO_82 (O_82,N_2889,N_2476);
nand UO_83 (O_83,N_2770,N_2988);
nor UO_84 (O_84,N_2668,N_2795);
and UO_85 (O_85,N_2781,N_2406);
and UO_86 (O_86,N_2566,N_2922);
or UO_87 (O_87,N_2786,N_2851);
nor UO_88 (O_88,N_2565,N_2773);
or UO_89 (O_89,N_2705,N_2722);
and UO_90 (O_90,N_2911,N_2974);
and UO_91 (O_91,N_2863,N_2968);
nor UO_92 (O_92,N_2929,N_2784);
or UO_93 (O_93,N_2666,N_2856);
nand UO_94 (O_94,N_2761,N_2669);
nand UO_95 (O_95,N_2714,N_2901);
and UO_96 (O_96,N_2637,N_2792);
nor UO_97 (O_97,N_2804,N_2680);
nand UO_98 (O_98,N_2908,N_2796);
and UO_99 (O_99,N_2535,N_2883);
xnor UO_100 (O_100,N_2763,N_2613);
nand UO_101 (O_101,N_2711,N_2950);
or UO_102 (O_102,N_2721,N_2724);
or UO_103 (O_103,N_2682,N_2753);
nor UO_104 (O_104,N_2416,N_2815);
nor UO_105 (O_105,N_2667,N_2527);
xor UO_106 (O_106,N_2928,N_2896);
or UO_107 (O_107,N_2859,N_2820);
xor UO_108 (O_108,N_2584,N_2618);
and UO_109 (O_109,N_2621,N_2408);
nand UO_110 (O_110,N_2616,N_2614);
and UO_111 (O_111,N_2987,N_2460);
or UO_112 (O_112,N_2871,N_2800);
or UO_113 (O_113,N_2425,N_2836);
xor UO_114 (O_114,N_2642,N_2644);
nor UO_115 (O_115,N_2639,N_2708);
xor UO_116 (O_116,N_2731,N_2462);
xor UO_117 (O_117,N_2488,N_2910);
nand UO_118 (O_118,N_2510,N_2873);
nand UO_119 (O_119,N_2946,N_2444);
nand UO_120 (O_120,N_2611,N_2594);
and UO_121 (O_121,N_2528,N_2422);
or UO_122 (O_122,N_2493,N_2920);
nor UO_123 (O_123,N_2657,N_2733);
and UO_124 (O_124,N_2743,N_2992);
nand UO_125 (O_125,N_2749,N_2979);
nor UO_126 (O_126,N_2982,N_2699);
nand UO_127 (O_127,N_2587,N_2852);
xor UO_128 (O_128,N_2676,N_2603);
and UO_129 (O_129,N_2467,N_2478);
or UO_130 (O_130,N_2758,N_2626);
nor UO_131 (O_131,N_2673,N_2725);
and UO_132 (O_132,N_2599,N_2672);
nand UO_133 (O_133,N_2552,N_2971);
and UO_134 (O_134,N_2832,N_2688);
nand UO_135 (O_135,N_2878,N_2780);
and UO_136 (O_136,N_2783,N_2622);
xnor UO_137 (O_137,N_2477,N_2788);
or UO_138 (O_138,N_2798,N_2544);
nand UO_139 (O_139,N_2634,N_2464);
nor UO_140 (O_140,N_2802,N_2532);
or UO_141 (O_141,N_2475,N_2958);
and UO_142 (O_142,N_2400,N_2686);
nand UO_143 (O_143,N_2664,N_2943);
or UO_144 (O_144,N_2605,N_2866);
and UO_145 (O_145,N_2915,N_2582);
nand UO_146 (O_146,N_2945,N_2631);
and UO_147 (O_147,N_2825,N_2940);
xor UO_148 (O_148,N_2963,N_2756);
nor UO_149 (O_149,N_2606,N_2751);
nand UO_150 (O_150,N_2947,N_2665);
nand UO_151 (O_151,N_2683,N_2560);
nor UO_152 (O_152,N_2421,N_2516);
nor UO_153 (O_153,N_2923,N_2953);
nand UO_154 (O_154,N_2502,N_2692);
nor UO_155 (O_155,N_2850,N_2524);
nand UO_156 (O_156,N_2842,N_2442);
nand UO_157 (O_157,N_2580,N_2409);
nor UO_158 (O_158,N_2497,N_2670);
xnor UO_159 (O_159,N_2491,N_2925);
or UO_160 (O_160,N_2537,N_2463);
and UO_161 (O_161,N_2459,N_2677);
xnor UO_162 (O_162,N_2729,N_2551);
or UO_163 (O_163,N_2500,N_2769);
nand UO_164 (O_164,N_2707,N_2541);
xor UO_165 (O_165,N_2771,N_2581);
and UO_166 (O_166,N_2494,N_2441);
or UO_167 (O_167,N_2870,N_2748);
xnor UO_168 (O_168,N_2980,N_2961);
xor UO_169 (O_169,N_2402,N_2994);
and UO_170 (O_170,N_2834,N_2831);
or UO_171 (O_171,N_2755,N_2960);
nor UO_172 (O_172,N_2984,N_2742);
xor UO_173 (O_173,N_2697,N_2509);
nand UO_174 (O_174,N_2407,N_2853);
xnor UO_175 (O_175,N_2415,N_2955);
or UO_176 (O_176,N_2767,N_2512);
nand UO_177 (O_177,N_2466,N_2410);
or UO_178 (O_178,N_2430,N_2638);
xnor UO_179 (O_179,N_2585,N_2548);
nor UO_180 (O_180,N_2956,N_2935);
and UO_181 (O_181,N_2818,N_2801);
and UO_182 (O_182,N_2557,N_2429);
and UO_183 (O_183,N_2654,N_2841);
or UO_184 (O_184,N_2917,N_2571);
nand UO_185 (O_185,N_2766,N_2808);
xor UO_186 (O_186,N_2954,N_2546);
nor UO_187 (O_187,N_2716,N_2595);
xnor UO_188 (O_188,N_2966,N_2881);
nor UO_189 (O_189,N_2436,N_2822);
nand UO_190 (O_190,N_2695,N_2660);
nor UO_191 (O_191,N_2578,N_2899);
and UO_192 (O_192,N_2480,N_2891);
or UO_193 (O_193,N_2738,N_2765);
nand UO_194 (O_194,N_2995,N_2496);
or UO_195 (O_195,N_2487,N_2608);
and UO_196 (O_196,N_2583,N_2520);
xor UO_197 (O_197,N_2931,N_2860);
xnor UO_198 (O_198,N_2887,N_2448);
xor UO_199 (O_199,N_2972,N_2569);
nor UO_200 (O_200,N_2858,N_2744);
xnor UO_201 (O_201,N_2750,N_2562);
xor UO_202 (O_202,N_2741,N_2864);
or UO_203 (O_203,N_2542,N_2455);
nor UO_204 (O_204,N_2894,N_2531);
nor UO_205 (O_205,N_2857,N_2635);
xnor UO_206 (O_206,N_2453,N_2986);
nor UO_207 (O_207,N_2508,N_2506);
xor UO_208 (O_208,N_2775,N_2607);
nand UO_209 (O_209,N_2553,N_2970);
xor UO_210 (O_210,N_2645,N_2845);
nand UO_211 (O_211,N_2709,N_2507);
nand UO_212 (O_212,N_2718,N_2907);
xor UO_213 (O_213,N_2485,N_2884);
and UO_214 (O_214,N_2526,N_2484);
nand UO_215 (O_215,N_2625,N_2713);
nand UO_216 (O_216,N_2919,N_2757);
and UO_217 (O_217,N_2658,N_2779);
or UO_218 (O_218,N_2423,N_2811);
nor UO_219 (O_219,N_2427,N_2547);
xnor UO_220 (O_220,N_2600,N_2533);
nand UO_221 (O_221,N_2876,N_2471);
nand UO_222 (O_222,N_2862,N_2691);
xnor UO_223 (O_223,N_2515,N_2854);
xnor UO_224 (O_224,N_2965,N_2432);
nor UO_225 (O_225,N_2909,N_2679);
xor UO_226 (O_226,N_2540,N_2833);
xnor UO_227 (O_227,N_2633,N_2602);
nand UO_228 (O_228,N_2499,N_2900);
xor UO_229 (O_229,N_2701,N_2492);
and UO_230 (O_230,N_2952,N_2700);
and UO_231 (O_231,N_2433,N_2473);
xor UO_232 (O_232,N_2973,N_2450);
or UO_233 (O_233,N_2561,N_2403);
and UO_234 (O_234,N_2428,N_2934);
xor UO_235 (O_235,N_2840,N_2933);
nand UO_236 (O_236,N_2650,N_2879);
nand UO_237 (O_237,N_2868,N_2814);
nand UO_238 (O_238,N_2717,N_2469);
nor UO_239 (O_239,N_2964,N_2486);
xor UO_240 (O_240,N_2865,N_2989);
nand UO_241 (O_241,N_2913,N_2810);
xor UO_242 (O_242,N_2872,N_2895);
and UO_243 (O_243,N_2514,N_2405);
or UO_244 (O_244,N_2977,N_2612);
and UO_245 (O_245,N_2835,N_2844);
or UO_246 (O_246,N_2817,N_2772);
or UO_247 (O_247,N_2619,N_2482);
and UO_248 (O_248,N_2824,N_2942);
nand UO_249 (O_249,N_2760,N_2687);
or UO_250 (O_250,N_2474,N_2461);
xnor UO_251 (O_251,N_2888,N_2675);
nor UO_252 (O_252,N_2916,N_2777);
nand UO_253 (O_253,N_2454,N_2914);
nor UO_254 (O_254,N_2727,N_2905);
nor UO_255 (O_255,N_2723,N_2624);
xor UO_256 (O_256,N_2944,N_2446);
or UO_257 (O_257,N_2696,N_2503);
nand UO_258 (O_258,N_2903,N_2830);
nor UO_259 (O_259,N_2736,N_2906);
or UO_260 (O_260,N_2684,N_2745);
nand UO_261 (O_261,N_2549,N_2610);
or UO_262 (O_262,N_2797,N_2647);
or UO_263 (O_263,N_2490,N_2785);
nand UO_264 (O_264,N_2420,N_2924);
or UO_265 (O_265,N_2513,N_2930);
nor UO_266 (O_266,N_2685,N_2643);
xnor UO_267 (O_267,N_2867,N_2794);
and UO_268 (O_268,N_2799,N_2504);
and UO_269 (O_269,N_2806,N_2912);
and UO_270 (O_270,N_2452,N_2823);
or UO_271 (O_271,N_2948,N_2939);
nand UO_272 (O_272,N_2921,N_2828);
nor UO_273 (O_273,N_2656,N_2651);
nor UO_274 (O_274,N_2483,N_2999);
nand UO_275 (O_275,N_2590,N_2975);
xnor UO_276 (O_276,N_2536,N_2993);
and UO_277 (O_277,N_2655,N_2764);
xor UO_278 (O_278,N_2877,N_2414);
and UO_279 (O_279,N_2719,N_2518);
nor UO_280 (O_280,N_2630,N_2747);
xor UO_281 (O_281,N_2926,N_2591);
xnor UO_282 (O_282,N_2567,N_2996);
nand UO_283 (O_283,N_2652,N_2627);
nand UO_284 (O_284,N_2592,N_2538);
or UO_285 (O_285,N_2759,N_2847);
or UO_286 (O_286,N_2846,N_2529);
and UO_287 (O_287,N_2641,N_2689);
xor UO_288 (O_288,N_2530,N_2577);
nand UO_289 (O_289,N_2978,N_2501);
or UO_290 (O_290,N_2615,N_2576);
nand UO_291 (O_291,N_2932,N_2573);
or UO_292 (O_292,N_2523,N_2472);
and UO_293 (O_293,N_2807,N_2990);
and UO_294 (O_294,N_2690,N_2401);
nand UO_295 (O_295,N_2620,N_2962);
and UO_296 (O_296,N_2793,N_2730);
xnor UO_297 (O_297,N_2927,N_2768);
and UO_298 (O_298,N_2495,N_2880);
nand UO_299 (O_299,N_2969,N_2519);
and UO_300 (O_300,N_2844,N_2661);
xnor UO_301 (O_301,N_2998,N_2542);
and UO_302 (O_302,N_2854,N_2791);
or UO_303 (O_303,N_2949,N_2513);
xor UO_304 (O_304,N_2880,N_2708);
or UO_305 (O_305,N_2803,N_2757);
and UO_306 (O_306,N_2906,N_2614);
nand UO_307 (O_307,N_2856,N_2990);
nand UO_308 (O_308,N_2806,N_2627);
nand UO_309 (O_309,N_2838,N_2675);
and UO_310 (O_310,N_2449,N_2908);
or UO_311 (O_311,N_2482,N_2542);
or UO_312 (O_312,N_2456,N_2752);
nor UO_313 (O_313,N_2753,N_2582);
xnor UO_314 (O_314,N_2720,N_2631);
xor UO_315 (O_315,N_2743,N_2901);
or UO_316 (O_316,N_2574,N_2514);
nor UO_317 (O_317,N_2680,N_2967);
nor UO_318 (O_318,N_2853,N_2693);
xnor UO_319 (O_319,N_2665,N_2704);
nor UO_320 (O_320,N_2821,N_2469);
nand UO_321 (O_321,N_2836,N_2930);
nand UO_322 (O_322,N_2490,N_2449);
nand UO_323 (O_323,N_2451,N_2693);
nor UO_324 (O_324,N_2993,N_2840);
nand UO_325 (O_325,N_2510,N_2537);
and UO_326 (O_326,N_2745,N_2430);
and UO_327 (O_327,N_2720,N_2453);
nand UO_328 (O_328,N_2579,N_2405);
nand UO_329 (O_329,N_2782,N_2892);
nand UO_330 (O_330,N_2883,N_2812);
and UO_331 (O_331,N_2604,N_2546);
and UO_332 (O_332,N_2479,N_2470);
nand UO_333 (O_333,N_2445,N_2447);
xnor UO_334 (O_334,N_2682,N_2946);
nand UO_335 (O_335,N_2971,N_2473);
xnor UO_336 (O_336,N_2877,N_2600);
nand UO_337 (O_337,N_2997,N_2569);
or UO_338 (O_338,N_2870,N_2451);
and UO_339 (O_339,N_2781,N_2627);
xor UO_340 (O_340,N_2739,N_2798);
nand UO_341 (O_341,N_2756,N_2576);
nand UO_342 (O_342,N_2801,N_2857);
nor UO_343 (O_343,N_2979,N_2480);
and UO_344 (O_344,N_2531,N_2828);
nor UO_345 (O_345,N_2466,N_2503);
nor UO_346 (O_346,N_2784,N_2867);
xnor UO_347 (O_347,N_2732,N_2673);
or UO_348 (O_348,N_2972,N_2703);
nor UO_349 (O_349,N_2893,N_2819);
nand UO_350 (O_350,N_2862,N_2736);
nor UO_351 (O_351,N_2679,N_2688);
nand UO_352 (O_352,N_2750,N_2708);
nand UO_353 (O_353,N_2969,N_2480);
nand UO_354 (O_354,N_2866,N_2425);
and UO_355 (O_355,N_2998,N_2615);
and UO_356 (O_356,N_2579,N_2774);
or UO_357 (O_357,N_2740,N_2866);
or UO_358 (O_358,N_2712,N_2786);
nor UO_359 (O_359,N_2662,N_2974);
nor UO_360 (O_360,N_2818,N_2793);
nor UO_361 (O_361,N_2426,N_2579);
nand UO_362 (O_362,N_2568,N_2693);
and UO_363 (O_363,N_2522,N_2497);
and UO_364 (O_364,N_2845,N_2784);
and UO_365 (O_365,N_2733,N_2536);
xor UO_366 (O_366,N_2614,N_2647);
or UO_367 (O_367,N_2869,N_2720);
and UO_368 (O_368,N_2831,N_2576);
nand UO_369 (O_369,N_2943,N_2932);
or UO_370 (O_370,N_2441,N_2688);
nand UO_371 (O_371,N_2614,N_2669);
nor UO_372 (O_372,N_2813,N_2718);
or UO_373 (O_373,N_2969,N_2454);
and UO_374 (O_374,N_2867,N_2927);
or UO_375 (O_375,N_2790,N_2718);
nand UO_376 (O_376,N_2491,N_2488);
or UO_377 (O_377,N_2566,N_2484);
or UO_378 (O_378,N_2507,N_2977);
nor UO_379 (O_379,N_2569,N_2867);
xor UO_380 (O_380,N_2933,N_2475);
or UO_381 (O_381,N_2636,N_2505);
nor UO_382 (O_382,N_2793,N_2541);
nor UO_383 (O_383,N_2972,N_2861);
nor UO_384 (O_384,N_2919,N_2511);
nor UO_385 (O_385,N_2858,N_2488);
and UO_386 (O_386,N_2404,N_2920);
xor UO_387 (O_387,N_2810,N_2427);
and UO_388 (O_388,N_2888,N_2838);
nor UO_389 (O_389,N_2543,N_2710);
nor UO_390 (O_390,N_2602,N_2946);
xor UO_391 (O_391,N_2627,N_2786);
xnor UO_392 (O_392,N_2936,N_2837);
and UO_393 (O_393,N_2805,N_2520);
and UO_394 (O_394,N_2813,N_2436);
nor UO_395 (O_395,N_2757,N_2427);
xor UO_396 (O_396,N_2404,N_2768);
xnor UO_397 (O_397,N_2740,N_2975);
xnor UO_398 (O_398,N_2619,N_2407);
or UO_399 (O_399,N_2524,N_2602);
or UO_400 (O_400,N_2518,N_2896);
xnor UO_401 (O_401,N_2684,N_2482);
nor UO_402 (O_402,N_2581,N_2912);
nand UO_403 (O_403,N_2843,N_2485);
and UO_404 (O_404,N_2787,N_2497);
nor UO_405 (O_405,N_2967,N_2950);
or UO_406 (O_406,N_2413,N_2811);
nand UO_407 (O_407,N_2937,N_2501);
nor UO_408 (O_408,N_2414,N_2472);
xnor UO_409 (O_409,N_2930,N_2451);
nor UO_410 (O_410,N_2822,N_2513);
nor UO_411 (O_411,N_2639,N_2897);
and UO_412 (O_412,N_2430,N_2553);
xnor UO_413 (O_413,N_2570,N_2592);
nor UO_414 (O_414,N_2742,N_2927);
or UO_415 (O_415,N_2487,N_2779);
nand UO_416 (O_416,N_2615,N_2689);
nand UO_417 (O_417,N_2863,N_2561);
or UO_418 (O_418,N_2990,N_2684);
and UO_419 (O_419,N_2468,N_2612);
or UO_420 (O_420,N_2933,N_2682);
nand UO_421 (O_421,N_2734,N_2599);
or UO_422 (O_422,N_2836,N_2595);
or UO_423 (O_423,N_2456,N_2975);
and UO_424 (O_424,N_2447,N_2733);
xor UO_425 (O_425,N_2602,N_2761);
xor UO_426 (O_426,N_2428,N_2749);
and UO_427 (O_427,N_2843,N_2902);
and UO_428 (O_428,N_2959,N_2678);
nor UO_429 (O_429,N_2986,N_2889);
nor UO_430 (O_430,N_2449,N_2721);
or UO_431 (O_431,N_2721,N_2741);
nor UO_432 (O_432,N_2671,N_2795);
and UO_433 (O_433,N_2772,N_2494);
nor UO_434 (O_434,N_2693,N_2489);
and UO_435 (O_435,N_2411,N_2860);
and UO_436 (O_436,N_2645,N_2742);
xor UO_437 (O_437,N_2520,N_2958);
or UO_438 (O_438,N_2501,N_2731);
or UO_439 (O_439,N_2842,N_2913);
and UO_440 (O_440,N_2486,N_2683);
nand UO_441 (O_441,N_2829,N_2572);
nor UO_442 (O_442,N_2446,N_2465);
or UO_443 (O_443,N_2816,N_2931);
and UO_444 (O_444,N_2903,N_2820);
and UO_445 (O_445,N_2448,N_2892);
or UO_446 (O_446,N_2459,N_2676);
or UO_447 (O_447,N_2855,N_2422);
or UO_448 (O_448,N_2979,N_2791);
nand UO_449 (O_449,N_2772,N_2713);
nor UO_450 (O_450,N_2573,N_2639);
or UO_451 (O_451,N_2558,N_2978);
or UO_452 (O_452,N_2772,N_2846);
and UO_453 (O_453,N_2677,N_2675);
xor UO_454 (O_454,N_2680,N_2459);
nor UO_455 (O_455,N_2652,N_2766);
xor UO_456 (O_456,N_2930,N_2437);
nand UO_457 (O_457,N_2699,N_2967);
xnor UO_458 (O_458,N_2857,N_2619);
xnor UO_459 (O_459,N_2671,N_2673);
xnor UO_460 (O_460,N_2978,N_2508);
or UO_461 (O_461,N_2828,N_2561);
nand UO_462 (O_462,N_2472,N_2844);
nand UO_463 (O_463,N_2738,N_2707);
or UO_464 (O_464,N_2742,N_2673);
and UO_465 (O_465,N_2771,N_2522);
or UO_466 (O_466,N_2747,N_2725);
nor UO_467 (O_467,N_2911,N_2529);
nor UO_468 (O_468,N_2403,N_2682);
and UO_469 (O_469,N_2784,N_2636);
and UO_470 (O_470,N_2587,N_2654);
nand UO_471 (O_471,N_2878,N_2696);
and UO_472 (O_472,N_2885,N_2419);
xor UO_473 (O_473,N_2558,N_2469);
xnor UO_474 (O_474,N_2911,N_2990);
nand UO_475 (O_475,N_2760,N_2900);
nor UO_476 (O_476,N_2901,N_2417);
and UO_477 (O_477,N_2774,N_2897);
or UO_478 (O_478,N_2466,N_2911);
nor UO_479 (O_479,N_2522,N_2707);
nand UO_480 (O_480,N_2647,N_2618);
nand UO_481 (O_481,N_2841,N_2655);
or UO_482 (O_482,N_2836,N_2768);
or UO_483 (O_483,N_2922,N_2747);
nor UO_484 (O_484,N_2891,N_2973);
nor UO_485 (O_485,N_2420,N_2736);
and UO_486 (O_486,N_2803,N_2593);
xnor UO_487 (O_487,N_2532,N_2546);
nand UO_488 (O_488,N_2699,N_2743);
nand UO_489 (O_489,N_2695,N_2643);
nor UO_490 (O_490,N_2676,N_2412);
nand UO_491 (O_491,N_2440,N_2983);
and UO_492 (O_492,N_2761,N_2633);
nor UO_493 (O_493,N_2503,N_2469);
nor UO_494 (O_494,N_2782,N_2647);
nor UO_495 (O_495,N_2879,N_2830);
nand UO_496 (O_496,N_2463,N_2619);
xor UO_497 (O_497,N_2828,N_2966);
nand UO_498 (O_498,N_2858,N_2906);
nand UO_499 (O_499,N_2767,N_2930);
endmodule