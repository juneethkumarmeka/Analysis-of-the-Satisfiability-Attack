module basic_750_5000_1000_25_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_296,In_687);
xor U1 (N_1,In_178,In_591);
nor U2 (N_2,In_664,In_146);
nand U3 (N_3,In_733,In_278);
nor U4 (N_4,In_62,In_127);
and U5 (N_5,In_448,In_217);
or U6 (N_6,In_310,In_379);
and U7 (N_7,In_130,In_507);
nand U8 (N_8,In_395,In_245);
and U9 (N_9,In_414,In_588);
and U10 (N_10,In_315,In_299);
nor U11 (N_11,In_143,In_432);
nand U12 (N_12,In_51,In_479);
xnor U13 (N_13,In_439,In_242);
or U14 (N_14,In_698,In_558);
xor U15 (N_15,In_683,In_602);
and U16 (N_16,In_631,In_271);
nand U17 (N_17,In_19,In_89);
or U18 (N_18,In_576,In_684);
and U19 (N_19,In_605,In_304);
and U20 (N_20,In_616,In_423);
and U21 (N_21,In_489,In_279);
nand U22 (N_22,In_107,In_693);
and U23 (N_23,In_510,In_565);
nand U24 (N_24,In_390,In_167);
and U25 (N_25,In_206,In_343);
nand U26 (N_26,In_42,In_268);
or U27 (N_27,In_111,In_416);
nand U28 (N_28,In_313,In_524);
nand U29 (N_29,In_248,In_504);
xor U30 (N_30,In_728,In_727);
xnor U31 (N_31,In_531,In_476);
and U32 (N_32,In_338,In_696);
xor U33 (N_33,In_451,In_475);
nand U34 (N_34,In_653,In_282);
xor U35 (N_35,In_17,In_35);
nor U36 (N_36,In_73,In_166);
nor U37 (N_37,In_470,In_309);
xnor U38 (N_38,In_397,In_4);
nor U39 (N_39,In_205,In_411);
and U40 (N_40,In_552,In_610);
or U41 (N_41,In_612,In_140);
nand U42 (N_42,In_224,In_142);
nor U43 (N_43,In_615,In_695);
or U44 (N_44,In_704,In_240);
nand U45 (N_45,In_298,In_102);
xnor U46 (N_46,In_160,In_462);
and U47 (N_47,In_219,In_74);
nor U48 (N_48,In_368,In_287);
nand U49 (N_49,In_633,In_596);
nor U50 (N_50,In_52,In_699);
and U51 (N_51,In_460,In_503);
xnor U52 (N_52,In_163,In_720);
xor U53 (N_53,In_647,In_208);
nor U54 (N_54,In_125,In_77);
and U55 (N_55,In_98,In_274);
or U56 (N_56,In_276,In_249);
and U57 (N_57,In_63,In_294);
nand U58 (N_58,In_553,In_614);
nand U59 (N_59,In_133,In_64);
nor U60 (N_60,In_179,In_50);
and U61 (N_61,In_594,In_361);
or U62 (N_62,In_663,In_95);
or U63 (N_63,In_40,In_353);
xnor U64 (N_64,In_227,In_263);
nand U65 (N_65,In_480,In_275);
nand U66 (N_66,In_264,In_120);
and U67 (N_67,In_430,In_478);
nand U68 (N_68,In_20,In_185);
and U69 (N_69,In_141,In_690);
or U70 (N_70,In_86,In_376);
xnor U71 (N_71,In_446,In_642);
nor U72 (N_72,In_578,In_307);
nand U73 (N_73,In_444,In_60);
nor U74 (N_74,In_389,In_721);
xor U75 (N_75,In_466,In_449);
or U76 (N_76,In_237,In_54);
nand U77 (N_77,In_335,In_210);
or U78 (N_78,In_300,In_494);
xnor U79 (N_79,In_427,In_403);
nand U80 (N_80,In_247,In_732);
and U81 (N_81,In_169,In_593);
xor U82 (N_82,In_398,In_316);
and U83 (N_83,In_406,In_676);
nand U84 (N_84,In_260,In_600);
nand U85 (N_85,In_546,In_645);
nand U86 (N_86,In_168,In_628);
or U87 (N_87,In_221,In_649);
nor U88 (N_88,In_27,In_743);
xnor U89 (N_89,In_14,In_196);
xor U90 (N_90,In_291,In_41);
nor U91 (N_91,In_575,In_362);
or U92 (N_92,In_204,In_409);
nand U93 (N_93,In_380,In_270);
and U94 (N_94,In_155,In_584);
nor U95 (N_95,In_233,In_443);
or U96 (N_96,In_655,In_400);
nand U97 (N_97,In_289,In_528);
nor U98 (N_98,In_530,In_734);
nor U99 (N_99,In_746,In_378);
nand U100 (N_100,In_29,In_319);
xor U101 (N_101,In_738,In_30);
nor U102 (N_102,In_719,In_214);
nand U103 (N_103,In_486,In_230);
nand U104 (N_104,In_290,In_326);
or U105 (N_105,In_177,In_59);
and U106 (N_106,In_48,In_556);
and U107 (N_107,In_660,In_391);
xnor U108 (N_108,In_190,In_635);
and U109 (N_109,In_356,In_641);
xor U110 (N_110,In_691,In_547);
nand U111 (N_111,In_682,In_492);
nor U112 (N_112,In_648,In_405);
nand U113 (N_113,In_656,In_498);
and U114 (N_114,In_363,In_694);
and U115 (N_115,In_408,In_567);
nor U116 (N_116,In_535,In_350);
nor U117 (N_117,In_147,In_393);
and U118 (N_118,In_198,In_428);
or U119 (N_119,In_424,In_108);
nand U120 (N_120,In_659,In_372);
or U121 (N_121,In_78,In_212);
and U122 (N_122,In_105,In_110);
nor U123 (N_123,In_638,In_716);
or U124 (N_124,In_231,In_415);
xnor U125 (N_125,In_392,In_117);
nor U126 (N_126,In_500,In_717);
and U127 (N_127,In_550,In_261);
xor U128 (N_128,In_139,In_506);
xnor U129 (N_129,In_213,In_606);
and U130 (N_130,In_624,In_144);
xnor U131 (N_131,In_431,In_657);
nor U132 (N_132,In_562,In_164);
xnor U133 (N_133,In_170,In_99);
or U134 (N_134,In_417,In_65);
nor U135 (N_135,In_412,In_33);
xor U136 (N_136,In_202,In_297);
nand U137 (N_137,In_607,In_452);
or U138 (N_138,In_336,In_109);
nor U139 (N_139,In_548,In_92);
nand U140 (N_140,In_436,In_679);
or U141 (N_141,In_188,In_235);
and U142 (N_142,In_238,In_135);
xnor U143 (N_143,In_723,In_499);
xnor U144 (N_144,In_106,In_341);
nand U145 (N_145,In_345,In_21);
and U146 (N_146,In_288,In_228);
nand U147 (N_147,In_455,In_613);
and U148 (N_148,In_697,In_440);
or U149 (N_149,In_311,In_599);
xor U150 (N_150,In_467,In_129);
xnor U151 (N_151,In_515,In_75);
or U152 (N_152,In_103,In_673);
nor U153 (N_153,In_173,In_201);
and U154 (N_154,In_61,In_6);
and U155 (N_155,In_355,In_68);
nor U156 (N_156,In_601,In_465);
nor U157 (N_157,In_241,In_150);
nand U158 (N_158,In_239,In_364);
nor U159 (N_159,In_730,In_207);
xnor U160 (N_160,In_681,In_488);
nand U161 (N_161,In_484,In_737);
and U162 (N_162,In_722,In_573);
nand U163 (N_163,In_453,In_23);
nor U164 (N_164,In_72,In_555);
nand U165 (N_165,In_331,In_585);
and U166 (N_166,In_445,In_579);
or U167 (N_167,In_10,In_183);
and U168 (N_168,In_592,In_564);
xnor U169 (N_169,In_458,In_90);
nand U170 (N_170,In_113,In_273);
or U171 (N_171,In_124,In_701);
and U172 (N_172,In_158,In_323);
nand U173 (N_173,In_385,In_25);
and U174 (N_174,In_388,In_262);
nand U175 (N_175,In_157,In_182);
xor U176 (N_176,In_677,In_344);
nand U177 (N_177,In_570,In_623);
nand U178 (N_178,In_636,In_193);
nand U179 (N_179,In_724,In_327);
or U180 (N_180,In_748,In_561);
nand U181 (N_181,In_747,In_357);
and U182 (N_182,In_442,In_700);
nand U183 (N_183,In_454,In_303);
nand U184 (N_184,In_354,In_122);
and U185 (N_185,In_469,In_671);
or U186 (N_186,In_83,In_349);
nand U187 (N_187,In_666,In_640);
or U188 (N_188,In_580,In_121);
nand U189 (N_189,In_373,In_493);
or U190 (N_190,In_209,In_348);
xor U191 (N_191,In_46,In_496);
xnor U192 (N_192,In_662,In_726);
nor U193 (N_193,In_24,In_324);
xor U194 (N_194,In_587,In_710);
nor U195 (N_195,In_80,In_487);
nor U196 (N_196,In_292,In_251);
xnor U197 (N_197,In_330,In_329);
xnor U198 (N_198,In_149,In_401);
xnor U199 (N_199,In_554,In_632);
nand U200 (N_200,N_67,In_617);
xor U201 (N_201,N_191,N_74);
or U202 (N_202,N_89,In_200);
nor U203 (N_203,In_119,In_171);
or U204 (N_204,In_243,In_540);
and U205 (N_205,In_560,In_334);
and U206 (N_206,In_36,N_155);
nor U207 (N_207,N_54,In_386);
xnor U208 (N_208,N_110,In_429);
and U209 (N_209,In_96,N_85);
xor U210 (N_210,In_82,In_229);
or U211 (N_211,N_70,In_630);
nand U212 (N_212,N_186,In_661);
xnor U213 (N_213,In_351,In_384);
or U214 (N_214,In_598,In_172);
nand U215 (N_215,In_69,In_520);
nand U216 (N_216,N_190,In_277);
xnor U217 (N_217,N_197,In_250);
nor U218 (N_218,In_625,N_167);
nor U219 (N_219,N_195,In_57);
and U220 (N_220,In_162,In_367);
and U221 (N_221,N_150,In_670);
xnor U222 (N_222,In_634,In_337);
xnor U223 (N_223,In_123,N_5);
nor U224 (N_224,In_322,In_501);
or U225 (N_225,N_13,In_114);
xor U226 (N_226,In_32,In_218);
or U227 (N_227,In_513,In_340);
and U228 (N_228,In_518,In_739);
and U229 (N_229,In_609,N_108);
or U230 (N_230,N_68,In_132);
or U231 (N_231,In_643,In_740);
nand U232 (N_232,In_509,In_187);
or U233 (N_233,N_77,In_413);
xnor U234 (N_234,In_490,In_58);
xnor U235 (N_235,In_2,In_718);
xor U236 (N_236,In_269,N_21);
nand U237 (N_237,In_244,N_84);
nor U238 (N_238,In_749,In_101);
nor U239 (N_239,N_109,In_543);
nor U240 (N_240,In_136,In_549);
xor U241 (N_241,N_105,In_712);
nand U242 (N_242,N_174,In_474);
nor U243 (N_243,N_153,In_394);
and U244 (N_244,In_191,In_45);
and U245 (N_245,N_20,In_399);
xnor U246 (N_246,In_174,In_654);
and U247 (N_247,In_104,N_57);
and U248 (N_248,N_199,In_538);
nor U249 (N_249,N_114,In_468);
xnor U250 (N_250,N_137,N_160);
and U251 (N_251,N_158,In_708);
nand U252 (N_252,In_346,In_620);
nand U253 (N_253,N_187,In_665);
xor U254 (N_254,In_582,In_521);
nor U255 (N_255,N_128,N_151);
nand U256 (N_256,N_177,In_265);
nor U257 (N_257,In_450,In_280);
or U258 (N_258,In_175,N_168);
nand U259 (N_259,In_371,N_170);
nor U260 (N_260,In_745,In_321);
nand U261 (N_261,In_225,In_369);
and U262 (N_262,N_59,N_107);
nand U263 (N_263,In_541,In_539);
or U264 (N_264,In_502,N_61);
nand U265 (N_265,In_542,N_1);
and U266 (N_266,N_69,In_644);
and U267 (N_267,N_90,In_529);
nand U268 (N_268,In_590,In_159);
nand U269 (N_269,N_164,In_13);
xnor U270 (N_270,N_0,In_199);
and U271 (N_271,In_674,N_42);
nor U272 (N_272,In_472,In_646);
and U273 (N_273,In_669,In_161);
nand U274 (N_274,N_104,N_181);
nor U275 (N_275,In_544,In_258);
nor U276 (N_276,N_72,In_94);
and U277 (N_277,In_483,N_118);
or U278 (N_278,N_198,In_128);
or U279 (N_279,N_83,N_183);
nand U280 (N_280,In_464,In_627);
nand U281 (N_281,In_639,In_332);
xor U282 (N_282,N_75,In_203);
nand U283 (N_283,In_622,In_286);
nor U284 (N_284,In_744,In_482);
and U285 (N_285,In_195,In_481);
xor U286 (N_286,In_545,In_281);
nand U287 (N_287,N_119,In_381);
and U288 (N_288,N_166,In_581);
nor U289 (N_289,In_216,N_6);
and U290 (N_290,In_255,N_113);
nor U291 (N_291,In_537,In_595);
or U292 (N_292,In_477,In_688);
nor U293 (N_293,In_709,In_256);
or U294 (N_294,N_88,In_112);
and U295 (N_295,N_14,In_731);
and U296 (N_296,N_79,In_67);
nor U297 (N_297,In_49,N_26);
or U298 (N_298,N_65,N_97);
nor U299 (N_299,In_618,In_266);
nand U300 (N_300,N_162,In_320);
or U301 (N_301,N_71,N_34);
or U302 (N_302,N_11,In_729);
and U303 (N_303,In_715,N_98);
nand U304 (N_304,N_175,In_66);
nor U305 (N_305,In_88,In_586);
or U306 (N_306,In_713,In_735);
or U307 (N_307,In_360,In_736);
nor U308 (N_308,In_211,N_149);
and U309 (N_309,In_421,In_220);
and U310 (N_310,N_134,In_650);
xnor U311 (N_311,N_62,N_52);
nor U312 (N_312,N_133,In_28);
or U313 (N_313,In_253,In_418);
nand U314 (N_314,In_559,N_82);
or U315 (N_315,In_192,In_306);
and U316 (N_316,N_116,In_44);
or U317 (N_317,In_711,In_608);
or U318 (N_318,In_495,N_124);
nor U319 (N_319,In_151,In_404);
xnor U320 (N_320,In_680,In_437);
or U321 (N_321,In_226,In_689);
xor U322 (N_322,In_377,In_512);
nor U323 (N_323,N_95,In_370);
and U324 (N_324,In_153,In_55);
and U325 (N_325,N_185,N_148);
and U326 (N_326,N_171,In_145);
xor U327 (N_327,In_38,N_101);
or U328 (N_328,N_127,In_53);
xor U329 (N_329,N_178,N_152);
xnor U330 (N_330,In_569,N_45);
xnor U331 (N_331,In_16,N_86);
xnor U332 (N_332,N_23,N_56);
or U333 (N_333,N_92,N_51);
and U334 (N_334,N_120,N_46);
nor U335 (N_335,In_742,In_511);
nand U336 (N_336,N_49,In_246);
nor U337 (N_337,In_284,In_619);
or U338 (N_338,In_165,In_116);
or U339 (N_339,In_637,In_456);
and U340 (N_340,N_16,In_402);
nor U341 (N_341,N_136,In_115);
or U342 (N_342,N_100,In_47);
xor U343 (N_343,N_126,N_32);
nor U344 (N_344,N_138,In_508);
or U345 (N_345,In_222,In_525);
and U346 (N_346,In_7,N_180);
or U347 (N_347,In_604,In_197);
or U348 (N_348,N_163,N_40);
xor U349 (N_349,N_188,In_232);
nor U350 (N_350,N_142,N_29);
or U351 (N_351,N_4,In_447);
nand U352 (N_352,In_522,N_176);
nor U353 (N_353,N_81,In_534);
nor U354 (N_354,In_84,In_485);
and U355 (N_355,N_129,In_589);
nand U356 (N_356,In_705,In_497);
xor U357 (N_357,N_159,In_410);
nor U358 (N_358,N_55,N_154);
xnor U359 (N_359,In_473,N_172);
or U360 (N_360,In_37,In_312);
xor U361 (N_361,N_194,N_25);
and U362 (N_362,In_667,N_196);
xor U363 (N_363,In_56,In_523);
nor U364 (N_364,N_27,In_678);
and U365 (N_365,In_365,In_422);
nand U366 (N_366,In_31,In_505);
and U367 (N_367,In_741,N_161);
xor U368 (N_368,N_39,In_272);
or U369 (N_369,N_106,N_10);
xor U370 (N_370,In_22,In_305);
nand U371 (N_371,In_461,In_252);
nand U372 (N_372,N_24,N_165);
or U373 (N_373,N_94,N_31);
nor U374 (N_374,N_7,N_140);
xor U375 (N_375,In_574,In_257);
xnor U376 (N_376,In_184,In_533);
xor U377 (N_377,In_76,In_434);
and U378 (N_378,In_725,In_342);
nand U379 (N_379,N_173,In_134);
xnor U380 (N_380,N_38,N_103);
nor U381 (N_381,In_419,In_152);
or U382 (N_382,N_48,In_675);
xor U383 (N_383,In_176,N_135);
and U384 (N_384,In_1,In_15);
xor U385 (N_385,In_70,In_491);
xnor U386 (N_386,In_519,In_536);
and U387 (N_387,N_43,In_435);
nand U388 (N_388,In_532,In_426);
nand U389 (N_389,In_420,In_557);
or U390 (N_390,In_97,N_80);
or U391 (N_391,N_143,N_58);
nor U392 (N_392,In_626,N_130);
and U393 (N_393,In_9,In_156);
nand U394 (N_394,N_139,In_514);
nand U395 (N_395,N_179,N_145);
xor U396 (N_396,N_53,In_285);
or U397 (N_397,In_79,In_407);
nand U398 (N_398,In_375,In_18);
and U399 (N_399,In_267,In_39);
xor U400 (N_400,In_71,In_629);
nand U401 (N_401,N_131,N_325);
xnor U402 (N_402,N_182,N_339);
or U403 (N_403,N_318,N_392);
or U404 (N_404,N_353,N_327);
nor U405 (N_405,N_326,N_316);
nand U406 (N_406,N_393,N_269);
and U407 (N_407,N_245,N_300);
and U408 (N_408,In_471,In_571);
xnor U409 (N_409,N_337,In_180);
nand U410 (N_410,N_41,In_714);
nor U411 (N_411,N_141,N_382);
xor U412 (N_412,N_322,In_131);
xor U413 (N_413,N_303,N_351);
xor U414 (N_414,N_33,In_707);
nor U415 (N_415,N_364,N_380);
nand U416 (N_416,In_317,N_271);
and U417 (N_417,N_146,N_30);
nand U418 (N_418,In_382,In_181);
or U419 (N_419,N_347,N_125);
xor U420 (N_420,N_17,N_225);
and U421 (N_421,N_263,In_527);
nor U422 (N_422,N_201,N_367);
nor U423 (N_423,N_28,N_102);
nor U424 (N_424,N_76,N_144);
nor U425 (N_425,N_3,N_390);
xor U426 (N_426,In_118,N_329);
or U427 (N_427,N_214,In_441);
nor U428 (N_428,In_314,N_264);
nand U429 (N_429,N_284,N_292);
or U430 (N_430,N_206,N_233);
xnor U431 (N_431,In_672,In_283);
xnor U432 (N_432,N_12,N_267);
or U433 (N_433,N_239,N_247);
xor U434 (N_434,N_202,In_5);
nand U435 (N_435,In_702,N_213);
and U436 (N_436,In_100,N_352);
nor U437 (N_437,N_112,N_37);
or U438 (N_438,N_323,N_304);
nor U439 (N_439,In_658,N_223);
nor U440 (N_440,In_11,N_336);
or U441 (N_441,N_372,N_258);
xor U442 (N_442,N_246,N_276);
nand U443 (N_443,In_0,N_219);
xnor U444 (N_444,In_597,N_357);
nand U445 (N_445,In_577,N_47);
nor U446 (N_446,In_457,N_262);
and U447 (N_447,In_234,N_250);
and U448 (N_448,In_215,N_282);
and U449 (N_449,In_583,N_391);
nor U450 (N_450,N_272,N_63);
nand U451 (N_451,In_551,In_526);
and U452 (N_452,N_121,In_686);
nand U453 (N_453,N_8,N_273);
and U454 (N_454,N_240,N_231);
nor U455 (N_455,In_685,N_111);
or U456 (N_456,N_279,N_343);
or U457 (N_457,N_311,N_302);
nand U458 (N_458,N_294,N_365);
and U459 (N_459,N_312,N_342);
nor U460 (N_460,In_358,N_232);
or U461 (N_461,N_355,In_87);
xor U462 (N_462,N_259,N_338);
and U463 (N_463,N_346,In_236);
or U464 (N_464,In_301,N_78);
or U465 (N_465,N_189,N_288);
and U466 (N_466,N_50,N_257);
and U467 (N_467,In_359,N_394);
nand U468 (N_468,N_200,N_387);
or U469 (N_469,N_384,In_194);
nor U470 (N_470,In_563,N_370);
nand U471 (N_471,N_383,N_209);
nor U472 (N_472,N_243,In_568);
nor U473 (N_473,N_377,N_184);
nand U474 (N_474,N_331,N_235);
nand U475 (N_475,N_253,N_252);
and U476 (N_476,N_397,N_334);
nand U477 (N_477,In_295,N_275);
or U478 (N_478,N_374,N_360);
nand U479 (N_479,N_99,N_362);
nand U480 (N_480,N_255,In_259);
nand U481 (N_481,N_324,N_328);
xnor U482 (N_482,N_22,N_244);
xnor U483 (N_483,In_516,In_328);
nand U484 (N_484,In_366,In_463);
or U485 (N_485,N_283,N_216);
or U486 (N_486,N_96,In_651);
nor U487 (N_487,N_385,N_297);
nand U488 (N_488,In_293,In_396);
or U489 (N_489,N_280,In_387);
or U490 (N_490,N_93,N_317);
and U491 (N_491,N_295,N_251);
and U492 (N_492,N_217,N_345);
or U493 (N_493,N_132,N_36);
xor U494 (N_494,N_254,In_8);
nand U495 (N_495,N_375,N_386);
xor U496 (N_496,N_308,In_374);
or U497 (N_497,In_148,N_220);
or U498 (N_498,In_706,In_138);
nor U499 (N_499,N_291,N_274);
and U500 (N_500,In_85,In_137);
nor U501 (N_501,N_44,N_281);
nand U502 (N_502,In_308,N_147);
or U503 (N_503,N_289,N_237);
or U504 (N_504,In_347,N_379);
nor U505 (N_505,N_354,N_224);
or U506 (N_506,N_348,N_315);
nand U507 (N_507,In_126,N_277);
nand U508 (N_508,N_115,N_286);
or U509 (N_509,N_366,N_230);
nor U510 (N_510,N_285,N_398);
or U511 (N_511,N_301,N_330);
and U512 (N_512,N_361,In_566);
nand U513 (N_513,N_320,N_395);
xor U514 (N_514,In_186,N_376);
nor U515 (N_515,N_310,N_241);
xor U516 (N_516,N_396,N_91);
nand U517 (N_517,N_210,N_228);
or U518 (N_518,N_293,N_156);
xnor U519 (N_519,N_123,N_333);
and U520 (N_520,N_73,N_358);
xor U521 (N_521,N_321,N_60);
nand U522 (N_522,N_332,N_221);
nor U523 (N_523,N_211,N_2);
xnor U524 (N_524,In_517,N_205);
xnor U525 (N_525,In_333,N_169);
and U526 (N_526,In_26,In_572);
nor U527 (N_527,N_290,N_212);
and U528 (N_528,N_204,In_325);
and U529 (N_529,N_122,In_318);
xor U530 (N_530,N_287,N_238);
nor U531 (N_531,N_309,N_15);
nor U532 (N_532,N_35,In_12);
nor U533 (N_533,In_91,In_154);
xor U534 (N_534,N_234,N_319);
and U535 (N_535,N_249,In_425);
or U536 (N_536,In_383,In_3);
and U537 (N_537,N_359,In_302);
nor U538 (N_538,N_314,N_296);
nor U539 (N_539,In_339,N_260);
nand U540 (N_540,N_229,N_207);
nor U541 (N_541,N_270,N_389);
or U542 (N_542,In_34,N_222);
and U543 (N_543,N_335,N_349);
nor U544 (N_544,N_388,N_218);
and U545 (N_545,In_93,In_189);
nand U546 (N_546,N_371,In_668);
and U547 (N_547,N_192,N_307);
or U548 (N_548,N_193,N_299);
xor U549 (N_549,N_369,N_265);
and U550 (N_550,N_399,In_43);
nor U551 (N_551,N_344,N_340);
nor U552 (N_552,N_157,In_692);
or U553 (N_553,N_278,N_378);
or U554 (N_554,In_223,N_19);
xor U555 (N_555,N_256,N_363);
xor U556 (N_556,N_117,N_305);
or U557 (N_557,N_373,N_368);
xnor U558 (N_558,N_87,In_621);
xnor U559 (N_559,N_203,N_313);
nand U560 (N_560,N_64,N_341);
or U561 (N_561,N_350,N_381);
xnor U562 (N_562,In_433,N_66);
nor U563 (N_563,N_242,In_459);
nand U564 (N_564,In_603,In_703);
nand U565 (N_565,N_208,In_81);
or U566 (N_566,N_236,N_261);
nor U567 (N_567,N_9,N_298);
and U568 (N_568,In_652,N_268);
and U569 (N_569,N_18,In_352);
or U570 (N_570,N_266,In_611);
nor U571 (N_571,N_248,N_226);
or U572 (N_572,N_215,N_227);
nand U573 (N_573,N_306,N_356);
nand U574 (N_574,In_438,In_254);
nand U575 (N_575,N_221,N_333);
and U576 (N_576,In_566,N_307);
or U577 (N_577,N_259,N_60);
nor U578 (N_578,In_154,N_117);
or U579 (N_579,N_203,N_66);
xnor U580 (N_580,In_571,N_271);
nor U581 (N_581,N_316,N_231);
or U582 (N_582,N_381,N_348);
or U583 (N_583,In_366,In_137);
xnor U584 (N_584,N_50,N_373);
xor U585 (N_585,N_233,N_295);
and U586 (N_586,N_338,N_217);
or U587 (N_587,N_189,N_367);
nor U588 (N_588,N_112,In_583);
xor U589 (N_589,N_209,N_131);
and U590 (N_590,N_253,N_235);
nor U591 (N_591,N_394,N_376);
or U592 (N_592,N_93,In_551);
nand U593 (N_593,N_319,N_226);
xor U594 (N_594,N_358,N_201);
or U595 (N_595,N_37,N_279);
xor U596 (N_596,In_302,N_230);
or U597 (N_597,N_295,N_169);
nand U598 (N_598,N_264,N_322);
and U599 (N_599,N_33,N_373);
or U600 (N_600,N_413,N_492);
nand U601 (N_601,N_497,N_569);
xor U602 (N_602,N_488,N_504);
and U603 (N_603,N_559,N_468);
xnor U604 (N_604,N_484,N_563);
nand U605 (N_605,N_575,N_415);
nor U606 (N_606,N_580,N_477);
and U607 (N_607,N_576,N_452);
xnor U608 (N_608,N_540,N_402);
and U609 (N_609,N_574,N_500);
nand U610 (N_610,N_437,N_425);
and U611 (N_611,N_522,N_572);
nor U612 (N_612,N_419,N_403);
nand U613 (N_613,N_533,N_406);
xor U614 (N_614,N_471,N_463);
nand U615 (N_615,N_486,N_557);
xnor U616 (N_616,N_582,N_470);
or U617 (N_617,N_536,N_493);
or U618 (N_618,N_567,N_547);
and U619 (N_619,N_561,N_469);
and U620 (N_620,N_476,N_479);
nor U621 (N_621,N_515,N_573);
xnor U622 (N_622,N_441,N_458);
and U623 (N_623,N_495,N_583);
xnor U624 (N_624,N_592,N_496);
nor U625 (N_625,N_499,N_439);
nor U626 (N_626,N_581,N_404);
or U627 (N_627,N_435,N_475);
or U628 (N_628,N_528,N_598);
xnor U629 (N_629,N_412,N_445);
xnor U630 (N_630,N_498,N_487);
and U631 (N_631,N_449,N_448);
xnor U632 (N_632,N_570,N_537);
nor U633 (N_633,N_503,N_507);
or U634 (N_634,N_442,N_418);
and U635 (N_635,N_524,N_532);
or U636 (N_636,N_485,N_424);
xnor U637 (N_637,N_473,N_490);
nor U638 (N_638,N_599,N_446);
or U639 (N_639,N_467,N_544);
or U640 (N_640,N_502,N_541);
and U641 (N_641,N_508,N_505);
and U642 (N_642,N_593,N_506);
xor U643 (N_643,N_578,N_545);
nand U644 (N_644,N_440,N_595);
xnor U645 (N_645,N_564,N_512);
and U646 (N_646,N_494,N_480);
and U647 (N_647,N_405,N_552);
xor U648 (N_648,N_596,N_565);
or U649 (N_649,N_509,N_481);
and U650 (N_650,N_436,N_514);
nand U651 (N_651,N_417,N_450);
or U652 (N_652,N_411,N_579);
nor U653 (N_653,N_433,N_453);
nor U654 (N_654,N_516,N_531);
nor U655 (N_655,N_438,N_517);
xnor U656 (N_656,N_549,N_421);
nand U657 (N_657,N_428,N_482);
or U658 (N_658,N_401,N_529);
or U659 (N_659,N_587,N_414);
and U660 (N_660,N_423,N_597);
and U661 (N_661,N_427,N_555);
nor U662 (N_662,N_571,N_584);
nor U663 (N_663,N_556,N_489);
nand U664 (N_664,N_539,N_478);
or U665 (N_665,N_407,N_457);
nand U666 (N_666,N_543,N_594);
nand U667 (N_667,N_526,N_548);
xnor U668 (N_668,N_432,N_444);
nand U669 (N_669,N_461,N_525);
and U670 (N_670,N_429,N_562);
and U671 (N_671,N_520,N_410);
and U672 (N_672,N_542,N_586);
and U673 (N_673,N_568,N_523);
nand U674 (N_674,N_501,N_431);
and U675 (N_675,N_430,N_558);
or U676 (N_676,N_546,N_513);
or U677 (N_677,N_577,N_534);
and U678 (N_678,N_589,N_451);
or U679 (N_679,N_535,N_538);
and U680 (N_680,N_416,N_459);
nand U681 (N_681,N_551,N_462);
and U682 (N_682,N_519,N_426);
nand U683 (N_683,N_554,N_465);
and U684 (N_684,N_447,N_466);
xor U685 (N_685,N_518,N_527);
and U686 (N_686,N_483,N_422);
and U687 (N_687,N_454,N_511);
and U688 (N_688,N_464,N_460);
nor U689 (N_689,N_530,N_456);
and U690 (N_690,N_409,N_590);
xnor U691 (N_691,N_491,N_521);
nor U692 (N_692,N_400,N_510);
and U693 (N_693,N_591,N_553);
nor U694 (N_694,N_472,N_550);
nor U695 (N_695,N_420,N_560);
and U696 (N_696,N_434,N_588);
and U697 (N_697,N_566,N_443);
and U698 (N_698,N_474,N_455);
nand U699 (N_699,N_408,N_585);
xnor U700 (N_700,N_566,N_462);
or U701 (N_701,N_523,N_561);
or U702 (N_702,N_413,N_557);
xnor U703 (N_703,N_535,N_561);
nand U704 (N_704,N_434,N_445);
or U705 (N_705,N_572,N_575);
nand U706 (N_706,N_472,N_599);
nor U707 (N_707,N_412,N_516);
nand U708 (N_708,N_474,N_551);
and U709 (N_709,N_473,N_438);
or U710 (N_710,N_544,N_489);
nor U711 (N_711,N_518,N_547);
nor U712 (N_712,N_530,N_491);
and U713 (N_713,N_445,N_430);
nand U714 (N_714,N_518,N_427);
or U715 (N_715,N_427,N_477);
and U716 (N_716,N_584,N_557);
nand U717 (N_717,N_583,N_599);
nor U718 (N_718,N_543,N_479);
or U719 (N_719,N_495,N_408);
and U720 (N_720,N_406,N_544);
and U721 (N_721,N_584,N_425);
and U722 (N_722,N_460,N_480);
and U723 (N_723,N_568,N_597);
xnor U724 (N_724,N_409,N_442);
nand U725 (N_725,N_438,N_595);
and U726 (N_726,N_476,N_506);
nand U727 (N_727,N_460,N_583);
nor U728 (N_728,N_528,N_403);
or U729 (N_729,N_436,N_515);
nand U730 (N_730,N_484,N_460);
and U731 (N_731,N_565,N_571);
xor U732 (N_732,N_477,N_532);
and U733 (N_733,N_536,N_584);
or U734 (N_734,N_521,N_453);
nor U735 (N_735,N_544,N_402);
or U736 (N_736,N_556,N_460);
nor U737 (N_737,N_503,N_564);
nor U738 (N_738,N_557,N_429);
nor U739 (N_739,N_400,N_517);
or U740 (N_740,N_589,N_590);
nand U741 (N_741,N_414,N_447);
xor U742 (N_742,N_527,N_468);
or U743 (N_743,N_549,N_442);
or U744 (N_744,N_480,N_588);
nor U745 (N_745,N_595,N_416);
nand U746 (N_746,N_508,N_435);
xor U747 (N_747,N_475,N_513);
nand U748 (N_748,N_588,N_412);
nor U749 (N_749,N_523,N_502);
nor U750 (N_750,N_525,N_568);
nand U751 (N_751,N_431,N_453);
or U752 (N_752,N_407,N_419);
nor U753 (N_753,N_452,N_469);
nand U754 (N_754,N_577,N_475);
xnor U755 (N_755,N_420,N_458);
xor U756 (N_756,N_435,N_421);
and U757 (N_757,N_518,N_435);
xnor U758 (N_758,N_513,N_576);
and U759 (N_759,N_471,N_424);
and U760 (N_760,N_501,N_569);
or U761 (N_761,N_415,N_513);
nor U762 (N_762,N_407,N_469);
or U763 (N_763,N_473,N_422);
and U764 (N_764,N_404,N_432);
and U765 (N_765,N_581,N_449);
nor U766 (N_766,N_445,N_454);
and U767 (N_767,N_556,N_444);
nand U768 (N_768,N_530,N_490);
and U769 (N_769,N_438,N_579);
nand U770 (N_770,N_443,N_488);
or U771 (N_771,N_566,N_536);
xor U772 (N_772,N_574,N_530);
and U773 (N_773,N_434,N_529);
nor U774 (N_774,N_476,N_503);
nor U775 (N_775,N_450,N_510);
xor U776 (N_776,N_448,N_416);
xor U777 (N_777,N_408,N_574);
nor U778 (N_778,N_460,N_591);
and U779 (N_779,N_474,N_553);
nor U780 (N_780,N_585,N_557);
nand U781 (N_781,N_408,N_597);
xor U782 (N_782,N_403,N_473);
xor U783 (N_783,N_525,N_420);
nand U784 (N_784,N_538,N_577);
nand U785 (N_785,N_525,N_576);
and U786 (N_786,N_534,N_511);
nor U787 (N_787,N_506,N_488);
xor U788 (N_788,N_564,N_568);
nor U789 (N_789,N_512,N_416);
and U790 (N_790,N_436,N_510);
or U791 (N_791,N_468,N_448);
xor U792 (N_792,N_425,N_563);
or U793 (N_793,N_559,N_423);
and U794 (N_794,N_405,N_485);
and U795 (N_795,N_423,N_442);
nand U796 (N_796,N_432,N_454);
and U797 (N_797,N_509,N_559);
xor U798 (N_798,N_597,N_595);
nor U799 (N_799,N_454,N_563);
xnor U800 (N_800,N_700,N_722);
xnor U801 (N_801,N_713,N_690);
or U802 (N_802,N_710,N_738);
xnor U803 (N_803,N_782,N_624);
and U804 (N_804,N_795,N_612);
and U805 (N_805,N_625,N_770);
or U806 (N_806,N_608,N_666);
and U807 (N_807,N_771,N_615);
nand U808 (N_808,N_658,N_619);
nand U809 (N_809,N_693,N_662);
and U810 (N_810,N_628,N_652);
xnor U811 (N_811,N_670,N_725);
nor U812 (N_812,N_749,N_671);
nor U813 (N_813,N_681,N_794);
and U814 (N_814,N_702,N_616);
nand U815 (N_815,N_614,N_633);
nand U816 (N_816,N_783,N_793);
or U817 (N_817,N_768,N_760);
xnor U818 (N_818,N_689,N_778);
nor U819 (N_819,N_630,N_642);
nor U820 (N_820,N_779,N_692);
and U821 (N_821,N_684,N_744);
nor U822 (N_822,N_661,N_601);
xor U823 (N_823,N_660,N_635);
or U824 (N_824,N_643,N_672);
nor U825 (N_825,N_712,N_758);
xnor U826 (N_826,N_640,N_679);
nor U827 (N_827,N_664,N_605);
and U828 (N_828,N_634,N_762);
nand U829 (N_829,N_618,N_764);
and U830 (N_830,N_776,N_704);
or U831 (N_831,N_791,N_723);
xor U832 (N_832,N_638,N_650);
and U833 (N_833,N_604,N_737);
or U834 (N_834,N_680,N_743);
nand U835 (N_835,N_626,N_765);
xor U836 (N_836,N_777,N_766);
and U837 (N_837,N_657,N_789);
or U838 (N_838,N_707,N_715);
or U839 (N_839,N_622,N_687);
nor U840 (N_840,N_655,N_609);
and U841 (N_841,N_798,N_703);
xor U842 (N_842,N_797,N_726);
xor U843 (N_843,N_620,N_659);
nand U844 (N_844,N_646,N_675);
xnor U845 (N_845,N_735,N_781);
nand U846 (N_846,N_730,N_728);
or U847 (N_847,N_772,N_649);
nor U848 (N_848,N_756,N_716);
xor U849 (N_849,N_698,N_708);
nand U850 (N_850,N_603,N_641);
or U851 (N_851,N_740,N_632);
and U852 (N_852,N_606,N_688);
xnor U853 (N_853,N_623,N_668);
nor U854 (N_854,N_724,N_621);
and U855 (N_855,N_678,N_775);
or U856 (N_856,N_727,N_683);
nand U857 (N_857,N_645,N_750);
or U858 (N_858,N_602,N_709);
nor U859 (N_859,N_747,N_720);
or U860 (N_860,N_663,N_763);
and U861 (N_861,N_639,N_757);
nand U862 (N_862,N_733,N_685);
xnor U863 (N_863,N_706,N_651);
nor U864 (N_864,N_667,N_786);
xor U865 (N_865,N_755,N_711);
or U866 (N_866,N_769,N_617);
and U867 (N_867,N_673,N_686);
nand U868 (N_868,N_600,N_732);
or U869 (N_869,N_734,N_742);
or U870 (N_870,N_787,N_721);
and U871 (N_871,N_753,N_741);
or U872 (N_872,N_653,N_705);
and U873 (N_873,N_610,N_627);
xnor U874 (N_874,N_745,N_718);
xor U875 (N_875,N_607,N_746);
or U876 (N_876,N_774,N_648);
xor U877 (N_877,N_701,N_736);
and U878 (N_878,N_784,N_691);
and U879 (N_879,N_759,N_677);
xor U880 (N_880,N_796,N_761);
or U881 (N_881,N_799,N_697);
or U882 (N_882,N_731,N_682);
nand U883 (N_883,N_629,N_748);
and U884 (N_884,N_665,N_780);
nor U885 (N_885,N_767,N_695);
or U886 (N_886,N_719,N_773);
or U887 (N_887,N_611,N_792);
or U888 (N_888,N_656,N_788);
or U889 (N_889,N_696,N_647);
nor U890 (N_890,N_714,N_676);
nand U891 (N_891,N_637,N_694);
and U892 (N_892,N_739,N_644);
or U893 (N_893,N_785,N_674);
or U894 (N_894,N_754,N_654);
or U895 (N_895,N_717,N_790);
and U896 (N_896,N_699,N_751);
nand U897 (N_897,N_636,N_669);
nor U898 (N_898,N_752,N_613);
and U899 (N_899,N_631,N_729);
nand U900 (N_900,N_619,N_617);
or U901 (N_901,N_634,N_797);
xor U902 (N_902,N_674,N_746);
or U903 (N_903,N_684,N_680);
nor U904 (N_904,N_625,N_612);
nand U905 (N_905,N_716,N_612);
xor U906 (N_906,N_687,N_681);
or U907 (N_907,N_763,N_621);
and U908 (N_908,N_754,N_650);
or U909 (N_909,N_678,N_671);
and U910 (N_910,N_721,N_796);
xnor U911 (N_911,N_744,N_636);
or U912 (N_912,N_678,N_698);
and U913 (N_913,N_789,N_608);
xnor U914 (N_914,N_738,N_628);
nor U915 (N_915,N_604,N_664);
nand U916 (N_916,N_703,N_760);
and U917 (N_917,N_647,N_779);
or U918 (N_918,N_653,N_754);
and U919 (N_919,N_656,N_773);
nand U920 (N_920,N_613,N_709);
and U921 (N_921,N_799,N_761);
xnor U922 (N_922,N_799,N_603);
or U923 (N_923,N_732,N_698);
and U924 (N_924,N_741,N_625);
nor U925 (N_925,N_772,N_762);
xnor U926 (N_926,N_724,N_666);
xor U927 (N_927,N_648,N_668);
xnor U928 (N_928,N_786,N_604);
or U929 (N_929,N_739,N_712);
and U930 (N_930,N_786,N_697);
and U931 (N_931,N_734,N_652);
nand U932 (N_932,N_744,N_649);
and U933 (N_933,N_680,N_664);
and U934 (N_934,N_710,N_693);
or U935 (N_935,N_757,N_638);
or U936 (N_936,N_681,N_684);
or U937 (N_937,N_666,N_648);
nor U938 (N_938,N_698,N_692);
xnor U939 (N_939,N_656,N_655);
and U940 (N_940,N_780,N_674);
or U941 (N_941,N_770,N_775);
nand U942 (N_942,N_759,N_719);
and U943 (N_943,N_751,N_771);
or U944 (N_944,N_668,N_692);
nor U945 (N_945,N_754,N_755);
nand U946 (N_946,N_789,N_647);
and U947 (N_947,N_606,N_611);
and U948 (N_948,N_719,N_638);
xor U949 (N_949,N_770,N_606);
or U950 (N_950,N_789,N_656);
xnor U951 (N_951,N_647,N_649);
xor U952 (N_952,N_635,N_699);
or U953 (N_953,N_795,N_678);
and U954 (N_954,N_614,N_738);
or U955 (N_955,N_768,N_738);
xnor U956 (N_956,N_606,N_782);
and U957 (N_957,N_719,N_749);
nand U958 (N_958,N_784,N_797);
and U959 (N_959,N_675,N_795);
and U960 (N_960,N_692,N_751);
and U961 (N_961,N_783,N_747);
xnor U962 (N_962,N_781,N_616);
and U963 (N_963,N_663,N_624);
or U964 (N_964,N_660,N_701);
or U965 (N_965,N_633,N_677);
and U966 (N_966,N_669,N_763);
nand U967 (N_967,N_722,N_620);
and U968 (N_968,N_635,N_755);
xnor U969 (N_969,N_621,N_665);
and U970 (N_970,N_661,N_736);
and U971 (N_971,N_721,N_783);
nor U972 (N_972,N_657,N_751);
or U973 (N_973,N_651,N_636);
xnor U974 (N_974,N_760,N_690);
and U975 (N_975,N_793,N_651);
nor U976 (N_976,N_799,N_770);
xnor U977 (N_977,N_743,N_668);
nor U978 (N_978,N_695,N_734);
or U979 (N_979,N_656,N_670);
and U980 (N_980,N_604,N_776);
or U981 (N_981,N_796,N_689);
or U982 (N_982,N_650,N_709);
nand U983 (N_983,N_700,N_625);
or U984 (N_984,N_654,N_642);
nor U985 (N_985,N_705,N_620);
or U986 (N_986,N_654,N_669);
nand U987 (N_987,N_663,N_631);
nor U988 (N_988,N_772,N_783);
or U989 (N_989,N_655,N_727);
nor U990 (N_990,N_725,N_775);
and U991 (N_991,N_768,N_655);
or U992 (N_992,N_737,N_758);
nor U993 (N_993,N_783,N_690);
and U994 (N_994,N_731,N_646);
or U995 (N_995,N_707,N_615);
or U996 (N_996,N_707,N_794);
and U997 (N_997,N_756,N_793);
xnor U998 (N_998,N_677,N_628);
xnor U999 (N_999,N_792,N_778);
nand U1000 (N_1000,N_853,N_950);
or U1001 (N_1001,N_973,N_944);
nand U1002 (N_1002,N_889,N_834);
or U1003 (N_1003,N_811,N_959);
and U1004 (N_1004,N_979,N_879);
nor U1005 (N_1005,N_874,N_814);
xor U1006 (N_1006,N_887,N_808);
or U1007 (N_1007,N_957,N_929);
nand U1008 (N_1008,N_913,N_835);
nor U1009 (N_1009,N_988,N_820);
nand U1010 (N_1010,N_810,N_871);
and U1011 (N_1011,N_815,N_829);
xor U1012 (N_1012,N_948,N_843);
nor U1013 (N_1013,N_958,N_909);
nor U1014 (N_1014,N_809,N_857);
nand U1015 (N_1015,N_885,N_953);
nor U1016 (N_1016,N_895,N_920);
nor U1017 (N_1017,N_993,N_939);
and U1018 (N_1018,N_864,N_807);
or U1019 (N_1019,N_925,N_999);
xor U1020 (N_1020,N_892,N_947);
or U1021 (N_1021,N_990,N_997);
nor U1022 (N_1022,N_926,N_801);
or U1023 (N_1023,N_960,N_832);
nand U1024 (N_1024,N_823,N_995);
and U1025 (N_1025,N_983,N_934);
nor U1026 (N_1026,N_986,N_932);
nand U1027 (N_1027,N_850,N_949);
xnor U1028 (N_1028,N_846,N_851);
xor U1029 (N_1029,N_908,N_922);
or U1030 (N_1030,N_977,N_968);
nand U1031 (N_1031,N_903,N_992);
and U1032 (N_1032,N_854,N_927);
nor U1033 (N_1033,N_804,N_981);
or U1034 (N_1034,N_896,N_802);
xor U1035 (N_1035,N_914,N_978);
or U1036 (N_1036,N_898,N_826);
nor U1037 (N_1037,N_862,N_942);
xor U1038 (N_1038,N_985,N_901);
nor U1039 (N_1039,N_856,N_890);
xnor U1040 (N_1040,N_906,N_848);
or U1041 (N_1041,N_975,N_845);
and U1042 (N_1042,N_886,N_930);
or U1043 (N_1043,N_900,N_858);
nor U1044 (N_1044,N_855,N_964);
and U1045 (N_1045,N_951,N_924);
nand U1046 (N_1046,N_928,N_989);
or U1047 (N_1047,N_915,N_937);
or U1048 (N_1048,N_970,N_963);
nand U1049 (N_1049,N_994,N_805);
and U1050 (N_1050,N_881,N_821);
nand U1051 (N_1051,N_863,N_876);
nor U1052 (N_1052,N_800,N_847);
xnor U1053 (N_1053,N_984,N_865);
or U1054 (N_1054,N_936,N_987);
nand U1055 (N_1055,N_955,N_921);
nand U1056 (N_1056,N_910,N_962);
nand U1057 (N_1057,N_916,N_803);
and U1058 (N_1058,N_869,N_833);
or U1059 (N_1059,N_891,N_917);
xnor U1060 (N_1060,N_961,N_836);
nand U1061 (N_1061,N_972,N_806);
and U1062 (N_1062,N_897,N_827);
and U1063 (N_1063,N_911,N_974);
and U1064 (N_1064,N_861,N_952);
or U1065 (N_1065,N_888,N_816);
nand U1066 (N_1066,N_971,N_966);
nor U1067 (N_1067,N_867,N_842);
or U1068 (N_1068,N_894,N_980);
or U1069 (N_1069,N_938,N_840);
nand U1070 (N_1070,N_996,N_813);
nand U1071 (N_1071,N_872,N_878);
or U1072 (N_1072,N_945,N_976);
or U1073 (N_1073,N_965,N_969);
xnor U1074 (N_1074,N_893,N_839);
xor U1075 (N_1075,N_883,N_991);
nand U1076 (N_1076,N_902,N_852);
or U1077 (N_1077,N_812,N_825);
xnor U1078 (N_1078,N_873,N_982);
nand U1079 (N_1079,N_941,N_828);
nor U1080 (N_1080,N_899,N_919);
and U1081 (N_1081,N_956,N_912);
nor U1082 (N_1082,N_849,N_877);
nand U1083 (N_1083,N_904,N_933);
nor U1084 (N_1084,N_817,N_837);
nor U1085 (N_1085,N_931,N_824);
or U1086 (N_1086,N_859,N_940);
nand U1087 (N_1087,N_830,N_943);
xnor U1088 (N_1088,N_875,N_918);
or U1089 (N_1089,N_954,N_870);
and U1090 (N_1090,N_907,N_882);
xnor U1091 (N_1091,N_841,N_868);
nand U1092 (N_1092,N_905,N_838);
nor U1093 (N_1093,N_866,N_946);
nor U1094 (N_1094,N_818,N_935);
nand U1095 (N_1095,N_844,N_831);
xnor U1096 (N_1096,N_880,N_923);
nand U1097 (N_1097,N_998,N_822);
and U1098 (N_1098,N_884,N_967);
xor U1099 (N_1099,N_860,N_819);
or U1100 (N_1100,N_988,N_999);
and U1101 (N_1101,N_854,N_902);
xor U1102 (N_1102,N_967,N_825);
or U1103 (N_1103,N_883,N_834);
and U1104 (N_1104,N_932,N_893);
xnor U1105 (N_1105,N_982,N_892);
nor U1106 (N_1106,N_930,N_973);
xor U1107 (N_1107,N_810,N_850);
xnor U1108 (N_1108,N_863,N_850);
nor U1109 (N_1109,N_895,N_877);
xnor U1110 (N_1110,N_866,N_807);
or U1111 (N_1111,N_978,N_908);
xor U1112 (N_1112,N_979,N_986);
xnor U1113 (N_1113,N_829,N_888);
xor U1114 (N_1114,N_904,N_876);
or U1115 (N_1115,N_968,N_862);
xnor U1116 (N_1116,N_807,N_954);
nand U1117 (N_1117,N_980,N_889);
xnor U1118 (N_1118,N_964,N_982);
xnor U1119 (N_1119,N_976,N_891);
and U1120 (N_1120,N_924,N_831);
nor U1121 (N_1121,N_964,N_816);
xnor U1122 (N_1122,N_969,N_935);
xnor U1123 (N_1123,N_998,N_905);
xnor U1124 (N_1124,N_871,N_982);
and U1125 (N_1125,N_970,N_853);
xor U1126 (N_1126,N_802,N_817);
nor U1127 (N_1127,N_920,N_988);
and U1128 (N_1128,N_977,N_806);
and U1129 (N_1129,N_849,N_875);
or U1130 (N_1130,N_939,N_931);
nor U1131 (N_1131,N_899,N_833);
or U1132 (N_1132,N_808,N_967);
or U1133 (N_1133,N_876,N_844);
nand U1134 (N_1134,N_983,N_832);
and U1135 (N_1135,N_840,N_935);
xor U1136 (N_1136,N_995,N_831);
nand U1137 (N_1137,N_843,N_981);
nor U1138 (N_1138,N_848,N_945);
nor U1139 (N_1139,N_879,N_973);
nor U1140 (N_1140,N_816,N_880);
or U1141 (N_1141,N_934,N_974);
nand U1142 (N_1142,N_858,N_926);
xnor U1143 (N_1143,N_861,N_972);
or U1144 (N_1144,N_904,N_816);
and U1145 (N_1145,N_822,N_973);
nand U1146 (N_1146,N_851,N_952);
xnor U1147 (N_1147,N_988,N_828);
xor U1148 (N_1148,N_865,N_810);
and U1149 (N_1149,N_848,N_970);
or U1150 (N_1150,N_818,N_952);
and U1151 (N_1151,N_836,N_862);
nand U1152 (N_1152,N_817,N_863);
nor U1153 (N_1153,N_875,N_903);
or U1154 (N_1154,N_959,N_852);
and U1155 (N_1155,N_972,N_894);
nor U1156 (N_1156,N_855,N_941);
xor U1157 (N_1157,N_879,N_900);
xor U1158 (N_1158,N_984,N_816);
or U1159 (N_1159,N_859,N_950);
xor U1160 (N_1160,N_808,N_954);
and U1161 (N_1161,N_922,N_946);
nor U1162 (N_1162,N_815,N_835);
nor U1163 (N_1163,N_857,N_946);
and U1164 (N_1164,N_820,N_855);
nand U1165 (N_1165,N_864,N_919);
nor U1166 (N_1166,N_953,N_849);
nand U1167 (N_1167,N_910,N_842);
nand U1168 (N_1168,N_871,N_949);
or U1169 (N_1169,N_811,N_858);
nor U1170 (N_1170,N_931,N_838);
or U1171 (N_1171,N_816,N_882);
and U1172 (N_1172,N_861,N_857);
xor U1173 (N_1173,N_951,N_906);
and U1174 (N_1174,N_990,N_870);
and U1175 (N_1175,N_995,N_909);
nand U1176 (N_1176,N_920,N_852);
nand U1177 (N_1177,N_995,N_841);
xor U1178 (N_1178,N_979,N_981);
nor U1179 (N_1179,N_850,N_852);
nand U1180 (N_1180,N_878,N_882);
nand U1181 (N_1181,N_957,N_971);
xnor U1182 (N_1182,N_856,N_808);
xor U1183 (N_1183,N_841,N_942);
and U1184 (N_1184,N_833,N_935);
nor U1185 (N_1185,N_861,N_968);
nand U1186 (N_1186,N_969,N_954);
nand U1187 (N_1187,N_814,N_869);
and U1188 (N_1188,N_851,N_972);
nand U1189 (N_1189,N_915,N_928);
nor U1190 (N_1190,N_951,N_936);
xor U1191 (N_1191,N_826,N_905);
nand U1192 (N_1192,N_822,N_922);
nand U1193 (N_1193,N_848,N_887);
or U1194 (N_1194,N_909,N_978);
xor U1195 (N_1195,N_957,N_961);
and U1196 (N_1196,N_805,N_961);
or U1197 (N_1197,N_865,N_992);
nor U1198 (N_1198,N_859,N_815);
and U1199 (N_1199,N_807,N_955);
nand U1200 (N_1200,N_1041,N_1163);
nand U1201 (N_1201,N_1122,N_1119);
nand U1202 (N_1202,N_1042,N_1088);
and U1203 (N_1203,N_1120,N_1174);
nor U1204 (N_1204,N_1072,N_1144);
nor U1205 (N_1205,N_1195,N_1092);
and U1206 (N_1206,N_1115,N_1138);
or U1207 (N_1207,N_1027,N_1155);
xor U1208 (N_1208,N_1007,N_1015);
nand U1209 (N_1209,N_1183,N_1018);
xor U1210 (N_1210,N_1097,N_1020);
nand U1211 (N_1211,N_1182,N_1019);
xor U1212 (N_1212,N_1188,N_1178);
xor U1213 (N_1213,N_1171,N_1137);
nor U1214 (N_1214,N_1085,N_1108);
nand U1215 (N_1215,N_1073,N_1008);
nand U1216 (N_1216,N_1118,N_1051);
and U1217 (N_1217,N_1135,N_1198);
nand U1218 (N_1218,N_1117,N_1165);
and U1219 (N_1219,N_1169,N_1002);
xnor U1220 (N_1220,N_1030,N_1040);
nand U1221 (N_1221,N_1162,N_1159);
xor U1222 (N_1222,N_1187,N_1111);
and U1223 (N_1223,N_1047,N_1114);
nand U1224 (N_1224,N_1185,N_1134);
or U1225 (N_1225,N_1140,N_1036);
and U1226 (N_1226,N_1069,N_1121);
nor U1227 (N_1227,N_1065,N_1062);
and U1228 (N_1228,N_1035,N_1012);
nand U1229 (N_1229,N_1013,N_1161);
nor U1230 (N_1230,N_1074,N_1031);
or U1231 (N_1231,N_1017,N_1184);
nor U1232 (N_1232,N_1133,N_1179);
nand U1233 (N_1233,N_1004,N_1034);
nor U1234 (N_1234,N_1175,N_1166);
nand U1235 (N_1235,N_1089,N_1023);
xor U1236 (N_1236,N_1146,N_1000);
xor U1237 (N_1237,N_1100,N_1176);
nor U1238 (N_1238,N_1164,N_1186);
and U1239 (N_1239,N_1087,N_1160);
nand U1240 (N_1240,N_1196,N_1126);
and U1241 (N_1241,N_1049,N_1099);
and U1242 (N_1242,N_1180,N_1125);
nor U1243 (N_1243,N_1081,N_1001);
or U1244 (N_1244,N_1197,N_1014);
or U1245 (N_1245,N_1045,N_1039);
xnor U1246 (N_1246,N_1044,N_1091);
nor U1247 (N_1247,N_1066,N_1123);
or U1248 (N_1248,N_1101,N_1032);
and U1249 (N_1249,N_1006,N_1070);
or U1250 (N_1250,N_1055,N_1068);
xor U1251 (N_1251,N_1151,N_1060);
nand U1252 (N_1252,N_1177,N_1168);
xor U1253 (N_1253,N_1113,N_1154);
nand U1254 (N_1254,N_1152,N_1105);
nor U1255 (N_1255,N_1142,N_1024);
nor U1256 (N_1256,N_1116,N_1064);
nand U1257 (N_1257,N_1199,N_1038);
or U1258 (N_1258,N_1128,N_1153);
xor U1259 (N_1259,N_1094,N_1079);
or U1260 (N_1260,N_1033,N_1080);
nand U1261 (N_1261,N_1127,N_1095);
nor U1262 (N_1262,N_1191,N_1090);
nor U1263 (N_1263,N_1011,N_1147);
nand U1264 (N_1264,N_1173,N_1054);
xnor U1265 (N_1265,N_1037,N_1167);
xor U1266 (N_1266,N_1110,N_1086);
or U1267 (N_1267,N_1193,N_1124);
xor U1268 (N_1268,N_1084,N_1046);
xnor U1269 (N_1269,N_1053,N_1192);
nor U1270 (N_1270,N_1003,N_1052);
xor U1271 (N_1271,N_1028,N_1139);
xor U1272 (N_1272,N_1129,N_1063);
nor U1273 (N_1273,N_1157,N_1083);
xor U1274 (N_1274,N_1043,N_1130);
or U1275 (N_1275,N_1098,N_1061);
nand U1276 (N_1276,N_1056,N_1093);
and U1277 (N_1277,N_1009,N_1131);
or U1278 (N_1278,N_1194,N_1029);
nand U1279 (N_1279,N_1025,N_1158);
nand U1280 (N_1280,N_1143,N_1050);
xnor U1281 (N_1281,N_1071,N_1096);
nor U1282 (N_1282,N_1048,N_1170);
xor U1283 (N_1283,N_1109,N_1102);
xor U1284 (N_1284,N_1067,N_1106);
nor U1285 (N_1285,N_1059,N_1150);
nand U1286 (N_1286,N_1104,N_1057);
and U1287 (N_1287,N_1112,N_1077);
or U1288 (N_1288,N_1005,N_1107);
nand U1289 (N_1289,N_1149,N_1026);
xor U1290 (N_1290,N_1058,N_1189);
nand U1291 (N_1291,N_1181,N_1010);
and U1292 (N_1292,N_1172,N_1148);
or U1293 (N_1293,N_1078,N_1132);
xor U1294 (N_1294,N_1075,N_1141);
and U1295 (N_1295,N_1145,N_1103);
nand U1296 (N_1296,N_1156,N_1021);
and U1297 (N_1297,N_1016,N_1076);
and U1298 (N_1298,N_1022,N_1082);
xor U1299 (N_1299,N_1190,N_1136);
xor U1300 (N_1300,N_1162,N_1043);
nor U1301 (N_1301,N_1083,N_1128);
or U1302 (N_1302,N_1104,N_1086);
and U1303 (N_1303,N_1039,N_1072);
and U1304 (N_1304,N_1004,N_1006);
xnor U1305 (N_1305,N_1106,N_1190);
nand U1306 (N_1306,N_1060,N_1125);
nand U1307 (N_1307,N_1148,N_1161);
and U1308 (N_1308,N_1146,N_1083);
or U1309 (N_1309,N_1025,N_1172);
nand U1310 (N_1310,N_1027,N_1030);
nand U1311 (N_1311,N_1168,N_1151);
and U1312 (N_1312,N_1075,N_1104);
nand U1313 (N_1313,N_1100,N_1128);
nand U1314 (N_1314,N_1185,N_1079);
nor U1315 (N_1315,N_1116,N_1078);
and U1316 (N_1316,N_1098,N_1106);
nand U1317 (N_1317,N_1182,N_1111);
and U1318 (N_1318,N_1164,N_1025);
nor U1319 (N_1319,N_1072,N_1014);
xor U1320 (N_1320,N_1159,N_1004);
or U1321 (N_1321,N_1010,N_1191);
xor U1322 (N_1322,N_1111,N_1064);
xnor U1323 (N_1323,N_1116,N_1018);
xnor U1324 (N_1324,N_1105,N_1007);
nand U1325 (N_1325,N_1142,N_1135);
nor U1326 (N_1326,N_1119,N_1161);
nor U1327 (N_1327,N_1063,N_1037);
xor U1328 (N_1328,N_1106,N_1006);
xor U1329 (N_1329,N_1184,N_1046);
or U1330 (N_1330,N_1013,N_1061);
xor U1331 (N_1331,N_1140,N_1069);
and U1332 (N_1332,N_1137,N_1097);
nand U1333 (N_1333,N_1007,N_1058);
and U1334 (N_1334,N_1186,N_1085);
and U1335 (N_1335,N_1000,N_1013);
nor U1336 (N_1336,N_1155,N_1039);
nand U1337 (N_1337,N_1091,N_1169);
xor U1338 (N_1338,N_1190,N_1112);
and U1339 (N_1339,N_1053,N_1165);
and U1340 (N_1340,N_1086,N_1088);
nand U1341 (N_1341,N_1137,N_1183);
and U1342 (N_1342,N_1039,N_1180);
nand U1343 (N_1343,N_1157,N_1044);
or U1344 (N_1344,N_1194,N_1112);
xnor U1345 (N_1345,N_1190,N_1022);
nand U1346 (N_1346,N_1003,N_1169);
xnor U1347 (N_1347,N_1172,N_1084);
or U1348 (N_1348,N_1062,N_1171);
and U1349 (N_1349,N_1153,N_1193);
nand U1350 (N_1350,N_1045,N_1116);
and U1351 (N_1351,N_1077,N_1116);
xor U1352 (N_1352,N_1042,N_1071);
xor U1353 (N_1353,N_1125,N_1052);
nor U1354 (N_1354,N_1132,N_1094);
and U1355 (N_1355,N_1153,N_1124);
and U1356 (N_1356,N_1177,N_1071);
nand U1357 (N_1357,N_1193,N_1004);
nor U1358 (N_1358,N_1018,N_1050);
and U1359 (N_1359,N_1017,N_1100);
xor U1360 (N_1360,N_1139,N_1008);
and U1361 (N_1361,N_1034,N_1188);
nand U1362 (N_1362,N_1108,N_1115);
xor U1363 (N_1363,N_1154,N_1132);
or U1364 (N_1364,N_1168,N_1122);
xnor U1365 (N_1365,N_1048,N_1033);
nand U1366 (N_1366,N_1155,N_1175);
nor U1367 (N_1367,N_1032,N_1120);
nor U1368 (N_1368,N_1003,N_1175);
nand U1369 (N_1369,N_1181,N_1073);
xor U1370 (N_1370,N_1019,N_1086);
nand U1371 (N_1371,N_1122,N_1191);
nor U1372 (N_1372,N_1062,N_1059);
nor U1373 (N_1373,N_1131,N_1052);
and U1374 (N_1374,N_1072,N_1075);
nand U1375 (N_1375,N_1147,N_1135);
and U1376 (N_1376,N_1023,N_1111);
xor U1377 (N_1377,N_1166,N_1140);
xnor U1378 (N_1378,N_1137,N_1136);
or U1379 (N_1379,N_1176,N_1067);
or U1380 (N_1380,N_1075,N_1087);
nand U1381 (N_1381,N_1026,N_1071);
xnor U1382 (N_1382,N_1025,N_1092);
xnor U1383 (N_1383,N_1035,N_1175);
nand U1384 (N_1384,N_1192,N_1066);
xnor U1385 (N_1385,N_1166,N_1056);
xnor U1386 (N_1386,N_1144,N_1098);
xor U1387 (N_1387,N_1099,N_1004);
or U1388 (N_1388,N_1057,N_1071);
and U1389 (N_1389,N_1097,N_1152);
or U1390 (N_1390,N_1050,N_1084);
nand U1391 (N_1391,N_1188,N_1033);
and U1392 (N_1392,N_1166,N_1180);
and U1393 (N_1393,N_1020,N_1100);
or U1394 (N_1394,N_1146,N_1067);
and U1395 (N_1395,N_1072,N_1089);
or U1396 (N_1396,N_1034,N_1111);
xnor U1397 (N_1397,N_1087,N_1124);
or U1398 (N_1398,N_1187,N_1077);
or U1399 (N_1399,N_1038,N_1132);
nand U1400 (N_1400,N_1244,N_1386);
or U1401 (N_1401,N_1306,N_1269);
nor U1402 (N_1402,N_1224,N_1257);
nand U1403 (N_1403,N_1211,N_1264);
and U1404 (N_1404,N_1240,N_1307);
nor U1405 (N_1405,N_1382,N_1258);
nand U1406 (N_1406,N_1204,N_1241);
or U1407 (N_1407,N_1349,N_1256);
and U1408 (N_1408,N_1337,N_1252);
or U1409 (N_1409,N_1330,N_1321);
xor U1410 (N_1410,N_1215,N_1304);
nand U1411 (N_1411,N_1281,N_1276);
and U1412 (N_1412,N_1296,N_1372);
or U1413 (N_1413,N_1203,N_1270);
and U1414 (N_1414,N_1353,N_1345);
and U1415 (N_1415,N_1294,N_1359);
and U1416 (N_1416,N_1213,N_1314);
nor U1417 (N_1417,N_1229,N_1318);
nand U1418 (N_1418,N_1380,N_1346);
and U1419 (N_1419,N_1259,N_1384);
or U1420 (N_1420,N_1357,N_1338);
nand U1421 (N_1421,N_1396,N_1378);
or U1422 (N_1422,N_1363,N_1394);
nor U1423 (N_1423,N_1320,N_1327);
and U1424 (N_1424,N_1398,N_1260);
nand U1425 (N_1425,N_1308,N_1201);
nor U1426 (N_1426,N_1280,N_1364);
or U1427 (N_1427,N_1356,N_1212);
nor U1428 (N_1428,N_1319,N_1388);
nand U1429 (N_1429,N_1354,N_1262);
and U1430 (N_1430,N_1350,N_1347);
xnor U1431 (N_1431,N_1342,N_1253);
and U1432 (N_1432,N_1208,N_1210);
or U1433 (N_1433,N_1236,N_1218);
and U1434 (N_1434,N_1376,N_1272);
and U1435 (N_1435,N_1290,N_1329);
or U1436 (N_1436,N_1383,N_1371);
nand U1437 (N_1437,N_1341,N_1309);
and U1438 (N_1438,N_1232,N_1374);
xor U1439 (N_1439,N_1362,N_1324);
nand U1440 (N_1440,N_1302,N_1243);
nand U1441 (N_1441,N_1255,N_1273);
nand U1442 (N_1442,N_1246,N_1300);
and U1443 (N_1443,N_1293,N_1251);
nand U1444 (N_1444,N_1310,N_1322);
or U1445 (N_1445,N_1340,N_1331);
and U1446 (N_1446,N_1265,N_1266);
xnor U1447 (N_1447,N_1222,N_1344);
nand U1448 (N_1448,N_1263,N_1209);
nor U1449 (N_1449,N_1361,N_1312);
or U1450 (N_1450,N_1235,N_1288);
or U1451 (N_1451,N_1242,N_1278);
and U1452 (N_1452,N_1261,N_1219);
xnor U1453 (N_1453,N_1275,N_1231);
nand U1454 (N_1454,N_1200,N_1392);
xnor U1455 (N_1455,N_1247,N_1207);
and U1456 (N_1456,N_1360,N_1387);
and U1457 (N_1457,N_1289,N_1271);
nand U1458 (N_1458,N_1390,N_1305);
xnor U1459 (N_1459,N_1325,N_1279);
and U1460 (N_1460,N_1220,N_1355);
or U1461 (N_1461,N_1333,N_1223);
or U1462 (N_1462,N_1370,N_1336);
xor U1463 (N_1463,N_1348,N_1326);
xnor U1464 (N_1464,N_1217,N_1381);
nand U1465 (N_1465,N_1313,N_1214);
or U1466 (N_1466,N_1238,N_1254);
and U1467 (N_1467,N_1316,N_1366);
or U1468 (N_1468,N_1205,N_1297);
or U1469 (N_1469,N_1369,N_1389);
nor U1470 (N_1470,N_1239,N_1267);
nor U1471 (N_1471,N_1303,N_1277);
and U1472 (N_1472,N_1311,N_1301);
and U1473 (N_1473,N_1295,N_1317);
nor U1474 (N_1474,N_1284,N_1227);
nor U1475 (N_1475,N_1237,N_1202);
nand U1476 (N_1476,N_1352,N_1282);
nor U1477 (N_1477,N_1339,N_1323);
nand U1478 (N_1478,N_1233,N_1358);
nor U1479 (N_1479,N_1385,N_1245);
nor U1480 (N_1480,N_1332,N_1397);
nor U1481 (N_1481,N_1268,N_1248);
nor U1482 (N_1482,N_1286,N_1221);
and U1483 (N_1483,N_1249,N_1393);
nor U1484 (N_1484,N_1334,N_1287);
or U1485 (N_1485,N_1299,N_1226);
or U1486 (N_1486,N_1368,N_1367);
or U1487 (N_1487,N_1228,N_1216);
xor U1488 (N_1488,N_1351,N_1230);
nand U1489 (N_1489,N_1298,N_1377);
xnor U1490 (N_1490,N_1379,N_1283);
xor U1491 (N_1491,N_1274,N_1375);
nand U1492 (N_1492,N_1343,N_1234);
and U1493 (N_1493,N_1391,N_1365);
or U1494 (N_1494,N_1395,N_1285);
xor U1495 (N_1495,N_1399,N_1328);
or U1496 (N_1496,N_1315,N_1291);
nand U1497 (N_1497,N_1373,N_1250);
or U1498 (N_1498,N_1225,N_1335);
nand U1499 (N_1499,N_1206,N_1292);
or U1500 (N_1500,N_1376,N_1303);
or U1501 (N_1501,N_1236,N_1228);
and U1502 (N_1502,N_1372,N_1381);
nand U1503 (N_1503,N_1288,N_1345);
nor U1504 (N_1504,N_1294,N_1218);
nor U1505 (N_1505,N_1286,N_1300);
nor U1506 (N_1506,N_1397,N_1227);
nand U1507 (N_1507,N_1290,N_1297);
and U1508 (N_1508,N_1282,N_1346);
or U1509 (N_1509,N_1356,N_1288);
nor U1510 (N_1510,N_1225,N_1390);
nand U1511 (N_1511,N_1332,N_1392);
nor U1512 (N_1512,N_1286,N_1380);
nand U1513 (N_1513,N_1247,N_1327);
xor U1514 (N_1514,N_1379,N_1214);
or U1515 (N_1515,N_1201,N_1334);
and U1516 (N_1516,N_1367,N_1232);
nor U1517 (N_1517,N_1325,N_1222);
and U1518 (N_1518,N_1337,N_1367);
nand U1519 (N_1519,N_1249,N_1278);
nand U1520 (N_1520,N_1323,N_1279);
or U1521 (N_1521,N_1237,N_1397);
nand U1522 (N_1522,N_1249,N_1329);
nand U1523 (N_1523,N_1226,N_1285);
or U1524 (N_1524,N_1200,N_1282);
nand U1525 (N_1525,N_1313,N_1275);
nor U1526 (N_1526,N_1254,N_1376);
xnor U1527 (N_1527,N_1377,N_1205);
or U1528 (N_1528,N_1366,N_1238);
and U1529 (N_1529,N_1305,N_1274);
or U1530 (N_1530,N_1362,N_1213);
xor U1531 (N_1531,N_1310,N_1397);
or U1532 (N_1532,N_1235,N_1301);
nand U1533 (N_1533,N_1340,N_1253);
and U1534 (N_1534,N_1296,N_1312);
and U1535 (N_1535,N_1305,N_1356);
xor U1536 (N_1536,N_1332,N_1221);
and U1537 (N_1537,N_1249,N_1335);
or U1538 (N_1538,N_1250,N_1388);
and U1539 (N_1539,N_1385,N_1359);
nor U1540 (N_1540,N_1356,N_1294);
nor U1541 (N_1541,N_1249,N_1377);
nand U1542 (N_1542,N_1319,N_1249);
xnor U1543 (N_1543,N_1362,N_1387);
nor U1544 (N_1544,N_1390,N_1361);
and U1545 (N_1545,N_1351,N_1237);
nand U1546 (N_1546,N_1343,N_1303);
or U1547 (N_1547,N_1261,N_1260);
xor U1548 (N_1548,N_1371,N_1392);
nand U1549 (N_1549,N_1370,N_1387);
xor U1550 (N_1550,N_1322,N_1245);
or U1551 (N_1551,N_1203,N_1288);
xnor U1552 (N_1552,N_1360,N_1349);
or U1553 (N_1553,N_1370,N_1341);
nand U1554 (N_1554,N_1235,N_1335);
nand U1555 (N_1555,N_1240,N_1301);
nand U1556 (N_1556,N_1326,N_1365);
or U1557 (N_1557,N_1280,N_1243);
and U1558 (N_1558,N_1382,N_1215);
nor U1559 (N_1559,N_1374,N_1224);
nor U1560 (N_1560,N_1244,N_1298);
xor U1561 (N_1561,N_1398,N_1293);
nand U1562 (N_1562,N_1259,N_1215);
nor U1563 (N_1563,N_1396,N_1399);
nand U1564 (N_1564,N_1235,N_1343);
xnor U1565 (N_1565,N_1316,N_1326);
nand U1566 (N_1566,N_1335,N_1308);
and U1567 (N_1567,N_1322,N_1209);
nor U1568 (N_1568,N_1304,N_1296);
or U1569 (N_1569,N_1332,N_1320);
or U1570 (N_1570,N_1245,N_1234);
and U1571 (N_1571,N_1370,N_1292);
xor U1572 (N_1572,N_1214,N_1261);
nand U1573 (N_1573,N_1258,N_1233);
nor U1574 (N_1574,N_1339,N_1395);
nand U1575 (N_1575,N_1250,N_1344);
nand U1576 (N_1576,N_1291,N_1283);
nand U1577 (N_1577,N_1221,N_1344);
xnor U1578 (N_1578,N_1357,N_1392);
xnor U1579 (N_1579,N_1371,N_1361);
nor U1580 (N_1580,N_1381,N_1298);
and U1581 (N_1581,N_1281,N_1202);
xor U1582 (N_1582,N_1241,N_1318);
xor U1583 (N_1583,N_1267,N_1316);
and U1584 (N_1584,N_1399,N_1355);
or U1585 (N_1585,N_1383,N_1261);
and U1586 (N_1586,N_1208,N_1340);
xnor U1587 (N_1587,N_1317,N_1229);
nand U1588 (N_1588,N_1289,N_1226);
or U1589 (N_1589,N_1280,N_1354);
nand U1590 (N_1590,N_1246,N_1303);
and U1591 (N_1591,N_1228,N_1342);
nand U1592 (N_1592,N_1264,N_1297);
nor U1593 (N_1593,N_1289,N_1263);
xor U1594 (N_1594,N_1252,N_1304);
or U1595 (N_1595,N_1241,N_1348);
nor U1596 (N_1596,N_1289,N_1288);
or U1597 (N_1597,N_1231,N_1246);
xor U1598 (N_1598,N_1204,N_1225);
or U1599 (N_1599,N_1225,N_1243);
or U1600 (N_1600,N_1513,N_1543);
and U1601 (N_1601,N_1438,N_1554);
and U1602 (N_1602,N_1528,N_1464);
nor U1603 (N_1603,N_1485,N_1500);
nand U1604 (N_1604,N_1588,N_1442);
nor U1605 (N_1605,N_1467,N_1561);
nor U1606 (N_1606,N_1558,N_1576);
nor U1607 (N_1607,N_1466,N_1566);
or U1608 (N_1608,N_1518,N_1544);
xnor U1609 (N_1609,N_1538,N_1510);
nand U1610 (N_1610,N_1534,N_1560);
and U1611 (N_1611,N_1497,N_1527);
or U1612 (N_1612,N_1526,N_1409);
or U1613 (N_1613,N_1580,N_1480);
xnor U1614 (N_1614,N_1489,N_1508);
and U1615 (N_1615,N_1476,N_1559);
and U1616 (N_1616,N_1516,N_1515);
xnor U1617 (N_1617,N_1540,N_1475);
or U1618 (N_1618,N_1573,N_1551);
or U1619 (N_1619,N_1595,N_1571);
xor U1620 (N_1620,N_1450,N_1522);
nand U1621 (N_1621,N_1530,N_1499);
or U1622 (N_1622,N_1448,N_1597);
or U1623 (N_1623,N_1536,N_1470);
xnor U1624 (N_1624,N_1550,N_1401);
and U1625 (N_1625,N_1492,N_1445);
nand U1626 (N_1626,N_1491,N_1407);
xnor U1627 (N_1627,N_1494,N_1549);
nand U1628 (N_1628,N_1472,N_1574);
nor U1629 (N_1629,N_1565,N_1598);
or U1630 (N_1630,N_1456,N_1596);
nand U1631 (N_1631,N_1408,N_1562);
nor U1632 (N_1632,N_1542,N_1557);
nand U1633 (N_1633,N_1463,N_1507);
nand U1634 (N_1634,N_1412,N_1582);
nor U1635 (N_1635,N_1457,N_1462);
nand U1636 (N_1636,N_1553,N_1414);
nand U1637 (N_1637,N_1477,N_1441);
nor U1638 (N_1638,N_1584,N_1465);
nor U1639 (N_1639,N_1493,N_1535);
nand U1640 (N_1640,N_1583,N_1437);
and U1641 (N_1641,N_1577,N_1403);
and U1642 (N_1642,N_1454,N_1433);
or U1643 (N_1643,N_1453,N_1423);
and U1644 (N_1644,N_1451,N_1478);
or U1645 (N_1645,N_1434,N_1468);
or U1646 (N_1646,N_1599,N_1531);
and U1647 (N_1647,N_1420,N_1427);
xor U1648 (N_1648,N_1479,N_1471);
and U1649 (N_1649,N_1504,N_1490);
nor U1650 (N_1650,N_1512,N_1590);
xnor U1651 (N_1651,N_1594,N_1488);
or U1652 (N_1652,N_1581,N_1587);
or U1653 (N_1653,N_1405,N_1459);
nand U1654 (N_1654,N_1586,N_1525);
nand U1655 (N_1655,N_1517,N_1417);
nor U1656 (N_1656,N_1404,N_1402);
nand U1657 (N_1657,N_1496,N_1421);
xor U1658 (N_1658,N_1555,N_1503);
or U1659 (N_1659,N_1529,N_1439);
or U1660 (N_1660,N_1593,N_1410);
nor U1661 (N_1661,N_1570,N_1432);
or U1662 (N_1662,N_1422,N_1519);
nand U1663 (N_1663,N_1487,N_1533);
or U1664 (N_1664,N_1473,N_1400);
xnor U1665 (N_1665,N_1418,N_1426);
nor U1666 (N_1666,N_1501,N_1579);
nor U1667 (N_1667,N_1482,N_1430);
or U1668 (N_1668,N_1431,N_1569);
nor U1669 (N_1669,N_1548,N_1449);
nor U1670 (N_1670,N_1567,N_1419);
or U1671 (N_1671,N_1547,N_1546);
nand U1672 (N_1672,N_1425,N_1428);
and U1673 (N_1673,N_1498,N_1532);
nor U1674 (N_1674,N_1455,N_1460);
xnor U1675 (N_1675,N_1444,N_1483);
xnor U1676 (N_1676,N_1443,N_1447);
nand U1677 (N_1677,N_1484,N_1552);
nor U1678 (N_1678,N_1461,N_1481);
nand U1679 (N_1679,N_1511,N_1545);
or U1680 (N_1680,N_1474,N_1506);
or U1681 (N_1681,N_1585,N_1424);
nor U1682 (N_1682,N_1458,N_1486);
nor U1683 (N_1683,N_1415,N_1502);
xor U1684 (N_1684,N_1520,N_1509);
xnor U1685 (N_1685,N_1541,N_1564);
nand U1686 (N_1686,N_1469,N_1592);
and U1687 (N_1687,N_1514,N_1539);
nor U1688 (N_1688,N_1436,N_1411);
nor U1689 (N_1689,N_1505,N_1563);
nand U1690 (N_1690,N_1556,N_1589);
nor U1691 (N_1691,N_1429,N_1575);
xor U1692 (N_1692,N_1524,N_1406);
nor U1693 (N_1693,N_1495,N_1521);
or U1694 (N_1694,N_1440,N_1452);
xnor U1695 (N_1695,N_1413,N_1537);
and U1696 (N_1696,N_1416,N_1435);
or U1697 (N_1697,N_1578,N_1591);
or U1698 (N_1698,N_1523,N_1568);
nand U1699 (N_1699,N_1446,N_1572);
nand U1700 (N_1700,N_1453,N_1418);
nor U1701 (N_1701,N_1552,N_1485);
xnor U1702 (N_1702,N_1581,N_1417);
and U1703 (N_1703,N_1525,N_1569);
nand U1704 (N_1704,N_1536,N_1407);
nor U1705 (N_1705,N_1474,N_1418);
nand U1706 (N_1706,N_1599,N_1475);
or U1707 (N_1707,N_1462,N_1438);
nand U1708 (N_1708,N_1469,N_1471);
xor U1709 (N_1709,N_1550,N_1578);
or U1710 (N_1710,N_1574,N_1527);
or U1711 (N_1711,N_1558,N_1504);
or U1712 (N_1712,N_1549,N_1520);
nand U1713 (N_1713,N_1464,N_1517);
xnor U1714 (N_1714,N_1433,N_1415);
or U1715 (N_1715,N_1595,N_1515);
nor U1716 (N_1716,N_1523,N_1444);
nand U1717 (N_1717,N_1559,N_1426);
or U1718 (N_1718,N_1545,N_1466);
nand U1719 (N_1719,N_1523,N_1423);
and U1720 (N_1720,N_1426,N_1544);
or U1721 (N_1721,N_1471,N_1563);
nand U1722 (N_1722,N_1544,N_1585);
nor U1723 (N_1723,N_1425,N_1541);
and U1724 (N_1724,N_1583,N_1457);
xnor U1725 (N_1725,N_1524,N_1577);
xnor U1726 (N_1726,N_1468,N_1416);
nor U1727 (N_1727,N_1462,N_1447);
nand U1728 (N_1728,N_1581,N_1462);
nor U1729 (N_1729,N_1586,N_1592);
and U1730 (N_1730,N_1583,N_1416);
nor U1731 (N_1731,N_1465,N_1558);
nor U1732 (N_1732,N_1556,N_1409);
and U1733 (N_1733,N_1454,N_1445);
or U1734 (N_1734,N_1405,N_1472);
xnor U1735 (N_1735,N_1521,N_1565);
and U1736 (N_1736,N_1451,N_1498);
xnor U1737 (N_1737,N_1592,N_1438);
nand U1738 (N_1738,N_1419,N_1559);
or U1739 (N_1739,N_1489,N_1522);
nor U1740 (N_1740,N_1559,N_1562);
nand U1741 (N_1741,N_1541,N_1502);
xnor U1742 (N_1742,N_1422,N_1534);
nand U1743 (N_1743,N_1439,N_1473);
xnor U1744 (N_1744,N_1405,N_1442);
or U1745 (N_1745,N_1463,N_1533);
xor U1746 (N_1746,N_1482,N_1534);
nor U1747 (N_1747,N_1514,N_1460);
xnor U1748 (N_1748,N_1434,N_1451);
nand U1749 (N_1749,N_1408,N_1581);
and U1750 (N_1750,N_1455,N_1474);
or U1751 (N_1751,N_1538,N_1573);
and U1752 (N_1752,N_1464,N_1422);
nand U1753 (N_1753,N_1453,N_1470);
nor U1754 (N_1754,N_1466,N_1474);
xnor U1755 (N_1755,N_1445,N_1417);
and U1756 (N_1756,N_1521,N_1575);
and U1757 (N_1757,N_1496,N_1575);
nor U1758 (N_1758,N_1554,N_1477);
xnor U1759 (N_1759,N_1415,N_1584);
nand U1760 (N_1760,N_1420,N_1451);
nor U1761 (N_1761,N_1531,N_1555);
nand U1762 (N_1762,N_1552,N_1575);
or U1763 (N_1763,N_1532,N_1476);
xor U1764 (N_1764,N_1418,N_1483);
xnor U1765 (N_1765,N_1486,N_1591);
xnor U1766 (N_1766,N_1464,N_1596);
nand U1767 (N_1767,N_1420,N_1568);
xnor U1768 (N_1768,N_1535,N_1559);
nor U1769 (N_1769,N_1587,N_1405);
or U1770 (N_1770,N_1459,N_1556);
nand U1771 (N_1771,N_1547,N_1490);
xnor U1772 (N_1772,N_1575,N_1514);
nand U1773 (N_1773,N_1440,N_1578);
and U1774 (N_1774,N_1439,N_1513);
or U1775 (N_1775,N_1530,N_1586);
or U1776 (N_1776,N_1400,N_1570);
nand U1777 (N_1777,N_1540,N_1515);
and U1778 (N_1778,N_1476,N_1580);
or U1779 (N_1779,N_1563,N_1422);
nand U1780 (N_1780,N_1553,N_1445);
nand U1781 (N_1781,N_1512,N_1583);
nand U1782 (N_1782,N_1423,N_1540);
and U1783 (N_1783,N_1554,N_1445);
nand U1784 (N_1784,N_1499,N_1473);
and U1785 (N_1785,N_1441,N_1588);
nor U1786 (N_1786,N_1425,N_1476);
nand U1787 (N_1787,N_1540,N_1500);
nand U1788 (N_1788,N_1481,N_1466);
or U1789 (N_1789,N_1439,N_1527);
or U1790 (N_1790,N_1553,N_1514);
nor U1791 (N_1791,N_1403,N_1420);
and U1792 (N_1792,N_1529,N_1515);
or U1793 (N_1793,N_1411,N_1569);
nor U1794 (N_1794,N_1401,N_1582);
xor U1795 (N_1795,N_1456,N_1468);
nor U1796 (N_1796,N_1435,N_1486);
or U1797 (N_1797,N_1540,N_1444);
and U1798 (N_1798,N_1555,N_1401);
or U1799 (N_1799,N_1517,N_1569);
xor U1800 (N_1800,N_1633,N_1709);
and U1801 (N_1801,N_1605,N_1636);
or U1802 (N_1802,N_1708,N_1769);
nand U1803 (N_1803,N_1785,N_1701);
xor U1804 (N_1804,N_1675,N_1750);
or U1805 (N_1805,N_1726,N_1614);
xnor U1806 (N_1806,N_1639,N_1642);
nand U1807 (N_1807,N_1753,N_1608);
or U1808 (N_1808,N_1719,N_1770);
and U1809 (N_1809,N_1745,N_1733);
xnor U1810 (N_1810,N_1667,N_1681);
xor U1811 (N_1811,N_1660,N_1654);
and U1812 (N_1812,N_1786,N_1629);
nand U1813 (N_1813,N_1649,N_1673);
or U1814 (N_1814,N_1656,N_1603);
nor U1815 (N_1815,N_1742,N_1775);
nand U1816 (N_1816,N_1662,N_1706);
or U1817 (N_1817,N_1645,N_1665);
nand U1818 (N_1818,N_1694,N_1641);
and U1819 (N_1819,N_1778,N_1657);
nor U1820 (N_1820,N_1621,N_1781);
nand U1821 (N_1821,N_1628,N_1680);
nand U1822 (N_1822,N_1692,N_1679);
or U1823 (N_1823,N_1748,N_1626);
and U1824 (N_1824,N_1682,N_1620);
or U1825 (N_1825,N_1615,N_1691);
nand U1826 (N_1826,N_1686,N_1767);
nor U1827 (N_1827,N_1702,N_1723);
nor U1828 (N_1828,N_1796,N_1666);
and U1829 (N_1829,N_1794,N_1722);
nor U1830 (N_1830,N_1631,N_1793);
nand U1831 (N_1831,N_1610,N_1768);
xnor U1832 (N_1832,N_1711,N_1618);
xor U1833 (N_1833,N_1655,N_1779);
and U1834 (N_1834,N_1650,N_1652);
and U1835 (N_1835,N_1715,N_1765);
xor U1836 (N_1836,N_1772,N_1735);
xor U1837 (N_1837,N_1713,N_1670);
xnor U1838 (N_1838,N_1617,N_1717);
xnor U1839 (N_1839,N_1634,N_1700);
or U1840 (N_1840,N_1787,N_1728);
nand U1841 (N_1841,N_1622,N_1710);
xor U1842 (N_1842,N_1724,N_1688);
nand U1843 (N_1843,N_1799,N_1703);
or U1844 (N_1844,N_1697,N_1782);
nand U1845 (N_1845,N_1795,N_1611);
nand U1846 (N_1846,N_1734,N_1741);
nor U1847 (N_1847,N_1749,N_1647);
nand U1848 (N_1848,N_1612,N_1774);
nand U1849 (N_1849,N_1630,N_1725);
and U1850 (N_1850,N_1658,N_1606);
nor U1851 (N_1851,N_1689,N_1676);
nor U1852 (N_1852,N_1671,N_1672);
xnor U1853 (N_1853,N_1627,N_1766);
nor U1854 (N_1854,N_1721,N_1747);
nand U1855 (N_1855,N_1777,N_1632);
nand U1856 (N_1856,N_1684,N_1637);
and U1857 (N_1857,N_1714,N_1659);
xor U1858 (N_1858,N_1600,N_1685);
nor U1859 (N_1859,N_1616,N_1613);
nand U1860 (N_1860,N_1755,N_1623);
and U1861 (N_1861,N_1698,N_1643);
nand U1862 (N_1862,N_1687,N_1690);
and U1863 (N_1863,N_1788,N_1789);
xnor U1864 (N_1864,N_1661,N_1635);
nor U1865 (N_1865,N_1696,N_1727);
and U1866 (N_1866,N_1764,N_1695);
xor U1867 (N_1867,N_1602,N_1607);
xnor U1868 (N_1868,N_1797,N_1798);
and U1869 (N_1869,N_1761,N_1754);
nand U1870 (N_1870,N_1646,N_1699);
and U1871 (N_1871,N_1773,N_1730);
and U1872 (N_1872,N_1752,N_1663);
nand U1873 (N_1873,N_1678,N_1758);
and U1874 (N_1874,N_1731,N_1762);
nor U1875 (N_1875,N_1792,N_1780);
and U1876 (N_1876,N_1737,N_1677);
nand U1877 (N_1877,N_1791,N_1732);
and U1878 (N_1878,N_1648,N_1609);
or U1879 (N_1879,N_1729,N_1693);
nand U1880 (N_1880,N_1668,N_1716);
nand U1881 (N_1881,N_1653,N_1743);
xnor U1882 (N_1882,N_1739,N_1740);
or U1883 (N_1883,N_1718,N_1601);
and U1884 (N_1884,N_1771,N_1720);
and U1885 (N_1885,N_1705,N_1783);
and U1886 (N_1886,N_1744,N_1738);
and U1887 (N_1887,N_1604,N_1736);
nand U1888 (N_1888,N_1776,N_1669);
or U1889 (N_1889,N_1757,N_1640);
or U1890 (N_1890,N_1707,N_1674);
xnor U1891 (N_1891,N_1790,N_1683);
and U1892 (N_1892,N_1751,N_1712);
nand U1893 (N_1893,N_1638,N_1756);
or U1894 (N_1894,N_1651,N_1704);
xnor U1895 (N_1895,N_1746,N_1625);
and U1896 (N_1896,N_1619,N_1624);
nand U1897 (N_1897,N_1784,N_1664);
and U1898 (N_1898,N_1644,N_1760);
and U1899 (N_1899,N_1763,N_1759);
nand U1900 (N_1900,N_1761,N_1700);
xnor U1901 (N_1901,N_1677,N_1646);
and U1902 (N_1902,N_1670,N_1706);
nor U1903 (N_1903,N_1757,N_1627);
nor U1904 (N_1904,N_1683,N_1782);
and U1905 (N_1905,N_1799,N_1653);
xor U1906 (N_1906,N_1628,N_1677);
nor U1907 (N_1907,N_1766,N_1709);
xor U1908 (N_1908,N_1730,N_1716);
and U1909 (N_1909,N_1609,N_1703);
nor U1910 (N_1910,N_1714,N_1631);
nand U1911 (N_1911,N_1601,N_1734);
and U1912 (N_1912,N_1627,N_1760);
nand U1913 (N_1913,N_1794,N_1678);
xor U1914 (N_1914,N_1793,N_1645);
and U1915 (N_1915,N_1685,N_1601);
or U1916 (N_1916,N_1797,N_1616);
or U1917 (N_1917,N_1651,N_1785);
nand U1918 (N_1918,N_1692,N_1752);
nor U1919 (N_1919,N_1684,N_1784);
nor U1920 (N_1920,N_1719,N_1717);
nand U1921 (N_1921,N_1640,N_1662);
nand U1922 (N_1922,N_1760,N_1619);
and U1923 (N_1923,N_1720,N_1784);
nand U1924 (N_1924,N_1660,N_1705);
and U1925 (N_1925,N_1689,N_1723);
nor U1926 (N_1926,N_1610,N_1717);
and U1927 (N_1927,N_1775,N_1786);
nor U1928 (N_1928,N_1764,N_1600);
or U1929 (N_1929,N_1749,N_1659);
and U1930 (N_1930,N_1638,N_1662);
xor U1931 (N_1931,N_1746,N_1627);
xor U1932 (N_1932,N_1742,N_1638);
nand U1933 (N_1933,N_1735,N_1649);
or U1934 (N_1934,N_1733,N_1735);
xor U1935 (N_1935,N_1745,N_1791);
nand U1936 (N_1936,N_1665,N_1684);
and U1937 (N_1937,N_1670,N_1720);
nand U1938 (N_1938,N_1697,N_1663);
nand U1939 (N_1939,N_1622,N_1632);
xnor U1940 (N_1940,N_1619,N_1770);
nand U1941 (N_1941,N_1700,N_1649);
nand U1942 (N_1942,N_1691,N_1642);
and U1943 (N_1943,N_1732,N_1652);
or U1944 (N_1944,N_1645,N_1640);
nor U1945 (N_1945,N_1729,N_1648);
or U1946 (N_1946,N_1610,N_1601);
and U1947 (N_1947,N_1661,N_1749);
nor U1948 (N_1948,N_1611,N_1600);
nand U1949 (N_1949,N_1776,N_1702);
nor U1950 (N_1950,N_1621,N_1741);
and U1951 (N_1951,N_1730,N_1637);
xor U1952 (N_1952,N_1647,N_1738);
nor U1953 (N_1953,N_1786,N_1684);
nor U1954 (N_1954,N_1678,N_1608);
or U1955 (N_1955,N_1684,N_1712);
and U1956 (N_1956,N_1734,N_1767);
and U1957 (N_1957,N_1625,N_1775);
xnor U1958 (N_1958,N_1711,N_1642);
nor U1959 (N_1959,N_1626,N_1754);
nor U1960 (N_1960,N_1645,N_1762);
xor U1961 (N_1961,N_1709,N_1679);
and U1962 (N_1962,N_1734,N_1661);
xor U1963 (N_1963,N_1740,N_1702);
xor U1964 (N_1964,N_1790,N_1679);
xor U1965 (N_1965,N_1635,N_1682);
or U1966 (N_1966,N_1657,N_1647);
nand U1967 (N_1967,N_1738,N_1601);
nand U1968 (N_1968,N_1711,N_1606);
xnor U1969 (N_1969,N_1667,N_1798);
nand U1970 (N_1970,N_1678,N_1765);
xor U1971 (N_1971,N_1630,N_1703);
xnor U1972 (N_1972,N_1668,N_1739);
or U1973 (N_1973,N_1760,N_1710);
and U1974 (N_1974,N_1682,N_1632);
and U1975 (N_1975,N_1637,N_1713);
xnor U1976 (N_1976,N_1734,N_1653);
and U1977 (N_1977,N_1689,N_1719);
or U1978 (N_1978,N_1702,N_1666);
nand U1979 (N_1979,N_1794,N_1706);
or U1980 (N_1980,N_1722,N_1736);
and U1981 (N_1981,N_1746,N_1621);
nand U1982 (N_1982,N_1723,N_1712);
or U1983 (N_1983,N_1772,N_1750);
and U1984 (N_1984,N_1796,N_1616);
xnor U1985 (N_1985,N_1789,N_1628);
nand U1986 (N_1986,N_1735,N_1698);
or U1987 (N_1987,N_1752,N_1742);
nor U1988 (N_1988,N_1727,N_1708);
and U1989 (N_1989,N_1668,N_1690);
xor U1990 (N_1990,N_1628,N_1753);
nor U1991 (N_1991,N_1667,N_1753);
xnor U1992 (N_1992,N_1602,N_1659);
xor U1993 (N_1993,N_1649,N_1729);
nand U1994 (N_1994,N_1698,N_1771);
and U1995 (N_1995,N_1669,N_1772);
xnor U1996 (N_1996,N_1630,N_1709);
xnor U1997 (N_1997,N_1645,N_1749);
and U1998 (N_1998,N_1795,N_1768);
nor U1999 (N_1999,N_1672,N_1634);
xor U2000 (N_2000,N_1875,N_1923);
xnor U2001 (N_2001,N_1817,N_1819);
or U2002 (N_2002,N_1838,N_1834);
nand U2003 (N_2003,N_1927,N_1984);
nor U2004 (N_2004,N_1931,N_1874);
and U2005 (N_2005,N_1846,N_1805);
xor U2006 (N_2006,N_1993,N_1917);
and U2007 (N_2007,N_1866,N_1974);
nor U2008 (N_2008,N_1975,N_1926);
nand U2009 (N_2009,N_1899,N_1961);
nor U2010 (N_2010,N_1988,N_1954);
or U2011 (N_2011,N_1936,N_1980);
nand U2012 (N_2012,N_1895,N_1880);
nor U2013 (N_2013,N_1821,N_1890);
nor U2014 (N_2014,N_1893,N_1950);
xnor U2015 (N_2015,N_1892,N_1982);
xnor U2016 (N_2016,N_1887,N_1918);
nand U2017 (N_2017,N_1932,N_1983);
nor U2018 (N_2018,N_1889,N_1958);
or U2019 (N_2019,N_1946,N_1913);
nor U2020 (N_2020,N_1881,N_1904);
or U2021 (N_2021,N_1930,N_1940);
or U2022 (N_2022,N_1827,N_1815);
and U2023 (N_2023,N_1992,N_1990);
or U2024 (N_2024,N_1989,N_1909);
or U2025 (N_2025,N_1861,N_1951);
nand U2026 (N_2026,N_1920,N_1826);
xnor U2027 (N_2027,N_1891,N_1994);
nor U2028 (N_2028,N_1999,N_1832);
and U2029 (N_2029,N_1981,N_1929);
nand U2030 (N_2030,N_1841,N_1911);
xor U2031 (N_2031,N_1970,N_1850);
nor U2032 (N_2032,N_1823,N_1908);
xor U2033 (N_2033,N_1901,N_1803);
nor U2034 (N_2034,N_1860,N_1977);
or U2035 (N_2035,N_1806,N_1877);
nand U2036 (N_2036,N_1822,N_1998);
and U2037 (N_2037,N_1828,N_1844);
or U2038 (N_2038,N_1949,N_1839);
nor U2039 (N_2039,N_1804,N_1955);
or U2040 (N_2040,N_1863,N_1813);
nor U2041 (N_2041,N_1985,N_1944);
nand U2042 (N_2042,N_1856,N_1915);
or U2043 (N_2043,N_1964,N_1959);
and U2044 (N_2044,N_1972,N_1808);
or U2045 (N_2045,N_1830,N_1816);
or U2046 (N_2046,N_1888,N_1829);
nand U2047 (N_2047,N_1870,N_1924);
and U2048 (N_2048,N_1845,N_1953);
nor U2049 (N_2049,N_1818,N_1995);
or U2050 (N_2050,N_1840,N_1968);
xor U2051 (N_2051,N_1802,N_1945);
and U2052 (N_2052,N_1810,N_1836);
nand U2053 (N_2053,N_1871,N_1935);
nand U2054 (N_2054,N_1962,N_1987);
and U2055 (N_2055,N_1878,N_1801);
or U2056 (N_2056,N_1842,N_1865);
nand U2057 (N_2057,N_1922,N_1848);
xor U2058 (N_2058,N_1948,N_1978);
and U2059 (N_2059,N_1885,N_1837);
and U2060 (N_2060,N_1900,N_1857);
nor U2061 (N_2061,N_1869,N_1824);
nand U2062 (N_2062,N_1854,N_1876);
xor U2063 (N_2063,N_1973,N_1835);
xor U2064 (N_2064,N_1898,N_1905);
or U2065 (N_2065,N_1872,N_1941);
xnor U2066 (N_2066,N_1965,N_1912);
and U2067 (N_2067,N_1903,N_1939);
nand U2068 (N_2068,N_1896,N_1879);
or U2069 (N_2069,N_1938,N_1979);
and U2070 (N_2070,N_1966,N_1886);
nor U2071 (N_2071,N_1858,N_1925);
nand U2072 (N_2072,N_1910,N_1969);
nand U2073 (N_2073,N_1942,N_1807);
and U2074 (N_2074,N_1934,N_1947);
xnor U2075 (N_2075,N_1897,N_1967);
nand U2076 (N_2076,N_1867,N_1921);
nand U2077 (N_2077,N_1957,N_1812);
or U2078 (N_2078,N_1919,N_1825);
nor U2079 (N_2079,N_1963,N_1882);
nor U2080 (N_2080,N_1902,N_1831);
nor U2081 (N_2081,N_1843,N_1956);
xnor U2082 (N_2082,N_1849,N_1859);
and U2083 (N_2083,N_1933,N_1907);
and U2084 (N_2084,N_1883,N_1800);
xnor U2085 (N_2085,N_1991,N_1906);
nor U2086 (N_2086,N_1811,N_1894);
xnor U2087 (N_2087,N_1864,N_1833);
and U2088 (N_2088,N_1855,N_1952);
xnor U2089 (N_2089,N_1873,N_1852);
xnor U2090 (N_2090,N_1928,N_1851);
or U2091 (N_2091,N_1853,N_1868);
or U2092 (N_2092,N_1997,N_1814);
nand U2093 (N_2093,N_1976,N_1847);
or U2094 (N_2094,N_1937,N_1884);
xnor U2095 (N_2095,N_1820,N_1862);
nor U2096 (N_2096,N_1809,N_1916);
or U2097 (N_2097,N_1996,N_1971);
nand U2098 (N_2098,N_1986,N_1943);
and U2099 (N_2099,N_1914,N_1960);
or U2100 (N_2100,N_1918,N_1865);
and U2101 (N_2101,N_1892,N_1916);
nor U2102 (N_2102,N_1856,N_1877);
nand U2103 (N_2103,N_1960,N_1921);
or U2104 (N_2104,N_1910,N_1857);
xnor U2105 (N_2105,N_1823,N_1950);
xor U2106 (N_2106,N_1831,N_1835);
xnor U2107 (N_2107,N_1828,N_1813);
or U2108 (N_2108,N_1962,N_1864);
and U2109 (N_2109,N_1897,N_1904);
xnor U2110 (N_2110,N_1851,N_1888);
and U2111 (N_2111,N_1818,N_1987);
nand U2112 (N_2112,N_1944,N_1858);
and U2113 (N_2113,N_1923,N_1874);
and U2114 (N_2114,N_1966,N_1972);
nand U2115 (N_2115,N_1860,N_1975);
nor U2116 (N_2116,N_1813,N_1874);
nor U2117 (N_2117,N_1896,N_1849);
nor U2118 (N_2118,N_1871,N_1829);
nor U2119 (N_2119,N_1872,N_1961);
xor U2120 (N_2120,N_1958,N_1850);
and U2121 (N_2121,N_1839,N_1861);
and U2122 (N_2122,N_1973,N_1836);
xnor U2123 (N_2123,N_1872,N_1962);
or U2124 (N_2124,N_1900,N_1948);
xor U2125 (N_2125,N_1872,N_1923);
xnor U2126 (N_2126,N_1964,N_1869);
nor U2127 (N_2127,N_1938,N_1989);
or U2128 (N_2128,N_1937,N_1913);
nor U2129 (N_2129,N_1801,N_1800);
and U2130 (N_2130,N_1805,N_1892);
nand U2131 (N_2131,N_1980,N_1819);
xnor U2132 (N_2132,N_1975,N_1809);
or U2133 (N_2133,N_1905,N_1881);
and U2134 (N_2134,N_1850,N_1896);
nand U2135 (N_2135,N_1807,N_1990);
or U2136 (N_2136,N_1865,N_1988);
and U2137 (N_2137,N_1948,N_1856);
or U2138 (N_2138,N_1800,N_1947);
xnor U2139 (N_2139,N_1947,N_1892);
xor U2140 (N_2140,N_1949,N_1968);
nand U2141 (N_2141,N_1932,N_1810);
xnor U2142 (N_2142,N_1897,N_1968);
nor U2143 (N_2143,N_1834,N_1930);
nor U2144 (N_2144,N_1889,N_1980);
nand U2145 (N_2145,N_1850,N_1943);
nand U2146 (N_2146,N_1967,N_1814);
nor U2147 (N_2147,N_1971,N_1801);
xnor U2148 (N_2148,N_1890,N_1856);
or U2149 (N_2149,N_1981,N_1837);
nor U2150 (N_2150,N_1814,N_1935);
nor U2151 (N_2151,N_1849,N_1945);
or U2152 (N_2152,N_1819,N_1813);
nand U2153 (N_2153,N_1858,N_1819);
or U2154 (N_2154,N_1805,N_1843);
and U2155 (N_2155,N_1826,N_1841);
nor U2156 (N_2156,N_1891,N_1924);
nand U2157 (N_2157,N_1897,N_1909);
and U2158 (N_2158,N_1891,N_1960);
and U2159 (N_2159,N_1832,N_1856);
and U2160 (N_2160,N_1966,N_1863);
and U2161 (N_2161,N_1870,N_1820);
or U2162 (N_2162,N_1929,N_1844);
or U2163 (N_2163,N_1992,N_1965);
nor U2164 (N_2164,N_1844,N_1967);
and U2165 (N_2165,N_1866,N_1917);
and U2166 (N_2166,N_1838,N_1969);
or U2167 (N_2167,N_1856,N_1928);
nand U2168 (N_2168,N_1854,N_1845);
nor U2169 (N_2169,N_1801,N_1924);
and U2170 (N_2170,N_1914,N_1825);
nand U2171 (N_2171,N_1956,N_1976);
nand U2172 (N_2172,N_1872,N_1943);
nand U2173 (N_2173,N_1844,N_1996);
xnor U2174 (N_2174,N_1985,N_1927);
xor U2175 (N_2175,N_1813,N_1848);
nor U2176 (N_2176,N_1902,N_1962);
and U2177 (N_2177,N_1833,N_1918);
or U2178 (N_2178,N_1886,N_1935);
nor U2179 (N_2179,N_1818,N_1833);
or U2180 (N_2180,N_1968,N_1819);
nand U2181 (N_2181,N_1948,N_1980);
nor U2182 (N_2182,N_1911,N_1849);
or U2183 (N_2183,N_1802,N_1865);
nor U2184 (N_2184,N_1891,N_1915);
and U2185 (N_2185,N_1950,N_1904);
and U2186 (N_2186,N_1880,N_1840);
nor U2187 (N_2187,N_1806,N_1866);
and U2188 (N_2188,N_1942,N_1961);
and U2189 (N_2189,N_1945,N_1939);
or U2190 (N_2190,N_1880,N_1936);
nand U2191 (N_2191,N_1843,N_1872);
and U2192 (N_2192,N_1957,N_1985);
xor U2193 (N_2193,N_1949,N_1951);
or U2194 (N_2194,N_1854,N_1853);
and U2195 (N_2195,N_1983,N_1837);
nor U2196 (N_2196,N_1853,N_1831);
nor U2197 (N_2197,N_1814,N_1861);
nand U2198 (N_2198,N_1933,N_1987);
or U2199 (N_2199,N_1844,N_1887);
or U2200 (N_2200,N_2171,N_2179);
and U2201 (N_2201,N_2020,N_2033);
nand U2202 (N_2202,N_2009,N_2100);
nor U2203 (N_2203,N_2012,N_2156);
or U2204 (N_2204,N_2099,N_2070);
nand U2205 (N_2205,N_2154,N_2076);
and U2206 (N_2206,N_2178,N_2136);
nor U2207 (N_2207,N_2101,N_2132);
nand U2208 (N_2208,N_2087,N_2198);
nand U2209 (N_2209,N_2022,N_2174);
nor U2210 (N_2210,N_2073,N_2196);
nand U2211 (N_2211,N_2036,N_2180);
nand U2212 (N_2212,N_2108,N_2181);
nand U2213 (N_2213,N_2029,N_2123);
nand U2214 (N_2214,N_2089,N_2008);
and U2215 (N_2215,N_2106,N_2096);
or U2216 (N_2216,N_2090,N_2064);
nand U2217 (N_2217,N_2169,N_2110);
xnor U2218 (N_2218,N_2151,N_2142);
or U2219 (N_2219,N_2030,N_2117);
nor U2220 (N_2220,N_2015,N_2148);
xnor U2221 (N_2221,N_2121,N_2134);
xnor U2222 (N_2222,N_2042,N_2043);
nor U2223 (N_2223,N_2027,N_2160);
and U2224 (N_2224,N_2000,N_2054);
nand U2225 (N_2225,N_2102,N_2082);
or U2226 (N_2226,N_2086,N_2112);
nand U2227 (N_2227,N_2140,N_2092);
or U2228 (N_2228,N_2126,N_2039);
and U2229 (N_2229,N_2056,N_2115);
nand U2230 (N_2230,N_2113,N_2053);
xnor U2231 (N_2231,N_2135,N_2028);
nand U2232 (N_2232,N_2044,N_2195);
or U2233 (N_2233,N_2010,N_2111);
nor U2234 (N_2234,N_2062,N_2018);
nand U2235 (N_2235,N_2078,N_2159);
or U2236 (N_2236,N_2164,N_2122);
and U2237 (N_2237,N_2193,N_2048);
and U2238 (N_2238,N_2003,N_2093);
nor U2239 (N_2239,N_2023,N_2107);
xor U2240 (N_2240,N_2130,N_2055);
nand U2241 (N_2241,N_2167,N_2016);
and U2242 (N_2242,N_2041,N_2128);
nand U2243 (N_2243,N_2103,N_2095);
nand U2244 (N_2244,N_2131,N_2066);
xnor U2245 (N_2245,N_2119,N_2185);
xnor U2246 (N_2246,N_2035,N_2158);
nor U2247 (N_2247,N_2147,N_2186);
xnor U2248 (N_2248,N_2081,N_2137);
nand U2249 (N_2249,N_2125,N_2072);
nand U2250 (N_2250,N_2155,N_2138);
xnor U2251 (N_2251,N_2077,N_2060);
xnor U2252 (N_2252,N_2014,N_2192);
and U2253 (N_2253,N_2091,N_2045);
xnor U2254 (N_2254,N_2046,N_2040);
xnor U2255 (N_2255,N_2176,N_2047);
nand U2256 (N_2256,N_2133,N_2005);
nor U2257 (N_2257,N_2032,N_2199);
and U2258 (N_2258,N_2004,N_2157);
and U2259 (N_2259,N_2061,N_2166);
nand U2260 (N_2260,N_2050,N_2197);
xnor U2261 (N_2261,N_2172,N_2168);
nand U2262 (N_2262,N_2191,N_2145);
xor U2263 (N_2263,N_2001,N_2094);
nand U2264 (N_2264,N_2074,N_2083);
nor U2265 (N_2265,N_2052,N_2031);
nand U2266 (N_2266,N_2051,N_2165);
and U2267 (N_2267,N_2127,N_2071);
nand U2268 (N_2268,N_2170,N_2105);
xor U2269 (N_2269,N_2065,N_2175);
nand U2270 (N_2270,N_2184,N_2152);
and U2271 (N_2271,N_2057,N_2129);
xor U2272 (N_2272,N_2058,N_2049);
or U2273 (N_2273,N_2002,N_2024);
xor U2274 (N_2274,N_2189,N_2013);
or U2275 (N_2275,N_2080,N_2084);
or U2276 (N_2276,N_2124,N_2187);
xnor U2277 (N_2277,N_2085,N_2162);
or U2278 (N_2278,N_2067,N_2007);
nor U2279 (N_2279,N_2017,N_2109);
and U2280 (N_2280,N_2026,N_2161);
or U2281 (N_2281,N_2097,N_2182);
xnor U2282 (N_2282,N_2063,N_2011);
or U2283 (N_2283,N_2163,N_2021);
nor U2284 (N_2284,N_2141,N_2150);
nor U2285 (N_2285,N_2143,N_2006);
nand U2286 (N_2286,N_2144,N_2088);
xor U2287 (N_2287,N_2183,N_2069);
xnor U2288 (N_2288,N_2149,N_2120);
or U2289 (N_2289,N_2098,N_2188);
xor U2290 (N_2290,N_2173,N_2019);
xnor U2291 (N_2291,N_2038,N_2037);
nor U2292 (N_2292,N_2116,N_2114);
or U2293 (N_2293,N_2075,N_2118);
or U2294 (N_2294,N_2194,N_2153);
or U2295 (N_2295,N_2068,N_2104);
and U2296 (N_2296,N_2034,N_2177);
nand U2297 (N_2297,N_2146,N_2139);
xor U2298 (N_2298,N_2025,N_2059);
xor U2299 (N_2299,N_2190,N_2079);
or U2300 (N_2300,N_2180,N_2140);
xnor U2301 (N_2301,N_2068,N_2065);
nor U2302 (N_2302,N_2022,N_2082);
or U2303 (N_2303,N_2148,N_2173);
or U2304 (N_2304,N_2047,N_2033);
nor U2305 (N_2305,N_2190,N_2064);
and U2306 (N_2306,N_2135,N_2146);
nor U2307 (N_2307,N_2020,N_2035);
nor U2308 (N_2308,N_2145,N_2090);
and U2309 (N_2309,N_2069,N_2188);
or U2310 (N_2310,N_2177,N_2077);
xor U2311 (N_2311,N_2127,N_2184);
xnor U2312 (N_2312,N_2030,N_2063);
or U2313 (N_2313,N_2009,N_2007);
nand U2314 (N_2314,N_2079,N_2177);
nand U2315 (N_2315,N_2113,N_2073);
and U2316 (N_2316,N_2130,N_2196);
or U2317 (N_2317,N_2148,N_2143);
nor U2318 (N_2318,N_2199,N_2050);
or U2319 (N_2319,N_2066,N_2114);
xor U2320 (N_2320,N_2156,N_2068);
nor U2321 (N_2321,N_2091,N_2141);
or U2322 (N_2322,N_2164,N_2160);
or U2323 (N_2323,N_2039,N_2159);
nor U2324 (N_2324,N_2053,N_2106);
nor U2325 (N_2325,N_2056,N_2144);
nor U2326 (N_2326,N_2014,N_2152);
nor U2327 (N_2327,N_2172,N_2186);
and U2328 (N_2328,N_2080,N_2003);
or U2329 (N_2329,N_2174,N_2198);
xnor U2330 (N_2330,N_2111,N_2159);
nand U2331 (N_2331,N_2067,N_2033);
xnor U2332 (N_2332,N_2012,N_2009);
and U2333 (N_2333,N_2112,N_2039);
nand U2334 (N_2334,N_2040,N_2032);
nor U2335 (N_2335,N_2148,N_2049);
and U2336 (N_2336,N_2130,N_2014);
nand U2337 (N_2337,N_2030,N_2133);
or U2338 (N_2338,N_2002,N_2153);
and U2339 (N_2339,N_2150,N_2112);
nand U2340 (N_2340,N_2015,N_2095);
nor U2341 (N_2341,N_2041,N_2061);
nand U2342 (N_2342,N_2160,N_2136);
nand U2343 (N_2343,N_2189,N_2099);
or U2344 (N_2344,N_2034,N_2022);
nor U2345 (N_2345,N_2098,N_2177);
nand U2346 (N_2346,N_2085,N_2119);
and U2347 (N_2347,N_2053,N_2190);
and U2348 (N_2348,N_2160,N_2057);
nand U2349 (N_2349,N_2068,N_2186);
xnor U2350 (N_2350,N_2090,N_2078);
nand U2351 (N_2351,N_2048,N_2058);
or U2352 (N_2352,N_2187,N_2130);
or U2353 (N_2353,N_2000,N_2077);
and U2354 (N_2354,N_2185,N_2190);
nor U2355 (N_2355,N_2024,N_2096);
nand U2356 (N_2356,N_2160,N_2199);
and U2357 (N_2357,N_2049,N_2195);
and U2358 (N_2358,N_2104,N_2124);
nor U2359 (N_2359,N_2069,N_2107);
and U2360 (N_2360,N_2147,N_2102);
or U2361 (N_2361,N_2054,N_2013);
nor U2362 (N_2362,N_2160,N_2081);
or U2363 (N_2363,N_2133,N_2024);
nor U2364 (N_2364,N_2035,N_2092);
and U2365 (N_2365,N_2142,N_2039);
and U2366 (N_2366,N_2099,N_2065);
nand U2367 (N_2367,N_2080,N_2119);
nand U2368 (N_2368,N_2064,N_2108);
nand U2369 (N_2369,N_2134,N_2093);
nor U2370 (N_2370,N_2041,N_2100);
xor U2371 (N_2371,N_2164,N_2112);
nand U2372 (N_2372,N_2057,N_2087);
nand U2373 (N_2373,N_2028,N_2110);
nand U2374 (N_2374,N_2108,N_2027);
nor U2375 (N_2375,N_2132,N_2129);
and U2376 (N_2376,N_2018,N_2057);
nor U2377 (N_2377,N_2035,N_2087);
xnor U2378 (N_2378,N_2062,N_2169);
or U2379 (N_2379,N_2013,N_2000);
and U2380 (N_2380,N_2039,N_2027);
or U2381 (N_2381,N_2025,N_2191);
and U2382 (N_2382,N_2085,N_2147);
xnor U2383 (N_2383,N_2035,N_2101);
xnor U2384 (N_2384,N_2097,N_2132);
and U2385 (N_2385,N_2184,N_2078);
nor U2386 (N_2386,N_2150,N_2006);
and U2387 (N_2387,N_2006,N_2151);
nand U2388 (N_2388,N_2006,N_2067);
nor U2389 (N_2389,N_2179,N_2168);
and U2390 (N_2390,N_2179,N_2066);
xor U2391 (N_2391,N_2152,N_2059);
xnor U2392 (N_2392,N_2126,N_2017);
xor U2393 (N_2393,N_2081,N_2108);
nand U2394 (N_2394,N_2150,N_2191);
nand U2395 (N_2395,N_2079,N_2040);
nor U2396 (N_2396,N_2146,N_2013);
or U2397 (N_2397,N_2142,N_2165);
and U2398 (N_2398,N_2051,N_2090);
xor U2399 (N_2399,N_2192,N_2007);
and U2400 (N_2400,N_2325,N_2366);
nor U2401 (N_2401,N_2248,N_2215);
or U2402 (N_2402,N_2254,N_2285);
or U2403 (N_2403,N_2329,N_2290);
or U2404 (N_2404,N_2397,N_2211);
xnor U2405 (N_2405,N_2362,N_2288);
and U2406 (N_2406,N_2357,N_2392);
nor U2407 (N_2407,N_2244,N_2220);
xnor U2408 (N_2408,N_2260,N_2353);
xnor U2409 (N_2409,N_2365,N_2330);
or U2410 (N_2410,N_2286,N_2289);
xor U2411 (N_2411,N_2270,N_2359);
xor U2412 (N_2412,N_2210,N_2371);
nor U2413 (N_2413,N_2219,N_2367);
xor U2414 (N_2414,N_2204,N_2318);
and U2415 (N_2415,N_2275,N_2389);
nor U2416 (N_2416,N_2320,N_2292);
and U2417 (N_2417,N_2280,N_2282);
and U2418 (N_2418,N_2317,N_2276);
or U2419 (N_2419,N_2242,N_2377);
xor U2420 (N_2420,N_2373,N_2298);
or U2421 (N_2421,N_2247,N_2202);
or U2422 (N_2422,N_2201,N_2296);
and U2423 (N_2423,N_2370,N_2229);
nand U2424 (N_2424,N_2213,N_2251);
and U2425 (N_2425,N_2338,N_2256);
or U2426 (N_2426,N_2360,N_2295);
nand U2427 (N_2427,N_2235,N_2369);
nor U2428 (N_2428,N_2343,N_2200);
nor U2429 (N_2429,N_2283,N_2245);
nor U2430 (N_2430,N_2203,N_2223);
nor U2431 (N_2431,N_2249,N_2393);
xor U2432 (N_2432,N_2305,N_2316);
nand U2433 (N_2433,N_2307,N_2272);
xnor U2434 (N_2434,N_2314,N_2333);
nor U2435 (N_2435,N_2304,N_2206);
or U2436 (N_2436,N_2252,N_2354);
nand U2437 (N_2437,N_2340,N_2299);
and U2438 (N_2438,N_2351,N_2238);
xnor U2439 (N_2439,N_2394,N_2375);
nand U2440 (N_2440,N_2342,N_2246);
xnor U2441 (N_2441,N_2355,N_2216);
xor U2442 (N_2442,N_2291,N_2390);
or U2443 (N_2443,N_2380,N_2271);
nor U2444 (N_2444,N_2266,N_2207);
xor U2445 (N_2445,N_2384,N_2332);
and U2446 (N_2446,N_2279,N_2269);
or U2447 (N_2447,N_2278,N_2230);
nor U2448 (N_2448,N_2372,N_2225);
or U2449 (N_2449,N_2261,N_2311);
or U2450 (N_2450,N_2396,N_2381);
or U2451 (N_2451,N_2335,N_2234);
or U2452 (N_2452,N_2258,N_2301);
nor U2453 (N_2453,N_2217,N_2358);
nand U2454 (N_2454,N_2387,N_2265);
and U2455 (N_2455,N_2331,N_2221);
and U2456 (N_2456,N_2239,N_2374);
nand U2457 (N_2457,N_2300,N_2209);
nor U2458 (N_2458,N_2344,N_2293);
nor U2459 (N_2459,N_2297,N_2341);
nand U2460 (N_2460,N_2257,N_2259);
nor U2461 (N_2461,N_2321,N_2347);
nand U2462 (N_2462,N_2339,N_2364);
or U2463 (N_2463,N_2326,N_2262);
nand U2464 (N_2464,N_2334,N_2336);
or U2465 (N_2465,N_2356,N_2264);
and U2466 (N_2466,N_2228,N_2287);
nand U2467 (N_2467,N_2227,N_2263);
nor U2468 (N_2468,N_2391,N_2323);
and U2469 (N_2469,N_2383,N_2205);
and U2470 (N_2470,N_2319,N_2303);
xnor U2471 (N_2471,N_2231,N_2379);
or U2472 (N_2472,N_2218,N_2310);
nand U2473 (N_2473,N_2250,N_2281);
nand U2474 (N_2474,N_2337,N_2232);
or U2475 (N_2475,N_2352,N_2368);
nand U2476 (N_2476,N_2268,N_2386);
and U2477 (N_2477,N_2322,N_2345);
or U2478 (N_2478,N_2243,N_2388);
or U2479 (N_2479,N_2399,N_2306);
nor U2480 (N_2480,N_2240,N_2294);
nand U2481 (N_2481,N_2255,N_2222);
nand U2482 (N_2482,N_2214,N_2324);
and U2483 (N_2483,N_2363,N_2208);
nor U2484 (N_2484,N_2309,N_2308);
nand U2485 (N_2485,N_2346,N_2236);
nor U2486 (N_2486,N_2302,N_2376);
and U2487 (N_2487,N_2237,N_2398);
nand U2488 (N_2488,N_2267,N_2224);
or U2489 (N_2489,N_2253,N_2315);
nand U2490 (N_2490,N_2350,N_2348);
nor U2491 (N_2491,N_2274,N_2328);
xnor U2492 (N_2492,N_2395,N_2313);
xor U2493 (N_2493,N_2273,N_2378);
or U2494 (N_2494,N_2349,N_2361);
or U2495 (N_2495,N_2382,N_2226);
and U2496 (N_2496,N_2312,N_2385);
nand U2497 (N_2497,N_2277,N_2284);
nor U2498 (N_2498,N_2212,N_2327);
nor U2499 (N_2499,N_2241,N_2233);
xor U2500 (N_2500,N_2278,N_2248);
nor U2501 (N_2501,N_2234,N_2261);
nand U2502 (N_2502,N_2253,N_2235);
nor U2503 (N_2503,N_2332,N_2302);
or U2504 (N_2504,N_2356,N_2310);
nor U2505 (N_2505,N_2376,N_2342);
nor U2506 (N_2506,N_2222,N_2374);
and U2507 (N_2507,N_2272,N_2344);
or U2508 (N_2508,N_2202,N_2256);
and U2509 (N_2509,N_2306,N_2212);
nand U2510 (N_2510,N_2359,N_2240);
or U2511 (N_2511,N_2310,N_2252);
or U2512 (N_2512,N_2200,N_2379);
nand U2513 (N_2513,N_2236,N_2239);
xor U2514 (N_2514,N_2279,N_2220);
xor U2515 (N_2515,N_2320,N_2332);
and U2516 (N_2516,N_2249,N_2336);
nand U2517 (N_2517,N_2291,N_2268);
and U2518 (N_2518,N_2394,N_2207);
nor U2519 (N_2519,N_2304,N_2276);
nor U2520 (N_2520,N_2383,N_2233);
nand U2521 (N_2521,N_2311,N_2227);
and U2522 (N_2522,N_2240,N_2246);
nand U2523 (N_2523,N_2267,N_2203);
xnor U2524 (N_2524,N_2327,N_2313);
nand U2525 (N_2525,N_2375,N_2310);
xor U2526 (N_2526,N_2242,N_2232);
and U2527 (N_2527,N_2358,N_2270);
xor U2528 (N_2528,N_2339,N_2272);
nand U2529 (N_2529,N_2340,N_2283);
nor U2530 (N_2530,N_2313,N_2355);
xnor U2531 (N_2531,N_2260,N_2270);
and U2532 (N_2532,N_2230,N_2311);
and U2533 (N_2533,N_2239,N_2324);
nor U2534 (N_2534,N_2221,N_2259);
or U2535 (N_2535,N_2263,N_2300);
and U2536 (N_2536,N_2264,N_2393);
nand U2537 (N_2537,N_2277,N_2265);
nand U2538 (N_2538,N_2230,N_2308);
nand U2539 (N_2539,N_2305,N_2257);
and U2540 (N_2540,N_2350,N_2232);
or U2541 (N_2541,N_2236,N_2307);
xor U2542 (N_2542,N_2318,N_2367);
nor U2543 (N_2543,N_2237,N_2359);
nor U2544 (N_2544,N_2261,N_2218);
and U2545 (N_2545,N_2307,N_2380);
or U2546 (N_2546,N_2229,N_2283);
nand U2547 (N_2547,N_2301,N_2351);
or U2548 (N_2548,N_2219,N_2250);
and U2549 (N_2549,N_2207,N_2314);
nor U2550 (N_2550,N_2284,N_2336);
and U2551 (N_2551,N_2392,N_2329);
nor U2552 (N_2552,N_2295,N_2381);
nand U2553 (N_2553,N_2206,N_2335);
or U2554 (N_2554,N_2344,N_2222);
nor U2555 (N_2555,N_2347,N_2293);
nor U2556 (N_2556,N_2213,N_2353);
xnor U2557 (N_2557,N_2261,N_2256);
nand U2558 (N_2558,N_2303,N_2301);
or U2559 (N_2559,N_2264,N_2325);
nand U2560 (N_2560,N_2280,N_2240);
nor U2561 (N_2561,N_2399,N_2257);
nor U2562 (N_2562,N_2345,N_2320);
or U2563 (N_2563,N_2315,N_2272);
and U2564 (N_2564,N_2291,N_2284);
nor U2565 (N_2565,N_2359,N_2289);
xnor U2566 (N_2566,N_2263,N_2319);
and U2567 (N_2567,N_2355,N_2373);
nand U2568 (N_2568,N_2249,N_2398);
nor U2569 (N_2569,N_2388,N_2278);
and U2570 (N_2570,N_2216,N_2243);
xnor U2571 (N_2571,N_2207,N_2330);
xnor U2572 (N_2572,N_2389,N_2241);
nand U2573 (N_2573,N_2265,N_2272);
xor U2574 (N_2574,N_2390,N_2203);
and U2575 (N_2575,N_2341,N_2288);
xor U2576 (N_2576,N_2279,N_2233);
nand U2577 (N_2577,N_2395,N_2296);
xnor U2578 (N_2578,N_2288,N_2278);
nand U2579 (N_2579,N_2342,N_2317);
or U2580 (N_2580,N_2370,N_2351);
and U2581 (N_2581,N_2254,N_2392);
nor U2582 (N_2582,N_2340,N_2374);
xor U2583 (N_2583,N_2348,N_2363);
xnor U2584 (N_2584,N_2364,N_2286);
and U2585 (N_2585,N_2267,N_2321);
nor U2586 (N_2586,N_2357,N_2281);
and U2587 (N_2587,N_2326,N_2398);
or U2588 (N_2588,N_2393,N_2254);
nor U2589 (N_2589,N_2352,N_2259);
and U2590 (N_2590,N_2332,N_2228);
or U2591 (N_2591,N_2285,N_2301);
nor U2592 (N_2592,N_2342,N_2345);
nand U2593 (N_2593,N_2352,N_2345);
nand U2594 (N_2594,N_2395,N_2212);
and U2595 (N_2595,N_2262,N_2294);
nor U2596 (N_2596,N_2280,N_2364);
or U2597 (N_2597,N_2240,N_2203);
or U2598 (N_2598,N_2347,N_2341);
nand U2599 (N_2599,N_2289,N_2223);
and U2600 (N_2600,N_2577,N_2409);
nor U2601 (N_2601,N_2499,N_2418);
and U2602 (N_2602,N_2517,N_2401);
nor U2603 (N_2603,N_2501,N_2591);
and U2604 (N_2604,N_2573,N_2562);
and U2605 (N_2605,N_2415,N_2527);
and U2606 (N_2606,N_2525,N_2444);
xor U2607 (N_2607,N_2479,N_2496);
and U2608 (N_2608,N_2585,N_2426);
nand U2609 (N_2609,N_2436,N_2572);
nor U2610 (N_2610,N_2464,N_2542);
nand U2611 (N_2611,N_2400,N_2476);
nand U2612 (N_2612,N_2534,N_2469);
nand U2613 (N_2613,N_2557,N_2554);
nor U2614 (N_2614,N_2462,N_2402);
nand U2615 (N_2615,N_2404,N_2471);
nand U2616 (N_2616,N_2536,N_2595);
nor U2617 (N_2617,N_2410,N_2455);
nand U2618 (N_2618,N_2553,N_2488);
and U2619 (N_2619,N_2457,N_2569);
nor U2620 (N_2620,N_2495,N_2434);
xor U2621 (N_2621,N_2526,N_2508);
and U2622 (N_2622,N_2543,N_2505);
xor U2623 (N_2623,N_2438,N_2592);
xor U2624 (N_2624,N_2506,N_2458);
nand U2625 (N_2625,N_2448,N_2437);
xor U2626 (N_2626,N_2502,N_2578);
xnor U2627 (N_2627,N_2538,N_2452);
or U2628 (N_2628,N_2579,N_2568);
or U2629 (N_2629,N_2419,N_2587);
nand U2630 (N_2630,N_2477,N_2561);
nand U2631 (N_2631,N_2531,N_2430);
xor U2632 (N_2632,N_2441,N_2582);
and U2633 (N_2633,N_2445,N_2483);
xor U2634 (N_2634,N_2588,N_2412);
nor U2635 (N_2635,N_2449,N_2580);
nor U2636 (N_2636,N_2484,N_2551);
or U2637 (N_2637,N_2432,N_2552);
and U2638 (N_2638,N_2407,N_2451);
nand U2639 (N_2639,N_2498,N_2431);
nand U2640 (N_2640,N_2529,N_2514);
xnor U2641 (N_2641,N_2428,N_2593);
and U2642 (N_2642,N_2468,N_2541);
and U2643 (N_2643,N_2490,N_2439);
nor U2644 (N_2644,N_2465,N_2533);
nand U2645 (N_2645,N_2416,N_2540);
and U2646 (N_2646,N_2544,N_2467);
nand U2647 (N_2647,N_2598,N_2559);
nor U2648 (N_2648,N_2516,N_2481);
nor U2649 (N_2649,N_2513,N_2403);
nand U2650 (N_2650,N_2589,N_2548);
nor U2651 (N_2651,N_2466,N_2443);
or U2652 (N_2652,N_2475,N_2509);
nor U2653 (N_2653,N_2493,N_2480);
or U2654 (N_2654,N_2567,N_2522);
nor U2655 (N_2655,N_2532,N_2523);
or U2656 (N_2656,N_2420,N_2459);
nand U2657 (N_2657,N_2425,N_2470);
and U2658 (N_2658,N_2442,N_2507);
xnor U2659 (N_2659,N_2492,N_2427);
or U2660 (N_2660,N_2596,N_2560);
or U2661 (N_2661,N_2421,N_2535);
nand U2662 (N_2662,N_2406,N_2504);
and U2663 (N_2663,N_2539,N_2446);
or U2664 (N_2664,N_2474,N_2494);
nor U2665 (N_2665,N_2586,N_2429);
or U2666 (N_2666,N_2571,N_2460);
nand U2667 (N_2667,N_2515,N_2574);
or U2668 (N_2668,N_2500,N_2583);
nor U2669 (N_2669,N_2581,N_2417);
or U2670 (N_2670,N_2491,N_2435);
or U2671 (N_2671,N_2594,N_2497);
or U2672 (N_2672,N_2511,N_2456);
nand U2673 (N_2673,N_2450,N_2570);
nand U2674 (N_2674,N_2411,N_2546);
nor U2675 (N_2675,N_2521,N_2472);
xnor U2676 (N_2676,N_2510,N_2566);
xnor U2677 (N_2677,N_2590,N_2482);
and U2678 (N_2678,N_2413,N_2520);
and U2679 (N_2679,N_2576,N_2486);
xor U2680 (N_2680,N_2422,N_2564);
nand U2681 (N_2681,N_2489,N_2524);
or U2682 (N_2682,N_2487,N_2565);
and U2683 (N_2683,N_2556,N_2447);
nand U2684 (N_2684,N_2599,N_2537);
nor U2685 (N_2685,N_2597,N_2512);
nand U2686 (N_2686,N_2528,N_2530);
nand U2687 (N_2687,N_2549,N_2545);
xnor U2688 (N_2688,N_2405,N_2547);
nor U2689 (N_2689,N_2485,N_2478);
xnor U2690 (N_2690,N_2453,N_2440);
or U2691 (N_2691,N_2414,N_2518);
and U2692 (N_2692,N_2550,N_2408);
xor U2693 (N_2693,N_2423,N_2503);
or U2694 (N_2694,N_2519,N_2563);
xor U2695 (N_2695,N_2584,N_2454);
and U2696 (N_2696,N_2558,N_2463);
nor U2697 (N_2697,N_2461,N_2424);
xnor U2698 (N_2698,N_2433,N_2575);
xnor U2699 (N_2699,N_2555,N_2473);
xnor U2700 (N_2700,N_2550,N_2434);
nor U2701 (N_2701,N_2586,N_2444);
xnor U2702 (N_2702,N_2505,N_2539);
nand U2703 (N_2703,N_2495,N_2532);
and U2704 (N_2704,N_2424,N_2462);
nand U2705 (N_2705,N_2480,N_2551);
or U2706 (N_2706,N_2422,N_2533);
nor U2707 (N_2707,N_2483,N_2490);
nor U2708 (N_2708,N_2561,N_2524);
or U2709 (N_2709,N_2555,N_2533);
xnor U2710 (N_2710,N_2509,N_2403);
nor U2711 (N_2711,N_2549,N_2440);
nand U2712 (N_2712,N_2475,N_2593);
or U2713 (N_2713,N_2543,N_2536);
xnor U2714 (N_2714,N_2447,N_2580);
xor U2715 (N_2715,N_2593,N_2581);
or U2716 (N_2716,N_2545,N_2553);
nand U2717 (N_2717,N_2424,N_2528);
and U2718 (N_2718,N_2500,N_2499);
and U2719 (N_2719,N_2495,N_2566);
xnor U2720 (N_2720,N_2471,N_2407);
or U2721 (N_2721,N_2461,N_2503);
nor U2722 (N_2722,N_2491,N_2490);
and U2723 (N_2723,N_2447,N_2470);
and U2724 (N_2724,N_2519,N_2474);
xor U2725 (N_2725,N_2522,N_2561);
or U2726 (N_2726,N_2591,N_2475);
xnor U2727 (N_2727,N_2448,N_2499);
or U2728 (N_2728,N_2567,N_2413);
nor U2729 (N_2729,N_2494,N_2599);
nand U2730 (N_2730,N_2423,N_2516);
xor U2731 (N_2731,N_2438,N_2529);
or U2732 (N_2732,N_2531,N_2457);
or U2733 (N_2733,N_2495,N_2564);
nor U2734 (N_2734,N_2508,N_2563);
nor U2735 (N_2735,N_2563,N_2443);
nor U2736 (N_2736,N_2433,N_2476);
and U2737 (N_2737,N_2480,N_2518);
xnor U2738 (N_2738,N_2552,N_2415);
nand U2739 (N_2739,N_2587,N_2491);
and U2740 (N_2740,N_2495,N_2576);
nand U2741 (N_2741,N_2596,N_2591);
nand U2742 (N_2742,N_2409,N_2482);
and U2743 (N_2743,N_2581,N_2453);
and U2744 (N_2744,N_2455,N_2434);
nor U2745 (N_2745,N_2503,N_2527);
and U2746 (N_2746,N_2476,N_2432);
nor U2747 (N_2747,N_2482,N_2432);
xnor U2748 (N_2748,N_2402,N_2464);
nand U2749 (N_2749,N_2446,N_2487);
and U2750 (N_2750,N_2569,N_2478);
or U2751 (N_2751,N_2507,N_2477);
nand U2752 (N_2752,N_2407,N_2479);
nand U2753 (N_2753,N_2429,N_2517);
nor U2754 (N_2754,N_2429,N_2573);
nand U2755 (N_2755,N_2568,N_2509);
and U2756 (N_2756,N_2527,N_2422);
nand U2757 (N_2757,N_2466,N_2574);
or U2758 (N_2758,N_2437,N_2562);
nand U2759 (N_2759,N_2530,N_2585);
and U2760 (N_2760,N_2594,N_2451);
nor U2761 (N_2761,N_2435,N_2444);
and U2762 (N_2762,N_2573,N_2487);
or U2763 (N_2763,N_2413,N_2465);
nand U2764 (N_2764,N_2424,N_2539);
xnor U2765 (N_2765,N_2517,N_2579);
or U2766 (N_2766,N_2538,N_2498);
nor U2767 (N_2767,N_2589,N_2556);
and U2768 (N_2768,N_2552,N_2439);
nor U2769 (N_2769,N_2462,N_2598);
xnor U2770 (N_2770,N_2592,N_2448);
nand U2771 (N_2771,N_2593,N_2446);
xnor U2772 (N_2772,N_2520,N_2509);
nand U2773 (N_2773,N_2570,N_2405);
or U2774 (N_2774,N_2521,N_2541);
xor U2775 (N_2775,N_2516,N_2438);
xnor U2776 (N_2776,N_2494,N_2592);
nand U2777 (N_2777,N_2562,N_2485);
or U2778 (N_2778,N_2593,N_2422);
nand U2779 (N_2779,N_2555,N_2512);
nand U2780 (N_2780,N_2456,N_2519);
xor U2781 (N_2781,N_2494,N_2447);
nor U2782 (N_2782,N_2592,N_2474);
nor U2783 (N_2783,N_2543,N_2581);
nand U2784 (N_2784,N_2543,N_2568);
nor U2785 (N_2785,N_2530,N_2574);
xor U2786 (N_2786,N_2444,N_2493);
nor U2787 (N_2787,N_2412,N_2427);
or U2788 (N_2788,N_2501,N_2534);
or U2789 (N_2789,N_2540,N_2491);
nand U2790 (N_2790,N_2570,N_2572);
nand U2791 (N_2791,N_2519,N_2472);
and U2792 (N_2792,N_2407,N_2584);
or U2793 (N_2793,N_2410,N_2417);
or U2794 (N_2794,N_2478,N_2400);
nand U2795 (N_2795,N_2592,N_2596);
and U2796 (N_2796,N_2469,N_2554);
xor U2797 (N_2797,N_2529,N_2537);
nand U2798 (N_2798,N_2567,N_2409);
and U2799 (N_2799,N_2503,N_2455);
nand U2800 (N_2800,N_2719,N_2603);
or U2801 (N_2801,N_2727,N_2779);
and U2802 (N_2802,N_2652,N_2608);
and U2803 (N_2803,N_2620,N_2758);
and U2804 (N_2804,N_2692,N_2734);
xnor U2805 (N_2805,N_2761,N_2743);
nand U2806 (N_2806,N_2666,N_2646);
or U2807 (N_2807,N_2637,N_2775);
nand U2808 (N_2808,N_2639,N_2686);
or U2809 (N_2809,N_2760,N_2694);
nor U2810 (N_2810,N_2755,N_2752);
nand U2811 (N_2811,N_2757,N_2685);
nand U2812 (N_2812,N_2650,N_2713);
xor U2813 (N_2813,N_2628,N_2661);
and U2814 (N_2814,N_2684,N_2705);
or U2815 (N_2815,N_2768,N_2682);
or U2816 (N_2816,N_2662,N_2701);
or U2817 (N_2817,N_2740,N_2785);
nand U2818 (N_2818,N_2640,N_2712);
and U2819 (N_2819,N_2674,N_2792);
and U2820 (N_2820,N_2716,N_2633);
nand U2821 (N_2821,N_2797,N_2624);
nand U2822 (N_2822,N_2625,N_2714);
xor U2823 (N_2823,N_2651,N_2645);
or U2824 (N_2824,N_2749,N_2765);
and U2825 (N_2825,N_2638,N_2704);
and U2826 (N_2826,N_2750,N_2790);
nand U2827 (N_2827,N_2618,N_2711);
xnor U2828 (N_2828,N_2723,N_2626);
and U2829 (N_2829,N_2776,N_2722);
nor U2830 (N_2830,N_2798,N_2751);
nand U2831 (N_2831,N_2673,N_2641);
and U2832 (N_2832,N_2663,N_2770);
or U2833 (N_2833,N_2655,N_2700);
nor U2834 (N_2834,N_2709,N_2720);
nand U2835 (N_2835,N_2616,N_2738);
xnor U2836 (N_2836,N_2613,N_2617);
and U2837 (N_2837,N_2724,N_2676);
and U2838 (N_2838,N_2605,N_2794);
nand U2839 (N_2839,N_2687,N_2693);
or U2840 (N_2840,N_2781,N_2683);
nor U2841 (N_2841,N_2799,N_2621);
xnor U2842 (N_2842,N_2600,N_2767);
and U2843 (N_2843,N_2773,N_2609);
nand U2844 (N_2844,N_2707,N_2644);
and U2845 (N_2845,N_2736,N_2690);
nand U2846 (N_2846,N_2632,N_2680);
and U2847 (N_2847,N_2715,N_2622);
or U2848 (N_2848,N_2766,N_2677);
xor U2849 (N_2849,N_2664,N_2729);
and U2850 (N_2850,N_2699,N_2759);
or U2851 (N_2851,N_2631,N_2656);
xor U2852 (N_2852,N_2745,N_2654);
xor U2853 (N_2853,N_2610,N_2726);
and U2854 (N_2854,N_2703,N_2630);
nor U2855 (N_2855,N_2706,N_2737);
and U2856 (N_2856,N_2748,N_2691);
nor U2857 (N_2857,N_2717,N_2636);
and U2858 (N_2858,N_2791,N_2702);
xor U2859 (N_2859,N_2718,N_2754);
nand U2860 (N_2860,N_2777,N_2787);
nor U2861 (N_2861,N_2698,N_2739);
xor U2862 (N_2862,N_2774,N_2606);
nor U2863 (N_2863,N_2614,N_2764);
nand U2864 (N_2864,N_2753,N_2681);
nor U2865 (N_2865,N_2695,N_2769);
or U2866 (N_2866,N_2629,N_2782);
nand U2867 (N_2867,N_2601,N_2667);
or U2868 (N_2868,N_2619,N_2733);
nor U2869 (N_2869,N_2643,N_2710);
and U2870 (N_2870,N_2658,N_2762);
nor U2871 (N_2871,N_2789,N_2642);
xnor U2872 (N_2872,N_2786,N_2730);
nand U2873 (N_2873,N_2611,N_2756);
nand U2874 (N_2874,N_2689,N_2742);
or U2875 (N_2875,N_2649,N_2725);
or U2876 (N_2876,N_2602,N_2635);
nor U2877 (N_2877,N_2697,N_2795);
and U2878 (N_2878,N_2772,N_2778);
xnor U2879 (N_2879,N_2688,N_2627);
and U2880 (N_2880,N_2744,N_2678);
or U2881 (N_2881,N_2623,N_2657);
or U2882 (N_2882,N_2747,N_2728);
nand U2883 (N_2883,N_2671,N_2653);
and U2884 (N_2884,N_2612,N_2746);
nor U2885 (N_2885,N_2607,N_2670);
nor U2886 (N_2886,N_2780,N_2660);
nor U2887 (N_2887,N_2665,N_2696);
and U2888 (N_2888,N_2679,N_2735);
xnor U2889 (N_2889,N_2659,N_2741);
or U2890 (N_2890,N_2731,N_2672);
xor U2891 (N_2891,N_2668,N_2763);
nor U2892 (N_2892,N_2708,N_2647);
xnor U2893 (N_2893,N_2771,N_2784);
nand U2894 (N_2894,N_2604,N_2648);
and U2895 (N_2895,N_2675,N_2793);
xnor U2896 (N_2896,N_2783,N_2732);
or U2897 (N_2897,N_2721,N_2796);
xor U2898 (N_2898,N_2634,N_2788);
and U2899 (N_2899,N_2669,N_2615);
xnor U2900 (N_2900,N_2688,N_2680);
and U2901 (N_2901,N_2754,N_2611);
nor U2902 (N_2902,N_2699,N_2697);
nand U2903 (N_2903,N_2663,N_2647);
or U2904 (N_2904,N_2785,N_2722);
nor U2905 (N_2905,N_2681,N_2748);
xor U2906 (N_2906,N_2761,N_2636);
nor U2907 (N_2907,N_2610,N_2664);
or U2908 (N_2908,N_2771,N_2674);
and U2909 (N_2909,N_2659,N_2660);
nor U2910 (N_2910,N_2659,N_2760);
nand U2911 (N_2911,N_2611,N_2660);
nand U2912 (N_2912,N_2613,N_2647);
or U2913 (N_2913,N_2716,N_2698);
xnor U2914 (N_2914,N_2642,N_2652);
nor U2915 (N_2915,N_2662,N_2707);
or U2916 (N_2916,N_2635,N_2606);
xnor U2917 (N_2917,N_2768,N_2623);
or U2918 (N_2918,N_2725,N_2744);
xor U2919 (N_2919,N_2782,N_2604);
or U2920 (N_2920,N_2624,N_2710);
nand U2921 (N_2921,N_2652,N_2664);
or U2922 (N_2922,N_2604,N_2662);
and U2923 (N_2923,N_2685,N_2794);
or U2924 (N_2924,N_2601,N_2694);
and U2925 (N_2925,N_2738,N_2786);
or U2926 (N_2926,N_2622,N_2671);
and U2927 (N_2927,N_2622,N_2731);
or U2928 (N_2928,N_2748,N_2616);
or U2929 (N_2929,N_2683,N_2663);
and U2930 (N_2930,N_2671,N_2638);
nand U2931 (N_2931,N_2652,N_2749);
nor U2932 (N_2932,N_2732,N_2799);
and U2933 (N_2933,N_2784,N_2794);
nor U2934 (N_2934,N_2757,N_2719);
xnor U2935 (N_2935,N_2633,N_2730);
nand U2936 (N_2936,N_2713,N_2640);
nor U2937 (N_2937,N_2633,N_2744);
xnor U2938 (N_2938,N_2656,N_2607);
nor U2939 (N_2939,N_2612,N_2695);
or U2940 (N_2940,N_2737,N_2686);
nand U2941 (N_2941,N_2766,N_2774);
xnor U2942 (N_2942,N_2665,N_2703);
xor U2943 (N_2943,N_2724,N_2787);
xnor U2944 (N_2944,N_2619,N_2762);
nor U2945 (N_2945,N_2604,N_2762);
xor U2946 (N_2946,N_2795,N_2709);
and U2947 (N_2947,N_2798,N_2722);
or U2948 (N_2948,N_2713,N_2648);
nor U2949 (N_2949,N_2772,N_2750);
or U2950 (N_2950,N_2696,N_2686);
nor U2951 (N_2951,N_2757,N_2606);
xnor U2952 (N_2952,N_2691,N_2751);
nor U2953 (N_2953,N_2788,N_2731);
nor U2954 (N_2954,N_2683,N_2601);
nand U2955 (N_2955,N_2749,N_2783);
xor U2956 (N_2956,N_2684,N_2678);
nor U2957 (N_2957,N_2656,N_2782);
nor U2958 (N_2958,N_2788,N_2745);
xnor U2959 (N_2959,N_2772,N_2620);
nand U2960 (N_2960,N_2783,N_2651);
nor U2961 (N_2961,N_2754,N_2650);
and U2962 (N_2962,N_2615,N_2701);
or U2963 (N_2963,N_2646,N_2730);
xnor U2964 (N_2964,N_2765,N_2623);
nor U2965 (N_2965,N_2719,N_2768);
or U2966 (N_2966,N_2758,N_2798);
and U2967 (N_2967,N_2680,N_2733);
nor U2968 (N_2968,N_2743,N_2633);
xor U2969 (N_2969,N_2783,N_2786);
xor U2970 (N_2970,N_2715,N_2642);
or U2971 (N_2971,N_2721,N_2642);
xnor U2972 (N_2972,N_2744,N_2654);
nor U2973 (N_2973,N_2755,N_2651);
nand U2974 (N_2974,N_2710,N_2655);
nor U2975 (N_2975,N_2615,N_2666);
and U2976 (N_2976,N_2704,N_2648);
nand U2977 (N_2977,N_2627,N_2710);
nor U2978 (N_2978,N_2606,N_2756);
or U2979 (N_2979,N_2702,N_2660);
and U2980 (N_2980,N_2746,N_2642);
nand U2981 (N_2981,N_2659,N_2700);
or U2982 (N_2982,N_2746,N_2782);
xnor U2983 (N_2983,N_2756,N_2722);
or U2984 (N_2984,N_2779,N_2701);
xnor U2985 (N_2985,N_2733,N_2757);
or U2986 (N_2986,N_2710,N_2626);
nor U2987 (N_2987,N_2617,N_2644);
and U2988 (N_2988,N_2785,N_2792);
nor U2989 (N_2989,N_2646,N_2760);
and U2990 (N_2990,N_2755,N_2689);
and U2991 (N_2991,N_2734,N_2602);
nand U2992 (N_2992,N_2792,N_2666);
and U2993 (N_2993,N_2753,N_2616);
nor U2994 (N_2994,N_2742,N_2683);
xnor U2995 (N_2995,N_2759,N_2666);
nand U2996 (N_2996,N_2754,N_2738);
nor U2997 (N_2997,N_2678,N_2659);
or U2998 (N_2998,N_2658,N_2754);
xnor U2999 (N_2999,N_2768,N_2672);
nand U3000 (N_3000,N_2927,N_2909);
or U3001 (N_3001,N_2844,N_2967);
and U3002 (N_3002,N_2925,N_2980);
nor U3003 (N_3003,N_2889,N_2839);
and U3004 (N_3004,N_2881,N_2929);
nand U3005 (N_3005,N_2876,N_2880);
xnor U3006 (N_3006,N_2862,N_2851);
xnor U3007 (N_3007,N_2823,N_2986);
nand U3008 (N_3008,N_2838,N_2883);
or U3009 (N_3009,N_2928,N_2933);
nand U3010 (N_3010,N_2841,N_2902);
nor U3011 (N_3011,N_2951,N_2935);
nand U3012 (N_3012,N_2979,N_2907);
nor U3013 (N_3013,N_2975,N_2891);
nor U3014 (N_3014,N_2842,N_2898);
xor U3015 (N_3015,N_2906,N_2895);
and U3016 (N_3016,N_2957,N_2830);
and U3017 (N_3017,N_2988,N_2859);
xnor U3018 (N_3018,N_2805,N_2807);
or U3019 (N_3019,N_2977,N_2853);
or U3020 (N_3020,N_2854,N_2834);
and U3021 (N_3021,N_2921,N_2952);
nand U3022 (N_3022,N_2912,N_2843);
xor U3023 (N_3023,N_2845,N_2824);
or U3024 (N_3024,N_2917,N_2972);
nor U3025 (N_3025,N_2829,N_2875);
and U3026 (N_3026,N_2802,N_2865);
and U3027 (N_3027,N_2885,N_2899);
and U3028 (N_3028,N_2837,N_2870);
or U3029 (N_3029,N_2835,N_2945);
and U3030 (N_3030,N_2825,N_2950);
and U3031 (N_3031,N_2846,N_2993);
nor U3032 (N_3032,N_2874,N_2857);
nor U3033 (N_3033,N_2827,N_2888);
and U3034 (N_3034,N_2974,N_2913);
nand U3035 (N_3035,N_2966,N_2908);
or U3036 (N_3036,N_2813,N_2978);
xor U3037 (N_3037,N_2811,N_2984);
nor U3038 (N_3038,N_2878,N_2848);
and U3039 (N_3039,N_2969,N_2937);
nor U3040 (N_3040,N_2812,N_2996);
or U3041 (N_3041,N_2953,N_2948);
nand U3042 (N_3042,N_2954,N_2814);
and U3043 (N_3043,N_2926,N_2923);
nor U3044 (N_3044,N_2867,N_2970);
nand U3045 (N_3045,N_2973,N_2915);
nand U3046 (N_3046,N_2877,N_2801);
nand U3047 (N_3047,N_2817,N_2855);
nand U3048 (N_3048,N_2956,N_2965);
and U3049 (N_3049,N_2882,N_2968);
nand U3050 (N_3050,N_2871,N_2916);
and U3051 (N_3051,N_2866,N_2941);
xnor U3052 (N_3052,N_2836,N_2868);
or U3053 (N_3053,N_2920,N_2987);
and U3054 (N_3054,N_2803,N_2959);
or U3055 (N_3055,N_2997,N_2903);
nor U3056 (N_3056,N_2858,N_2860);
nor U3057 (N_3057,N_2893,N_2924);
and U3058 (N_3058,N_2991,N_2936);
xnor U3059 (N_3059,N_2905,N_2861);
nand U3060 (N_3060,N_2989,N_2810);
xnor U3061 (N_3061,N_2892,N_2897);
nand U3062 (N_3062,N_2822,N_2938);
xnor U3063 (N_3063,N_2981,N_2890);
xor U3064 (N_3064,N_2849,N_2808);
nor U3065 (N_3065,N_2955,N_2960);
and U3066 (N_3066,N_2832,N_2863);
nand U3067 (N_3067,N_2961,N_2911);
nor U3068 (N_3068,N_2943,N_2939);
or U3069 (N_3069,N_2963,N_2922);
nor U3070 (N_3070,N_2930,N_2932);
or U3071 (N_3071,N_2850,N_2982);
and U3072 (N_3072,N_2872,N_2949);
or U3073 (N_3073,N_2840,N_2934);
xor U3074 (N_3074,N_2809,N_2879);
nand U3075 (N_3075,N_2833,N_2919);
xnor U3076 (N_3076,N_2820,N_2821);
xor U3077 (N_3077,N_2819,N_2964);
nor U3078 (N_3078,N_2958,N_2887);
and U3079 (N_3079,N_2990,N_2896);
or U3080 (N_3080,N_2901,N_2998);
xnor U3081 (N_3081,N_2999,N_2804);
nand U3082 (N_3082,N_2847,N_2918);
xnor U3083 (N_3083,N_2962,N_2904);
and U3084 (N_3084,N_2971,N_2884);
or U3085 (N_3085,N_2947,N_2992);
xor U3086 (N_3086,N_2852,N_2826);
and U3087 (N_3087,N_2864,N_2985);
nor U3088 (N_3088,N_2931,N_2856);
or U3089 (N_3089,N_2946,N_2869);
nor U3090 (N_3090,N_2873,N_2815);
and U3091 (N_3091,N_2800,N_2828);
and U3092 (N_3092,N_2816,N_2995);
xnor U3093 (N_3093,N_2886,N_2894);
nand U3094 (N_3094,N_2994,N_2914);
nand U3095 (N_3095,N_2940,N_2983);
xor U3096 (N_3096,N_2818,N_2910);
nor U3097 (N_3097,N_2831,N_2976);
or U3098 (N_3098,N_2942,N_2944);
and U3099 (N_3099,N_2900,N_2806);
and U3100 (N_3100,N_2805,N_2893);
or U3101 (N_3101,N_2939,N_2937);
nand U3102 (N_3102,N_2962,N_2804);
xor U3103 (N_3103,N_2837,N_2889);
or U3104 (N_3104,N_2961,N_2827);
or U3105 (N_3105,N_2992,N_2957);
nand U3106 (N_3106,N_2995,N_2992);
and U3107 (N_3107,N_2840,N_2953);
xor U3108 (N_3108,N_2968,N_2996);
xnor U3109 (N_3109,N_2914,N_2875);
or U3110 (N_3110,N_2919,N_2807);
xor U3111 (N_3111,N_2967,N_2909);
nor U3112 (N_3112,N_2923,N_2918);
xnor U3113 (N_3113,N_2839,N_2946);
or U3114 (N_3114,N_2868,N_2992);
nand U3115 (N_3115,N_2888,N_2854);
nor U3116 (N_3116,N_2837,N_2817);
xnor U3117 (N_3117,N_2934,N_2904);
nand U3118 (N_3118,N_2839,N_2988);
nand U3119 (N_3119,N_2800,N_2920);
and U3120 (N_3120,N_2833,N_2819);
xor U3121 (N_3121,N_2923,N_2917);
or U3122 (N_3122,N_2840,N_2952);
and U3123 (N_3123,N_2960,N_2886);
or U3124 (N_3124,N_2911,N_2816);
or U3125 (N_3125,N_2908,N_2887);
and U3126 (N_3126,N_2847,N_2821);
nand U3127 (N_3127,N_2877,N_2977);
nand U3128 (N_3128,N_2880,N_2824);
and U3129 (N_3129,N_2938,N_2832);
and U3130 (N_3130,N_2922,N_2888);
nor U3131 (N_3131,N_2874,N_2971);
or U3132 (N_3132,N_2973,N_2928);
nor U3133 (N_3133,N_2902,N_2804);
and U3134 (N_3134,N_2875,N_2953);
xor U3135 (N_3135,N_2833,N_2905);
nand U3136 (N_3136,N_2903,N_2820);
or U3137 (N_3137,N_2805,N_2988);
or U3138 (N_3138,N_2857,N_2847);
xor U3139 (N_3139,N_2915,N_2972);
or U3140 (N_3140,N_2946,N_2940);
and U3141 (N_3141,N_2992,N_2876);
or U3142 (N_3142,N_2984,N_2968);
xor U3143 (N_3143,N_2818,N_2877);
or U3144 (N_3144,N_2898,N_2956);
nor U3145 (N_3145,N_2852,N_2973);
and U3146 (N_3146,N_2933,N_2865);
xor U3147 (N_3147,N_2988,N_2947);
nor U3148 (N_3148,N_2827,N_2963);
or U3149 (N_3149,N_2845,N_2825);
or U3150 (N_3150,N_2864,N_2959);
nand U3151 (N_3151,N_2902,N_2900);
nand U3152 (N_3152,N_2978,N_2998);
nand U3153 (N_3153,N_2903,N_2975);
or U3154 (N_3154,N_2892,N_2929);
xnor U3155 (N_3155,N_2873,N_2853);
or U3156 (N_3156,N_2844,N_2948);
or U3157 (N_3157,N_2955,N_2983);
nor U3158 (N_3158,N_2999,N_2951);
or U3159 (N_3159,N_2934,N_2989);
xor U3160 (N_3160,N_2909,N_2905);
nand U3161 (N_3161,N_2887,N_2994);
nor U3162 (N_3162,N_2942,N_2872);
nand U3163 (N_3163,N_2848,N_2840);
nand U3164 (N_3164,N_2954,N_2856);
nand U3165 (N_3165,N_2865,N_2966);
and U3166 (N_3166,N_2932,N_2949);
and U3167 (N_3167,N_2895,N_2896);
and U3168 (N_3168,N_2927,N_2800);
nor U3169 (N_3169,N_2919,N_2887);
nand U3170 (N_3170,N_2949,N_2867);
xnor U3171 (N_3171,N_2834,N_2976);
or U3172 (N_3172,N_2873,N_2880);
nand U3173 (N_3173,N_2860,N_2827);
xnor U3174 (N_3174,N_2845,N_2878);
and U3175 (N_3175,N_2924,N_2922);
or U3176 (N_3176,N_2816,N_2897);
xnor U3177 (N_3177,N_2909,N_2965);
nand U3178 (N_3178,N_2952,N_2814);
xnor U3179 (N_3179,N_2877,N_2939);
and U3180 (N_3180,N_2813,N_2823);
nand U3181 (N_3181,N_2821,N_2872);
nand U3182 (N_3182,N_2997,N_2830);
nand U3183 (N_3183,N_2910,N_2922);
nor U3184 (N_3184,N_2981,N_2938);
nand U3185 (N_3185,N_2972,N_2824);
nand U3186 (N_3186,N_2934,N_2906);
or U3187 (N_3187,N_2844,N_2975);
and U3188 (N_3188,N_2803,N_2851);
or U3189 (N_3189,N_2956,N_2910);
xor U3190 (N_3190,N_2965,N_2885);
and U3191 (N_3191,N_2862,N_2885);
nand U3192 (N_3192,N_2884,N_2832);
nor U3193 (N_3193,N_2975,N_2832);
nor U3194 (N_3194,N_2997,N_2928);
xnor U3195 (N_3195,N_2924,N_2879);
and U3196 (N_3196,N_2925,N_2809);
or U3197 (N_3197,N_2890,N_2938);
xnor U3198 (N_3198,N_2978,N_2909);
xor U3199 (N_3199,N_2927,N_2996);
nor U3200 (N_3200,N_3029,N_3127);
and U3201 (N_3201,N_3084,N_3147);
xor U3202 (N_3202,N_3038,N_3122);
xor U3203 (N_3203,N_3021,N_3003);
or U3204 (N_3204,N_3106,N_3110);
and U3205 (N_3205,N_3009,N_3166);
and U3206 (N_3206,N_3102,N_3027);
and U3207 (N_3207,N_3082,N_3019);
nor U3208 (N_3208,N_3006,N_3103);
nand U3209 (N_3209,N_3061,N_3186);
and U3210 (N_3210,N_3070,N_3154);
or U3211 (N_3211,N_3077,N_3173);
and U3212 (N_3212,N_3091,N_3044);
xnor U3213 (N_3213,N_3025,N_3118);
and U3214 (N_3214,N_3020,N_3151);
xnor U3215 (N_3215,N_3133,N_3159);
xor U3216 (N_3216,N_3040,N_3036);
or U3217 (N_3217,N_3113,N_3011);
or U3218 (N_3218,N_3188,N_3046);
nor U3219 (N_3219,N_3041,N_3194);
or U3220 (N_3220,N_3042,N_3178);
or U3221 (N_3221,N_3049,N_3158);
xor U3222 (N_3222,N_3071,N_3139);
or U3223 (N_3223,N_3123,N_3179);
nand U3224 (N_3224,N_3004,N_3140);
xnor U3225 (N_3225,N_3191,N_3066);
and U3226 (N_3226,N_3030,N_3115);
or U3227 (N_3227,N_3086,N_3169);
nand U3228 (N_3228,N_3056,N_3051);
or U3229 (N_3229,N_3058,N_3120);
nand U3230 (N_3230,N_3063,N_3007);
xor U3231 (N_3231,N_3012,N_3059);
or U3232 (N_3232,N_3095,N_3187);
or U3233 (N_3233,N_3176,N_3002);
and U3234 (N_3234,N_3060,N_3050);
nor U3235 (N_3235,N_3013,N_3161);
nor U3236 (N_3236,N_3185,N_3093);
or U3237 (N_3237,N_3190,N_3101);
nand U3238 (N_3238,N_3068,N_3171);
and U3239 (N_3239,N_3144,N_3016);
and U3240 (N_3240,N_3045,N_3163);
xnor U3241 (N_3241,N_3145,N_3132);
xnor U3242 (N_3242,N_3097,N_3087);
or U3243 (N_3243,N_3034,N_3054);
and U3244 (N_3244,N_3150,N_3053);
and U3245 (N_3245,N_3043,N_3094);
xnor U3246 (N_3246,N_3064,N_3170);
and U3247 (N_3247,N_3117,N_3076);
xnor U3248 (N_3248,N_3081,N_3080);
or U3249 (N_3249,N_3000,N_3174);
nor U3250 (N_3250,N_3099,N_3177);
nand U3251 (N_3251,N_3073,N_3198);
nor U3252 (N_3252,N_3183,N_3130);
or U3253 (N_3253,N_3114,N_3121);
and U3254 (N_3254,N_3105,N_3155);
nor U3255 (N_3255,N_3098,N_3075);
nor U3256 (N_3256,N_3037,N_3181);
nor U3257 (N_3257,N_3039,N_3109);
xor U3258 (N_3258,N_3078,N_3138);
and U3259 (N_3259,N_3189,N_3143);
nand U3260 (N_3260,N_3172,N_3195);
or U3261 (N_3261,N_3065,N_3196);
nor U3262 (N_3262,N_3135,N_3014);
or U3263 (N_3263,N_3052,N_3033);
or U3264 (N_3264,N_3074,N_3085);
and U3265 (N_3265,N_3197,N_3015);
nand U3266 (N_3266,N_3108,N_3026);
nand U3267 (N_3267,N_3125,N_3112);
nand U3268 (N_3268,N_3035,N_3156);
nand U3269 (N_3269,N_3146,N_3090);
nor U3270 (N_3270,N_3164,N_3116);
nor U3271 (N_3271,N_3079,N_3023);
and U3272 (N_3272,N_3168,N_3124);
or U3273 (N_3273,N_3089,N_3031);
and U3274 (N_3274,N_3100,N_3005);
nor U3275 (N_3275,N_3129,N_3157);
nor U3276 (N_3276,N_3184,N_3111);
or U3277 (N_3277,N_3008,N_3119);
and U3278 (N_3278,N_3131,N_3141);
nand U3279 (N_3279,N_3057,N_3022);
nor U3280 (N_3280,N_3092,N_3175);
xnor U3281 (N_3281,N_3162,N_3149);
nand U3282 (N_3282,N_3126,N_3010);
or U3283 (N_3283,N_3048,N_3137);
xnor U3284 (N_3284,N_3001,N_3062);
nand U3285 (N_3285,N_3180,N_3193);
nand U3286 (N_3286,N_3104,N_3182);
nor U3287 (N_3287,N_3024,N_3055);
nor U3288 (N_3288,N_3136,N_3107);
nand U3289 (N_3289,N_3165,N_3032);
nand U3290 (N_3290,N_3128,N_3199);
and U3291 (N_3291,N_3152,N_3153);
nor U3292 (N_3292,N_3083,N_3167);
and U3293 (N_3293,N_3069,N_3072);
xnor U3294 (N_3294,N_3160,N_3088);
nand U3295 (N_3295,N_3096,N_3142);
nand U3296 (N_3296,N_3047,N_3192);
nand U3297 (N_3297,N_3134,N_3018);
nor U3298 (N_3298,N_3067,N_3148);
nand U3299 (N_3299,N_3017,N_3028);
or U3300 (N_3300,N_3168,N_3103);
xnor U3301 (N_3301,N_3027,N_3035);
nor U3302 (N_3302,N_3194,N_3092);
or U3303 (N_3303,N_3038,N_3175);
or U3304 (N_3304,N_3142,N_3125);
xnor U3305 (N_3305,N_3193,N_3130);
or U3306 (N_3306,N_3139,N_3010);
or U3307 (N_3307,N_3072,N_3152);
nor U3308 (N_3308,N_3114,N_3108);
nand U3309 (N_3309,N_3039,N_3030);
and U3310 (N_3310,N_3197,N_3010);
xnor U3311 (N_3311,N_3068,N_3007);
or U3312 (N_3312,N_3179,N_3009);
nor U3313 (N_3313,N_3122,N_3024);
xor U3314 (N_3314,N_3169,N_3050);
nor U3315 (N_3315,N_3171,N_3096);
xor U3316 (N_3316,N_3088,N_3148);
and U3317 (N_3317,N_3034,N_3000);
or U3318 (N_3318,N_3190,N_3019);
xnor U3319 (N_3319,N_3148,N_3022);
or U3320 (N_3320,N_3196,N_3188);
xnor U3321 (N_3321,N_3113,N_3031);
nand U3322 (N_3322,N_3049,N_3163);
nor U3323 (N_3323,N_3074,N_3025);
nor U3324 (N_3324,N_3054,N_3189);
and U3325 (N_3325,N_3164,N_3195);
nand U3326 (N_3326,N_3192,N_3051);
and U3327 (N_3327,N_3032,N_3128);
nand U3328 (N_3328,N_3170,N_3075);
nor U3329 (N_3329,N_3183,N_3088);
or U3330 (N_3330,N_3017,N_3158);
and U3331 (N_3331,N_3088,N_3035);
nand U3332 (N_3332,N_3145,N_3073);
xnor U3333 (N_3333,N_3049,N_3065);
or U3334 (N_3334,N_3180,N_3199);
and U3335 (N_3335,N_3185,N_3189);
nor U3336 (N_3336,N_3020,N_3034);
nor U3337 (N_3337,N_3100,N_3121);
nor U3338 (N_3338,N_3190,N_3161);
nand U3339 (N_3339,N_3153,N_3018);
nand U3340 (N_3340,N_3166,N_3078);
or U3341 (N_3341,N_3197,N_3178);
xnor U3342 (N_3342,N_3055,N_3145);
xor U3343 (N_3343,N_3133,N_3033);
nand U3344 (N_3344,N_3186,N_3028);
or U3345 (N_3345,N_3081,N_3121);
nand U3346 (N_3346,N_3181,N_3154);
or U3347 (N_3347,N_3089,N_3180);
and U3348 (N_3348,N_3094,N_3061);
nor U3349 (N_3349,N_3012,N_3187);
and U3350 (N_3350,N_3146,N_3117);
and U3351 (N_3351,N_3126,N_3074);
nand U3352 (N_3352,N_3100,N_3119);
nor U3353 (N_3353,N_3065,N_3013);
nand U3354 (N_3354,N_3030,N_3000);
nand U3355 (N_3355,N_3023,N_3046);
and U3356 (N_3356,N_3156,N_3105);
xnor U3357 (N_3357,N_3170,N_3101);
nand U3358 (N_3358,N_3086,N_3120);
or U3359 (N_3359,N_3030,N_3097);
nand U3360 (N_3360,N_3040,N_3138);
nand U3361 (N_3361,N_3199,N_3045);
or U3362 (N_3362,N_3043,N_3025);
or U3363 (N_3363,N_3151,N_3027);
and U3364 (N_3364,N_3131,N_3014);
and U3365 (N_3365,N_3101,N_3075);
nand U3366 (N_3366,N_3081,N_3195);
nor U3367 (N_3367,N_3091,N_3142);
and U3368 (N_3368,N_3051,N_3087);
and U3369 (N_3369,N_3038,N_3130);
or U3370 (N_3370,N_3023,N_3029);
nor U3371 (N_3371,N_3143,N_3102);
nand U3372 (N_3372,N_3019,N_3097);
xor U3373 (N_3373,N_3147,N_3002);
or U3374 (N_3374,N_3099,N_3189);
and U3375 (N_3375,N_3101,N_3063);
nand U3376 (N_3376,N_3144,N_3149);
nand U3377 (N_3377,N_3094,N_3196);
nand U3378 (N_3378,N_3063,N_3137);
or U3379 (N_3379,N_3087,N_3110);
or U3380 (N_3380,N_3080,N_3079);
and U3381 (N_3381,N_3166,N_3100);
and U3382 (N_3382,N_3080,N_3194);
or U3383 (N_3383,N_3090,N_3127);
and U3384 (N_3384,N_3002,N_3104);
xnor U3385 (N_3385,N_3148,N_3166);
nand U3386 (N_3386,N_3045,N_3122);
or U3387 (N_3387,N_3098,N_3065);
or U3388 (N_3388,N_3089,N_3080);
or U3389 (N_3389,N_3128,N_3188);
xor U3390 (N_3390,N_3008,N_3063);
nor U3391 (N_3391,N_3190,N_3189);
nand U3392 (N_3392,N_3094,N_3163);
or U3393 (N_3393,N_3141,N_3135);
or U3394 (N_3394,N_3152,N_3186);
nand U3395 (N_3395,N_3066,N_3029);
and U3396 (N_3396,N_3163,N_3101);
and U3397 (N_3397,N_3025,N_3135);
xnor U3398 (N_3398,N_3124,N_3008);
and U3399 (N_3399,N_3129,N_3021);
xnor U3400 (N_3400,N_3288,N_3389);
or U3401 (N_3401,N_3323,N_3361);
nor U3402 (N_3402,N_3303,N_3321);
or U3403 (N_3403,N_3229,N_3248);
nand U3404 (N_3404,N_3234,N_3262);
and U3405 (N_3405,N_3383,N_3271);
nand U3406 (N_3406,N_3379,N_3336);
or U3407 (N_3407,N_3284,N_3231);
xor U3408 (N_3408,N_3382,N_3224);
and U3409 (N_3409,N_3399,N_3283);
and U3410 (N_3410,N_3264,N_3245);
nor U3411 (N_3411,N_3255,N_3330);
xnor U3412 (N_3412,N_3362,N_3356);
nor U3413 (N_3413,N_3228,N_3393);
and U3414 (N_3414,N_3285,N_3201);
or U3415 (N_3415,N_3225,N_3392);
nor U3416 (N_3416,N_3265,N_3202);
nand U3417 (N_3417,N_3390,N_3360);
nand U3418 (N_3418,N_3378,N_3259);
or U3419 (N_3419,N_3354,N_3205);
xnor U3420 (N_3420,N_3329,N_3312);
nor U3421 (N_3421,N_3351,N_3344);
and U3422 (N_3422,N_3310,N_3366);
or U3423 (N_3423,N_3297,N_3396);
nand U3424 (N_3424,N_3219,N_3308);
nor U3425 (N_3425,N_3215,N_3217);
and U3426 (N_3426,N_3306,N_3302);
xnor U3427 (N_3427,N_3358,N_3391);
or U3428 (N_3428,N_3221,N_3200);
nor U3429 (N_3429,N_3258,N_3307);
and U3430 (N_3430,N_3220,N_3289);
nor U3431 (N_3431,N_3273,N_3210);
and U3432 (N_3432,N_3328,N_3387);
nor U3433 (N_3433,N_3233,N_3287);
nor U3434 (N_3434,N_3216,N_3236);
xor U3435 (N_3435,N_3278,N_3300);
nor U3436 (N_3436,N_3293,N_3213);
and U3437 (N_3437,N_3296,N_3277);
xor U3438 (N_3438,N_3397,N_3208);
nor U3439 (N_3439,N_3367,N_3280);
or U3440 (N_3440,N_3207,N_3291);
xor U3441 (N_3441,N_3334,N_3230);
nand U3442 (N_3442,N_3333,N_3279);
nor U3443 (N_3443,N_3286,N_3365);
xor U3444 (N_3444,N_3342,N_3348);
xor U3445 (N_3445,N_3212,N_3359);
or U3446 (N_3446,N_3341,N_3332);
and U3447 (N_3447,N_3240,N_3272);
and U3448 (N_3448,N_3314,N_3320);
and U3449 (N_3449,N_3270,N_3276);
nand U3450 (N_3450,N_3395,N_3261);
or U3451 (N_3451,N_3385,N_3326);
nand U3452 (N_3452,N_3305,N_3246);
or U3453 (N_3453,N_3352,N_3238);
nand U3454 (N_3454,N_3347,N_3239);
nor U3455 (N_3455,N_3384,N_3313);
and U3456 (N_3456,N_3337,N_3325);
nor U3457 (N_3457,N_3223,N_3232);
xor U3458 (N_3458,N_3357,N_3298);
or U3459 (N_3459,N_3204,N_3263);
nor U3460 (N_3460,N_3251,N_3311);
nor U3461 (N_3461,N_3398,N_3243);
or U3462 (N_3462,N_3275,N_3376);
xnor U3463 (N_3463,N_3252,N_3335);
xor U3464 (N_3464,N_3250,N_3260);
and U3465 (N_3465,N_3350,N_3373);
and U3466 (N_3466,N_3237,N_3209);
nor U3467 (N_3467,N_3331,N_3317);
xnor U3468 (N_3468,N_3309,N_3214);
nand U3469 (N_3469,N_3368,N_3206);
or U3470 (N_3470,N_3294,N_3247);
nand U3471 (N_3471,N_3227,N_3338);
or U3472 (N_3472,N_3340,N_3327);
nand U3473 (N_3473,N_3295,N_3290);
nand U3474 (N_3474,N_3241,N_3253);
nand U3475 (N_3475,N_3203,N_3242);
or U3476 (N_3476,N_3380,N_3257);
xor U3477 (N_3477,N_3364,N_3304);
nand U3478 (N_3478,N_3211,N_3343);
or U3479 (N_3479,N_3381,N_3281);
nand U3480 (N_3480,N_3339,N_3244);
and U3481 (N_3481,N_3299,N_3319);
and U3482 (N_3482,N_3375,N_3256);
and U3483 (N_3483,N_3267,N_3218);
and U3484 (N_3484,N_3353,N_3226);
and U3485 (N_3485,N_3316,N_3254);
nand U3486 (N_3486,N_3249,N_3388);
nand U3487 (N_3487,N_3315,N_3370);
xnor U3488 (N_3488,N_3372,N_3324);
xor U3489 (N_3489,N_3346,N_3269);
nand U3490 (N_3490,N_3363,N_3274);
nand U3491 (N_3491,N_3322,N_3377);
nand U3492 (N_3492,N_3292,N_3222);
nand U3493 (N_3493,N_3394,N_3266);
or U3494 (N_3494,N_3235,N_3349);
or U3495 (N_3495,N_3282,N_3301);
or U3496 (N_3496,N_3369,N_3355);
xor U3497 (N_3497,N_3371,N_3318);
xnor U3498 (N_3498,N_3386,N_3345);
and U3499 (N_3499,N_3374,N_3268);
nor U3500 (N_3500,N_3260,N_3357);
xor U3501 (N_3501,N_3346,N_3278);
nand U3502 (N_3502,N_3346,N_3220);
xor U3503 (N_3503,N_3323,N_3242);
xnor U3504 (N_3504,N_3211,N_3259);
nand U3505 (N_3505,N_3228,N_3300);
and U3506 (N_3506,N_3337,N_3232);
nand U3507 (N_3507,N_3322,N_3211);
or U3508 (N_3508,N_3355,N_3343);
nor U3509 (N_3509,N_3299,N_3364);
nor U3510 (N_3510,N_3342,N_3249);
nand U3511 (N_3511,N_3254,N_3213);
nor U3512 (N_3512,N_3322,N_3392);
nand U3513 (N_3513,N_3353,N_3210);
nand U3514 (N_3514,N_3358,N_3333);
nor U3515 (N_3515,N_3304,N_3263);
nand U3516 (N_3516,N_3388,N_3314);
xnor U3517 (N_3517,N_3293,N_3209);
or U3518 (N_3518,N_3269,N_3304);
nor U3519 (N_3519,N_3323,N_3246);
xnor U3520 (N_3520,N_3303,N_3218);
or U3521 (N_3521,N_3288,N_3234);
xnor U3522 (N_3522,N_3264,N_3269);
and U3523 (N_3523,N_3267,N_3328);
and U3524 (N_3524,N_3319,N_3242);
nor U3525 (N_3525,N_3232,N_3238);
xor U3526 (N_3526,N_3291,N_3284);
or U3527 (N_3527,N_3334,N_3355);
and U3528 (N_3528,N_3346,N_3395);
or U3529 (N_3529,N_3231,N_3202);
and U3530 (N_3530,N_3388,N_3280);
nor U3531 (N_3531,N_3254,N_3313);
xor U3532 (N_3532,N_3338,N_3373);
nor U3533 (N_3533,N_3259,N_3380);
xor U3534 (N_3534,N_3354,N_3242);
xor U3535 (N_3535,N_3244,N_3243);
or U3536 (N_3536,N_3267,N_3260);
or U3537 (N_3537,N_3241,N_3326);
nor U3538 (N_3538,N_3323,N_3266);
xnor U3539 (N_3539,N_3241,N_3345);
or U3540 (N_3540,N_3372,N_3362);
nand U3541 (N_3541,N_3272,N_3238);
nand U3542 (N_3542,N_3352,N_3207);
or U3543 (N_3543,N_3215,N_3332);
or U3544 (N_3544,N_3240,N_3281);
and U3545 (N_3545,N_3349,N_3287);
xor U3546 (N_3546,N_3331,N_3349);
xnor U3547 (N_3547,N_3263,N_3305);
or U3548 (N_3548,N_3209,N_3228);
nand U3549 (N_3549,N_3361,N_3327);
and U3550 (N_3550,N_3325,N_3355);
or U3551 (N_3551,N_3223,N_3343);
xor U3552 (N_3552,N_3327,N_3373);
nor U3553 (N_3553,N_3237,N_3338);
nand U3554 (N_3554,N_3243,N_3271);
nand U3555 (N_3555,N_3261,N_3243);
or U3556 (N_3556,N_3209,N_3373);
or U3557 (N_3557,N_3368,N_3372);
or U3558 (N_3558,N_3346,N_3392);
nor U3559 (N_3559,N_3305,N_3359);
and U3560 (N_3560,N_3202,N_3222);
nor U3561 (N_3561,N_3358,N_3319);
nor U3562 (N_3562,N_3382,N_3204);
nand U3563 (N_3563,N_3295,N_3322);
xnor U3564 (N_3564,N_3365,N_3228);
and U3565 (N_3565,N_3295,N_3362);
xor U3566 (N_3566,N_3234,N_3305);
and U3567 (N_3567,N_3268,N_3222);
xor U3568 (N_3568,N_3244,N_3270);
nand U3569 (N_3569,N_3398,N_3321);
and U3570 (N_3570,N_3375,N_3355);
nand U3571 (N_3571,N_3238,N_3268);
nor U3572 (N_3572,N_3327,N_3213);
or U3573 (N_3573,N_3258,N_3249);
and U3574 (N_3574,N_3364,N_3260);
nand U3575 (N_3575,N_3342,N_3256);
nor U3576 (N_3576,N_3268,N_3278);
or U3577 (N_3577,N_3343,N_3201);
and U3578 (N_3578,N_3372,N_3329);
nor U3579 (N_3579,N_3204,N_3217);
nand U3580 (N_3580,N_3343,N_3375);
or U3581 (N_3581,N_3279,N_3209);
xnor U3582 (N_3582,N_3368,N_3243);
nor U3583 (N_3583,N_3329,N_3313);
and U3584 (N_3584,N_3296,N_3397);
or U3585 (N_3585,N_3275,N_3308);
nand U3586 (N_3586,N_3285,N_3304);
nand U3587 (N_3587,N_3200,N_3285);
nand U3588 (N_3588,N_3239,N_3305);
and U3589 (N_3589,N_3279,N_3307);
xnor U3590 (N_3590,N_3261,N_3251);
xor U3591 (N_3591,N_3385,N_3348);
or U3592 (N_3592,N_3356,N_3211);
and U3593 (N_3593,N_3358,N_3267);
xnor U3594 (N_3594,N_3240,N_3250);
and U3595 (N_3595,N_3232,N_3336);
nor U3596 (N_3596,N_3337,N_3334);
xor U3597 (N_3597,N_3313,N_3383);
or U3598 (N_3598,N_3294,N_3391);
xnor U3599 (N_3599,N_3232,N_3237);
nand U3600 (N_3600,N_3592,N_3475);
or U3601 (N_3601,N_3406,N_3501);
or U3602 (N_3602,N_3534,N_3476);
or U3603 (N_3603,N_3550,N_3429);
xor U3604 (N_3604,N_3559,N_3434);
nand U3605 (N_3605,N_3486,N_3439);
nand U3606 (N_3606,N_3588,N_3479);
nor U3607 (N_3607,N_3535,N_3504);
xnor U3608 (N_3608,N_3503,N_3453);
xnor U3609 (N_3609,N_3540,N_3482);
nor U3610 (N_3610,N_3594,N_3548);
and U3611 (N_3611,N_3510,N_3581);
nor U3612 (N_3612,N_3575,N_3539);
or U3613 (N_3613,N_3502,N_3564);
nand U3614 (N_3614,N_3425,N_3473);
or U3615 (N_3615,N_3537,N_3565);
nand U3616 (N_3616,N_3527,N_3428);
and U3617 (N_3617,N_3528,N_3420);
nor U3618 (N_3618,N_3493,N_3487);
and U3619 (N_3619,N_3505,N_3485);
nor U3620 (N_3620,N_3508,N_3579);
and U3621 (N_3621,N_3595,N_3597);
nor U3622 (N_3622,N_3571,N_3468);
nor U3623 (N_3623,N_3496,N_3526);
xor U3624 (N_3624,N_3408,N_3586);
xnor U3625 (N_3625,N_3438,N_3415);
nor U3626 (N_3626,N_3490,N_3531);
xnor U3627 (N_3627,N_3402,N_3462);
or U3628 (N_3628,N_3566,N_3536);
and U3629 (N_3629,N_3511,N_3497);
and U3630 (N_3630,N_3585,N_3444);
and U3631 (N_3631,N_3584,N_3523);
or U3632 (N_3632,N_3498,N_3403);
nor U3633 (N_3633,N_3541,N_3572);
or U3634 (N_3634,N_3587,N_3472);
or U3635 (N_3635,N_3495,N_3546);
xnor U3636 (N_3636,N_3449,N_3448);
or U3637 (N_3637,N_3570,N_3405);
xnor U3638 (N_3638,N_3421,N_3418);
nor U3639 (N_3639,N_3517,N_3513);
or U3640 (N_3640,N_3443,N_3480);
nor U3641 (N_3641,N_3404,N_3542);
and U3642 (N_3642,N_3471,N_3436);
xor U3643 (N_3643,N_3488,N_3477);
nor U3644 (N_3644,N_3437,N_3562);
nand U3645 (N_3645,N_3481,N_3553);
nor U3646 (N_3646,N_3409,N_3529);
or U3647 (N_3647,N_3569,N_3442);
nor U3648 (N_3648,N_3491,N_3589);
nand U3649 (N_3649,N_3593,N_3568);
xnor U3650 (N_3650,N_3576,N_3544);
nand U3651 (N_3651,N_3560,N_3555);
xor U3652 (N_3652,N_3474,N_3557);
nand U3653 (N_3653,N_3543,N_3547);
nand U3654 (N_3654,N_3552,N_3411);
or U3655 (N_3655,N_3596,N_3525);
nor U3656 (N_3656,N_3469,N_3466);
nand U3657 (N_3657,N_3483,N_3431);
or U3658 (N_3658,N_3426,N_3478);
and U3659 (N_3659,N_3538,N_3450);
or U3660 (N_3660,N_3407,N_3412);
and U3661 (N_3661,N_3573,N_3530);
nor U3662 (N_3662,N_3512,N_3556);
xor U3663 (N_3663,N_3577,N_3457);
nand U3664 (N_3664,N_3598,N_3467);
or U3665 (N_3665,N_3563,N_3509);
and U3666 (N_3666,N_3400,N_3551);
and U3667 (N_3667,N_3401,N_3451);
or U3668 (N_3668,N_3424,N_3516);
and U3669 (N_3669,N_3514,N_3545);
xnor U3670 (N_3670,N_3427,N_3574);
and U3671 (N_3671,N_3567,N_3549);
or U3672 (N_3672,N_3422,N_3447);
and U3673 (N_3673,N_3489,N_3441);
and U3674 (N_3674,N_3590,N_3519);
and U3675 (N_3675,N_3432,N_3518);
and U3676 (N_3676,N_3532,N_3463);
nand U3677 (N_3677,N_3515,N_3419);
and U3678 (N_3678,N_3460,N_3520);
or U3679 (N_3679,N_3413,N_3458);
nand U3680 (N_3680,N_3446,N_3484);
or U3681 (N_3681,N_3452,N_3455);
xor U3682 (N_3682,N_3522,N_3456);
nor U3683 (N_3683,N_3464,N_3561);
or U3684 (N_3684,N_3494,N_3533);
nand U3685 (N_3685,N_3454,N_3554);
xor U3686 (N_3686,N_3583,N_3521);
and U3687 (N_3687,N_3492,N_3416);
xnor U3688 (N_3688,N_3410,N_3445);
xnor U3689 (N_3689,N_3461,N_3558);
or U3690 (N_3690,N_3580,N_3417);
and U3691 (N_3691,N_3506,N_3507);
nor U3692 (N_3692,N_3500,N_3582);
or U3693 (N_3693,N_3599,N_3423);
and U3694 (N_3694,N_3499,N_3440);
xnor U3695 (N_3695,N_3465,N_3524);
or U3696 (N_3696,N_3414,N_3435);
nor U3697 (N_3697,N_3459,N_3578);
nor U3698 (N_3698,N_3591,N_3430);
nor U3699 (N_3699,N_3433,N_3470);
xor U3700 (N_3700,N_3588,N_3516);
xnor U3701 (N_3701,N_3553,N_3513);
xor U3702 (N_3702,N_3455,N_3557);
or U3703 (N_3703,N_3492,N_3531);
and U3704 (N_3704,N_3451,N_3452);
nor U3705 (N_3705,N_3582,N_3548);
and U3706 (N_3706,N_3547,N_3454);
nand U3707 (N_3707,N_3520,N_3434);
or U3708 (N_3708,N_3451,N_3457);
or U3709 (N_3709,N_3424,N_3463);
nand U3710 (N_3710,N_3591,N_3472);
nand U3711 (N_3711,N_3590,N_3451);
nor U3712 (N_3712,N_3491,N_3526);
or U3713 (N_3713,N_3539,N_3598);
xnor U3714 (N_3714,N_3476,N_3438);
or U3715 (N_3715,N_3582,N_3440);
nand U3716 (N_3716,N_3531,N_3560);
nor U3717 (N_3717,N_3556,N_3597);
xor U3718 (N_3718,N_3550,N_3578);
nand U3719 (N_3719,N_3595,N_3451);
nand U3720 (N_3720,N_3511,N_3589);
nor U3721 (N_3721,N_3570,N_3453);
nor U3722 (N_3722,N_3435,N_3495);
and U3723 (N_3723,N_3562,N_3430);
or U3724 (N_3724,N_3472,N_3492);
nor U3725 (N_3725,N_3577,N_3426);
or U3726 (N_3726,N_3466,N_3560);
and U3727 (N_3727,N_3425,N_3431);
or U3728 (N_3728,N_3409,N_3455);
or U3729 (N_3729,N_3498,N_3580);
nor U3730 (N_3730,N_3475,N_3419);
or U3731 (N_3731,N_3444,N_3438);
and U3732 (N_3732,N_3471,N_3535);
nand U3733 (N_3733,N_3498,N_3538);
xnor U3734 (N_3734,N_3547,N_3421);
nor U3735 (N_3735,N_3442,N_3590);
and U3736 (N_3736,N_3435,N_3547);
and U3737 (N_3737,N_3554,N_3581);
xor U3738 (N_3738,N_3446,N_3406);
or U3739 (N_3739,N_3582,N_3505);
xnor U3740 (N_3740,N_3521,N_3497);
nand U3741 (N_3741,N_3408,N_3500);
and U3742 (N_3742,N_3479,N_3599);
xor U3743 (N_3743,N_3585,N_3418);
or U3744 (N_3744,N_3489,N_3550);
nor U3745 (N_3745,N_3552,N_3413);
and U3746 (N_3746,N_3419,N_3402);
nor U3747 (N_3747,N_3565,N_3445);
and U3748 (N_3748,N_3414,N_3484);
xnor U3749 (N_3749,N_3430,N_3576);
nand U3750 (N_3750,N_3532,N_3422);
or U3751 (N_3751,N_3437,N_3440);
or U3752 (N_3752,N_3541,N_3495);
nor U3753 (N_3753,N_3498,N_3581);
and U3754 (N_3754,N_3414,N_3553);
xor U3755 (N_3755,N_3528,N_3401);
nor U3756 (N_3756,N_3410,N_3547);
xor U3757 (N_3757,N_3512,N_3543);
nand U3758 (N_3758,N_3458,N_3425);
xor U3759 (N_3759,N_3470,N_3467);
nor U3760 (N_3760,N_3444,N_3485);
or U3761 (N_3761,N_3555,N_3481);
or U3762 (N_3762,N_3462,N_3474);
xnor U3763 (N_3763,N_3523,N_3504);
nor U3764 (N_3764,N_3482,N_3550);
and U3765 (N_3765,N_3502,N_3547);
and U3766 (N_3766,N_3435,N_3474);
or U3767 (N_3767,N_3524,N_3412);
nor U3768 (N_3768,N_3493,N_3422);
nand U3769 (N_3769,N_3523,N_3510);
nor U3770 (N_3770,N_3444,N_3548);
and U3771 (N_3771,N_3534,N_3494);
or U3772 (N_3772,N_3561,N_3429);
or U3773 (N_3773,N_3475,N_3481);
xor U3774 (N_3774,N_3511,N_3449);
nand U3775 (N_3775,N_3419,N_3467);
or U3776 (N_3776,N_3546,N_3551);
nand U3777 (N_3777,N_3504,N_3415);
nand U3778 (N_3778,N_3518,N_3492);
nand U3779 (N_3779,N_3406,N_3452);
xor U3780 (N_3780,N_3554,N_3586);
or U3781 (N_3781,N_3486,N_3595);
nor U3782 (N_3782,N_3493,N_3506);
nand U3783 (N_3783,N_3461,N_3576);
or U3784 (N_3784,N_3485,N_3413);
or U3785 (N_3785,N_3403,N_3558);
and U3786 (N_3786,N_3456,N_3476);
xor U3787 (N_3787,N_3488,N_3494);
and U3788 (N_3788,N_3508,N_3462);
and U3789 (N_3789,N_3495,N_3444);
nor U3790 (N_3790,N_3479,N_3521);
nor U3791 (N_3791,N_3460,N_3477);
nand U3792 (N_3792,N_3492,N_3549);
or U3793 (N_3793,N_3536,N_3546);
or U3794 (N_3794,N_3408,N_3494);
nor U3795 (N_3795,N_3581,N_3549);
or U3796 (N_3796,N_3595,N_3481);
xor U3797 (N_3797,N_3443,N_3429);
or U3798 (N_3798,N_3493,N_3410);
or U3799 (N_3799,N_3469,N_3419);
nor U3800 (N_3800,N_3726,N_3631);
xnor U3801 (N_3801,N_3691,N_3759);
xnor U3802 (N_3802,N_3633,N_3790);
or U3803 (N_3803,N_3650,N_3752);
and U3804 (N_3804,N_3601,N_3714);
xnor U3805 (N_3805,N_3765,N_3782);
nand U3806 (N_3806,N_3732,N_3699);
nand U3807 (N_3807,N_3705,N_3624);
and U3808 (N_3808,N_3763,N_3674);
nor U3809 (N_3809,N_3670,N_3608);
nor U3810 (N_3810,N_3652,N_3687);
nand U3811 (N_3811,N_3700,N_3671);
or U3812 (N_3812,N_3749,N_3640);
nor U3813 (N_3813,N_3792,N_3745);
nor U3814 (N_3814,N_3753,N_3647);
nor U3815 (N_3815,N_3764,N_3701);
xor U3816 (N_3816,N_3612,N_3794);
nand U3817 (N_3817,N_3657,N_3659);
xor U3818 (N_3818,N_3731,N_3677);
and U3819 (N_3819,N_3791,N_3754);
nand U3820 (N_3820,N_3716,N_3751);
nor U3821 (N_3821,N_3773,N_3797);
nand U3822 (N_3822,N_3696,N_3686);
nor U3823 (N_3823,N_3741,N_3621);
or U3824 (N_3824,N_3638,N_3632);
and U3825 (N_3825,N_3643,N_3747);
nand U3826 (N_3826,N_3793,N_3679);
nor U3827 (N_3827,N_3762,N_3777);
xnor U3828 (N_3828,N_3708,N_3680);
nand U3829 (N_3829,N_3746,N_3727);
nand U3830 (N_3830,N_3799,N_3798);
nand U3831 (N_3831,N_3616,N_3786);
nand U3832 (N_3832,N_3618,N_3723);
nor U3833 (N_3833,N_3689,N_3766);
nor U3834 (N_3834,N_3738,N_3703);
nor U3835 (N_3835,N_3636,N_3669);
or U3836 (N_3836,N_3779,N_3729);
nand U3837 (N_3837,N_3625,N_3718);
nor U3838 (N_3838,N_3715,N_3644);
xor U3839 (N_3839,N_3774,N_3663);
nand U3840 (N_3840,N_3645,N_3617);
nor U3841 (N_3841,N_3653,N_3622);
xor U3842 (N_3842,N_3690,N_3771);
nand U3843 (N_3843,N_3743,N_3744);
and U3844 (N_3844,N_3675,N_3755);
nand U3845 (N_3845,N_3613,N_3694);
or U3846 (N_3846,N_3628,N_3626);
nor U3847 (N_3847,N_3681,N_3728);
nand U3848 (N_3848,N_3783,N_3610);
nor U3849 (N_3849,N_3627,N_3717);
nor U3850 (N_3850,N_3767,N_3619);
xnor U3851 (N_3851,N_3684,N_3721);
and U3852 (N_3852,N_3634,N_3615);
nor U3853 (N_3853,N_3688,N_3676);
and U3854 (N_3854,N_3656,N_3602);
and U3855 (N_3855,N_3736,N_3611);
nor U3856 (N_3856,N_3713,N_3607);
nor U3857 (N_3857,N_3635,N_3666);
or U3858 (N_3858,N_3702,N_3685);
or U3859 (N_3859,N_3654,N_3682);
and U3860 (N_3860,N_3795,N_3665);
nor U3861 (N_3861,N_3646,N_3796);
or U3862 (N_3862,N_3664,N_3672);
or U3863 (N_3863,N_3735,N_3630);
nor U3864 (N_3864,N_3642,N_3768);
nor U3865 (N_3865,N_3648,N_3789);
and U3866 (N_3866,N_3707,N_3757);
nor U3867 (N_3867,N_3761,N_3600);
and U3868 (N_3868,N_3742,N_3734);
nand U3869 (N_3869,N_3649,N_3604);
nand U3870 (N_3870,N_3722,N_3712);
or U3871 (N_3871,N_3603,N_3673);
nor U3872 (N_3872,N_3606,N_3693);
or U3873 (N_3873,N_3695,N_3641);
nor U3874 (N_3874,N_3668,N_3623);
xnor U3875 (N_3875,N_3750,N_3724);
or U3876 (N_3876,N_3651,N_3758);
nand U3877 (N_3877,N_3748,N_3683);
nand U3878 (N_3878,N_3769,N_3737);
xor U3879 (N_3879,N_3775,N_3658);
or U3880 (N_3880,N_3637,N_3711);
or U3881 (N_3881,N_3706,N_3719);
nor U3882 (N_3882,N_3620,N_3787);
nor U3883 (N_3883,N_3678,N_3739);
and U3884 (N_3884,N_3639,N_3710);
or U3885 (N_3885,N_3772,N_3698);
xor U3886 (N_3886,N_3667,N_3660);
nor U3887 (N_3887,N_3740,N_3785);
and U3888 (N_3888,N_3730,N_3697);
xor U3889 (N_3889,N_3655,N_3788);
xnor U3890 (N_3890,N_3720,N_3609);
or U3891 (N_3891,N_3725,N_3709);
and U3892 (N_3892,N_3760,N_3784);
nand U3893 (N_3893,N_3780,N_3733);
or U3894 (N_3894,N_3781,N_3662);
and U3895 (N_3895,N_3776,N_3605);
xnor U3896 (N_3896,N_3770,N_3704);
nand U3897 (N_3897,N_3661,N_3756);
and U3898 (N_3898,N_3614,N_3778);
xnor U3899 (N_3899,N_3692,N_3629);
nand U3900 (N_3900,N_3642,N_3699);
nand U3901 (N_3901,N_3727,N_3678);
nand U3902 (N_3902,N_3736,N_3765);
or U3903 (N_3903,N_3672,N_3743);
or U3904 (N_3904,N_3774,N_3752);
xnor U3905 (N_3905,N_3716,N_3725);
and U3906 (N_3906,N_3667,N_3756);
nor U3907 (N_3907,N_3780,N_3799);
or U3908 (N_3908,N_3706,N_3726);
and U3909 (N_3909,N_3798,N_3769);
nor U3910 (N_3910,N_3788,N_3649);
and U3911 (N_3911,N_3617,N_3712);
nor U3912 (N_3912,N_3737,N_3605);
nor U3913 (N_3913,N_3637,N_3662);
or U3914 (N_3914,N_3736,N_3663);
xnor U3915 (N_3915,N_3761,N_3693);
or U3916 (N_3916,N_3713,N_3743);
or U3917 (N_3917,N_3782,N_3762);
xor U3918 (N_3918,N_3785,N_3630);
nor U3919 (N_3919,N_3761,N_3785);
or U3920 (N_3920,N_3762,N_3712);
nor U3921 (N_3921,N_3691,N_3704);
nand U3922 (N_3922,N_3730,N_3617);
or U3923 (N_3923,N_3634,N_3712);
and U3924 (N_3924,N_3653,N_3704);
or U3925 (N_3925,N_3625,N_3799);
nor U3926 (N_3926,N_3750,N_3651);
nand U3927 (N_3927,N_3657,N_3676);
xor U3928 (N_3928,N_3788,N_3787);
and U3929 (N_3929,N_3762,N_3736);
xnor U3930 (N_3930,N_3760,N_3775);
nor U3931 (N_3931,N_3621,N_3767);
xnor U3932 (N_3932,N_3672,N_3711);
xor U3933 (N_3933,N_3717,N_3776);
or U3934 (N_3934,N_3617,N_3735);
or U3935 (N_3935,N_3715,N_3776);
or U3936 (N_3936,N_3729,N_3798);
nand U3937 (N_3937,N_3702,N_3681);
or U3938 (N_3938,N_3610,N_3728);
and U3939 (N_3939,N_3775,N_3673);
nor U3940 (N_3940,N_3720,N_3707);
nor U3941 (N_3941,N_3790,N_3644);
and U3942 (N_3942,N_3635,N_3685);
xor U3943 (N_3943,N_3761,N_3725);
xor U3944 (N_3944,N_3708,N_3796);
nand U3945 (N_3945,N_3601,N_3603);
nand U3946 (N_3946,N_3663,N_3687);
nand U3947 (N_3947,N_3742,N_3757);
nand U3948 (N_3948,N_3652,N_3665);
or U3949 (N_3949,N_3716,N_3623);
and U3950 (N_3950,N_3681,N_3796);
nand U3951 (N_3951,N_3745,N_3717);
nor U3952 (N_3952,N_3772,N_3666);
or U3953 (N_3953,N_3611,N_3612);
nor U3954 (N_3954,N_3701,N_3629);
and U3955 (N_3955,N_3777,N_3758);
and U3956 (N_3956,N_3773,N_3771);
nor U3957 (N_3957,N_3619,N_3675);
or U3958 (N_3958,N_3770,N_3671);
and U3959 (N_3959,N_3797,N_3704);
nand U3960 (N_3960,N_3734,N_3704);
and U3961 (N_3961,N_3769,N_3771);
or U3962 (N_3962,N_3752,N_3607);
nor U3963 (N_3963,N_3663,N_3741);
nor U3964 (N_3964,N_3725,N_3655);
or U3965 (N_3965,N_3755,N_3678);
xor U3966 (N_3966,N_3778,N_3709);
or U3967 (N_3967,N_3706,N_3746);
or U3968 (N_3968,N_3672,N_3705);
and U3969 (N_3969,N_3702,N_3753);
and U3970 (N_3970,N_3761,N_3638);
nand U3971 (N_3971,N_3723,N_3713);
or U3972 (N_3972,N_3763,N_3798);
xor U3973 (N_3973,N_3742,N_3719);
xnor U3974 (N_3974,N_3671,N_3669);
nand U3975 (N_3975,N_3622,N_3607);
or U3976 (N_3976,N_3776,N_3603);
or U3977 (N_3977,N_3702,N_3757);
and U3978 (N_3978,N_3736,N_3628);
xnor U3979 (N_3979,N_3646,N_3773);
nor U3980 (N_3980,N_3685,N_3724);
and U3981 (N_3981,N_3735,N_3778);
or U3982 (N_3982,N_3648,N_3657);
and U3983 (N_3983,N_3664,N_3752);
nand U3984 (N_3984,N_3732,N_3779);
and U3985 (N_3985,N_3667,N_3733);
or U3986 (N_3986,N_3715,N_3696);
or U3987 (N_3987,N_3766,N_3606);
nand U3988 (N_3988,N_3666,N_3657);
and U3989 (N_3989,N_3764,N_3768);
and U3990 (N_3990,N_3660,N_3636);
and U3991 (N_3991,N_3672,N_3605);
and U3992 (N_3992,N_3723,N_3664);
and U3993 (N_3993,N_3693,N_3778);
and U3994 (N_3994,N_3652,N_3729);
and U3995 (N_3995,N_3623,N_3785);
and U3996 (N_3996,N_3698,N_3751);
and U3997 (N_3997,N_3668,N_3782);
nor U3998 (N_3998,N_3642,N_3676);
and U3999 (N_3999,N_3667,N_3609);
and U4000 (N_4000,N_3810,N_3919);
nor U4001 (N_4001,N_3830,N_3869);
nand U4002 (N_4002,N_3860,N_3958);
xor U4003 (N_4003,N_3903,N_3970);
nor U4004 (N_4004,N_3898,N_3972);
nor U4005 (N_4005,N_3896,N_3878);
and U4006 (N_4006,N_3847,N_3971);
xor U4007 (N_4007,N_3921,N_3881);
nand U4008 (N_4008,N_3858,N_3888);
xnor U4009 (N_4009,N_3901,N_3899);
and U4010 (N_4010,N_3845,N_3889);
nand U4011 (N_4011,N_3998,N_3907);
xnor U4012 (N_4012,N_3838,N_3989);
and U4013 (N_4013,N_3916,N_3859);
or U4014 (N_4014,N_3976,N_3846);
nand U4015 (N_4015,N_3884,N_3984);
and U4016 (N_4016,N_3886,N_3947);
nor U4017 (N_4017,N_3874,N_3939);
or U4018 (N_4018,N_3908,N_3816);
xor U4019 (N_4019,N_3988,N_3904);
xor U4020 (N_4020,N_3802,N_3946);
nand U4021 (N_4021,N_3920,N_3880);
and U4022 (N_4022,N_3887,N_3915);
xor U4023 (N_4023,N_3806,N_3829);
or U4024 (N_4024,N_3814,N_3955);
nand U4025 (N_4025,N_3926,N_3934);
or U4026 (N_4026,N_3841,N_3807);
and U4027 (N_4027,N_3892,N_3876);
nor U4028 (N_4028,N_3909,N_3905);
and U4029 (N_4029,N_3821,N_3959);
nor U4030 (N_4030,N_3834,N_3922);
and U4031 (N_4031,N_3914,N_3817);
nand U4032 (N_4032,N_3995,N_3818);
and U4033 (N_4033,N_3969,N_3891);
nor U4034 (N_4034,N_3911,N_3831);
nor U4035 (N_4035,N_3918,N_3912);
xor U4036 (N_4036,N_3862,N_3820);
nor U4037 (N_4037,N_3986,N_3835);
nand U4038 (N_4038,N_3963,N_3966);
xor U4039 (N_4039,N_3864,N_3804);
and U4040 (N_4040,N_3942,N_3941);
xor U4041 (N_4041,N_3879,N_3932);
and U4042 (N_4042,N_3953,N_3945);
nor U4043 (N_4043,N_3882,N_3935);
nand U4044 (N_4044,N_3848,N_3877);
nor U4045 (N_4045,N_3993,N_3973);
xor U4046 (N_4046,N_3872,N_3923);
and U4047 (N_4047,N_3819,N_3885);
or U4048 (N_4048,N_3960,N_3965);
nor U4049 (N_4049,N_3990,N_3843);
xor U4050 (N_4050,N_3893,N_3956);
or U4051 (N_4051,N_3983,N_3928);
nand U4052 (N_4052,N_3933,N_3854);
or U4053 (N_4053,N_3937,N_3803);
nor U4054 (N_4054,N_3824,N_3873);
or U4055 (N_4055,N_3936,N_3894);
nand U4056 (N_4056,N_3844,N_3865);
or U4057 (N_4057,N_3897,N_3801);
xnor U4058 (N_4058,N_3883,N_3855);
or U4059 (N_4059,N_3943,N_3991);
nor U4060 (N_4060,N_3827,N_3842);
and U4061 (N_4061,N_3868,N_3805);
xor U4062 (N_4062,N_3967,N_3851);
nor U4063 (N_4063,N_3852,N_3875);
and U4064 (N_4064,N_3828,N_3861);
nand U4065 (N_4065,N_3974,N_3800);
xor U4066 (N_4066,N_3930,N_3968);
and U4067 (N_4067,N_3867,N_3826);
or U4068 (N_4068,N_3811,N_3825);
nor U4069 (N_4069,N_3977,N_3954);
nand U4070 (N_4070,N_3871,N_3863);
nand U4071 (N_4071,N_3961,N_3840);
and U4072 (N_4072,N_3813,N_3987);
xnor U4073 (N_4073,N_3931,N_3964);
xor U4074 (N_4074,N_3980,N_3938);
nand U4075 (N_4075,N_3815,N_3962);
or U4076 (N_4076,N_3906,N_3924);
nand U4077 (N_4077,N_3996,N_3978);
nand U4078 (N_4078,N_3890,N_3832);
nand U4079 (N_4079,N_3927,N_3910);
nand U4080 (N_4080,N_3940,N_3870);
xor U4081 (N_4081,N_3975,N_3902);
nand U4082 (N_4082,N_3837,N_3982);
and U4083 (N_4083,N_3985,N_3857);
xnor U4084 (N_4084,N_3992,N_3979);
nand U4085 (N_4085,N_3866,N_3836);
nand U4086 (N_4086,N_3917,N_3948);
and U4087 (N_4087,N_3895,N_3853);
nor U4088 (N_4088,N_3822,N_3849);
and U4089 (N_4089,N_3981,N_3809);
nand U4090 (N_4090,N_3957,N_3839);
xor U4091 (N_4091,N_3950,N_3944);
nand U4092 (N_4092,N_3823,N_3808);
nand U4093 (N_4093,N_3994,N_3999);
nor U4094 (N_4094,N_3952,N_3850);
nand U4095 (N_4095,N_3913,N_3900);
nor U4096 (N_4096,N_3951,N_3997);
xor U4097 (N_4097,N_3812,N_3925);
or U4098 (N_4098,N_3833,N_3929);
or U4099 (N_4099,N_3856,N_3949);
nand U4100 (N_4100,N_3927,N_3944);
xor U4101 (N_4101,N_3952,N_3953);
or U4102 (N_4102,N_3811,N_3971);
and U4103 (N_4103,N_3843,N_3816);
xor U4104 (N_4104,N_3858,N_3872);
nand U4105 (N_4105,N_3926,N_3907);
or U4106 (N_4106,N_3968,N_3898);
and U4107 (N_4107,N_3866,N_3804);
nor U4108 (N_4108,N_3888,N_3926);
xor U4109 (N_4109,N_3821,N_3892);
or U4110 (N_4110,N_3854,N_3814);
or U4111 (N_4111,N_3802,N_3971);
or U4112 (N_4112,N_3807,N_3858);
xnor U4113 (N_4113,N_3903,N_3931);
or U4114 (N_4114,N_3882,N_3985);
and U4115 (N_4115,N_3911,N_3834);
xor U4116 (N_4116,N_3968,N_3965);
nand U4117 (N_4117,N_3948,N_3816);
and U4118 (N_4118,N_3834,N_3912);
xnor U4119 (N_4119,N_3803,N_3981);
or U4120 (N_4120,N_3998,N_3848);
nand U4121 (N_4121,N_3811,N_3932);
nand U4122 (N_4122,N_3857,N_3992);
or U4123 (N_4123,N_3889,N_3868);
nand U4124 (N_4124,N_3815,N_3981);
xor U4125 (N_4125,N_3850,N_3803);
nand U4126 (N_4126,N_3875,N_3905);
nand U4127 (N_4127,N_3908,N_3988);
xor U4128 (N_4128,N_3943,N_3931);
or U4129 (N_4129,N_3846,N_3934);
or U4130 (N_4130,N_3923,N_3985);
nor U4131 (N_4131,N_3867,N_3860);
and U4132 (N_4132,N_3810,N_3875);
xnor U4133 (N_4133,N_3982,N_3973);
or U4134 (N_4134,N_3941,N_3962);
or U4135 (N_4135,N_3969,N_3911);
xor U4136 (N_4136,N_3802,N_3949);
nor U4137 (N_4137,N_3991,N_3952);
nor U4138 (N_4138,N_3945,N_3943);
or U4139 (N_4139,N_3830,N_3934);
xor U4140 (N_4140,N_3824,N_3860);
xor U4141 (N_4141,N_3859,N_3802);
nand U4142 (N_4142,N_3855,N_3874);
xnor U4143 (N_4143,N_3819,N_3841);
xor U4144 (N_4144,N_3977,N_3811);
and U4145 (N_4145,N_3807,N_3853);
xor U4146 (N_4146,N_3966,N_3930);
nand U4147 (N_4147,N_3881,N_3847);
nor U4148 (N_4148,N_3921,N_3889);
xor U4149 (N_4149,N_3875,N_3944);
and U4150 (N_4150,N_3953,N_3933);
or U4151 (N_4151,N_3898,N_3870);
nor U4152 (N_4152,N_3972,N_3869);
and U4153 (N_4153,N_3871,N_3977);
or U4154 (N_4154,N_3976,N_3963);
nor U4155 (N_4155,N_3957,N_3996);
and U4156 (N_4156,N_3911,N_3891);
and U4157 (N_4157,N_3965,N_3910);
and U4158 (N_4158,N_3826,N_3835);
xnor U4159 (N_4159,N_3991,N_3850);
or U4160 (N_4160,N_3992,N_3835);
and U4161 (N_4161,N_3966,N_3955);
nand U4162 (N_4162,N_3881,N_3863);
or U4163 (N_4163,N_3939,N_3958);
xnor U4164 (N_4164,N_3805,N_3856);
or U4165 (N_4165,N_3922,N_3944);
nor U4166 (N_4166,N_3922,N_3845);
nor U4167 (N_4167,N_3860,N_3978);
nor U4168 (N_4168,N_3804,N_3913);
and U4169 (N_4169,N_3806,N_3938);
nor U4170 (N_4170,N_3912,N_3813);
and U4171 (N_4171,N_3867,N_3897);
nand U4172 (N_4172,N_3835,N_3972);
or U4173 (N_4173,N_3917,N_3811);
or U4174 (N_4174,N_3958,N_3825);
or U4175 (N_4175,N_3993,N_3958);
and U4176 (N_4176,N_3935,N_3809);
nor U4177 (N_4177,N_3946,N_3853);
nand U4178 (N_4178,N_3838,N_3867);
or U4179 (N_4179,N_3822,N_3960);
and U4180 (N_4180,N_3914,N_3972);
and U4181 (N_4181,N_3974,N_3946);
or U4182 (N_4182,N_3919,N_3925);
or U4183 (N_4183,N_3904,N_3870);
and U4184 (N_4184,N_3938,N_3935);
and U4185 (N_4185,N_3975,N_3925);
or U4186 (N_4186,N_3956,N_3826);
xnor U4187 (N_4187,N_3952,N_3941);
nor U4188 (N_4188,N_3813,N_3935);
or U4189 (N_4189,N_3891,N_3920);
and U4190 (N_4190,N_3836,N_3832);
or U4191 (N_4191,N_3819,N_3941);
xor U4192 (N_4192,N_3876,N_3882);
or U4193 (N_4193,N_3903,N_3904);
xnor U4194 (N_4194,N_3904,N_3898);
nand U4195 (N_4195,N_3959,N_3808);
and U4196 (N_4196,N_3873,N_3864);
nand U4197 (N_4197,N_3918,N_3844);
nor U4198 (N_4198,N_3947,N_3938);
and U4199 (N_4199,N_3998,N_3915);
nor U4200 (N_4200,N_4075,N_4191);
nand U4201 (N_4201,N_4161,N_4083);
nor U4202 (N_4202,N_4045,N_4085);
and U4203 (N_4203,N_4029,N_4046);
nand U4204 (N_4204,N_4089,N_4016);
or U4205 (N_4205,N_4010,N_4130);
nor U4206 (N_4206,N_4023,N_4117);
and U4207 (N_4207,N_4095,N_4040);
and U4208 (N_4208,N_4155,N_4019);
or U4209 (N_4209,N_4113,N_4140);
nand U4210 (N_4210,N_4074,N_4011);
or U4211 (N_4211,N_4056,N_4096);
nand U4212 (N_4212,N_4171,N_4157);
xor U4213 (N_4213,N_4104,N_4060);
nand U4214 (N_4214,N_4091,N_4017);
nand U4215 (N_4215,N_4057,N_4195);
nor U4216 (N_4216,N_4153,N_4000);
or U4217 (N_4217,N_4167,N_4077);
nand U4218 (N_4218,N_4124,N_4193);
xor U4219 (N_4219,N_4135,N_4047);
or U4220 (N_4220,N_4072,N_4165);
nor U4221 (N_4221,N_4038,N_4169);
and U4222 (N_4222,N_4014,N_4173);
or U4223 (N_4223,N_4149,N_4110);
or U4224 (N_4224,N_4128,N_4189);
xor U4225 (N_4225,N_4184,N_4129);
nor U4226 (N_4226,N_4094,N_4177);
or U4227 (N_4227,N_4101,N_4027);
or U4228 (N_4228,N_4194,N_4020);
and U4229 (N_4229,N_4133,N_4035);
xor U4230 (N_4230,N_4145,N_4059);
and U4231 (N_4231,N_4150,N_4061);
xor U4232 (N_4232,N_4190,N_4136);
or U4233 (N_4233,N_4030,N_4097);
or U4234 (N_4234,N_4007,N_4141);
or U4235 (N_4235,N_4116,N_4158);
nor U4236 (N_4236,N_4071,N_4179);
and U4237 (N_4237,N_4032,N_4028);
nor U4238 (N_4238,N_4044,N_4144);
or U4239 (N_4239,N_4152,N_4002);
or U4240 (N_4240,N_4178,N_4005);
or U4241 (N_4241,N_4049,N_4121);
nand U4242 (N_4242,N_4070,N_4119);
nor U4243 (N_4243,N_4086,N_4185);
xnor U4244 (N_4244,N_4127,N_4118);
or U4245 (N_4245,N_4122,N_4031);
and U4246 (N_4246,N_4092,N_4143);
nor U4247 (N_4247,N_4142,N_4114);
xor U4248 (N_4248,N_4034,N_4079);
or U4249 (N_4249,N_4001,N_4013);
nor U4250 (N_4250,N_4058,N_4131);
or U4251 (N_4251,N_4112,N_4053);
or U4252 (N_4252,N_4054,N_4088);
nand U4253 (N_4253,N_4115,N_4093);
xor U4254 (N_4254,N_4036,N_4164);
or U4255 (N_4255,N_4111,N_4103);
xnor U4256 (N_4256,N_4139,N_4174);
or U4257 (N_4257,N_4162,N_4106);
nor U4258 (N_4258,N_4098,N_4182);
nand U4259 (N_4259,N_4062,N_4105);
or U4260 (N_4260,N_4187,N_4125);
nor U4261 (N_4261,N_4082,N_4163);
and U4262 (N_4262,N_4022,N_4196);
nor U4263 (N_4263,N_4154,N_4048);
nor U4264 (N_4264,N_4024,N_4069);
and U4265 (N_4265,N_4175,N_4134);
nor U4266 (N_4266,N_4197,N_4004);
xor U4267 (N_4267,N_4084,N_4108);
and U4268 (N_4268,N_4050,N_4076);
and U4269 (N_4269,N_4160,N_4021);
and U4270 (N_4270,N_4102,N_4041);
nand U4271 (N_4271,N_4052,N_4015);
or U4272 (N_4272,N_4073,N_4166);
xor U4273 (N_4273,N_4026,N_4176);
xnor U4274 (N_4274,N_4078,N_4064);
xor U4275 (N_4275,N_4018,N_4065);
xnor U4276 (N_4276,N_4181,N_4199);
xor U4277 (N_4277,N_4159,N_4067);
or U4278 (N_4278,N_4037,N_4090);
or U4279 (N_4279,N_4051,N_4039);
and U4280 (N_4280,N_4066,N_4151);
nand U4281 (N_4281,N_4192,N_4180);
nand U4282 (N_4282,N_4081,N_4033);
and U4283 (N_4283,N_4168,N_4188);
or U4284 (N_4284,N_4126,N_4012);
and U4285 (N_4285,N_4009,N_4107);
nand U4286 (N_4286,N_4042,N_4080);
xor U4287 (N_4287,N_4138,N_4146);
nor U4288 (N_4288,N_4170,N_4043);
or U4289 (N_4289,N_4068,N_4123);
nand U4290 (N_4290,N_4198,N_4055);
or U4291 (N_4291,N_4148,N_4147);
nand U4292 (N_4292,N_4132,N_4006);
nor U4293 (N_4293,N_4087,N_4003);
xor U4294 (N_4294,N_4137,N_4109);
and U4295 (N_4295,N_4183,N_4156);
and U4296 (N_4296,N_4100,N_4120);
nor U4297 (N_4297,N_4008,N_4025);
nand U4298 (N_4298,N_4099,N_4172);
and U4299 (N_4299,N_4186,N_4063);
and U4300 (N_4300,N_4171,N_4044);
and U4301 (N_4301,N_4198,N_4037);
nor U4302 (N_4302,N_4182,N_4188);
nand U4303 (N_4303,N_4096,N_4193);
nor U4304 (N_4304,N_4047,N_4041);
and U4305 (N_4305,N_4028,N_4187);
nand U4306 (N_4306,N_4171,N_4194);
xor U4307 (N_4307,N_4068,N_4146);
nor U4308 (N_4308,N_4197,N_4181);
or U4309 (N_4309,N_4039,N_4048);
or U4310 (N_4310,N_4096,N_4184);
or U4311 (N_4311,N_4092,N_4075);
or U4312 (N_4312,N_4111,N_4104);
or U4313 (N_4313,N_4109,N_4096);
nand U4314 (N_4314,N_4065,N_4137);
xor U4315 (N_4315,N_4044,N_4147);
nand U4316 (N_4316,N_4124,N_4076);
and U4317 (N_4317,N_4100,N_4045);
nor U4318 (N_4318,N_4186,N_4149);
and U4319 (N_4319,N_4172,N_4010);
xor U4320 (N_4320,N_4159,N_4011);
nand U4321 (N_4321,N_4109,N_4157);
xnor U4322 (N_4322,N_4042,N_4191);
xnor U4323 (N_4323,N_4019,N_4114);
or U4324 (N_4324,N_4061,N_4102);
xor U4325 (N_4325,N_4069,N_4017);
nand U4326 (N_4326,N_4061,N_4153);
xnor U4327 (N_4327,N_4096,N_4016);
xnor U4328 (N_4328,N_4174,N_4010);
or U4329 (N_4329,N_4039,N_4005);
nand U4330 (N_4330,N_4000,N_4019);
or U4331 (N_4331,N_4090,N_4035);
xnor U4332 (N_4332,N_4039,N_4118);
xnor U4333 (N_4333,N_4199,N_4098);
and U4334 (N_4334,N_4063,N_4174);
and U4335 (N_4335,N_4131,N_4144);
and U4336 (N_4336,N_4075,N_4028);
and U4337 (N_4337,N_4019,N_4065);
or U4338 (N_4338,N_4041,N_4150);
or U4339 (N_4339,N_4165,N_4142);
and U4340 (N_4340,N_4085,N_4096);
and U4341 (N_4341,N_4164,N_4021);
xor U4342 (N_4342,N_4014,N_4036);
and U4343 (N_4343,N_4128,N_4065);
xnor U4344 (N_4344,N_4107,N_4178);
and U4345 (N_4345,N_4193,N_4083);
and U4346 (N_4346,N_4084,N_4082);
xor U4347 (N_4347,N_4063,N_4151);
and U4348 (N_4348,N_4112,N_4100);
or U4349 (N_4349,N_4198,N_4144);
nor U4350 (N_4350,N_4166,N_4149);
xor U4351 (N_4351,N_4159,N_4059);
nor U4352 (N_4352,N_4142,N_4107);
nand U4353 (N_4353,N_4179,N_4009);
and U4354 (N_4354,N_4102,N_4111);
xor U4355 (N_4355,N_4115,N_4036);
nand U4356 (N_4356,N_4124,N_4117);
nor U4357 (N_4357,N_4129,N_4163);
nor U4358 (N_4358,N_4003,N_4016);
and U4359 (N_4359,N_4151,N_4174);
or U4360 (N_4360,N_4050,N_4162);
or U4361 (N_4361,N_4193,N_4163);
nand U4362 (N_4362,N_4147,N_4038);
xor U4363 (N_4363,N_4169,N_4074);
nor U4364 (N_4364,N_4019,N_4035);
xnor U4365 (N_4365,N_4195,N_4017);
nor U4366 (N_4366,N_4060,N_4134);
or U4367 (N_4367,N_4127,N_4062);
nand U4368 (N_4368,N_4125,N_4150);
or U4369 (N_4369,N_4095,N_4029);
and U4370 (N_4370,N_4123,N_4156);
or U4371 (N_4371,N_4158,N_4110);
nand U4372 (N_4372,N_4027,N_4114);
nor U4373 (N_4373,N_4078,N_4074);
or U4374 (N_4374,N_4195,N_4000);
xnor U4375 (N_4375,N_4012,N_4113);
nand U4376 (N_4376,N_4024,N_4092);
and U4377 (N_4377,N_4023,N_4018);
xnor U4378 (N_4378,N_4018,N_4055);
and U4379 (N_4379,N_4121,N_4037);
xor U4380 (N_4380,N_4024,N_4107);
or U4381 (N_4381,N_4101,N_4123);
or U4382 (N_4382,N_4169,N_4016);
or U4383 (N_4383,N_4057,N_4186);
nand U4384 (N_4384,N_4056,N_4060);
xnor U4385 (N_4385,N_4039,N_4104);
and U4386 (N_4386,N_4167,N_4013);
nor U4387 (N_4387,N_4132,N_4144);
or U4388 (N_4388,N_4021,N_4112);
and U4389 (N_4389,N_4098,N_4123);
nand U4390 (N_4390,N_4161,N_4120);
and U4391 (N_4391,N_4022,N_4127);
nand U4392 (N_4392,N_4121,N_4021);
nor U4393 (N_4393,N_4055,N_4095);
nand U4394 (N_4394,N_4065,N_4187);
and U4395 (N_4395,N_4045,N_4129);
nand U4396 (N_4396,N_4071,N_4003);
nand U4397 (N_4397,N_4033,N_4167);
nand U4398 (N_4398,N_4000,N_4016);
or U4399 (N_4399,N_4159,N_4070);
nand U4400 (N_4400,N_4362,N_4254);
xor U4401 (N_4401,N_4220,N_4335);
nor U4402 (N_4402,N_4355,N_4367);
xor U4403 (N_4403,N_4295,N_4292);
nand U4404 (N_4404,N_4307,N_4365);
or U4405 (N_4405,N_4380,N_4265);
nand U4406 (N_4406,N_4269,N_4356);
nand U4407 (N_4407,N_4350,N_4353);
nor U4408 (N_4408,N_4397,N_4309);
nor U4409 (N_4409,N_4261,N_4256);
nand U4410 (N_4410,N_4347,N_4332);
nand U4411 (N_4411,N_4334,N_4203);
nor U4412 (N_4412,N_4234,N_4391);
or U4413 (N_4413,N_4373,N_4349);
and U4414 (N_4414,N_4246,N_4341);
and U4415 (N_4415,N_4399,N_4238);
xor U4416 (N_4416,N_4210,N_4329);
and U4417 (N_4417,N_4308,N_4320);
nor U4418 (N_4418,N_4323,N_4363);
xnor U4419 (N_4419,N_4226,N_4326);
and U4420 (N_4420,N_4230,N_4227);
nor U4421 (N_4421,N_4303,N_4392);
and U4422 (N_4422,N_4384,N_4272);
xnor U4423 (N_4423,N_4263,N_4276);
xnor U4424 (N_4424,N_4270,N_4333);
and U4425 (N_4425,N_4288,N_4213);
or U4426 (N_4426,N_4337,N_4346);
or U4427 (N_4427,N_4340,N_4286);
and U4428 (N_4428,N_4374,N_4240);
or U4429 (N_4429,N_4376,N_4232);
and U4430 (N_4430,N_4275,N_4354);
nand U4431 (N_4431,N_4360,N_4242);
xor U4432 (N_4432,N_4321,N_4398);
or U4433 (N_4433,N_4236,N_4214);
and U4434 (N_4434,N_4388,N_4372);
and U4435 (N_4435,N_4218,N_4330);
and U4436 (N_4436,N_4248,N_4211);
or U4437 (N_4437,N_4268,N_4378);
nand U4438 (N_4438,N_4395,N_4369);
and U4439 (N_4439,N_4304,N_4207);
nor U4440 (N_4440,N_4316,N_4385);
nor U4441 (N_4441,N_4312,N_4260);
and U4442 (N_4442,N_4302,N_4318);
and U4443 (N_4443,N_4390,N_4361);
and U4444 (N_4444,N_4249,N_4208);
and U4445 (N_4445,N_4221,N_4215);
nor U4446 (N_4446,N_4257,N_4244);
or U4447 (N_4447,N_4206,N_4271);
xor U4448 (N_4448,N_4331,N_4239);
xor U4449 (N_4449,N_4294,N_4383);
and U4450 (N_4450,N_4216,N_4267);
nand U4451 (N_4451,N_4351,N_4322);
and U4452 (N_4452,N_4357,N_4262);
nand U4453 (N_4453,N_4219,N_4342);
nand U4454 (N_4454,N_4313,N_4223);
nand U4455 (N_4455,N_4387,N_4358);
xnor U4456 (N_4456,N_4379,N_4299);
nor U4457 (N_4457,N_4317,N_4325);
or U4458 (N_4458,N_4310,N_4297);
xor U4459 (N_4459,N_4389,N_4235);
nor U4460 (N_4460,N_4266,N_4345);
xnor U4461 (N_4461,N_4306,N_4328);
and U4462 (N_4462,N_4375,N_4370);
or U4463 (N_4463,N_4247,N_4282);
nand U4464 (N_4464,N_4280,N_4339);
nor U4465 (N_4465,N_4301,N_4291);
or U4466 (N_4466,N_4289,N_4277);
xor U4467 (N_4467,N_4336,N_4396);
or U4468 (N_4468,N_4348,N_4217);
nor U4469 (N_4469,N_4382,N_4287);
nand U4470 (N_4470,N_4264,N_4212);
nand U4471 (N_4471,N_4352,N_4381);
or U4472 (N_4472,N_4255,N_4314);
nand U4473 (N_4473,N_4241,N_4386);
nor U4474 (N_4474,N_4201,N_4368);
or U4475 (N_4475,N_4237,N_4202);
xnor U4476 (N_4476,N_4224,N_4359);
nand U4477 (N_4477,N_4258,N_4366);
and U4478 (N_4478,N_4298,N_4205);
xnor U4479 (N_4479,N_4296,N_4259);
xnor U4480 (N_4480,N_4377,N_4209);
and U4481 (N_4481,N_4343,N_4300);
nand U4482 (N_4482,N_4245,N_4293);
nor U4483 (N_4483,N_4393,N_4284);
nor U4484 (N_4484,N_4233,N_4281);
and U4485 (N_4485,N_4290,N_4229);
xnor U4486 (N_4486,N_4252,N_4319);
nor U4487 (N_4487,N_4222,N_4285);
nand U4488 (N_4488,N_4228,N_4204);
and U4489 (N_4489,N_4251,N_4305);
nand U4490 (N_4490,N_4283,N_4243);
or U4491 (N_4491,N_4279,N_4274);
nand U4492 (N_4492,N_4344,N_4324);
xor U4493 (N_4493,N_4394,N_4364);
or U4494 (N_4494,N_4315,N_4225);
xnor U4495 (N_4495,N_4371,N_4327);
or U4496 (N_4496,N_4200,N_4273);
nand U4497 (N_4497,N_4231,N_4278);
nand U4498 (N_4498,N_4311,N_4253);
nor U4499 (N_4499,N_4250,N_4338);
xnor U4500 (N_4500,N_4221,N_4366);
or U4501 (N_4501,N_4373,N_4201);
or U4502 (N_4502,N_4365,N_4385);
or U4503 (N_4503,N_4360,N_4251);
or U4504 (N_4504,N_4328,N_4302);
and U4505 (N_4505,N_4216,N_4311);
xor U4506 (N_4506,N_4219,N_4256);
or U4507 (N_4507,N_4336,N_4288);
nand U4508 (N_4508,N_4373,N_4392);
nand U4509 (N_4509,N_4394,N_4333);
or U4510 (N_4510,N_4244,N_4378);
nor U4511 (N_4511,N_4332,N_4317);
and U4512 (N_4512,N_4224,N_4201);
nor U4513 (N_4513,N_4258,N_4353);
or U4514 (N_4514,N_4306,N_4395);
xnor U4515 (N_4515,N_4310,N_4293);
xor U4516 (N_4516,N_4321,N_4243);
nand U4517 (N_4517,N_4202,N_4206);
and U4518 (N_4518,N_4328,N_4279);
nor U4519 (N_4519,N_4300,N_4264);
and U4520 (N_4520,N_4203,N_4290);
nor U4521 (N_4521,N_4263,N_4380);
xnor U4522 (N_4522,N_4268,N_4247);
or U4523 (N_4523,N_4397,N_4373);
nor U4524 (N_4524,N_4357,N_4286);
or U4525 (N_4525,N_4214,N_4395);
and U4526 (N_4526,N_4232,N_4216);
nand U4527 (N_4527,N_4358,N_4359);
xor U4528 (N_4528,N_4253,N_4329);
and U4529 (N_4529,N_4319,N_4363);
and U4530 (N_4530,N_4288,N_4399);
nor U4531 (N_4531,N_4202,N_4269);
nand U4532 (N_4532,N_4326,N_4348);
and U4533 (N_4533,N_4332,N_4253);
or U4534 (N_4534,N_4386,N_4278);
and U4535 (N_4535,N_4207,N_4294);
or U4536 (N_4536,N_4284,N_4365);
nand U4537 (N_4537,N_4248,N_4297);
nand U4538 (N_4538,N_4254,N_4305);
nor U4539 (N_4539,N_4363,N_4303);
nand U4540 (N_4540,N_4351,N_4245);
nand U4541 (N_4541,N_4346,N_4246);
nor U4542 (N_4542,N_4283,N_4342);
and U4543 (N_4543,N_4232,N_4369);
nor U4544 (N_4544,N_4278,N_4319);
nor U4545 (N_4545,N_4244,N_4282);
and U4546 (N_4546,N_4386,N_4200);
or U4547 (N_4547,N_4387,N_4392);
and U4548 (N_4548,N_4331,N_4254);
nand U4549 (N_4549,N_4226,N_4358);
or U4550 (N_4550,N_4340,N_4347);
or U4551 (N_4551,N_4319,N_4253);
and U4552 (N_4552,N_4260,N_4396);
nand U4553 (N_4553,N_4243,N_4302);
or U4554 (N_4554,N_4301,N_4223);
xor U4555 (N_4555,N_4377,N_4228);
nand U4556 (N_4556,N_4326,N_4363);
nor U4557 (N_4557,N_4320,N_4302);
or U4558 (N_4558,N_4378,N_4232);
nor U4559 (N_4559,N_4321,N_4327);
nor U4560 (N_4560,N_4213,N_4307);
nand U4561 (N_4561,N_4372,N_4225);
nand U4562 (N_4562,N_4328,N_4240);
nand U4563 (N_4563,N_4201,N_4209);
nand U4564 (N_4564,N_4320,N_4337);
and U4565 (N_4565,N_4325,N_4352);
xnor U4566 (N_4566,N_4308,N_4228);
nand U4567 (N_4567,N_4384,N_4341);
and U4568 (N_4568,N_4242,N_4397);
or U4569 (N_4569,N_4321,N_4288);
and U4570 (N_4570,N_4312,N_4293);
or U4571 (N_4571,N_4296,N_4323);
nand U4572 (N_4572,N_4380,N_4239);
or U4573 (N_4573,N_4318,N_4226);
and U4574 (N_4574,N_4281,N_4333);
nand U4575 (N_4575,N_4200,N_4360);
and U4576 (N_4576,N_4272,N_4300);
nand U4577 (N_4577,N_4350,N_4392);
and U4578 (N_4578,N_4232,N_4390);
nand U4579 (N_4579,N_4236,N_4362);
nand U4580 (N_4580,N_4331,N_4325);
nor U4581 (N_4581,N_4314,N_4239);
xnor U4582 (N_4582,N_4320,N_4381);
and U4583 (N_4583,N_4335,N_4367);
and U4584 (N_4584,N_4288,N_4218);
or U4585 (N_4585,N_4219,N_4236);
xor U4586 (N_4586,N_4319,N_4360);
and U4587 (N_4587,N_4224,N_4367);
and U4588 (N_4588,N_4280,N_4205);
xor U4589 (N_4589,N_4279,N_4224);
and U4590 (N_4590,N_4385,N_4248);
nand U4591 (N_4591,N_4236,N_4340);
or U4592 (N_4592,N_4350,N_4236);
nor U4593 (N_4593,N_4243,N_4260);
xor U4594 (N_4594,N_4283,N_4382);
or U4595 (N_4595,N_4344,N_4228);
nor U4596 (N_4596,N_4290,N_4333);
and U4597 (N_4597,N_4256,N_4353);
nor U4598 (N_4598,N_4280,N_4200);
and U4599 (N_4599,N_4243,N_4245);
nand U4600 (N_4600,N_4555,N_4570);
xor U4601 (N_4601,N_4411,N_4418);
nand U4602 (N_4602,N_4547,N_4559);
and U4603 (N_4603,N_4569,N_4489);
nor U4604 (N_4604,N_4575,N_4542);
nor U4605 (N_4605,N_4476,N_4430);
nand U4606 (N_4606,N_4456,N_4447);
and U4607 (N_4607,N_4409,N_4593);
and U4608 (N_4608,N_4518,N_4498);
xnor U4609 (N_4609,N_4434,N_4545);
nor U4610 (N_4610,N_4460,N_4455);
nor U4611 (N_4611,N_4468,N_4532);
nand U4612 (N_4612,N_4412,N_4470);
nor U4613 (N_4613,N_4452,N_4515);
xnor U4614 (N_4614,N_4502,N_4562);
nand U4615 (N_4615,N_4513,N_4438);
nand U4616 (N_4616,N_4481,N_4501);
xor U4617 (N_4617,N_4487,N_4488);
nand U4618 (N_4618,N_4568,N_4520);
or U4619 (N_4619,N_4473,N_4403);
or U4620 (N_4620,N_4554,N_4478);
or U4621 (N_4621,N_4553,N_4537);
nor U4622 (N_4622,N_4509,N_4529);
and U4623 (N_4623,N_4400,N_4408);
xnor U4624 (N_4624,N_4424,N_4457);
nor U4625 (N_4625,N_4578,N_4466);
nor U4626 (N_4626,N_4469,N_4508);
and U4627 (N_4627,N_4480,N_4504);
nand U4628 (N_4628,N_4591,N_4528);
xor U4629 (N_4629,N_4448,N_4477);
nor U4630 (N_4630,N_4556,N_4436);
nand U4631 (N_4631,N_4486,N_4552);
nand U4632 (N_4632,N_4546,N_4527);
nand U4633 (N_4633,N_4482,N_4566);
nor U4634 (N_4634,N_4439,N_4597);
and U4635 (N_4635,N_4541,N_4573);
and U4636 (N_4636,N_4490,N_4450);
and U4637 (N_4637,N_4505,N_4415);
or U4638 (N_4638,N_4420,N_4596);
or U4639 (N_4639,N_4428,N_4453);
or U4640 (N_4640,N_4405,N_4407);
xor U4641 (N_4641,N_4565,N_4531);
nand U4642 (N_4642,N_4592,N_4497);
and U4643 (N_4643,N_4503,N_4581);
and U4644 (N_4644,N_4521,N_4494);
or U4645 (N_4645,N_4514,N_4406);
or U4646 (N_4646,N_4423,N_4574);
xnor U4647 (N_4647,N_4493,N_4516);
xnor U4648 (N_4648,N_4417,N_4451);
and U4649 (N_4649,N_4576,N_4454);
or U4650 (N_4650,N_4594,N_4491);
xnor U4651 (N_4651,N_4524,N_4425);
xor U4652 (N_4652,N_4538,N_4485);
nand U4653 (N_4653,N_4464,N_4401);
nor U4654 (N_4654,N_4551,N_4465);
nand U4655 (N_4655,N_4558,N_4462);
nor U4656 (N_4656,N_4442,N_4484);
nor U4657 (N_4657,N_4422,N_4441);
nand U4658 (N_4658,N_4461,N_4530);
nor U4659 (N_4659,N_4584,N_4571);
nor U4660 (N_4660,N_4586,N_4599);
and U4661 (N_4661,N_4517,N_4421);
or U4662 (N_4662,N_4427,N_4572);
nor U4663 (N_4663,N_4522,N_4444);
nand U4664 (N_4664,N_4431,N_4540);
nand U4665 (N_4665,N_4402,N_4589);
or U4666 (N_4666,N_4496,N_4507);
nand U4667 (N_4667,N_4419,N_4426);
xnor U4668 (N_4668,N_4588,N_4413);
nand U4669 (N_4669,N_4432,N_4445);
nor U4670 (N_4670,N_4583,N_4533);
or U4671 (N_4671,N_4467,N_4410);
xor U4672 (N_4672,N_4510,N_4544);
or U4673 (N_4673,N_4526,N_4506);
nand U4674 (N_4674,N_4564,N_4474);
and U4675 (N_4675,N_4577,N_4475);
xor U4676 (N_4676,N_4483,N_4525);
nor U4677 (N_4677,N_4440,N_4560);
or U4678 (N_4678,N_4443,N_4561);
nand U4679 (N_4679,N_4587,N_4512);
or U4680 (N_4680,N_4459,N_4416);
nor U4681 (N_4681,N_4500,N_4414);
or U4682 (N_4682,N_4523,N_4472);
or U4683 (N_4683,N_4548,N_4535);
or U4684 (N_4684,N_4437,N_4471);
nand U4685 (N_4685,N_4433,N_4429);
or U4686 (N_4686,N_4519,N_4404);
or U4687 (N_4687,N_4595,N_4579);
and U4688 (N_4688,N_4492,N_4567);
xnor U4689 (N_4689,N_4499,N_4543);
nor U4690 (N_4690,N_4557,N_4479);
and U4691 (N_4691,N_4536,N_4463);
xnor U4692 (N_4692,N_4495,N_4582);
xnor U4693 (N_4693,N_4539,N_4549);
or U4694 (N_4694,N_4580,N_4458);
nor U4695 (N_4695,N_4511,N_4435);
and U4696 (N_4696,N_4590,N_4534);
nor U4697 (N_4697,N_4550,N_4585);
nand U4698 (N_4698,N_4446,N_4598);
or U4699 (N_4699,N_4449,N_4563);
or U4700 (N_4700,N_4473,N_4431);
xor U4701 (N_4701,N_4585,N_4503);
nand U4702 (N_4702,N_4474,N_4467);
and U4703 (N_4703,N_4527,N_4573);
or U4704 (N_4704,N_4591,N_4406);
or U4705 (N_4705,N_4507,N_4467);
and U4706 (N_4706,N_4503,N_4497);
or U4707 (N_4707,N_4511,N_4493);
xnor U4708 (N_4708,N_4591,N_4451);
xor U4709 (N_4709,N_4465,N_4540);
or U4710 (N_4710,N_4461,N_4465);
nor U4711 (N_4711,N_4586,N_4447);
nand U4712 (N_4712,N_4411,N_4431);
nand U4713 (N_4713,N_4444,N_4495);
nand U4714 (N_4714,N_4455,N_4508);
nand U4715 (N_4715,N_4455,N_4501);
nand U4716 (N_4716,N_4427,N_4504);
nand U4717 (N_4717,N_4472,N_4506);
or U4718 (N_4718,N_4586,N_4427);
nor U4719 (N_4719,N_4594,N_4443);
nand U4720 (N_4720,N_4413,N_4469);
xor U4721 (N_4721,N_4436,N_4492);
nor U4722 (N_4722,N_4482,N_4569);
nor U4723 (N_4723,N_4587,N_4545);
xor U4724 (N_4724,N_4416,N_4400);
xnor U4725 (N_4725,N_4539,N_4435);
xnor U4726 (N_4726,N_4500,N_4549);
and U4727 (N_4727,N_4410,N_4521);
or U4728 (N_4728,N_4478,N_4493);
xnor U4729 (N_4729,N_4561,N_4450);
nand U4730 (N_4730,N_4443,N_4598);
nand U4731 (N_4731,N_4588,N_4576);
nor U4732 (N_4732,N_4404,N_4597);
or U4733 (N_4733,N_4454,N_4422);
and U4734 (N_4734,N_4590,N_4440);
nand U4735 (N_4735,N_4431,N_4429);
xnor U4736 (N_4736,N_4450,N_4554);
and U4737 (N_4737,N_4528,N_4576);
xnor U4738 (N_4738,N_4400,N_4424);
nand U4739 (N_4739,N_4586,N_4433);
nor U4740 (N_4740,N_4581,N_4415);
nand U4741 (N_4741,N_4559,N_4437);
nand U4742 (N_4742,N_4458,N_4474);
xnor U4743 (N_4743,N_4444,N_4466);
nand U4744 (N_4744,N_4430,N_4576);
nor U4745 (N_4745,N_4491,N_4417);
xor U4746 (N_4746,N_4562,N_4509);
or U4747 (N_4747,N_4403,N_4544);
xnor U4748 (N_4748,N_4455,N_4548);
nand U4749 (N_4749,N_4562,N_4539);
nor U4750 (N_4750,N_4444,N_4416);
or U4751 (N_4751,N_4589,N_4586);
nand U4752 (N_4752,N_4503,N_4578);
xor U4753 (N_4753,N_4401,N_4565);
nand U4754 (N_4754,N_4539,N_4401);
nand U4755 (N_4755,N_4436,N_4477);
xor U4756 (N_4756,N_4448,N_4536);
nand U4757 (N_4757,N_4440,N_4485);
xnor U4758 (N_4758,N_4503,N_4548);
and U4759 (N_4759,N_4474,N_4413);
nor U4760 (N_4760,N_4532,N_4471);
and U4761 (N_4761,N_4453,N_4536);
nand U4762 (N_4762,N_4589,N_4597);
xnor U4763 (N_4763,N_4599,N_4570);
or U4764 (N_4764,N_4517,N_4481);
nand U4765 (N_4765,N_4417,N_4517);
nor U4766 (N_4766,N_4549,N_4568);
or U4767 (N_4767,N_4509,N_4416);
and U4768 (N_4768,N_4599,N_4412);
or U4769 (N_4769,N_4504,N_4576);
and U4770 (N_4770,N_4554,N_4485);
or U4771 (N_4771,N_4444,N_4419);
xnor U4772 (N_4772,N_4457,N_4569);
and U4773 (N_4773,N_4509,N_4485);
or U4774 (N_4774,N_4465,N_4470);
nor U4775 (N_4775,N_4590,N_4587);
nor U4776 (N_4776,N_4416,N_4479);
xnor U4777 (N_4777,N_4579,N_4428);
nor U4778 (N_4778,N_4523,N_4411);
nor U4779 (N_4779,N_4523,N_4574);
nor U4780 (N_4780,N_4452,N_4532);
and U4781 (N_4781,N_4493,N_4577);
xnor U4782 (N_4782,N_4553,N_4437);
nor U4783 (N_4783,N_4436,N_4592);
and U4784 (N_4784,N_4511,N_4486);
or U4785 (N_4785,N_4451,N_4526);
nand U4786 (N_4786,N_4597,N_4533);
nor U4787 (N_4787,N_4525,N_4418);
nor U4788 (N_4788,N_4418,N_4465);
nor U4789 (N_4789,N_4539,N_4565);
nand U4790 (N_4790,N_4536,N_4430);
xnor U4791 (N_4791,N_4590,N_4486);
and U4792 (N_4792,N_4430,N_4584);
and U4793 (N_4793,N_4581,N_4536);
or U4794 (N_4794,N_4408,N_4454);
or U4795 (N_4795,N_4580,N_4509);
xnor U4796 (N_4796,N_4497,N_4548);
nand U4797 (N_4797,N_4408,N_4517);
nor U4798 (N_4798,N_4463,N_4516);
or U4799 (N_4799,N_4552,N_4494);
or U4800 (N_4800,N_4746,N_4782);
nor U4801 (N_4801,N_4674,N_4623);
xor U4802 (N_4802,N_4644,N_4734);
and U4803 (N_4803,N_4751,N_4744);
and U4804 (N_4804,N_4667,N_4688);
nor U4805 (N_4805,N_4698,N_4686);
nor U4806 (N_4806,N_4666,N_4645);
and U4807 (N_4807,N_4671,N_4743);
nor U4808 (N_4808,N_4778,N_4723);
nor U4809 (N_4809,N_4607,N_4772);
nor U4810 (N_4810,N_4601,N_4610);
or U4811 (N_4811,N_4770,N_4745);
nand U4812 (N_4812,N_4689,N_4619);
nand U4813 (N_4813,N_4609,N_4614);
nor U4814 (N_4814,N_4629,N_4694);
and U4815 (N_4815,N_4718,N_4780);
or U4816 (N_4816,N_4732,N_4640);
and U4817 (N_4817,N_4706,N_4720);
nor U4818 (N_4818,N_4792,N_4652);
nand U4819 (N_4819,N_4765,N_4649);
and U4820 (N_4820,N_4626,N_4632);
nor U4821 (N_4821,N_4710,N_4736);
xnor U4822 (N_4822,N_4794,N_4657);
or U4823 (N_4823,N_4625,N_4722);
or U4824 (N_4824,N_4750,N_4799);
xor U4825 (N_4825,N_4662,N_4781);
nor U4826 (N_4826,N_4753,N_4687);
nor U4827 (N_4827,N_4615,N_4642);
and U4828 (N_4828,N_4774,N_4775);
nor U4829 (N_4829,N_4779,N_4622);
or U4830 (N_4830,N_4768,N_4664);
or U4831 (N_4831,N_4633,N_4691);
and U4832 (N_4832,N_4679,N_4740);
xor U4833 (N_4833,N_4643,N_4697);
nand U4834 (N_4834,N_4647,N_4630);
or U4835 (N_4835,N_4795,N_4798);
or U4836 (N_4836,N_4729,N_4635);
xnor U4837 (N_4837,N_4758,N_4637);
nand U4838 (N_4838,N_4721,N_4767);
or U4839 (N_4839,N_4608,N_4748);
xor U4840 (N_4840,N_4762,N_4787);
xor U4841 (N_4841,N_4764,N_4719);
nand U4842 (N_4842,N_4604,N_4788);
nor U4843 (N_4843,N_4757,N_4651);
and U4844 (N_4844,N_4755,N_4716);
and U4845 (N_4845,N_4760,N_4747);
nand U4846 (N_4846,N_4634,N_4702);
nor U4847 (N_4847,N_4650,N_4661);
nand U4848 (N_4848,N_4678,N_4638);
or U4849 (N_4849,N_4715,N_4646);
nor U4850 (N_4850,N_4703,N_4683);
or U4851 (N_4851,N_4654,N_4704);
nand U4852 (N_4852,N_4611,N_4725);
nor U4853 (N_4853,N_4738,N_4612);
and U4854 (N_4854,N_4685,N_4620);
or U4855 (N_4855,N_4696,N_4659);
or U4856 (N_4856,N_4766,N_4684);
nor U4857 (N_4857,N_4669,N_4700);
or U4858 (N_4858,N_4695,N_4724);
and U4859 (N_4859,N_4693,N_4737);
nand U4860 (N_4860,N_4648,N_4728);
and U4861 (N_4861,N_4769,N_4754);
xnor U4862 (N_4862,N_4699,N_4714);
nor U4863 (N_4863,N_4786,N_4790);
nand U4864 (N_4864,N_4656,N_4712);
nor U4865 (N_4865,N_4776,N_4713);
and U4866 (N_4866,N_4773,N_4761);
xor U4867 (N_4867,N_4791,N_4658);
xor U4868 (N_4868,N_4628,N_4600);
and U4869 (N_4869,N_4739,N_4705);
nand U4870 (N_4870,N_4735,N_4785);
nand U4871 (N_4871,N_4771,N_4639);
xor U4872 (N_4872,N_4707,N_4681);
nand U4873 (N_4873,N_4606,N_4665);
xor U4874 (N_4874,N_4730,N_4677);
nand U4875 (N_4875,N_4655,N_4676);
or U4876 (N_4876,N_4660,N_4627);
nor U4877 (N_4877,N_4613,N_4777);
nand U4878 (N_4878,N_4741,N_4617);
nor U4879 (N_4879,N_4701,N_4668);
or U4880 (N_4880,N_4663,N_4752);
nand U4881 (N_4881,N_4756,N_4759);
nor U4882 (N_4882,N_4784,N_4675);
nand U4883 (N_4883,N_4727,N_4682);
nor U4884 (N_4884,N_4670,N_4717);
xor U4885 (N_4885,N_4763,N_4796);
or U4886 (N_4886,N_4742,N_4631);
or U4887 (N_4887,N_4673,N_4641);
nor U4888 (N_4888,N_4733,N_4603);
or U4889 (N_4889,N_4783,N_4624);
and U4890 (N_4890,N_4797,N_4731);
xnor U4891 (N_4891,N_4692,N_4621);
and U4892 (N_4892,N_4726,N_4749);
nand U4893 (N_4893,N_4672,N_4618);
xnor U4894 (N_4894,N_4709,N_4653);
nand U4895 (N_4895,N_4789,N_4605);
xor U4896 (N_4896,N_4711,N_4690);
xor U4897 (N_4897,N_4708,N_4793);
and U4898 (N_4898,N_4636,N_4602);
or U4899 (N_4899,N_4616,N_4680);
nand U4900 (N_4900,N_4777,N_4646);
nand U4901 (N_4901,N_4670,N_4760);
and U4902 (N_4902,N_4784,N_4701);
xor U4903 (N_4903,N_4735,N_4634);
and U4904 (N_4904,N_4760,N_4771);
and U4905 (N_4905,N_4769,N_4708);
nand U4906 (N_4906,N_4720,N_4627);
or U4907 (N_4907,N_4657,N_4796);
nand U4908 (N_4908,N_4698,N_4757);
nor U4909 (N_4909,N_4765,N_4645);
nand U4910 (N_4910,N_4659,N_4702);
xnor U4911 (N_4911,N_4642,N_4652);
nor U4912 (N_4912,N_4646,N_4655);
or U4913 (N_4913,N_4614,N_4706);
nand U4914 (N_4914,N_4605,N_4767);
nand U4915 (N_4915,N_4770,N_4710);
xor U4916 (N_4916,N_4665,N_4626);
nand U4917 (N_4917,N_4619,N_4750);
nand U4918 (N_4918,N_4697,N_4705);
and U4919 (N_4919,N_4747,N_4754);
xor U4920 (N_4920,N_4655,N_4612);
xnor U4921 (N_4921,N_4664,N_4618);
nand U4922 (N_4922,N_4716,N_4746);
or U4923 (N_4923,N_4694,N_4696);
nand U4924 (N_4924,N_4728,N_4663);
xnor U4925 (N_4925,N_4635,N_4642);
xor U4926 (N_4926,N_4687,N_4660);
and U4927 (N_4927,N_4705,N_4693);
nor U4928 (N_4928,N_4618,N_4756);
nand U4929 (N_4929,N_4734,N_4704);
and U4930 (N_4930,N_4712,N_4703);
nor U4931 (N_4931,N_4604,N_4709);
nor U4932 (N_4932,N_4614,N_4725);
and U4933 (N_4933,N_4732,N_4645);
xor U4934 (N_4934,N_4759,N_4601);
xnor U4935 (N_4935,N_4638,N_4600);
or U4936 (N_4936,N_4652,N_4776);
nor U4937 (N_4937,N_4737,N_4604);
xor U4938 (N_4938,N_4613,N_4634);
xnor U4939 (N_4939,N_4601,N_4746);
nor U4940 (N_4940,N_4689,N_4637);
or U4941 (N_4941,N_4631,N_4784);
xnor U4942 (N_4942,N_4644,N_4745);
or U4943 (N_4943,N_4611,N_4663);
xor U4944 (N_4944,N_4695,N_4635);
nand U4945 (N_4945,N_4756,N_4750);
xor U4946 (N_4946,N_4745,N_4681);
and U4947 (N_4947,N_4718,N_4781);
and U4948 (N_4948,N_4737,N_4727);
and U4949 (N_4949,N_4678,N_4775);
xor U4950 (N_4950,N_4775,N_4604);
or U4951 (N_4951,N_4659,N_4641);
xnor U4952 (N_4952,N_4779,N_4667);
xor U4953 (N_4953,N_4706,N_4726);
nand U4954 (N_4954,N_4753,N_4718);
and U4955 (N_4955,N_4665,N_4673);
nand U4956 (N_4956,N_4670,N_4713);
nor U4957 (N_4957,N_4740,N_4675);
and U4958 (N_4958,N_4711,N_4669);
and U4959 (N_4959,N_4741,N_4772);
nand U4960 (N_4960,N_4790,N_4773);
or U4961 (N_4961,N_4728,N_4688);
xnor U4962 (N_4962,N_4781,N_4739);
nand U4963 (N_4963,N_4663,N_4602);
or U4964 (N_4964,N_4703,N_4781);
xnor U4965 (N_4965,N_4778,N_4745);
xor U4966 (N_4966,N_4634,N_4792);
or U4967 (N_4967,N_4753,N_4729);
nor U4968 (N_4968,N_4699,N_4626);
or U4969 (N_4969,N_4734,N_4631);
and U4970 (N_4970,N_4655,N_4781);
and U4971 (N_4971,N_4617,N_4740);
or U4972 (N_4972,N_4680,N_4744);
or U4973 (N_4973,N_4619,N_4621);
and U4974 (N_4974,N_4658,N_4709);
or U4975 (N_4975,N_4752,N_4799);
xor U4976 (N_4976,N_4616,N_4747);
nor U4977 (N_4977,N_4729,N_4658);
xnor U4978 (N_4978,N_4714,N_4711);
or U4979 (N_4979,N_4709,N_4766);
and U4980 (N_4980,N_4651,N_4737);
or U4981 (N_4981,N_4771,N_4619);
nand U4982 (N_4982,N_4708,N_4761);
nor U4983 (N_4983,N_4765,N_4640);
or U4984 (N_4984,N_4600,N_4723);
nand U4985 (N_4985,N_4732,N_4624);
nand U4986 (N_4986,N_4788,N_4692);
nand U4987 (N_4987,N_4666,N_4705);
nand U4988 (N_4988,N_4747,N_4638);
nor U4989 (N_4989,N_4628,N_4603);
nor U4990 (N_4990,N_4766,N_4748);
nor U4991 (N_4991,N_4628,N_4668);
or U4992 (N_4992,N_4786,N_4681);
nor U4993 (N_4993,N_4685,N_4624);
and U4994 (N_4994,N_4640,N_4625);
xnor U4995 (N_4995,N_4788,N_4752);
nand U4996 (N_4996,N_4714,N_4702);
xor U4997 (N_4997,N_4614,N_4684);
and U4998 (N_4998,N_4753,N_4758);
nor U4999 (N_4999,N_4652,N_4727);
xor UO_0 (O_0,N_4826,N_4885);
nand UO_1 (O_1,N_4933,N_4883);
nand UO_2 (O_2,N_4954,N_4907);
or UO_3 (O_3,N_4924,N_4974);
nand UO_4 (O_4,N_4937,N_4972);
nor UO_5 (O_5,N_4947,N_4876);
and UO_6 (O_6,N_4807,N_4917);
nand UO_7 (O_7,N_4943,N_4966);
xor UO_8 (O_8,N_4875,N_4898);
xnor UO_9 (O_9,N_4940,N_4890);
nand UO_10 (O_10,N_4993,N_4889);
xor UO_11 (O_11,N_4997,N_4989);
xnor UO_12 (O_12,N_4874,N_4801);
and UO_13 (O_13,N_4845,N_4920);
and UO_14 (O_14,N_4867,N_4922);
or UO_15 (O_15,N_4870,N_4970);
and UO_16 (O_16,N_4976,N_4809);
nor UO_17 (O_17,N_4873,N_4855);
xnor UO_18 (O_18,N_4952,N_4858);
nor UO_19 (O_19,N_4834,N_4900);
xnor UO_20 (O_20,N_4909,N_4854);
and UO_21 (O_21,N_4916,N_4880);
nor UO_22 (O_22,N_4981,N_4992);
nor UO_23 (O_23,N_4872,N_4859);
or UO_24 (O_24,N_4946,N_4939);
or UO_25 (O_25,N_4823,N_4921);
and UO_26 (O_26,N_4913,N_4914);
xor UO_27 (O_27,N_4986,N_4819);
xor UO_28 (O_28,N_4896,N_4948);
nand UO_29 (O_29,N_4848,N_4863);
and UO_30 (O_30,N_4959,N_4804);
xor UO_31 (O_31,N_4805,N_4886);
nor UO_32 (O_32,N_4967,N_4808);
nor UO_33 (O_33,N_4908,N_4864);
nor UO_34 (O_34,N_4998,N_4816);
nor UO_35 (O_35,N_4971,N_4847);
xnor UO_36 (O_36,N_4950,N_4868);
or UO_37 (O_37,N_4827,N_4911);
nor UO_38 (O_38,N_4927,N_4926);
nand UO_39 (O_39,N_4990,N_4860);
xor UO_40 (O_40,N_4892,N_4965);
or UO_41 (O_41,N_4824,N_4815);
nand UO_42 (O_42,N_4831,N_4853);
and UO_43 (O_43,N_4821,N_4849);
xnor UO_44 (O_44,N_4802,N_4983);
and UO_45 (O_45,N_4958,N_4929);
and UO_46 (O_46,N_4904,N_4811);
and UO_47 (O_47,N_4918,N_4931);
xor UO_48 (O_48,N_4941,N_4832);
or UO_49 (O_49,N_4882,N_4810);
or UO_50 (O_50,N_4866,N_4945);
nor UO_51 (O_51,N_4979,N_4957);
nand UO_52 (O_52,N_4961,N_4951);
xnor UO_53 (O_53,N_4830,N_4995);
xnor UO_54 (O_54,N_4835,N_4841);
xor UO_55 (O_55,N_4818,N_4894);
or UO_56 (O_56,N_4893,N_4851);
xor UO_57 (O_57,N_4915,N_4843);
nand UO_58 (O_58,N_4871,N_4846);
and UO_59 (O_59,N_4968,N_4923);
nand UO_60 (O_60,N_4985,N_4850);
xnor UO_61 (O_61,N_4852,N_4996);
xor UO_62 (O_62,N_4938,N_4991);
or UO_63 (O_63,N_4812,N_4833);
xor UO_64 (O_64,N_4877,N_4806);
xnor UO_65 (O_65,N_4865,N_4902);
nor UO_66 (O_66,N_4928,N_4964);
nor UO_67 (O_67,N_4925,N_4901);
nand UO_68 (O_68,N_4932,N_4977);
and UO_69 (O_69,N_4919,N_4978);
nand UO_70 (O_70,N_4973,N_4838);
xnor UO_71 (O_71,N_4839,N_4953);
or UO_72 (O_72,N_4905,N_4869);
nor UO_73 (O_73,N_4817,N_4829);
nand UO_74 (O_74,N_4862,N_4982);
and UO_75 (O_75,N_4857,N_4984);
xor UO_76 (O_76,N_4942,N_4844);
nor UO_77 (O_77,N_4969,N_4955);
nor UO_78 (O_78,N_4975,N_4814);
and UO_79 (O_79,N_4999,N_4912);
xor UO_80 (O_80,N_4856,N_4861);
and UO_81 (O_81,N_4836,N_4895);
nor UO_82 (O_82,N_4888,N_4891);
and UO_83 (O_83,N_4960,N_4879);
xor UO_84 (O_84,N_4837,N_4822);
nand UO_85 (O_85,N_4878,N_4994);
xor UO_86 (O_86,N_4987,N_4887);
nor UO_87 (O_87,N_4881,N_4825);
nand UO_88 (O_88,N_4903,N_4949);
nand UO_89 (O_89,N_4820,N_4963);
and UO_90 (O_90,N_4956,N_4897);
or UO_91 (O_91,N_4906,N_4884);
xor UO_92 (O_92,N_4899,N_4980);
or UO_93 (O_93,N_4840,N_4944);
nand UO_94 (O_94,N_4935,N_4800);
nor UO_95 (O_95,N_4962,N_4813);
nor UO_96 (O_96,N_4803,N_4934);
nand UO_97 (O_97,N_4842,N_4930);
or UO_98 (O_98,N_4988,N_4936);
nand UO_99 (O_99,N_4910,N_4828);
nand UO_100 (O_100,N_4813,N_4860);
nand UO_101 (O_101,N_4856,N_4870);
or UO_102 (O_102,N_4975,N_4939);
nand UO_103 (O_103,N_4914,N_4891);
nand UO_104 (O_104,N_4849,N_4840);
nor UO_105 (O_105,N_4993,N_4972);
and UO_106 (O_106,N_4860,N_4948);
nor UO_107 (O_107,N_4913,N_4806);
and UO_108 (O_108,N_4916,N_4984);
nand UO_109 (O_109,N_4807,N_4897);
nor UO_110 (O_110,N_4822,N_4828);
and UO_111 (O_111,N_4906,N_4971);
nand UO_112 (O_112,N_4883,N_4806);
xor UO_113 (O_113,N_4834,N_4970);
or UO_114 (O_114,N_4827,N_4988);
nand UO_115 (O_115,N_4980,N_4920);
nand UO_116 (O_116,N_4947,N_4992);
xor UO_117 (O_117,N_4835,N_4808);
and UO_118 (O_118,N_4982,N_4905);
or UO_119 (O_119,N_4841,N_4996);
nand UO_120 (O_120,N_4995,N_4897);
nand UO_121 (O_121,N_4855,N_4833);
nand UO_122 (O_122,N_4961,N_4882);
nor UO_123 (O_123,N_4904,N_4862);
or UO_124 (O_124,N_4880,N_4929);
xor UO_125 (O_125,N_4830,N_4902);
xor UO_126 (O_126,N_4929,N_4966);
nand UO_127 (O_127,N_4859,N_4889);
nor UO_128 (O_128,N_4973,N_4940);
or UO_129 (O_129,N_4810,N_4877);
or UO_130 (O_130,N_4842,N_4997);
nand UO_131 (O_131,N_4973,N_4981);
xor UO_132 (O_132,N_4813,N_4815);
xor UO_133 (O_133,N_4968,N_4819);
nor UO_134 (O_134,N_4915,N_4963);
nor UO_135 (O_135,N_4970,N_4934);
nand UO_136 (O_136,N_4857,N_4967);
and UO_137 (O_137,N_4800,N_4839);
or UO_138 (O_138,N_4895,N_4977);
and UO_139 (O_139,N_4804,N_4812);
xnor UO_140 (O_140,N_4843,N_4976);
xnor UO_141 (O_141,N_4892,N_4909);
or UO_142 (O_142,N_4981,N_4996);
nor UO_143 (O_143,N_4842,N_4869);
and UO_144 (O_144,N_4924,N_4837);
nor UO_145 (O_145,N_4955,N_4993);
or UO_146 (O_146,N_4920,N_4983);
and UO_147 (O_147,N_4844,N_4917);
and UO_148 (O_148,N_4980,N_4947);
nor UO_149 (O_149,N_4862,N_4827);
nand UO_150 (O_150,N_4978,N_4813);
xor UO_151 (O_151,N_4923,N_4854);
nand UO_152 (O_152,N_4984,N_4940);
or UO_153 (O_153,N_4847,N_4966);
or UO_154 (O_154,N_4805,N_4875);
nor UO_155 (O_155,N_4944,N_4963);
nor UO_156 (O_156,N_4885,N_4856);
nor UO_157 (O_157,N_4811,N_4926);
and UO_158 (O_158,N_4824,N_4858);
and UO_159 (O_159,N_4812,N_4967);
or UO_160 (O_160,N_4854,N_4829);
and UO_161 (O_161,N_4897,N_4870);
or UO_162 (O_162,N_4911,N_4886);
nand UO_163 (O_163,N_4824,N_4969);
xor UO_164 (O_164,N_4889,N_4981);
nor UO_165 (O_165,N_4866,N_4911);
nor UO_166 (O_166,N_4860,N_4941);
nand UO_167 (O_167,N_4935,N_4896);
xnor UO_168 (O_168,N_4897,N_4951);
or UO_169 (O_169,N_4961,N_4860);
or UO_170 (O_170,N_4842,N_4801);
and UO_171 (O_171,N_4992,N_4948);
xnor UO_172 (O_172,N_4818,N_4832);
or UO_173 (O_173,N_4944,N_4953);
nand UO_174 (O_174,N_4960,N_4911);
or UO_175 (O_175,N_4811,N_4825);
nor UO_176 (O_176,N_4849,N_4902);
or UO_177 (O_177,N_4804,N_4969);
or UO_178 (O_178,N_4898,N_4924);
nand UO_179 (O_179,N_4843,N_4831);
nand UO_180 (O_180,N_4976,N_4931);
nand UO_181 (O_181,N_4912,N_4867);
nor UO_182 (O_182,N_4964,N_4853);
and UO_183 (O_183,N_4980,N_4901);
xnor UO_184 (O_184,N_4891,N_4824);
nand UO_185 (O_185,N_4980,N_4846);
nor UO_186 (O_186,N_4868,N_4958);
and UO_187 (O_187,N_4806,N_4949);
nor UO_188 (O_188,N_4873,N_4991);
or UO_189 (O_189,N_4927,N_4921);
nand UO_190 (O_190,N_4850,N_4834);
or UO_191 (O_191,N_4936,N_4882);
and UO_192 (O_192,N_4917,N_4855);
or UO_193 (O_193,N_4891,N_4825);
or UO_194 (O_194,N_4802,N_4988);
or UO_195 (O_195,N_4878,N_4987);
or UO_196 (O_196,N_4856,N_4891);
or UO_197 (O_197,N_4994,N_4811);
xor UO_198 (O_198,N_4973,N_4909);
xnor UO_199 (O_199,N_4992,N_4881);
nor UO_200 (O_200,N_4877,N_4837);
nand UO_201 (O_201,N_4872,N_4878);
or UO_202 (O_202,N_4912,N_4820);
nand UO_203 (O_203,N_4814,N_4968);
nand UO_204 (O_204,N_4906,N_4902);
or UO_205 (O_205,N_4923,N_4941);
xor UO_206 (O_206,N_4980,N_4880);
nor UO_207 (O_207,N_4918,N_4917);
nor UO_208 (O_208,N_4989,N_4856);
nand UO_209 (O_209,N_4905,N_4908);
and UO_210 (O_210,N_4920,N_4851);
nor UO_211 (O_211,N_4811,N_4886);
or UO_212 (O_212,N_4805,N_4966);
or UO_213 (O_213,N_4836,N_4935);
xnor UO_214 (O_214,N_4961,N_4842);
nor UO_215 (O_215,N_4982,N_4896);
and UO_216 (O_216,N_4807,N_4836);
nand UO_217 (O_217,N_4919,N_4850);
nor UO_218 (O_218,N_4807,N_4948);
nand UO_219 (O_219,N_4914,N_4804);
nor UO_220 (O_220,N_4805,N_4870);
nand UO_221 (O_221,N_4869,N_4821);
and UO_222 (O_222,N_4826,N_4830);
and UO_223 (O_223,N_4817,N_4856);
and UO_224 (O_224,N_4860,N_4991);
xnor UO_225 (O_225,N_4834,N_4860);
xor UO_226 (O_226,N_4825,N_4863);
nand UO_227 (O_227,N_4801,N_4999);
and UO_228 (O_228,N_4955,N_4904);
nand UO_229 (O_229,N_4858,N_4862);
and UO_230 (O_230,N_4961,N_4806);
xnor UO_231 (O_231,N_4952,N_4878);
nor UO_232 (O_232,N_4973,N_4819);
or UO_233 (O_233,N_4877,N_4929);
xnor UO_234 (O_234,N_4963,N_4824);
and UO_235 (O_235,N_4964,N_4997);
or UO_236 (O_236,N_4815,N_4975);
nand UO_237 (O_237,N_4994,N_4881);
nor UO_238 (O_238,N_4843,N_4916);
or UO_239 (O_239,N_4893,N_4889);
and UO_240 (O_240,N_4828,N_4938);
or UO_241 (O_241,N_4835,N_4800);
and UO_242 (O_242,N_4900,N_4982);
and UO_243 (O_243,N_4871,N_4932);
nor UO_244 (O_244,N_4816,N_4885);
xnor UO_245 (O_245,N_4819,N_4938);
xor UO_246 (O_246,N_4910,N_4885);
xor UO_247 (O_247,N_4988,N_4925);
and UO_248 (O_248,N_4932,N_4873);
and UO_249 (O_249,N_4989,N_4909);
and UO_250 (O_250,N_4860,N_4821);
nand UO_251 (O_251,N_4931,N_4977);
or UO_252 (O_252,N_4856,N_4910);
xor UO_253 (O_253,N_4892,N_4882);
nand UO_254 (O_254,N_4983,N_4870);
xnor UO_255 (O_255,N_4924,N_4903);
xor UO_256 (O_256,N_4885,N_4835);
and UO_257 (O_257,N_4832,N_4964);
and UO_258 (O_258,N_4940,N_4821);
nor UO_259 (O_259,N_4800,N_4954);
nand UO_260 (O_260,N_4966,N_4836);
nor UO_261 (O_261,N_4953,N_4879);
and UO_262 (O_262,N_4808,N_4828);
xor UO_263 (O_263,N_4961,N_4832);
xnor UO_264 (O_264,N_4928,N_4949);
and UO_265 (O_265,N_4960,N_4941);
nor UO_266 (O_266,N_4889,N_4843);
and UO_267 (O_267,N_4905,N_4828);
nand UO_268 (O_268,N_4989,N_4836);
nor UO_269 (O_269,N_4852,N_4949);
nand UO_270 (O_270,N_4966,N_4865);
and UO_271 (O_271,N_4872,N_4991);
nor UO_272 (O_272,N_4819,N_4999);
nand UO_273 (O_273,N_4902,N_4919);
xnor UO_274 (O_274,N_4928,N_4954);
or UO_275 (O_275,N_4981,N_4972);
and UO_276 (O_276,N_4943,N_4956);
xnor UO_277 (O_277,N_4841,N_4891);
nor UO_278 (O_278,N_4956,N_4987);
xor UO_279 (O_279,N_4941,N_4954);
xnor UO_280 (O_280,N_4819,N_4936);
and UO_281 (O_281,N_4975,N_4805);
nand UO_282 (O_282,N_4960,N_4987);
nor UO_283 (O_283,N_4860,N_4981);
nor UO_284 (O_284,N_4945,N_4802);
nor UO_285 (O_285,N_4944,N_4868);
xnor UO_286 (O_286,N_4938,N_4942);
nor UO_287 (O_287,N_4852,N_4923);
nand UO_288 (O_288,N_4823,N_4889);
nand UO_289 (O_289,N_4837,N_4942);
or UO_290 (O_290,N_4838,N_4898);
nand UO_291 (O_291,N_4865,N_4973);
or UO_292 (O_292,N_4811,N_4814);
nor UO_293 (O_293,N_4859,N_4979);
nor UO_294 (O_294,N_4833,N_4938);
xnor UO_295 (O_295,N_4950,N_4808);
or UO_296 (O_296,N_4990,N_4804);
xnor UO_297 (O_297,N_4864,N_4898);
or UO_298 (O_298,N_4983,N_4949);
nand UO_299 (O_299,N_4950,N_4882);
and UO_300 (O_300,N_4817,N_4961);
nand UO_301 (O_301,N_4967,N_4935);
nand UO_302 (O_302,N_4941,N_4887);
nand UO_303 (O_303,N_4958,N_4883);
and UO_304 (O_304,N_4888,N_4980);
xnor UO_305 (O_305,N_4915,N_4904);
nand UO_306 (O_306,N_4841,N_4865);
and UO_307 (O_307,N_4869,N_4868);
or UO_308 (O_308,N_4967,N_4989);
nor UO_309 (O_309,N_4916,N_4898);
nand UO_310 (O_310,N_4969,N_4925);
or UO_311 (O_311,N_4812,N_4939);
xor UO_312 (O_312,N_4894,N_4918);
and UO_313 (O_313,N_4952,N_4911);
xnor UO_314 (O_314,N_4800,N_4947);
nand UO_315 (O_315,N_4968,N_4938);
xnor UO_316 (O_316,N_4968,N_4832);
nor UO_317 (O_317,N_4829,N_4943);
or UO_318 (O_318,N_4929,N_4995);
and UO_319 (O_319,N_4986,N_4927);
nor UO_320 (O_320,N_4841,N_4934);
nand UO_321 (O_321,N_4908,N_4888);
nand UO_322 (O_322,N_4862,N_4884);
xnor UO_323 (O_323,N_4874,N_4850);
nor UO_324 (O_324,N_4986,N_4834);
or UO_325 (O_325,N_4872,N_4892);
or UO_326 (O_326,N_4948,N_4856);
xnor UO_327 (O_327,N_4960,N_4917);
xor UO_328 (O_328,N_4933,N_4918);
or UO_329 (O_329,N_4891,N_4800);
or UO_330 (O_330,N_4810,N_4845);
nand UO_331 (O_331,N_4927,N_4939);
xnor UO_332 (O_332,N_4812,N_4872);
nand UO_333 (O_333,N_4864,N_4892);
nand UO_334 (O_334,N_4806,N_4832);
nand UO_335 (O_335,N_4883,N_4929);
and UO_336 (O_336,N_4946,N_4866);
or UO_337 (O_337,N_4812,N_4911);
nor UO_338 (O_338,N_4809,N_4963);
and UO_339 (O_339,N_4890,N_4930);
nor UO_340 (O_340,N_4990,N_4841);
xor UO_341 (O_341,N_4835,N_4872);
nor UO_342 (O_342,N_4817,N_4998);
xor UO_343 (O_343,N_4902,N_4961);
xor UO_344 (O_344,N_4836,N_4823);
xor UO_345 (O_345,N_4937,N_4924);
nand UO_346 (O_346,N_4870,N_4940);
nor UO_347 (O_347,N_4853,N_4930);
xor UO_348 (O_348,N_4826,N_4969);
nor UO_349 (O_349,N_4905,N_4916);
xor UO_350 (O_350,N_4810,N_4901);
xnor UO_351 (O_351,N_4811,N_4800);
xor UO_352 (O_352,N_4999,N_4811);
nand UO_353 (O_353,N_4930,N_4997);
nand UO_354 (O_354,N_4875,N_4849);
or UO_355 (O_355,N_4870,N_4945);
and UO_356 (O_356,N_4917,N_4819);
nand UO_357 (O_357,N_4907,N_4824);
nand UO_358 (O_358,N_4891,N_4973);
or UO_359 (O_359,N_4913,N_4829);
nor UO_360 (O_360,N_4947,N_4849);
or UO_361 (O_361,N_4883,N_4962);
xnor UO_362 (O_362,N_4824,N_4881);
xnor UO_363 (O_363,N_4978,N_4808);
xnor UO_364 (O_364,N_4920,N_4817);
nand UO_365 (O_365,N_4994,N_4852);
xnor UO_366 (O_366,N_4910,N_4845);
and UO_367 (O_367,N_4857,N_4916);
nor UO_368 (O_368,N_4867,N_4971);
nor UO_369 (O_369,N_4819,N_4969);
nor UO_370 (O_370,N_4933,N_4910);
nor UO_371 (O_371,N_4871,N_4907);
or UO_372 (O_372,N_4987,N_4805);
xor UO_373 (O_373,N_4864,N_4928);
and UO_374 (O_374,N_4859,N_4861);
or UO_375 (O_375,N_4896,N_4964);
nor UO_376 (O_376,N_4988,N_4904);
nor UO_377 (O_377,N_4936,N_4979);
nand UO_378 (O_378,N_4855,N_4822);
nand UO_379 (O_379,N_4948,N_4836);
or UO_380 (O_380,N_4909,N_4801);
or UO_381 (O_381,N_4851,N_4948);
xor UO_382 (O_382,N_4866,N_4931);
or UO_383 (O_383,N_4884,N_4895);
nand UO_384 (O_384,N_4865,N_4924);
nor UO_385 (O_385,N_4888,N_4813);
nand UO_386 (O_386,N_4979,N_4853);
xnor UO_387 (O_387,N_4810,N_4832);
or UO_388 (O_388,N_4829,N_4805);
nor UO_389 (O_389,N_4992,N_4885);
xnor UO_390 (O_390,N_4883,N_4997);
and UO_391 (O_391,N_4928,N_4847);
nand UO_392 (O_392,N_4929,N_4815);
and UO_393 (O_393,N_4837,N_4862);
nand UO_394 (O_394,N_4953,N_4888);
nand UO_395 (O_395,N_4857,N_4997);
nor UO_396 (O_396,N_4890,N_4921);
nor UO_397 (O_397,N_4973,N_4980);
nand UO_398 (O_398,N_4997,N_4918);
nor UO_399 (O_399,N_4867,N_4857);
nor UO_400 (O_400,N_4997,N_4992);
and UO_401 (O_401,N_4988,N_4919);
or UO_402 (O_402,N_4863,N_4943);
xnor UO_403 (O_403,N_4816,N_4962);
xor UO_404 (O_404,N_4881,N_4808);
or UO_405 (O_405,N_4968,N_4935);
and UO_406 (O_406,N_4807,N_4989);
or UO_407 (O_407,N_4863,N_4940);
or UO_408 (O_408,N_4810,N_4820);
or UO_409 (O_409,N_4942,N_4985);
xor UO_410 (O_410,N_4821,N_4968);
or UO_411 (O_411,N_4894,N_4806);
or UO_412 (O_412,N_4889,N_4983);
nand UO_413 (O_413,N_4934,N_4984);
and UO_414 (O_414,N_4850,N_4978);
nor UO_415 (O_415,N_4876,N_4820);
or UO_416 (O_416,N_4873,N_4836);
nand UO_417 (O_417,N_4859,N_4915);
nor UO_418 (O_418,N_4832,N_4809);
nand UO_419 (O_419,N_4940,N_4942);
and UO_420 (O_420,N_4858,N_4930);
nor UO_421 (O_421,N_4931,N_4912);
or UO_422 (O_422,N_4961,N_4920);
nor UO_423 (O_423,N_4860,N_4847);
nand UO_424 (O_424,N_4957,N_4811);
nor UO_425 (O_425,N_4834,N_4895);
xor UO_426 (O_426,N_4955,N_4911);
xor UO_427 (O_427,N_4812,N_4941);
xnor UO_428 (O_428,N_4957,N_4848);
nand UO_429 (O_429,N_4805,N_4971);
nor UO_430 (O_430,N_4834,N_4905);
nor UO_431 (O_431,N_4933,N_4834);
nor UO_432 (O_432,N_4853,N_4860);
and UO_433 (O_433,N_4963,N_4979);
nand UO_434 (O_434,N_4811,N_4818);
or UO_435 (O_435,N_4941,N_4805);
xor UO_436 (O_436,N_4920,N_4810);
nor UO_437 (O_437,N_4868,N_4824);
nor UO_438 (O_438,N_4894,N_4962);
nand UO_439 (O_439,N_4804,N_4995);
nor UO_440 (O_440,N_4843,N_4817);
nor UO_441 (O_441,N_4857,N_4877);
or UO_442 (O_442,N_4974,N_4877);
and UO_443 (O_443,N_4966,N_4963);
nor UO_444 (O_444,N_4897,N_4844);
and UO_445 (O_445,N_4935,N_4913);
and UO_446 (O_446,N_4955,N_4963);
nand UO_447 (O_447,N_4810,N_4937);
xor UO_448 (O_448,N_4847,N_4921);
and UO_449 (O_449,N_4946,N_4982);
nand UO_450 (O_450,N_4808,N_4937);
nand UO_451 (O_451,N_4851,N_4825);
and UO_452 (O_452,N_4901,N_4806);
or UO_453 (O_453,N_4872,N_4814);
or UO_454 (O_454,N_4836,N_4986);
or UO_455 (O_455,N_4959,N_4985);
nand UO_456 (O_456,N_4851,N_4876);
nand UO_457 (O_457,N_4946,N_4949);
or UO_458 (O_458,N_4805,N_4822);
nand UO_459 (O_459,N_4879,N_4965);
nor UO_460 (O_460,N_4883,N_4800);
and UO_461 (O_461,N_4987,N_4968);
xor UO_462 (O_462,N_4857,N_4887);
and UO_463 (O_463,N_4875,N_4986);
and UO_464 (O_464,N_4992,N_4967);
xor UO_465 (O_465,N_4990,N_4959);
nor UO_466 (O_466,N_4812,N_4801);
xor UO_467 (O_467,N_4862,N_4939);
nand UO_468 (O_468,N_4942,N_4859);
nor UO_469 (O_469,N_4866,N_4985);
xor UO_470 (O_470,N_4969,N_4844);
nand UO_471 (O_471,N_4944,N_4839);
nor UO_472 (O_472,N_4911,N_4873);
nand UO_473 (O_473,N_4930,N_4957);
xor UO_474 (O_474,N_4966,N_4992);
and UO_475 (O_475,N_4934,N_4891);
and UO_476 (O_476,N_4873,N_4999);
or UO_477 (O_477,N_4810,N_4874);
and UO_478 (O_478,N_4952,N_4922);
nor UO_479 (O_479,N_4910,N_4837);
and UO_480 (O_480,N_4970,N_4991);
nor UO_481 (O_481,N_4855,N_4987);
nand UO_482 (O_482,N_4820,N_4971);
and UO_483 (O_483,N_4924,N_4834);
xnor UO_484 (O_484,N_4937,N_4928);
and UO_485 (O_485,N_4976,N_4973);
nand UO_486 (O_486,N_4865,N_4925);
and UO_487 (O_487,N_4886,N_4906);
and UO_488 (O_488,N_4903,N_4890);
and UO_489 (O_489,N_4916,N_4802);
and UO_490 (O_490,N_4926,N_4866);
or UO_491 (O_491,N_4839,N_4811);
and UO_492 (O_492,N_4832,N_4875);
nand UO_493 (O_493,N_4819,N_4817);
and UO_494 (O_494,N_4844,N_4866);
nor UO_495 (O_495,N_4863,N_4894);
or UO_496 (O_496,N_4841,N_4827);
nand UO_497 (O_497,N_4946,N_4997);
nand UO_498 (O_498,N_4837,N_4933);
nor UO_499 (O_499,N_4977,N_4919);
and UO_500 (O_500,N_4892,N_4931);
or UO_501 (O_501,N_4950,N_4905);
xnor UO_502 (O_502,N_4966,N_4919);
and UO_503 (O_503,N_4914,N_4828);
nor UO_504 (O_504,N_4903,N_4827);
nor UO_505 (O_505,N_4803,N_4861);
nand UO_506 (O_506,N_4931,N_4848);
nand UO_507 (O_507,N_4998,N_4920);
nor UO_508 (O_508,N_4807,N_4854);
nor UO_509 (O_509,N_4850,N_4951);
or UO_510 (O_510,N_4859,N_4812);
nor UO_511 (O_511,N_4825,N_4937);
xnor UO_512 (O_512,N_4903,N_4950);
nor UO_513 (O_513,N_4959,N_4922);
or UO_514 (O_514,N_4983,N_4821);
or UO_515 (O_515,N_4882,N_4918);
xnor UO_516 (O_516,N_4928,N_4957);
or UO_517 (O_517,N_4938,N_4887);
nand UO_518 (O_518,N_4879,N_4860);
and UO_519 (O_519,N_4882,N_4836);
nand UO_520 (O_520,N_4832,N_4853);
xor UO_521 (O_521,N_4845,N_4870);
or UO_522 (O_522,N_4956,N_4991);
or UO_523 (O_523,N_4899,N_4936);
or UO_524 (O_524,N_4979,N_4836);
nand UO_525 (O_525,N_4966,N_4876);
and UO_526 (O_526,N_4988,N_4930);
or UO_527 (O_527,N_4929,N_4930);
nand UO_528 (O_528,N_4957,N_4838);
nand UO_529 (O_529,N_4840,N_4853);
and UO_530 (O_530,N_4811,N_4829);
nor UO_531 (O_531,N_4868,N_4853);
or UO_532 (O_532,N_4959,N_4930);
or UO_533 (O_533,N_4891,N_4910);
nand UO_534 (O_534,N_4960,N_4840);
xnor UO_535 (O_535,N_4803,N_4863);
nand UO_536 (O_536,N_4892,N_4920);
and UO_537 (O_537,N_4822,N_4905);
or UO_538 (O_538,N_4915,N_4822);
or UO_539 (O_539,N_4820,N_4822);
and UO_540 (O_540,N_4911,N_4917);
nor UO_541 (O_541,N_4866,N_4864);
nor UO_542 (O_542,N_4970,N_4967);
or UO_543 (O_543,N_4868,N_4941);
nor UO_544 (O_544,N_4804,N_4874);
or UO_545 (O_545,N_4970,N_4948);
nor UO_546 (O_546,N_4899,N_4986);
or UO_547 (O_547,N_4901,N_4986);
and UO_548 (O_548,N_4830,N_4920);
or UO_549 (O_549,N_4861,N_4983);
nand UO_550 (O_550,N_4925,N_4946);
and UO_551 (O_551,N_4887,N_4825);
xnor UO_552 (O_552,N_4902,N_4867);
xor UO_553 (O_553,N_4823,N_4991);
xor UO_554 (O_554,N_4889,N_4973);
xnor UO_555 (O_555,N_4871,N_4976);
nor UO_556 (O_556,N_4950,N_4949);
xnor UO_557 (O_557,N_4829,N_4816);
xnor UO_558 (O_558,N_4940,N_4944);
or UO_559 (O_559,N_4816,N_4887);
xor UO_560 (O_560,N_4830,N_4862);
nor UO_561 (O_561,N_4968,N_4936);
nor UO_562 (O_562,N_4999,N_4970);
nand UO_563 (O_563,N_4835,N_4856);
nand UO_564 (O_564,N_4922,N_4850);
xnor UO_565 (O_565,N_4811,N_4983);
xnor UO_566 (O_566,N_4961,N_4878);
or UO_567 (O_567,N_4816,N_4981);
and UO_568 (O_568,N_4915,N_4945);
nand UO_569 (O_569,N_4897,N_4874);
and UO_570 (O_570,N_4926,N_4879);
or UO_571 (O_571,N_4991,N_4818);
nor UO_572 (O_572,N_4874,N_4957);
and UO_573 (O_573,N_4958,N_4904);
and UO_574 (O_574,N_4804,N_4823);
and UO_575 (O_575,N_4949,N_4936);
xor UO_576 (O_576,N_4956,N_4955);
xnor UO_577 (O_577,N_4985,N_4926);
xnor UO_578 (O_578,N_4959,N_4925);
nand UO_579 (O_579,N_4975,N_4931);
nor UO_580 (O_580,N_4819,N_4984);
or UO_581 (O_581,N_4997,N_4926);
or UO_582 (O_582,N_4906,N_4929);
nor UO_583 (O_583,N_4958,N_4989);
nand UO_584 (O_584,N_4892,N_4993);
nand UO_585 (O_585,N_4819,N_4976);
nand UO_586 (O_586,N_4897,N_4816);
nand UO_587 (O_587,N_4923,N_4915);
nand UO_588 (O_588,N_4830,N_4900);
nand UO_589 (O_589,N_4932,N_4840);
or UO_590 (O_590,N_4868,N_4986);
nor UO_591 (O_591,N_4862,N_4969);
nand UO_592 (O_592,N_4823,N_4849);
nor UO_593 (O_593,N_4906,N_4935);
and UO_594 (O_594,N_4814,N_4866);
and UO_595 (O_595,N_4969,N_4894);
nor UO_596 (O_596,N_4935,N_4843);
nor UO_597 (O_597,N_4863,N_4950);
nor UO_598 (O_598,N_4914,N_4888);
or UO_599 (O_599,N_4836,N_4820);
nor UO_600 (O_600,N_4865,N_4904);
and UO_601 (O_601,N_4815,N_4820);
or UO_602 (O_602,N_4887,N_4885);
xor UO_603 (O_603,N_4819,N_4837);
nor UO_604 (O_604,N_4913,N_4862);
and UO_605 (O_605,N_4959,N_4940);
or UO_606 (O_606,N_4875,N_4868);
and UO_607 (O_607,N_4976,N_4874);
xnor UO_608 (O_608,N_4881,N_4815);
xor UO_609 (O_609,N_4991,N_4920);
xor UO_610 (O_610,N_4838,N_4978);
or UO_611 (O_611,N_4803,N_4883);
or UO_612 (O_612,N_4863,N_4946);
or UO_613 (O_613,N_4855,N_4967);
or UO_614 (O_614,N_4826,N_4919);
and UO_615 (O_615,N_4919,N_4805);
and UO_616 (O_616,N_4943,N_4808);
xnor UO_617 (O_617,N_4964,N_4890);
or UO_618 (O_618,N_4932,N_4969);
xnor UO_619 (O_619,N_4801,N_4951);
nand UO_620 (O_620,N_4901,N_4851);
nand UO_621 (O_621,N_4836,N_4808);
and UO_622 (O_622,N_4881,N_4897);
or UO_623 (O_623,N_4954,N_4963);
and UO_624 (O_624,N_4871,N_4926);
or UO_625 (O_625,N_4953,N_4805);
nor UO_626 (O_626,N_4978,N_4844);
and UO_627 (O_627,N_4975,N_4875);
nor UO_628 (O_628,N_4826,N_4837);
or UO_629 (O_629,N_4830,N_4943);
or UO_630 (O_630,N_4825,N_4894);
nor UO_631 (O_631,N_4815,N_4985);
xnor UO_632 (O_632,N_4804,N_4955);
and UO_633 (O_633,N_4927,N_4897);
nor UO_634 (O_634,N_4887,N_4976);
nand UO_635 (O_635,N_4874,N_4838);
or UO_636 (O_636,N_4969,N_4956);
and UO_637 (O_637,N_4802,N_4824);
and UO_638 (O_638,N_4830,N_4871);
nor UO_639 (O_639,N_4940,N_4826);
or UO_640 (O_640,N_4864,N_4834);
or UO_641 (O_641,N_4924,N_4867);
nor UO_642 (O_642,N_4815,N_4811);
xor UO_643 (O_643,N_4820,N_4808);
and UO_644 (O_644,N_4993,N_4876);
nand UO_645 (O_645,N_4883,N_4963);
nand UO_646 (O_646,N_4991,N_4808);
xor UO_647 (O_647,N_4957,N_4924);
nor UO_648 (O_648,N_4921,N_4977);
nor UO_649 (O_649,N_4963,N_4913);
nand UO_650 (O_650,N_4849,N_4950);
and UO_651 (O_651,N_4970,N_4922);
or UO_652 (O_652,N_4859,N_4958);
nand UO_653 (O_653,N_4979,N_4807);
nand UO_654 (O_654,N_4958,N_4937);
nor UO_655 (O_655,N_4963,N_4947);
and UO_656 (O_656,N_4932,N_4949);
or UO_657 (O_657,N_4829,N_4865);
nand UO_658 (O_658,N_4853,N_4928);
xor UO_659 (O_659,N_4885,N_4935);
nor UO_660 (O_660,N_4885,N_4805);
nand UO_661 (O_661,N_4983,N_4914);
nor UO_662 (O_662,N_4840,N_4966);
xor UO_663 (O_663,N_4903,N_4871);
xor UO_664 (O_664,N_4887,N_4876);
nand UO_665 (O_665,N_4810,N_4834);
xnor UO_666 (O_666,N_4987,N_4963);
or UO_667 (O_667,N_4989,N_4861);
or UO_668 (O_668,N_4994,N_4954);
nor UO_669 (O_669,N_4828,N_4923);
nand UO_670 (O_670,N_4813,N_4870);
or UO_671 (O_671,N_4830,N_4827);
nor UO_672 (O_672,N_4829,N_4864);
nand UO_673 (O_673,N_4836,N_4805);
or UO_674 (O_674,N_4848,N_4940);
or UO_675 (O_675,N_4918,N_4995);
and UO_676 (O_676,N_4907,N_4890);
and UO_677 (O_677,N_4961,N_4924);
xor UO_678 (O_678,N_4921,N_4986);
and UO_679 (O_679,N_4823,N_4884);
nor UO_680 (O_680,N_4858,N_4821);
and UO_681 (O_681,N_4987,N_4954);
nand UO_682 (O_682,N_4913,N_4921);
nor UO_683 (O_683,N_4923,N_4974);
or UO_684 (O_684,N_4962,N_4943);
nand UO_685 (O_685,N_4864,N_4852);
nor UO_686 (O_686,N_4914,N_4901);
and UO_687 (O_687,N_4937,N_4866);
xor UO_688 (O_688,N_4983,N_4972);
xor UO_689 (O_689,N_4996,N_4926);
or UO_690 (O_690,N_4850,N_4806);
or UO_691 (O_691,N_4877,N_4848);
nand UO_692 (O_692,N_4895,N_4864);
nand UO_693 (O_693,N_4992,N_4904);
nor UO_694 (O_694,N_4829,N_4924);
xnor UO_695 (O_695,N_4899,N_4985);
nand UO_696 (O_696,N_4913,N_4865);
nand UO_697 (O_697,N_4862,N_4953);
xor UO_698 (O_698,N_4816,N_4963);
and UO_699 (O_699,N_4973,N_4907);
nand UO_700 (O_700,N_4811,N_4856);
and UO_701 (O_701,N_4964,N_4972);
nand UO_702 (O_702,N_4854,N_4963);
xor UO_703 (O_703,N_4901,N_4896);
or UO_704 (O_704,N_4905,N_4918);
nor UO_705 (O_705,N_4991,N_4907);
nand UO_706 (O_706,N_4867,N_4861);
or UO_707 (O_707,N_4947,N_4890);
and UO_708 (O_708,N_4874,N_4960);
nand UO_709 (O_709,N_4939,N_4895);
or UO_710 (O_710,N_4900,N_4864);
nand UO_711 (O_711,N_4976,N_4853);
or UO_712 (O_712,N_4918,N_4996);
nand UO_713 (O_713,N_4804,N_4999);
nor UO_714 (O_714,N_4967,N_4860);
and UO_715 (O_715,N_4907,N_4914);
and UO_716 (O_716,N_4813,N_4862);
nand UO_717 (O_717,N_4973,N_4960);
nand UO_718 (O_718,N_4907,N_4996);
xor UO_719 (O_719,N_4842,N_4858);
xnor UO_720 (O_720,N_4886,N_4933);
and UO_721 (O_721,N_4848,N_4932);
and UO_722 (O_722,N_4910,N_4941);
or UO_723 (O_723,N_4877,N_4911);
xnor UO_724 (O_724,N_4860,N_4952);
nor UO_725 (O_725,N_4898,N_4856);
nor UO_726 (O_726,N_4892,N_4806);
nor UO_727 (O_727,N_4908,N_4915);
nand UO_728 (O_728,N_4982,N_4870);
nand UO_729 (O_729,N_4922,N_4842);
and UO_730 (O_730,N_4871,N_4952);
or UO_731 (O_731,N_4988,N_4880);
and UO_732 (O_732,N_4883,N_4828);
nor UO_733 (O_733,N_4896,N_4840);
nand UO_734 (O_734,N_4939,N_4873);
xnor UO_735 (O_735,N_4924,N_4917);
nand UO_736 (O_736,N_4989,N_4896);
nor UO_737 (O_737,N_4914,N_4930);
xnor UO_738 (O_738,N_4816,N_4832);
or UO_739 (O_739,N_4953,N_4820);
and UO_740 (O_740,N_4886,N_4968);
xnor UO_741 (O_741,N_4918,N_4907);
or UO_742 (O_742,N_4903,N_4948);
nor UO_743 (O_743,N_4889,N_4985);
xor UO_744 (O_744,N_4892,N_4848);
or UO_745 (O_745,N_4978,N_4848);
nor UO_746 (O_746,N_4855,N_4970);
and UO_747 (O_747,N_4959,N_4807);
nor UO_748 (O_748,N_4838,N_4853);
or UO_749 (O_749,N_4976,N_4810);
or UO_750 (O_750,N_4808,N_4935);
or UO_751 (O_751,N_4972,N_4958);
nand UO_752 (O_752,N_4886,N_4841);
or UO_753 (O_753,N_4832,N_4811);
xnor UO_754 (O_754,N_4885,N_4811);
nand UO_755 (O_755,N_4944,N_4802);
xor UO_756 (O_756,N_4869,N_4985);
nand UO_757 (O_757,N_4952,N_4853);
and UO_758 (O_758,N_4966,N_4944);
nor UO_759 (O_759,N_4982,N_4927);
nand UO_760 (O_760,N_4900,N_4804);
or UO_761 (O_761,N_4994,N_4894);
or UO_762 (O_762,N_4926,N_4880);
or UO_763 (O_763,N_4838,N_4862);
and UO_764 (O_764,N_4924,N_4955);
nand UO_765 (O_765,N_4986,N_4912);
or UO_766 (O_766,N_4968,N_4895);
xor UO_767 (O_767,N_4909,N_4940);
nor UO_768 (O_768,N_4902,N_4989);
nand UO_769 (O_769,N_4971,N_4902);
or UO_770 (O_770,N_4966,N_4980);
nor UO_771 (O_771,N_4812,N_4995);
nor UO_772 (O_772,N_4979,N_4843);
and UO_773 (O_773,N_4980,N_4910);
nor UO_774 (O_774,N_4927,N_4878);
and UO_775 (O_775,N_4987,N_4971);
nor UO_776 (O_776,N_4901,N_4918);
nor UO_777 (O_777,N_4938,N_4927);
xnor UO_778 (O_778,N_4812,N_4860);
xor UO_779 (O_779,N_4829,N_4933);
xnor UO_780 (O_780,N_4918,N_4908);
nor UO_781 (O_781,N_4881,N_4987);
and UO_782 (O_782,N_4990,N_4840);
xnor UO_783 (O_783,N_4983,N_4855);
or UO_784 (O_784,N_4878,N_4856);
nand UO_785 (O_785,N_4918,N_4990);
nor UO_786 (O_786,N_4897,N_4818);
nand UO_787 (O_787,N_4910,N_4871);
nor UO_788 (O_788,N_4823,N_4914);
and UO_789 (O_789,N_4834,N_4910);
and UO_790 (O_790,N_4865,N_4937);
nor UO_791 (O_791,N_4868,N_4862);
and UO_792 (O_792,N_4967,N_4895);
or UO_793 (O_793,N_4883,N_4805);
nand UO_794 (O_794,N_4887,N_4898);
and UO_795 (O_795,N_4954,N_4876);
or UO_796 (O_796,N_4857,N_4830);
or UO_797 (O_797,N_4849,N_4866);
xnor UO_798 (O_798,N_4944,N_4943);
nand UO_799 (O_799,N_4851,N_4871);
nand UO_800 (O_800,N_4977,N_4924);
and UO_801 (O_801,N_4962,N_4915);
nor UO_802 (O_802,N_4950,N_4876);
nand UO_803 (O_803,N_4811,N_4914);
and UO_804 (O_804,N_4965,N_4849);
and UO_805 (O_805,N_4931,N_4982);
nor UO_806 (O_806,N_4990,N_4829);
nor UO_807 (O_807,N_4811,N_4860);
nor UO_808 (O_808,N_4893,N_4811);
nor UO_809 (O_809,N_4805,N_4994);
or UO_810 (O_810,N_4819,N_4865);
or UO_811 (O_811,N_4972,N_4907);
xor UO_812 (O_812,N_4967,N_4891);
or UO_813 (O_813,N_4862,N_4981);
nand UO_814 (O_814,N_4931,N_4864);
nor UO_815 (O_815,N_4852,N_4866);
nand UO_816 (O_816,N_4851,N_4956);
and UO_817 (O_817,N_4967,N_4914);
and UO_818 (O_818,N_4891,N_4928);
xor UO_819 (O_819,N_4922,N_4861);
nor UO_820 (O_820,N_4959,N_4839);
and UO_821 (O_821,N_4903,N_4852);
or UO_822 (O_822,N_4924,N_4991);
nand UO_823 (O_823,N_4835,N_4868);
xnor UO_824 (O_824,N_4822,N_4863);
nor UO_825 (O_825,N_4904,N_4882);
xor UO_826 (O_826,N_4962,N_4856);
nor UO_827 (O_827,N_4839,N_4828);
nor UO_828 (O_828,N_4946,N_4948);
and UO_829 (O_829,N_4996,N_4847);
nor UO_830 (O_830,N_4853,N_4960);
nand UO_831 (O_831,N_4823,N_4957);
or UO_832 (O_832,N_4858,N_4991);
nand UO_833 (O_833,N_4913,N_4888);
nor UO_834 (O_834,N_4918,N_4831);
nor UO_835 (O_835,N_4836,N_4826);
and UO_836 (O_836,N_4841,N_4822);
and UO_837 (O_837,N_4874,N_4919);
xnor UO_838 (O_838,N_4809,N_4918);
or UO_839 (O_839,N_4977,N_4926);
and UO_840 (O_840,N_4923,N_4839);
and UO_841 (O_841,N_4980,N_4832);
and UO_842 (O_842,N_4931,N_4890);
nor UO_843 (O_843,N_4855,N_4854);
and UO_844 (O_844,N_4878,N_4908);
nand UO_845 (O_845,N_4930,N_4933);
xor UO_846 (O_846,N_4890,N_4924);
xor UO_847 (O_847,N_4853,N_4922);
or UO_848 (O_848,N_4818,N_4884);
and UO_849 (O_849,N_4846,N_4996);
xnor UO_850 (O_850,N_4839,N_4922);
nand UO_851 (O_851,N_4986,N_4807);
or UO_852 (O_852,N_4959,N_4978);
or UO_853 (O_853,N_4901,N_4842);
nor UO_854 (O_854,N_4922,N_4857);
nor UO_855 (O_855,N_4998,N_4865);
nand UO_856 (O_856,N_4817,N_4852);
or UO_857 (O_857,N_4954,N_4887);
or UO_858 (O_858,N_4961,N_4863);
xor UO_859 (O_859,N_4833,N_4940);
nand UO_860 (O_860,N_4879,N_4899);
and UO_861 (O_861,N_4947,N_4935);
and UO_862 (O_862,N_4993,N_4853);
nor UO_863 (O_863,N_4835,N_4960);
xnor UO_864 (O_864,N_4832,N_4967);
nand UO_865 (O_865,N_4887,N_4951);
xnor UO_866 (O_866,N_4835,N_4880);
nor UO_867 (O_867,N_4978,N_4801);
or UO_868 (O_868,N_4935,N_4841);
nor UO_869 (O_869,N_4944,N_4850);
or UO_870 (O_870,N_4800,N_4958);
and UO_871 (O_871,N_4800,N_4869);
nor UO_872 (O_872,N_4915,N_4833);
and UO_873 (O_873,N_4968,N_4826);
nor UO_874 (O_874,N_4987,N_4843);
nand UO_875 (O_875,N_4989,N_4995);
nor UO_876 (O_876,N_4849,N_4844);
or UO_877 (O_877,N_4859,N_4874);
xor UO_878 (O_878,N_4874,N_4814);
nand UO_879 (O_879,N_4991,N_4983);
nor UO_880 (O_880,N_4952,N_4954);
nand UO_881 (O_881,N_4832,N_4886);
or UO_882 (O_882,N_4892,N_4899);
or UO_883 (O_883,N_4835,N_4908);
and UO_884 (O_884,N_4958,N_4878);
or UO_885 (O_885,N_4841,N_4877);
xnor UO_886 (O_886,N_4954,N_4835);
nand UO_887 (O_887,N_4917,N_4954);
xor UO_888 (O_888,N_4821,N_4967);
nor UO_889 (O_889,N_4927,N_4947);
nand UO_890 (O_890,N_4898,N_4834);
and UO_891 (O_891,N_4976,N_4938);
or UO_892 (O_892,N_4974,N_4878);
nor UO_893 (O_893,N_4850,N_4881);
and UO_894 (O_894,N_4899,N_4849);
xor UO_895 (O_895,N_4965,N_4954);
xor UO_896 (O_896,N_4974,N_4945);
and UO_897 (O_897,N_4863,N_4873);
and UO_898 (O_898,N_4914,N_4996);
nand UO_899 (O_899,N_4920,N_4929);
xnor UO_900 (O_900,N_4883,N_4824);
xnor UO_901 (O_901,N_4975,N_4823);
or UO_902 (O_902,N_4881,N_4915);
nor UO_903 (O_903,N_4901,N_4911);
nor UO_904 (O_904,N_4896,N_4999);
nand UO_905 (O_905,N_4876,N_4829);
nand UO_906 (O_906,N_4931,N_4891);
nand UO_907 (O_907,N_4912,N_4858);
nor UO_908 (O_908,N_4996,N_4901);
xor UO_909 (O_909,N_4881,N_4839);
nand UO_910 (O_910,N_4935,N_4824);
nand UO_911 (O_911,N_4929,N_4942);
or UO_912 (O_912,N_4862,N_4930);
and UO_913 (O_913,N_4974,N_4839);
xnor UO_914 (O_914,N_4928,N_4983);
xnor UO_915 (O_915,N_4821,N_4941);
nand UO_916 (O_916,N_4804,N_4847);
and UO_917 (O_917,N_4886,N_4971);
and UO_918 (O_918,N_4842,N_4834);
xnor UO_919 (O_919,N_4814,N_4887);
nand UO_920 (O_920,N_4895,N_4890);
nor UO_921 (O_921,N_4993,N_4909);
or UO_922 (O_922,N_4948,N_4942);
and UO_923 (O_923,N_4991,N_4871);
nand UO_924 (O_924,N_4805,N_4804);
or UO_925 (O_925,N_4845,N_4868);
nor UO_926 (O_926,N_4875,N_4847);
or UO_927 (O_927,N_4859,N_4807);
xnor UO_928 (O_928,N_4911,N_4897);
xnor UO_929 (O_929,N_4952,N_4988);
xor UO_930 (O_930,N_4822,N_4803);
xor UO_931 (O_931,N_4872,N_4851);
or UO_932 (O_932,N_4919,N_4839);
nor UO_933 (O_933,N_4933,N_4959);
nand UO_934 (O_934,N_4963,N_4880);
xor UO_935 (O_935,N_4919,N_4908);
nor UO_936 (O_936,N_4869,N_4870);
and UO_937 (O_937,N_4914,N_4851);
nand UO_938 (O_938,N_4869,N_4986);
and UO_939 (O_939,N_4874,N_4956);
or UO_940 (O_940,N_4885,N_4823);
or UO_941 (O_941,N_4800,N_4911);
and UO_942 (O_942,N_4918,N_4873);
nand UO_943 (O_943,N_4963,N_4855);
and UO_944 (O_944,N_4995,N_4955);
xor UO_945 (O_945,N_4980,N_4854);
and UO_946 (O_946,N_4831,N_4935);
xnor UO_947 (O_947,N_4830,N_4969);
xor UO_948 (O_948,N_4847,N_4923);
nand UO_949 (O_949,N_4800,N_4907);
or UO_950 (O_950,N_4946,N_4825);
nor UO_951 (O_951,N_4948,N_4982);
xor UO_952 (O_952,N_4927,N_4856);
nor UO_953 (O_953,N_4907,N_4848);
nor UO_954 (O_954,N_4832,N_4913);
nor UO_955 (O_955,N_4868,N_4884);
xnor UO_956 (O_956,N_4809,N_4909);
nand UO_957 (O_957,N_4970,N_4952);
and UO_958 (O_958,N_4948,N_4925);
nor UO_959 (O_959,N_4830,N_4808);
and UO_960 (O_960,N_4878,N_4805);
nor UO_961 (O_961,N_4886,N_4935);
nand UO_962 (O_962,N_4950,N_4806);
or UO_963 (O_963,N_4952,N_4828);
xor UO_964 (O_964,N_4818,N_4952);
nor UO_965 (O_965,N_4856,N_4859);
nor UO_966 (O_966,N_4804,N_4814);
xnor UO_967 (O_967,N_4812,N_4977);
nand UO_968 (O_968,N_4906,N_4821);
nor UO_969 (O_969,N_4883,N_4995);
xor UO_970 (O_970,N_4952,N_4893);
nand UO_971 (O_971,N_4861,N_4929);
and UO_972 (O_972,N_4982,N_4800);
nor UO_973 (O_973,N_4920,N_4889);
xor UO_974 (O_974,N_4835,N_4822);
or UO_975 (O_975,N_4867,N_4892);
xor UO_976 (O_976,N_4834,N_4996);
nand UO_977 (O_977,N_4933,N_4832);
or UO_978 (O_978,N_4852,N_4940);
nor UO_979 (O_979,N_4883,N_4886);
nor UO_980 (O_980,N_4806,N_4842);
and UO_981 (O_981,N_4998,N_4800);
and UO_982 (O_982,N_4924,N_4920);
or UO_983 (O_983,N_4802,N_4937);
nor UO_984 (O_984,N_4944,N_4975);
nand UO_985 (O_985,N_4953,N_4983);
nand UO_986 (O_986,N_4848,N_4800);
and UO_987 (O_987,N_4914,N_4800);
and UO_988 (O_988,N_4860,N_4964);
nand UO_989 (O_989,N_4815,N_4902);
or UO_990 (O_990,N_4932,N_4899);
nor UO_991 (O_991,N_4915,N_4890);
or UO_992 (O_992,N_4952,N_4931);
xnor UO_993 (O_993,N_4861,N_4909);
nand UO_994 (O_994,N_4965,N_4989);
nand UO_995 (O_995,N_4851,N_4836);
or UO_996 (O_996,N_4903,N_4952);
and UO_997 (O_997,N_4936,N_4961);
xor UO_998 (O_998,N_4813,N_4852);
or UO_999 (O_999,N_4923,N_4858);
endmodule