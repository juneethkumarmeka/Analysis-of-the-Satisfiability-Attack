module basic_3000_30000_3500_25_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_163,In_1267);
nor U1 (N_1,In_2667,In_236);
xor U2 (N_2,In_2059,In_957);
and U3 (N_3,In_2570,In_616);
nor U4 (N_4,In_2226,In_1236);
nand U5 (N_5,In_2680,In_2674);
xnor U6 (N_6,In_1810,In_842);
nor U7 (N_7,In_2678,In_1685);
xor U8 (N_8,In_2320,In_1582);
nor U9 (N_9,In_1822,In_2697);
nand U10 (N_10,In_1596,In_1655);
and U11 (N_11,In_978,In_1766);
xor U12 (N_12,In_643,In_2445);
xnor U13 (N_13,In_1371,In_1790);
xnor U14 (N_14,In_412,In_1748);
nand U15 (N_15,In_594,In_2301);
and U16 (N_16,In_2143,In_1797);
or U17 (N_17,In_503,In_883);
xnor U18 (N_18,In_2398,In_2677);
nand U19 (N_19,In_2189,In_1778);
and U20 (N_20,In_2275,In_1800);
nand U21 (N_21,In_2400,In_2103);
or U22 (N_22,In_1681,In_683);
xor U23 (N_23,In_2425,In_2050);
xnor U24 (N_24,In_2018,In_2240);
nand U25 (N_25,In_623,In_2638);
or U26 (N_26,In_1429,In_1974);
or U27 (N_27,In_1498,In_1409);
and U28 (N_28,In_2549,In_2187);
xor U29 (N_29,In_231,In_1883);
nand U30 (N_30,In_411,In_2727);
xnor U31 (N_31,In_2604,In_2192);
and U32 (N_32,In_2666,In_1437);
nor U33 (N_33,In_521,In_1198);
and U34 (N_34,In_53,In_155);
or U35 (N_35,In_34,In_180);
and U36 (N_36,In_0,In_2113);
and U37 (N_37,In_456,In_644);
nor U38 (N_38,In_637,In_580);
and U39 (N_39,In_119,In_221);
xor U40 (N_40,In_906,In_2941);
xnor U41 (N_41,In_914,In_1093);
nor U42 (N_42,In_1297,In_1895);
xnor U43 (N_43,In_1721,In_426);
nor U44 (N_44,In_2183,In_2536);
or U45 (N_45,In_543,In_125);
nor U46 (N_46,In_800,In_2860);
nor U47 (N_47,In_1204,In_559);
nand U48 (N_48,In_2816,In_1563);
nor U49 (N_49,In_312,In_2488);
nand U50 (N_50,In_112,In_2648);
nand U51 (N_51,In_463,In_1641);
or U52 (N_52,In_2831,In_1570);
or U53 (N_53,In_2055,In_81);
nand U54 (N_54,In_2950,In_2938);
and U55 (N_55,In_361,In_63);
xnor U56 (N_56,In_573,In_2136);
or U57 (N_57,In_550,In_628);
or U58 (N_58,In_586,In_1406);
or U59 (N_59,In_2498,In_2151);
or U60 (N_60,In_4,In_1849);
or U61 (N_61,In_1864,In_1359);
and U62 (N_62,In_868,In_294);
and U63 (N_63,In_28,In_2550);
nand U64 (N_64,In_1009,In_1287);
or U65 (N_65,In_67,In_1414);
nand U66 (N_66,In_1842,In_1456);
nand U67 (N_67,In_2042,In_513);
nand U68 (N_68,In_590,In_38);
xnor U69 (N_69,In_2568,In_1256);
nand U70 (N_70,In_2842,In_2758);
and U71 (N_71,In_2595,In_494);
xor U72 (N_72,In_2464,In_1686);
or U73 (N_73,In_760,In_2813);
or U74 (N_74,In_1179,In_187);
and U75 (N_75,In_2646,In_2088);
or U76 (N_76,In_871,In_2476);
xnor U77 (N_77,In_753,In_735);
and U78 (N_78,In_2991,In_1891);
nand U79 (N_79,In_2807,In_1869);
and U80 (N_80,In_296,In_2964);
nand U81 (N_81,In_1909,In_799);
or U82 (N_82,In_624,In_416);
xor U83 (N_83,In_2242,In_1464);
and U84 (N_84,In_2659,In_1283);
nand U85 (N_85,In_2628,In_828);
nand U86 (N_86,In_876,In_1615);
nand U87 (N_87,In_424,In_1779);
nand U88 (N_88,In_2021,In_1701);
or U89 (N_89,In_2267,In_1759);
nor U90 (N_90,In_2499,In_94);
or U91 (N_91,In_2695,In_757);
and U92 (N_92,In_1704,In_583);
or U93 (N_93,In_572,In_659);
or U94 (N_94,In_227,In_2120);
nor U95 (N_95,In_62,In_529);
or U96 (N_96,In_452,In_425);
xor U97 (N_97,In_266,In_2041);
nor U98 (N_98,In_1330,In_154);
or U99 (N_99,In_1404,In_2717);
nor U100 (N_100,In_2401,In_913);
or U101 (N_101,In_1194,In_1460);
and U102 (N_102,In_1938,In_2794);
xnor U103 (N_103,In_1426,In_2539);
or U104 (N_104,In_2239,In_158);
or U105 (N_105,In_1657,In_390);
or U106 (N_106,In_540,In_556);
nand U107 (N_107,In_1059,In_1774);
and U108 (N_108,In_974,In_2161);
and U109 (N_109,In_1934,In_863);
xnor U110 (N_110,In_304,In_866);
nor U111 (N_111,In_1033,In_2289);
nor U112 (N_112,In_2959,In_339);
nor U113 (N_113,In_1691,In_1226);
or U114 (N_114,In_2204,In_2116);
and U115 (N_115,In_164,In_1468);
nand U116 (N_116,In_2428,In_781);
or U117 (N_117,In_1591,In_332);
or U118 (N_118,In_1408,In_2332);
xor U119 (N_119,In_1858,In_1699);
and U120 (N_120,In_551,In_912);
nand U121 (N_121,In_2034,In_496);
nor U122 (N_122,In_2821,In_2869);
or U123 (N_123,In_1875,In_171);
xnor U124 (N_124,In_442,In_1967);
nor U125 (N_125,In_1035,In_2708);
nor U126 (N_126,In_1863,In_1567);
nand U127 (N_127,In_2827,In_310);
xnor U128 (N_128,In_1162,In_1343);
nor U129 (N_129,In_208,In_1061);
xor U130 (N_130,In_1036,In_2736);
xor U131 (N_131,In_83,In_405);
xor U132 (N_132,In_1474,In_629);
nor U133 (N_133,In_1349,In_2764);
and U134 (N_134,In_2801,In_1525);
or U135 (N_135,In_1131,In_1542);
nand U136 (N_136,In_2981,In_2925);
or U137 (N_137,In_1240,In_2494);
or U138 (N_138,In_730,In_734);
nor U139 (N_139,In_2265,In_141);
xnor U140 (N_140,In_1105,In_609);
nor U141 (N_141,In_273,In_1140);
or U142 (N_142,In_1756,In_1451);
and U143 (N_143,In_718,In_2802);
nor U144 (N_144,In_2343,In_1788);
xnor U145 (N_145,In_2026,In_277);
xor U146 (N_146,In_1363,In_2507);
nand U147 (N_147,In_545,In_1928);
nand U148 (N_148,In_89,In_1682);
or U149 (N_149,In_1002,In_2745);
nand U150 (N_150,In_1637,In_2729);
xnor U151 (N_151,In_432,In_2030);
xnor U152 (N_152,In_2641,In_2215);
nand U153 (N_153,In_1167,In_2109);
nand U154 (N_154,In_832,In_1357);
or U155 (N_155,In_1802,In_938);
and U156 (N_156,In_697,In_2993);
or U157 (N_157,In_2108,In_2490);
nand U158 (N_158,In_2027,In_2791);
and U159 (N_159,In_449,In_1975);
xnor U160 (N_160,In_2497,In_1234);
and U161 (N_161,In_1344,In_1057);
and U162 (N_162,In_809,In_2255);
xnor U163 (N_163,In_2538,In_998);
and U164 (N_164,In_1811,In_33);
and U165 (N_165,In_2773,In_2508);
xnor U166 (N_166,In_1830,In_910);
and U167 (N_167,In_126,In_2923);
or U168 (N_168,In_1430,In_1558);
nor U169 (N_169,In_1207,In_380);
nor U170 (N_170,In_554,In_2503);
and U171 (N_171,In_2890,In_387);
or U172 (N_172,In_983,In_1051);
nand U173 (N_173,In_363,In_2790);
nand U174 (N_174,In_245,In_2062);
and U175 (N_175,In_627,In_1834);
or U176 (N_176,In_585,In_2184);
xnor U177 (N_177,In_2412,In_2430);
nor U178 (N_178,In_1049,In_2954);
xnor U179 (N_179,In_2943,In_1719);
nor U180 (N_180,In_896,In_2937);
nor U181 (N_181,In_2312,In_74);
and U182 (N_182,In_473,In_1702);
xnor U183 (N_183,In_1076,In_996);
nor U184 (N_184,In_860,In_2979);
xor U185 (N_185,In_2098,In_2714);
nor U186 (N_186,In_2968,In_1614);
and U187 (N_187,In_2087,In_885);
xnor U188 (N_188,In_2838,In_1754);
nand U189 (N_189,In_2957,In_1020);
and U190 (N_190,In_1899,In_1770);
nand U191 (N_191,In_861,In_691);
or U192 (N_192,In_2453,In_2721);
or U193 (N_193,In_2726,In_10);
nor U194 (N_194,In_2894,In_1878);
nand U195 (N_195,In_981,In_640);
or U196 (N_196,In_2160,In_1042);
nor U197 (N_197,In_140,In_2367);
nor U198 (N_198,In_688,In_1218);
and U199 (N_199,In_1262,In_929);
nor U200 (N_200,In_2602,In_1116);
and U201 (N_201,In_143,In_936);
nor U202 (N_202,In_2610,In_531);
or U203 (N_203,In_642,In_1106);
or U204 (N_204,In_1896,In_462);
nand U205 (N_205,In_2107,In_232);
xnor U206 (N_206,In_127,In_2075);
and U207 (N_207,In_1734,In_104);
nor U208 (N_208,In_530,In_1978);
nor U209 (N_209,In_2211,In_1643);
nor U210 (N_210,In_490,In_2715);
or U211 (N_211,In_2933,In_2693);
xnor U212 (N_212,In_142,In_173);
nand U213 (N_213,In_2070,In_1543);
nor U214 (N_214,In_2371,In_1271);
xnor U215 (N_215,In_2156,In_2663);
xor U216 (N_216,In_536,In_1238);
or U217 (N_217,In_2634,In_88);
nand U218 (N_218,In_2895,In_409);
xor U219 (N_219,In_2148,In_1177);
nand U220 (N_220,In_1332,In_907);
xor U221 (N_221,In_2482,In_1765);
or U222 (N_222,In_1160,In_1624);
nor U223 (N_223,In_2295,In_1399);
or U224 (N_224,In_1170,In_1027);
xor U225 (N_225,In_1744,In_2131);
nand U226 (N_226,In_93,In_1239);
and U227 (N_227,In_1016,In_570);
nand U228 (N_228,In_2125,In_737);
and U229 (N_229,In_909,In_1678);
xor U230 (N_230,In_2571,In_565);
nand U231 (N_231,In_774,In_618);
nand U232 (N_232,In_631,In_2);
or U233 (N_233,In_2718,In_450);
and U234 (N_234,In_1783,In_2637);
and U235 (N_235,In_1620,In_1769);
nand U236 (N_236,In_859,In_2334);
nand U237 (N_237,In_2118,In_2313);
nand U238 (N_238,In_2661,In_373);
nor U239 (N_239,In_2649,In_2228);
xor U240 (N_240,In_1861,In_87);
or U241 (N_241,In_2783,In_2232);
or U242 (N_242,In_2540,In_1361);
and U243 (N_243,In_1416,In_698);
nand U244 (N_244,In_1443,In_1631);
or U245 (N_245,In_1044,In_2284);
nor U246 (N_246,In_2878,In_24);
or U247 (N_247,In_502,In_612);
xor U248 (N_248,In_96,In_1987);
or U249 (N_249,In_877,In_2603);
and U250 (N_250,In_1155,In_2734);
xnor U251 (N_251,In_862,In_635);
nor U252 (N_252,In_962,In_1174);
nor U253 (N_253,In_162,In_775);
nor U254 (N_254,In_2947,In_2493);
nand U255 (N_255,In_2974,In_2071);
and U256 (N_256,In_2287,In_2362);
and U257 (N_257,In_1605,In_1901);
xnor U258 (N_258,In_135,In_695);
xor U259 (N_259,In_1755,In_2505);
nand U260 (N_260,In_898,In_1821);
or U261 (N_261,In_2913,In_354);
nor U262 (N_262,In_546,In_761);
or U263 (N_263,In_2961,In_749);
or U264 (N_264,In_1868,In_1599);
xor U265 (N_265,In_1289,In_1336);
nor U266 (N_266,In_1396,In_1841);
nor U267 (N_267,In_1927,In_2236);
and U268 (N_268,In_680,In_1006);
nor U269 (N_269,In_486,In_1480);
xor U270 (N_270,In_2031,In_1139);
nor U271 (N_271,In_340,In_1254);
nor U272 (N_272,In_120,In_2960);
nand U273 (N_273,In_2133,In_134);
and U274 (N_274,In_1041,In_2624);
and U275 (N_275,In_2902,In_1613);
and U276 (N_276,In_1690,In_2618);
and U277 (N_277,In_19,In_2365);
or U278 (N_278,In_2079,In_2441);
nand U279 (N_279,In_1164,In_1181);
nand U280 (N_280,In_2281,In_2939);
xor U281 (N_281,In_2496,In_113);
or U282 (N_282,In_2009,In_1202);
and U283 (N_283,In_552,In_2326);
or U284 (N_284,In_2779,In_2525);
nor U285 (N_285,In_1219,In_64);
nand U286 (N_286,In_2205,In_2951);
nor U287 (N_287,In_258,In_14);
nor U288 (N_288,In_1860,In_283);
nand U289 (N_289,In_1946,In_1902);
or U290 (N_290,In_1710,In_1529);
and U291 (N_291,In_1130,In_700);
xnor U292 (N_292,In_524,In_1998);
or U293 (N_293,In_1192,In_395);
nand U294 (N_294,In_1676,In_2137);
xor U295 (N_295,In_884,In_1183);
and U296 (N_296,In_217,In_2864);
and U297 (N_297,In_70,In_1593);
nand U298 (N_298,In_1887,In_1876);
and U299 (N_299,In_2158,In_1884);
and U300 (N_300,In_61,In_2376);
nand U301 (N_301,In_923,In_2179);
xor U302 (N_302,In_2528,In_670);
nand U303 (N_303,In_2378,In_2065);
nor U304 (N_304,In_1838,In_1339);
nand U305 (N_305,In_693,In_538);
or U306 (N_306,In_207,In_2599);
xor U307 (N_307,In_1530,In_169);
nand U308 (N_308,In_652,In_5);
nand U309 (N_309,In_2681,In_1089);
nand U310 (N_310,In_812,In_1165);
or U311 (N_311,In_769,In_951);
and U312 (N_312,In_2977,In_2209);
nor U313 (N_313,In_1751,In_2351);
nand U314 (N_314,In_1188,In_804);
and U315 (N_315,In_686,In_1309);
xor U316 (N_316,In_1325,In_1794);
nor U317 (N_317,In_1885,In_469);
or U318 (N_318,In_1232,In_2164);
or U319 (N_319,In_2825,In_2360);
xnor U320 (N_320,In_1293,In_2749);
xor U321 (N_321,In_2713,In_2173);
or U322 (N_322,In_2559,In_579);
xnor U323 (N_323,In_2145,In_1261);
nand U324 (N_324,In_1196,In_1879);
nor U325 (N_325,In_79,In_2439);
nor U326 (N_326,In_2562,In_1038);
or U327 (N_327,In_979,In_2958);
and U328 (N_328,In_772,In_708);
nor U329 (N_329,In_944,In_1644);
nor U330 (N_330,In_1251,In_2052);
or U331 (N_331,In_2983,In_459);
xnor U332 (N_332,In_1825,In_2245);
or U333 (N_333,In_2590,In_444);
xnor U334 (N_334,In_830,In_1229);
nor U335 (N_335,In_453,In_890);
nor U336 (N_336,In_35,In_2433);
nor U337 (N_337,In_2516,In_2848);
and U338 (N_338,In_1465,In_982);
nand U339 (N_339,In_520,In_2870);
nand U340 (N_340,In_771,In_1865);
and U341 (N_341,In_1609,In_2944);
nor U342 (N_342,In_2421,In_2517);
or U343 (N_343,In_216,In_66);
and U344 (N_344,In_1535,In_1067);
or U345 (N_345,In_1812,In_505);
and U346 (N_346,In_1942,In_384);
xor U347 (N_347,In_2193,In_1556);
nand U348 (N_348,In_886,In_1126);
nand U349 (N_349,In_2887,In_2303);
xor U350 (N_350,In_1992,In_2694);
nor U351 (N_351,In_2345,In_1786);
nand U352 (N_352,In_1971,In_1918);
xnor U353 (N_353,In_1713,In_651);
nor U354 (N_354,In_2669,In_1551);
nand U355 (N_355,In_466,In_2952);
or U356 (N_356,In_2480,In_2238);
nand U357 (N_357,In_1032,In_582);
nor U358 (N_358,In_1365,In_2483);
xnor U359 (N_359,In_1286,In_254);
and U360 (N_360,In_1421,In_2846);
and U361 (N_361,In_2155,In_1904);
or U362 (N_362,In_2001,In_2537);
nand U363 (N_363,In_2310,In_894);
xor U364 (N_364,In_835,In_1237);
nor U365 (N_365,In_1532,In_2003);
nand U366 (N_366,In_2700,In_858);
or U367 (N_367,In_1101,In_2440);
or U368 (N_368,In_941,In_479);
and U369 (N_369,In_1499,In_1172);
or U370 (N_370,In_2199,In_1082);
and U371 (N_371,In_555,In_2399);
nor U372 (N_372,In_2467,In_2366);
nand U373 (N_373,In_926,In_1201);
nand U374 (N_374,In_2573,In_1080);
nor U375 (N_375,In_292,In_791);
xnor U376 (N_376,In_2391,In_233);
xor U377 (N_377,In_73,In_1117);
nor U378 (N_378,In_1505,In_2554);
xor U379 (N_379,In_2893,In_2668);
and U380 (N_380,In_1266,In_588);
or U381 (N_381,In_255,In_32);
xor U382 (N_382,In_2578,In_2501);
nand U383 (N_383,In_1922,In_1724);
and U384 (N_384,In_2930,In_2642);
nor U385 (N_385,In_1182,In_903);
nand U386 (N_386,In_1388,In_916);
nand U387 (N_387,In_1511,In_86);
xnor U388 (N_388,In_1642,In_1768);
nor U389 (N_389,In_1110,In_1476);
nor U390 (N_390,In_1804,In_2548);
or U391 (N_391,In_676,In_2920);
and U392 (N_392,In_677,In_795);
and U393 (N_393,In_1011,In_1536);
and U394 (N_394,In_2218,In_2220);
nand U395 (N_395,In_535,In_228);
xnor U396 (N_396,In_2545,In_2200);
nor U397 (N_397,In_2805,In_2989);
or U398 (N_398,In_1275,In_2627);
nand U399 (N_399,In_2796,In_1670);
and U400 (N_400,In_2502,In_2147);
or U401 (N_401,In_902,In_240);
xnor U402 (N_402,In_2407,In_1957);
nand U403 (N_403,In_2778,In_2405);
and U404 (N_404,In_2763,In_1141);
xor U405 (N_405,In_1230,In_1146);
and U406 (N_406,In_639,In_1425);
nand U407 (N_407,In_1827,In_338);
nand U408 (N_408,In_601,In_1438);
or U409 (N_409,In_765,In_2686);
and U410 (N_410,In_17,In_1763);
xnor U411 (N_411,In_2591,In_2307);
nand U412 (N_412,In_1952,In_1985);
xnor U413 (N_413,In_964,In_904);
or U414 (N_414,In_324,In_897);
xnor U415 (N_415,In_853,In_475);
nor U416 (N_416,In_1461,In_1279);
or U417 (N_417,In_423,In_2866);
nor U418 (N_418,In_366,In_307);
nand U419 (N_419,In_2432,In_2374);
xor U420 (N_420,In_710,In_658);
nor U421 (N_421,In_985,In_591);
xnor U422 (N_422,In_782,In_1300);
or U423 (N_423,In_1435,In_2940);
and U424 (N_424,In_880,In_2389);
or U425 (N_425,In_2038,In_280);
or U426 (N_426,In_2725,In_2814);
nand U427 (N_427,In_2260,In_2100);
nand U428 (N_428,In_1738,In_1948);
and U429 (N_429,In_2168,In_2132);
nand U430 (N_430,In_1999,In_1882);
nand U431 (N_431,In_1616,In_2077);
or U432 (N_432,In_2884,In_2664);
or U433 (N_433,In_1886,In_561);
nor U434 (N_434,In_418,In_403);
nor U435 (N_435,In_2975,In_1128);
xnor U436 (N_436,In_1488,In_1069);
nor U437 (N_437,In_220,In_1193);
and U438 (N_438,In_2770,In_1574);
nand U439 (N_439,In_437,In_934);
xnor U440 (N_440,In_1152,In_2462);
and U441 (N_441,In_1555,In_249);
or U442 (N_442,In_1355,In_1004);
xor U443 (N_443,In_1533,In_1705);
nand U444 (N_444,In_1651,In_298);
xnor U445 (N_445,In_1298,In_2297);
nor U446 (N_446,In_987,In_1337);
and U447 (N_447,In_1583,In_2596);
xnor U448 (N_448,In_2774,In_2613);
xnor U449 (N_449,In_599,In_1466);
nor U450 (N_450,In_370,In_1921);
xor U451 (N_451,In_1516,In_2942);
nor U452 (N_452,In_2512,In_2737);
or U453 (N_453,In_675,In_1197);
or U454 (N_454,In_615,In_1305);
nor U455 (N_455,In_1222,In_958);
xor U456 (N_456,In_2542,In_537);
nor U457 (N_457,In_2853,In_489);
nand U458 (N_458,In_397,In_150);
xor U459 (N_459,In_1784,In_2475);
and U460 (N_460,In_1626,In_2066);
nor U461 (N_461,In_1813,In_2355);
nand U462 (N_462,In_1220,In_823);
nand U463 (N_463,In_584,In_641);
nand U464 (N_464,In_85,In_2328);
nor U465 (N_465,In_2454,In_1565);
xnor U466 (N_466,In_1398,In_1351);
nor U467 (N_467,In_1689,In_813);
nor U468 (N_468,In_702,In_129);
nand U469 (N_469,In_1837,In_2420);
nand U470 (N_470,In_2300,In_2875);
nor U471 (N_471,In_2575,In_2580);
and U472 (N_472,In_932,In_855);
xnor U473 (N_473,In_574,In_833);
and U474 (N_474,In_2818,In_1598);
nand U475 (N_475,In_2033,In_223);
nand U476 (N_476,In_2043,In_2427);
xnor U477 (N_477,In_440,In_2533);
xnor U478 (N_478,In_337,In_454);
nor U479 (N_479,In_899,In_1716);
nand U480 (N_480,In_1374,In_1276);
or U481 (N_481,In_2682,In_653);
and U482 (N_482,In_965,In_2175);
and U483 (N_483,In_1394,In_1427);
nand U484 (N_484,In_389,In_719);
xor U485 (N_485,In_250,In_2459);
nor U486 (N_486,In_2180,In_256);
xor U487 (N_487,In_966,In_845);
or U488 (N_488,In_2317,In_1216);
and U489 (N_489,In_399,In_2254);
xnor U490 (N_490,In_748,In_2410);
nor U491 (N_491,In_117,In_1845);
xnor U492 (N_492,In_1761,In_2110);
or U493 (N_493,In_2344,In_1013);
and U494 (N_494,In_2198,In_2515);
xnor U495 (N_495,In_1411,In_1071);
nand U496 (N_496,In_2781,In_1650);
xnor U497 (N_497,In_388,In_1334);
nand U498 (N_498,In_1494,In_1687);
xnor U499 (N_499,In_1114,In_45);
nand U500 (N_500,In_2601,In_516);
and U501 (N_501,In_439,In_2593);
xnor U502 (N_502,In_1500,In_2150);
or U503 (N_503,In_182,In_2728);
and U504 (N_504,In_2305,In_334);
nand U505 (N_505,In_1648,In_1531);
and U506 (N_506,In_840,In_1272);
nor U507 (N_507,In_269,In_874);
and U508 (N_508,In_1653,In_785);
or U509 (N_509,In_650,In_206);
nand U510 (N_510,In_410,In_2202);
xor U511 (N_511,In_1718,In_869);
nand U512 (N_512,In_952,In_2388);
or U513 (N_513,In_1415,In_553);
xnor U514 (N_514,In_1818,In_2948);
nand U515 (N_515,In_1075,In_2044);
xnor U516 (N_516,In_1538,In_165);
nand U517 (N_517,In_1608,In_1294);
nand U518 (N_518,In_2247,In_971);
xnor U519 (N_519,In_645,In_329);
and U520 (N_520,In_1315,In_2903);
or U521 (N_521,In_726,In_548);
and U522 (N_522,In_52,In_1677);
or U523 (N_523,In_2629,In_393);
and U524 (N_524,In_419,In_2521);
nor U525 (N_525,In_1955,In_918);
nand U526 (N_526,In_2619,In_209);
or U527 (N_527,In_2561,In_1652);
and U528 (N_528,In_2274,In_168);
or U529 (N_529,In_1669,In_1149);
nor U530 (N_530,In_90,In_272);
nor U531 (N_531,In_2206,In_1814);
or U532 (N_532,In_1163,In_2862);
nand U533 (N_533,In_264,In_2309);
xnor U534 (N_534,In_648,In_2369);
nand U535 (N_535,In_1725,In_1798);
xnor U536 (N_536,In_1731,In_2169);
nand U537 (N_537,In_2191,In_2980);
xor U538 (N_538,In_420,In_1703);
and U539 (N_539,In_2623,In_2847);
or U540 (N_540,In_820,In_308);
or U541 (N_541,In_1472,In_1742);
and U542 (N_542,In_1354,In_602);
or U543 (N_543,In_2861,In_1475);
xnor U544 (N_544,In_2841,In_321);
nand U545 (N_545,In_2017,In_661);
nor U546 (N_546,In_1440,In_768);
nor U547 (N_547,In_1022,In_131);
nor U548 (N_548,In_175,In_76);
nand U549 (N_549,In_1175,In_2858);
or U550 (N_550,In_2073,In_1215);
nor U551 (N_551,In_767,In_2817);
nor U552 (N_552,In_2611,In_1977);
nor U553 (N_553,In_2785,In_1439);
or U554 (N_554,In_1111,In_291);
or U555 (N_555,In_928,In_2472);
and U556 (N_556,In_878,In_1923);
or U557 (N_557,In_1431,In_299);
nor U558 (N_558,In_1288,In_1995);
and U559 (N_559,In_1168,In_2359);
or U560 (N_560,In_600,In_667);
or U561 (N_561,In_2868,In_2928);
and U562 (N_562,In_649,In_2823);
nor U563 (N_563,In_1303,In_1595);
xor U564 (N_564,In_919,In_1692);
or U565 (N_565,In_1980,In_1278);
nor U566 (N_566,In_925,In_668);
and U567 (N_567,In_2556,In_2670);
nand U568 (N_568,In_2258,In_1907);
nand U569 (N_569,In_2182,In_1950);
or U570 (N_570,In_1154,In_1025);
nor U571 (N_571,In_1600,In_498);
and U572 (N_572,In_1125,In_870);
xnor U573 (N_573,In_1741,In_829);
or U574 (N_574,In_1012,In_1135);
and U575 (N_575,In_2832,In_367);
nor U576 (N_576,In_317,In_2911);
xor U577 (N_577,In_1282,In_2471);
nor U578 (N_578,In_1078,In_2264);
nor U579 (N_579,In_689,In_816);
or U580 (N_580,In_2243,In_2789);
or U581 (N_581,In_1989,In_1866);
nand U582 (N_582,In_194,In_1241);
nor U583 (N_583,In_1840,In_446);
or U584 (N_584,In_2759,In_2986);
xnor U585 (N_585,In_672,In_200);
nor U586 (N_586,In_2268,In_2186);
or U587 (N_587,In_414,In_1019);
or U588 (N_588,In_1835,In_2560);
and U589 (N_589,In_1277,In_122);
and U590 (N_590,In_1656,In_522);
xnor U591 (N_591,In_476,In_2705);
nand U592 (N_592,In_1450,In_1495);
and U593 (N_593,In_1781,In_2455);
or U594 (N_594,In_933,In_1377);
and U595 (N_595,In_468,In_1870);
and U596 (N_596,In_1178,In_1385);
and U597 (N_597,In_873,In_549);
nand U598 (N_598,In_2965,In_606);
and U599 (N_599,In_2426,In_2810);
xnor U600 (N_600,In_1789,In_2196);
and U601 (N_601,In_2701,In_986);
nand U602 (N_602,In_2976,In_2849);
or U603 (N_603,In_2970,In_2935);
nor U604 (N_604,In_755,In_501);
nor U605 (N_605,In_2082,In_2857);
or U606 (N_606,In_1515,In_2089);
nor U607 (N_607,In_1233,In_211);
xor U608 (N_608,In_2278,In_1449);
or U609 (N_609,In_970,In_1323);
or U610 (N_610,In_13,In_1520);
nand U611 (N_611,In_2896,In_1217);
or U612 (N_612,In_499,In_1112);
nand U613 (N_613,In_1688,In_2640);
xnor U614 (N_614,In_993,In_2567);
nand U615 (N_615,In_638,In_2385);
xnor U616 (N_616,In_576,In_603);
xnor U617 (N_617,In_2879,In_2616);
and U618 (N_618,In_684,In_568);
nand U619 (N_619,In_2889,In_1509);
nor U620 (N_620,In_879,In_2743);
nand U621 (N_621,In_2165,In_1663);
and U622 (N_622,In_369,In_634);
nand U623 (N_623,In_1143,In_547);
and U624 (N_624,In_2583,In_1335);
and U625 (N_625,In_544,In_43);
or U626 (N_626,In_2134,In_360);
or U627 (N_627,In_770,In_2111);
nand U628 (N_628,In_1579,In_2152);
nor U629 (N_629,In_128,In_1214);
nor U630 (N_630,In_1347,In_1791);
nor U631 (N_631,In_300,In_386);
nor U632 (N_632,In_1119,In_6);
xnor U633 (N_633,In_391,In_776);
or U634 (N_634,In_2724,In_2340);
or U635 (N_635,In_1424,In_1491);
xor U636 (N_636,In_109,In_2123);
nand U637 (N_637,In_2064,In_29);
nand U638 (N_638,In_219,In_2529);
and U639 (N_639,In_318,In_1510);
and U640 (N_640,In_2029,In_1805);
xnor U641 (N_641,In_1161,In_243);
or U642 (N_642,In_428,In_1939);
or U643 (N_643,In_2555,In_2058);
or U644 (N_644,In_1228,In_2711);
or U645 (N_645,In_1470,In_124);
or U646 (N_646,In_47,In_2675);
nor U647 (N_647,In_1782,In_2443);
xnor U648 (N_648,In_2076,In_392);
nor U649 (N_649,In_1212,In_179);
and U650 (N_650,In_915,In_319);
nor U651 (N_651,In_2178,In_1991);
and U652 (N_652,In_2936,In_2306);
and U653 (N_653,In_1968,In_844);
nand U654 (N_654,In_344,In_2122);
xor U655 (N_655,In_1562,In_729);
nand U656 (N_656,In_1906,In_483);
nand U657 (N_657,In_1054,In_891);
or U658 (N_658,In_491,In_151);
nand U659 (N_659,In_1065,In_2535);
and U660 (N_660,In_1730,In_197);
or U661 (N_661,In_2000,In_564);
nand U662 (N_662,In_2354,In_1121);
and U663 (N_663,In_1693,In_1047);
and U664 (N_664,In_2403,In_1607);
or U665 (N_665,In_2534,In_1210);
nor U666 (N_666,In_972,In_1873);
nand U667 (N_667,In_2716,In_1338);
and U668 (N_668,In_1521,In_1133);
xnor U669 (N_669,In_1554,In_2104);
nor U670 (N_670,In_230,In_2479);
nand U671 (N_671,In_750,In_1284);
and U672 (N_672,In_2854,In_2921);
and U673 (N_673,In_1268,In_924);
nor U674 (N_674,In_948,In_1250);
and U675 (N_675,In_1263,In_474);
and U676 (N_676,In_229,In_528);
xor U677 (N_677,In_1073,In_116);
or U678 (N_678,In_1954,In_348);
or U679 (N_679,In_1034,In_2654);
nor U680 (N_680,In_2689,In_560);
nor U681 (N_681,In_810,In_2748);
nand U682 (N_682,In_2793,In_2452);
and U683 (N_683,In_2800,In_472);
and U684 (N_684,In_2900,In_740);
and U685 (N_685,In_239,In_1548);
xor U686 (N_686,In_2576,In_2738);
nor U687 (N_687,In_110,In_1248);
and U688 (N_688,In_1569,In_1085);
nand U689 (N_689,In_2396,In_493);
and U690 (N_690,In_1199,In_2356);
xnor U691 (N_691,In_2653,In_2352);
nand U692 (N_692,In_1667,In_1880);
nand U693 (N_693,In_2585,In_481);
xor U694 (N_694,In_662,In_132);
and U695 (N_695,In_2093,In_2292);
nand U696 (N_696,In_849,In_711);
and U697 (N_697,In_525,In_1544);
xnor U698 (N_698,In_1381,In_969);
and U699 (N_699,In_2815,In_945);
nor U700 (N_700,In_2691,In_892);
nand U701 (N_701,In_534,In_2806);
or U702 (N_702,In_305,In_1709);
nand U703 (N_703,In_1851,In_2754);
and U704 (N_704,In_1859,In_458);
xnor U705 (N_705,In_2235,In_51);
xor U706 (N_706,In_2484,In_2910);
nand U707 (N_707,In_2377,In_2510);
and U708 (N_708,In_2978,In_7);
nand U709 (N_709,In_2409,In_2709);
nand U710 (N_710,In_1862,In_2651);
nor U711 (N_711,In_764,In_2995);
and U712 (N_712,In_1735,In_1058);
nor U713 (N_713,In_436,In_445);
nor U714 (N_714,In_1932,In_15);
nand U715 (N_715,In_2451,In_663);
nand U716 (N_716,In_1373,In_2908);
and U717 (N_717,In_1855,In_1935);
xor U718 (N_718,In_214,In_1321);
nand U719 (N_719,In_893,In_2096);
xor U720 (N_720,In_56,In_805);
nand U721 (N_721,In_1252,In_1743);
or U722 (N_722,In_1370,In_2144);
and U723 (N_723,In_1587,In_1937);
or U724 (N_724,In_212,In_1636);
or U725 (N_725,In_1988,In_1962);
or U726 (N_726,In_1717,In_725);
and U727 (N_727,In_2509,In_1773);
xnor U728 (N_728,In_2101,In_55);
or U729 (N_729,In_1096,In_2370);
xor U730 (N_730,In_2587,In_1206);
xnor U731 (N_731,In_2319,In_2270);
nand U732 (N_732,In_1045,In_1311);
xor U733 (N_733,In_2230,In_1929);
and U734 (N_734,In_2330,In_1668);
xor U735 (N_735,In_374,In_2207);
or U736 (N_736,In_864,In_372);
nor U737 (N_737,In_1850,In_2324);
nand U738 (N_738,In_504,In_2159);
and U739 (N_739,In_2277,In_2897);
nor U740 (N_740,In_1107,In_1043);
nor U741 (N_741,In_1949,In_2712);
and U742 (N_742,In_99,In_1740);
nor U743 (N_743,In_1750,In_2347);
or U744 (N_744,In_716,In_417);
nor U745 (N_745,In_2929,In_482);
nand U746 (N_746,In_2170,In_2163);
nor U747 (N_747,In_811,In_2617);
and U748 (N_748,In_2966,In_968);
nor U749 (N_749,In_464,In_2102);
nor U750 (N_750,In_1115,In_2581);
and U751 (N_751,In_1048,In_145);
or U752 (N_752,In_2916,In_377);
nor U753 (N_753,In_137,In_267);
and U754 (N_754,In_707,In_848);
or U755 (N_755,In_1836,In_2308);
or U756 (N_756,In_1568,In_1448);
and U757 (N_757,In_443,In_1015);
xnor U758 (N_758,In_1382,In_21);
nand U759 (N_759,In_210,In_1618);
and U760 (N_760,In_655,In_57);
or U761 (N_761,In_2149,In_2068);
nor U762 (N_762,In_2671,In_279);
nand U763 (N_763,In_2083,In_1752);
nand U764 (N_764,In_2272,In_2722);
nor U765 (N_765,In_364,In_1745);
and U766 (N_766,In_1350,In_1490);
xor U767 (N_767,In_1584,In_1081);
or U768 (N_768,In_105,In_2660);
nand U769 (N_769,In_2016,In_581);
xnor U770 (N_770,In_37,In_92);
and U771 (N_771,In_2035,In_2885);
xnor U772 (N_772,In_441,In_1072);
and U773 (N_773,In_1299,In_613);
and U774 (N_774,In_357,In_2600);
or U775 (N_775,In_1308,In_1384);
xor U776 (N_776,In_327,In_107);
and U777 (N_777,In_201,In_2532);
and U778 (N_778,In_1697,In_1539);
and U779 (N_779,In_939,In_1098);
nor U780 (N_780,In_2237,In_815);
nand U781 (N_781,In_2316,In_2447);
and U782 (N_782,In_378,In_1635);
or U783 (N_783,In_621,In_2212);
and U784 (N_784,In_1578,In_2167);
or U785 (N_785,In_2106,In_2608);
or U786 (N_786,In_148,In_2639);
nand U787 (N_787,In_2350,In_510);
xor U788 (N_788,In_260,In_2074);
nand U789 (N_789,In_694,In_2037);
nand U790 (N_790,In_988,In_1943);
or U791 (N_791,In_276,In_567);
or U792 (N_792,In_287,In_1318);
nand U793 (N_793,In_1008,In_1393);
and U794 (N_794,In_2322,In_1319);
or U795 (N_795,In_511,In_1809);
nor U796 (N_796,In_647,In_1247);
xnor U797 (N_797,In_790,In_872);
or U798 (N_798,In_2157,In_2337);
xnor U799 (N_799,In_2262,In_796);
and U800 (N_800,In_1242,In_1046);
nand U801 (N_801,In_2598,In_1302);
or U802 (N_802,In_257,In_673);
nand U803 (N_803,In_1793,In_743);
xnor U804 (N_804,In_850,In_2799);
and U805 (N_805,In_2495,In_2054);
nor U806 (N_806,In_955,In_2105);
nor U807 (N_807,In_656,In_248);
xnor U808 (N_808,In_1507,In_199);
nand U809 (N_809,In_1453,In_138);
or U810 (N_810,In_2219,In_106);
and U811 (N_811,In_1559,In_736);
nor U812 (N_812,In_2531,In_2543);
or U813 (N_813,In_1074,In_242);
and U814 (N_814,In_2967,In_1503);
xnor U815 (N_815,In_1479,In_461);
nor U816 (N_816,In_587,In_1285);
nor U817 (N_817,In_1208,In_315);
xnor U818 (N_818,In_2392,In_2782);
xor U819 (N_819,In_1244,In_259);
xor U820 (N_820,In_123,In_1982);
xor U821 (N_821,In_630,In_1187);
nor U822 (N_822,In_2450,In_1964);
and U823 (N_823,In_752,In_139);
xor U824 (N_824,In_394,In_1024);
nand U825 (N_825,In_666,In_1348);
nand U826 (N_826,In_2626,In_2811);
xor U827 (N_827,In_1136,In_2004);
nand U828 (N_828,In_721,In_2520);
nor U829 (N_829,In_2609,In_1005);
nor U830 (N_830,In_196,In_960);
and U831 (N_831,In_115,In_1872);
nor U832 (N_832,In_2886,In_626);
xor U833 (N_833,In_18,In_690);
nand U834 (N_834,In_604,In_2892);
xor U835 (N_835,In_470,In_487);
and U836 (N_836,In_1654,In_69);
nor U837 (N_837,In_1758,In_121);
or U838 (N_838,In_2006,In_2325);
nor U839 (N_839,In_1469,In_1623);
xor U840 (N_840,In_1673,In_2760);
or U841 (N_841,In_157,In_188);
and U842 (N_842,In_492,In_857);
and U843 (N_843,In_1169,In_2698);
nand U844 (N_844,In_262,In_1760);
or U845 (N_845,In_2063,In_927);
and U846 (N_846,In_2750,In_1604);
nand U847 (N_847,In_36,In_251);
nand U848 (N_848,In_806,In_114);
or U849 (N_849,In_1698,In_8);
or U850 (N_850,In_947,In_834);
nand U851 (N_851,In_2788,In_1737);
xor U852 (N_852,In_1571,In_2898);
xor U853 (N_853,In_2380,In_2011);
and U854 (N_854,In_2092,In_2302);
nor U855 (N_855,In_2057,In_16);
and U856 (N_856,In_1958,In_1062);
or U857 (N_857,In_1342,In_950);
nor U858 (N_858,In_1547,In_2852);
or U859 (N_859,In_1097,In_331);
nand U860 (N_860,In_2645,In_289);
nor U861 (N_861,In_2855,In_2506);
or U862 (N_862,In_2304,In_1264);
nand U863 (N_863,In_1184,In_2039);
or U864 (N_864,In_2997,In_917);
or U865 (N_865,In_713,In_234);
and U866 (N_866,In_2449,In_1736);
xnor U867 (N_867,In_2112,In_376);
nand U868 (N_868,In_2197,In_2276);
and U869 (N_869,In_11,In_2835);
nor U870 (N_870,In_2845,In_1983);
nor U871 (N_871,In_1903,In_2222);
xor U872 (N_872,In_1159,In_2418);
nand U873 (N_873,In_2294,In_2829);
nor U874 (N_874,In_1874,In_2474);
nand U875 (N_875,In_2883,In_1483);
xnor U876 (N_876,In_398,In_341);
xor U877 (N_877,In_202,In_1843);
and U878 (N_878,In_2739,In_1993);
nand U879 (N_879,In_1944,In_2614);
or U880 (N_880,In_2138,In_1589);
or U881 (N_881,In_314,In_95);
and U882 (N_882,In_1145,In_39);
nand U883 (N_883,In_2953,In_2839);
or U884 (N_884,In_2253,In_2339);
nand U885 (N_885,In_2061,In_2408);
and U886 (N_886,In_2673,In_2266);
and U887 (N_887,In_1796,In_976);
nor U888 (N_888,In_1227,In_2588);
xor U889 (N_889,In_1372,In_1645);
xor U890 (N_890,In_2171,In_413);
xor U891 (N_891,In_2558,In_1007);
and U892 (N_892,In_2402,In_2704);
and U893 (N_893,In_2915,In_607);
and U894 (N_894,In_2419,In_1996);
nand U895 (N_895,In_2676,In_1889);
or U896 (N_896,In_189,In_1540);
or U897 (N_897,In_404,In_714);
xor U898 (N_898,In_2524,In_383);
nor U899 (N_899,In_786,In_447);
or U900 (N_900,In_400,In_1675);
and U901 (N_901,In_2513,In_2630);
xnor U902 (N_902,In_1200,In_1091);
or U903 (N_903,In_792,In_732);
nand U904 (N_904,In_777,In_2139);
nor U905 (N_905,In_2466,In_2917);
or U906 (N_906,In_2435,In_1077);
or U907 (N_907,In_1413,In_2901);
nand U908 (N_908,In_149,In_2423);
and U909 (N_909,In_2955,In_2621);
xor U910 (N_910,In_477,In_422);
and U911 (N_911,In_2569,In_2756);
xnor U912 (N_912,In_22,In_2919);
xor U913 (N_913,In_1340,In_2395);
and U914 (N_914,In_808,In_836);
nand U915 (N_915,In_186,In_1028);
and U916 (N_916,In_994,In_237);
nor U917 (N_917,In_865,In_427);
or U918 (N_918,In_1273,In_1103);
nor U919 (N_919,In_2241,In_343);
or U920 (N_920,In_851,In_1147);
xor U921 (N_921,In_1728,In_65);
xnor U922 (N_922,In_253,In_1523);
and U923 (N_923,In_2615,In_1723);
nand U924 (N_924,In_1881,In_1364);
nand U925 (N_925,In_2644,In_514);
or U926 (N_926,In_2259,In_235);
nor U927 (N_927,In_1867,In_27);
or U928 (N_928,In_1757,In_2314);
or U929 (N_929,In_342,In_533);
xnor U930 (N_930,In_1405,In_741);
nand U931 (N_931,In_2379,In_2720);
nand U932 (N_932,In_1580,In_2971);
and U933 (N_933,In_2876,In_345);
or U934 (N_934,In_1722,In_2491);
xor U935 (N_935,In_611,In_2566);
nand U936 (N_936,In_571,In_2358);
xor U937 (N_937,In_1951,In_2458);
and U938 (N_938,In_1446,In_605);
xor U939 (N_939,In_252,In_2522);
or U940 (N_940,In_1331,In_1326);
nand U941 (N_941,In_1269,In_97);
xnor U942 (N_942,In_1243,In_2795);
and U943 (N_943,In_2424,In_2867);
and U944 (N_944,In_1576,In_2081);
and U945 (N_945,In_1912,In_671);
or U946 (N_946,In_181,In_2776);
nand U947 (N_947,In_1225,In_598);
and U948 (N_948,In_854,In_2672);
and U949 (N_949,In_2286,In_1646);
nor U950 (N_950,In_759,In_819);
or U951 (N_951,In_185,In_9);
nor U952 (N_952,In_1171,In_678);
and U953 (N_953,In_2195,In_1662);
or U954 (N_954,In_1026,In_198);
xnor U955 (N_955,In_270,In_1801);
xor U956 (N_956,In_1700,In_274);
xor U957 (N_957,In_2130,In_1660);
or U958 (N_958,In_1517,In_1255);
and U959 (N_959,In_84,In_783);
xnor U960 (N_960,In_2227,In_213);
and U961 (N_961,In_1661,In_632);
or U962 (N_962,In_100,In_433);
or U963 (N_963,In_2771,In_636);
xor U964 (N_964,In_1671,In_706);
nand U965 (N_965,In_2014,In_563);
xor U966 (N_966,In_589,In_2747);
nor U967 (N_967,In_322,In_146);
xor U968 (N_968,In_681,In_295);
xor U969 (N_969,In_1581,In_1327);
or U970 (N_970,In_2456,In_91);
xnor U971 (N_971,In_1888,In_802);
nand U972 (N_972,In_2348,In_1395);
xnor U973 (N_973,In_184,In_2934);
xnor U974 (N_974,In_1407,In_225);
and U975 (N_975,In_2757,In_1186);
nor U976 (N_976,In_1258,In_1419);
and U977 (N_977,In_1166,In_622);
nor U978 (N_978,In_953,In_1940);
or U979 (N_979,In_2153,In_1916);
nor U980 (N_980,In_40,In_2135);
and U981 (N_981,In_779,In_1316);
nand U982 (N_982,In_995,In_1680);
and U983 (N_983,In_1281,In_2045);
nor U984 (N_984,In_1454,In_226);
xor U985 (N_985,In_2025,In_12);
xnor U986 (N_986,In_1970,In_2633);
nor U987 (N_987,In_2787,In_687);
or U988 (N_988,In_2803,In_167);
nand U989 (N_989,In_2945,In_1513);
and U990 (N_990,In_2744,In_1732);
nor U991 (N_991,In_2249,In_1138);
xor U992 (N_992,In_2765,In_1749);
nand U993 (N_993,In_2761,In_1056);
xnor U994 (N_994,In_935,In_1423);
or U995 (N_995,In_2772,In_2932);
or U996 (N_996,In_620,In_2703);
nor U997 (N_997,In_2210,In_1189);
nor U998 (N_998,In_136,In_177);
nor U999 (N_999,In_2250,In_657);
or U1000 (N_1000,In_1060,In_1833);
and U1001 (N_1001,In_712,In_2820);
and U1002 (N_1002,In_1848,In_2056);
nor U1003 (N_1003,In_654,In_1053);
and U1004 (N_1004,In_2086,In_2840);
and U1005 (N_1005,In_1442,In_2719);
and U1006 (N_1006,In_288,In_385);
xnor U1007 (N_1007,In_1090,In_71);
and U1008 (N_1008,In_946,In_887);
or U1009 (N_1009,In_2767,In_1467);
xor U1010 (N_1010,In_2926,In_1753);
nand U1011 (N_1011,In_2019,In_2257);
or U1012 (N_1012,In_2084,In_2994);
nand U1013 (N_1013,In_1560,In_1630);
nand U1014 (N_1014,In_2662,In_1010);
and U1015 (N_1015,In_2413,In_2162);
xor U1016 (N_1016,In_2688,In_1894);
xnor U1017 (N_1017,In_2650,In_2023);
xnor U1018 (N_1018,In_2468,In_371);
nand U1019 (N_1019,In_1023,In_1223);
or U1020 (N_1020,In_2126,In_2487);
and U1021 (N_1021,In_2444,In_2546);
nand U1022 (N_1022,In_1037,In_512);
nand U1023 (N_1023,In_1961,In_963);
xor U1024 (N_1024,In_2072,In_328);
nor U1025 (N_1025,In_41,In_2461);
nand U1026 (N_1026,In_1050,In_788);
xnor U1027 (N_1027,In_1379,In_2809);
and U1028 (N_1028,In_2740,In_2741);
nor U1029 (N_1029,In_745,In_625);
and U1030 (N_1030,In_1933,In_1205);
and U1031 (N_1031,In_2172,In_1625);
nand U1032 (N_1032,In_1068,In_153);
nand U1033 (N_1033,In_2658,In_1221);
nand U1034 (N_1034,In_335,In_701);
or U1035 (N_1035,In_784,In_2323);
xnor U1036 (N_1036,In_2234,In_2683);
and U1037 (N_1037,In_1706,In_1930);
xnor U1038 (N_1038,In_1088,In_2336);
nand U1039 (N_1039,In_2188,In_682);
nor U1040 (N_1040,In_1444,In_728);
xor U1041 (N_1041,In_807,In_778);
nor U1042 (N_1042,In_959,In_2564);
xnor U1043 (N_1043,In_244,In_330);
nor U1044 (N_1044,In_457,In_1501);
nor U1045 (N_1045,In_2592,In_1209);
and U1046 (N_1046,In_2129,In_2216);
or U1047 (N_1047,In_2381,In_75);
and U1048 (N_1048,In_2956,In_2457);
nand U1049 (N_1049,In_130,In_1666);
xnor U1050 (N_1050,In_2085,In_2221);
nand U1051 (N_1051,In_794,In_1508);
xnor U1052 (N_1052,In_2684,In_2504);
nor U1053 (N_1053,In_1606,In_1966);
xor U1054 (N_1054,In_1619,In_2692);
xor U1055 (N_1055,In_2190,In_2060);
nor U1056 (N_1056,In_756,In_101);
nand U1057 (N_1057,In_2094,In_1621);
nor U1058 (N_1058,In_1346,In_1224);
and U1059 (N_1059,In_1176,In_519);
and U1060 (N_1060,In_888,In_1854);
nor U1061 (N_1061,In_1376,In_990);
xnor U1062 (N_1062,In_1553,In_2002);
or U1063 (N_1063,In_1485,In_1960);
nand U1064 (N_1064,In_2460,In_1647);
xnor U1065 (N_1065,In_2830,In_346);
and U1066 (N_1066,In_2406,In_977);
and U1067 (N_1067,In_152,In_2985);
xnor U1068 (N_1068,In_2819,In_2766);
xnor U1069 (N_1069,In_2288,In_1712);
xnor U1070 (N_1070,In_1314,In_2114);
xnor U1071 (N_1071,In_1819,In_1857);
nor U1072 (N_1072,In_2448,In_401);
and U1073 (N_1073,In_2291,In_1506);
and U1074 (N_1074,In_1679,In_984);
and U1075 (N_1075,In_25,In_218);
nor U1076 (N_1076,In_1301,In_2477);
xnor U1077 (N_1077,In_2685,In_166);
nor U1078 (N_1078,In_408,In_1390);
xnor U1079 (N_1079,In_1392,In_2393);
nand U1080 (N_1080,In_751,In_59);
or U1081 (N_1081,In_2526,In_911);
or U1082 (N_1082,In_2625,In_1913);
or U1083 (N_1083,In_1524,In_2891);
xor U1084 (N_1084,In_174,In_1541);
nor U1085 (N_1085,In_679,In_2998);
and U1086 (N_1086,In_2880,In_2996);
nor U1087 (N_1087,In_455,In_975);
nand U1088 (N_1088,In_297,In_1994);
nor U1089 (N_1089,In_1526,In_2769);
and U1090 (N_1090,In_1492,In_1823);
nor U1091 (N_1091,In_696,In_1064);
nand U1092 (N_1092,In_1905,In_2372);
or U1093 (N_1093,In_1322,In_1897);
and U1094 (N_1094,In_350,In_1792);
or U1095 (N_1095,In_2256,In_80);
or U1096 (N_1096,In_396,In_1828);
nand U1097 (N_1097,In_578,In_2208);
and U1098 (N_1098,In_2181,In_2311);
and U1099 (N_1099,In_973,In_1853);
xnor U1100 (N_1100,In_2194,In_2333);
and U1101 (N_1101,In_1803,In_1956);
and U1102 (N_1102,In_1777,In_542);
or U1103 (N_1103,In_359,In_1632);
nand U1104 (N_1104,In_375,In_1979);
xnor U1105 (N_1105,In_1917,In_2028);
or U1106 (N_1106,In_2280,In_727);
xor U1107 (N_1107,In_2873,In_2775);
or U1108 (N_1108,In_1990,In_831);
nand U1109 (N_1109,In_1148,In_2024);
nor U1110 (N_1110,In_2177,In_431);
and U1111 (N_1111,In_1259,In_2224);
xnor U1112 (N_1112,In_1249,In_313);
xor U1113 (N_1113,In_2315,In_421);
xnor U1114 (N_1114,In_1597,In_1447);
nand U1115 (N_1115,In_2523,In_739);
and U1116 (N_1116,In_1561,In_2687);
and U1117 (N_1117,In_1358,In_1577);
and U1118 (N_1118,In_2586,In_1296);
nor U1119 (N_1119,In_1203,In_284);
or U1120 (N_1120,In_1707,In_1157);
xor U1121 (N_1121,In_2612,In_358);
and U1122 (N_1122,In_1714,In_798);
nand U1123 (N_1123,In_1785,In_2261);
or U1124 (N_1124,In_1156,In_558);
nor U1125 (N_1125,In_1352,In_1292);
and U1126 (N_1126,In_320,In_500);
and U1127 (N_1127,In_881,In_2828);
and U1128 (N_1128,In_1100,In_992);
nor U1129 (N_1129,In_309,In_1775);
and U1130 (N_1130,In_415,In_2282);
nand U1131 (N_1131,In_1118,In_1087);
nor U1132 (N_1132,In_2470,In_2384);
or U1133 (N_1133,In_31,In_193);
xor U1134 (N_1134,In_780,In_1925);
xnor U1135 (N_1135,In_2463,In_2015);
nand U1136 (N_1136,In_1375,In_2036);
and U1137 (N_1137,In_1806,In_715);
xnor U1138 (N_1138,In_311,In_1312);
and U1139 (N_1139,In_1592,In_841);
or U1140 (N_1140,In_1633,In_2012);
nand U1141 (N_1141,In_1622,In_1017);
and U1142 (N_1142,In_2473,In_1496);
or U1143 (N_1143,In_2710,In_102);
xnor U1144 (N_1144,In_1367,In_2999);
nand U1145 (N_1145,In_1084,In_1387);
xor U1146 (N_1146,In_2856,In_23);
nor U1147 (N_1147,In_1549,In_2373);
nand U1148 (N_1148,In_1628,In_1129);
or U1149 (N_1149,In_967,In_827);
xnor U1150 (N_1150,In_2293,In_1104);
nor U1151 (N_1151,In_1900,In_2154);
xnor U1152 (N_1152,In_961,In_1099);
nor U1153 (N_1153,In_532,In_1612);
nor U1154 (N_1154,In_1113,In_2665);
xor U1155 (N_1155,In_699,In_1403);
nor U1156 (N_1156,In_1856,In_241);
or U1157 (N_1157,In_2053,In_1459);
and U1158 (N_1158,In_843,In_1369);
or U1159 (N_1159,In_1764,In_2755);
and U1160 (N_1160,In_290,In_190);
and U1161 (N_1161,In_2922,In_1877);
or U1162 (N_1162,In_1733,In_485);
nor U1163 (N_1163,In_2912,In_669);
nand U1164 (N_1164,In_2622,In_1457);
xor U1165 (N_1165,In_2931,In_2246);
nand U1166 (N_1166,In_1345,In_922);
nor U1167 (N_1167,In_1537,In_349);
nor U1168 (N_1168,In_2013,In_1386);
nand U1169 (N_1169,In_1428,In_1304);
and U1170 (N_1170,In_2833,In_1482);
xor U1171 (N_1171,In_303,In_709);
nor U1172 (N_1172,In_754,In_839);
xnor U1173 (N_1173,In_1852,In_2751);
and U1174 (N_1174,In_991,In_1659);
nand U1175 (N_1175,In_2099,In_2485);
nor U1176 (N_1176,In_78,In_541);
xor U1177 (N_1177,In_2252,In_1973);
or U1178 (N_1178,In_1066,In_1366);
xnor U1179 (N_1179,In_900,In_2962);
and U1180 (N_1180,In_2223,In_1095);
and U1181 (N_1181,In_1191,In_382);
and U1182 (N_1182,In_365,In_2335);
xor U1183 (N_1183,In_118,In_2918);
xor U1184 (N_1184,In_103,In_281);
xnor U1185 (N_1185,In_517,In_2551);
nor U1186 (N_1186,In_2203,In_515);
nand U1187 (N_1187,In_2990,In_1564);
nand U1188 (N_1188,In_2874,In_930);
and U1189 (N_1189,In_2519,In_2834);
nor U1190 (N_1190,In_2871,In_2632);
nand U1191 (N_1191,In_1083,In_1324);
xnor U1192 (N_1192,In_664,In_821);
or U1193 (N_1193,In_1573,In_2696);
nor U1194 (N_1194,In_509,In_1545);
or U1195 (N_1195,In_1150,In_2753);
nand U1196 (N_1196,In_527,In_1926);
xor U1197 (N_1197,In_172,In_215);
nor U1198 (N_1198,In_1109,In_2733);
or U1199 (N_1199,In_20,In_1518);
and U1200 (N_1200,N_204,N_924);
or U1201 (N_1201,N_1151,N_488);
and U1202 (N_1202,In_286,N_1041);
nor U1203 (N_1203,N_405,In_1040);
xor U1204 (N_1204,N_148,N_942);
or U1205 (N_1205,In_1486,In_2656);
xnor U1206 (N_1206,N_1129,N_401);
or U1207 (N_1207,N_963,In_610);
nor U1208 (N_1208,N_939,N_1140);
nand U1209 (N_1209,In_2166,N_851);
nor U1210 (N_1210,N_1037,In_2434);
or U1211 (N_1211,In_133,N_123);
or U1212 (N_1212,N_409,In_2383);
or U1213 (N_1213,N_139,In_2909);
xnor U1214 (N_1214,N_660,In_2429);
nor U1215 (N_1215,N_663,In_1137);
nand U1216 (N_1216,N_549,N_526);
nand U1217 (N_1217,N_1146,N_99);
nand U1218 (N_1218,N_674,N_837);
or U1219 (N_1219,N_442,N_1088);
xnor U1220 (N_1220,N_840,In_2486);
and U1221 (N_1221,N_66,In_1715);
nor U1222 (N_1222,N_772,In_170);
xor U1223 (N_1223,N_1178,N_1032);
nand U1224 (N_1224,N_627,N_949);
xnor U1225 (N_1225,N_625,N_359);
or U1226 (N_1226,N_358,N_1170);
and U1227 (N_1227,N_1158,N_867);
xnor U1228 (N_1228,N_361,In_1094);
nand U1229 (N_1229,N_749,N_191);
and U1230 (N_1230,In_575,N_599);
xnor U1231 (N_1231,N_936,N_1034);
nor U1232 (N_1232,N_1007,N_441);
and U1233 (N_1233,In_46,N_845);
and U1234 (N_1234,N_803,In_336);
or U1235 (N_1235,N_1031,N_452);
nand U1236 (N_1236,N_1061,In_1919);
nor U1237 (N_1237,In_908,In_720);
or U1238 (N_1238,In_1185,N_703);
and U1239 (N_1239,N_246,N_1114);
xor U1240 (N_1240,N_834,N_450);
or U1241 (N_1241,N_883,N_1120);
and U1242 (N_1242,N_31,In_2140);
xor U1243 (N_1243,In_847,In_465);
or U1244 (N_1244,N_614,In_2010);
nand U1245 (N_1245,N_1195,In_2541);
xor U1246 (N_1246,N_186,N_486);
and U1247 (N_1247,N_317,N_708);
nand U1248 (N_1248,N_220,In_895);
nand U1249 (N_1249,N_241,In_2481);
or U1250 (N_1250,In_1787,N_1123);
nor U1251 (N_1251,N_1119,N_21);
nand U1252 (N_1252,In_595,N_997);
or U1253 (N_1253,N_1164,N_189);
or U1254 (N_1254,N_820,N_567);
or U1255 (N_1255,N_1067,In_2273);
xnor U1256 (N_1256,N_106,N_465);
and U1257 (N_1257,N_208,N_298);
xor U1258 (N_1258,N_278,N_713);
or U1259 (N_1259,N_748,In_2824);
or U1260 (N_1260,N_305,N_383);
and U1261 (N_1261,In_355,N_906);
nand U1262 (N_1262,N_438,N_47);
or U1263 (N_1263,N_583,In_2804);
or U1264 (N_1264,N_711,In_1306);
or U1265 (N_1265,N_929,N_798);
xor U1266 (N_1266,In_183,N_373);
nand U1267 (N_1267,In_793,N_770);
nor U1268 (N_1268,N_454,N_1045);
or U1269 (N_1269,In_205,N_1000);
nor U1270 (N_1270,In_356,N_291);
xor U1271 (N_1271,In_1213,In_1122);
nor U1272 (N_1272,In_26,In_2597);
xor U1273 (N_1273,N_982,N_652);
xor U1274 (N_1274,N_257,In_2269);
nor U1275 (N_1275,N_805,N_194);
nor U1276 (N_1276,N_641,In_2051);
nand U1277 (N_1277,N_722,N_1128);
or U1278 (N_1278,N_113,N_118);
nor U1279 (N_1279,N_1106,N_1005);
or U1280 (N_1280,N_376,N_558);
nor U1281 (N_1281,In_2442,In_2859);
nand U1282 (N_1282,N_607,N_744);
nand U1283 (N_1283,N_615,N_456);
xor U1284 (N_1284,N_1153,N_385);
or U1285 (N_1285,N_461,In_2963);
nand U1286 (N_1286,N_6,In_949);
or U1287 (N_1287,N_1132,In_191);
xor U1288 (N_1288,N_679,N_789);
nor U1289 (N_1289,In_2574,N_1144);
nor U1290 (N_1290,N_13,In_2127);
nand U1291 (N_1291,N_969,N_993);
xnor U1292 (N_1292,N_1115,In_818);
nor U1293 (N_1293,N_143,N_90);
nand U1294 (N_1294,N_530,In_838);
and U1295 (N_1295,N_80,N_691);
xor U1296 (N_1296,N_433,In_2201);
nor U1297 (N_1297,N_842,N_408);
nand U1298 (N_1298,N_374,N_1161);
or U1299 (N_1299,N_823,N_362);
nor U1300 (N_1300,In_703,In_1893);
nand U1301 (N_1301,N_219,N_480);
or U1302 (N_1302,In_1550,N_76);
or U1303 (N_1303,N_0,In_467);
xnor U1304 (N_1304,N_349,N_224);
and U1305 (N_1305,N_616,N_619);
and U1306 (N_1306,In_368,N_554);
and U1307 (N_1307,N_288,N_1121);
nand U1308 (N_1308,N_64,N_618);
nand U1309 (N_1309,In_937,N_821);
and U1310 (N_1310,In_435,N_1087);
nand U1311 (N_1311,N_782,In_646);
nand U1312 (N_1312,N_161,N_345);
xor U1313 (N_1313,N_1077,In_1649);
nand U1314 (N_1314,In_593,N_109);
and U1315 (N_1315,In_1772,N_1069);
nor U1316 (N_1316,N_854,N_910);
nand U1317 (N_1317,N_459,In_1963);
xnor U1318 (N_1318,In_2342,N_1042);
nand U1319 (N_1319,In_478,N_743);
and U1320 (N_1320,N_9,In_2251);
or U1321 (N_1321,N_495,N_694);
and U1322 (N_1322,N_552,In_1947);
and U1323 (N_1323,N_318,N_395);
and U1324 (N_1324,N_17,N_977);
and U1325 (N_1325,In_1739,In_1527);
and U1326 (N_1326,N_518,N_233);
nand U1327 (N_1327,In_1945,N_878);
nand U1328 (N_1328,In_1776,In_2115);
and U1329 (N_1329,In_323,N_42);
nor U1330 (N_1330,N_296,In_1890);
and U1331 (N_1331,N_212,N_890);
and U1332 (N_1332,N_135,In_2394);
xnor U1333 (N_1333,In_921,In_2589);
xnor U1334 (N_1334,In_1695,N_275);
nand U1335 (N_1335,In_2544,N_387);
or U1336 (N_1336,In_1892,N_792);
xnor U1337 (N_1337,N_697,N_1191);
or U1338 (N_1338,N_600,In_2702);
nand U1339 (N_1339,In_2387,N_1075);
nor U1340 (N_1340,In_1102,N_768);
or U1341 (N_1341,N_578,N_508);
nand U1342 (N_1342,N_1029,N_440);
and U1343 (N_1343,N_1073,N_150);
xnor U1344 (N_1344,In_2647,N_574);
nor U1345 (N_1345,In_2500,N_861);
nand U1346 (N_1346,N_1184,N_1142);
nand U1347 (N_1347,N_1112,N_751);
nor U1348 (N_1348,N_863,N_584);
nand U1349 (N_1349,N_263,N_170);
nand U1350 (N_1350,N_357,N_755);
and U1351 (N_1351,N_728,N_475);
nand U1352 (N_1352,N_737,N_669);
nand U1353 (N_1353,In_2735,N_481);
and U1354 (N_1354,N_166,In_2285);
nand U1355 (N_1355,In_1432,In_1055);
or U1356 (N_1356,N_402,N_315);
nor U1357 (N_1357,In_1601,N_24);
or U1358 (N_1358,In_2808,In_2214);
xnor U1359 (N_1359,N_1072,In_1976);
nand U1360 (N_1360,N_1166,N_683);
and U1361 (N_1361,In_82,N_717);
or U1362 (N_1362,N_432,In_1380);
nor U1363 (N_1363,N_689,N_1199);
and U1364 (N_1364,N_302,N_1193);
or U1365 (N_1365,N_44,N_532);
xnor U1366 (N_1366,N_1185,In_692);
xor U1367 (N_1367,N_211,N_436);
nand U1368 (N_1368,N_828,N_1063);
nor U1369 (N_1369,N_180,In_1720);
xor U1370 (N_1370,N_85,N_569);
nor U1371 (N_1371,N_328,N_1126);
and U1372 (N_1372,In_2530,In_2174);
nand U1373 (N_1373,N_739,In_2290);
or U1374 (N_1374,N_1091,N_134);
xor U1375 (N_1375,N_912,In_2020);
xnor U1376 (N_1376,In_1586,In_817);
and U1377 (N_1377,In_2067,N_868);
or U1378 (N_1378,N_494,In_1473);
and U1379 (N_1379,N_427,N_188);
nor U1380 (N_1380,N_754,N_1188);
and U1381 (N_1381,N_701,In_1173);
nor U1382 (N_1382,N_827,N_681);
nor U1383 (N_1383,N_671,In_2142);
nand U1384 (N_1384,In_2636,In_824);
nand U1385 (N_1385,N_88,N_187);
nand U1386 (N_1386,In_1936,N_294);
and U1387 (N_1387,N_629,N_172);
and U1388 (N_1388,In_2987,N_477);
or U1389 (N_1389,N_152,N_921);
or U1390 (N_1390,In_1092,N_418);
and U1391 (N_1391,N_709,In_2279);
nor U1392 (N_1392,N_223,In_665);
or U1393 (N_1393,N_225,N_1025);
and U1394 (N_1394,In_2233,N_1049);
xor U1395 (N_1395,N_237,In_1400);
nor U1396 (N_1396,In_1497,In_1153);
nor U1397 (N_1397,In_407,In_592);
or U1398 (N_1398,N_253,N_455);
nand U1399 (N_1399,In_1585,In_882);
nor U1400 (N_1400,N_561,N_158);
or U1401 (N_1401,In_429,In_1826);
nand U1402 (N_1402,In_619,N_230);
nor U1403 (N_1403,In_1402,In_2863);
or U1404 (N_1404,In_2047,N_1141);
or U1405 (N_1405,N_425,N_699);
xor U1406 (N_1406,In_2415,In_2411);
or U1407 (N_1407,In_1455,N_1165);
and U1408 (N_1408,In_1180,N_758);
nor U1409 (N_1409,N_876,N_661);
and U1410 (N_1410,In_1039,In_1726);
xor U1411 (N_1411,N_1081,N_1033);
nor U1412 (N_1412,In_2489,In_1477);
xnor U1413 (N_1413,In_285,N_375);
or U1414 (N_1414,In_1871,N_1113);
and U1415 (N_1415,N_412,In_1658);
or U1416 (N_1416,N_655,N_724);
xnor U1417 (N_1417,In_2768,In_2690);
and U1418 (N_1418,N_133,In_1711);
or U1419 (N_1419,In_822,N_882);
and U1420 (N_1420,N_1076,N_18);
or U1421 (N_1421,N_502,N_326);
and U1422 (N_1422,N_280,In_381);
nor U1423 (N_1423,N_115,N_103);
xnor U1424 (N_1424,N_593,N_37);
or U1425 (N_1425,N_704,In_1463);
and U1426 (N_1426,In_222,In_1001);
nand U1427 (N_1427,In_2097,In_1235);
nor U1428 (N_1428,N_543,N_469);
nor U1429 (N_1429,N_147,N_382);
xnor U1430 (N_1430,N_444,N_467);
and U1431 (N_1431,In_451,N_946);
and U1432 (N_1432,In_1696,N_637);
xor U1433 (N_1433,N_830,N_1194);
and U1434 (N_1434,In_2984,N_531);
nor U1435 (N_1435,N_544,In_596);
xor U1436 (N_1436,N_283,N_331);
nor U1437 (N_1437,N_706,N_227);
xnor U1438 (N_1438,N_389,N_1026);
nand U1439 (N_1439,N_873,In_943);
and U1440 (N_1440,N_510,N_52);
or U1441 (N_1441,N_853,N_1163);
nor U1442 (N_1442,In_1422,N_1101);
and U1443 (N_1443,N_363,N_206);
nand U1444 (N_1444,N_865,In_2553);
nor U1445 (N_1445,In_797,N_864);
xor U1446 (N_1446,N_261,In_247);
nor U1447 (N_1447,N_991,N_260);
xnor U1448 (N_1448,N_267,In_2732);
xor U1449 (N_1449,In_2907,In_1378);
nor U1450 (N_1450,In_1832,N_644);
nand U1451 (N_1451,N_996,N_301);
nor U1452 (N_1452,N_299,N_285);
nor U1453 (N_1453,N_466,N_738);
nand U1454 (N_1454,N_82,In_2069);
or U1455 (N_1455,In_674,N_682);
nor U1456 (N_1456,N_423,In_837);
nand U1457 (N_1457,In_1445,In_1972);
nor U1458 (N_1458,N_891,N_372);
or U1459 (N_1459,N_229,N_1186);
xor U1460 (N_1460,In_2299,N_50);
xnor U1461 (N_1461,In_1552,N_862);
or U1462 (N_1462,In_1815,N_948);
or U1463 (N_1463,N_396,N_84);
xor U1464 (N_1464,In_723,N_122);
or U1465 (N_1465,In_526,In_2679);
and U1466 (N_1466,N_342,In_1274);
or U1467 (N_1467,N_960,In_2888);
and U1468 (N_1468,In_2655,N_951);
and U1469 (N_1469,N_892,N_506);
nor U1470 (N_1470,N_995,N_228);
nor U1471 (N_1471,N_390,N_588);
and U1472 (N_1472,In_2635,N_841);
xor U1473 (N_1473,N_156,In_2465);
nand U1474 (N_1474,N_742,In_333);
nand U1475 (N_1475,N_1017,N_848);
xnor U1476 (N_1476,N_1071,In_2826);
or U1477 (N_1477,N_364,N_72);
nand U1478 (N_1478,N_781,N_15);
and U1479 (N_1479,N_55,N_643);
nand U1480 (N_1480,In_733,N_448);
xor U1481 (N_1481,N_26,N_276);
and U1482 (N_1482,N_664,N_1100);
nand U1483 (N_1483,In_2321,N_872);
or U1484 (N_1484,N_716,N_1098);
nand U1485 (N_1485,N_355,N_881);
xnor U1486 (N_1486,N_1187,N_888);
nand U1487 (N_1487,In_539,N_40);
and U1488 (N_1488,N_1192,N_877);
and U1489 (N_1489,In_717,N_507);
or U1490 (N_1490,In_1898,In_2527);
nand U1491 (N_1491,N_117,N_757);
nor U1492 (N_1492,In_1683,N_1150);
or U1493 (N_1493,N_333,N_1043);
xnor U1494 (N_1494,N_1117,In_1063);
and U1495 (N_1495,N_551,N_886);
nand U1496 (N_1496,N_934,In_557);
xnor U1497 (N_1497,N_295,N_492);
nor U1498 (N_1498,N_541,N_340);
or U1499 (N_1499,N_988,N_710);
nand U1500 (N_1500,N_210,N_656);
and U1501 (N_1501,N_130,N_1137);
nand U1502 (N_1502,N_48,In_176);
xnor U1503 (N_1503,In_2657,N_175);
nor U1504 (N_1504,N_752,N_591);
nand U1505 (N_1505,N_1001,N_849);
xor U1506 (N_1506,In_608,In_2988);
nand U1507 (N_1507,N_329,N_1109);
or U1508 (N_1508,In_406,In_278);
nand U1509 (N_1509,N_1086,N_516);
and U1510 (N_1510,N_309,In_704);
or U1511 (N_1511,In_1627,In_434);
and U1512 (N_1512,In_1333,In_803);
or U1513 (N_1513,N_816,N_491);
nand U1514 (N_1514,In_2478,In_826);
nand U1515 (N_1515,In_867,In_742);
or U1516 (N_1516,In_506,In_1829);
and U1517 (N_1517,N_404,In_2518);
xnor U1518 (N_1518,In_246,N_902);
or U1519 (N_1519,In_1844,In_160);
nor U1520 (N_1520,In_2969,N_1108);
nor U1521 (N_1521,N_611,N_1162);
and U1522 (N_1522,N_795,N_514);
and U1523 (N_1523,N_799,In_2341);
nor U1524 (N_1524,N_595,N_916);
xor U1525 (N_1525,N_824,N_1054);
or U1526 (N_1526,In_302,In_2390);
and U1527 (N_1527,N_952,In_1);
xor U1528 (N_1528,N_142,N_528);
xor U1529 (N_1529,In_1914,N_741);
or U1530 (N_1530,N_176,In_507);
and U1531 (N_1531,N_182,N_248);
nor U1532 (N_1532,N_468,N_769);
nor U1533 (N_1533,N_68,N_174);
xnor U1534 (N_1534,In_1158,In_1417);
and U1535 (N_1535,In_2229,In_2946);
nand U1536 (N_1536,N_1019,N_1182);
xor U1537 (N_1537,N_164,In_1329);
xor U1538 (N_1538,In_1602,In_2982);
and U1539 (N_1539,N_905,N_25);
xor U1540 (N_1540,N_831,N_610);
or U1541 (N_1541,N_534,In_2437);
and U1542 (N_1542,N_489,N_972);
nor U1543 (N_1543,In_1052,N_1175);
xor U1544 (N_1544,In_60,N_406);
xor U1545 (N_1545,N_693,N_527);
xnor U1546 (N_1546,N_110,N_132);
nand U1547 (N_1547,In_2363,N_380);
nor U1548 (N_1548,N_145,N_310);
nand U1549 (N_1549,In_2005,N_866);
xnor U1550 (N_1550,N_903,In_746);
and U1551 (N_1551,In_2124,N_915);
or U1552 (N_1552,N_259,N_1051);
and U1553 (N_1553,In_2565,N_719);
and U1554 (N_1554,N_967,In_2329);
nand U1555 (N_1555,N_925,N_662);
and U1556 (N_1556,N_1046,In_2431);
xor U1557 (N_1557,N_415,In_1634);
xnor U1558 (N_1558,N_857,N_684);
and U1559 (N_1559,In_1368,N_1111);
nand U1560 (N_1560,N_1083,N_1052);
or U1561 (N_1561,N_57,In_1031);
and U1562 (N_1562,N_91,N_1102);
or U1563 (N_1563,In_614,In_2375);
nor U1564 (N_1564,N_829,N_1116);
or U1565 (N_1565,N_87,In_161);
xnor U1566 (N_1566,N_483,In_2511);
nand U1567 (N_1567,N_240,N_95);
nand U1568 (N_1568,N_282,In_2992);
and U1569 (N_1569,N_965,In_1808);
nand U1570 (N_1570,N_157,In_1014);
and U1571 (N_1571,N_344,In_1931);
xnor U1572 (N_1572,N_1023,N_353);
or U1573 (N_1573,N_417,N_67);
and U1574 (N_1574,In_1246,In_2225);
and U1575 (N_1575,N_193,N_102);
and U1576 (N_1576,N_1130,N_343);
nor U1577 (N_1577,N_381,N_736);
and U1578 (N_1578,N_564,In_48);
xor U1579 (N_1579,In_1522,N_568);
xor U1580 (N_1580,In_326,N_485);
or U1581 (N_1581,N_424,In_1672);
xnor U1582 (N_1582,In_2318,N_451);
nand U1583 (N_1583,N_1085,N_844);
or U1584 (N_1584,In_1123,N_630);
or U1585 (N_1585,N_1159,N_105);
nand U1586 (N_1586,N_732,In_2514);
or U1587 (N_1587,N_1058,N_539);
xor U1588 (N_1588,N_1068,In_44);
nand U1589 (N_1589,N_984,N_121);
xor U1590 (N_1590,In_144,N_623);
nand U1591 (N_1591,N_478,In_2836);
nor U1592 (N_1592,N_761,In_1397);
nand U1593 (N_1593,N_457,N_1059);
nor U1594 (N_1594,N_247,N_970);
or U1595 (N_1595,N_35,N_760);
nand U1596 (N_1596,N_54,N_806);
and U1597 (N_1597,N_501,N_493);
xor U1598 (N_1598,In_2080,N_617);
and U1599 (N_1599,N_980,In_1629);
and U1600 (N_1600,N_426,N_1148);
and U1601 (N_1601,In_1502,N_75);
nor U1602 (N_1602,In_566,N_559);
or U1603 (N_1603,In_111,N_860);
nor U1604 (N_1604,N_413,N_334);
or U1605 (N_1605,In_2446,N_513);
or U1606 (N_1606,N_81,In_1353);
xnor U1607 (N_1607,N_753,N_416);
and U1608 (N_1608,In_263,N_974);
or U1609 (N_1609,N_153,N_521);
and U1610 (N_1610,N_356,N_287);
or U1611 (N_1611,In_2346,In_1120);
or U1612 (N_1612,In_1391,N_104);
or U1613 (N_1613,N_1143,N_1139);
nand U1614 (N_1614,N_926,N_243);
nand U1615 (N_1615,N_571,N_750);
nand U1616 (N_1616,N_1149,In_1478);
or U1617 (N_1617,N_1030,In_2091);
xnor U1618 (N_1618,In_42,N_1124);
nor U1619 (N_1619,In_2730,N_394);
nand U1620 (N_1620,N_580,In_1639);
and U1621 (N_1621,N_476,N_435);
and U1622 (N_1622,In_633,N_954);
nand U1623 (N_1623,In_508,N_885);
xor U1624 (N_1624,N_633,N_286);
nand U1625 (N_1625,N_794,N_62);
nand U1626 (N_1626,N_814,N_650);
nor U1627 (N_1627,In_2850,N_378);
or U1628 (N_1628,N_86,N_177);
xnor U1629 (N_1629,N_264,In_1003);
xnor U1630 (N_1630,N_522,N_893);
xor U1631 (N_1631,N_1080,N_127);
nor U1632 (N_1632,N_596,N_330);
xor U1633 (N_1633,N_730,N_918);
nand U1634 (N_1634,N_790,N_41);
or U1635 (N_1635,In_1260,In_1401);
nor U1636 (N_1636,N_178,N_300);
and U1637 (N_1637,In_68,N_348);
or U1638 (N_1638,N_151,In_2382);
or U1639 (N_1639,In_747,N_920);
and U1640 (N_1640,N_245,In_2032);
nand U1641 (N_1641,N_1127,N_961);
nand U1642 (N_1642,In_1142,In_1356);
or U1643 (N_1643,In_1132,In_1727);
xor U1644 (N_1644,N_1133,In_1458);
or U1645 (N_1645,In_1924,In_1831);
xnor U1646 (N_1646,N_238,In_1708);
and U1647 (N_1647,N_256,In_2128);
nor U1648 (N_1648,N_1196,In_2851);
nor U1649 (N_1649,In_2972,N_973);
or U1650 (N_1650,N_765,In_940);
nand U1651 (N_1651,N_520,N_810);
or U1652 (N_1652,In_1847,In_2973);
nor U1653 (N_1653,In_1588,N_1079);
and U1654 (N_1654,N_832,N_658);
or U1655 (N_1655,N_731,N_943);
xor U1656 (N_1656,N_702,N_850);
nand U1657 (N_1657,N_1110,N_97);
nand U1658 (N_1658,N_654,N_195);
xor U1659 (N_1659,N_707,N_303);
or U1660 (N_1660,N_313,N_92);
nor U1661 (N_1661,In_787,In_2881);
xor U1662 (N_1662,N_428,In_204);
xnor U1663 (N_1663,In_275,N_524);
xnor U1664 (N_1664,N_1096,N_308);
nor U1665 (N_1665,N_529,N_165);
xnor U1666 (N_1666,In_2723,N_1036);
nand U1667 (N_1667,N_632,N_1172);
nand U1668 (N_1668,In_1684,N_490);
nor U1669 (N_1669,N_154,N_602);
nand U1670 (N_1670,In_2327,In_724);
and U1671 (N_1671,N_657,N_397);
and U1672 (N_1672,N_430,N_346);
nand U1673 (N_1673,N_1062,In_2882);
and U1674 (N_1674,In_2048,N_1035);
nor U1675 (N_1675,In_347,In_2563);
or U1676 (N_1676,N_649,In_1807);
xnor U1677 (N_1677,In_1280,N_100);
and U1678 (N_1678,In_801,In_1514);
nor U1679 (N_1679,In_178,N_726);
or U1680 (N_1680,N_570,In_773);
xnor U1681 (N_1681,In_282,N_140);
nor U1682 (N_1682,N_819,In_1487);
or U1683 (N_1683,N_471,N_463);
nand U1684 (N_1684,N_258,N_962);
and U1685 (N_1685,N_512,N_399);
nor U1686 (N_1686,In_2731,N_89);
or U1687 (N_1687,N_1095,N_575);
xnor U1688 (N_1688,N_911,In_766);
xnor U1689 (N_1689,N_265,N_909);
xnor U1690 (N_1690,N_1134,N_843);
nor U1691 (N_1691,N_989,In_1079);
nor U1692 (N_1692,In_2416,In_825);
or U1693 (N_1693,In_1124,N_937);
or U1694 (N_1694,N_101,N_197);
xor U1695 (N_1695,N_30,N_780);
nand U1696 (N_1696,N_365,N_1010);
xor U1697 (N_1697,N_335,In_488);
and U1698 (N_1698,N_74,In_2786);
and U1699 (N_1699,N_370,In_301);
xor U1700 (N_1700,In_2422,In_316);
and U1701 (N_1701,N_563,N_1160);
nand U1702 (N_1702,N_901,N_453);
nand U1703 (N_1703,N_367,In_1911);
or U1704 (N_1704,N_712,In_2797);
and U1705 (N_1705,N_339,In_999);
or U1706 (N_1706,In_2008,N_826);
and U1707 (N_1707,N_1181,In_1190);
or U1708 (N_1708,N_146,In_980);
or U1709 (N_1709,In_2822,N_411);
nor U1710 (N_1710,N_352,In_1018);
nor U1711 (N_1711,N_690,In_1328);
nand U1712 (N_1712,N_927,N_16);
and U1713 (N_1713,N_589,N_56);
nand U1714 (N_1714,N_1006,N_45);
or U1715 (N_1715,N_11,N_1047);
xnor U1716 (N_1716,In_2784,N_1039);
nand U1717 (N_1717,N_729,N_899);
xnor U1718 (N_1718,N_533,N_137);
or U1719 (N_1719,N_587,N_218);
or U1720 (N_1720,In_30,In_2906);
nand U1721 (N_1721,N_771,N_96);
and U1722 (N_1722,N_214,N_639);
and U1723 (N_1723,N_293,N_1197);
nand U1724 (N_1724,In_1310,N_721);
nand U1725 (N_1725,N_801,N_203);
xnor U1726 (N_1726,In_577,N_1074);
nand U1727 (N_1727,N_192,N_605);
xnor U1728 (N_1728,N_266,N_1168);
or U1729 (N_1729,N_403,N_398);
nor U1730 (N_1730,N_636,N_98);
or U1731 (N_1731,N_696,In_2872);
and U1732 (N_1732,In_1086,In_617);
nor U1733 (N_1733,N_884,N_431);
and U1734 (N_1734,In_2296,N_289);
xnor U1735 (N_1735,In_1816,N_149);
nor U1736 (N_1736,N_1078,In_2706);
or U1737 (N_1737,N_307,N_778);
or U1738 (N_1738,N_777,N_268);
nor U1739 (N_1739,In_1313,N_38);
nor U1740 (N_1740,N_273,N_290);
nand U1741 (N_1741,In_353,N_78);
nand U1742 (N_1742,N_978,In_1127);
nand U1743 (N_1743,N_833,N_767);
nor U1744 (N_1744,In_265,In_2572);
xor U1745 (N_1745,In_497,N_941);
nand U1746 (N_1746,In_1546,N_1136);
xor U1747 (N_1747,N_419,N_608);
or U1748 (N_1748,N_205,In_789);
nand U1749 (N_1749,In_2762,In_1504);
nor U1750 (N_1750,N_613,In_293);
nor U1751 (N_1751,N_945,In_2244);
or U1752 (N_1752,In_2579,N_226);
nand U1753 (N_1753,N_536,N_1057);
xor U1754 (N_1754,In_2022,In_1362);
nor U1755 (N_1755,N_449,In_147);
xor U1756 (N_1756,N_262,In_261);
and U1757 (N_1757,N_366,In_1824);
nor U1758 (N_1758,N_817,N_985);
nand U1759 (N_1759,N_766,N_562);
nand U1760 (N_1760,N_1008,N_673);
and U1761 (N_1761,N_635,N_560);
nand U1762 (N_1762,In_956,N_434);
xor U1763 (N_1763,In_920,In_1290);
or U1764 (N_1764,N_793,In_1452);
or U1765 (N_1765,N_114,N_168);
xor U1766 (N_1766,N_429,N_791);
nor U1767 (N_1767,N_959,In_1029);
nand U1768 (N_1768,N_621,N_626);
or U1769 (N_1769,N_1024,N_852);
nor U1770 (N_1770,N_160,N_446);
nand U1771 (N_1771,In_480,N_692);
nor U1772 (N_1772,In_1674,N_124);
nand U1773 (N_1773,N_590,N_1021);
or U1774 (N_1774,In_2594,In_58);
xor U1775 (N_1775,N_73,N_1056);
and U1776 (N_1776,In_1665,In_856);
nor U1777 (N_1777,In_49,In_2905);
and U1778 (N_1778,N_470,N_686);
xnor U1779 (N_1779,In_2007,N_1013);
nor U1780 (N_1780,N_338,N_213);
nor U1781 (N_1781,In_1910,N_880);
nand U1782 (N_1782,N_668,N_138);
and U1783 (N_1783,In_2364,In_1575);
nand U1784 (N_1784,N_125,N_20);
xnor U1785 (N_1785,N_131,In_731);
nand U1786 (N_1786,In_2557,N_553);
or U1787 (N_1787,N_594,In_2607);
and U1788 (N_1788,N_445,In_1134);
nand U1789 (N_1789,In_271,N_61);
and U1790 (N_1790,In_2792,In_1317);
nor U1791 (N_1791,In_562,N_460);
nand U1792 (N_1792,In_2368,In_2707);
nand U1793 (N_1793,N_547,N_953);
nor U1794 (N_1794,N_351,N_538);
nand U1795 (N_1795,In_1638,N_734);
nand U1796 (N_1796,In_1341,N_474);
nor U1797 (N_1797,N_1179,N_270);
and U1798 (N_1798,N_695,N_955);
nor U1799 (N_1799,N_128,N_1169);
and U1800 (N_1800,N_825,N_1012);
nor U1801 (N_1801,N_354,In_1434);
xnor U1802 (N_1802,N_762,N_931);
nor U1803 (N_1803,N_976,N_162);
or U1804 (N_1804,In_989,N_179);
nor U1805 (N_1805,N_879,N_548);
xor U1806 (N_1806,N_190,N_49);
nor U1807 (N_1807,N_720,N_628);
and U1808 (N_1808,In_159,N_63);
or U1809 (N_1809,N_19,In_1617);
and U1810 (N_1810,N_640,In_2078);
or U1811 (N_1811,In_2812,N_775);
xor U1812 (N_1812,N_297,N_371);
nand U1813 (N_1813,N_8,N_645);
nand U1814 (N_1814,N_818,N_1);
xor U1815 (N_1815,In_54,N_316);
nor U1816 (N_1816,N_503,In_569);
or U1817 (N_1817,N_968,N_271);
and U1818 (N_1818,N_1015,In_1747);
xor U1819 (N_1819,In_875,N_1135);
or U1820 (N_1820,In_2843,N_447);
or U1821 (N_1821,N_69,N_874);
xnor U1822 (N_1822,N_198,In_2606);
and U1823 (N_1823,N_1055,N_400);
or U1824 (N_1824,N_39,In_744);
nor U1825 (N_1825,N_347,In_1694);
nor U1826 (N_1826,N_422,N_647);
nand U1827 (N_1827,N_217,N_201);
nor U1828 (N_1828,N_620,N_234);
nand U1829 (N_1829,N_252,In_889);
xor U1830 (N_1830,N_847,N_4);
nor U1831 (N_1831,N_1089,N_65);
nor U1832 (N_1832,N_169,In_901);
and U1833 (N_1833,N_908,In_814);
nor U1834 (N_1834,In_2119,N_28);
or U1835 (N_1835,N_200,N_51);
nand U1836 (N_1836,N_839,In_1000);
xor U1837 (N_1837,N_32,N_685);
or U1838 (N_1838,In_50,N_155);
nand U1839 (N_1839,In_2046,N_320);
nor U1840 (N_1840,In_997,In_2331);
nand U1841 (N_1841,In_1144,In_2090);
or U1842 (N_1842,In_762,N_482);
and U1843 (N_1843,N_497,N_958);
nor U1844 (N_1844,N_897,In_1410);
nand U1845 (N_1845,In_72,N_70);
and U1846 (N_1846,In_2361,In_2746);
and U1847 (N_1847,In_2643,In_2040);
xor U1848 (N_1848,In_1986,In_597);
and U1849 (N_1849,In_448,In_2605);
xor U1850 (N_1850,In_2117,N_108);
nand U1851 (N_1851,N_504,N_1177);
and U1852 (N_1852,N_1103,N_207);
nand U1853 (N_1853,In_1846,In_1211);
nor U1854 (N_1854,N_718,N_1183);
xor U1855 (N_1855,N_648,N_43);
xnor U1856 (N_1856,N_1097,N_964);
xor U1857 (N_1857,In_1799,In_1820);
xnor U1858 (N_1858,N_386,In_2699);
nand U1859 (N_1859,N_1048,N_577);
xnor U1860 (N_1860,In_1493,N_975);
nand U1861 (N_1861,N_500,N_573);
nand U1862 (N_1862,In_2582,N_472);
nor U1863 (N_1863,N_196,In_352);
nor U1864 (N_1864,In_2584,N_239);
and U1865 (N_1865,In_1519,In_1780);
nor U1866 (N_1866,In_460,N_1190);
nand U1867 (N_1867,N_557,In_108);
xnor U1868 (N_1868,In_660,N_22);
nand U1869 (N_1869,N_1066,N_1065);
or U1870 (N_1870,N_279,In_1566);
and U1871 (N_1871,N_998,N_622);
or U1872 (N_1872,In_1795,In_1959);
xnor U1873 (N_1873,In_351,In_306);
nor U1874 (N_1874,N_871,N_479);
or U1875 (N_1875,In_852,N_350);
xor U1876 (N_1876,N_323,In_1231);
xnor U1877 (N_1877,In_1418,N_887);
and U1878 (N_1878,N_1022,In_1729);
or U1879 (N_1879,N_537,N_1125);
xor U1880 (N_1880,In_2577,In_2414);
or U1881 (N_1881,N_822,In_1360);
or U1882 (N_1882,N_421,N_312);
or U1883 (N_1883,N_540,N_116);
nand U1884 (N_1884,N_746,N_277);
xor U1885 (N_1885,In_2547,N_944);
and U1886 (N_1886,N_272,N_957);
or U1887 (N_1887,N_1122,N_796);
xor U1888 (N_1888,N_525,N_1189);
xor U1889 (N_1889,N_236,N_1018);
or U1890 (N_1890,N_1154,N_1176);
nand U1891 (N_1891,N_144,N_1131);
and U1892 (N_1892,N_733,N_231);
xnor U1893 (N_1893,In_705,In_1611);
or U1894 (N_1894,N_802,N_987);
xnor U1895 (N_1895,N_384,N_1104);
nor U1896 (N_1896,N_27,N_856);
nand U1897 (N_1897,N_938,N_59);
nor U1898 (N_1898,In_2752,N_458);
or U1899 (N_1899,N_838,N_747);
nor U1900 (N_1900,N_222,N_2);
or U1901 (N_1901,N_1064,N_904);
and U1902 (N_1902,N_776,In_2837);
nand U1903 (N_1903,N_604,N_269);
nand U1904 (N_1904,N_606,In_2338);
nor U1905 (N_1905,N_1118,N_499);
or U1906 (N_1906,In_738,In_1436);
nand U1907 (N_1907,N_700,N_496);
and U1908 (N_1908,N_807,N_5);
xor U1909 (N_1909,N_1050,N_919);
or U1910 (N_1910,N_368,N_1082);
xor U1911 (N_1911,In_2924,N_517);
and U1912 (N_1912,N_1173,N_437);
xnor U1913 (N_1913,In_1070,In_1965);
nor U1914 (N_1914,In_2386,N_917);
nand U1915 (N_1915,N_907,N_665);
and U1916 (N_1916,In_2780,In_192);
xor U1917 (N_1917,N_785,N_1040);
and U1918 (N_1918,N_443,N_1167);
nor U1919 (N_1919,N_727,N_58);
xnor U1920 (N_1920,N_232,N_555);
nor U1921 (N_1921,N_603,N_542);
nor U1922 (N_1922,N_932,N_609);
xor U1923 (N_1923,N_1094,N_1028);
and U1924 (N_1924,N_858,In_518);
or U1925 (N_1925,In_905,In_1462);
and U1926 (N_1926,In_1420,N_33);
nand U1927 (N_1927,N_12,In_1291);
or U1928 (N_1928,In_1389,In_2492);
nor U1929 (N_1929,N_1053,N_487);
and U1930 (N_1930,N_535,In_484);
and U1931 (N_1931,N_94,In_3);
xor U1932 (N_1932,N_1038,N_725);
xnor U1933 (N_1933,N_979,In_1441);
xnor U1934 (N_1934,N_813,N_1070);
xnor U1935 (N_1935,In_722,N_585);
and U1936 (N_1936,In_1915,N_129);
or U1937 (N_1937,In_2417,In_1640);
xnor U1938 (N_1938,N_439,N_914);
xor U1939 (N_1939,In_156,N_159);
and U1940 (N_1940,In_2552,In_1839);
xnor U1941 (N_1941,N_940,N_835);
and U1942 (N_1942,N_774,N_651);
or U1943 (N_1943,In_98,N_947);
and U1944 (N_1944,In_1534,In_1151);
or U1945 (N_1945,In_2844,In_2865);
nor U1946 (N_1946,N_1099,In_1528);
xnor U1947 (N_1947,In_2213,N_462);
or U1948 (N_1948,In_1265,N_473);
and U1949 (N_1949,N_1027,In_1920);
xnor U1950 (N_1950,In_2095,N_255);
or U1951 (N_1951,N_107,N_183);
or U1952 (N_1952,N_119,In_471);
nand U1953 (N_1953,In_1594,N_498);
xor U1954 (N_1954,N_759,N_202);
nor U1955 (N_1955,N_1020,N_1004);
xnor U1956 (N_1956,N_1093,N_875);
and U1957 (N_1957,N_322,N_1105);
or U1958 (N_1958,N_519,In_2397);
or U1959 (N_1959,N_249,N_1180);
xnor U1960 (N_1960,In_1603,In_2248);
nor U1961 (N_1961,N_1003,N_788);
nand U1962 (N_1962,In_2798,N_410);
nand U1963 (N_1963,N_950,In_2298);
and U1964 (N_1964,N_391,N_667);
nand U1965 (N_1965,N_332,N_141);
nand U1966 (N_1966,N_846,In_2185);
and U1967 (N_1967,N_800,N_675);
nand U1968 (N_1968,N_981,N_1107);
and U1969 (N_1969,N_855,N_688);
nor U1970 (N_1970,N_36,In_495);
xnor U1971 (N_1971,N_815,In_1969);
nor U1972 (N_1972,N_898,N_723);
or U1973 (N_1973,N_631,N_136);
nand U1974 (N_1974,N_244,In_846);
xor U1975 (N_1975,N_999,In_1817);
and U1976 (N_1976,N_209,N_1157);
nand U1977 (N_1977,N_928,In_1108);
nand U1978 (N_1978,N_120,N_745);
nand U1979 (N_1979,N_1155,N_171);
or U1980 (N_1980,N_784,In_2141);
and U1981 (N_1981,N_680,N_281);
xnor U1982 (N_1982,In_268,In_1021);
nand U1983 (N_1983,In_942,N_672);
nand U1984 (N_1984,N_546,N_763);
and U1985 (N_1985,N_111,N_1009);
nand U1986 (N_1986,In_2271,N_306);
and U1987 (N_1987,N_388,In_2877);
xnor U1988 (N_1988,N_274,In_430);
and U1989 (N_1989,In_1610,In_224);
xnor U1990 (N_1990,In_195,N_379);
xor U1991 (N_1991,In_2949,N_687);
and U1992 (N_1992,In_2263,N_321);
nand U1993 (N_1993,N_173,N_592);
nand U1994 (N_1994,In_1320,In_931);
or U1995 (N_1995,N_992,N_60);
and U1996 (N_1996,N_740,N_515);
nor U1997 (N_1997,N_933,N_185);
nor U1998 (N_1998,N_811,N_254);
nand U1999 (N_1999,N_250,N_14);
and U2000 (N_2000,In_1767,In_2620);
and U2001 (N_2001,N_894,In_1512);
and U2002 (N_2002,N_505,N_1156);
and U2003 (N_2003,N_634,N_653);
or U2004 (N_2004,N_393,N_336);
nor U2005 (N_2005,N_666,N_242);
nand U2006 (N_2006,In_402,In_2349);
nand U2007 (N_2007,N_735,N_1014);
nor U2008 (N_2008,In_1908,N_930);
and U2009 (N_2009,N_1044,N_235);
xor U2010 (N_2010,In_379,In_2357);
nand U2011 (N_2011,In_238,N_971);
nand U2012 (N_2012,In_1981,In_1270);
xor U2013 (N_2013,In_1030,N_1060);
xnor U2014 (N_2014,In_1590,N_678);
nand U2015 (N_2015,N_896,In_1557);
and U2016 (N_2016,N_787,In_1471);
nand U2017 (N_2017,In_2904,N_550);
nand U2018 (N_2018,In_2353,In_2176);
and U2019 (N_2019,In_1746,In_2049);
nand U2020 (N_2020,In_2777,N_889);
nor U2021 (N_2021,N_360,N_484);
xor U2022 (N_2022,N_324,N_199);
nand U2023 (N_2023,In_2146,N_509);
xnor U2024 (N_2024,N_311,N_126);
and U2025 (N_2025,N_836,N_677);
xnor U2026 (N_2026,N_808,N_956);
nand U2027 (N_2027,N_638,N_181);
and U2028 (N_2028,In_2927,N_545);
xor U2029 (N_2029,In_1295,N_579);
and U2030 (N_2030,N_337,N_29);
nand U2031 (N_2031,N_642,N_1174);
and U2032 (N_2032,N_715,In_685);
nor U2033 (N_2033,N_565,N_900);
nand U2034 (N_2034,N_809,N_1152);
or U2035 (N_2035,N_34,N_1198);
and U2036 (N_2036,N_1147,In_2121);
xor U2037 (N_2037,N_407,N_1011);
xor U2038 (N_2038,N_377,N_1171);
and U2039 (N_2039,N_698,N_773);
xnor U2040 (N_2040,In_1253,N_53);
and U2041 (N_2041,In_1307,In_1664);
and U2042 (N_2042,N_251,In_2231);
nand U2043 (N_2043,In_1953,In_2652);
or U2044 (N_2044,N_582,N_646);
nand U2045 (N_2045,N_319,In_77);
and U2046 (N_2046,N_1138,N_923);
xor U2047 (N_2047,N_779,N_325);
xor U2048 (N_2048,N_71,In_1997);
or U2049 (N_2049,In_1771,In_758);
or U2050 (N_2050,N_572,In_1984);
nor U2051 (N_2051,N_597,In_325);
nor U2052 (N_2052,N_895,N_624);
nand U2053 (N_2053,In_763,N_215);
nor U2054 (N_2054,In_2436,N_705);
nor U2055 (N_2055,In_203,In_2217);
nor U2056 (N_2056,N_77,N_392);
or U2057 (N_2057,N_783,In_1941);
xnor U2058 (N_2058,N_797,In_1481);
and U2059 (N_2059,N_990,In_1572);
nor U2060 (N_2060,N_983,N_581);
nand U2061 (N_2061,In_1433,N_292);
xnor U2062 (N_2062,In_2899,N_523);
nand U2063 (N_2063,In_2438,N_314);
nor U2064 (N_2064,N_756,N_369);
and U2065 (N_2065,In_1484,N_556);
nor U2066 (N_2066,N_7,In_2631);
nor U2067 (N_2067,N_764,N_1016);
nor U2068 (N_2068,N_612,N_93);
nor U2069 (N_2069,In_1245,N_1092);
xor U2070 (N_2070,N_786,N_922);
nor U2071 (N_2071,N_859,N_869);
and U2072 (N_2072,In_954,In_1412);
nand U2073 (N_2073,N_1002,N_586);
nand U2074 (N_2074,N_464,N_304);
xnor U2075 (N_2075,N_284,N_676);
nor U2076 (N_2076,N_1084,In_1195);
xor U2077 (N_2077,N_112,N_79);
and U2078 (N_2078,N_804,N_167);
xor U2079 (N_2079,N_216,In_1257);
xor U2080 (N_2080,N_659,In_1383);
and U2081 (N_2081,N_341,In_2404);
nand U2082 (N_2082,In_438,N_420);
or U2083 (N_2083,N_966,N_994);
and U2084 (N_2084,N_598,In_2469);
or U2085 (N_2085,In_2742,N_935);
xor U2086 (N_2086,N_414,In_523);
or U2087 (N_2087,N_327,N_1090);
nor U2088 (N_2088,N_221,N_714);
xnor U2089 (N_2089,In_1762,N_163);
or U2090 (N_2090,N_1145,N_812);
or U2091 (N_2091,In_2914,N_23);
nand U2092 (N_2092,N_10,N_184);
or U2093 (N_2093,In_2283,N_913);
or U2094 (N_2094,N_670,In_362);
and U2095 (N_2095,N_3,N_46);
nand U2096 (N_2096,In_1489,N_576);
nor U2097 (N_2097,N_511,N_566);
or U2098 (N_2098,N_870,N_601);
or U2099 (N_2099,N_986,N_83);
nor U2100 (N_2100,N_549,N_597);
xor U2101 (N_2101,N_1110,N_664);
nand U2102 (N_2102,N_22,N_919);
and U2103 (N_2103,N_716,N_1159);
xor U2104 (N_2104,In_2553,In_2742);
nand U2105 (N_2105,In_1123,N_138);
and U2106 (N_2106,N_720,N_845);
or U2107 (N_2107,In_1420,N_502);
nand U2108 (N_2108,In_2010,N_1071);
xor U2109 (N_2109,N_1000,N_554);
nand U2110 (N_2110,In_326,N_397);
or U2111 (N_2111,N_981,In_2914);
nor U2112 (N_2112,In_2361,N_534);
or U2113 (N_2113,N_1178,N_1094);
nor U2114 (N_2114,N_350,In_2115);
nand U2115 (N_2115,In_2904,N_138);
nor U2116 (N_2116,N_147,In_1391);
nand U2117 (N_2117,N_509,In_2097);
nor U2118 (N_2118,N_642,In_246);
xor U2119 (N_2119,N_478,N_991);
xor U2120 (N_2120,N_806,In_2557);
nand U2121 (N_2121,N_287,In_1919);
and U2122 (N_2122,N_707,N_58);
nand U2123 (N_2123,In_147,N_349);
and U2124 (N_2124,In_58,N_32);
and U2125 (N_2125,N_920,N_193);
xor U2126 (N_2126,N_866,N_1121);
nor U2127 (N_2127,N_1010,N_765);
nor U2128 (N_2128,In_1486,N_372);
and U2129 (N_2129,N_8,N_654);
nor U2130 (N_2130,In_766,N_1009);
or U2131 (N_2131,N_648,In_1463);
or U2132 (N_2132,N_1136,N_279);
nand U2133 (N_2133,In_1003,In_2746);
nand U2134 (N_2134,N_115,N_70);
and U2135 (N_2135,N_950,N_179);
or U2136 (N_2136,N_1196,N_714);
nand U2137 (N_2137,In_1320,N_1180);
or U2138 (N_2138,N_743,In_2872);
and U2139 (N_2139,N_212,N_507);
xor U2140 (N_2140,N_422,N_882);
nor U2141 (N_2141,N_1193,N_638);
nor U2142 (N_2142,In_720,N_7);
nor U2143 (N_2143,In_2127,N_773);
xnor U2144 (N_2144,N_1047,N_946);
xor U2145 (N_2145,In_1984,N_522);
nor U2146 (N_2146,In_2353,N_220);
or U2147 (N_2147,N_866,N_789);
and U2148 (N_2148,N_762,In_1893);
or U2149 (N_2149,In_2882,N_105);
nor U2150 (N_2150,N_135,N_398);
and U2151 (N_2151,In_2387,N_571);
and U2152 (N_2152,In_325,N_778);
nor U2153 (N_2153,In_2577,In_2273);
and U2154 (N_2154,N_685,N_391);
or U2155 (N_2155,N_419,In_2907);
or U2156 (N_2156,N_1047,In_2217);
xor U2157 (N_2157,N_445,N_289);
xor U2158 (N_2158,N_897,N_1086);
and U2159 (N_2159,N_505,N_616);
or U2160 (N_2160,In_1487,N_336);
xor U2161 (N_2161,In_480,N_920);
or U2162 (N_2162,In_2777,N_1009);
or U2163 (N_2163,In_30,N_567);
nor U2164 (N_2164,N_500,N_714);
and U2165 (N_2165,In_942,In_2414);
nand U2166 (N_2166,In_2090,In_1471);
or U2167 (N_2167,In_1504,N_1034);
or U2168 (N_2168,N_1070,N_45);
or U2169 (N_2169,N_689,N_821);
or U2170 (N_2170,N_724,N_842);
and U2171 (N_2171,In_1328,N_72);
nand U2172 (N_2172,N_594,N_984);
and U2173 (N_2173,N_1073,N_1145);
and U2174 (N_2174,In_999,N_666);
nand U2175 (N_2175,In_2735,N_722);
and U2176 (N_2176,In_1557,N_758);
xor U2177 (N_2177,N_390,In_2091);
xor U2178 (N_2178,N_346,N_302);
and U2179 (N_2179,N_680,In_2478);
nand U2180 (N_2180,N_643,In_895);
xnor U2181 (N_2181,In_1063,N_546);
nor U2182 (N_2182,N_284,N_563);
or U2183 (N_2183,In_2607,In_665);
and U2184 (N_2184,N_1159,In_1452);
nand U2185 (N_2185,In_1965,N_501);
nor U2186 (N_2186,N_84,N_143);
and U2187 (N_2187,N_97,In_762);
xnor U2188 (N_2188,In_353,N_1020);
xnor U2189 (N_2189,N_1125,In_1031);
xnor U2190 (N_2190,N_105,In_1772);
and U2191 (N_2191,In_1458,N_689);
xnor U2192 (N_2192,N_1014,In_203);
nand U2193 (N_2193,N_670,N_901);
xnor U2194 (N_2194,In_608,N_806);
or U2195 (N_2195,N_351,In_1747);
xnor U2196 (N_2196,In_2394,In_178);
xnor U2197 (N_2197,In_1190,N_1161);
and U2198 (N_2198,In_1235,N_606);
nand U2199 (N_2199,In_2836,N_550);
nor U2200 (N_2200,In_2657,In_1422);
xor U2201 (N_2201,N_984,N_49);
or U2202 (N_2202,N_951,In_1514);
xor U2203 (N_2203,N_575,In_26);
xor U2204 (N_2204,In_610,In_1684);
xnor U2205 (N_2205,N_803,N_33);
nand U2206 (N_2206,N_308,N_994);
xnor U2207 (N_2207,N_1142,N_549);
and U2208 (N_2208,N_932,N_558);
nor U2209 (N_2209,N_101,N_1018);
nor U2210 (N_2210,N_270,N_798);
nand U2211 (N_2211,N_903,N_219);
or U2212 (N_2212,N_674,In_723);
nor U2213 (N_2213,In_381,N_618);
and U2214 (N_2214,In_882,N_819);
or U2215 (N_2215,N_120,In_2383);
xnor U2216 (N_2216,N_1172,N_883);
nor U2217 (N_2217,N_657,N_1119);
or U2218 (N_2218,N_963,N_1032);
or U2219 (N_2219,N_486,N_172);
nand U2220 (N_2220,N_1103,N_106);
nand U2221 (N_2221,N_134,N_800);
nor U2222 (N_2222,N_350,N_694);
xnor U2223 (N_2223,N_1062,N_749);
nor U2224 (N_2224,N_886,N_1086);
xor U2225 (N_2225,N_993,N_998);
or U2226 (N_2226,N_133,N_91);
nor U2227 (N_2227,N_922,In_2547);
or U2228 (N_2228,N_1083,N_1018);
xnor U2229 (N_2229,In_2843,N_144);
nor U2230 (N_2230,N_897,N_40);
nor U2231 (N_2231,In_2636,In_2271);
and U2232 (N_2232,In_704,N_261);
and U2233 (N_2233,N_306,N_913);
and U2234 (N_2234,N_439,N_8);
nand U2235 (N_2235,In_1746,N_1103);
or U2236 (N_2236,In_557,N_263);
or U2237 (N_2237,N_88,N_300);
or U2238 (N_2238,N_334,N_711);
nor U2239 (N_2239,N_745,N_363);
or U2240 (N_2240,N_221,N_254);
nand U2241 (N_2241,In_2397,N_1144);
and U2242 (N_2242,N_23,In_2949);
nor U2243 (N_2243,N_1102,N_72);
nor U2244 (N_2244,N_499,In_1190);
xnor U2245 (N_2245,N_290,N_852);
and U2246 (N_2246,N_783,N_354);
nor U2247 (N_2247,N_654,In_1173);
nor U2248 (N_2248,In_2481,In_2046);
nand U2249 (N_2249,N_103,In_1981);
nand U2250 (N_2250,N_442,In_2327);
nor U2251 (N_2251,N_614,N_842);
nor U2252 (N_2252,In_747,In_1601);
nand U2253 (N_2253,N_103,In_2022);
xnor U2254 (N_2254,In_2364,N_80);
xor U2255 (N_2255,In_1070,In_2233);
and U2256 (N_2256,N_260,N_287);
nor U2257 (N_2257,In_895,N_521);
and U2258 (N_2258,N_419,N_910);
or U2259 (N_2259,N_113,In_1039);
xor U2260 (N_2260,N_330,N_291);
nand U2261 (N_2261,N_1196,N_416);
or U2262 (N_2262,In_2826,In_82);
or U2263 (N_2263,In_2655,In_1986);
nand U2264 (N_2264,In_2527,N_300);
nand U2265 (N_2265,In_1727,N_920);
xnor U2266 (N_2266,In_2924,N_976);
nand U2267 (N_2267,N_183,N_459);
or U2268 (N_2268,In_147,N_244);
or U2269 (N_2269,N_640,N_786);
and U2270 (N_2270,In_1795,In_1634);
or U2271 (N_2271,N_425,N_710);
xnor U2272 (N_2272,In_1003,In_471);
nor U2273 (N_2273,N_100,N_532);
xnor U2274 (N_2274,N_607,N_876);
and U2275 (N_2275,N_516,N_488);
and U2276 (N_2276,In_989,N_509);
nor U2277 (N_2277,N_1056,N_178);
or U2278 (N_2278,In_2233,In_1433);
nand U2279 (N_2279,N_425,N_1032);
xor U2280 (N_2280,N_473,N_87);
and U2281 (N_2281,N_508,N_908);
xor U2282 (N_2282,N_798,In_2364);
and U2283 (N_2283,N_442,N_124);
and U2284 (N_2284,In_1672,N_981);
nand U2285 (N_2285,N_41,N_1051);
or U2286 (N_2286,N_641,N_987);
nand U2287 (N_2287,In_2904,N_744);
nand U2288 (N_2288,In_2047,In_931);
nand U2289 (N_2289,N_85,N_722);
nor U2290 (N_2290,In_261,N_1119);
or U2291 (N_2291,N_223,N_873);
xor U2292 (N_2292,In_569,N_691);
or U2293 (N_2293,N_849,N_246);
and U2294 (N_2294,N_1072,In_2514);
xnor U2295 (N_2295,In_746,N_411);
nor U2296 (N_2296,N_7,N_1043);
xor U2297 (N_2297,N_743,In_1001);
xnor U2298 (N_2298,N_114,In_2730);
nor U2299 (N_2299,N_941,In_997);
and U2300 (N_2300,N_521,N_412);
or U2301 (N_2301,In_2386,In_497);
or U2302 (N_2302,N_176,N_258);
and U2303 (N_2303,In_1029,N_864);
or U2304 (N_2304,N_536,In_838);
nor U2305 (N_2305,N_948,N_931);
xnor U2306 (N_2306,N_910,In_2124);
nor U2307 (N_2307,N_881,In_368);
nand U2308 (N_2308,N_963,N_309);
and U2309 (N_2309,In_920,N_778);
xnor U2310 (N_2310,In_1715,In_1585);
and U2311 (N_2311,N_450,N_258);
nor U2312 (N_2312,N_471,In_1328);
xor U2313 (N_2313,N_761,N_98);
or U2314 (N_2314,N_557,In_2346);
xor U2315 (N_2315,In_58,N_1145);
nor U2316 (N_2316,N_1104,N_1030);
and U2317 (N_2317,N_882,N_263);
xor U2318 (N_2318,N_1124,In_608);
nand U2319 (N_2319,N_815,In_205);
nand U2320 (N_2320,N_940,In_2225);
nand U2321 (N_2321,N_367,In_766);
xnor U2322 (N_2322,N_729,In_2762);
and U2323 (N_2323,N_795,In_1672);
or U2324 (N_2324,N_1052,N_955);
and U2325 (N_2325,N_438,N_886);
or U2326 (N_2326,In_1816,In_2489);
or U2327 (N_2327,N_1009,N_1150);
nor U2328 (N_2328,N_631,In_577);
nand U2329 (N_2329,N_510,In_908);
and U2330 (N_2330,In_2047,In_633);
nand U2331 (N_2331,N_1017,N_975);
xor U2332 (N_2332,N_640,N_779);
xor U2333 (N_2333,N_986,In_758);
or U2334 (N_2334,In_2321,N_11);
or U2335 (N_2335,In_2786,In_1180);
or U2336 (N_2336,N_361,N_588);
nand U2337 (N_2337,N_350,N_779);
xnor U2338 (N_2338,N_14,N_761);
or U2339 (N_2339,N_833,N_911);
nand U2340 (N_2340,In_506,N_1084);
and U2341 (N_2341,N_318,N_93);
and U2342 (N_2342,N_920,N_1128);
nand U2343 (N_2343,N_378,N_162);
and U2344 (N_2344,N_1021,In_1497);
or U2345 (N_2345,N_118,N_870);
xor U2346 (N_2346,In_2279,N_998);
nor U2347 (N_2347,N_596,N_418);
nand U2348 (N_2348,In_1534,In_2907);
nand U2349 (N_2349,N_567,N_385);
nand U2350 (N_2350,In_2699,In_495);
nand U2351 (N_2351,N_394,In_435);
nor U2352 (N_2352,N_446,In_1602);
xnor U2353 (N_2353,N_433,N_648);
nor U2354 (N_2354,N_5,N_932);
and U2355 (N_2355,N_1118,N_386);
nor U2356 (N_2356,N_687,N_558);
and U2357 (N_2357,N_792,N_598);
nor U2358 (N_2358,In_2730,N_321);
and U2359 (N_2359,N_831,In_733);
or U2360 (N_2360,In_2331,N_106);
and U2361 (N_2361,N_1018,N_228);
xnor U2362 (N_2362,N_1040,In_2969);
or U2363 (N_2363,N_1131,In_1493);
or U2364 (N_2364,In_2090,In_2851);
nor U2365 (N_2365,In_1452,N_1151);
or U2366 (N_2366,In_1070,In_1462);
or U2367 (N_2367,In_161,N_697);
or U2368 (N_2368,N_972,In_58);
xor U2369 (N_2369,In_2798,N_59);
and U2370 (N_2370,N_429,N_1057);
xor U2371 (N_2371,N_1016,N_597);
and U2372 (N_2372,N_700,N_1039);
nand U2373 (N_2373,N_118,In_1389);
xor U2374 (N_2374,In_1291,N_425);
nor U2375 (N_2375,In_1418,N_901);
and U2376 (N_2376,N_20,N_556);
xnor U2377 (N_2377,N_1036,N_101);
nor U2378 (N_2378,In_2338,N_313);
nor U2379 (N_2379,N_380,N_838);
nor U2380 (N_2380,N_992,N_837);
and U2381 (N_2381,N_660,N_825);
nand U2382 (N_2382,N_525,N_10);
nor U2383 (N_2383,N_1123,N_259);
or U2384 (N_2384,N_1107,N_295);
and U2385 (N_2385,N_547,In_2318);
and U2386 (N_2386,N_590,In_2382);
xnor U2387 (N_2387,N_860,N_885);
and U2388 (N_2388,In_1694,In_2008);
xor U2389 (N_2389,N_1086,In_434);
or U2390 (N_2390,N_37,In_2518);
and U2391 (N_2391,N_1153,In_285);
or U2392 (N_2392,In_2655,In_2078);
nand U2393 (N_2393,In_2357,N_279);
or U2394 (N_2394,N_141,In_1455);
or U2395 (N_2395,N_48,N_86);
and U2396 (N_2396,In_1014,In_2244);
xnor U2397 (N_2397,N_694,N_441);
nand U2398 (N_2398,In_2882,N_1009);
nand U2399 (N_2399,N_1025,In_1412);
nand U2400 (N_2400,N_2299,N_2220);
xor U2401 (N_2401,N_2095,N_1760);
nand U2402 (N_2402,N_1448,N_1294);
and U2403 (N_2403,N_2312,N_1851);
and U2404 (N_2404,N_1256,N_1346);
and U2405 (N_2405,N_1451,N_2208);
xor U2406 (N_2406,N_1633,N_1685);
nand U2407 (N_2407,N_2301,N_2025);
nor U2408 (N_2408,N_1690,N_1849);
or U2409 (N_2409,N_2257,N_1663);
or U2410 (N_2410,N_1489,N_1657);
or U2411 (N_2411,N_2329,N_1427);
or U2412 (N_2412,N_2189,N_1513);
or U2413 (N_2413,N_1988,N_1579);
xnor U2414 (N_2414,N_1970,N_1512);
nor U2415 (N_2415,N_1485,N_1818);
or U2416 (N_2416,N_1942,N_1321);
or U2417 (N_2417,N_1403,N_2170);
and U2418 (N_2418,N_1552,N_1302);
and U2419 (N_2419,N_1859,N_2196);
and U2420 (N_2420,N_1777,N_2260);
nor U2421 (N_2421,N_2010,N_1536);
nand U2422 (N_2422,N_1282,N_1644);
nor U2423 (N_2423,N_1244,N_1484);
or U2424 (N_2424,N_2123,N_2294);
nor U2425 (N_2425,N_1532,N_1406);
and U2426 (N_2426,N_2380,N_1903);
or U2427 (N_2427,N_1698,N_1259);
and U2428 (N_2428,N_1637,N_1430);
xor U2429 (N_2429,N_2079,N_1695);
nor U2430 (N_2430,N_1857,N_1841);
xnor U2431 (N_2431,N_2321,N_2387);
nand U2432 (N_2432,N_1213,N_1531);
or U2433 (N_2433,N_2336,N_1215);
and U2434 (N_2434,N_2323,N_2143);
nor U2435 (N_2435,N_2087,N_1589);
or U2436 (N_2436,N_1959,N_1895);
or U2437 (N_2437,N_2050,N_1993);
nand U2438 (N_2438,N_1207,N_1928);
or U2439 (N_2439,N_2287,N_2304);
nor U2440 (N_2440,N_1673,N_1968);
nand U2441 (N_2441,N_1904,N_1470);
nand U2442 (N_2442,N_1697,N_2221);
and U2443 (N_2443,N_1774,N_2113);
nand U2444 (N_2444,N_1208,N_2376);
nand U2445 (N_2445,N_2334,N_2177);
or U2446 (N_2446,N_1630,N_1655);
and U2447 (N_2447,N_1803,N_2291);
nand U2448 (N_2448,N_2204,N_1212);
nor U2449 (N_2449,N_1844,N_1845);
and U2450 (N_2450,N_2031,N_2057);
nand U2451 (N_2451,N_1323,N_2328);
xor U2452 (N_2452,N_1709,N_2111);
and U2453 (N_2453,N_2256,N_1548);
xor U2454 (N_2454,N_1705,N_1924);
and U2455 (N_2455,N_2053,N_1665);
nor U2456 (N_2456,N_2049,N_1370);
or U2457 (N_2457,N_1814,N_2001);
nand U2458 (N_2458,N_1361,N_1574);
xor U2459 (N_2459,N_2349,N_1347);
and U2460 (N_2460,N_1925,N_1262);
nand U2461 (N_2461,N_1396,N_2385);
and U2462 (N_2462,N_2180,N_1964);
xor U2463 (N_2463,N_1413,N_2035);
and U2464 (N_2464,N_1433,N_2076);
nand U2465 (N_2465,N_1234,N_1599);
nor U2466 (N_2466,N_2185,N_1375);
nor U2467 (N_2467,N_1758,N_2373);
or U2468 (N_2468,N_1704,N_2018);
or U2469 (N_2469,N_2141,N_2102);
or U2470 (N_2470,N_1965,N_1738);
nor U2471 (N_2471,N_2078,N_1303);
nand U2472 (N_2472,N_1488,N_1566);
nor U2473 (N_2473,N_1251,N_1807);
and U2474 (N_2474,N_1722,N_1986);
xor U2475 (N_2475,N_2274,N_1821);
or U2476 (N_2476,N_1671,N_1969);
or U2477 (N_2477,N_1737,N_2259);
nor U2478 (N_2478,N_1486,N_2290);
xnor U2479 (N_2479,N_1525,N_1809);
nor U2480 (N_2480,N_1874,N_2152);
or U2481 (N_2481,N_1624,N_2393);
and U2482 (N_2482,N_1373,N_1463);
xor U2483 (N_2483,N_1983,N_2390);
nor U2484 (N_2484,N_1931,N_1628);
or U2485 (N_2485,N_1992,N_1352);
or U2486 (N_2486,N_2003,N_1640);
xor U2487 (N_2487,N_2162,N_2014);
and U2488 (N_2488,N_1483,N_1977);
or U2489 (N_2489,N_2222,N_1940);
nand U2490 (N_2490,N_1668,N_1391);
nor U2491 (N_2491,N_1712,N_1586);
and U2492 (N_2492,N_1257,N_1409);
nor U2493 (N_2493,N_1538,N_1639);
or U2494 (N_2494,N_1242,N_1870);
or U2495 (N_2495,N_1223,N_1847);
nor U2496 (N_2496,N_1674,N_1675);
nor U2497 (N_2497,N_1820,N_2369);
nor U2498 (N_2498,N_1260,N_2013);
or U2499 (N_2499,N_1500,N_1756);
or U2500 (N_2500,N_2121,N_1692);
nor U2501 (N_2501,N_1998,N_2354);
nand U2502 (N_2502,N_1881,N_1832);
nand U2503 (N_2503,N_1336,N_1591);
nand U2504 (N_2504,N_1434,N_2075);
nand U2505 (N_2505,N_2335,N_2302);
nor U2506 (N_2506,N_1775,N_2339);
or U2507 (N_2507,N_2131,N_1752);
or U2508 (N_2508,N_1919,N_2364);
or U2509 (N_2509,N_2273,N_1353);
xor U2510 (N_2510,N_1779,N_2359);
nand U2511 (N_2511,N_1985,N_1827);
xor U2512 (N_2512,N_1476,N_2231);
and U2513 (N_2513,N_2343,N_2205);
xnor U2514 (N_2514,N_1474,N_1773);
nor U2515 (N_2515,N_1647,N_2389);
xnor U2516 (N_2516,N_1506,N_1499);
xnor U2517 (N_2517,N_1748,N_2316);
nand U2518 (N_2518,N_1581,N_1437);
or U2519 (N_2519,N_2397,N_1417);
nor U2520 (N_2520,N_2080,N_2388);
xor U2521 (N_2521,N_2247,N_2324);
nand U2522 (N_2522,N_2178,N_2396);
and U2523 (N_2523,N_2155,N_1364);
and U2524 (N_2524,N_2101,N_1585);
nor U2525 (N_2525,N_1801,N_2174);
xor U2526 (N_2526,N_1562,N_1740);
and U2527 (N_2527,N_2238,N_1263);
nand U2528 (N_2528,N_1862,N_2167);
or U2529 (N_2529,N_1984,N_1209);
nand U2530 (N_2530,N_1226,N_1508);
or U2531 (N_2531,N_2214,N_1271);
or U2532 (N_2532,N_2097,N_2129);
nand U2533 (N_2533,N_1309,N_1570);
or U2534 (N_2534,N_2068,N_2094);
or U2535 (N_2535,N_1299,N_2194);
and U2536 (N_2536,N_1629,N_1460);
nand U2537 (N_2537,N_1443,N_2156);
xnor U2538 (N_2538,N_1472,N_2024);
nand U2539 (N_2539,N_1785,N_2346);
and U2540 (N_2540,N_1292,N_1727);
nand U2541 (N_2541,N_1613,N_2252);
nor U2542 (N_2542,N_1677,N_1627);
and U2543 (N_2543,N_1455,N_1333);
or U2544 (N_2544,N_1478,N_1368);
xor U2545 (N_2545,N_1381,N_1468);
xnor U2546 (N_2546,N_2292,N_1219);
nand U2547 (N_2547,N_2073,N_1349);
or U2548 (N_2548,N_1252,N_1838);
nor U2549 (N_2549,N_1345,N_1363);
nor U2550 (N_2550,N_1782,N_1441);
nor U2551 (N_2551,N_1432,N_1929);
or U2552 (N_2552,N_2008,N_2392);
nand U2553 (N_2553,N_1431,N_1355);
and U2554 (N_2554,N_1461,N_2303);
nand U2555 (N_2555,N_1576,N_1643);
and U2556 (N_2556,N_1887,N_1405);
nand U2557 (N_2557,N_1715,N_1702);
and U2558 (N_2558,N_1781,N_2117);
and U2559 (N_2559,N_1314,N_1313);
or U2560 (N_2560,N_1535,N_1201);
and U2561 (N_2561,N_1392,N_1635);
nor U2562 (N_2562,N_1235,N_1923);
nand U2563 (N_2563,N_1603,N_1795);
and U2564 (N_2564,N_1742,N_2348);
nor U2565 (N_2565,N_1595,N_1955);
xnor U2566 (N_2566,N_2148,N_2203);
or U2567 (N_2567,N_1240,N_1274);
nand U2568 (N_2568,N_2071,N_1686);
or U2569 (N_2569,N_1997,N_1854);
and U2570 (N_2570,N_1232,N_2004);
nand U2571 (N_2571,N_1654,N_2210);
nor U2572 (N_2572,N_2229,N_2042);
xor U2573 (N_2573,N_1735,N_2037);
or U2574 (N_2574,N_1961,N_2358);
and U2575 (N_2575,N_1202,N_1516);
xnor U2576 (N_2576,N_1407,N_2319);
nor U2577 (N_2577,N_1253,N_1337);
and U2578 (N_2578,N_1596,N_2352);
and U2579 (N_2579,N_2060,N_2065);
xor U2580 (N_2580,N_2258,N_2000);
xnor U2581 (N_2581,N_1941,N_1217);
nand U2582 (N_2582,N_2310,N_1944);
and U2583 (N_2583,N_1880,N_1906);
and U2584 (N_2584,N_1708,N_2158);
nor U2585 (N_2585,N_1926,N_1469);
nor U2586 (N_2586,N_1289,N_2093);
and U2587 (N_2587,N_2173,N_2026);
xnor U2588 (N_2588,N_1823,N_1759);
and U2589 (N_2589,N_1527,N_1878);
or U2590 (N_2590,N_2127,N_1645);
xnor U2591 (N_2591,N_1334,N_1605);
and U2592 (N_2592,N_2384,N_1855);
or U2593 (N_2593,N_1688,N_2293);
xor U2594 (N_2594,N_1689,N_1534);
xor U2595 (N_2595,N_1399,N_2240);
xnor U2596 (N_2596,N_2379,N_1385);
xor U2597 (N_2597,N_1730,N_1575);
xor U2598 (N_2598,N_1281,N_1388);
and U2599 (N_2599,N_1568,N_1320);
or U2600 (N_2600,N_2020,N_2032);
or U2601 (N_2601,N_1864,N_1280);
nand U2602 (N_2602,N_1962,N_1357);
nand U2603 (N_2603,N_1684,N_1691);
nand U2604 (N_2604,N_1794,N_1636);
xnor U2605 (N_2605,N_1249,N_1721);
or U2606 (N_2606,N_2046,N_1806);
nor U2607 (N_2607,N_2126,N_1446);
nand U2608 (N_2608,N_1598,N_1293);
or U2609 (N_2609,N_1703,N_1418);
xor U2610 (N_2610,N_2153,N_1651);
nor U2611 (N_2611,N_1245,N_1416);
nand U2612 (N_2612,N_1236,N_1800);
or U2613 (N_2613,N_2040,N_1482);
and U2614 (N_2614,N_1543,N_2184);
nand U2615 (N_2615,N_1679,N_1400);
nand U2616 (N_2616,N_1764,N_1848);
xnor U2617 (N_2617,N_1401,N_1393);
nor U2618 (N_2618,N_1344,N_1846);
xnor U2619 (N_2619,N_1348,N_2186);
nand U2620 (N_2620,N_2367,N_1772);
and U2621 (N_2621,N_2043,N_1545);
nand U2622 (N_2622,N_2146,N_2070);
nand U2623 (N_2623,N_2241,N_2021);
and U2624 (N_2624,N_1739,N_2253);
and U2625 (N_2625,N_1815,N_2382);
and U2626 (N_2626,N_1780,N_2331);
or U2627 (N_2627,N_1338,N_1277);
and U2628 (N_2628,N_1354,N_2016);
or U2629 (N_2629,N_1826,N_2201);
and U2630 (N_2630,N_2326,N_1790);
and U2631 (N_2631,N_2019,N_1793);
nand U2632 (N_2632,N_1971,N_1222);
and U2633 (N_2633,N_2022,N_1475);
nand U2634 (N_2634,N_2395,N_1350);
xnor U2635 (N_2635,N_2098,N_1852);
xor U2636 (N_2636,N_1641,N_1544);
or U2637 (N_2637,N_1533,N_1560);
nand U2638 (N_2638,N_2118,N_2107);
nor U2639 (N_2639,N_1593,N_2219);
nand U2640 (N_2640,N_1957,N_1725);
nor U2641 (N_2641,N_1699,N_2104);
or U2642 (N_2642,N_1853,N_2181);
xnor U2643 (N_2643,N_2267,N_2134);
xor U2644 (N_2644,N_2317,N_2378);
xor U2645 (N_2645,N_2047,N_1952);
xnor U2646 (N_2646,N_1776,N_1732);
xor U2647 (N_2647,N_1731,N_1830);
and U2648 (N_2648,N_1204,N_1408);
or U2649 (N_2649,N_1948,N_1746);
nor U2650 (N_2650,N_1558,N_1376);
nor U2651 (N_2651,N_1652,N_2182);
or U2652 (N_2652,N_2172,N_2213);
xor U2653 (N_2653,N_2216,N_1250);
nor U2654 (N_2654,N_1541,N_2171);
xnor U2655 (N_2655,N_1642,N_2038);
nor U2656 (N_2656,N_1729,N_1224);
or U2657 (N_2657,N_1519,N_1907);
and U2658 (N_2658,N_1255,N_2226);
xnor U2659 (N_2659,N_1565,N_1723);
nand U2660 (N_2660,N_2135,N_1920);
and U2661 (N_2661,N_1398,N_1411);
xor U2662 (N_2662,N_1680,N_2375);
nor U2663 (N_2663,N_1386,N_1933);
nand U2664 (N_2664,N_2305,N_1741);
xor U2665 (N_2665,N_2307,N_2136);
and U2666 (N_2666,N_1656,N_1956);
and U2667 (N_2667,N_1310,N_1395);
nand U2668 (N_2668,N_1382,N_1367);
and U2669 (N_2669,N_2313,N_1233);
nand U2670 (N_2670,N_1205,N_1745);
nor U2671 (N_2671,N_1587,N_2041);
or U2672 (N_2672,N_1511,N_1380);
nand U2673 (N_2673,N_2157,N_1218);
xor U2674 (N_2674,N_2325,N_1927);
nor U2675 (N_2675,N_2202,N_1750);
or U2676 (N_2676,N_1318,N_1267);
xor U2677 (N_2677,N_1521,N_2399);
or U2678 (N_2678,N_2309,N_2059);
and U2679 (N_2679,N_2054,N_1799);
nand U2680 (N_2680,N_1297,N_1938);
and U2681 (N_2681,N_1912,N_1917);
xnor U2682 (N_2682,N_2218,N_1648);
or U2683 (N_2683,N_1307,N_2191);
or U2684 (N_2684,N_1632,N_1863);
nand U2685 (N_2685,N_2361,N_1991);
nand U2686 (N_2686,N_1664,N_2066);
nor U2687 (N_2687,N_1770,N_2144);
and U2688 (N_2688,N_2193,N_2027);
xor U2689 (N_2689,N_1840,N_1808);
and U2690 (N_2690,N_2233,N_1888);
nand U2691 (N_2691,N_2183,N_2282);
and U2692 (N_2692,N_1530,N_1425);
nor U2693 (N_2693,N_2289,N_2278);
nand U2694 (N_2694,N_1296,N_2298);
xnor U2695 (N_2695,N_2391,N_1362);
or U2696 (N_2696,N_2009,N_2138);
nand U2697 (N_2697,N_1372,N_1214);
nand U2698 (N_2698,N_2333,N_1711);
nand U2699 (N_2699,N_1378,N_1701);
nand U2700 (N_2700,N_1834,N_1584);
and U2701 (N_2701,N_2264,N_1428);
or U2702 (N_2702,N_2083,N_1442);
or U2703 (N_2703,N_2002,N_1424);
xor U2704 (N_2704,N_1877,N_1900);
xnor U2705 (N_2705,N_1556,N_1916);
xor U2706 (N_2706,N_1377,N_1649);
xnor U2707 (N_2707,N_1551,N_1200);
xor U2708 (N_2708,N_2088,N_1466);
xor U2709 (N_2709,N_2356,N_1891);
and U2710 (N_2710,N_2074,N_1762);
xnor U2711 (N_2711,N_2338,N_1285);
nor U2712 (N_2712,N_1369,N_1546);
or U2713 (N_2713,N_1898,N_1528);
nor U2714 (N_2714,N_1327,N_1829);
and U2715 (N_2715,N_2197,N_1618);
nand U2716 (N_2716,N_1414,N_2245);
nor U2717 (N_2717,N_2199,N_1600);
xor U2718 (N_2718,N_1659,N_2058);
xor U2719 (N_2719,N_1620,N_1272);
nand U2720 (N_2720,N_1753,N_2314);
xnor U2721 (N_2721,N_1526,N_1331);
xor U2722 (N_2722,N_1899,N_1203);
xnor U2723 (N_2723,N_1206,N_1974);
nand U2724 (N_2724,N_1945,N_1819);
and U2725 (N_2725,N_1445,N_2090);
nand U2726 (N_2726,N_1561,N_1305);
nand U2727 (N_2727,N_1812,N_1835);
or U2728 (N_2728,N_1265,N_2320);
or U2729 (N_2729,N_1578,N_1456);
or U2730 (N_2730,N_1871,N_1831);
and U2731 (N_2731,N_1426,N_2342);
nand U2732 (N_2732,N_1902,N_2232);
nand U2733 (N_2733,N_2377,N_2268);
nor U2734 (N_2734,N_1588,N_1876);
nor U2735 (N_2735,N_1311,N_2159);
and U2736 (N_2736,N_2340,N_1477);
or U2737 (N_2737,N_2085,N_1850);
and U2738 (N_2738,N_1278,N_1622);
or U2739 (N_2739,N_1670,N_2366);
xor U2740 (N_2740,N_1230,N_1554);
nor U2741 (N_2741,N_1867,N_1550);
or U2742 (N_2742,N_1910,N_1279);
xor U2743 (N_2743,N_1619,N_2266);
or U2744 (N_2744,N_1473,N_2362);
and U2745 (N_2745,N_2261,N_1341);
nand U2746 (N_2746,N_1608,N_2106);
nand U2747 (N_2747,N_2212,N_1423);
nand U2748 (N_2748,N_1617,N_1733);
xnor U2749 (N_2749,N_2308,N_1946);
nand U2750 (N_2750,N_1861,N_1567);
and U2751 (N_2751,N_1342,N_1439);
and U2752 (N_2752,N_1537,N_1322);
xor U2753 (N_2753,N_2363,N_1435);
or U2754 (N_2754,N_1238,N_1389);
and U2755 (N_2755,N_1967,N_1868);
nand U2756 (N_2756,N_1975,N_1514);
nor U2757 (N_2757,N_2089,N_2033);
nor U2758 (N_2758,N_2350,N_1356);
or U2759 (N_2759,N_1319,N_1743);
and U2760 (N_2760,N_1247,N_1761);
nor U2761 (N_2761,N_1607,N_2322);
nor U2762 (N_2762,N_2275,N_2341);
nand U2763 (N_2763,N_1996,N_2011);
nand U2764 (N_2764,N_1231,N_1429);
and U2765 (N_2765,N_2006,N_2300);
nand U2766 (N_2766,N_1707,N_1493);
nor U2767 (N_2767,N_1481,N_2355);
or U2768 (N_2768,N_1394,N_1749);
or U2769 (N_2769,N_1797,N_1947);
or U2770 (N_2770,N_1710,N_1787);
and U2771 (N_2771,N_2139,N_2372);
xor U2772 (N_2772,N_1609,N_1555);
nor U2773 (N_2773,N_2142,N_1918);
nor U2774 (N_2774,N_1496,N_1713);
nand U2775 (N_2775,N_2255,N_1865);
and U2776 (N_2776,N_1275,N_2108);
nand U2777 (N_2777,N_1783,N_2034);
and U2778 (N_2778,N_1879,N_1572);
xor U2779 (N_2779,N_2224,N_1883);
and U2780 (N_2780,N_2077,N_2056);
nand U2781 (N_2781,N_2069,N_1495);
and U2782 (N_2782,N_1842,N_1872);
xnor U2783 (N_2783,N_1497,N_1653);
xor U2784 (N_2784,N_1540,N_1509);
xnor U2785 (N_2785,N_2029,N_1935);
or U2786 (N_2786,N_2250,N_1374);
nor U2787 (N_2787,N_1683,N_2383);
nor U2788 (N_2788,N_2165,N_1706);
and U2789 (N_2789,N_2288,N_1681);
or U2790 (N_2790,N_1505,N_1804);
or U2791 (N_2791,N_1365,N_2311);
nand U2792 (N_2792,N_2092,N_1360);
or U2793 (N_2793,N_1896,N_1366);
nand U2794 (N_2794,N_1911,N_1634);
xor U2795 (N_2795,N_2284,N_2195);
and U2796 (N_2796,N_1306,N_1590);
or U2797 (N_2797,N_1471,N_2271);
nor U2798 (N_2798,N_2045,N_1958);
nor U2799 (N_2799,N_1577,N_2176);
nor U2800 (N_2800,N_1592,N_1606);
and U2801 (N_2801,N_1615,N_2154);
nor U2802 (N_2802,N_1805,N_1553);
and U2803 (N_2803,N_1465,N_2179);
or U2804 (N_2804,N_2242,N_1908);
or U2805 (N_2805,N_1248,N_1228);
nand U2806 (N_2806,N_2140,N_1410);
xnor U2807 (N_2807,N_1751,N_2332);
and U2808 (N_2808,N_1905,N_1700);
xor U2809 (N_2809,N_2200,N_2270);
and U2810 (N_2810,N_1922,N_1682);
nor U2811 (N_2811,N_1616,N_2286);
or U2812 (N_2812,N_1980,N_1501);
nand U2813 (N_2813,N_1494,N_1676);
or U2814 (N_2814,N_2160,N_1457);
xor U2815 (N_2815,N_2132,N_1464);
or U2816 (N_2816,N_2281,N_2244);
xor U2817 (N_2817,N_2130,N_1583);
or U2818 (N_2818,N_1315,N_2217);
nand U2819 (N_2819,N_1332,N_1765);
nor U2820 (N_2820,N_1978,N_2161);
or U2821 (N_2821,N_2265,N_1239);
nor U2822 (N_2822,N_1884,N_1650);
or U2823 (N_2823,N_2109,N_1754);
or U2824 (N_2824,N_2122,N_2081);
nand U2825 (N_2825,N_1454,N_1221);
and U2826 (N_2826,N_2052,N_1325);
nor U2827 (N_2827,N_1778,N_1359);
or U2828 (N_2828,N_1211,N_1440);
nor U2829 (N_2829,N_1943,N_2064);
and U2830 (N_2830,N_1734,N_2169);
or U2831 (N_2831,N_2133,N_2055);
xor U2832 (N_2832,N_1547,N_1422);
nor U2833 (N_2833,N_2234,N_1989);
and U2834 (N_2834,N_1421,N_1972);
or U2835 (N_2835,N_1510,N_1963);
nor U2836 (N_2836,N_1953,N_1914);
or U2837 (N_2837,N_1273,N_1825);
xor U2838 (N_2838,N_2099,N_2353);
nand U2839 (N_2839,N_1890,N_1934);
xor U2840 (N_2840,N_1573,N_2237);
nor U2841 (N_2841,N_2091,N_1726);
xnor U2842 (N_2842,N_2103,N_1316);
xor U2843 (N_2843,N_1932,N_2295);
and U2844 (N_2844,N_1412,N_1611);
nand U2845 (N_2845,N_2039,N_1792);
xnor U2846 (N_2846,N_2283,N_1458);
and U2847 (N_2847,N_2345,N_1771);
or U2848 (N_2848,N_1667,N_1504);
and U2849 (N_2849,N_1270,N_1889);
xor U2850 (N_2850,N_1351,N_1909);
and U2851 (N_2851,N_2067,N_2017);
and U2852 (N_2852,N_2227,N_2072);
and U2853 (N_2853,N_2084,N_2368);
nor U2854 (N_2854,N_1873,N_1339);
or U2855 (N_2855,N_1419,N_1981);
nor U2856 (N_2856,N_1802,N_1921);
nor U2857 (N_2857,N_2236,N_1288);
nor U2858 (N_2858,N_2347,N_1658);
and U2859 (N_2859,N_1987,N_2168);
nor U2860 (N_2860,N_1340,N_1716);
or U2861 (N_2861,N_1843,N_2166);
or U2862 (N_2862,N_2086,N_1858);
xnor U2863 (N_2863,N_1300,N_1875);
or U2864 (N_2864,N_2188,N_2228);
xor U2865 (N_2865,N_1856,N_1995);
nand U2866 (N_2866,N_1717,N_2149);
and U2867 (N_2867,N_1893,N_1860);
nor U2868 (N_2868,N_1326,N_1747);
xnor U2869 (N_2869,N_1766,N_2351);
and U2870 (N_2870,N_1523,N_2285);
and U2871 (N_2871,N_1237,N_1696);
and U2872 (N_2872,N_1714,N_1438);
and U2873 (N_2873,N_1520,N_1243);
and U2874 (N_2874,N_1930,N_1791);
and U2875 (N_2875,N_1882,N_2344);
nor U2876 (N_2876,N_1950,N_1811);
or U2877 (N_2877,N_1724,N_1261);
xor U2878 (N_2878,N_1559,N_1447);
nor U2879 (N_2879,N_1216,N_2137);
and U2880 (N_2880,N_2296,N_1660);
xor U2881 (N_2881,N_2036,N_1324);
nand U2882 (N_2882,N_2230,N_2119);
and U2883 (N_2883,N_1415,N_1982);
xor U2884 (N_2884,N_1915,N_1789);
nand U2885 (N_2885,N_2272,N_2012);
and U2886 (N_2886,N_1502,N_1669);
and U2887 (N_2887,N_1491,N_1295);
and U2888 (N_2888,N_1736,N_1828);
or U2889 (N_2889,N_2327,N_2215);
and U2890 (N_2890,N_2048,N_1227);
nor U2891 (N_2891,N_1913,N_1768);
and U2892 (N_2892,N_1264,N_1824);
or U2893 (N_2893,N_1444,N_1678);
nand U2894 (N_2894,N_1604,N_1755);
xor U2895 (N_2895,N_2023,N_2128);
and U2896 (N_2896,N_1594,N_1796);
nand U2897 (N_2897,N_2223,N_1631);
xnor U2898 (N_2898,N_2192,N_1390);
nor U2899 (N_2899,N_1949,N_1693);
or U2900 (N_2900,N_1241,N_1718);
xnor U2901 (N_2901,N_1503,N_2357);
or U2902 (N_2902,N_1480,N_2263);
xnor U2903 (N_2903,N_2209,N_2280);
nor U2904 (N_2904,N_1258,N_1597);
nand U2905 (N_2905,N_1966,N_1268);
xnor U2906 (N_2906,N_1479,N_1973);
xor U2907 (N_2907,N_1625,N_1459);
or U2908 (N_2908,N_2246,N_2164);
nor U2909 (N_2909,N_2243,N_2370);
or U2910 (N_2910,N_1788,N_2318);
xnor U2911 (N_2911,N_1763,N_1330);
nand U2912 (N_2912,N_1767,N_1582);
xnor U2913 (N_2913,N_2251,N_2330);
and U2914 (N_2914,N_1524,N_1990);
and U2915 (N_2915,N_1539,N_1312);
and U2916 (N_2916,N_1936,N_1436);
nand U2917 (N_2917,N_2297,N_1467);
xnor U2918 (N_2918,N_1661,N_1646);
and U2919 (N_2919,N_2105,N_1564);
nand U2920 (N_2920,N_1254,N_2386);
or U2921 (N_2921,N_1979,N_2114);
xor U2922 (N_2922,N_2239,N_1894);
or U2923 (N_2923,N_2120,N_1301);
and U2924 (N_2924,N_1329,N_2028);
and U2925 (N_2925,N_1951,N_1220);
and U2926 (N_2926,N_1798,N_1308);
nand U2927 (N_2927,N_1328,N_1549);
xor U2928 (N_2928,N_1286,N_1210);
nor U2929 (N_2929,N_1225,N_1976);
xnor U2930 (N_2930,N_1450,N_2211);
and U2931 (N_2931,N_1358,N_1839);
nand U2932 (N_2932,N_1420,N_2206);
nand U2933 (N_2933,N_2381,N_1744);
or U2934 (N_2934,N_1994,N_2262);
nor U2935 (N_2935,N_1786,N_1886);
and U2936 (N_2936,N_1518,N_1269);
nor U2937 (N_2937,N_1557,N_1284);
or U2938 (N_2938,N_1379,N_1728);
nor U2939 (N_2939,N_1623,N_2277);
xnor U2940 (N_2940,N_2163,N_1885);
nor U2941 (N_2941,N_2100,N_1769);
or U2942 (N_2942,N_1335,N_1626);
nor U2943 (N_2943,N_1939,N_2279);
xor U2944 (N_2944,N_2082,N_1229);
xor U2945 (N_2945,N_1387,N_1869);
xnor U2946 (N_2946,N_2175,N_1901);
nor U2947 (N_2947,N_2315,N_1492);
nor U2948 (N_2948,N_1638,N_1960);
or U2949 (N_2949,N_2051,N_1816);
nand U2950 (N_2950,N_1866,N_2096);
nand U2951 (N_2951,N_2371,N_1621);
xor U2952 (N_2952,N_1614,N_1601);
xnor U2953 (N_2953,N_2063,N_1563);
nor U2954 (N_2954,N_2030,N_2115);
or U2955 (N_2955,N_1542,N_2007);
nand U2956 (N_2956,N_2269,N_1999);
xnor U2957 (N_2957,N_1298,N_2337);
and U2958 (N_2958,N_1580,N_2225);
xor U2959 (N_2959,N_2147,N_1515);
and U2960 (N_2960,N_2394,N_1836);
and U2961 (N_2961,N_1612,N_1937);
xnor U2962 (N_2962,N_2062,N_1837);
and U2963 (N_2963,N_2150,N_1813);
xor U2964 (N_2964,N_2110,N_1757);
xnor U2965 (N_2965,N_1666,N_1462);
nand U2966 (N_2966,N_1687,N_2151);
nand U2967 (N_2967,N_2248,N_1276);
nor U2968 (N_2968,N_2190,N_1384);
or U2969 (N_2969,N_2276,N_1522);
nor U2970 (N_2970,N_2116,N_1571);
xor U2971 (N_2971,N_1897,N_1343);
nand U2972 (N_2972,N_1507,N_1719);
nand U2973 (N_2973,N_1810,N_1291);
or U2974 (N_2974,N_2306,N_1402);
nand U2975 (N_2975,N_2124,N_2044);
nor U2976 (N_2976,N_1672,N_2005);
and U2977 (N_2977,N_1602,N_1833);
xnor U2978 (N_2978,N_1954,N_1304);
and U2979 (N_2979,N_2145,N_2374);
xor U2980 (N_2980,N_1517,N_1371);
nand U2981 (N_2981,N_1498,N_1610);
nand U2982 (N_2982,N_1246,N_1290);
nor U2983 (N_2983,N_1383,N_1452);
and U2984 (N_2984,N_1720,N_2125);
or U2985 (N_2985,N_1283,N_2015);
xor U2986 (N_2986,N_1287,N_2112);
xnor U2987 (N_2987,N_1892,N_1569);
nand U2988 (N_2988,N_1662,N_1449);
nor U2989 (N_2989,N_1266,N_2249);
xor U2990 (N_2990,N_1490,N_1784);
and U2991 (N_2991,N_1397,N_1404);
and U2992 (N_2992,N_1694,N_2365);
and U2993 (N_2993,N_1822,N_1453);
or U2994 (N_2994,N_1529,N_2235);
xor U2995 (N_2995,N_1487,N_2061);
and U2996 (N_2996,N_2398,N_2207);
nand U2997 (N_2997,N_2187,N_1817);
nand U2998 (N_2998,N_1317,N_2254);
xor U2999 (N_2999,N_2198,N_2360);
nand U3000 (N_3000,N_1852,N_1951);
nor U3001 (N_3001,N_1755,N_2282);
or U3002 (N_3002,N_2271,N_1600);
xnor U3003 (N_3003,N_1861,N_1473);
or U3004 (N_3004,N_1437,N_1308);
xnor U3005 (N_3005,N_1360,N_1381);
nand U3006 (N_3006,N_1260,N_1978);
or U3007 (N_3007,N_1529,N_1907);
xnor U3008 (N_3008,N_1723,N_1868);
or U3009 (N_3009,N_1605,N_2072);
xnor U3010 (N_3010,N_1394,N_1527);
nand U3011 (N_3011,N_1624,N_1843);
nand U3012 (N_3012,N_2340,N_2330);
and U3013 (N_3013,N_1510,N_2292);
or U3014 (N_3014,N_2258,N_1438);
or U3015 (N_3015,N_2278,N_1970);
xor U3016 (N_3016,N_1717,N_1872);
xor U3017 (N_3017,N_2206,N_1209);
and U3018 (N_3018,N_2032,N_1432);
nand U3019 (N_3019,N_2345,N_1690);
nand U3020 (N_3020,N_2114,N_1323);
nor U3021 (N_3021,N_2034,N_2107);
xor U3022 (N_3022,N_1734,N_1301);
or U3023 (N_3023,N_2368,N_2130);
and U3024 (N_3024,N_1709,N_1874);
and U3025 (N_3025,N_1790,N_1965);
xor U3026 (N_3026,N_1470,N_1566);
xor U3027 (N_3027,N_2310,N_2165);
or U3028 (N_3028,N_2269,N_2111);
and U3029 (N_3029,N_2222,N_1210);
xnor U3030 (N_3030,N_2093,N_2006);
and U3031 (N_3031,N_1400,N_1273);
xor U3032 (N_3032,N_1243,N_1283);
nor U3033 (N_3033,N_1377,N_2205);
nor U3034 (N_3034,N_2150,N_1739);
and U3035 (N_3035,N_2334,N_1940);
xor U3036 (N_3036,N_1680,N_1317);
nor U3037 (N_3037,N_2330,N_2378);
nand U3038 (N_3038,N_2059,N_1236);
nand U3039 (N_3039,N_2393,N_1996);
xor U3040 (N_3040,N_1650,N_1277);
or U3041 (N_3041,N_1518,N_1405);
nor U3042 (N_3042,N_1932,N_1994);
nor U3043 (N_3043,N_1349,N_1332);
nor U3044 (N_3044,N_1513,N_2343);
and U3045 (N_3045,N_2181,N_1711);
and U3046 (N_3046,N_1228,N_1361);
or U3047 (N_3047,N_1278,N_1753);
or U3048 (N_3048,N_2054,N_2308);
nand U3049 (N_3049,N_1617,N_1711);
and U3050 (N_3050,N_1240,N_1384);
or U3051 (N_3051,N_1716,N_1843);
or U3052 (N_3052,N_1749,N_2117);
or U3053 (N_3053,N_2298,N_1521);
nand U3054 (N_3054,N_2215,N_1334);
or U3055 (N_3055,N_2106,N_2249);
xor U3056 (N_3056,N_1271,N_1738);
and U3057 (N_3057,N_1817,N_1652);
xor U3058 (N_3058,N_1765,N_2337);
nand U3059 (N_3059,N_1477,N_1375);
nand U3060 (N_3060,N_1776,N_1673);
or U3061 (N_3061,N_2043,N_1788);
and U3062 (N_3062,N_1944,N_1774);
nor U3063 (N_3063,N_1924,N_1895);
xor U3064 (N_3064,N_2225,N_1466);
nand U3065 (N_3065,N_1358,N_1986);
or U3066 (N_3066,N_1200,N_1530);
xnor U3067 (N_3067,N_1538,N_1467);
nor U3068 (N_3068,N_1953,N_1599);
nand U3069 (N_3069,N_1370,N_2209);
nor U3070 (N_3070,N_1251,N_1494);
or U3071 (N_3071,N_1478,N_1805);
nand U3072 (N_3072,N_1793,N_1511);
nor U3073 (N_3073,N_1299,N_2033);
and U3074 (N_3074,N_1357,N_1977);
or U3075 (N_3075,N_1738,N_1315);
xnor U3076 (N_3076,N_1479,N_2140);
nor U3077 (N_3077,N_1888,N_1526);
and U3078 (N_3078,N_1931,N_1812);
xnor U3079 (N_3079,N_1578,N_1674);
xnor U3080 (N_3080,N_2190,N_2287);
nand U3081 (N_3081,N_1909,N_1616);
or U3082 (N_3082,N_1752,N_2341);
and U3083 (N_3083,N_1326,N_2023);
and U3084 (N_3084,N_1302,N_2393);
and U3085 (N_3085,N_1316,N_1555);
nor U3086 (N_3086,N_2009,N_1807);
xor U3087 (N_3087,N_2276,N_1495);
nand U3088 (N_3088,N_2394,N_2177);
and U3089 (N_3089,N_2373,N_1248);
nand U3090 (N_3090,N_1254,N_2221);
xnor U3091 (N_3091,N_2363,N_2288);
nand U3092 (N_3092,N_1854,N_1332);
xnor U3093 (N_3093,N_2240,N_1356);
or U3094 (N_3094,N_1619,N_1622);
xor U3095 (N_3095,N_1766,N_1219);
and U3096 (N_3096,N_1463,N_1507);
xnor U3097 (N_3097,N_2336,N_2198);
or U3098 (N_3098,N_2076,N_1492);
xnor U3099 (N_3099,N_1736,N_1481);
nor U3100 (N_3100,N_2163,N_1575);
and U3101 (N_3101,N_2172,N_2359);
nor U3102 (N_3102,N_2346,N_1964);
nand U3103 (N_3103,N_1911,N_1307);
nor U3104 (N_3104,N_1961,N_2131);
nand U3105 (N_3105,N_1396,N_2022);
or U3106 (N_3106,N_2389,N_1949);
xor U3107 (N_3107,N_1243,N_2055);
and U3108 (N_3108,N_1698,N_1755);
and U3109 (N_3109,N_1776,N_2234);
nor U3110 (N_3110,N_1715,N_2184);
nand U3111 (N_3111,N_1543,N_1456);
and U3112 (N_3112,N_2036,N_1360);
nand U3113 (N_3113,N_1831,N_1245);
nand U3114 (N_3114,N_2226,N_1345);
and U3115 (N_3115,N_1894,N_2360);
nand U3116 (N_3116,N_1790,N_1700);
nor U3117 (N_3117,N_1221,N_2106);
nor U3118 (N_3118,N_1576,N_1435);
and U3119 (N_3119,N_1612,N_1708);
xnor U3120 (N_3120,N_1755,N_1217);
nor U3121 (N_3121,N_1512,N_2294);
nor U3122 (N_3122,N_2286,N_1443);
and U3123 (N_3123,N_2171,N_1346);
nor U3124 (N_3124,N_1801,N_1797);
nor U3125 (N_3125,N_1486,N_2302);
nand U3126 (N_3126,N_2315,N_2238);
and U3127 (N_3127,N_2134,N_1725);
or U3128 (N_3128,N_1292,N_1885);
xor U3129 (N_3129,N_1417,N_1994);
or U3130 (N_3130,N_2222,N_1674);
nand U3131 (N_3131,N_1923,N_2283);
or U3132 (N_3132,N_2350,N_1796);
nand U3133 (N_3133,N_1287,N_2188);
nor U3134 (N_3134,N_2394,N_2032);
nor U3135 (N_3135,N_2373,N_1860);
nor U3136 (N_3136,N_2266,N_1311);
or U3137 (N_3137,N_2056,N_1920);
nand U3138 (N_3138,N_1294,N_1406);
nor U3139 (N_3139,N_2228,N_1735);
and U3140 (N_3140,N_1504,N_1465);
nand U3141 (N_3141,N_1625,N_1718);
xor U3142 (N_3142,N_1208,N_1315);
or U3143 (N_3143,N_2287,N_1716);
or U3144 (N_3144,N_1332,N_1601);
xnor U3145 (N_3145,N_1522,N_1839);
and U3146 (N_3146,N_1956,N_1215);
nor U3147 (N_3147,N_1712,N_1917);
or U3148 (N_3148,N_1748,N_2347);
or U3149 (N_3149,N_1259,N_2271);
or U3150 (N_3150,N_2089,N_1902);
xor U3151 (N_3151,N_1715,N_2136);
and U3152 (N_3152,N_2354,N_1320);
and U3153 (N_3153,N_1909,N_1621);
nor U3154 (N_3154,N_1672,N_1859);
nand U3155 (N_3155,N_1535,N_1841);
or U3156 (N_3156,N_1297,N_1339);
nand U3157 (N_3157,N_1778,N_2229);
nor U3158 (N_3158,N_2027,N_1347);
nand U3159 (N_3159,N_2160,N_2278);
xnor U3160 (N_3160,N_1997,N_1492);
xnor U3161 (N_3161,N_1333,N_2186);
nor U3162 (N_3162,N_1440,N_1325);
xor U3163 (N_3163,N_1583,N_1906);
nand U3164 (N_3164,N_1422,N_2064);
xor U3165 (N_3165,N_2365,N_2284);
nand U3166 (N_3166,N_2109,N_1305);
and U3167 (N_3167,N_2004,N_1494);
and U3168 (N_3168,N_1532,N_2052);
nor U3169 (N_3169,N_1324,N_2039);
nand U3170 (N_3170,N_2173,N_1221);
or U3171 (N_3171,N_1880,N_1603);
nand U3172 (N_3172,N_1207,N_1815);
or U3173 (N_3173,N_2060,N_1907);
nor U3174 (N_3174,N_1702,N_1478);
or U3175 (N_3175,N_1403,N_1422);
xor U3176 (N_3176,N_1755,N_1356);
xnor U3177 (N_3177,N_1678,N_1393);
xnor U3178 (N_3178,N_2281,N_2331);
and U3179 (N_3179,N_2168,N_1446);
nor U3180 (N_3180,N_1261,N_2010);
xor U3181 (N_3181,N_1920,N_1979);
and U3182 (N_3182,N_2139,N_1268);
or U3183 (N_3183,N_1940,N_1222);
nor U3184 (N_3184,N_2295,N_2115);
and U3185 (N_3185,N_1484,N_1457);
nor U3186 (N_3186,N_1975,N_1826);
nand U3187 (N_3187,N_1322,N_1305);
nand U3188 (N_3188,N_1348,N_1583);
xnor U3189 (N_3189,N_1862,N_1697);
or U3190 (N_3190,N_1502,N_2248);
nand U3191 (N_3191,N_1486,N_1268);
or U3192 (N_3192,N_1879,N_1815);
and U3193 (N_3193,N_1632,N_1596);
nor U3194 (N_3194,N_1358,N_1399);
or U3195 (N_3195,N_1987,N_2192);
and U3196 (N_3196,N_1369,N_2365);
or U3197 (N_3197,N_2194,N_1432);
nor U3198 (N_3198,N_2111,N_1219);
nand U3199 (N_3199,N_1751,N_2010);
nand U3200 (N_3200,N_1804,N_2211);
xor U3201 (N_3201,N_1518,N_2009);
and U3202 (N_3202,N_1790,N_2180);
or U3203 (N_3203,N_2312,N_1402);
or U3204 (N_3204,N_1875,N_1658);
and U3205 (N_3205,N_2312,N_1610);
and U3206 (N_3206,N_2063,N_1793);
xor U3207 (N_3207,N_1739,N_1708);
or U3208 (N_3208,N_1697,N_2282);
xor U3209 (N_3209,N_1719,N_1312);
nand U3210 (N_3210,N_1948,N_2309);
nor U3211 (N_3211,N_2246,N_2260);
or U3212 (N_3212,N_1677,N_1406);
and U3213 (N_3213,N_1348,N_2127);
nor U3214 (N_3214,N_2310,N_1984);
nor U3215 (N_3215,N_1686,N_2355);
nand U3216 (N_3216,N_1369,N_2217);
nor U3217 (N_3217,N_1579,N_1413);
and U3218 (N_3218,N_1795,N_1439);
and U3219 (N_3219,N_1356,N_1913);
xor U3220 (N_3220,N_1756,N_1225);
xor U3221 (N_3221,N_2184,N_1552);
xor U3222 (N_3222,N_1597,N_1599);
nand U3223 (N_3223,N_2347,N_1383);
xor U3224 (N_3224,N_2156,N_2251);
xor U3225 (N_3225,N_2164,N_1228);
nand U3226 (N_3226,N_2256,N_2088);
xor U3227 (N_3227,N_1402,N_1379);
or U3228 (N_3228,N_1502,N_1830);
and U3229 (N_3229,N_1752,N_2129);
or U3230 (N_3230,N_1440,N_1589);
xnor U3231 (N_3231,N_1837,N_1431);
xor U3232 (N_3232,N_2070,N_1964);
nand U3233 (N_3233,N_1384,N_1359);
nand U3234 (N_3234,N_1573,N_2358);
xnor U3235 (N_3235,N_1556,N_2159);
nor U3236 (N_3236,N_2371,N_1204);
nand U3237 (N_3237,N_2193,N_1554);
or U3238 (N_3238,N_1550,N_2334);
and U3239 (N_3239,N_1560,N_2351);
nand U3240 (N_3240,N_1609,N_2104);
or U3241 (N_3241,N_2259,N_2132);
xnor U3242 (N_3242,N_1365,N_1759);
xor U3243 (N_3243,N_2347,N_1783);
or U3244 (N_3244,N_2387,N_2236);
and U3245 (N_3245,N_2381,N_2338);
nand U3246 (N_3246,N_2214,N_1889);
or U3247 (N_3247,N_2029,N_1788);
nand U3248 (N_3248,N_1503,N_2136);
nand U3249 (N_3249,N_1743,N_1236);
or U3250 (N_3250,N_2205,N_2015);
and U3251 (N_3251,N_2160,N_1876);
and U3252 (N_3252,N_1247,N_1240);
nor U3253 (N_3253,N_2219,N_2383);
and U3254 (N_3254,N_2307,N_1746);
nand U3255 (N_3255,N_1460,N_1522);
or U3256 (N_3256,N_1554,N_1954);
and U3257 (N_3257,N_1249,N_1856);
xor U3258 (N_3258,N_2024,N_1943);
nor U3259 (N_3259,N_1801,N_2301);
nand U3260 (N_3260,N_2380,N_2079);
or U3261 (N_3261,N_2291,N_1885);
nand U3262 (N_3262,N_2353,N_1599);
xor U3263 (N_3263,N_1656,N_1499);
nor U3264 (N_3264,N_1855,N_1271);
nand U3265 (N_3265,N_1208,N_1666);
nor U3266 (N_3266,N_2193,N_2047);
nand U3267 (N_3267,N_2014,N_1710);
or U3268 (N_3268,N_2361,N_1967);
nor U3269 (N_3269,N_1891,N_2306);
nor U3270 (N_3270,N_1393,N_1758);
xnor U3271 (N_3271,N_1576,N_1432);
or U3272 (N_3272,N_2348,N_1456);
nor U3273 (N_3273,N_1337,N_1953);
and U3274 (N_3274,N_1220,N_2354);
nor U3275 (N_3275,N_2173,N_2072);
or U3276 (N_3276,N_1817,N_1464);
xnor U3277 (N_3277,N_1321,N_1447);
or U3278 (N_3278,N_2053,N_2392);
nor U3279 (N_3279,N_1245,N_1216);
and U3280 (N_3280,N_2333,N_1227);
nand U3281 (N_3281,N_1334,N_1861);
nor U3282 (N_3282,N_1842,N_2035);
or U3283 (N_3283,N_2063,N_1820);
or U3284 (N_3284,N_2013,N_1484);
nand U3285 (N_3285,N_2272,N_1833);
and U3286 (N_3286,N_2341,N_1855);
nor U3287 (N_3287,N_1248,N_2339);
nand U3288 (N_3288,N_2120,N_1441);
or U3289 (N_3289,N_1517,N_2323);
nor U3290 (N_3290,N_2134,N_2017);
or U3291 (N_3291,N_2050,N_1226);
or U3292 (N_3292,N_2211,N_1692);
xnor U3293 (N_3293,N_1823,N_1254);
nor U3294 (N_3294,N_1927,N_1404);
nor U3295 (N_3295,N_2390,N_1338);
and U3296 (N_3296,N_1804,N_2007);
and U3297 (N_3297,N_1630,N_1665);
or U3298 (N_3298,N_2016,N_1356);
and U3299 (N_3299,N_2251,N_2338);
and U3300 (N_3300,N_1723,N_2326);
nor U3301 (N_3301,N_2260,N_2355);
nor U3302 (N_3302,N_1812,N_1832);
nor U3303 (N_3303,N_1361,N_1933);
nor U3304 (N_3304,N_1849,N_2064);
nand U3305 (N_3305,N_1868,N_1961);
nor U3306 (N_3306,N_1479,N_1958);
xnor U3307 (N_3307,N_2330,N_1214);
nor U3308 (N_3308,N_2101,N_1644);
xnor U3309 (N_3309,N_1354,N_1681);
nor U3310 (N_3310,N_1764,N_1794);
nand U3311 (N_3311,N_1923,N_2295);
and U3312 (N_3312,N_1691,N_2245);
nand U3313 (N_3313,N_1404,N_2308);
nor U3314 (N_3314,N_1643,N_1283);
xnor U3315 (N_3315,N_1727,N_1867);
or U3316 (N_3316,N_2197,N_1980);
xor U3317 (N_3317,N_1684,N_1896);
nand U3318 (N_3318,N_1696,N_1384);
and U3319 (N_3319,N_2188,N_1800);
nand U3320 (N_3320,N_1700,N_1999);
and U3321 (N_3321,N_1774,N_1251);
nor U3322 (N_3322,N_1516,N_1362);
and U3323 (N_3323,N_2092,N_1832);
nand U3324 (N_3324,N_2039,N_1615);
or U3325 (N_3325,N_1353,N_1905);
nor U3326 (N_3326,N_2394,N_1751);
nand U3327 (N_3327,N_1717,N_2119);
nor U3328 (N_3328,N_1750,N_2181);
nor U3329 (N_3329,N_2078,N_2059);
xor U3330 (N_3330,N_2393,N_1864);
or U3331 (N_3331,N_1283,N_1650);
nand U3332 (N_3332,N_2133,N_2089);
xnor U3333 (N_3333,N_1322,N_1966);
xnor U3334 (N_3334,N_2089,N_1550);
nand U3335 (N_3335,N_1333,N_1464);
or U3336 (N_3336,N_1646,N_1697);
xor U3337 (N_3337,N_1959,N_2397);
or U3338 (N_3338,N_1303,N_1640);
nand U3339 (N_3339,N_2079,N_1963);
nor U3340 (N_3340,N_2366,N_1497);
or U3341 (N_3341,N_2170,N_1287);
nor U3342 (N_3342,N_1665,N_1777);
and U3343 (N_3343,N_1451,N_1424);
and U3344 (N_3344,N_1220,N_1379);
nor U3345 (N_3345,N_1973,N_2319);
nand U3346 (N_3346,N_1475,N_2049);
and U3347 (N_3347,N_1473,N_1405);
xor U3348 (N_3348,N_1502,N_1464);
or U3349 (N_3349,N_1226,N_2370);
and U3350 (N_3350,N_1730,N_1450);
and U3351 (N_3351,N_1296,N_1920);
and U3352 (N_3352,N_1953,N_1656);
and U3353 (N_3353,N_1749,N_1563);
xor U3354 (N_3354,N_2144,N_2131);
nand U3355 (N_3355,N_2295,N_1256);
nor U3356 (N_3356,N_1992,N_2207);
nand U3357 (N_3357,N_1250,N_1914);
nor U3358 (N_3358,N_2199,N_1530);
or U3359 (N_3359,N_2383,N_2033);
xor U3360 (N_3360,N_1212,N_1316);
or U3361 (N_3361,N_1294,N_2082);
and U3362 (N_3362,N_1781,N_1399);
nand U3363 (N_3363,N_1425,N_1397);
or U3364 (N_3364,N_1318,N_1704);
and U3365 (N_3365,N_1260,N_1958);
nor U3366 (N_3366,N_1289,N_1990);
and U3367 (N_3367,N_1512,N_1559);
and U3368 (N_3368,N_2148,N_1463);
or U3369 (N_3369,N_1379,N_1657);
and U3370 (N_3370,N_1513,N_2006);
xor U3371 (N_3371,N_1821,N_1559);
or U3372 (N_3372,N_1275,N_1702);
nor U3373 (N_3373,N_2229,N_1516);
nand U3374 (N_3374,N_1349,N_1314);
nand U3375 (N_3375,N_1900,N_1921);
and U3376 (N_3376,N_1336,N_1666);
nor U3377 (N_3377,N_2380,N_1868);
nor U3378 (N_3378,N_1959,N_2296);
and U3379 (N_3379,N_1856,N_1205);
and U3380 (N_3380,N_1985,N_2024);
nor U3381 (N_3381,N_1201,N_2099);
nand U3382 (N_3382,N_2287,N_2028);
nor U3383 (N_3383,N_2102,N_1467);
and U3384 (N_3384,N_1897,N_1346);
nand U3385 (N_3385,N_1573,N_2340);
or U3386 (N_3386,N_1692,N_1765);
or U3387 (N_3387,N_1685,N_2293);
or U3388 (N_3388,N_1865,N_1345);
xnor U3389 (N_3389,N_2290,N_1600);
xnor U3390 (N_3390,N_1273,N_1976);
and U3391 (N_3391,N_2120,N_1718);
or U3392 (N_3392,N_2114,N_1410);
and U3393 (N_3393,N_1823,N_2127);
or U3394 (N_3394,N_2355,N_1617);
nand U3395 (N_3395,N_1980,N_1395);
or U3396 (N_3396,N_1396,N_1355);
xor U3397 (N_3397,N_2353,N_1680);
xor U3398 (N_3398,N_2290,N_1252);
nor U3399 (N_3399,N_1535,N_1719);
and U3400 (N_3400,N_1272,N_1762);
xor U3401 (N_3401,N_1544,N_2373);
nand U3402 (N_3402,N_2273,N_1655);
xor U3403 (N_3403,N_1982,N_1931);
nand U3404 (N_3404,N_1737,N_1871);
nand U3405 (N_3405,N_1672,N_1561);
xnor U3406 (N_3406,N_2367,N_1816);
or U3407 (N_3407,N_1273,N_1581);
or U3408 (N_3408,N_2144,N_1999);
nand U3409 (N_3409,N_1270,N_2132);
or U3410 (N_3410,N_1513,N_1539);
xnor U3411 (N_3411,N_1924,N_1912);
and U3412 (N_3412,N_1565,N_1658);
or U3413 (N_3413,N_1945,N_1671);
and U3414 (N_3414,N_2229,N_1963);
and U3415 (N_3415,N_1288,N_2008);
or U3416 (N_3416,N_2359,N_1215);
nor U3417 (N_3417,N_1622,N_2347);
nor U3418 (N_3418,N_1626,N_2082);
xnor U3419 (N_3419,N_2148,N_2394);
xor U3420 (N_3420,N_1687,N_1644);
xnor U3421 (N_3421,N_1644,N_2263);
nand U3422 (N_3422,N_2324,N_1853);
and U3423 (N_3423,N_1791,N_1670);
nand U3424 (N_3424,N_1929,N_1738);
and U3425 (N_3425,N_1538,N_2256);
nand U3426 (N_3426,N_1996,N_1203);
xnor U3427 (N_3427,N_1634,N_1434);
and U3428 (N_3428,N_2286,N_1219);
xnor U3429 (N_3429,N_1403,N_2249);
nand U3430 (N_3430,N_2260,N_2031);
xor U3431 (N_3431,N_1339,N_2255);
nand U3432 (N_3432,N_1992,N_1943);
or U3433 (N_3433,N_2232,N_2118);
nor U3434 (N_3434,N_1321,N_1259);
nand U3435 (N_3435,N_1758,N_1286);
xnor U3436 (N_3436,N_1627,N_1837);
and U3437 (N_3437,N_1846,N_1339);
nor U3438 (N_3438,N_1803,N_1354);
and U3439 (N_3439,N_1324,N_1592);
or U3440 (N_3440,N_2181,N_1959);
nand U3441 (N_3441,N_1522,N_2364);
xnor U3442 (N_3442,N_1946,N_1912);
nor U3443 (N_3443,N_1725,N_1873);
nor U3444 (N_3444,N_1478,N_1550);
nor U3445 (N_3445,N_1849,N_2094);
nand U3446 (N_3446,N_1236,N_1873);
nand U3447 (N_3447,N_1218,N_1699);
and U3448 (N_3448,N_1775,N_2063);
or U3449 (N_3449,N_1326,N_1610);
and U3450 (N_3450,N_2253,N_1522);
nand U3451 (N_3451,N_1335,N_2262);
and U3452 (N_3452,N_2141,N_1454);
xor U3453 (N_3453,N_1570,N_2221);
nor U3454 (N_3454,N_2101,N_2111);
nand U3455 (N_3455,N_1319,N_2386);
nor U3456 (N_3456,N_1608,N_2191);
xor U3457 (N_3457,N_1504,N_1540);
and U3458 (N_3458,N_1650,N_1767);
nand U3459 (N_3459,N_1318,N_1885);
or U3460 (N_3460,N_1829,N_2133);
or U3461 (N_3461,N_1632,N_1920);
or U3462 (N_3462,N_2325,N_1534);
and U3463 (N_3463,N_2196,N_1206);
xor U3464 (N_3464,N_1362,N_2180);
and U3465 (N_3465,N_1628,N_1632);
xor U3466 (N_3466,N_1490,N_2135);
and U3467 (N_3467,N_1585,N_2382);
nand U3468 (N_3468,N_1445,N_1902);
nand U3469 (N_3469,N_2083,N_2097);
nand U3470 (N_3470,N_2263,N_1841);
and U3471 (N_3471,N_2350,N_2297);
or U3472 (N_3472,N_2348,N_1587);
nand U3473 (N_3473,N_2249,N_1774);
xor U3474 (N_3474,N_1898,N_1632);
nor U3475 (N_3475,N_1517,N_1924);
or U3476 (N_3476,N_1629,N_1604);
or U3477 (N_3477,N_1590,N_2070);
nor U3478 (N_3478,N_1724,N_1896);
and U3479 (N_3479,N_2241,N_1723);
and U3480 (N_3480,N_1480,N_1661);
nor U3481 (N_3481,N_1445,N_1651);
nand U3482 (N_3482,N_1373,N_1256);
nor U3483 (N_3483,N_1278,N_1913);
nor U3484 (N_3484,N_1750,N_1258);
and U3485 (N_3485,N_1798,N_1481);
xor U3486 (N_3486,N_1498,N_1944);
nor U3487 (N_3487,N_1334,N_1203);
nor U3488 (N_3488,N_2221,N_2397);
nor U3489 (N_3489,N_1890,N_2259);
nor U3490 (N_3490,N_1870,N_1307);
and U3491 (N_3491,N_1820,N_1992);
or U3492 (N_3492,N_1702,N_1227);
and U3493 (N_3493,N_2265,N_2165);
or U3494 (N_3494,N_2357,N_2225);
nor U3495 (N_3495,N_2209,N_1309);
or U3496 (N_3496,N_2266,N_2135);
nor U3497 (N_3497,N_1644,N_2177);
nor U3498 (N_3498,N_1978,N_1953);
and U3499 (N_3499,N_1944,N_1833);
and U3500 (N_3500,N_1397,N_1294);
nand U3501 (N_3501,N_1910,N_1552);
nor U3502 (N_3502,N_1868,N_1793);
and U3503 (N_3503,N_2104,N_1365);
xor U3504 (N_3504,N_1389,N_1954);
or U3505 (N_3505,N_2306,N_1811);
nor U3506 (N_3506,N_2124,N_1953);
or U3507 (N_3507,N_1456,N_1901);
xor U3508 (N_3508,N_1719,N_1437);
and U3509 (N_3509,N_1826,N_1646);
and U3510 (N_3510,N_1229,N_1261);
nand U3511 (N_3511,N_2280,N_1820);
and U3512 (N_3512,N_1591,N_2384);
or U3513 (N_3513,N_1992,N_1792);
xor U3514 (N_3514,N_2320,N_1645);
and U3515 (N_3515,N_1500,N_2368);
or U3516 (N_3516,N_1735,N_1823);
and U3517 (N_3517,N_2386,N_1867);
xor U3518 (N_3518,N_2094,N_1425);
nor U3519 (N_3519,N_1915,N_2037);
xor U3520 (N_3520,N_1485,N_1457);
or U3521 (N_3521,N_1211,N_1447);
nor U3522 (N_3522,N_1746,N_1911);
nor U3523 (N_3523,N_1832,N_2012);
nand U3524 (N_3524,N_2380,N_1298);
and U3525 (N_3525,N_2231,N_1805);
xnor U3526 (N_3526,N_2205,N_2291);
or U3527 (N_3527,N_1807,N_1415);
xnor U3528 (N_3528,N_1950,N_1202);
or U3529 (N_3529,N_1671,N_2124);
nor U3530 (N_3530,N_1656,N_1935);
and U3531 (N_3531,N_1890,N_2353);
xnor U3532 (N_3532,N_2122,N_1439);
xnor U3533 (N_3533,N_2392,N_1227);
and U3534 (N_3534,N_1254,N_1221);
nor U3535 (N_3535,N_2231,N_1758);
nor U3536 (N_3536,N_2326,N_1917);
nor U3537 (N_3537,N_1696,N_2243);
or U3538 (N_3538,N_1386,N_1953);
or U3539 (N_3539,N_1636,N_2388);
or U3540 (N_3540,N_1666,N_1641);
xnor U3541 (N_3541,N_1809,N_1816);
nand U3542 (N_3542,N_2193,N_1383);
or U3543 (N_3543,N_2379,N_1255);
nand U3544 (N_3544,N_1744,N_1829);
xor U3545 (N_3545,N_2224,N_2053);
xnor U3546 (N_3546,N_1280,N_1248);
xor U3547 (N_3547,N_2175,N_1218);
or U3548 (N_3548,N_2237,N_1211);
xnor U3549 (N_3549,N_1518,N_1413);
nor U3550 (N_3550,N_1283,N_1524);
or U3551 (N_3551,N_2050,N_2158);
and U3552 (N_3552,N_2305,N_2371);
nor U3553 (N_3553,N_2199,N_2252);
xor U3554 (N_3554,N_1622,N_1236);
xnor U3555 (N_3555,N_1694,N_1260);
xor U3556 (N_3556,N_1522,N_1323);
nor U3557 (N_3557,N_1436,N_1605);
or U3558 (N_3558,N_1202,N_1838);
and U3559 (N_3559,N_1998,N_1391);
nor U3560 (N_3560,N_1981,N_2040);
or U3561 (N_3561,N_2272,N_1710);
and U3562 (N_3562,N_2397,N_2029);
nand U3563 (N_3563,N_1989,N_1916);
nor U3564 (N_3564,N_2238,N_2167);
or U3565 (N_3565,N_1249,N_1978);
and U3566 (N_3566,N_2375,N_1462);
xor U3567 (N_3567,N_2191,N_1410);
nor U3568 (N_3568,N_1591,N_1964);
nor U3569 (N_3569,N_1399,N_1920);
nand U3570 (N_3570,N_1381,N_1331);
and U3571 (N_3571,N_1622,N_2391);
nand U3572 (N_3572,N_1479,N_1996);
nand U3573 (N_3573,N_1624,N_1390);
xor U3574 (N_3574,N_2216,N_2235);
nand U3575 (N_3575,N_1478,N_2324);
or U3576 (N_3576,N_2325,N_1712);
nand U3577 (N_3577,N_2253,N_1417);
and U3578 (N_3578,N_2255,N_1870);
nor U3579 (N_3579,N_1591,N_1373);
and U3580 (N_3580,N_2129,N_1495);
nor U3581 (N_3581,N_1455,N_1982);
nor U3582 (N_3582,N_2000,N_1943);
nand U3583 (N_3583,N_1428,N_1357);
nand U3584 (N_3584,N_1348,N_1573);
xor U3585 (N_3585,N_2394,N_1749);
nor U3586 (N_3586,N_1367,N_2202);
and U3587 (N_3587,N_1392,N_2398);
xor U3588 (N_3588,N_1741,N_1355);
nand U3589 (N_3589,N_1900,N_2217);
and U3590 (N_3590,N_1910,N_2162);
and U3591 (N_3591,N_1247,N_1258);
or U3592 (N_3592,N_1427,N_1324);
nor U3593 (N_3593,N_1477,N_2229);
and U3594 (N_3594,N_1295,N_1829);
nand U3595 (N_3595,N_1854,N_1849);
xnor U3596 (N_3596,N_1250,N_1560);
nand U3597 (N_3597,N_1338,N_1350);
nand U3598 (N_3598,N_1763,N_2264);
nor U3599 (N_3599,N_1224,N_2024);
nor U3600 (N_3600,N_3189,N_2529);
and U3601 (N_3601,N_3163,N_2671);
nor U3602 (N_3602,N_3494,N_3431);
and U3603 (N_3603,N_3266,N_2567);
nand U3604 (N_3604,N_2993,N_2771);
or U3605 (N_3605,N_3288,N_2592);
nor U3606 (N_3606,N_3523,N_2604);
or U3607 (N_3607,N_2984,N_3243);
nor U3608 (N_3608,N_2721,N_2576);
and U3609 (N_3609,N_3521,N_2920);
nor U3610 (N_3610,N_2698,N_2942);
and U3611 (N_3611,N_2875,N_3184);
xor U3612 (N_3612,N_3109,N_3096);
or U3613 (N_3613,N_2645,N_2553);
and U3614 (N_3614,N_3472,N_3107);
nor U3615 (N_3615,N_2407,N_3596);
and U3616 (N_3616,N_3457,N_2850);
nand U3617 (N_3617,N_3597,N_2620);
xnor U3618 (N_3618,N_2663,N_2437);
and U3619 (N_3619,N_2523,N_2445);
and U3620 (N_3620,N_3347,N_3415);
xor U3621 (N_3621,N_3402,N_2968);
and U3622 (N_3622,N_3139,N_2848);
nor U3623 (N_3623,N_2624,N_3587);
or U3624 (N_3624,N_3204,N_3039);
nor U3625 (N_3625,N_3337,N_3529);
xor U3626 (N_3626,N_2908,N_3146);
and U3627 (N_3627,N_2644,N_2625);
or U3628 (N_3628,N_2999,N_3191);
and U3629 (N_3629,N_3537,N_2651);
nor U3630 (N_3630,N_2737,N_2617);
xnor U3631 (N_3631,N_3501,N_2820);
xnor U3632 (N_3632,N_3065,N_2494);
nand U3633 (N_3633,N_2809,N_3125);
nand U3634 (N_3634,N_3103,N_3242);
and U3635 (N_3635,N_2686,N_2932);
nand U3636 (N_3636,N_3187,N_3100);
or U3637 (N_3637,N_2889,N_2923);
nor U3638 (N_3638,N_2898,N_2668);
nor U3639 (N_3639,N_2454,N_2715);
xnor U3640 (N_3640,N_3438,N_2697);
xor U3641 (N_3641,N_3018,N_2703);
or U3642 (N_3642,N_3250,N_2521);
and U3643 (N_3643,N_3376,N_3491);
and U3644 (N_3644,N_3366,N_2425);
and U3645 (N_3645,N_3442,N_3154);
and U3646 (N_3646,N_3225,N_3031);
and U3647 (N_3647,N_3538,N_3573);
nor U3648 (N_3648,N_2650,N_3594);
nand U3649 (N_3649,N_2824,N_2404);
nor U3650 (N_3650,N_2777,N_2902);
and U3651 (N_3651,N_3291,N_3240);
nand U3652 (N_3652,N_2467,N_3554);
nor U3653 (N_3653,N_2803,N_3540);
xnor U3654 (N_3654,N_3256,N_2863);
xnor U3655 (N_3655,N_2545,N_2796);
nand U3656 (N_3656,N_3008,N_3492);
or U3657 (N_3657,N_2989,N_3598);
xnor U3658 (N_3658,N_3053,N_3413);
xor U3659 (N_3659,N_2979,N_2856);
xor U3660 (N_3660,N_3434,N_2912);
or U3661 (N_3661,N_2688,N_2519);
nand U3662 (N_3662,N_2716,N_2955);
and U3663 (N_3663,N_2720,N_3002);
and U3664 (N_3664,N_3326,N_2974);
xor U3665 (N_3665,N_2578,N_2757);
and U3666 (N_3666,N_2776,N_3268);
nor U3667 (N_3667,N_3003,N_2699);
xor U3668 (N_3668,N_3206,N_2866);
xor U3669 (N_3669,N_3112,N_3421);
or U3670 (N_3670,N_2452,N_3576);
or U3671 (N_3671,N_2988,N_3488);
nor U3672 (N_3672,N_2951,N_3270);
nor U3673 (N_3673,N_2954,N_3228);
or U3674 (N_3674,N_2556,N_2832);
nor U3675 (N_3675,N_2732,N_3176);
nor U3676 (N_3676,N_2901,N_2774);
nor U3677 (N_3677,N_3387,N_3244);
nor U3678 (N_3678,N_2543,N_2835);
xor U3679 (N_3679,N_3528,N_2925);
and U3680 (N_3680,N_3482,N_2441);
and U3681 (N_3681,N_2655,N_2811);
and U3682 (N_3682,N_2963,N_2797);
nand U3683 (N_3683,N_2411,N_2939);
xor U3684 (N_3684,N_2829,N_2591);
and U3685 (N_3685,N_2563,N_3060);
and U3686 (N_3686,N_3114,N_3199);
or U3687 (N_3687,N_2477,N_3503);
and U3688 (N_3688,N_3033,N_3271);
nand U3689 (N_3689,N_3302,N_3247);
and U3690 (N_3690,N_2432,N_3422);
or U3691 (N_3691,N_3460,N_2930);
nand U3692 (N_3692,N_2682,N_2630);
nand U3693 (N_3693,N_2983,N_2990);
nand U3694 (N_3694,N_3052,N_2507);
nor U3695 (N_3695,N_2967,N_2742);
nand U3696 (N_3696,N_3452,N_2847);
xnor U3697 (N_3697,N_2778,N_3339);
nand U3698 (N_3698,N_3177,N_2730);
nor U3699 (N_3699,N_2938,N_2472);
and U3700 (N_3700,N_2540,N_2812);
or U3701 (N_3701,N_3294,N_2665);
and U3702 (N_3702,N_2548,N_3577);
and U3703 (N_3703,N_3304,N_3589);
xnor U3704 (N_3704,N_2457,N_2729);
nand U3705 (N_3705,N_2428,N_3511);
or U3706 (N_3706,N_2629,N_2915);
and U3707 (N_3707,N_2957,N_2568);
and U3708 (N_3708,N_3128,N_2570);
nor U3709 (N_3709,N_2561,N_3314);
or U3710 (N_3710,N_2450,N_2637);
xor U3711 (N_3711,N_2936,N_3106);
nor U3712 (N_3712,N_3217,N_3440);
nand U3713 (N_3713,N_2818,N_3553);
nor U3714 (N_3714,N_3175,N_2764);
nand U3715 (N_3715,N_3526,N_3342);
nor U3716 (N_3716,N_2622,N_2470);
or U3717 (N_3717,N_2836,N_2631);
nand U3718 (N_3718,N_3080,N_2634);
nand U3719 (N_3719,N_3162,N_2653);
and U3720 (N_3720,N_3433,N_2572);
xnor U3721 (N_3721,N_3298,N_2654);
nor U3722 (N_3722,N_3325,N_3098);
or U3723 (N_3723,N_2734,N_2941);
and U3724 (N_3724,N_2804,N_2887);
or U3725 (N_3725,N_3513,N_2892);
and U3726 (N_3726,N_3129,N_2897);
xnor U3727 (N_3727,N_3439,N_3332);
xnor U3728 (N_3728,N_3520,N_3500);
nand U3729 (N_3729,N_2858,N_3370);
xor U3730 (N_3730,N_2577,N_3470);
or U3731 (N_3731,N_3046,N_2891);
or U3732 (N_3732,N_2869,N_2439);
xor U3733 (N_3733,N_3006,N_2790);
xor U3734 (N_3734,N_3159,N_2746);
xor U3735 (N_3735,N_2792,N_2642);
nand U3736 (N_3736,N_3093,N_2985);
xnor U3737 (N_3737,N_2594,N_2574);
and U3738 (N_3738,N_2408,N_2962);
and U3739 (N_3739,N_2934,N_2751);
nand U3740 (N_3740,N_3481,N_3341);
nand U3741 (N_3741,N_2557,N_2659);
and U3742 (N_3742,N_2909,N_3144);
or U3743 (N_3743,N_2621,N_2530);
nor U3744 (N_3744,N_3135,N_2471);
xor U3745 (N_3745,N_2406,N_3253);
or U3746 (N_3746,N_3531,N_3336);
nand U3747 (N_3747,N_3059,N_3581);
nor U3748 (N_3748,N_2768,N_2843);
nand U3749 (N_3749,N_3280,N_3547);
and U3750 (N_3750,N_2597,N_2596);
nand U3751 (N_3751,N_3149,N_3077);
nor U3752 (N_3752,N_3377,N_2464);
or U3753 (N_3753,N_3373,N_3113);
xor U3754 (N_3754,N_3216,N_3117);
and U3755 (N_3755,N_3444,N_3365);
nor U3756 (N_3756,N_3049,N_2602);
and U3757 (N_3757,N_3075,N_3207);
nor U3758 (N_3758,N_2943,N_3374);
nor U3759 (N_3759,N_3548,N_2788);
and U3760 (N_3760,N_3475,N_3382);
xnor U3761 (N_3761,N_3131,N_2834);
nor U3762 (N_3762,N_3557,N_3512);
or U3763 (N_3763,N_2773,N_3579);
or U3764 (N_3764,N_2695,N_3289);
nor U3765 (N_3765,N_3168,N_3561);
or U3766 (N_3766,N_2462,N_3388);
xor U3767 (N_3767,N_3023,N_2640);
or U3768 (N_3768,N_2899,N_2724);
or U3769 (N_3769,N_3478,N_3248);
and U3770 (N_3770,N_2722,N_2485);
and U3771 (N_3771,N_3297,N_3156);
nand U3772 (N_3772,N_2833,N_2917);
nor U3773 (N_3773,N_2853,N_3563);
nand U3774 (N_3774,N_2460,N_2584);
nand U3775 (N_3775,N_3405,N_2403);
xnor U3776 (N_3776,N_3510,N_2839);
xor U3777 (N_3777,N_3437,N_3132);
xor U3778 (N_3778,N_2753,N_2517);
nor U3779 (N_3779,N_3036,N_2633);
xor U3780 (N_3780,N_3122,N_2546);
nor U3781 (N_3781,N_2501,N_2965);
nand U3782 (N_3782,N_2489,N_3185);
nand U3783 (N_3783,N_3322,N_2518);
or U3784 (N_3784,N_3571,N_3447);
or U3785 (N_3785,N_2453,N_3186);
or U3786 (N_3786,N_3200,N_2515);
xnor U3787 (N_3787,N_2958,N_2918);
nor U3788 (N_3788,N_2947,N_3264);
and U3789 (N_3789,N_3467,N_3476);
and U3790 (N_3790,N_2800,N_3272);
nand U3791 (N_3791,N_3234,N_3198);
nor U3792 (N_3792,N_2550,N_2717);
nand U3793 (N_3793,N_2924,N_2613);
nor U3794 (N_3794,N_2646,N_3195);
nand U3795 (N_3795,N_2440,N_3153);
xnor U3796 (N_3796,N_2708,N_3284);
xnor U3797 (N_3797,N_2883,N_3543);
nor U3798 (N_3798,N_3121,N_2880);
and U3799 (N_3799,N_2490,N_3340);
nand U3800 (N_3800,N_3315,N_3252);
and U3801 (N_3801,N_3172,N_2527);
nand U3802 (N_3802,N_2718,N_2614);
or U3803 (N_3803,N_2881,N_3427);
or U3804 (N_3804,N_2693,N_3221);
or U3805 (N_3805,N_2844,N_2973);
or U3806 (N_3806,N_3222,N_2714);
xor U3807 (N_3807,N_3567,N_2615);
nand U3808 (N_3808,N_3285,N_2483);
nor U3809 (N_3809,N_2535,N_3585);
xor U3810 (N_3810,N_3260,N_2429);
nor U3811 (N_3811,N_3044,N_3559);
xor U3812 (N_3812,N_3353,N_3164);
or U3813 (N_3813,N_3335,N_3257);
and U3814 (N_3814,N_2652,N_3454);
nand U3815 (N_3815,N_3130,N_2735);
and U3816 (N_3816,N_3527,N_2493);
or U3817 (N_3817,N_2632,N_3108);
nand U3818 (N_3818,N_2444,N_3517);
nor U3819 (N_3819,N_3180,N_2799);
nor U3820 (N_3820,N_3010,N_2598);
nor U3821 (N_3821,N_2896,N_2745);
or U3822 (N_3822,N_2435,N_2571);
nor U3823 (N_3823,N_3102,N_2784);
or U3824 (N_3824,N_3487,N_2562);
nand U3825 (N_3825,N_2770,N_3522);
or U3826 (N_3826,N_2935,N_2443);
and U3827 (N_3827,N_2595,N_3351);
or U3828 (N_3828,N_3533,N_3534);
nor U3829 (N_3829,N_2558,N_2961);
and U3830 (N_3830,N_2786,N_3011);
xor U3831 (N_3831,N_3329,N_2551);
and U3832 (N_3832,N_2420,N_2914);
and U3833 (N_3833,N_3094,N_2674);
and U3834 (N_3834,N_2959,N_3231);
nand U3835 (N_3835,N_3530,N_2903);
and U3836 (N_3836,N_3568,N_3138);
or U3837 (N_3837,N_2672,N_3518);
nand U3838 (N_3838,N_2952,N_2638);
xnor U3839 (N_3839,N_2667,N_2566);
nor U3840 (N_3840,N_2760,N_3550);
nor U3841 (N_3841,N_3319,N_3480);
xor U3842 (N_3842,N_2680,N_2534);
and U3843 (N_3843,N_3165,N_3014);
or U3844 (N_3844,N_2775,N_3566);
xnor U3845 (N_3845,N_3028,N_2612);
and U3846 (N_3846,N_2492,N_3582);
nand U3847 (N_3847,N_2884,N_3083);
xor U3848 (N_3848,N_2929,N_2877);
and U3849 (N_3849,N_3384,N_2678);
and U3850 (N_3850,N_3495,N_3073);
nor U3851 (N_3851,N_2451,N_3197);
nor U3852 (N_3852,N_2861,N_3506);
nor U3853 (N_3853,N_2639,N_3095);
and U3854 (N_3854,N_3593,N_2971);
or U3855 (N_3855,N_2755,N_3355);
or U3856 (N_3856,N_2830,N_3258);
nand U3857 (N_3857,N_2673,N_3430);
nand U3858 (N_3858,N_3147,N_2458);
or U3859 (N_3859,N_3432,N_3292);
xnor U3860 (N_3860,N_2821,N_3343);
nand U3861 (N_3861,N_3082,N_2750);
xor U3862 (N_3862,N_2991,N_3544);
and U3863 (N_3863,N_2749,N_2748);
or U3864 (N_3864,N_3461,N_3140);
and U3865 (N_3865,N_3532,N_2660);
or U3866 (N_3866,N_2484,N_3215);
nor U3867 (N_3867,N_3323,N_2867);
xor U3868 (N_3868,N_2826,N_2763);
nand U3869 (N_3869,N_2498,N_2502);
or U3870 (N_3870,N_2948,N_2785);
or U3871 (N_3871,N_3090,N_2427);
or U3872 (N_3872,N_2499,N_3584);
xnor U3873 (N_3873,N_3352,N_3182);
xnor U3874 (N_3874,N_2906,N_2400);
and U3875 (N_3875,N_3330,N_2446);
and U3876 (N_3876,N_2879,N_3359);
and U3877 (N_3877,N_2669,N_2780);
xnor U3878 (N_3878,N_2831,N_3212);
or U3879 (N_3879,N_3290,N_3265);
or U3880 (N_3880,N_2656,N_3552);
and U3881 (N_3881,N_3001,N_2414);
nand U3882 (N_3882,N_3193,N_3473);
nand U3883 (N_3883,N_2946,N_2463);
nand U3884 (N_3884,N_2433,N_3118);
nor U3885 (N_3885,N_2738,N_3443);
xnor U3886 (N_3886,N_2536,N_2878);
nand U3887 (N_3887,N_2468,N_2982);
nand U3888 (N_3888,N_2998,N_2560);
or U3889 (N_3889,N_2418,N_3397);
nand U3890 (N_3890,N_2419,N_2661);
or U3891 (N_3891,N_2580,N_2476);
and U3892 (N_3892,N_2933,N_3262);
nand U3893 (N_3893,N_2859,N_3371);
and U3894 (N_3894,N_2694,N_2825);
xnor U3895 (N_3895,N_2459,N_2506);
xnor U3896 (N_3896,N_2793,N_2713);
nand U3897 (N_3897,N_2872,N_3578);
nand U3898 (N_3898,N_2554,N_3309);
nor U3899 (N_3899,N_3205,N_3562);
xnor U3900 (N_3900,N_3456,N_3145);
and U3901 (N_3901,N_3338,N_3219);
or U3902 (N_3902,N_3084,N_2508);
nand U3903 (N_3903,N_3378,N_2685);
nand U3904 (N_3904,N_3591,N_3246);
xor U3905 (N_3905,N_2913,N_3004);
and U3906 (N_3906,N_2975,N_2565);
nor U3907 (N_3907,N_2945,N_2977);
nor U3908 (N_3908,N_2658,N_2588);
nor U3909 (N_3909,N_3190,N_2772);
nand U3910 (N_3910,N_2416,N_3201);
nor U3911 (N_3911,N_3555,N_2648);
nand U3912 (N_3912,N_2728,N_3091);
nand U3913 (N_3913,N_2607,N_2865);
or U3914 (N_3914,N_3392,N_2806);
and U3915 (N_3915,N_2860,N_3043);
nor U3916 (N_3916,N_3462,N_2705);
nand U3917 (N_3917,N_3345,N_3465);
and U3918 (N_3918,N_2449,N_3021);
and U3919 (N_3919,N_3072,N_2854);
or U3920 (N_3920,N_2928,N_3275);
nand U3921 (N_3921,N_3574,N_2417);
or U3922 (N_3922,N_3549,N_2618);
and U3923 (N_3923,N_3070,N_2885);
or U3924 (N_3924,N_3545,N_3398);
or U3925 (N_3925,N_2497,N_2926);
xor U3926 (N_3926,N_2744,N_3054);
nor U3927 (N_3927,N_3391,N_2766);
and U3928 (N_3928,N_2995,N_3237);
xnor U3929 (N_3929,N_3403,N_3572);
or U3930 (N_3930,N_2978,N_3312);
nand U3931 (N_3931,N_2845,N_3167);
xor U3932 (N_3932,N_2816,N_3029);
nand U3933 (N_3933,N_2849,N_3287);
nor U3934 (N_3934,N_2949,N_3379);
xnor U3935 (N_3935,N_3399,N_3061);
and U3936 (N_3936,N_3375,N_2600);
nor U3937 (N_3937,N_2992,N_2402);
or U3938 (N_3938,N_3469,N_3241);
or U3939 (N_3939,N_2616,N_2681);
nand U3940 (N_3940,N_2707,N_3045);
or U3941 (N_3941,N_3181,N_2609);
and U3942 (N_3942,N_2711,N_2731);
and U3943 (N_3943,N_2552,N_3344);
and U3944 (N_3944,N_3441,N_3306);
or U3945 (N_3945,N_2538,N_3238);
nor U3946 (N_3946,N_3449,N_3435);
and U3947 (N_3947,N_3227,N_2692);
nand U3948 (N_3948,N_2469,N_3000);
or U3949 (N_3949,N_2904,N_3356);
nand U3950 (N_3950,N_2813,N_3064);
and U3951 (N_3951,N_2549,N_2657);
nor U3952 (N_3952,N_3068,N_3224);
xor U3953 (N_3953,N_3569,N_3024);
and U3954 (N_3954,N_2481,N_3448);
nor U3955 (N_3955,N_2670,N_3453);
and U3956 (N_3956,N_2666,N_3575);
nand U3957 (N_3957,N_2555,N_3389);
or U3958 (N_3958,N_3551,N_2805);
nand U3959 (N_3959,N_2868,N_2542);
and U3960 (N_3960,N_2579,N_2505);
nand U3961 (N_3961,N_3499,N_2593);
nand U3962 (N_3962,N_2987,N_3396);
or U3963 (N_3963,N_2430,N_2514);
nor U3964 (N_3964,N_2662,N_3174);
or U3965 (N_3965,N_3069,N_3411);
or U3966 (N_3966,N_2886,N_2465);
nand U3967 (N_3967,N_3120,N_2921);
nand U3968 (N_3968,N_3474,N_3286);
xor U3969 (N_3969,N_2496,N_2761);
and U3970 (N_3970,N_2611,N_2478);
nand U3971 (N_3971,N_2851,N_2931);
nor U3972 (N_3972,N_2423,N_3299);
and U3973 (N_3973,N_2559,N_2413);
nand U3974 (N_3974,N_2964,N_2480);
nor U3975 (N_3975,N_3136,N_2422);
or U3976 (N_3976,N_2544,N_3025);
nand U3977 (N_3977,N_3141,N_3542);
and U3978 (N_3978,N_2706,N_2976);
xor U3979 (N_3979,N_3560,N_2725);
or U3980 (N_3980,N_3087,N_3005);
or U3981 (N_3981,N_2719,N_2573);
or U3982 (N_3982,N_3358,N_3196);
and U3983 (N_3983,N_2726,N_3362);
nand U3984 (N_3984,N_2838,N_2828);
xnor U3985 (N_3985,N_3179,N_2405);
and U3986 (N_3986,N_3079,N_2980);
xnor U3987 (N_3987,N_2599,N_2910);
or U3988 (N_3988,N_2564,N_3386);
and U3989 (N_3989,N_2736,N_2700);
nor U3990 (N_3990,N_3160,N_3493);
or U3991 (N_3991,N_2819,N_3307);
xnor U3992 (N_3992,N_3328,N_3209);
and U3993 (N_3993,N_2873,N_2511);
or U3994 (N_3994,N_3171,N_3331);
xnor U3995 (N_3995,N_3081,N_2922);
and U3996 (N_3996,N_2798,N_3426);
or U3997 (N_3997,N_3220,N_2937);
xor U3998 (N_3998,N_3058,N_3541);
and U3999 (N_3999,N_2525,N_2894);
nor U4000 (N_4000,N_2676,N_2767);
xor U4001 (N_4001,N_2996,N_3047);
nand U4002 (N_4002,N_3498,N_3514);
xor U4003 (N_4003,N_3283,N_2474);
xnor U4004 (N_4004,N_2664,N_3295);
or U4005 (N_4005,N_2628,N_2743);
or U4006 (N_4006,N_3126,N_3111);
xor U4007 (N_4007,N_3502,N_3213);
nor U4008 (N_4008,N_3170,N_3274);
or U4009 (N_4009,N_3278,N_2782);
and U4010 (N_4010,N_3229,N_3394);
or U4011 (N_4011,N_2704,N_3468);
nand U4012 (N_4012,N_2575,N_2972);
nor U4013 (N_4013,N_2807,N_3183);
xor U4014 (N_4014,N_3477,N_2758);
and U4015 (N_4015,N_3458,N_3048);
and U4016 (N_4016,N_3074,N_3590);
nor U4017 (N_4017,N_2608,N_3369);
nor U4018 (N_4018,N_3419,N_3418);
and U4019 (N_4019,N_3214,N_3305);
nor U4020 (N_4020,N_3363,N_2619);
and U4021 (N_4021,N_3055,N_3105);
or U4022 (N_4022,N_3150,N_3595);
nor U4023 (N_4023,N_3414,N_3208);
xnor U4024 (N_4024,N_3504,N_3393);
nand U4025 (N_4025,N_2586,N_3158);
and U4026 (N_4026,N_3486,N_3515);
or U4027 (N_4027,N_2814,N_3311);
xnor U4028 (N_4028,N_3255,N_2635);
and U4029 (N_4029,N_3428,N_3484);
nand U4030 (N_4030,N_3556,N_3279);
or U4031 (N_4031,N_3211,N_2410);
and U4032 (N_4032,N_2475,N_3203);
nor U4033 (N_4033,N_3483,N_2966);
xor U4034 (N_4034,N_3032,N_3202);
or U4035 (N_4035,N_2781,N_2907);
or U4036 (N_4036,N_3509,N_3233);
and U4037 (N_4037,N_3583,N_3037);
nor U4038 (N_4038,N_3019,N_3056);
nand U4039 (N_4039,N_3381,N_3066);
and U4040 (N_4040,N_2723,N_2986);
and U4041 (N_4041,N_3261,N_3218);
and U4042 (N_4042,N_3310,N_3321);
xor U4043 (N_4043,N_3259,N_2900);
xor U4044 (N_4044,N_2882,N_3042);
xor U4045 (N_4045,N_3350,N_3599);
xnor U4046 (N_4046,N_3301,N_2520);
xnor U4047 (N_4047,N_3143,N_2857);
xnor U4048 (N_4048,N_3346,N_2495);
nor U4049 (N_4049,N_3115,N_3116);
nor U4050 (N_4050,N_2582,N_2456);
nor U4051 (N_4051,N_3592,N_3463);
and U4052 (N_4052,N_2895,N_3565);
or U4053 (N_4053,N_2532,N_2815);
or U4054 (N_4054,N_2531,N_3360);
xor U4055 (N_4055,N_2862,N_2684);
xnor U4056 (N_4056,N_3016,N_3429);
xor U4057 (N_4057,N_2970,N_3027);
nor U4058 (N_4058,N_2919,N_3249);
nand U4059 (N_4059,N_3099,N_3507);
and U4060 (N_4060,N_3546,N_3137);
xor U4061 (N_4061,N_2687,N_3409);
and U4062 (N_4062,N_2769,N_3071);
nand U4063 (N_4063,N_2754,N_2759);
nor U4064 (N_4064,N_3089,N_2626);
and U4065 (N_4065,N_2822,N_3536);
nor U4066 (N_4066,N_3152,N_3110);
xnor U4067 (N_4067,N_3178,N_3327);
nand U4068 (N_4068,N_2794,N_2528);
nand U4069 (N_4069,N_3026,N_2436);
xnor U4070 (N_4070,N_2956,N_2739);
nor U4071 (N_4071,N_2509,N_3239);
or U4072 (N_4072,N_2569,N_2583);
or U4073 (N_4073,N_3151,N_3235);
or U4074 (N_4074,N_3230,N_3007);
nand U4075 (N_4075,N_3119,N_2679);
nand U4076 (N_4076,N_3086,N_2916);
xor U4077 (N_4077,N_3067,N_3017);
or U4078 (N_4078,N_2969,N_3210);
and U4079 (N_4079,N_3400,N_2482);
xor U4080 (N_4080,N_2756,N_2512);
or U4081 (N_4081,N_3148,N_2997);
and U4082 (N_4082,N_3505,N_2733);
nor U4083 (N_4083,N_3063,N_3564);
nor U4084 (N_4084,N_3316,N_2606);
nand U4085 (N_4085,N_2855,N_2712);
nand U4086 (N_4086,N_2533,N_3535);
xnor U4087 (N_4087,N_2636,N_3455);
or U4088 (N_4088,N_3009,N_3124);
xnor U4089 (N_4089,N_3088,N_2649);
xnor U4090 (N_4090,N_3404,N_3303);
nand U4091 (N_4091,N_2846,N_3097);
xor U4092 (N_4092,N_3308,N_3570);
nor U4093 (N_4093,N_3236,N_3334);
nor U4094 (N_4094,N_2709,N_2466);
or U4095 (N_4095,N_2401,N_3580);
xor U4096 (N_4096,N_3194,N_3318);
nand U4097 (N_4097,N_3519,N_3408);
or U4098 (N_4098,N_3296,N_3436);
xor U4099 (N_4099,N_2701,N_3076);
nor U4100 (N_4100,N_2752,N_2643);
and U4101 (N_4101,N_3416,N_2415);
nor U4102 (N_4102,N_3263,N_2448);
or U4103 (N_4103,N_2808,N_2940);
nor U4104 (N_4104,N_3364,N_2409);
nand U4105 (N_4105,N_3226,N_2981);
or U4106 (N_4106,N_2431,N_3104);
xor U4107 (N_4107,N_2641,N_3524);
nand U4108 (N_4108,N_2727,N_3057);
and U4109 (N_4109,N_2953,N_3281);
nand U4110 (N_4110,N_2696,N_2888);
nand U4111 (N_4111,N_3357,N_3155);
xor U4112 (N_4112,N_3348,N_2791);
xor U4113 (N_4113,N_2442,N_3277);
and U4114 (N_4114,N_3267,N_3051);
and U4115 (N_4115,N_3192,N_2871);
nand U4116 (N_4116,N_3423,N_3038);
or U4117 (N_4117,N_3245,N_2864);
xor U4118 (N_4118,N_2810,N_2601);
or U4119 (N_4119,N_3232,N_2827);
nand U4120 (N_4120,N_3078,N_3142);
and U4121 (N_4121,N_3169,N_2516);
and U4122 (N_4122,N_3383,N_3349);
or U4123 (N_4123,N_2890,N_3406);
or U4124 (N_4124,N_3489,N_2852);
and U4125 (N_4125,N_3127,N_2547);
and U4126 (N_4126,N_2500,N_3516);
xor U4127 (N_4127,N_2455,N_3223);
xnor U4128 (N_4128,N_2424,N_2741);
nor U4129 (N_4129,N_3293,N_2504);
nor U4130 (N_4130,N_3471,N_2447);
nand U4131 (N_4131,N_3022,N_3133);
nand U4132 (N_4132,N_2817,N_2675);
or U4133 (N_4133,N_2927,N_2539);
and U4134 (N_4134,N_2905,N_2590);
and U4135 (N_4135,N_3368,N_2438);
and U4136 (N_4136,N_3015,N_2487);
nand U4137 (N_4137,N_3251,N_2762);
and U4138 (N_4138,N_2689,N_2627);
nor U4139 (N_4139,N_3035,N_3020);
and U4140 (N_4140,N_3085,N_3390);
or U4141 (N_4141,N_3276,N_2479);
nand U4142 (N_4142,N_2581,N_3525);
nand U4143 (N_4143,N_3558,N_3372);
xor U4144 (N_4144,N_3012,N_3173);
xnor U4145 (N_4145,N_3485,N_3123);
nor U4146 (N_4146,N_2541,N_3385);
or U4147 (N_4147,N_3466,N_2876);
nand U4148 (N_4148,N_2840,N_2683);
nor U4149 (N_4149,N_2647,N_2587);
xnor U4150 (N_4150,N_3539,N_2837);
and U4151 (N_4151,N_3354,N_2522);
nor U4152 (N_4152,N_2823,N_3062);
nand U4153 (N_4153,N_2434,N_3420);
and U4154 (N_4154,N_2801,N_3451);
or U4155 (N_4155,N_2691,N_3367);
nand U4156 (N_4156,N_3588,N_2874);
nand U4157 (N_4157,N_3050,N_2537);
nand U4158 (N_4158,N_2787,N_3410);
and U4159 (N_4159,N_2421,N_2960);
nor U4160 (N_4160,N_3034,N_2491);
or U4161 (N_4161,N_2690,N_2526);
nor U4162 (N_4162,N_3040,N_3254);
nor U4163 (N_4163,N_3300,N_2841);
nor U4164 (N_4164,N_3161,N_3166);
and U4165 (N_4165,N_3464,N_3401);
nor U4166 (N_4166,N_3445,N_3412);
or U4167 (N_4167,N_2524,N_2426);
xor U4168 (N_4168,N_2893,N_2412);
xor U4169 (N_4169,N_2589,N_2603);
nor U4170 (N_4170,N_2510,N_3188);
xnor U4171 (N_4171,N_2842,N_3496);
xnor U4172 (N_4172,N_2585,N_3361);
and U4173 (N_4173,N_2503,N_2795);
nand U4174 (N_4174,N_2623,N_2783);
and U4175 (N_4175,N_2702,N_2473);
nor U4176 (N_4176,N_2513,N_3269);
or U4177 (N_4177,N_3030,N_3013);
nor U4178 (N_4178,N_3320,N_2870);
or U4179 (N_4179,N_2486,N_3273);
nand U4180 (N_4180,N_3407,N_3586);
nand U4181 (N_4181,N_3459,N_3333);
or U4182 (N_4182,N_3092,N_3446);
xnor U4183 (N_4183,N_3041,N_2911);
xor U4184 (N_4184,N_3282,N_2610);
xnor U4185 (N_4185,N_3313,N_2461);
nand U4186 (N_4186,N_3317,N_3395);
or U4187 (N_4187,N_3324,N_2779);
nand U4188 (N_4188,N_2488,N_2950);
nor U4189 (N_4189,N_2789,N_2605);
or U4190 (N_4190,N_2944,N_3417);
nand U4191 (N_4191,N_3450,N_2765);
and U4192 (N_4192,N_2747,N_3424);
nand U4193 (N_4193,N_2802,N_2677);
xor U4194 (N_4194,N_3134,N_3157);
nor U4195 (N_4195,N_2710,N_3497);
nand U4196 (N_4196,N_3425,N_3380);
nand U4197 (N_4197,N_3508,N_3101);
nor U4198 (N_4198,N_3490,N_3479);
xor U4199 (N_4199,N_2994,N_2740);
xnor U4200 (N_4200,N_3335,N_3221);
nand U4201 (N_4201,N_3147,N_2464);
xnor U4202 (N_4202,N_3105,N_3584);
nor U4203 (N_4203,N_3537,N_3023);
xor U4204 (N_4204,N_3099,N_3287);
or U4205 (N_4205,N_2661,N_2449);
or U4206 (N_4206,N_3561,N_2817);
and U4207 (N_4207,N_2558,N_2852);
nor U4208 (N_4208,N_2636,N_3453);
nor U4209 (N_4209,N_3006,N_2570);
or U4210 (N_4210,N_2425,N_2879);
nand U4211 (N_4211,N_3253,N_3565);
nand U4212 (N_4212,N_2661,N_2802);
or U4213 (N_4213,N_2644,N_2906);
or U4214 (N_4214,N_3424,N_2923);
nor U4215 (N_4215,N_3531,N_3502);
nand U4216 (N_4216,N_2783,N_3173);
or U4217 (N_4217,N_3096,N_2914);
nand U4218 (N_4218,N_3019,N_3173);
or U4219 (N_4219,N_2602,N_2608);
or U4220 (N_4220,N_2555,N_2985);
nand U4221 (N_4221,N_2838,N_3454);
nand U4222 (N_4222,N_2676,N_3571);
xnor U4223 (N_4223,N_2636,N_2529);
nand U4224 (N_4224,N_3551,N_2754);
nand U4225 (N_4225,N_3509,N_3339);
nand U4226 (N_4226,N_3592,N_3386);
xor U4227 (N_4227,N_3146,N_2822);
xnor U4228 (N_4228,N_3105,N_3570);
or U4229 (N_4229,N_3580,N_2431);
nor U4230 (N_4230,N_3262,N_2837);
or U4231 (N_4231,N_2628,N_2853);
nand U4232 (N_4232,N_3231,N_2906);
or U4233 (N_4233,N_3541,N_3529);
and U4234 (N_4234,N_2781,N_3208);
nor U4235 (N_4235,N_3536,N_3186);
nor U4236 (N_4236,N_3555,N_3477);
nor U4237 (N_4237,N_2456,N_2555);
and U4238 (N_4238,N_3072,N_3543);
or U4239 (N_4239,N_3492,N_2592);
and U4240 (N_4240,N_2759,N_2873);
or U4241 (N_4241,N_3566,N_2652);
or U4242 (N_4242,N_2959,N_3534);
xnor U4243 (N_4243,N_2940,N_3448);
or U4244 (N_4244,N_3248,N_3101);
nor U4245 (N_4245,N_2628,N_2691);
nand U4246 (N_4246,N_2469,N_2506);
xnor U4247 (N_4247,N_2704,N_2951);
nand U4248 (N_4248,N_3138,N_3144);
and U4249 (N_4249,N_3336,N_2893);
nor U4250 (N_4250,N_3461,N_3453);
xor U4251 (N_4251,N_2976,N_2497);
nor U4252 (N_4252,N_2434,N_2909);
nand U4253 (N_4253,N_2528,N_3428);
nand U4254 (N_4254,N_3553,N_2665);
nor U4255 (N_4255,N_3159,N_2535);
xnor U4256 (N_4256,N_2625,N_2423);
and U4257 (N_4257,N_2788,N_2879);
nor U4258 (N_4258,N_3485,N_2807);
or U4259 (N_4259,N_3479,N_2824);
and U4260 (N_4260,N_3490,N_2962);
nand U4261 (N_4261,N_3151,N_2548);
or U4262 (N_4262,N_3390,N_3243);
xnor U4263 (N_4263,N_2779,N_3080);
xnor U4264 (N_4264,N_3523,N_3361);
or U4265 (N_4265,N_3294,N_2834);
xor U4266 (N_4266,N_3301,N_3317);
or U4267 (N_4267,N_3561,N_3386);
xor U4268 (N_4268,N_3412,N_2465);
nor U4269 (N_4269,N_3267,N_2801);
nor U4270 (N_4270,N_3457,N_3470);
or U4271 (N_4271,N_3359,N_3511);
nor U4272 (N_4272,N_2744,N_2755);
nor U4273 (N_4273,N_2464,N_2413);
and U4274 (N_4274,N_2910,N_3172);
xor U4275 (N_4275,N_2772,N_2960);
nor U4276 (N_4276,N_3540,N_2683);
and U4277 (N_4277,N_2636,N_2774);
and U4278 (N_4278,N_3238,N_2418);
and U4279 (N_4279,N_3126,N_2914);
nand U4280 (N_4280,N_3106,N_2586);
xor U4281 (N_4281,N_3255,N_3354);
xor U4282 (N_4282,N_3569,N_2904);
or U4283 (N_4283,N_2730,N_3200);
or U4284 (N_4284,N_2913,N_2808);
nand U4285 (N_4285,N_3583,N_3132);
or U4286 (N_4286,N_3324,N_2594);
nor U4287 (N_4287,N_3288,N_2447);
xnor U4288 (N_4288,N_2806,N_3453);
nand U4289 (N_4289,N_3541,N_3144);
and U4290 (N_4290,N_3251,N_2432);
xnor U4291 (N_4291,N_3130,N_2971);
or U4292 (N_4292,N_3072,N_3588);
and U4293 (N_4293,N_3215,N_2739);
and U4294 (N_4294,N_2600,N_2848);
xnor U4295 (N_4295,N_3462,N_2615);
nand U4296 (N_4296,N_2561,N_3354);
xnor U4297 (N_4297,N_3572,N_2444);
or U4298 (N_4298,N_2548,N_2793);
nand U4299 (N_4299,N_2783,N_3582);
nand U4300 (N_4300,N_3532,N_2497);
nor U4301 (N_4301,N_3391,N_2772);
or U4302 (N_4302,N_2960,N_2924);
or U4303 (N_4303,N_2749,N_3210);
nor U4304 (N_4304,N_2496,N_2598);
nand U4305 (N_4305,N_2908,N_3038);
and U4306 (N_4306,N_2463,N_3158);
xor U4307 (N_4307,N_3574,N_3169);
or U4308 (N_4308,N_2931,N_3095);
and U4309 (N_4309,N_3383,N_3416);
xor U4310 (N_4310,N_3431,N_3230);
and U4311 (N_4311,N_3434,N_2605);
xor U4312 (N_4312,N_3405,N_3150);
nand U4313 (N_4313,N_3337,N_2684);
nand U4314 (N_4314,N_3337,N_3418);
nand U4315 (N_4315,N_3239,N_3594);
nor U4316 (N_4316,N_3402,N_3069);
xor U4317 (N_4317,N_3278,N_2743);
or U4318 (N_4318,N_3262,N_2966);
nand U4319 (N_4319,N_3451,N_3354);
xnor U4320 (N_4320,N_3597,N_2869);
xnor U4321 (N_4321,N_3360,N_3201);
and U4322 (N_4322,N_2451,N_3101);
xnor U4323 (N_4323,N_2492,N_2705);
nor U4324 (N_4324,N_3355,N_2686);
and U4325 (N_4325,N_2885,N_2666);
nor U4326 (N_4326,N_2645,N_3564);
and U4327 (N_4327,N_2855,N_2921);
nand U4328 (N_4328,N_3582,N_2984);
nand U4329 (N_4329,N_3445,N_3028);
nand U4330 (N_4330,N_2470,N_2541);
nor U4331 (N_4331,N_3367,N_3454);
and U4332 (N_4332,N_3272,N_3340);
xor U4333 (N_4333,N_2535,N_2957);
xnor U4334 (N_4334,N_3376,N_2647);
xor U4335 (N_4335,N_3522,N_2941);
or U4336 (N_4336,N_3565,N_3453);
or U4337 (N_4337,N_3304,N_3233);
nand U4338 (N_4338,N_3458,N_2421);
xnor U4339 (N_4339,N_3103,N_3278);
or U4340 (N_4340,N_3327,N_3426);
xor U4341 (N_4341,N_3259,N_2970);
or U4342 (N_4342,N_3567,N_3160);
nand U4343 (N_4343,N_3462,N_2523);
nand U4344 (N_4344,N_2924,N_3195);
xnor U4345 (N_4345,N_3513,N_3562);
nor U4346 (N_4346,N_2902,N_3245);
and U4347 (N_4347,N_2946,N_3590);
or U4348 (N_4348,N_2680,N_3325);
or U4349 (N_4349,N_3466,N_3160);
nor U4350 (N_4350,N_2534,N_2582);
or U4351 (N_4351,N_2408,N_2739);
nand U4352 (N_4352,N_2427,N_3267);
and U4353 (N_4353,N_3040,N_3104);
nor U4354 (N_4354,N_2948,N_2583);
or U4355 (N_4355,N_2681,N_3510);
xnor U4356 (N_4356,N_2934,N_3531);
nand U4357 (N_4357,N_3407,N_3006);
xnor U4358 (N_4358,N_3255,N_2667);
nor U4359 (N_4359,N_2998,N_3395);
nor U4360 (N_4360,N_3136,N_3558);
xnor U4361 (N_4361,N_3404,N_3229);
nor U4362 (N_4362,N_3219,N_2671);
nor U4363 (N_4363,N_3514,N_3563);
nand U4364 (N_4364,N_2547,N_2558);
xor U4365 (N_4365,N_2739,N_3116);
xnor U4366 (N_4366,N_2732,N_3322);
xor U4367 (N_4367,N_2728,N_3188);
or U4368 (N_4368,N_2527,N_3070);
nor U4369 (N_4369,N_3201,N_3451);
nor U4370 (N_4370,N_2815,N_2534);
and U4371 (N_4371,N_2821,N_2940);
xnor U4372 (N_4372,N_2634,N_2678);
and U4373 (N_4373,N_2872,N_2907);
nor U4374 (N_4374,N_2471,N_3423);
or U4375 (N_4375,N_3004,N_3351);
nand U4376 (N_4376,N_3095,N_3250);
nand U4377 (N_4377,N_3577,N_2422);
or U4378 (N_4378,N_3431,N_3302);
xor U4379 (N_4379,N_3307,N_3227);
nand U4380 (N_4380,N_3237,N_2456);
nor U4381 (N_4381,N_3199,N_3443);
nand U4382 (N_4382,N_2400,N_3020);
nand U4383 (N_4383,N_3006,N_2457);
or U4384 (N_4384,N_2518,N_2621);
or U4385 (N_4385,N_2720,N_2834);
nor U4386 (N_4386,N_3599,N_3322);
or U4387 (N_4387,N_3240,N_2740);
and U4388 (N_4388,N_3255,N_3185);
nor U4389 (N_4389,N_3509,N_2809);
nand U4390 (N_4390,N_3412,N_2833);
nor U4391 (N_4391,N_3267,N_2466);
and U4392 (N_4392,N_2776,N_2857);
xnor U4393 (N_4393,N_2752,N_3526);
nand U4394 (N_4394,N_2649,N_3118);
or U4395 (N_4395,N_3104,N_3391);
xor U4396 (N_4396,N_2672,N_3082);
or U4397 (N_4397,N_2665,N_2800);
and U4398 (N_4398,N_3515,N_2725);
or U4399 (N_4399,N_3571,N_3435);
nor U4400 (N_4400,N_3534,N_3123);
nand U4401 (N_4401,N_2911,N_2411);
xnor U4402 (N_4402,N_2569,N_2826);
xor U4403 (N_4403,N_2438,N_3112);
nor U4404 (N_4404,N_2931,N_3361);
nor U4405 (N_4405,N_2579,N_2704);
and U4406 (N_4406,N_2438,N_2889);
and U4407 (N_4407,N_2891,N_3442);
nand U4408 (N_4408,N_3581,N_3446);
nand U4409 (N_4409,N_3165,N_3413);
nor U4410 (N_4410,N_3541,N_3378);
xor U4411 (N_4411,N_3169,N_2712);
and U4412 (N_4412,N_3347,N_2619);
nor U4413 (N_4413,N_2420,N_2773);
xor U4414 (N_4414,N_2432,N_2498);
and U4415 (N_4415,N_2481,N_2598);
xor U4416 (N_4416,N_3266,N_2995);
or U4417 (N_4417,N_3028,N_2579);
or U4418 (N_4418,N_2534,N_3164);
and U4419 (N_4419,N_2695,N_2953);
or U4420 (N_4420,N_2662,N_3021);
nor U4421 (N_4421,N_2847,N_2831);
nor U4422 (N_4422,N_2809,N_3296);
xnor U4423 (N_4423,N_2486,N_2862);
xor U4424 (N_4424,N_2680,N_3159);
or U4425 (N_4425,N_3184,N_2810);
and U4426 (N_4426,N_2849,N_3414);
xor U4427 (N_4427,N_3538,N_2693);
or U4428 (N_4428,N_2524,N_3595);
nor U4429 (N_4429,N_3137,N_3251);
and U4430 (N_4430,N_2553,N_2649);
and U4431 (N_4431,N_3120,N_2867);
and U4432 (N_4432,N_3519,N_2612);
nand U4433 (N_4433,N_3386,N_3544);
or U4434 (N_4434,N_3574,N_3437);
and U4435 (N_4435,N_2583,N_2998);
and U4436 (N_4436,N_2420,N_2966);
nor U4437 (N_4437,N_3526,N_2577);
xor U4438 (N_4438,N_2762,N_2673);
nor U4439 (N_4439,N_3453,N_2992);
or U4440 (N_4440,N_3595,N_3182);
nand U4441 (N_4441,N_2521,N_2650);
nor U4442 (N_4442,N_3161,N_3014);
nand U4443 (N_4443,N_2976,N_3216);
and U4444 (N_4444,N_3119,N_3012);
or U4445 (N_4445,N_3280,N_3455);
nor U4446 (N_4446,N_3570,N_3290);
nor U4447 (N_4447,N_3009,N_3035);
nand U4448 (N_4448,N_2651,N_3293);
and U4449 (N_4449,N_3225,N_3021);
nor U4450 (N_4450,N_2871,N_2433);
or U4451 (N_4451,N_2799,N_3551);
xor U4452 (N_4452,N_3227,N_3174);
nor U4453 (N_4453,N_2573,N_2807);
nor U4454 (N_4454,N_3375,N_2999);
nor U4455 (N_4455,N_2677,N_3242);
nor U4456 (N_4456,N_2839,N_2575);
and U4457 (N_4457,N_3598,N_3433);
nand U4458 (N_4458,N_3599,N_3550);
nand U4459 (N_4459,N_2675,N_2669);
and U4460 (N_4460,N_3575,N_2942);
nand U4461 (N_4461,N_2847,N_2826);
nor U4462 (N_4462,N_2455,N_2624);
nand U4463 (N_4463,N_3260,N_2421);
nand U4464 (N_4464,N_3409,N_2595);
or U4465 (N_4465,N_3314,N_3062);
xor U4466 (N_4466,N_3181,N_3179);
nand U4467 (N_4467,N_2892,N_3444);
xnor U4468 (N_4468,N_2774,N_2979);
and U4469 (N_4469,N_2511,N_3561);
or U4470 (N_4470,N_3282,N_3068);
or U4471 (N_4471,N_2804,N_3119);
and U4472 (N_4472,N_2687,N_2953);
xnor U4473 (N_4473,N_3076,N_3580);
nor U4474 (N_4474,N_3089,N_3385);
or U4475 (N_4475,N_3522,N_2503);
or U4476 (N_4476,N_3193,N_3557);
and U4477 (N_4477,N_3267,N_2808);
and U4478 (N_4478,N_2587,N_2926);
nand U4479 (N_4479,N_3083,N_3187);
nand U4480 (N_4480,N_2987,N_2567);
or U4481 (N_4481,N_2429,N_2816);
nand U4482 (N_4482,N_3599,N_3077);
or U4483 (N_4483,N_2728,N_2645);
and U4484 (N_4484,N_3109,N_3200);
nand U4485 (N_4485,N_3518,N_2589);
xor U4486 (N_4486,N_2437,N_3054);
or U4487 (N_4487,N_2971,N_3293);
nor U4488 (N_4488,N_2976,N_3560);
or U4489 (N_4489,N_3532,N_2897);
or U4490 (N_4490,N_2465,N_3536);
nand U4491 (N_4491,N_3546,N_3483);
xnor U4492 (N_4492,N_3182,N_2856);
or U4493 (N_4493,N_2417,N_2853);
or U4494 (N_4494,N_2734,N_2660);
nand U4495 (N_4495,N_3383,N_3313);
nor U4496 (N_4496,N_2876,N_3405);
and U4497 (N_4497,N_2965,N_3050);
xnor U4498 (N_4498,N_3259,N_2708);
and U4499 (N_4499,N_3447,N_2435);
xor U4500 (N_4500,N_2616,N_3150);
nor U4501 (N_4501,N_2461,N_2765);
or U4502 (N_4502,N_3263,N_3559);
xnor U4503 (N_4503,N_3041,N_2765);
nand U4504 (N_4504,N_2595,N_3388);
or U4505 (N_4505,N_3208,N_3288);
and U4506 (N_4506,N_3367,N_2777);
or U4507 (N_4507,N_3073,N_2411);
nor U4508 (N_4508,N_3414,N_2838);
nand U4509 (N_4509,N_2830,N_2951);
nor U4510 (N_4510,N_3210,N_3372);
nor U4511 (N_4511,N_3578,N_3581);
nor U4512 (N_4512,N_3513,N_3310);
or U4513 (N_4513,N_3580,N_2694);
nand U4514 (N_4514,N_3200,N_2541);
nor U4515 (N_4515,N_3469,N_2851);
nor U4516 (N_4516,N_3002,N_2925);
and U4517 (N_4517,N_2662,N_2539);
or U4518 (N_4518,N_2408,N_2935);
nor U4519 (N_4519,N_2724,N_2722);
xnor U4520 (N_4520,N_3069,N_2914);
or U4521 (N_4521,N_3408,N_3114);
xnor U4522 (N_4522,N_3347,N_3435);
or U4523 (N_4523,N_2690,N_2750);
and U4524 (N_4524,N_2747,N_3401);
nor U4525 (N_4525,N_2584,N_2887);
xnor U4526 (N_4526,N_3043,N_2657);
and U4527 (N_4527,N_3134,N_2958);
or U4528 (N_4528,N_2963,N_3305);
xor U4529 (N_4529,N_3124,N_3275);
or U4530 (N_4530,N_2537,N_3404);
nand U4531 (N_4531,N_3137,N_3587);
xor U4532 (N_4532,N_2601,N_3011);
nand U4533 (N_4533,N_2805,N_2622);
xor U4534 (N_4534,N_2893,N_3146);
and U4535 (N_4535,N_2635,N_2892);
xor U4536 (N_4536,N_2696,N_2940);
and U4537 (N_4537,N_2698,N_2514);
or U4538 (N_4538,N_2512,N_2780);
nor U4539 (N_4539,N_2914,N_3578);
nor U4540 (N_4540,N_3553,N_2686);
nand U4541 (N_4541,N_2552,N_2782);
nand U4542 (N_4542,N_3465,N_3437);
and U4543 (N_4543,N_3137,N_2856);
nor U4544 (N_4544,N_2652,N_2764);
xnor U4545 (N_4545,N_2505,N_3326);
or U4546 (N_4546,N_3185,N_2796);
xnor U4547 (N_4547,N_2901,N_3087);
nand U4548 (N_4548,N_3282,N_3335);
xor U4549 (N_4549,N_3381,N_2759);
xnor U4550 (N_4550,N_2631,N_3326);
and U4551 (N_4551,N_3404,N_3405);
nand U4552 (N_4552,N_3529,N_3063);
xor U4553 (N_4553,N_3261,N_3543);
nor U4554 (N_4554,N_2496,N_2835);
or U4555 (N_4555,N_3140,N_3385);
nor U4556 (N_4556,N_2603,N_2717);
nor U4557 (N_4557,N_3439,N_2624);
and U4558 (N_4558,N_2878,N_2976);
nand U4559 (N_4559,N_3121,N_3227);
or U4560 (N_4560,N_2508,N_2938);
and U4561 (N_4561,N_3116,N_2893);
nor U4562 (N_4562,N_3475,N_3521);
or U4563 (N_4563,N_2618,N_2565);
nand U4564 (N_4564,N_3349,N_3015);
and U4565 (N_4565,N_3023,N_3437);
nor U4566 (N_4566,N_2460,N_2872);
nand U4567 (N_4567,N_2820,N_3304);
xnor U4568 (N_4568,N_3364,N_3241);
xor U4569 (N_4569,N_2802,N_2513);
nor U4570 (N_4570,N_3155,N_2491);
nor U4571 (N_4571,N_2731,N_3126);
xor U4572 (N_4572,N_3290,N_2500);
and U4573 (N_4573,N_2851,N_2518);
or U4574 (N_4574,N_2714,N_3486);
and U4575 (N_4575,N_3310,N_3496);
nand U4576 (N_4576,N_3546,N_2909);
and U4577 (N_4577,N_2995,N_3278);
xnor U4578 (N_4578,N_3020,N_2946);
and U4579 (N_4579,N_2656,N_3108);
xnor U4580 (N_4580,N_2488,N_2427);
and U4581 (N_4581,N_3216,N_2822);
and U4582 (N_4582,N_3263,N_2891);
or U4583 (N_4583,N_3295,N_3269);
nor U4584 (N_4584,N_2414,N_2512);
and U4585 (N_4585,N_2887,N_2908);
nor U4586 (N_4586,N_3063,N_3272);
xnor U4587 (N_4587,N_2438,N_2713);
and U4588 (N_4588,N_2622,N_2481);
xnor U4589 (N_4589,N_2874,N_3416);
xnor U4590 (N_4590,N_3138,N_2980);
nor U4591 (N_4591,N_2773,N_2548);
nor U4592 (N_4592,N_3385,N_2581);
nor U4593 (N_4593,N_3371,N_2809);
nor U4594 (N_4594,N_3590,N_3179);
nor U4595 (N_4595,N_2594,N_3586);
or U4596 (N_4596,N_3282,N_3571);
xor U4597 (N_4597,N_3033,N_2765);
xor U4598 (N_4598,N_2849,N_3072);
xor U4599 (N_4599,N_2822,N_3161);
xor U4600 (N_4600,N_2825,N_2645);
or U4601 (N_4601,N_2507,N_2898);
nand U4602 (N_4602,N_2914,N_3166);
and U4603 (N_4603,N_3200,N_2499);
nor U4604 (N_4604,N_3597,N_3082);
or U4605 (N_4605,N_2612,N_3084);
and U4606 (N_4606,N_3101,N_3542);
xnor U4607 (N_4607,N_2466,N_3370);
nor U4608 (N_4608,N_2519,N_2626);
or U4609 (N_4609,N_3152,N_3567);
nor U4610 (N_4610,N_3317,N_3148);
nand U4611 (N_4611,N_2886,N_2413);
or U4612 (N_4612,N_3077,N_2658);
nor U4613 (N_4613,N_3434,N_3407);
nor U4614 (N_4614,N_2926,N_3345);
nand U4615 (N_4615,N_2618,N_3239);
xnor U4616 (N_4616,N_3175,N_2600);
nand U4617 (N_4617,N_3118,N_3548);
nand U4618 (N_4618,N_2834,N_2549);
xor U4619 (N_4619,N_2709,N_3467);
nand U4620 (N_4620,N_2463,N_3324);
or U4621 (N_4621,N_2575,N_3125);
nand U4622 (N_4622,N_2978,N_2753);
nand U4623 (N_4623,N_2566,N_3109);
nor U4624 (N_4624,N_2534,N_2822);
nor U4625 (N_4625,N_3356,N_3279);
xor U4626 (N_4626,N_3593,N_2901);
or U4627 (N_4627,N_2567,N_3147);
and U4628 (N_4628,N_3579,N_3455);
and U4629 (N_4629,N_2802,N_3206);
and U4630 (N_4630,N_3579,N_3448);
and U4631 (N_4631,N_2495,N_2429);
xor U4632 (N_4632,N_2706,N_3117);
or U4633 (N_4633,N_2539,N_3056);
nand U4634 (N_4634,N_3284,N_2883);
xor U4635 (N_4635,N_2417,N_2569);
nor U4636 (N_4636,N_2857,N_3356);
and U4637 (N_4637,N_2691,N_3239);
and U4638 (N_4638,N_2447,N_3126);
xnor U4639 (N_4639,N_3471,N_3389);
and U4640 (N_4640,N_2473,N_3419);
or U4641 (N_4641,N_3336,N_2485);
xnor U4642 (N_4642,N_3245,N_2749);
nand U4643 (N_4643,N_2977,N_3413);
xor U4644 (N_4644,N_3036,N_2555);
nor U4645 (N_4645,N_2406,N_3166);
nor U4646 (N_4646,N_2918,N_3062);
nor U4647 (N_4647,N_3563,N_3365);
or U4648 (N_4648,N_3089,N_3544);
nand U4649 (N_4649,N_3459,N_3133);
nand U4650 (N_4650,N_2877,N_2859);
nor U4651 (N_4651,N_3194,N_3043);
and U4652 (N_4652,N_3074,N_3017);
or U4653 (N_4653,N_2669,N_3118);
or U4654 (N_4654,N_3105,N_2725);
nand U4655 (N_4655,N_3115,N_2672);
xnor U4656 (N_4656,N_3497,N_2607);
nand U4657 (N_4657,N_2589,N_3547);
xnor U4658 (N_4658,N_3428,N_3396);
or U4659 (N_4659,N_2737,N_2916);
and U4660 (N_4660,N_3464,N_3200);
and U4661 (N_4661,N_3395,N_2719);
and U4662 (N_4662,N_2731,N_3574);
xnor U4663 (N_4663,N_2638,N_2568);
and U4664 (N_4664,N_3222,N_3316);
and U4665 (N_4665,N_3262,N_2751);
nor U4666 (N_4666,N_2794,N_2986);
nor U4667 (N_4667,N_2546,N_3119);
or U4668 (N_4668,N_3246,N_3547);
or U4669 (N_4669,N_3222,N_2471);
xnor U4670 (N_4670,N_2780,N_3407);
nand U4671 (N_4671,N_3365,N_3259);
and U4672 (N_4672,N_2803,N_2845);
and U4673 (N_4673,N_2915,N_2778);
or U4674 (N_4674,N_2661,N_2570);
and U4675 (N_4675,N_2568,N_3588);
or U4676 (N_4676,N_3545,N_2692);
and U4677 (N_4677,N_3535,N_2762);
or U4678 (N_4678,N_2699,N_2898);
xnor U4679 (N_4679,N_2538,N_3471);
and U4680 (N_4680,N_2632,N_2589);
nor U4681 (N_4681,N_2825,N_3074);
nor U4682 (N_4682,N_3397,N_3134);
and U4683 (N_4683,N_3263,N_3109);
nor U4684 (N_4684,N_3232,N_2803);
and U4685 (N_4685,N_3146,N_2878);
nand U4686 (N_4686,N_3359,N_3535);
or U4687 (N_4687,N_2486,N_2801);
xor U4688 (N_4688,N_2978,N_3554);
xor U4689 (N_4689,N_3439,N_3173);
nand U4690 (N_4690,N_3332,N_3170);
or U4691 (N_4691,N_2961,N_3587);
and U4692 (N_4692,N_2928,N_3239);
or U4693 (N_4693,N_2669,N_3586);
xnor U4694 (N_4694,N_3080,N_3468);
xnor U4695 (N_4695,N_2978,N_2872);
xor U4696 (N_4696,N_2525,N_3430);
and U4697 (N_4697,N_2502,N_2426);
nor U4698 (N_4698,N_2497,N_3301);
nand U4699 (N_4699,N_2478,N_2872);
nand U4700 (N_4700,N_3517,N_2741);
xnor U4701 (N_4701,N_3406,N_3566);
or U4702 (N_4702,N_3434,N_3432);
or U4703 (N_4703,N_2701,N_2952);
nor U4704 (N_4704,N_3547,N_3588);
and U4705 (N_4705,N_2899,N_2791);
or U4706 (N_4706,N_2591,N_2926);
xor U4707 (N_4707,N_3208,N_2569);
nand U4708 (N_4708,N_2492,N_3326);
nor U4709 (N_4709,N_3170,N_2432);
nor U4710 (N_4710,N_3297,N_3227);
xnor U4711 (N_4711,N_3055,N_3093);
nor U4712 (N_4712,N_2455,N_2416);
nor U4713 (N_4713,N_2700,N_2779);
xor U4714 (N_4714,N_3492,N_2687);
xor U4715 (N_4715,N_3385,N_2561);
xnor U4716 (N_4716,N_3284,N_3487);
and U4717 (N_4717,N_2989,N_2781);
or U4718 (N_4718,N_2979,N_3358);
nor U4719 (N_4719,N_3089,N_3162);
nand U4720 (N_4720,N_3167,N_2515);
and U4721 (N_4721,N_3416,N_2419);
xnor U4722 (N_4722,N_2833,N_3200);
or U4723 (N_4723,N_2756,N_2639);
or U4724 (N_4724,N_2863,N_3547);
nor U4725 (N_4725,N_3347,N_3296);
and U4726 (N_4726,N_2413,N_2752);
nor U4727 (N_4727,N_3010,N_2464);
nand U4728 (N_4728,N_3432,N_3205);
xnor U4729 (N_4729,N_3025,N_2989);
or U4730 (N_4730,N_2738,N_2910);
nand U4731 (N_4731,N_3184,N_3434);
nor U4732 (N_4732,N_2593,N_2942);
or U4733 (N_4733,N_2923,N_2800);
xnor U4734 (N_4734,N_3361,N_2593);
or U4735 (N_4735,N_3363,N_2687);
or U4736 (N_4736,N_3293,N_2783);
or U4737 (N_4737,N_2616,N_2486);
or U4738 (N_4738,N_2568,N_2911);
nand U4739 (N_4739,N_2546,N_3069);
or U4740 (N_4740,N_2858,N_2831);
nand U4741 (N_4741,N_3137,N_2657);
xnor U4742 (N_4742,N_3431,N_3033);
and U4743 (N_4743,N_2987,N_2660);
and U4744 (N_4744,N_2555,N_3167);
xor U4745 (N_4745,N_2875,N_3276);
nor U4746 (N_4746,N_2638,N_3574);
xor U4747 (N_4747,N_3203,N_2404);
nor U4748 (N_4748,N_2458,N_2673);
nor U4749 (N_4749,N_3249,N_3236);
nor U4750 (N_4750,N_2879,N_2859);
nor U4751 (N_4751,N_2456,N_3426);
nand U4752 (N_4752,N_3489,N_3381);
xnor U4753 (N_4753,N_3138,N_2557);
nor U4754 (N_4754,N_2653,N_3429);
nand U4755 (N_4755,N_2529,N_2762);
nand U4756 (N_4756,N_2897,N_2498);
nand U4757 (N_4757,N_2909,N_2739);
and U4758 (N_4758,N_3193,N_2855);
or U4759 (N_4759,N_2899,N_2938);
and U4760 (N_4760,N_2404,N_2740);
and U4761 (N_4761,N_2769,N_2594);
xnor U4762 (N_4762,N_2617,N_2499);
nor U4763 (N_4763,N_3348,N_3468);
and U4764 (N_4764,N_3087,N_3353);
and U4765 (N_4765,N_3566,N_2522);
nor U4766 (N_4766,N_2914,N_3531);
or U4767 (N_4767,N_2785,N_2701);
and U4768 (N_4768,N_3211,N_3079);
and U4769 (N_4769,N_3552,N_3161);
and U4770 (N_4770,N_3431,N_3338);
nor U4771 (N_4771,N_2831,N_2990);
nand U4772 (N_4772,N_2476,N_2990);
nand U4773 (N_4773,N_3524,N_3412);
nor U4774 (N_4774,N_3112,N_3273);
or U4775 (N_4775,N_2653,N_2885);
nor U4776 (N_4776,N_3327,N_2546);
nor U4777 (N_4777,N_3289,N_3346);
and U4778 (N_4778,N_3502,N_2976);
xnor U4779 (N_4779,N_3555,N_3237);
and U4780 (N_4780,N_2529,N_2519);
nand U4781 (N_4781,N_3397,N_3130);
xor U4782 (N_4782,N_2565,N_3404);
nor U4783 (N_4783,N_2830,N_3306);
nand U4784 (N_4784,N_3347,N_2572);
and U4785 (N_4785,N_2976,N_3313);
and U4786 (N_4786,N_2725,N_2428);
and U4787 (N_4787,N_3399,N_2814);
nor U4788 (N_4788,N_3241,N_3431);
nor U4789 (N_4789,N_3259,N_3088);
or U4790 (N_4790,N_3261,N_2494);
or U4791 (N_4791,N_2971,N_3005);
and U4792 (N_4792,N_2715,N_3228);
nor U4793 (N_4793,N_3419,N_2933);
nor U4794 (N_4794,N_3041,N_3447);
xnor U4795 (N_4795,N_3014,N_3043);
xnor U4796 (N_4796,N_3174,N_3033);
or U4797 (N_4797,N_2965,N_2742);
nor U4798 (N_4798,N_3093,N_3583);
and U4799 (N_4799,N_3204,N_3371);
xor U4800 (N_4800,N_4240,N_4182);
or U4801 (N_4801,N_4107,N_4367);
nor U4802 (N_4802,N_4102,N_3710);
nand U4803 (N_4803,N_3784,N_3687);
xnor U4804 (N_4804,N_4328,N_4311);
or U4805 (N_4805,N_4478,N_4692);
nor U4806 (N_4806,N_4363,N_4700);
xnor U4807 (N_4807,N_4072,N_3847);
nor U4808 (N_4808,N_4030,N_4390);
or U4809 (N_4809,N_4529,N_4040);
nand U4810 (N_4810,N_4783,N_3898);
nor U4811 (N_4811,N_4320,N_4526);
nor U4812 (N_4812,N_4049,N_4354);
nor U4813 (N_4813,N_4743,N_4649);
nor U4814 (N_4814,N_4680,N_3693);
xnor U4815 (N_4815,N_4042,N_4460);
nor U4816 (N_4816,N_4154,N_3837);
nand U4817 (N_4817,N_4751,N_3826);
nand U4818 (N_4818,N_4343,N_3631);
nand U4819 (N_4819,N_3995,N_3769);
xnor U4820 (N_4820,N_4604,N_3609);
and U4821 (N_4821,N_4357,N_4229);
xor U4822 (N_4822,N_3854,N_3922);
nand U4823 (N_4823,N_4274,N_4114);
and U4824 (N_4824,N_3732,N_4790);
and U4825 (N_4825,N_3997,N_4732);
nor U4826 (N_4826,N_4246,N_4704);
and U4827 (N_4827,N_4200,N_3985);
nor U4828 (N_4828,N_4537,N_4319);
or U4829 (N_4829,N_4546,N_4406);
nand U4830 (N_4830,N_3750,N_3872);
or U4831 (N_4831,N_4148,N_4631);
and U4832 (N_4832,N_4323,N_4186);
and U4833 (N_4833,N_4395,N_4681);
nand U4834 (N_4834,N_4206,N_4738);
nor U4835 (N_4835,N_4192,N_4270);
nor U4836 (N_4836,N_3634,N_3718);
nor U4837 (N_4837,N_4639,N_3856);
nand U4838 (N_4838,N_3917,N_4400);
xor U4839 (N_4839,N_4247,N_4541);
and U4840 (N_4840,N_4257,N_3734);
or U4841 (N_4841,N_4401,N_4022);
or U4842 (N_4842,N_4483,N_3787);
nor U4843 (N_4843,N_3881,N_3741);
nor U4844 (N_4844,N_4497,N_4194);
nor U4845 (N_4845,N_3870,N_4342);
or U4846 (N_4846,N_4686,N_3657);
xor U4847 (N_4847,N_4255,N_4368);
nand U4848 (N_4848,N_4238,N_3941);
nor U4849 (N_4849,N_4446,N_4134);
and U4850 (N_4850,N_3793,N_3629);
nor U4851 (N_4851,N_4643,N_4112);
or U4852 (N_4852,N_4004,N_3675);
nor U4853 (N_4853,N_4178,N_4447);
nand U4854 (N_4854,N_3960,N_4531);
nor U4855 (N_4855,N_4211,N_3803);
xor U4856 (N_4856,N_3866,N_3776);
nand U4857 (N_4857,N_3984,N_4325);
xor U4858 (N_4858,N_4348,N_4669);
xnor U4859 (N_4859,N_3983,N_3933);
and U4860 (N_4860,N_4794,N_4737);
or U4861 (N_4861,N_3999,N_4095);
xor U4862 (N_4862,N_4777,N_4451);
xor U4863 (N_4863,N_4252,N_4745);
xor U4864 (N_4864,N_3831,N_4124);
nor U4865 (N_4865,N_4678,N_4570);
and U4866 (N_4866,N_4027,N_4766);
and U4867 (N_4867,N_3660,N_3619);
and U4868 (N_4868,N_3781,N_4002);
nand U4869 (N_4869,N_3827,N_3825);
nor U4870 (N_4870,N_3664,N_3622);
nor U4871 (N_4871,N_4322,N_4793);
or U4872 (N_4872,N_4286,N_4679);
nand U4873 (N_4873,N_3646,N_4167);
and U4874 (N_4874,N_3773,N_4518);
and U4875 (N_4875,N_3968,N_3939);
or U4876 (N_4876,N_4415,N_4054);
nand U4877 (N_4877,N_3865,N_4550);
nand U4878 (N_4878,N_4025,N_4410);
xnor U4879 (N_4879,N_4340,N_4043);
xnor U4880 (N_4880,N_3877,N_4032);
nand U4881 (N_4881,N_3814,N_3757);
or U4882 (N_4882,N_4315,N_4113);
xnor U4883 (N_4883,N_4553,N_3615);
nand U4884 (N_4884,N_3864,N_4591);
and U4885 (N_4885,N_4509,N_4076);
nor U4886 (N_4886,N_4377,N_3740);
and U4887 (N_4887,N_4207,N_3943);
and U4888 (N_4888,N_4352,N_4157);
xnor U4889 (N_4889,N_3655,N_4662);
nand U4890 (N_4890,N_3681,N_4689);
and U4891 (N_4891,N_4729,N_4621);
and U4892 (N_4892,N_4261,N_4047);
or U4893 (N_4893,N_3860,N_4624);
xnor U4894 (N_4894,N_4472,N_4103);
nor U4895 (N_4895,N_4673,N_4119);
or U4896 (N_4896,N_4058,N_3930);
and U4897 (N_4897,N_4273,N_4302);
and U4898 (N_4898,N_3835,N_3852);
nand U4899 (N_4899,N_3715,N_4771);
or U4900 (N_4900,N_3954,N_4135);
nand U4901 (N_4901,N_4122,N_4228);
xor U4902 (N_4902,N_4608,N_3802);
and U4903 (N_4903,N_4241,N_4272);
xnor U4904 (N_4904,N_4569,N_3915);
nand U4905 (N_4905,N_4575,N_4005);
or U4906 (N_4906,N_3752,N_3706);
nand U4907 (N_4907,N_4219,N_4747);
and U4908 (N_4908,N_3643,N_3709);
or U4909 (N_4909,N_4339,N_4693);
or U4910 (N_4910,N_3962,N_4517);
nand U4911 (N_4911,N_3976,N_3610);
and U4912 (N_4912,N_3952,N_3747);
nor U4913 (N_4913,N_3788,N_4011);
xor U4914 (N_4914,N_3697,N_4660);
and U4915 (N_4915,N_4431,N_4403);
and U4916 (N_4916,N_3958,N_4330);
or U4917 (N_4917,N_3691,N_3978);
xnor U4918 (N_4918,N_4547,N_4007);
nand U4919 (N_4919,N_4374,N_4152);
nand U4920 (N_4920,N_3974,N_4199);
nand U4921 (N_4921,N_3987,N_4699);
nor U4922 (N_4922,N_3830,N_4720);
and U4923 (N_4923,N_4191,N_4379);
or U4924 (N_4924,N_4236,N_4768);
or U4925 (N_4925,N_4503,N_4445);
nand U4926 (N_4926,N_4064,N_4594);
xor U4927 (N_4927,N_4727,N_4079);
and U4928 (N_4928,N_4346,N_4131);
xnor U4929 (N_4929,N_4023,N_3948);
and U4930 (N_4930,N_4414,N_4539);
xor U4931 (N_4931,N_3973,N_4012);
nor U4932 (N_4932,N_4000,N_4017);
nand U4933 (N_4933,N_4232,N_4574);
nand U4934 (N_4934,N_3716,N_3925);
xnor U4935 (N_4935,N_3833,N_4278);
xor U4936 (N_4936,N_3677,N_3867);
nand U4937 (N_4937,N_4237,N_4034);
xnor U4938 (N_4938,N_3703,N_4770);
xnor U4939 (N_4939,N_3820,N_4314);
xnor U4940 (N_4940,N_4335,N_3824);
and U4941 (N_4941,N_4615,N_3671);
nor U4942 (N_4942,N_4016,N_4312);
xor U4943 (N_4943,N_4703,N_4417);
xor U4944 (N_4944,N_3724,N_4773);
xor U4945 (N_4945,N_4317,N_4640);
nand U4946 (N_4946,N_3810,N_3931);
nand U4947 (N_4947,N_4196,N_4694);
and U4948 (N_4948,N_4494,N_4021);
nand U4949 (N_4949,N_4502,N_4069);
nand U4950 (N_4950,N_3994,N_4430);
or U4951 (N_4951,N_4092,N_3882);
and U4952 (N_4952,N_3690,N_3818);
and U4953 (N_4953,N_3971,N_4398);
xnor U4954 (N_4954,N_4600,N_3908);
xnor U4955 (N_4955,N_4622,N_3678);
nor U4956 (N_4956,N_4426,N_3606);
nor U4957 (N_4957,N_3947,N_4653);
and U4958 (N_4958,N_4056,N_3990);
and U4959 (N_4959,N_3808,N_4209);
or U4960 (N_4960,N_3726,N_3604);
xor U4961 (N_4961,N_4077,N_4256);
xor U4962 (N_4962,N_4656,N_4293);
nand U4963 (N_4963,N_4501,N_4099);
nor U4964 (N_4964,N_4698,N_3725);
or U4965 (N_4965,N_4612,N_4180);
nand U4966 (N_4966,N_3673,N_4650);
nor U4967 (N_4967,N_3696,N_3910);
and U4968 (N_4968,N_4630,N_3745);
and U4969 (N_4969,N_4545,N_4020);
or U4970 (N_4970,N_4746,N_4036);
or U4971 (N_4971,N_4670,N_3886);
or U4972 (N_4972,N_3923,N_4279);
xnor U4973 (N_4973,N_4506,N_3654);
nor U4974 (N_4974,N_3907,N_4602);
xnor U4975 (N_4975,N_4087,N_4037);
and U4976 (N_4976,N_4397,N_3708);
nor U4977 (N_4977,N_3955,N_4225);
xnor U4978 (N_4978,N_4577,N_4373);
nand U4979 (N_4979,N_4111,N_4475);
and U4980 (N_4980,N_4734,N_4128);
nand U4981 (N_4981,N_3961,N_3705);
or U4982 (N_4982,N_3938,N_3763);
nor U4983 (N_4983,N_3937,N_4776);
xnor U4984 (N_4984,N_4333,N_4583);
nor U4985 (N_4985,N_4419,N_4633);
nand U4986 (N_4986,N_4175,N_4696);
xor U4987 (N_4987,N_4587,N_4461);
nor U4988 (N_4988,N_4068,N_4781);
xor U4989 (N_4989,N_4231,N_3662);
or U4990 (N_4990,N_3875,N_4318);
nor U4991 (N_4991,N_4603,N_3775);
or U4992 (N_4992,N_4080,N_3861);
xor U4993 (N_4993,N_4418,N_3707);
nand U4994 (N_4994,N_3608,N_3729);
nand U4995 (N_4995,N_3642,N_4364);
and U4996 (N_4996,N_4589,N_3772);
nor U4997 (N_4997,N_4074,N_4722);
nand U4998 (N_4998,N_3892,N_4299);
nand U4999 (N_4999,N_4062,N_4730);
nor U5000 (N_5000,N_3765,N_4070);
nor U5001 (N_5001,N_4285,N_4636);
nor U5002 (N_5002,N_4691,N_4227);
or U5003 (N_5003,N_3602,N_3921);
nand U5004 (N_5004,N_4504,N_3627);
nor U5005 (N_5005,N_3653,N_4712);
xor U5006 (N_5006,N_3884,N_4792);
xnor U5007 (N_5007,N_4752,N_4565);
nand U5008 (N_5008,N_3628,N_4090);
xor U5009 (N_5009,N_3695,N_4083);
nor U5010 (N_5010,N_4297,N_4146);
and U5011 (N_5011,N_4533,N_3644);
xnor U5012 (N_5012,N_4337,N_4276);
xor U5013 (N_5013,N_4761,N_4088);
xor U5014 (N_5014,N_3766,N_4571);
nor U5015 (N_5015,N_3737,N_4300);
xnor U5016 (N_5016,N_3887,N_3603);
nand U5017 (N_5017,N_3713,N_4728);
xor U5018 (N_5018,N_4439,N_4269);
and U5019 (N_5019,N_3748,N_4165);
or U5020 (N_5020,N_3893,N_4674);
xnor U5021 (N_5021,N_4404,N_4138);
nor U5022 (N_5022,N_4581,N_4310);
nor U5023 (N_5023,N_4166,N_4073);
xnor U5024 (N_5024,N_4201,N_3640);
and U5025 (N_5025,N_4251,N_3848);
nand U5026 (N_5026,N_3876,N_4380);
or U5027 (N_5027,N_3945,N_4651);
nand U5028 (N_5028,N_3899,N_4671);
xnor U5029 (N_5029,N_3873,N_4632);
nor U5030 (N_5030,N_3620,N_4427);
xor U5031 (N_5031,N_3767,N_4489);
nand U5032 (N_5032,N_3813,N_4764);
nor U5033 (N_5033,N_4634,N_3844);
nand U5034 (N_5034,N_4006,N_4029);
and U5035 (N_5035,N_4234,N_4324);
or U5036 (N_5036,N_4564,N_4492);
or U5037 (N_5037,N_4481,N_4283);
nand U5038 (N_5038,N_4024,N_4215);
nand U5039 (N_5039,N_3746,N_4378);
xnor U5040 (N_5040,N_4376,N_4051);
or U5041 (N_5041,N_3819,N_4797);
or U5042 (N_5042,N_3680,N_3953);
nand U5043 (N_5043,N_3723,N_4567);
and U5044 (N_5044,N_3699,N_4421);
xnor U5045 (N_5045,N_3863,N_3704);
xnor U5046 (N_5046,N_4697,N_4249);
xor U5047 (N_5047,N_4579,N_4578);
nor U5048 (N_5048,N_4353,N_4218);
or U5049 (N_5049,N_4303,N_4795);
nor U5050 (N_5050,N_4733,N_4641);
and U5051 (N_5051,N_3674,N_3883);
xor U5052 (N_5052,N_4384,N_4668);
nor U5053 (N_5053,N_4396,N_4635);
nor U5054 (N_5054,N_3749,N_4785);
nor U5055 (N_5055,N_4125,N_4658);
nand U5056 (N_5056,N_3849,N_3714);
nor U5057 (N_5057,N_3770,N_3730);
nand U5058 (N_5058,N_4476,N_3601);
nand U5059 (N_5059,N_3946,N_4026);
and U5060 (N_5060,N_4149,N_4361);
nor U5061 (N_5061,N_3834,N_4362);
xnor U5062 (N_5062,N_4144,N_4520);
xnor U5063 (N_5063,N_4391,N_4637);
or U5064 (N_5064,N_3742,N_3889);
nand U5065 (N_5065,N_4796,N_3649);
xor U5066 (N_5066,N_4477,N_4757);
nor U5067 (N_5067,N_3896,N_4100);
or U5068 (N_5068,N_3845,N_4713);
nor U5069 (N_5069,N_4061,N_3659);
and U5070 (N_5070,N_4437,N_4078);
nor U5071 (N_5071,N_4326,N_4726);
nand U5072 (N_5072,N_4126,N_3841);
nor U5073 (N_5073,N_4760,N_4242);
xnor U5074 (N_5074,N_3846,N_4652);
nand U5075 (N_5075,N_3605,N_4482);
nand U5076 (N_5076,N_3638,N_3991);
nand U5077 (N_5077,N_3904,N_4347);
or U5078 (N_5078,N_4055,N_4763);
nor U5079 (N_5079,N_4267,N_3840);
nand U5080 (N_5080,N_4749,N_4663);
nor U5081 (N_5081,N_3721,N_4627);
nand U5082 (N_5082,N_4514,N_4153);
and U5083 (N_5083,N_4221,N_4185);
and U5084 (N_5084,N_4556,N_4243);
nor U5085 (N_5085,N_4585,N_4101);
or U5086 (N_5086,N_4519,N_3782);
nand U5087 (N_5087,N_4405,N_4588);
or U5088 (N_5088,N_3927,N_4177);
and U5089 (N_5089,N_4687,N_4171);
nor U5090 (N_5090,N_3758,N_4540);
xnor U5091 (N_5091,N_4160,N_4505);
nor U5092 (N_5092,N_4287,N_4499);
nand U5093 (N_5093,N_4308,N_4508);
nor U5094 (N_5094,N_3735,N_4093);
xnor U5095 (N_5095,N_4108,N_4572);
and U5096 (N_5096,N_4375,N_4132);
and U5097 (N_5097,N_4609,N_3905);
or U5098 (N_5098,N_4204,N_4458);
xnor U5099 (N_5099,N_4513,N_4336);
nand U5100 (N_5100,N_4140,N_4263);
nor U5101 (N_5101,N_4762,N_4690);
and U5102 (N_5102,N_4266,N_3698);
or U5103 (N_5103,N_4466,N_4717);
nand U5104 (N_5104,N_4592,N_4098);
nor U5105 (N_5105,N_4222,N_4515);
or U5106 (N_5106,N_4511,N_4423);
nand U5107 (N_5107,N_4253,N_4601);
nand U5108 (N_5108,N_4035,N_4031);
nand U5109 (N_5109,N_4409,N_4360);
and U5110 (N_5110,N_3617,N_4695);
xnor U5111 (N_5111,N_3645,N_3868);
or U5112 (N_5112,N_3795,N_4216);
or U5113 (N_5113,N_4118,N_3993);
or U5114 (N_5114,N_4151,N_3981);
or U5115 (N_5115,N_4628,N_4018);
nor U5116 (N_5116,N_4522,N_4536);
nand U5117 (N_5117,N_3975,N_4089);
or U5118 (N_5118,N_3701,N_4611);
xor U5119 (N_5119,N_4224,N_4289);
and U5120 (N_5120,N_4561,N_3618);
nor U5121 (N_5121,N_4724,N_4606);
or U5122 (N_5122,N_3839,N_4782);
nand U5123 (N_5123,N_4718,N_4758);
nand U5124 (N_5124,N_3685,N_4065);
nand U5125 (N_5125,N_4332,N_4557);
nor U5126 (N_5126,N_3966,N_4413);
or U5127 (N_5127,N_4524,N_3760);
or U5128 (N_5128,N_4424,N_4702);
xor U5129 (N_5129,N_4682,N_4063);
and U5130 (N_5130,N_3901,N_3719);
nand U5131 (N_5131,N_4428,N_4321);
nor U5132 (N_5132,N_4210,N_4468);
xnor U5133 (N_5133,N_4542,N_3928);
nor U5134 (N_5134,N_4655,N_4597);
or U5135 (N_5135,N_4184,N_4009);
nand U5136 (N_5136,N_3891,N_4248);
or U5137 (N_5137,N_4471,N_4527);
and U5138 (N_5138,N_3720,N_4711);
xnor U5139 (N_5139,N_4052,N_4137);
xor U5140 (N_5140,N_4740,N_3843);
nand U5141 (N_5141,N_4217,N_3989);
xor U5142 (N_5142,N_4675,N_4168);
nor U5143 (N_5143,N_4731,N_4551);
nand U5144 (N_5144,N_3815,N_4203);
nand U5145 (N_5145,N_3733,N_4264);
nand U5146 (N_5146,N_4493,N_3736);
nor U5147 (N_5147,N_4644,N_4331);
and U5148 (N_5148,N_3669,N_3979);
xnor U5149 (N_5149,N_4189,N_4774);
and U5150 (N_5150,N_4143,N_3790);
and U5151 (N_5151,N_4350,N_4523);
nor U5152 (N_5152,N_4369,N_3918);
xnor U5153 (N_5153,N_3779,N_4590);
xnor U5154 (N_5154,N_4123,N_4484);
or U5155 (N_5155,N_4059,N_4701);
nor U5156 (N_5156,N_3679,N_3702);
and U5157 (N_5157,N_4094,N_4429);
nand U5158 (N_5158,N_3666,N_3625);
xor U5159 (N_5159,N_3959,N_4019);
or U5160 (N_5160,N_3822,N_3647);
and U5161 (N_5161,N_3878,N_4787);
or U5162 (N_5162,N_4530,N_4725);
nor U5163 (N_5163,N_4453,N_4096);
or U5164 (N_5164,N_3754,N_4327);
nand U5165 (N_5165,N_3641,N_3700);
xor U5166 (N_5166,N_4646,N_3780);
nor U5167 (N_5167,N_3909,N_3836);
nor U5168 (N_5168,N_4085,N_4488);
xnor U5169 (N_5169,N_4086,N_4195);
or U5170 (N_5170,N_3712,N_4586);
nand U5171 (N_5171,N_3850,N_4183);
nand U5172 (N_5172,N_4613,N_4127);
or U5173 (N_5173,N_3851,N_4197);
xor U5174 (N_5174,N_4685,N_4387);
or U5175 (N_5175,N_4459,N_4463);
xor U5176 (N_5176,N_4371,N_3751);
xor U5177 (N_5177,N_3753,N_4109);
xnor U5178 (N_5178,N_3874,N_4498);
or U5179 (N_5179,N_4097,N_4647);
nand U5180 (N_5180,N_3636,N_4338);
or U5181 (N_5181,N_4039,N_4765);
nor U5182 (N_5182,N_4791,N_3762);
or U5183 (N_5183,N_4316,N_4136);
xor U5184 (N_5184,N_4365,N_3940);
xnor U5185 (N_5185,N_4239,N_4543);
or U5186 (N_5186,N_4778,N_4296);
and U5187 (N_5187,N_3935,N_3963);
and U5188 (N_5188,N_4392,N_4355);
xnor U5189 (N_5189,N_3650,N_4133);
and U5190 (N_5190,N_4281,N_4081);
and U5191 (N_5191,N_4438,N_4449);
xor U5192 (N_5192,N_3684,N_4610);
xor U5193 (N_5193,N_4435,N_4301);
xnor U5194 (N_5194,N_3805,N_3964);
xor U5195 (N_5195,N_4748,N_4573);
and U5196 (N_5196,N_3688,N_4198);
xnor U5197 (N_5197,N_4174,N_4349);
or U5198 (N_5198,N_4576,N_4496);
xor U5199 (N_5199,N_4491,N_4708);
and U5200 (N_5200,N_3607,N_4465);
xor U5201 (N_5201,N_4455,N_4220);
or U5202 (N_5202,N_3624,N_4104);
and U5203 (N_5203,N_3743,N_4528);
and U5204 (N_5204,N_4190,N_4667);
or U5205 (N_5205,N_4659,N_4290);
nand U5206 (N_5206,N_4188,N_4046);
and U5207 (N_5207,N_4179,N_4170);
and U5208 (N_5208,N_3906,N_4193);
nor U5209 (N_5209,N_4159,N_4510);
nor U5210 (N_5210,N_3686,N_4334);
nand U5211 (N_5211,N_4741,N_4436);
nor U5212 (N_5212,N_3663,N_4495);
or U5213 (N_5213,N_3900,N_4014);
nand U5214 (N_5214,N_3774,N_4623);
and U5215 (N_5215,N_4010,N_4657);
xnor U5216 (N_5216,N_4735,N_4282);
nand U5217 (N_5217,N_4677,N_4554);
nor U5218 (N_5218,N_3785,N_4386);
nand U5219 (N_5219,N_3894,N_4723);
nor U5220 (N_5220,N_3949,N_3853);
or U5221 (N_5221,N_3982,N_4779);
and U5222 (N_5222,N_4648,N_4142);
and U5223 (N_5223,N_3934,N_4329);
nor U5224 (N_5224,N_3652,N_3916);
xor U5225 (N_5225,N_3902,N_4277);
and U5226 (N_5226,N_4305,N_4756);
nand U5227 (N_5227,N_4291,N_4259);
nand U5228 (N_5228,N_4145,N_4558);
xor U5229 (N_5229,N_4532,N_4434);
nor U5230 (N_5230,N_3616,N_3656);
xnor U5231 (N_5231,N_3897,N_3717);
and U5232 (N_5232,N_3890,N_3986);
nand U5233 (N_5233,N_4467,N_4448);
xnor U5234 (N_5234,N_3727,N_3744);
or U5235 (N_5235,N_4619,N_4599);
nand U5236 (N_5236,N_4075,N_3972);
xor U5237 (N_5237,N_4372,N_4208);
xor U5238 (N_5238,N_3838,N_4306);
and U5239 (N_5239,N_3911,N_4754);
nor U5240 (N_5240,N_3777,N_3689);
xor U5241 (N_5241,N_4440,N_4008);
xnor U5242 (N_5242,N_4433,N_3639);
xor U5243 (N_5243,N_4706,N_3614);
nand U5244 (N_5244,N_4607,N_4202);
or U5245 (N_5245,N_4470,N_4469);
nor U5246 (N_5246,N_4120,N_4304);
and U5247 (N_5247,N_4041,N_3880);
nand U5248 (N_5248,N_3665,N_3670);
nand U5249 (N_5249,N_3977,N_4714);
or U5250 (N_5250,N_4715,N_3842);
xnor U5251 (N_5251,N_4750,N_4512);
and U5252 (N_5252,N_4780,N_4626);
and U5253 (N_5253,N_4244,N_4265);
nor U5254 (N_5254,N_3621,N_4568);
or U5255 (N_5255,N_3816,N_3957);
or U5256 (N_5256,N_4214,N_4566);
or U5257 (N_5257,N_4130,N_3791);
nand U5258 (N_5258,N_4672,N_3600);
xor U5259 (N_5259,N_4262,N_4485);
xor U5260 (N_5260,N_3632,N_3885);
and U5261 (N_5261,N_4212,N_4716);
and U5262 (N_5262,N_3912,N_3817);
nand U5263 (N_5263,N_4060,N_3661);
nand U5264 (N_5264,N_4705,N_4163);
and U5265 (N_5265,N_3648,N_4038);
xor U5266 (N_5266,N_4742,N_4638);
nor U5267 (N_5267,N_4596,N_3832);
and U5268 (N_5268,N_3821,N_4593);
nand U5269 (N_5269,N_3823,N_4538);
and U5270 (N_5270,N_4187,N_4629);
xnor U5271 (N_5271,N_3778,N_3764);
xor U5272 (N_5272,N_4260,N_4158);
nor U5273 (N_5273,N_3728,N_4625);
xnor U5274 (N_5274,N_4233,N_4066);
nor U5275 (N_5275,N_3768,N_4798);
and U5276 (N_5276,N_3800,N_4559);
nand U5277 (N_5277,N_4176,N_4753);
and U5278 (N_5278,N_3859,N_3920);
nand U5279 (N_5279,N_4388,N_3967);
nand U5280 (N_5280,N_4688,N_3761);
nand U5281 (N_5281,N_4412,N_3903);
or U5282 (N_5282,N_4474,N_3924);
nand U5283 (N_5283,N_4110,N_3711);
nor U5284 (N_5284,N_3626,N_3858);
and U5285 (N_5285,N_4788,N_4454);
nand U5286 (N_5286,N_3857,N_3792);
nor U5287 (N_5287,N_4271,N_3739);
nand U5288 (N_5288,N_3786,N_4755);
xor U5289 (N_5289,N_4420,N_4050);
xor U5290 (N_5290,N_4617,N_4254);
xnor U5291 (N_5291,N_4172,N_3692);
nand U5292 (N_5292,N_4560,N_3828);
xnor U5293 (N_5293,N_4767,N_4359);
and U5294 (N_5294,N_3996,N_3970);
or U5295 (N_5295,N_4358,N_4444);
nand U5296 (N_5296,N_4181,N_4719);
or U5297 (N_5297,N_4684,N_4710);
and U5298 (N_5298,N_4356,N_4275);
and U5299 (N_5299,N_4389,N_3998);
and U5300 (N_5300,N_3797,N_4053);
nand U5301 (N_5301,N_4205,N_4250);
nand U5302 (N_5302,N_3623,N_4598);
nand U5303 (N_5303,N_4786,N_4150);
nor U5304 (N_5304,N_4676,N_4161);
xor U5305 (N_5305,N_3879,N_4769);
nor U5306 (N_5306,N_3919,N_4345);
nor U5307 (N_5307,N_4307,N_4155);
xnor U5308 (N_5308,N_4443,N_4408);
or U5309 (N_5309,N_4156,N_3694);
xor U5310 (N_5310,N_4230,N_4759);
nor U5311 (N_5311,N_4548,N_4245);
or U5312 (N_5312,N_3630,N_4048);
nand U5313 (N_5313,N_4487,N_4411);
nand U5314 (N_5314,N_3676,N_3658);
xnor U5315 (N_5315,N_3738,N_3635);
or U5316 (N_5316,N_4162,N_4344);
xor U5317 (N_5317,N_4584,N_4393);
nand U5318 (N_5318,N_3862,N_3951);
or U5319 (N_5319,N_3801,N_4616);
and U5320 (N_5320,N_4683,N_4618);
nor U5321 (N_5321,N_4642,N_4665);
or U5322 (N_5322,N_3799,N_4534);
nand U5323 (N_5323,N_4366,N_3913);
and U5324 (N_5324,N_4084,N_4516);
nor U5325 (N_5325,N_4500,N_4544);
nand U5326 (N_5326,N_4736,N_3804);
nor U5327 (N_5327,N_4169,N_4223);
xor U5328 (N_5328,N_4394,N_4549);
nor U5329 (N_5329,N_4666,N_3936);
nand U5330 (N_5330,N_4525,N_4407);
nor U5331 (N_5331,N_4457,N_4507);
and U5332 (N_5332,N_3722,N_3992);
nand U5333 (N_5333,N_4402,N_4121);
and U5334 (N_5334,N_4268,N_3871);
or U5335 (N_5335,N_3855,N_4129);
or U5336 (N_5336,N_4091,N_4288);
and U5337 (N_5337,N_4664,N_4789);
nand U5338 (N_5338,N_3944,N_4654);
and U5339 (N_5339,N_4399,N_4226);
and U5340 (N_5340,N_4370,N_3755);
nor U5341 (N_5341,N_3829,N_4452);
nand U5342 (N_5342,N_3956,N_3965);
or U5343 (N_5343,N_4721,N_4744);
or U5344 (N_5344,N_4709,N_4456);
nand U5345 (N_5345,N_4645,N_4521);
xnor U5346 (N_5346,N_4284,N_4555);
and U5347 (N_5347,N_3672,N_3756);
xor U5348 (N_5348,N_3969,N_3929);
xor U5349 (N_5349,N_4425,N_4535);
and U5350 (N_5350,N_4450,N_4441);
xnor U5351 (N_5351,N_3783,N_3869);
xnor U5352 (N_5352,N_4385,N_3812);
and U5353 (N_5353,N_3950,N_4001);
or U5354 (N_5354,N_3942,N_4147);
or U5355 (N_5355,N_4595,N_4552);
or U5356 (N_5356,N_4473,N_4381);
and U5357 (N_5357,N_4003,N_4480);
and U5358 (N_5358,N_3914,N_4115);
xnor U5359 (N_5359,N_4082,N_4105);
nand U5360 (N_5360,N_4139,N_4775);
and U5361 (N_5361,N_4117,N_3759);
nand U5362 (N_5362,N_3794,N_4071);
nor U5363 (N_5363,N_4116,N_4422);
and U5364 (N_5364,N_4141,N_3789);
or U5365 (N_5365,N_4490,N_4614);
nor U5366 (N_5366,N_4309,N_4620);
and U5367 (N_5367,N_4235,N_4341);
or U5368 (N_5368,N_3796,N_4280);
xor U5369 (N_5369,N_4313,N_3668);
xor U5370 (N_5370,N_4295,N_4033);
or U5371 (N_5371,N_4173,N_4563);
and U5372 (N_5372,N_3807,N_3651);
nand U5373 (N_5373,N_4562,N_4707);
nand U5374 (N_5374,N_4772,N_4045);
nor U5375 (N_5375,N_4028,N_3798);
xor U5376 (N_5376,N_4294,N_4383);
or U5377 (N_5377,N_3612,N_4013);
xor U5378 (N_5378,N_3637,N_4661);
and U5379 (N_5379,N_3683,N_3667);
and U5380 (N_5380,N_3806,N_3895);
xor U5381 (N_5381,N_4442,N_4015);
or U5382 (N_5382,N_4432,N_4739);
nand U5383 (N_5383,N_4258,N_4486);
and U5384 (N_5384,N_4292,N_4298);
xor U5385 (N_5385,N_3926,N_3809);
nand U5386 (N_5386,N_4044,N_4799);
nor U5387 (N_5387,N_3932,N_4057);
nand U5388 (N_5388,N_4464,N_3613);
nor U5389 (N_5389,N_4784,N_4479);
nand U5390 (N_5390,N_4351,N_3682);
nand U5391 (N_5391,N_4382,N_3988);
or U5392 (N_5392,N_3888,N_4416);
xor U5393 (N_5393,N_3771,N_4462);
or U5394 (N_5394,N_3811,N_4067);
or U5395 (N_5395,N_4106,N_3980);
nor U5396 (N_5396,N_4605,N_4580);
xnor U5397 (N_5397,N_3611,N_4213);
and U5398 (N_5398,N_4582,N_3633);
nand U5399 (N_5399,N_3731,N_4164);
xor U5400 (N_5400,N_4421,N_4253);
xnor U5401 (N_5401,N_4533,N_3651);
and U5402 (N_5402,N_4079,N_4203);
or U5403 (N_5403,N_4468,N_3667);
xnor U5404 (N_5404,N_3627,N_4176);
and U5405 (N_5405,N_3850,N_4205);
xor U5406 (N_5406,N_4696,N_4451);
or U5407 (N_5407,N_3726,N_4156);
or U5408 (N_5408,N_4424,N_4633);
or U5409 (N_5409,N_3788,N_4009);
xnor U5410 (N_5410,N_3692,N_4339);
or U5411 (N_5411,N_3850,N_4418);
xnor U5412 (N_5412,N_4715,N_4307);
nor U5413 (N_5413,N_4274,N_4128);
xor U5414 (N_5414,N_4712,N_4208);
nor U5415 (N_5415,N_4679,N_4696);
or U5416 (N_5416,N_4544,N_4162);
nor U5417 (N_5417,N_3921,N_3756);
and U5418 (N_5418,N_3681,N_4570);
and U5419 (N_5419,N_3946,N_4533);
xor U5420 (N_5420,N_4395,N_4187);
and U5421 (N_5421,N_4215,N_4014);
or U5422 (N_5422,N_4318,N_4779);
nor U5423 (N_5423,N_3700,N_3830);
or U5424 (N_5424,N_4792,N_4619);
xor U5425 (N_5425,N_4397,N_4070);
xor U5426 (N_5426,N_4243,N_4112);
nand U5427 (N_5427,N_4576,N_4299);
nor U5428 (N_5428,N_3813,N_4052);
and U5429 (N_5429,N_4030,N_4336);
or U5430 (N_5430,N_4536,N_4566);
and U5431 (N_5431,N_3984,N_3972);
or U5432 (N_5432,N_4201,N_3696);
nand U5433 (N_5433,N_3810,N_4315);
or U5434 (N_5434,N_4241,N_3875);
or U5435 (N_5435,N_4797,N_4264);
nor U5436 (N_5436,N_4086,N_4550);
nand U5437 (N_5437,N_4725,N_4033);
nor U5438 (N_5438,N_4411,N_4372);
and U5439 (N_5439,N_4243,N_4799);
xnor U5440 (N_5440,N_4404,N_3712);
nand U5441 (N_5441,N_3905,N_4284);
and U5442 (N_5442,N_4232,N_4156);
xor U5443 (N_5443,N_4242,N_4534);
or U5444 (N_5444,N_4532,N_4628);
and U5445 (N_5445,N_4083,N_3620);
nor U5446 (N_5446,N_4658,N_3964);
or U5447 (N_5447,N_4214,N_3796);
xnor U5448 (N_5448,N_4169,N_4707);
nand U5449 (N_5449,N_3647,N_4326);
xor U5450 (N_5450,N_4358,N_4560);
nand U5451 (N_5451,N_4521,N_3943);
nand U5452 (N_5452,N_3870,N_4103);
xor U5453 (N_5453,N_4215,N_4733);
nor U5454 (N_5454,N_4550,N_3640);
xnor U5455 (N_5455,N_3853,N_3729);
or U5456 (N_5456,N_4700,N_4240);
nor U5457 (N_5457,N_4416,N_4007);
or U5458 (N_5458,N_4339,N_4690);
or U5459 (N_5459,N_4005,N_4663);
or U5460 (N_5460,N_4205,N_4751);
or U5461 (N_5461,N_3770,N_4676);
nand U5462 (N_5462,N_3894,N_3673);
or U5463 (N_5463,N_4036,N_3707);
and U5464 (N_5464,N_4690,N_3611);
xnor U5465 (N_5465,N_4107,N_3892);
nor U5466 (N_5466,N_4021,N_4390);
or U5467 (N_5467,N_3871,N_3683);
or U5468 (N_5468,N_3778,N_4755);
nand U5469 (N_5469,N_3989,N_3766);
nor U5470 (N_5470,N_3756,N_3659);
xor U5471 (N_5471,N_4780,N_4264);
xor U5472 (N_5472,N_4275,N_3677);
nand U5473 (N_5473,N_4151,N_4267);
and U5474 (N_5474,N_3894,N_4157);
nor U5475 (N_5475,N_4028,N_4342);
xor U5476 (N_5476,N_3657,N_4025);
nor U5477 (N_5477,N_3615,N_4557);
xor U5478 (N_5478,N_4657,N_3641);
nor U5479 (N_5479,N_4108,N_4318);
nor U5480 (N_5480,N_4763,N_4488);
nor U5481 (N_5481,N_4756,N_4047);
or U5482 (N_5482,N_4152,N_4348);
xnor U5483 (N_5483,N_4527,N_3666);
or U5484 (N_5484,N_4459,N_4433);
nor U5485 (N_5485,N_4036,N_4427);
nand U5486 (N_5486,N_3635,N_4644);
and U5487 (N_5487,N_4072,N_4699);
xor U5488 (N_5488,N_4447,N_4086);
xor U5489 (N_5489,N_4255,N_4244);
or U5490 (N_5490,N_3603,N_4018);
xnor U5491 (N_5491,N_4625,N_4556);
nor U5492 (N_5492,N_3819,N_4389);
nor U5493 (N_5493,N_4194,N_4761);
nor U5494 (N_5494,N_4053,N_4109);
nor U5495 (N_5495,N_3863,N_4510);
and U5496 (N_5496,N_4752,N_4390);
nand U5497 (N_5497,N_4423,N_4004);
and U5498 (N_5498,N_4711,N_3636);
or U5499 (N_5499,N_4093,N_4063);
nand U5500 (N_5500,N_4091,N_4499);
nor U5501 (N_5501,N_4756,N_4475);
and U5502 (N_5502,N_4700,N_3952);
or U5503 (N_5503,N_3941,N_4522);
xor U5504 (N_5504,N_3961,N_4242);
or U5505 (N_5505,N_4623,N_4492);
nand U5506 (N_5506,N_4111,N_4461);
nor U5507 (N_5507,N_3796,N_4101);
and U5508 (N_5508,N_4712,N_3799);
and U5509 (N_5509,N_4353,N_4639);
xnor U5510 (N_5510,N_4442,N_3928);
or U5511 (N_5511,N_4784,N_4592);
xnor U5512 (N_5512,N_4690,N_3718);
or U5513 (N_5513,N_4498,N_3955);
nand U5514 (N_5514,N_4733,N_4317);
and U5515 (N_5515,N_4413,N_4158);
or U5516 (N_5516,N_4004,N_4249);
nor U5517 (N_5517,N_4185,N_3733);
nand U5518 (N_5518,N_4514,N_3775);
nand U5519 (N_5519,N_4744,N_4118);
and U5520 (N_5520,N_4142,N_4677);
and U5521 (N_5521,N_4297,N_4755);
nor U5522 (N_5522,N_4539,N_3685);
and U5523 (N_5523,N_4522,N_4149);
or U5524 (N_5524,N_4218,N_4203);
nor U5525 (N_5525,N_3887,N_4274);
nor U5526 (N_5526,N_3668,N_4353);
nor U5527 (N_5527,N_4113,N_4053);
xor U5528 (N_5528,N_4260,N_3870);
and U5529 (N_5529,N_3836,N_4304);
nor U5530 (N_5530,N_4008,N_4749);
or U5531 (N_5531,N_3760,N_4082);
and U5532 (N_5532,N_4523,N_4752);
and U5533 (N_5533,N_4106,N_4587);
nor U5534 (N_5534,N_3890,N_4343);
or U5535 (N_5535,N_4457,N_4021);
and U5536 (N_5536,N_4106,N_3626);
nand U5537 (N_5537,N_3789,N_3682);
or U5538 (N_5538,N_3828,N_4588);
xor U5539 (N_5539,N_4382,N_4248);
and U5540 (N_5540,N_4084,N_4748);
or U5541 (N_5541,N_4371,N_3866);
nor U5542 (N_5542,N_4741,N_4052);
nor U5543 (N_5543,N_4207,N_4707);
xnor U5544 (N_5544,N_4294,N_4663);
xor U5545 (N_5545,N_4356,N_3642);
and U5546 (N_5546,N_4433,N_3688);
or U5547 (N_5547,N_4045,N_3820);
nor U5548 (N_5548,N_3618,N_3896);
or U5549 (N_5549,N_3831,N_4493);
nand U5550 (N_5550,N_3847,N_4561);
or U5551 (N_5551,N_4641,N_4738);
nand U5552 (N_5552,N_4111,N_3889);
xnor U5553 (N_5553,N_4316,N_4305);
xor U5554 (N_5554,N_3684,N_3765);
and U5555 (N_5555,N_4117,N_4553);
xnor U5556 (N_5556,N_4752,N_4543);
nand U5557 (N_5557,N_4658,N_4696);
and U5558 (N_5558,N_4482,N_3668);
and U5559 (N_5559,N_4444,N_4748);
or U5560 (N_5560,N_3868,N_4017);
and U5561 (N_5561,N_4633,N_3967);
nand U5562 (N_5562,N_4532,N_4637);
xor U5563 (N_5563,N_4525,N_4215);
and U5564 (N_5564,N_3616,N_3704);
nand U5565 (N_5565,N_4289,N_4581);
xnor U5566 (N_5566,N_3767,N_4294);
nand U5567 (N_5567,N_3966,N_3732);
nand U5568 (N_5568,N_4242,N_4160);
xor U5569 (N_5569,N_3965,N_4589);
or U5570 (N_5570,N_4443,N_4656);
xor U5571 (N_5571,N_4176,N_4788);
nor U5572 (N_5572,N_3656,N_4750);
nor U5573 (N_5573,N_4644,N_3726);
nor U5574 (N_5574,N_3930,N_4697);
nand U5575 (N_5575,N_4229,N_4010);
and U5576 (N_5576,N_4534,N_4174);
nand U5577 (N_5577,N_3785,N_4454);
nand U5578 (N_5578,N_3866,N_4001);
nand U5579 (N_5579,N_3845,N_4629);
nor U5580 (N_5580,N_4156,N_3641);
nor U5581 (N_5581,N_4352,N_4798);
nand U5582 (N_5582,N_3611,N_4786);
nor U5583 (N_5583,N_4106,N_4487);
xor U5584 (N_5584,N_3813,N_4728);
or U5585 (N_5585,N_4167,N_4041);
or U5586 (N_5586,N_4605,N_4707);
xor U5587 (N_5587,N_3639,N_3696);
nor U5588 (N_5588,N_4621,N_4600);
and U5589 (N_5589,N_3954,N_4002);
and U5590 (N_5590,N_4783,N_3887);
and U5591 (N_5591,N_3817,N_4195);
or U5592 (N_5592,N_4369,N_4456);
and U5593 (N_5593,N_4014,N_4077);
nor U5594 (N_5594,N_4314,N_3715);
nor U5595 (N_5595,N_4677,N_4227);
xor U5596 (N_5596,N_4394,N_4287);
and U5597 (N_5597,N_3696,N_3969);
nor U5598 (N_5598,N_4323,N_3825);
and U5599 (N_5599,N_4383,N_4290);
or U5600 (N_5600,N_3975,N_4172);
nand U5601 (N_5601,N_4215,N_4533);
nand U5602 (N_5602,N_3603,N_4172);
nand U5603 (N_5603,N_4012,N_3823);
nor U5604 (N_5604,N_4021,N_4671);
nand U5605 (N_5605,N_4670,N_4329);
or U5606 (N_5606,N_3656,N_4250);
xnor U5607 (N_5607,N_3790,N_4289);
nand U5608 (N_5608,N_3720,N_3626);
or U5609 (N_5609,N_4607,N_4041);
xor U5610 (N_5610,N_4711,N_3704);
xnor U5611 (N_5611,N_4659,N_4280);
xor U5612 (N_5612,N_3930,N_4274);
or U5613 (N_5613,N_4314,N_4339);
and U5614 (N_5614,N_4435,N_4459);
or U5615 (N_5615,N_3794,N_4393);
and U5616 (N_5616,N_3920,N_4440);
or U5617 (N_5617,N_4368,N_3790);
nand U5618 (N_5618,N_4290,N_4542);
nor U5619 (N_5619,N_3926,N_4128);
nand U5620 (N_5620,N_4751,N_4618);
and U5621 (N_5621,N_4275,N_4454);
nand U5622 (N_5622,N_3839,N_3638);
xnor U5623 (N_5623,N_4681,N_3977);
or U5624 (N_5624,N_4470,N_3834);
xnor U5625 (N_5625,N_4504,N_4672);
nand U5626 (N_5626,N_4091,N_4057);
nand U5627 (N_5627,N_4478,N_3812);
or U5628 (N_5628,N_4311,N_4488);
nor U5629 (N_5629,N_4221,N_4637);
and U5630 (N_5630,N_4436,N_4657);
and U5631 (N_5631,N_3792,N_3807);
xor U5632 (N_5632,N_4670,N_4733);
nand U5633 (N_5633,N_3771,N_4479);
nor U5634 (N_5634,N_4332,N_3790);
or U5635 (N_5635,N_4100,N_4547);
nand U5636 (N_5636,N_4728,N_3698);
nor U5637 (N_5637,N_4092,N_4517);
and U5638 (N_5638,N_3824,N_3951);
nor U5639 (N_5639,N_4498,N_4256);
xnor U5640 (N_5640,N_4033,N_4782);
and U5641 (N_5641,N_3880,N_4423);
nand U5642 (N_5642,N_4764,N_4588);
or U5643 (N_5643,N_3707,N_3880);
and U5644 (N_5644,N_4002,N_4510);
and U5645 (N_5645,N_4643,N_3867);
nor U5646 (N_5646,N_3826,N_4500);
xnor U5647 (N_5647,N_4207,N_4557);
nor U5648 (N_5648,N_3900,N_4597);
or U5649 (N_5649,N_3694,N_3788);
or U5650 (N_5650,N_4464,N_4073);
and U5651 (N_5651,N_3994,N_4238);
and U5652 (N_5652,N_4150,N_4293);
nand U5653 (N_5653,N_4196,N_4796);
or U5654 (N_5654,N_4286,N_3808);
nor U5655 (N_5655,N_3946,N_4433);
or U5656 (N_5656,N_4402,N_4787);
nor U5657 (N_5657,N_4694,N_4626);
and U5658 (N_5658,N_3617,N_4116);
and U5659 (N_5659,N_4212,N_4049);
or U5660 (N_5660,N_3737,N_3702);
nor U5661 (N_5661,N_4748,N_4195);
xnor U5662 (N_5662,N_4529,N_3852);
nand U5663 (N_5663,N_4038,N_4270);
xnor U5664 (N_5664,N_4533,N_4096);
or U5665 (N_5665,N_3695,N_3656);
nand U5666 (N_5666,N_4609,N_4708);
xnor U5667 (N_5667,N_4687,N_4733);
nand U5668 (N_5668,N_4161,N_4756);
and U5669 (N_5669,N_4591,N_4264);
nor U5670 (N_5670,N_3697,N_4241);
xnor U5671 (N_5671,N_4775,N_4079);
nor U5672 (N_5672,N_4388,N_4404);
nor U5673 (N_5673,N_4036,N_3861);
xor U5674 (N_5674,N_3882,N_4490);
nand U5675 (N_5675,N_4320,N_4127);
nor U5676 (N_5676,N_4200,N_4623);
nor U5677 (N_5677,N_4056,N_4047);
or U5678 (N_5678,N_3702,N_4260);
nor U5679 (N_5679,N_4422,N_4079);
and U5680 (N_5680,N_4455,N_3881);
and U5681 (N_5681,N_3990,N_4699);
nor U5682 (N_5682,N_4656,N_3737);
nor U5683 (N_5683,N_4314,N_4186);
nor U5684 (N_5684,N_4536,N_4466);
nand U5685 (N_5685,N_4402,N_4175);
or U5686 (N_5686,N_4011,N_4035);
nand U5687 (N_5687,N_3887,N_4266);
xor U5688 (N_5688,N_4102,N_4295);
nand U5689 (N_5689,N_4701,N_3617);
nand U5690 (N_5690,N_3700,N_4576);
xor U5691 (N_5691,N_3925,N_4705);
and U5692 (N_5692,N_4482,N_4780);
nand U5693 (N_5693,N_4342,N_4619);
xor U5694 (N_5694,N_4477,N_3934);
and U5695 (N_5695,N_4021,N_4430);
nor U5696 (N_5696,N_4142,N_3914);
nand U5697 (N_5697,N_3964,N_4005);
and U5698 (N_5698,N_4258,N_4538);
or U5699 (N_5699,N_3847,N_3784);
nand U5700 (N_5700,N_3923,N_3963);
or U5701 (N_5701,N_4477,N_4503);
nand U5702 (N_5702,N_3610,N_4546);
xnor U5703 (N_5703,N_4756,N_3915);
xor U5704 (N_5704,N_3662,N_4028);
xnor U5705 (N_5705,N_4713,N_3983);
and U5706 (N_5706,N_4361,N_4547);
nand U5707 (N_5707,N_3860,N_4378);
or U5708 (N_5708,N_4754,N_3695);
and U5709 (N_5709,N_4489,N_4753);
nand U5710 (N_5710,N_3789,N_4493);
and U5711 (N_5711,N_4729,N_4570);
and U5712 (N_5712,N_4134,N_4160);
nand U5713 (N_5713,N_4381,N_4211);
nand U5714 (N_5714,N_4200,N_3875);
xnor U5715 (N_5715,N_3913,N_4253);
or U5716 (N_5716,N_4649,N_4655);
nor U5717 (N_5717,N_4089,N_4291);
nor U5718 (N_5718,N_3799,N_4304);
xnor U5719 (N_5719,N_4223,N_4550);
and U5720 (N_5720,N_4420,N_3995);
and U5721 (N_5721,N_4752,N_3650);
and U5722 (N_5722,N_3800,N_4562);
xnor U5723 (N_5723,N_3866,N_4268);
nand U5724 (N_5724,N_3658,N_4267);
nor U5725 (N_5725,N_4202,N_4026);
xor U5726 (N_5726,N_3792,N_3906);
nand U5727 (N_5727,N_4154,N_4689);
or U5728 (N_5728,N_3606,N_3962);
nand U5729 (N_5729,N_4426,N_4384);
nor U5730 (N_5730,N_3889,N_3656);
and U5731 (N_5731,N_4777,N_4646);
nor U5732 (N_5732,N_3825,N_4160);
xnor U5733 (N_5733,N_4408,N_3751);
and U5734 (N_5734,N_3944,N_4294);
xnor U5735 (N_5735,N_4478,N_3925);
or U5736 (N_5736,N_4526,N_4681);
nor U5737 (N_5737,N_4681,N_4192);
or U5738 (N_5738,N_4697,N_3954);
nand U5739 (N_5739,N_3780,N_3887);
and U5740 (N_5740,N_4576,N_4480);
or U5741 (N_5741,N_3606,N_4664);
xor U5742 (N_5742,N_4234,N_3908);
xnor U5743 (N_5743,N_3974,N_4726);
and U5744 (N_5744,N_4171,N_4593);
xnor U5745 (N_5745,N_4168,N_4340);
xor U5746 (N_5746,N_3930,N_3627);
xnor U5747 (N_5747,N_3691,N_4267);
xor U5748 (N_5748,N_3778,N_4643);
nand U5749 (N_5749,N_3862,N_3991);
or U5750 (N_5750,N_4742,N_4136);
nor U5751 (N_5751,N_4030,N_3939);
nand U5752 (N_5752,N_4237,N_4161);
or U5753 (N_5753,N_4332,N_4518);
xnor U5754 (N_5754,N_4208,N_4593);
nor U5755 (N_5755,N_3882,N_4608);
nor U5756 (N_5756,N_3970,N_4787);
xor U5757 (N_5757,N_4608,N_4713);
nor U5758 (N_5758,N_4070,N_3659);
nand U5759 (N_5759,N_3776,N_3625);
or U5760 (N_5760,N_3930,N_4260);
or U5761 (N_5761,N_4007,N_3717);
nor U5762 (N_5762,N_4622,N_4624);
xor U5763 (N_5763,N_3616,N_4078);
and U5764 (N_5764,N_4173,N_4590);
or U5765 (N_5765,N_4451,N_3924);
nor U5766 (N_5766,N_4349,N_3809);
or U5767 (N_5767,N_3960,N_4070);
nor U5768 (N_5768,N_3693,N_4298);
nor U5769 (N_5769,N_3889,N_3837);
and U5770 (N_5770,N_4240,N_4344);
or U5771 (N_5771,N_4091,N_4197);
xor U5772 (N_5772,N_3662,N_4279);
xnor U5773 (N_5773,N_4450,N_4484);
nand U5774 (N_5774,N_4209,N_3759);
nand U5775 (N_5775,N_3740,N_4409);
xor U5776 (N_5776,N_4155,N_4308);
and U5777 (N_5777,N_3770,N_4153);
or U5778 (N_5778,N_4008,N_4198);
nand U5779 (N_5779,N_3989,N_4360);
and U5780 (N_5780,N_3681,N_4457);
xor U5781 (N_5781,N_4273,N_4380);
xnor U5782 (N_5782,N_3838,N_4272);
xor U5783 (N_5783,N_4364,N_3658);
xnor U5784 (N_5784,N_4117,N_4681);
or U5785 (N_5785,N_4305,N_3635);
nor U5786 (N_5786,N_4507,N_4222);
or U5787 (N_5787,N_4014,N_4651);
nor U5788 (N_5788,N_3600,N_4391);
nand U5789 (N_5789,N_4736,N_4467);
and U5790 (N_5790,N_4037,N_3687);
nor U5791 (N_5791,N_4235,N_4064);
and U5792 (N_5792,N_3667,N_4362);
and U5793 (N_5793,N_4607,N_4515);
xor U5794 (N_5794,N_4443,N_4618);
and U5795 (N_5795,N_3928,N_3728);
nand U5796 (N_5796,N_4223,N_4447);
xor U5797 (N_5797,N_4263,N_3760);
nor U5798 (N_5798,N_4346,N_4201);
or U5799 (N_5799,N_4382,N_4302);
xnor U5800 (N_5800,N_3992,N_4688);
nor U5801 (N_5801,N_3747,N_3933);
xnor U5802 (N_5802,N_4615,N_4674);
xor U5803 (N_5803,N_3624,N_4398);
or U5804 (N_5804,N_3932,N_4078);
and U5805 (N_5805,N_4265,N_4422);
xor U5806 (N_5806,N_3948,N_4296);
and U5807 (N_5807,N_3807,N_4136);
nor U5808 (N_5808,N_4294,N_4426);
and U5809 (N_5809,N_4204,N_3950);
and U5810 (N_5810,N_4079,N_4729);
or U5811 (N_5811,N_4188,N_4135);
or U5812 (N_5812,N_4565,N_4048);
and U5813 (N_5813,N_3653,N_3915);
and U5814 (N_5814,N_3801,N_4758);
and U5815 (N_5815,N_4484,N_4364);
nor U5816 (N_5816,N_4772,N_4220);
xor U5817 (N_5817,N_4234,N_3659);
and U5818 (N_5818,N_3832,N_4366);
and U5819 (N_5819,N_4006,N_3728);
or U5820 (N_5820,N_3996,N_3879);
and U5821 (N_5821,N_4733,N_4296);
nor U5822 (N_5822,N_4198,N_4490);
xnor U5823 (N_5823,N_3852,N_4282);
or U5824 (N_5824,N_3971,N_4069);
nand U5825 (N_5825,N_4632,N_4539);
nand U5826 (N_5826,N_3634,N_4318);
xor U5827 (N_5827,N_3934,N_4455);
and U5828 (N_5828,N_4311,N_4261);
or U5829 (N_5829,N_4077,N_4183);
nand U5830 (N_5830,N_4305,N_3939);
nand U5831 (N_5831,N_4695,N_3906);
nor U5832 (N_5832,N_3665,N_4174);
and U5833 (N_5833,N_3643,N_4168);
nand U5834 (N_5834,N_4017,N_3759);
nor U5835 (N_5835,N_4223,N_4429);
and U5836 (N_5836,N_4519,N_3796);
and U5837 (N_5837,N_4363,N_4344);
xor U5838 (N_5838,N_4098,N_3828);
and U5839 (N_5839,N_4131,N_4032);
xor U5840 (N_5840,N_4723,N_4624);
xor U5841 (N_5841,N_4529,N_4733);
xnor U5842 (N_5842,N_3931,N_4391);
nand U5843 (N_5843,N_4259,N_4729);
nor U5844 (N_5844,N_3632,N_4171);
xnor U5845 (N_5845,N_3637,N_3609);
nor U5846 (N_5846,N_3698,N_4308);
xor U5847 (N_5847,N_4778,N_4414);
nor U5848 (N_5848,N_4135,N_4581);
xor U5849 (N_5849,N_3768,N_4512);
or U5850 (N_5850,N_3892,N_3721);
nor U5851 (N_5851,N_3741,N_4355);
nand U5852 (N_5852,N_3768,N_3727);
xor U5853 (N_5853,N_4424,N_4331);
nand U5854 (N_5854,N_3950,N_4730);
and U5855 (N_5855,N_3982,N_3720);
xnor U5856 (N_5856,N_4388,N_3674);
nand U5857 (N_5857,N_4029,N_3791);
xnor U5858 (N_5858,N_4131,N_3971);
or U5859 (N_5859,N_3963,N_4719);
nand U5860 (N_5860,N_4789,N_4267);
and U5861 (N_5861,N_3800,N_4576);
nand U5862 (N_5862,N_3934,N_3987);
xnor U5863 (N_5863,N_3692,N_4411);
xnor U5864 (N_5864,N_4268,N_4233);
nand U5865 (N_5865,N_4404,N_3661);
nor U5866 (N_5866,N_3864,N_4726);
and U5867 (N_5867,N_4118,N_4063);
xor U5868 (N_5868,N_4615,N_4758);
or U5869 (N_5869,N_3807,N_4000);
nand U5870 (N_5870,N_4319,N_4448);
or U5871 (N_5871,N_4207,N_4267);
nand U5872 (N_5872,N_4266,N_4179);
nand U5873 (N_5873,N_4440,N_4267);
or U5874 (N_5874,N_4595,N_3797);
nand U5875 (N_5875,N_4476,N_4364);
nand U5876 (N_5876,N_4658,N_4555);
xor U5877 (N_5877,N_4128,N_3885);
xor U5878 (N_5878,N_3708,N_3785);
nand U5879 (N_5879,N_4375,N_3823);
nor U5880 (N_5880,N_3729,N_4011);
nand U5881 (N_5881,N_4095,N_4388);
and U5882 (N_5882,N_3926,N_4244);
nand U5883 (N_5883,N_4488,N_4475);
nor U5884 (N_5884,N_4176,N_4718);
or U5885 (N_5885,N_3965,N_4415);
and U5886 (N_5886,N_4723,N_3703);
nand U5887 (N_5887,N_4529,N_4364);
and U5888 (N_5888,N_4339,N_4487);
nor U5889 (N_5889,N_3684,N_4791);
or U5890 (N_5890,N_4753,N_3624);
and U5891 (N_5891,N_3773,N_3715);
xnor U5892 (N_5892,N_4533,N_3827);
and U5893 (N_5893,N_4557,N_4086);
nor U5894 (N_5894,N_3825,N_3886);
and U5895 (N_5895,N_3878,N_3844);
xnor U5896 (N_5896,N_3644,N_4035);
xor U5897 (N_5897,N_4439,N_4098);
xnor U5898 (N_5898,N_3761,N_3640);
and U5899 (N_5899,N_4206,N_3956);
and U5900 (N_5900,N_3684,N_3868);
or U5901 (N_5901,N_4505,N_4577);
or U5902 (N_5902,N_3780,N_4364);
nand U5903 (N_5903,N_4480,N_4699);
or U5904 (N_5904,N_3981,N_4445);
xnor U5905 (N_5905,N_3630,N_4529);
or U5906 (N_5906,N_4053,N_3842);
or U5907 (N_5907,N_4641,N_4701);
nand U5908 (N_5908,N_3987,N_3806);
and U5909 (N_5909,N_3621,N_4530);
and U5910 (N_5910,N_3617,N_4550);
or U5911 (N_5911,N_4575,N_3920);
xor U5912 (N_5912,N_4143,N_4488);
and U5913 (N_5913,N_4233,N_4606);
nor U5914 (N_5914,N_4648,N_4405);
xnor U5915 (N_5915,N_3638,N_4446);
or U5916 (N_5916,N_4365,N_3728);
nand U5917 (N_5917,N_4527,N_3709);
or U5918 (N_5918,N_3888,N_4681);
nand U5919 (N_5919,N_4708,N_3732);
xor U5920 (N_5920,N_4158,N_3737);
nor U5921 (N_5921,N_4290,N_4698);
nand U5922 (N_5922,N_4714,N_4599);
nand U5923 (N_5923,N_4600,N_4757);
nor U5924 (N_5924,N_4077,N_4781);
xor U5925 (N_5925,N_4228,N_4077);
xor U5926 (N_5926,N_3880,N_3750);
nand U5927 (N_5927,N_4677,N_4083);
or U5928 (N_5928,N_4043,N_3957);
nor U5929 (N_5929,N_3687,N_4282);
xnor U5930 (N_5930,N_3601,N_3703);
nand U5931 (N_5931,N_3766,N_3908);
nand U5932 (N_5932,N_3806,N_3743);
nand U5933 (N_5933,N_4597,N_4602);
and U5934 (N_5934,N_4331,N_4535);
xnor U5935 (N_5935,N_3738,N_4263);
nor U5936 (N_5936,N_4526,N_4210);
or U5937 (N_5937,N_3932,N_3967);
xnor U5938 (N_5938,N_3698,N_4445);
and U5939 (N_5939,N_3838,N_4748);
nor U5940 (N_5940,N_4652,N_4177);
nand U5941 (N_5941,N_3889,N_4787);
nand U5942 (N_5942,N_4349,N_4668);
xnor U5943 (N_5943,N_4101,N_4280);
nand U5944 (N_5944,N_4317,N_3686);
or U5945 (N_5945,N_3952,N_4162);
and U5946 (N_5946,N_3612,N_4036);
nor U5947 (N_5947,N_4319,N_3885);
or U5948 (N_5948,N_4368,N_4732);
xnor U5949 (N_5949,N_3967,N_4456);
nor U5950 (N_5950,N_4171,N_4361);
xor U5951 (N_5951,N_4395,N_4242);
and U5952 (N_5952,N_4294,N_3615);
nand U5953 (N_5953,N_3924,N_3946);
or U5954 (N_5954,N_4192,N_4430);
nor U5955 (N_5955,N_4138,N_3980);
or U5956 (N_5956,N_4434,N_4744);
nand U5957 (N_5957,N_4544,N_4263);
xor U5958 (N_5958,N_4341,N_4140);
or U5959 (N_5959,N_4505,N_3752);
nor U5960 (N_5960,N_4656,N_4149);
nand U5961 (N_5961,N_3924,N_4218);
nor U5962 (N_5962,N_4156,N_4157);
xor U5963 (N_5963,N_3651,N_3870);
nand U5964 (N_5964,N_4750,N_4314);
xnor U5965 (N_5965,N_4667,N_4060);
and U5966 (N_5966,N_3657,N_4047);
nor U5967 (N_5967,N_4494,N_4054);
nor U5968 (N_5968,N_4612,N_4537);
nand U5969 (N_5969,N_4033,N_4779);
nand U5970 (N_5970,N_4537,N_4395);
nand U5971 (N_5971,N_4183,N_3678);
and U5972 (N_5972,N_4129,N_4605);
or U5973 (N_5973,N_4709,N_4705);
nand U5974 (N_5974,N_4000,N_3833);
or U5975 (N_5975,N_4097,N_3902);
or U5976 (N_5976,N_4716,N_4627);
nand U5977 (N_5977,N_3937,N_4744);
nand U5978 (N_5978,N_4080,N_3952);
nand U5979 (N_5979,N_3642,N_4133);
nand U5980 (N_5980,N_4735,N_4059);
nand U5981 (N_5981,N_3857,N_4072);
xor U5982 (N_5982,N_3876,N_3660);
and U5983 (N_5983,N_3934,N_4395);
nor U5984 (N_5984,N_3621,N_3730);
or U5985 (N_5985,N_3731,N_3840);
nand U5986 (N_5986,N_4045,N_4224);
nor U5987 (N_5987,N_4034,N_3694);
nand U5988 (N_5988,N_4201,N_3810);
or U5989 (N_5989,N_4220,N_3852);
nand U5990 (N_5990,N_4431,N_4256);
nor U5991 (N_5991,N_3778,N_4422);
xor U5992 (N_5992,N_4220,N_4488);
nor U5993 (N_5993,N_4476,N_4723);
and U5994 (N_5994,N_4699,N_3768);
nand U5995 (N_5995,N_3851,N_4159);
nor U5996 (N_5996,N_4001,N_4482);
nor U5997 (N_5997,N_4380,N_3689);
and U5998 (N_5998,N_4296,N_3803);
nor U5999 (N_5999,N_4700,N_4696);
nand U6000 (N_6000,N_5313,N_5103);
or U6001 (N_6001,N_4914,N_5218);
xor U6002 (N_6002,N_4955,N_4923);
xnor U6003 (N_6003,N_5944,N_5807);
xnor U6004 (N_6004,N_5511,N_5893);
and U6005 (N_6005,N_5651,N_5362);
nor U6006 (N_6006,N_4962,N_4998);
nor U6007 (N_6007,N_5181,N_5478);
xnor U6008 (N_6008,N_5413,N_4970);
nand U6009 (N_6009,N_5395,N_5404);
or U6010 (N_6010,N_5906,N_4941);
xnor U6011 (N_6011,N_5668,N_4950);
and U6012 (N_6012,N_5577,N_5914);
or U6013 (N_6013,N_5846,N_5912);
or U6014 (N_6014,N_5001,N_5843);
and U6015 (N_6015,N_5146,N_4869);
nand U6016 (N_6016,N_5054,N_5081);
or U6017 (N_6017,N_5245,N_5141);
and U6018 (N_6018,N_5255,N_5350);
and U6019 (N_6019,N_5080,N_5215);
nor U6020 (N_6020,N_5832,N_4885);
nand U6021 (N_6021,N_5004,N_5866);
nor U6022 (N_6022,N_4992,N_5749);
xor U6023 (N_6023,N_4937,N_5370);
nand U6024 (N_6024,N_5780,N_5116);
nor U6025 (N_6025,N_5879,N_5382);
and U6026 (N_6026,N_5674,N_5186);
and U6027 (N_6027,N_5620,N_5208);
nand U6028 (N_6028,N_5176,N_5910);
nor U6029 (N_6029,N_5718,N_5018);
xnor U6030 (N_6030,N_5751,N_5451);
xnor U6031 (N_6031,N_5529,N_5528);
nand U6032 (N_6032,N_4908,N_5641);
and U6033 (N_6033,N_5523,N_5840);
nor U6034 (N_6034,N_5226,N_5729);
and U6035 (N_6035,N_5934,N_4911);
nand U6036 (N_6036,N_5995,N_5360);
and U6037 (N_6037,N_4919,N_5073);
nand U6038 (N_6038,N_5688,N_4929);
xor U6039 (N_6039,N_5170,N_4975);
nor U6040 (N_6040,N_5785,N_4991);
nor U6041 (N_6041,N_4823,N_5712);
nor U6042 (N_6042,N_5924,N_5050);
xnor U6043 (N_6043,N_5761,N_5673);
xor U6044 (N_6044,N_5069,N_5857);
nor U6045 (N_6045,N_5051,N_5822);
nor U6046 (N_6046,N_5532,N_5762);
nor U6047 (N_6047,N_5006,N_5939);
nand U6048 (N_6048,N_4898,N_4857);
and U6049 (N_6049,N_5294,N_5514);
xnor U6050 (N_6050,N_5520,N_5166);
xnor U6051 (N_6051,N_5450,N_5991);
and U6052 (N_6052,N_5479,N_5827);
nand U6053 (N_6053,N_5396,N_5072);
xnor U6054 (N_6054,N_5689,N_5552);
xnor U6055 (N_6055,N_5950,N_5896);
xor U6056 (N_6056,N_4932,N_5344);
and U6057 (N_6057,N_5766,N_5682);
xor U6058 (N_6058,N_5587,N_5562);
nor U6059 (N_6059,N_5709,N_5206);
and U6060 (N_6060,N_5379,N_5639);
xnor U6061 (N_6061,N_5687,N_5329);
nand U6062 (N_6062,N_5195,N_5736);
and U6063 (N_6063,N_5610,N_5560);
nand U6064 (N_6064,N_5868,N_5873);
xnor U6065 (N_6065,N_5284,N_4895);
or U6066 (N_6066,N_5459,N_5767);
and U6067 (N_6067,N_5618,N_5568);
nor U6068 (N_6068,N_5371,N_5745);
nor U6069 (N_6069,N_4994,N_4920);
nand U6070 (N_6070,N_4814,N_5183);
and U6071 (N_6071,N_5772,N_5209);
xor U6072 (N_6072,N_5306,N_5207);
xor U6073 (N_6073,N_5515,N_5854);
or U6074 (N_6074,N_5096,N_5229);
or U6075 (N_6075,N_5897,N_5653);
xor U6076 (N_6076,N_5647,N_5829);
or U6077 (N_6077,N_5128,N_5900);
xnor U6078 (N_6078,N_5833,N_4935);
and U6079 (N_6079,N_5999,N_5569);
and U6080 (N_6080,N_5929,N_4806);
nor U6081 (N_6081,N_5996,N_5440);
or U6082 (N_6082,N_5022,N_5037);
and U6083 (N_6083,N_5596,N_5706);
xnor U6084 (N_6084,N_5364,N_4847);
nor U6085 (N_6085,N_5608,N_5928);
nor U6086 (N_6086,N_5118,N_4948);
xor U6087 (N_6087,N_5115,N_5705);
nor U6088 (N_6088,N_5352,N_5921);
nor U6089 (N_6089,N_5679,N_5984);
and U6090 (N_6090,N_5010,N_5519);
and U6091 (N_6091,N_5769,N_5269);
nor U6092 (N_6092,N_4901,N_4800);
xnor U6093 (N_6093,N_5325,N_5919);
and U6094 (N_6094,N_5889,N_4853);
xnor U6095 (N_6095,N_4931,N_5390);
nor U6096 (N_6096,N_5951,N_5424);
nand U6097 (N_6097,N_5825,N_5504);
nor U6098 (N_6098,N_5828,N_5804);
nor U6099 (N_6099,N_5499,N_5722);
nand U6100 (N_6100,N_4968,N_4933);
xor U6101 (N_6101,N_5714,N_5506);
nand U6102 (N_6102,N_4995,N_5292);
or U6103 (N_6103,N_5266,N_5261);
nor U6104 (N_6104,N_5161,N_5711);
or U6105 (N_6105,N_5916,N_5606);
nor U6106 (N_6106,N_5727,N_5017);
or U6107 (N_6107,N_5310,N_5332);
or U6108 (N_6108,N_4876,N_4945);
or U6109 (N_6109,N_5730,N_5578);
and U6110 (N_6110,N_4934,N_5252);
or U6111 (N_6111,N_5631,N_5307);
or U6112 (N_6112,N_5923,N_5881);
and U6113 (N_6113,N_4839,N_5592);
nor U6114 (N_6114,N_5095,N_4969);
or U6115 (N_6115,N_4871,N_5091);
nor U6116 (N_6116,N_5263,N_5258);
and U6117 (N_6117,N_5342,N_4827);
and U6118 (N_6118,N_5670,N_5898);
nor U6119 (N_6119,N_4826,N_5955);
xor U6120 (N_6120,N_5223,N_5156);
nor U6121 (N_6121,N_4805,N_5940);
nor U6122 (N_6122,N_5537,N_5216);
or U6123 (N_6123,N_5801,N_4884);
or U6124 (N_6124,N_5628,N_5401);
nor U6125 (N_6125,N_4974,N_5811);
nor U6126 (N_6126,N_5861,N_5957);
or U6127 (N_6127,N_5633,N_4952);
and U6128 (N_6128,N_5570,N_5427);
nand U6129 (N_6129,N_5715,N_5199);
xnor U6130 (N_6130,N_5544,N_5841);
nand U6131 (N_6131,N_5244,N_5271);
and U6132 (N_6132,N_5009,N_5160);
and U6133 (N_6133,N_5474,N_5844);
xnor U6134 (N_6134,N_5201,N_5100);
nor U6135 (N_6135,N_5075,N_5556);
nand U6136 (N_6136,N_5510,N_5876);
nor U6137 (N_6137,N_5421,N_5959);
and U6138 (N_6138,N_5667,N_4821);
nor U6139 (N_6139,N_5129,N_5656);
nor U6140 (N_6140,N_5036,N_5473);
nor U6141 (N_6141,N_4822,N_5131);
nand U6142 (N_6142,N_5227,N_5301);
xnor U6143 (N_6143,N_5475,N_5085);
or U6144 (N_6144,N_5287,N_4907);
xnor U6145 (N_6145,N_5782,N_5402);
and U6146 (N_6146,N_5487,N_5591);
nand U6147 (N_6147,N_5792,N_5649);
nor U6148 (N_6148,N_5589,N_5175);
and U6149 (N_6149,N_5423,N_5806);
xor U6150 (N_6150,N_5717,N_5016);
and U6151 (N_6151,N_5977,N_4852);
xnor U6152 (N_6152,N_5617,N_5583);
xor U6153 (N_6153,N_5970,N_5978);
nand U6154 (N_6154,N_5071,N_5340);
or U6155 (N_6155,N_5627,N_4987);
nor U6156 (N_6156,N_5481,N_5905);
xnor U6157 (N_6157,N_5975,N_5174);
and U6158 (N_6158,N_5490,N_5874);
and U6159 (N_6159,N_5455,N_5860);
xnor U6160 (N_6160,N_5575,N_5613);
nor U6161 (N_6161,N_5400,N_5927);
nand U6162 (N_6162,N_5406,N_5045);
nor U6163 (N_6163,N_4926,N_5911);
nor U6164 (N_6164,N_5441,N_5983);
nor U6165 (N_6165,N_4858,N_5847);
xnor U6166 (N_6166,N_4928,N_5965);
xor U6167 (N_6167,N_5783,N_5661);
xnor U6168 (N_6168,N_5738,N_5856);
nor U6169 (N_6169,N_5025,N_5770);
nand U6170 (N_6170,N_5431,N_5005);
and U6171 (N_6171,N_5590,N_4954);
xnor U6172 (N_6172,N_4918,N_4832);
and U6173 (N_6173,N_5665,N_5937);
and U6174 (N_6174,N_5979,N_5925);
or U6175 (N_6175,N_5225,N_4836);
nand U6176 (N_6176,N_5849,N_5077);
nand U6177 (N_6177,N_5164,N_5626);
nor U6178 (N_6178,N_5147,N_4875);
nand U6179 (N_6179,N_5445,N_5657);
or U6180 (N_6180,N_5264,N_5611);
xor U6181 (N_6181,N_4803,N_5558);
nor U6182 (N_6182,N_5602,N_4840);
nand U6183 (N_6183,N_5132,N_5039);
xnor U6184 (N_6184,N_5391,N_5331);
nor U6185 (N_6185,N_5823,N_5040);
nand U6186 (N_6186,N_5437,N_5594);
xor U6187 (N_6187,N_5411,N_5138);
and U6188 (N_6188,N_5795,N_5581);
and U6189 (N_6189,N_5660,N_5148);
and U6190 (N_6190,N_5887,N_5516);
and U6191 (N_6191,N_5343,N_5677);
or U6192 (N_6192,N_5457,N_5047);
nand U6193 (N_6193,N_4925,N_5130);
nand U6194 (N_6194,N_5810,N_4837);
and U6195 (N_6195,N_5716,N_5632);
or U6196 (N_6196,N_5824,N_5752);
nor U6197 (N_6197,N_5742,N_5086);
and U6198 (N_6198,N_5399,N_5277);
nand U6199 (N_6199,N_4889,N_5774);
nor U6200 (N_6200,N_5328,N_5855);
nor U6201 (N_6201,N_5393,N_5470);
nor U6202 (N_6202,N_5802,N_5623);
xnor U6203 (N_6203,N_5852,N_5820);
nand U6204 (N_6204,N_5374,N_5540);
nand U6205 (N_6205,N_5865,N_5961);
and U6206 (N_6206,N_5122,N_4942);
or U6207 (N_6207,N_4881,N_5188);
and U6208 (N_6208,N_4855,N_5296);
nand U6209 (N_6209,N_5065,N_5638);
xnor U6210 (N_6210,N_5491,N_5737);
and U6211 (N_6211,N_5488,N_5375);
nand U6212 (N_6212,N_5253,N_5121);
or U6213 (N_6213,N_5388,N_5410);
xnor U6214 (N_6214,N_5755,N_5178);
or U6215 (N_6215,N_4978,N_5456);
xnor U6216 (N_6216,N_5068,N_5376);
nand U6217 (N_6217,N_5538,N_5011);
xor U6218 (N_6218,N_4862,N_5601);
xor U6219 (N_6219,N_5859,N_5463);
xnor U6220 (N_6220,N_5707,N_5561);
and U6221 (N_6221,N_5259,N_5798);
nor U6222 (N_6222,N_5312,N_5214);
nor U6223 (N_6223,N_4873,N_5980);
or U6224 (N_6224,N_4812,N_5526);
nor U6225 (N_6225,N_5584,N_5576);
nor U6226 (N_6226,N_4940,N_5619);
and U6227 (N_6227,N_5434,N_5527);
and U6228 (N_6228,N_5713,N_5298);
or U6229 (N_6229,N_4838,N_5694);
or U6230 (N_6230,N_5438,N_5383);
xnor U6231 (N_6231,N_5143,N_5177);
xor U6232 (N_6232,N_5685,N_4865);
xor U6233 (N_6233,N_5165,N_5875);
and U6234 (N_6234,N_5759,N_5358);
or U6235 (N_6235,N_4880,N_5436);
xor U6236 (N_6236,N_5405,N_5056);
and U6237 (N_6237,N_5797,N_5321);
or U6238 (N_6238,N_5407,N_5880);
nor U6239 (N_6239,N_4820,N_5947);
and U6240 (N_6240,N_5337,N_5369);
nand U6241 (N_6241,N_5235,N_4984);
xnor U6242 (N_6242,N_5744,N_5239);
nand U6243 (N_6243,N_5636,N_5468);
xor U6244 (N_6244,N_4807,N_5748);
xor U6245 (N_6245,N_4924,N_5192);
or U6246 (N_6246,N_5741,N_5913);
xor U6247 (N_6247,N_5327,N_5543);
or U6248 (N_6248,N_5200,N_5243);
and U6249 (N_6249,N_5120,N_4867);
nand U6250 (N_6250,N_5884,N_5734);
nor U6251 (N_6251,N_4859,N_5886);
and U6252 (N_6252,N_4927,N_5942);
nand U6253 (N_6253,N_5270,N_5816);
nand U6254 (N_6254,N_5791,N_5163);
xnor U6255 (N_6255,N_5593,N_5835);
nand U6256 (N_6256,N_4834,N_5052);
and U6257 (N_6257,N_5347,N_4996);
or U6258 (N_6258,N_5548,N_5439);
xnor U6259 (N_6259,N_4891,N_5691);
xnor U6260 (N_6260,N_5972,N_4999);
and U6261 (N_6261,N_5461,N_5267);
and U6262 (N_6262,N_5728,N_5671);
and U6263 (N_6263,N_5151,N_5184);
and U6264 (N_6264,N_5162,N_5142);
and U6265 (N_6265,N_4828,N_5700);
or U6266 (N_6266,N_5669,N_4964);
and U6267 (N_6267,N_5988,N_5559);
or U6268 (N_6268,N_5278,N_4808);
nand U6269 (N_6269,N_5140,N_5126);
xnor U6270 (N_6270,N_5197,N_5571);
nor U6271 (N_6271,N_5397,N_5877);
xor U6272 (N_6272,N_5501,N_5172);
nor U6273 (N_6273,N_4872,N_5830);
xnor U6274 (N_6274,N_5837,N_4843);
xnor U6275 (N_6275,N_5029,N_5850);
or U6276 (N_6276,N_5265,N_4982);
and U6277 (N_6277,N_5724,N_5013);
xor U6278 (N_6278,N_5318,N_5813);
nor U6279 (N_6279,N_5864,N_5609);
nand U6280 (N_6280,N_4897,N_5346);
and U6281 (N_6281,N_5469,N_5534);
nor U6282 (N_6282,N_5871,N_5027);
nand U6283 (N_6283,N_4985,N_5720);
or U6284 (N_6284,N_5974,N_5221);
xnor U6285 (N_6285,N_5895,N_4811);
or U6286 (N_6286,N_5546,N_5842);
xor U6287 (N_6287,N_5251,N_5680);
and U6288 (N_6288,N_4888,N_5471);
and U6289 (N_6289,N_5189,N_5135);
xor U6290 (N_6290,N_5675,N_5426);
xnor U6291 (N_6291,N_5786,N_5599);
and U6292 (N_6292,N_5361,N_5489);
nor U6293 (N_6293,N_5224,N_4902);
and U6294 (N_6294,N_5721,N_5775);
nor U6295 (N_6295,N_5309,N_5708);
nand U6296 (N_6296,N_4893,N_5987);
nand U6297 (N_6297,N_5595,N_4883);
or U6298 (N_6298,N_4943,N_5926);
and U6299 (N_6299,N_5454,N_5113);
and U6300 (N_6300,N_5735,N_5418);
xor U6301 (N_6301,N_4906,N_5088);
or U6302 (N_6302,N_5392,N_5918);
xnor U6303 (N_6303,N_5153,N_5028);
and U6304 (N_6304,N_5789,N_5026);
or U6305 (N_6305,N_5863,N_4956);
nor U6306 (N_6306,N_5291,N_4863);
nor U6307 (N_6307,N_5588,N_5483);
nand U6308 (N_6308,N_5422,N_4815);
nand U6309 (N_6309,N_5845,N_5363);
nand U6310 (N_6310,N_5563,N_5003);
nor U6311 (N_6311,N_5458,N_5535);
nand U6312 (N_6312,N_5366,N_5787);
or U6313 (N_6313,N_5373,N_5064);
nand U6314 (N_6314,N_5779,N_4961);
xor U6315 (N_6315,N_5629,N_5986);
xnor U6316 (N_6316,N_5645,N_5725);
xnor U6317 (N_6317,N_5272,N_5597);
or U6318 (N_6318,N_4848,N_4809);
or U6319 (N_6319,N_5958,N_5182);
nor U6320 (N_6320,N_4949,N_5948);
and U6321 (N_6321,N_5903,N_5092);
xnor U6322 (N_6322,N_5681,N_5211);
nor U6323 (N_6323,N_5099,N_5449);
nand U6324 (N_6324,N_4993,N_5247);
nor U6325 (N_6325,N_4890,N_4856);
or U6326 (N_6326,N_5477,N_5368);
nor U6327 (N_6327,N_5196,N_4841);
nor U6328 (N_6328,N_5125,N_5696);
or U6329 (N_6329,N_5853,N_4813);
or U6330 (N_6330,N_5701,N_5960);
nor U6331 (N_6331,N_5354,N_5848);
nor U6332 (N_6332,N_5063,N_5317);
and U6333 (N_6333,N_5262,N_5981);
nor U6334 (N_6334,N_5746,N_5155);
xnor U6335 (N_6335,N_5268,N_5333);
or U6336 (N_6336,N_5624,N_5339);
nand U6337 (N_6337,N_5758,N_5892);
or U6338 (N_6338,N_5697,N_5585);
nand U6339 (N_6339,N_5019,N_5600);
nor U6340 (N_6340,N_5952,N_4971);
or U6341 (N_6341,N_4909,N_5992);
xnor U6342 (N_6342,N_5964,N_5324);
or U6343 (N_6343,N_4874,N_4844);
or U6344 (N_6344,N_5316,N_5008);
xor U6345 (N_6345,N_5812,N_4916);
or U6346 (N_6346,N_5232,N_4951);
and U6347 (N_6347,N_5607,N_5743);
xnor U6348 (N_6348,N_5090,N_5079);
nor U6349 (N_6349,N_4912,N_5238);
xnor U6350 (N_6350,N_5330,N_5582);
nor U6351 (N_6351,N_4966,N_5799);
nor U6352 (N_6352,N_5756,N_5664);
xnor U6353 (N_6353,N_5231,N_5462);
or U6354 (N_6354,N_5943,N_5930);
xnor U6355 (N_6355,N_5447,N_5137);
or U6356 (N_6356,N_4989,N_5521);
nor U6357 (N_6357,N_5945,N_5435);
nand U6358 (N_6358,N_4900,N_5522);
or U6359 (N_6359,N_5280,N_5067);
or U6360 (N_6360,N_5518,N_5496);
and U6361 (N_6361,N_4802,N_4905);
and U6362 (N_6362,N_5356,N_5551);
nor U6363 (N_6363,N_5323,N_5351);
and U6364 (N_6364,N_5684,N_4922);
xnor U6365 (N_6365,N_4981,N_5603);
nand U6366 (N_6366,N_5464,N_5282);
xnor U6367 (N_6367,N_5127,N_5249);
xnor U6368 (N_6368,N_5283,N_5048);
nand U6369 (N_6369,N_5985,N_4980);
xor U6370 (N_6370,N_5250,N_5304);
and U6371 (N_6371,N_5650,N_5159);
and U6372 (N_6372,N_5179,N_5500);
nor U6373 (N_6373,N_5831,N_4959);
or U6374 (N_6374,N_5123,N_5541);
nand U6375 (N_6375,N_5030,N_5966);
nand U6376 (N_6376,N_5355,N_5190);
nand U6377 (N_6377,N_5902,N_4846);
or U6378 (N_6378,N_5042,N_4864);
or U6379 (N_6379,N_5429,N_5394);
and U6380 (N_6380,N_5335,N_5869);
and U6381 (N_6381,N_5035,N_4986);
xor U6382 (N_6382,N_4892,N_5119);
nand U6383 (N_6383,N_5187,N_4866);
xor U6384 (N_6384,N_5453,N_5425);
xnor U6385 (N_6385,N_5773,N_5084);
or U6386 (N_6386,N_5109,N_5031);
xor U6387 (N_6387,N_5203,N_5303);
or U6388 (N_6388,N_5891,N_5305);
xnor U6389 (N_6389,N_5150,N_5409);
xor U6390 (N_6390,N_4861,N_5111);
xor U6391 (N_6391,N_4913,N_5765);
and U6392 (N_6392,N_4921,N_5136);
and U6393 (N_6393,N_5794,N_5567);
and U6394 (N_6394,N_5246,N_5254);
nand U6395 (N_6395,N_5074,N_4957);
nand U6396 (N_6396,N_5976,N_5212);
or U6397 (N_6397,N_5104,N_5279);
xor U6398 (N_6398,N_4842,N_5415);
xnor U6399 (N_6399,N_5152,N_4910);
nand U6400 (N_6400,N_5554,N_5564);
nand U6401 (N_6401,N_5809,N_5698);
and U6402 (N_6402,N_4851,N_5288);
nand U6403 (N_6403,N_5452,N_5531);
nand U6404 (N_6404,N_5320,N_5776);
nor U6405 (N_6405,N_5295,N_5173);
nand U6406 (N_6406,N_5430,N_4849);
xnor U6407 (N_6407,N_5044,N_5171);
xor U6408 (N_6408,N_5338,N_5105);
or U6409 (N_6409,N_4817,N_5082);
xnor U6410 (N_6410,N_5525,N_5322);
and U6411 (N_6411,N_5763,N_5699);
nand U6412 (N_6412,N_5502,N_5530);
xnor U6413 (N_6413,N_4904,N_5533);
and U6414 (N_6414,N_5640,N_5771);
and U6415 (N_6415,N_4877,N_5145);
nor U6416 (N_6416,N_5777,N_5941);
or U6417 (N_6417,N_5637,N_5112);
or U6418 (N_6418,N_4938,N_5652);
nor U6419 (N_6419,N_5872,N_5750);
nand U6420 (N_6420,N_5646,N_5365);
xnor U6421 (N_6421,N_4854,N_5733);
nor U6422 (N_6422,N_5205,N_5542);
nand U6423 (N_6423,N_5899,N_4944);
and U6424 (N_6424,N_5107,N_5275);
nand U6425 (N_6425,N_5586,N_5041);
and U6426 (N_6426,N_5185,N_5154);
or U6427 (N_6427,N_5973,N_5878);
and U6428 (N_6428,N_5472,N_5648);
and U6429 (N_6429,N_5416,N_5579);
xor U6430 (N_6430,N_5883,N_5635);
xor U6431 (N_6431,N_5539,N_4983);
nor U6432 (N_6432,N_5241,N_5097);
or U6433 (N_6433,N_5784,N_5732);
and U6434 (N_6434,N_5169,N_5466);
or U6435 (N_6435,N_5790,N_5788);
and U6436 (N_6436,N_5139,N_5349);
xor U6437 (N_6437,N_5933,N_5300);
and U6438 (N_6438,N_5493,N_5222);
xor U6439 (N_6439,N_5760,N_5242);
nor U6440 (N_6440,N_5381,N_4979);
nand U6441 (N_6441,N_4939,N_5289);
xor U6442 (N_6442,N_5612,N_5007);
or U6443 (N_6443,N_5204,N_5290);
xor U6444 (N_6444,N_5034,N_5739);
and U6445 (N_6445,N_5061,N_5497);
nand U6446 (N_6446,N_5953,N_4830);
xnor U6447 (N_6447,N_5217,N_4953);
nand U6448 (N_6448,N_5882,N_5144);
or U6449 (N_6449,N_5020,N_5566);
nand U6450 (N_6450,N_5621,N_4829);
nand U6451 (N_6451,N_5348,N_5465);
xnor U6452 (N_6452,N_5821,N_5622);
nor U6453 (N_6453,N_5936,N_5678);
nand U6454 (N_6454,N_5862,N_4886);
or U6455 (N_6455,N_4930,N_5920);
xnor U6456 (N_6456,N_5101,N_5834);
and U6457 (N_6457,N_5553,N_5998);
nor U6458 (N_6458,N_5574,N_5917);
nor U6459 (N_6459,N_4831,N_5293);
or U6460 (N_6460,N_5803,N_5655);
nand U6461 (N_6461,N_5517,N_5962);
or U6462 (N_6462,N_5839,N_5315);
xnor U6463 (N_6463,N_5032,N_4946);
or U6464 (N_6464,N_5938,N_4977);
nor U6465 (N_6465,N_5634,N_5417);
nand U6466 (N_6466,N_5704,N_5060);
or U6467 (N_6467,N_5076,N_4915);
and U6468 (N_6468,N_5198,N_5202);
or U6469 (N_6469,N_5931,N_5710);
nor U6470 (N_6470,N_5644,N_5372);
nor U6471 (N_6471,N_5193,N_5719);
nor U6472 (N_6472,N_5157,N_5858);
and U6473 (N_6473,N_5731,N_5053);
and U6474 (N_6474,N_5385,N_5967);
nand U6475 (N_6475,N_5666,N_5753);
nand U6476 (N_6476,N_4801,N_5971);
xor U6477 (N_6477,N_5956,N_4816);
xor U6478 (N_6478,N_5693,N_5467);
xor U6479 (N_6479,N_5448,N_5686);
and U6480 (N_6480,N_5446,N_5219);
nand U6481 (N_6481,N_5066,N_5555);
nor U6482 (N_6482,N_5002,N_5768);
nand U6483 (N_6483,N_5747,N_5894);
nor U6484 (N_6484,N_5110,N_4960);
or U6485 (N_6485,N_4973,N_5630);
nand U6486 (N_6486,N_5089,N_5114);
xnor U6487 (N_6487,N_5419,N_5256);
xor U6488 (N_6488,N_5815,N_5994);
nand U6489 (N_6489,N_5726,N_4835);
nand U6490 (N_6490,N_4868,N_5547);
and U6491 (N_6491,N_5990,N_4845);
or U6492 (N_6492,N_5572,N_5389);
xor U6493 (N_6493,N_4882,N_4958);
or U6494 (N_6494,N_5257,N_5012);
nor U6495 (N_6495,N_5412,N_4833);
and U6496 (N_6496,N_5476,N_5403);
xor U6497 (N_6497,N_5909,N_5818);
or U6498 (N_6498,N_5826,N_5695);
nor U6499 (N_6499,N_5676,N_5851);
xor U6500 (N_6500,N_5228,N_5565);
or U6501 (N_6501,N_5683,N_5867);
or U6502 (N_6502,N_5311,N_5117);
and U6503 (N_6503,N_5285,N_5359);
or U6504 (N_6504,N_5486,N_4947);
or U6505 (N_6505,N_5124,N_5598);
and U6506 (N_6506,N_5377,N_5098);
or U6507 (N_6507,N_5167,N_5168);
and U6508 (N_6508,N_5276,N_5580);
xnor U6509 (N_6509,N_5055,N_5057);
xnor U6510 (N_6510,N_5021,N_4896);
nand U6511 (N_6511,N_5557,N_5408);
nor U6512 (N_6512,N_5605,N_5757);
nor U6513 (N_6513,N_4850,N_5341);
nor U6514 (N_6514,N_4936,N_5922);
nand U6515 (N_6515,N_5808,N_5692);
or U6516 (N_6516,N_5038,N_5484);
nor U6517 (N_6517,N_5260,N_5433);
xnor U6518 (N_6518,N_5485,N_5870);
and U6519 (N_6519,N_5494,N_5793);
and U6520 (N_6520,N_5024,N_5384);
and U6521 (N_6521,N_5663,N_5503);
and U6522 (N_6522,N_5482,N_4972);
or U6523 (N_6523,N_5046,N_5954);
and U6524 (N_6524,N_5888,N_5968);
xnor U6525 (N_6525,N_5654,N_5286);
xnor U6526 (N_6526,N_5658,N_5817);
or U6527 (N_6527,N_5615,N_5043);
or U6528 (N_6528,N_5740,N_5248);
nor U6529 (N_6529,N_4965,N_5015);
or U6530 (N_6530,N_5702,N_5102);
or U6531 (N_6531,N_5210,N_5969);
and U6532 (N_6532,N_5059,N_5460);
xor U6533 (N_6533,N_5549,N_5498);
nand U6534 (N_6534,N_4963,N_4903);
nor U6535 (N_6535,N_5106,N_5062);
xnor U6536 (N_6536,N_5378,N_5659);
nor U6537 (N_6537,N_5367,N_5778);
and U6538 (N_6538,N_5690,N_5314);
and U6539 (N_6539,N_5281,N_4825);
xor U6540 (N_6540,N_5949,N_5237);
xnor U6541 (N_6541,N_5915,N_5432);
and U6542 (N_6542,N_5616,N_5000);
xor U6543 (N_6543,N_5443,N_4860);
and U6544 (N_6544,N_5299,N_4917);
and U6545 (N_6545,N_5573,N_5083);
and U6546 (N_6546,N_5754,N_5508);
xor U6547 (N_6547,N_5319,N_5495);
xnor U6548 (N_6548,N_5058,N_5420);
xnor U6549 (N_6549,N_5781,N_5070);
and U6550 (N_6550,N_5838,N_4997);
nand U6551 (N_6551,N_5274,N_5194);
and U6552 (N_6552,N_5398,N_5191);
nand U6553 (N_6553,N_4988,N_5442);
and U6554 (N_6554,N_5033,N_5614);
nand U6555 (N_6555,N_4818,N_5078);
nor U6556 (N_6556,N_5982,N_5625);
or U6557 (N_6557,N_5345,N_5513);
nand U6558 (N_6558,N_5213,N_5989);
or U6559 (N_6559,N_5336,N_5935);
nand U6560 (N_6560,N_5819,N_5946);
xnor U6561 (N_6561,N_4810,N_5642);
and U6562 (N_6562,N_5800,N_5023);
nand U6563 (N_6563,N_5273,N_5297);
xor U6564 (N_6564,N_5386,N_5536);
and U6565 (N_6565,N_5885,N_5764);
xnor U6566 (N_6566,N_5094,N_5220);
xor U6567 (N_6567,N_5512,N_5444);
nand U6568 (N_6568,N_5932,N_5158);
xnor U6569 (N_6569,N_5353,N_5302);
or U6570 (N_6570,N_5414,N_5480);
xnor U6571 (N_6571,N_5334,N_5428);
nand U6572 (N_6572,N_5672,N_5093);
xnor U6573 (N_6573,N_5907,N_5014);
nand U6574 (N_6574,N_5662,N_5901);
or U6575 (N_6575,N_5904,N_5524);
nand U6576 (N_6576,N_5236,N_4804);
xor U6577 (N_6577,N_5108,N_4887);
nor U6578 (N_6578,N_5997,N_5805);
and U6579 (N_6579,N_5703,N_5133);
and U6580 (N_6580,N_5180,N_4967);
or U6581 (N_6581,N_5836,N_5604);
nand U6582 (N_6582,N_5890,N_5723);
or U6583 (N_6583,N_5505,N_4879);
and U6584 (N_6584,N_4878,N_5380);
or U6585 (N_6585,N_5087,N_5814);
nor U6586 (N_6586,N_5049,N_5240);
or U6587 (N_6587,N_5492,N_5643);
xnor U6588 (N_6588,N_5509,N_5230);
or U6589 (N_6589,N_5233,N_5796);
nand U6590 (N_6590,N_5357,N_4899);
nand U6591 (N_6591,N_4990,N_4894);
xnor U6592 (N_6592,N_5326,N_5545);
or U6593 (N_6593,N_5308,N_4976);
and U6594 (N_6594,N_5908,N_5550);
or U6595 (N_6595,N_5234,N_5507);
nor U6596 (N_6596,N_4819,N_4824);
nand U6597 (N_6597,N_5387,N_5134);
nor U6598 (N_6598,N_5963,N_5149);
nand U6599 (N_6599,N_5993,N_4870);
xnor U6600 (N_6600,N_5564,N_5002);
nand U6601 (N_6601,N_5277,N_4866);
nor U6602 (N_6602,N_5966,N_5742);
or U6603 (N_6603,N_5652,N_5708);
nand U6604 (N_6604,N_4934,N_5754);
and U6605 (N_6605,N_5738,N_4894);
or U6606 (N_6606,N_5021,N_5514);
and U6607 (N_6607,N_5381,N_5819);
or U6608 (N_6608,N_5716,N_5602);
nor U6609 (N_6609,N_5124,N_5739);
nand U6610 (N_6610,N_5842,N_5986);
xor U6611 (N_6611,N_5220,N_5229);
nand U6612 (N_6612,N_5817,N_5297);
xnor U6613 (N_6613,N_5408,N_5238);
nand U6614 (N_6614,N_5305,N_4904);
nor U6615 (N_6615,N_5522,N_5239);
nor U6616 (N_6616,N_5476,N_5897);
nand U6617 (N_6617,N_5837,N_5628);
and U6618 (N_6618,N_5508,N_5648);
xor U6619 (N_6619,N_5162,N_5845);
nand U6620 (N_6620,N_5357,N_5766);
or U6621 (N_6621,N_5210,N_5793);
nand U6622 (N_6622,N_5326,N_5885);
nor U6623 (N_6623,N_5698,N_5751);
and U6624 (N_6624,N_5346,N_5150);
xnor U6625 (N_6625,N_5283,N_5122);
nor U6626 (N_6626,N_4911,N_4954);
nor U6627 (N_6627,N_5732,N_5132);
nor U6628 (N_6628,N_5161,N_4912);
nand U6629 (N_6629,N_5731,N_5229);
and U6630 (N_6630,N_5684,N_4980);
xor U6631 (N_6631,N_5760,N_5978);
xnor U6632 (N_6632,N_5671,N_5957);
or U6633 (N_6633,N_5090,N_5948);
nand U6634 (N_6634,N_5967,N_5201);
or U6635 (N_6635,N_5680,N_5253);
or U6636 (N_6636,N_5316,N_5639);
xor U6637 (N_6637,N_5441,N_5256);
nand U6638 (N_6638,N_5238,N_5773);
nor U6639 (N_6639,N_4909,N_4990);
xnor U6640 (N_6640,N_5113,N_5997);
xor U6641 (N_6641,N_5291,N_5599);
or U6642 (N_6642,N_5423,N_5696);
or U6643 (N_6643,N_5749,N_5637);
xnor U6644 (N_6644,N_5282,N_4869);
and U6645 (N_6645,N_5255,N_5592);
nand U6646 (N_6646,N_5551,N_5230);
nor U6647 (N_6647,N_4856,N_5592);
and U6648 (N_6648,N_5434,N_5361);
or U6649 (N_6649,N_5957,N_5081);
or U6650 (N_6650,N_5035,N_5477);
xor U6651 (N_6651,N_5032,N_5309);
nand U6652 (N_6652,N_5304,N_5692);
or U6653 (N_6653,N_5639,N_5381);
xor U6654 (N_6654,N_4978,N_5689);
nand U6655 (N_6655,N_5791,N_5730);
nor U6656 (N_6656,N_5083,N_5001);
nand U6657 (N_6657,N_4915,N_5363);
or U6658 (N_6658,N_5707,N_4940);
nand U6659 (N_6659,N_4983,N_4832);
xor U6660 (N_6660,N_5734,N_5775);
and U6661 (N_6661,N_5710,N_4918);
nor U6662 (N_6662,N_5139,N_5172);
xnor U6663 (N_6663,N_5230,N_5638);
nor U6664 (N_6664,N_4864,N_4902);
and U6665 (N_6665,N_5747,N_5087);
nor U6666 (N_6666,N_5528,N_4859);
xnor U6667 (N_6667,N_5812,N_5623);
xor U6668 (N_6668,N_5202,N_5437);
and U6669 (N_6669,N_5380,N_5806);
and U6670 (N_6670,N_5875,N_5209);
or U6671 (N_6671,N_5360,N_5054);
nand U6672 (N_6672,N_5000,N_5642);
nand U6673 (N_6673,N_5780,N_5091);
nand U6674 (N_6674,N_4817,N_4969);
nor U6675 (N_6675,N_5335,N_5402);
xnor U6676 (N_6676,N_5814,N_4946);
nor U6677 (N_6677,N_5315,N_5999);
xnor U6678 (N_6678,N_4994,N_5404);
nor U6679 (N_6679,N_5875,N_5912);
nor U6680 (N_6680,N_5603,N_5549);
xnor U6681 (N_6681,N_5042,N_5998);
nor U6682 (N_6682,N_5284,N_5319);
and U6683 (N_6683,N_5525,N_5218);
xnor U6684 (N_6684,N_5770,N_5959);
nand U6685 (N_6685,N_4851,N_4982);
and U6686 (N_6686,N_5282,N_5505);
or U6687 (N_6687,N_5306,N_5330);
or U6688 (N_6688,N_5890,N_5984);
nor U6689 (N_6689,N_5196,N_4876);
nand U6690 (N_6690,N_5660,N_5427);
xnor U6691 (N_6691,N_5444,N_5557);
xor U6692 (N_6692,N_5220,N_4846);
xnor U6693 (N_6693,N_5024,N_5240);
or U6694 (N_6694,N_5015,N_4986);
nor U6695 (N_6695,N_5005,N_5130);
or U6696 (N_6696,N_5269,N_5125);
and U6697 (N_6697,N_5681,N_5351);
or U6698 (N_6698,N_5857,N_5413);
or U6699 (N_6699,N_5600,N_4910);
nor U6700 (N_6700,N_5781,N_5400);
nand U6701 (N_6701,N_5736,N_5158);
nand U6702 (N_6702,N_5598,N_5771);
nand U6703 (N_6703,N_4877,N_5577);
nand U6704 (N_6704,N_5751,N_5856);
or U6705 (N_6705,N_5832,N_5989);
nor U6706 (N_6706,N_5613,N_5092);
and U6707 (N_6707,N_5343,N_5676);
and U6708 (N_6708,N_5503,N_5649);
nand U6709 (N_6709,N_5983,N_5434);
nor U6710 (N_6710,N_5030,N_4862);
nand U6711 (N_6711,N_5246,N_5840);
nor U6712 (N_6712,N_5723,N_4934);
nand U6713 (N_6713,N_5561,N_5295);
or U6714 (N_6714,N_5428,N_5056);
nor U6715 (N_6715,N_5709,N_5065);
and U6716 (N_6716,N_4960,N_5604);
xnor U6717 (N_6717,N_5319,N_5441);
nor U6718 (N_6718,N_5564,N_5991);
or U6719 (N_6719,N_5213,N_5407);
xnor U6720 (N_6720,N_5049,N_5268);
or U6721 (N_6721,N_4855,N_5353);
nand U6722 (N_6722,N_4933,N_4950);
nand U6723 (N_6723,N_5149,N_5310);
or U6724 (N_6724,N_5575,N_5931);
or U6725 (N_6725,N_5877,N_5623);
xnor U6726 (N_6726,N_4955,N_4984);
nand U6727 (N_6727,N_5833,N_5956);
xor U6728 (N_6728,N_5410,N_5636);
nor U6729 (N_6729,N_5896,N_4951);
nand U6730 (N_6730,N_5757,N_5645);
and U6731 (N_6731,N_5917,N_5915);
and U6732 (N_6732,N_5679,N_5450);
or U6733 (N_6733,N_5951,N_4946);
nand U6734 (N_6734,N_5196,N_4978);
nand U6735 (N_6735,N_5591,N_5636);
nor U6736 (N_6736,N_5421,N_5651);
and U6737 (N_6737,N_5248,N_5712);
nand U6738 (N_6738,N_5934,N_4803);
nor U6739 (N_6739,N_5316,N_5416);
nand U6740 (N_6740,N_5978,N_5807);
xor U6741 (N_6741,N_5464,N_5135);
or U6742 (N_6742,N_5724,N_5423);
xor U6743 (N_6743,N_5772,N_5998);
and U6744 (N_6744,N_4914,N_5850);
xnor U6745 (N_6745,N_5568,N_4999);
nor U6746 (N_6746,N_5436,N_4903);
xor U6747 (N_6747,N_4932,N_5695);
and U6748 (N_6748,N_4964,N_5911);
and U6749 (N_6749,N_5727,N_4944);
nand U6750 (N_6750,N_5372,N_5613);
xnor U6751 (N_6751,N_5503,N_5947);
or U6752 (N_6752,N_5357,N_5866);
nor U6753 (N_6753,N_5316,N_5570);
nand U6754 (N_6754,N_4804,N_5010);
nor U6755 (N_6755,N_5485,N_5204);
and U6756 (N_6756,N_5928,N_5431);
and U6757 (N_6757,N_5312,N_5507);
nor U6758 (N_6758,N_5336,N_5838);
nand U6759 (N_6759,N_5815,N_5108);
nor U6760 (N_6760,N_5512,N_5866);
nor U6761 (N_6761,N_5044,N_5090);
xor U6762 (N_6762,N_5558,N_5937);
nor U6763 (N_6763,N_5757,N_4899);
and U6764 (N_6764,N_5980,N_5832);
nand U6765 (N_6765,N_5451,N_5948);
nand U6766 (N_6766,N_5845,N_5645);
nand U6767 (N_6767,N_5394,N_5279);
or U6768 (N_6768,N_5792,N_5638);
xnor U6769 (N_6769,N_5676,N_5703);
and U6770 (N_6770,N_5591,N_5457);
nand U6771 (N_6771,N_5129,N_4946);
and U6772 (N_6772,N_5896,N_5573);
nand U6773 (N_6773,N_5226,N_5506);
or U6774 (N_6774,N_4861,N_5880);
and U6775 (N_6775,N_5844,N_4959);
and U6776 (N_6776,N_5830,N_5094);
nand U6777 (N_6777,N_5734,N_5190);
xnor U6778 (N_6778,N_5134,N_5314);
xnor U6779 (N_6779,N_5632,N_4830);
or U6780 (N_6780,N_5328,N_5507);
or U6781 (N_6781,N_5589,N_5662);
and U6782 (N_6782,N_5778,N_5780);
xor U6783 (N_6783,N_4804,N_5131);
nand U6784 (N_6784,N_5287,N_5538);
nand U6785 (N_6785,N_4997,N_5834);
nor U6786 (N_6786,N_5828,N_5287);
and U6787 (N_6787,N_5954,N_5259);
xnor U6788 (N_6788,N_5139,N_4975);
and U6789 (N_6789,N_5676,N_5963);
or U6790 (N_6790,N_5065,N_5446);
or U6791 (N_6791,N_4985,N_5862);
or U6792 (N_6792,N_4825,N_5594);
xnor U6793 (N_6793,N_5487,N_5396);
or U6794 (N_6794,N_5767,N_5592);
xor U6795 (N_6795,N_5766,N_5851);
xnor U6796 (N_6796,N_5858,N_5013);
and U6797 (N_6797,N_4812,N_5662);
nand U6798 (N_6798,N_5314,N_4826);
nor U6799 (N_6799,N_5953,N_5884);
nand U6800 (N_6800,N_5745,N_5194);
nand U6801 (N_6801,N_5274,N_5264);
xor U6802 (N_6802,N_5299,N_4996);
nand U6803 (N_6803,N_5412,N_5545);
nor U6804 (N_6804,N_5019,N_5227);
xnor U6805 (N_6805,N_4875,N_4820);
nand U6806 (N_6806,N_5514,N_5070);
nand U6807 (N_6807,N_5162,N_5286);
nor U6808 (N_6808,N_5004,N_4846);
xnor U6809 (N_6809,N_4849,N_5005);
xnor U6810 (N_6810,N_4801,N_5953);
xor U6811 (N_6811,N_5453,N_5607);
or U6812 (N_6812,N_5867,N_5714);
and U6813 (N_6813,N_5918,N_5974);
nor U6814 (N_6814,N_4939,N_4810);
xnor U6815 (N_6815,N_5571,N_5712);
nand U6816 (N_6816,N_5084,N_5995);
xor U6817 (N_6817,N_5844,N_5340);
or U6818 (N_6818,N_5695,N_5186);
nor U6819 (N_6819,N_5123,N_5137);
xnor U6820 (N_6820,N_5228,N_5961);
nand U6821 (N_6821,N_4813,N_5692);
xnor U6822 (N_6822,N_5106,N_5815);
or U6823 (N_6823,N_5798,N_5362);
xnor U6824 (N_6824,N_5558,N_5506);
nand U6825 (N_6825,N_5266,N_5216);
and U6826 (N_6826,N_5157,N_5158);
xnor U6827 (N_6827,N_5271,N_5526);
and U6828 (N_6828,N_5254,N_5782);
or U6829 (N_6829,N_5013,N_5689);
xor U6830 (N_6830,N_4991,N_5185);
nor U6831 (N_6831,N_5285,N_5251);
nand U6832 (N_6832,N_5597,N_4901);
and U6833 (N_6833,N_5928,N_5114);
nor U6834 (N_6834,N_5155,N_5305);
xor U6835 (N_6835,N_5103,N_5866);
and U6836 (N_6836,N_5650,N_5535);
and U6837 (N_6837,N_5544,N_5818);
nor U6838 (N_6838,N_5974,N_5867);
nand U6839 (N_6839,N_5183,N_5043);
xor U6840 (N_6840,N_5266,N_5338);
and U6841 (N_6841,N_5618,N_4964);
xnor U6842 (N_6842,N_5147,N_5642);
xor U6843 (N_6843,N_5863,N_5020);
or U6844 (N_6844,N_5370,N_4803);
nand U6845 (N_6845,N_5256,N_5930);
and U6846 (N_6846,N_5081,N_5372);
nand U6847 (N_6847,N_5864,N_5903);
nor U6848 (N_6848,N_5541,N_5304);
xnor U6849 (N_6849,N_4890,N_5785);
xnor U6850 (N_6850,N_5029,N_5921);
and U6851 (N_6851,N_5957,N_5580);
nor U6852 (N_6852,N_5071,N_5090);
or U6853 (N_6853,N_4942,N_5995);
xor U6854 (N_6854,N_5019,N_5861);
nand U6855 (N_6855,N_5980,N_5849);
xnor U6856 (N_6856,N_5059,N_5575);
nand U6857 (N_6857,N_4912,N_5759);
or U6858 (N_6858,N_5632,N_5548);
and U6859 (N_6859,N_5399,N_4961);
or U6860 (N_6860,N_5186,N_5853);
nand U6861 (N_6861,N_5026,N_5213);
nor U6862 (N_6862,N_4953,N_5681);
and U6863 (N_6863,N_5584,N_5434);
xor U6864 (N_6864,N_5667,N_5825);
or U6865 (N_6865,N_5612,N_5168);
xnor U6866 (N_6866,N_4831,N_5662);
or U6867 (N_6867,N_5865,N_5489);
nor U6868 (N_6868,N_5077,N_4801);
and U6869 (N_6869,N_5218,N_5519);
or U6870 (N_6870,N_5379,N_5178);
or U6871 (N_6871,N_5961,N_5189);
nand U6872 (N_6872,N_5175,N_5700);
and U6873 (N_6873,N_5605,N_5705);
or U6874 (N_6874,N_5534,N_4963);
nand U6875 (N_6875,N_4946,N_4877);
and U6876 (N_6876,N_5713,N_5954);
or U6877 (N_6877,N_5116,N_5175);
nor U6878 (N_6878,N_5817,N_5736);
nand U6879 (N_6879,N_5173,N_5033);
and U6880 (N_6880,N_5951,N_5956);
or U6881 (N_6881,N_5727,N_5360);
nand U6882 (N_6882,N_5956,N_5617);
nand U6883 (N_6883,N_5945,N_5695);
nand U6884 (N_6884,N_5677,N_5992);
and U6885 (N_6885,N_4963,N_5701);
nand U6886 (N_6886,N_5437,N_5448);
or U6887 (N_6887,N_5220,N_5513);
nand U6888 (N_6888,N_5712,N_5665);
or U6889 (N_6889,N_5554,N_5714);
nand U6890 (N_6890,N_5522,N_4956);
nand U6891 (N_6891,N_5261,N_5518);
xor U6892 (N_6892,N_5776,N_5118);
nor U6893 (N_6893,N_4871,N_4902);
nand U6894 (N_6894,N_5038,N_5097);
and U6895 (N_6895,N_4887,N_5954);
nor U6896 (N_6896,N_5089,N_5688);
and U6897 (N_6897,N_5947,N_4905);
nor U6898 (N_6898,N_4969,N_5130);
nor U6899 (N_6899,N_5380,N_5415);
xnor U6900 (N_6900,N_5271,N_5659);
xnor U6901 (N_6901,N_5272,N_5805);
or U6902 (N_6902,N_5150,N_5927);
nor U6903 (N_6903,N_4987,N_5452);
or U6904 (N_6904,N_4829,N_5367);
or U6905 (N_6905,N_5099,N_5338);
or U6906 (N_6906,N_5096,N_5637);
nor U6907 (N_6907,N_4831,N_5924);
and U6908 (N_6908,N_5413,N_4894);
or U6909 (N_6909,N_5888,N_4931);
nor U6910 (N_6910,N_5773,N_5611);
and U6911 (N_6911,N_4932,N_5551);
or U6912 (N_6912,N_5073,N_5495);
xnor U6913 (N_6913,N_5705,N_5018);
or U6914 (N_6914,N_5907,N_5371);
xnor U6915 (N_6915,N_5793,N_5892);
nand U6916 (N_6916,N_4938,N_5212);
nor U6917 (N_6917,N_5801,N_5848);
and U6918 (N_6918,N_5716,N_4903);
xnor U6919 (N_6919,N_4955,N_5332);
nor U6920 (N_6920,N_5169,N_5122);
or U6921 (N_6921,N_4899,N_5279);
xnor U6922 (N_6922,N_5902,N_4951);
or U6923 (N_6923,N_5839,N_4913);
nor U6924 (N_6924,N_5426,N_5662);
xnor U6925 (N_6925,N_4859,N_5445);
xor U6926 (N_6926,N_5848,N_5168);
xnor U6927 (N_6927,N_5170,N_5448);
nand U6928 (N_6928,N_5025,N_5725);
nor U6929 (N_6929,N_5444,N_5927);
or U6930 (N_6930,N_4842,N_5682);
xnor U6931 (N_6931,N_5604,N_4886);
nand U6932 (N_6932,N_5196,N_5661);
xnor U6933 (N_6933,N_5235,N_5076);
or U6934 (N_6934,N_4857,N_5822);
nor U6935 (N_6935,N_5812,N_4835);
nand U6936 (N_6936,N_5986,N_5415);
nor U6937 (N_6937,N_5110,N_5842);
nor U6938 (N_6938,N_4964,N_5700);
nor U6939 (N_6939,N_5663,N_5318);
and U6940 (N_6940,N_5239,N_5011);
or U6941 (N_6941,N_5097,N_5320);
nor U6942 (N_6942,N_5919,N_5842);
xor U6943 (N_6943,N_5251,N_5331);
or U6944 (N_6944,N_4923,N_5816);
and U6945 (N_6945,N_5199,N_5960);
or U6946 (N_6946,N_4877,N_5785);
nor U6947 (N_6947,N_5297,N_4900);
and U6948 (N_6948,N_5164,N_5300);
and U6949 (N_6949,N_5826,N_5110);
nand U6950 (N_6950,N_5653,N_5191);
xor U6951 (N_6951,N_4854,N_5320);
and U6952 (N_6952,N_4918,N_5865);
or U6953 (N_6953,N_4814,N_5097);
and U6954 (N_6954,N_5257,N_5451);
nor U6955 (N_6955,N_5019,N_5985);
nor U6956 (N_6956,N_5115,N_5099);
and U6957 (N_6957,N_5514,N_5929);
or U6958 (N_6958,N_5213,N_5637);
nor U6959 (N_6959,N_5781,N_5713);
xnor U6960 (N_6960,N_5804,N_5242);
nor U6961 (N_6961,N_5151,N_5869);
nor U6962 (N_6962,N_4993,N_5576);
and U6963 (N_6963,N_5221,N_5483);
nand U6964 (N_6964,N_5458,N_4858);
nand U6965 (N_6965,N_5499,N_4896);
nor U6966 (N_6966,N_5514,N_5804);
or U6967 (N_6967,N_5721,N_5824);
nand U6968 (N_6968,N_5698,N_4913);
nand U6969 (N_6969,N_5987,N_5996);
xor U6970 (N_6970,N_5502,N_5001);
xnor U6971 (N_6971,N_5714,N_5343);
nor U6972 (N_6972,N_5416,N_5936);
xnor U6973 (N_6973,N_5758,N_5520);
xor U6974 (N_6974,N_5519,N_5064);
xnor U6975 (N_6975,N_5064,N_5076);
or U6976 (N_6976,N_5043,N_5862);
xor U6977 (N_6977,N_5348,N_5210);
and U6978 (N_6978,N_5557,N_5046);
xor U6979 (N_6979,N_4924,N_5703);
xor U6980 (N_6980,N_5012,N_5979);
xor U6981 (N_6981,N_5682,N_5650);
nand U6982 (N_6982,N_5433,N_5038);
xnor U6983 (N_6983,N_4814,N_5489);
and U6984 (N_6984,N_5337,N_5592);
and U6985 (N_6985,N_4856,N_5395);
nor U6986 (N_6986,N_4939,N_5565);
and U6987 (N_6987,N_5770,N_5481);
nand U6988 (N_6988,N_5526,N_5690);
and U6989 (N_6989,N_5928,N_4949);
xor U6990 (N_6990,N_5744,N_4853);
xor U6991 (N_6991,N_5257,N_5721);
and U6992 (N_6992,N_5609,N_5944);
nor U6993 (N_6993,N_5388,N_5030);
or U6994 (N_6994,N_5207,N_5254);
or U6995 (N_6995,N_5677,N_5006);
nand U6996 (N_6996,N_5805,N_5644);
or U6997 (N_6997,N_5751,N_5836);
and U6998 (N_6998,N_4807,N_5577);
nand U6999 (N_6999,N_5006,N_5269);
and U7000 (N_7000,N_4884,N_5485);
xnor U7001 (N_7001,N_5547,N_5793);
or U7002 (N_7002,N_5358,N_5178);
xor U7003 (N_7003,N_5798,N_5860);
xnor U7004 (N_7004,N_5248,N_5548);
and U7005 (N_7005,N_5039,N_5248);
and U7006 (N_7006,N_5732,N_4957);
and U7007 (N_7007,N_4991,N_5549);
xor U7008 (N_7008,N_4891,N_5553);
nor U7009 (N_7009,N_5050,N_5923);
and U7010 (N_7010,N_5751,N_5892);
nor U7011 (N_7011,N_5002,N_5221);
or U7012 (N_7012,N_5969,N_5233);
nor U7013 (N_7013,N_5165,N_5834);
and U7014 (N_7014,N_5584,N_5912);
nand U7015 (N_7015,N_5884,N_5017);
and U7016 (N_7016,N_5118,N_4840);
nand U7017 (N_7017,N_5643,N_5268);
xnor U7018 (N_7018,N_5421,N_5909);
or U7019 (N_7019,N_4993,N_4864);
and U7020 (N_7020,N_5894,N_5661);
and U7021 (N_7021,N_5747,N_5136);
xnor U7022 (N_7022,N_5254,N_5687);
or U7023 (N_7023,N_5337,N_5078);
xor U7024 (N_7024,N_5636,N_5748);
or U7025 (N_7025,N_5309,N_5373);
and U7026 (N_7026,N_5879,N_5554);
xor U7027 (N_7027,N_5283,N_5446);
or U7028 (N_7028,N_5613,N_5444);
xor U7029 (N_7029,N_5394,N_5146);
xor U7030 (N_7030,N_5218,N_5472);
xnor U7031 (N_7031,N_5190,N_5852);
nor U7032 (N_7032,N_5300,N_5954);
nor U7033 (N_7033,N_5615,N_5554);
nand U7034 (N_7034,N_5210,N_5734);
nor U7035 (N_7035,N_5219,N_5321);
nand U7036 (N_7036,N_5092,N_5827);
xor U7037 (N_7037,N_4814,N_5685);
nand U7038 (N_7038,N_5911,N_5824);
nor U7039 (N_7039,N_5891,N_5001);
nand U7040 (N_7040,N_5879,N_5015);
xor U7041 (N_7041,N_5440,N_4879);
nor U7042 (N_7042,N_5721,N_5570);
nor U7043 (N_7043,N_5272,N_5196);
or U7044 (N_7044,N_5686,N_5397);
nor U7045 (N_7045,N_4963,N_5560);
nand U7046 (N_7046,N_5667,N_5236);
or U7047 (N_7047,N_5636,N_5308);
nand U7048 (N_7048,N_4906,N_5633);
and U7049 (N_7049,N_5662,N_4932);
xor U7050 (N_7050,N_5962,N_5839);
xnor U7051 (N_7051,N_5228,N_5185);
nand U7052 (N_7052,N_5425,N_5905);
xor U7053 (N_7053,N_5286,N_5895);
nor U7054 (N_7054,N_5493,N_5571);
nor U7055 (N_7055,N_5713,N_5898);
nand U7056 (N_7056,N_5991,N_5735);
nand U7057 (N_7057,N_4829,N_4896);
xor U7058 (N_7058,N_5374,N_4824);
nor U7059 (N_7059,N_5986,N_5089);
and U7060 (N_7060,N_5650,N_5478);
nand U7061 (N_7061,N_4853,N_4872);
or U7062 (N_7062,N_5523,N_5082);
and U7063 (N_7063,N_5386,N_5550);
and U7064 (N_7064,N_5761,N_5654);
nor U7065 (N_7065,N_5411,N_5190);
or U7066 (N_7066,N_5426,N_5663);
nor U7067 (N_7067,N_5342,N_5694);
and U7068 (N_7068,N_5673,N_5161);
and U7069 (N_7069,N_4981,N_5120);
xor U7070 (N_7070,N_5838,N_5784);
and U7071 (N_7071,N_4934,N_5069);
xor U7072 (N_7072,N_5428,N_5481);
nor U7073 (N_7073,N_5876,N_5699);
xnor U7074 (N_7074,N_5348,N_4953);
xor U7075 (N_7075,N_5401,N_5476);
nand U7076 (N_7076,N_5585,N_5714);
xnor U7077 (N_7077,N_5037,N_5564);
and U7078 (N_7078,N_5237,N_5347);
nand U7079 (N_7079,N_5254,N_5294);
or U7080 (N_7080,N_5531,N_5494);
xor U7081 (N_7081,N_5607,N_5413);
nor U7082 (N_7082,N_5714,N_5028);
xnor U7083 (N_7083,N_4990,N_5460);
nor U7084 (N_7084,N_5376,N_5268);
or U7085 (N_7085,N_5889,N_5243);
nor U7086 (N_7086,N_5933,N_5944);
and U7087 (N_7087,N_4911,N_5369);
or U7088 (N_7088,N_5585,N_5732);
nor U7089 (N_7089,N_5632,N_5096);
xor U7090 (N_7090,N_4994,N_5753);
or U7091 (N_7091,N_4931,N_5923);
xnor U7092 (N_7092,N_4974,N_5453);
and U7093 (N_7093,N_5909,N_5934);
nor U7094 (N_7094,N_5361,N_5373);
and U7095 (N_7095,N_5109,N_5095);
or U7096 (N_7096,N_5967,N_5523);
xor U7097 (N_7097,N_5064,N_4936);
nor U7098 (N_7098,N_4864,N_4933);
and U7099 (N_7099,N_5026,N_5524);
nand U7100 (N_7100,N_5599,N_5030);
and U7101 (N_7101,N_5838,N_4814);
nand U7102 (N_7102,N_5623,N_5958);
xnor U7103 (N_7103,N_5747,N_5815);
and U7104 (N_7104,N_5284,N_5361);
and U7105 (N_7105,N_5215,N_5273);
nand U7106 (N_7106,N_5925,N_5468);
nor U7107 (N_7107,N_5661,N_4987);
or U7108 (N_7108,N_5471,N_4989);
or U7109 (N_7109,N_5336,N_5494);
and U7110 (N_7110,N_5385,N_5634);
nand U7111 (N_7111,N_5095,N_5635);
nand U7112 (N_7112,N_5390,N_5394);
nand U7113 (N_7113,N_5874,N_5562);
nand U7114 (N_7114,N_5563,N_4896);
xor U7115 (N_7115,N_5733,N_5030);
nand U7116 (N_7116,N_5800,N_5661);
nor U7117 (N_7117,N_5860,N_5801);
nand U7118 (N_7118,N_5254,N_4973);
and U7119 (N_7119,N_5392,N_5877);
xor U7120 (N_7120,N_5873,N_5413);
xnor U7121 (N_7121,N_5249,N_5634);
and U7122 (N_7122,N_5348,N_5646);
or U7123 (N_7123,N_5204,N_5492);
nor U7124 (N_7124,N_5595,N_5424);
nor U7125 (N_7125,N_5270,N_5123);
or U7126 (N_7126,N_5208,N_5764);
nand U7127 (N_7127,N_5382,N_5746);
nand U7128 (N_7128,N_5743,N_5314);
xnor U7129 (N_7129,N_5898,N_5012);
xor U7130 (N_7130,N_5183,N_5180);
and U7131 (N_7131,N_5360,N_5121);
xnor U7132 (N_7132,N_5881,N_5935);
nand U7133 (N_7133,N_5918,N_4907);
nand U7134 (N_7134,N_5483,N_5449);
nand U7135 (N_7135,N_5755,N_4837);
or U7136 (N_7136,N_5185,N_5311);
nor U7137 (N_7137,N_5090,N_5450);
nor U7138 (N_7138,N_5043,N_5607);
xor U7139 (N_7139,N_5569,N_5365);
or U7140 (N_7140,N_5232,N_5657);
xnor U7141 (N_7141,N_5299,N_4993);
nor U7142 (N_7142,N_5746,N_5839);
xnor U7143 (N_7143,N_5202,N_5743);
nor U7144 (N_7144,N_5833,N_5688);
xnor U7145 (N_7145,N_5118,N_5752);
nand U7146 (N_7146,N_5460,N_5087);
nor U7147 (N_7147,N_5463,N_5712);
and U7148 (N_7148,N_5083,N_5741);
nand U7149 (N_7149,N_5937,N_5988);
xor U7150 (N_7150,N_5035,N_5174);
nor U7151 (N_7151,N_5426,N_5408);
or U7152 (N_7152,N_5246,N_5116);
and U7153 (N_7153,N_5725,N_5632);
and U7154 (N_7154,N_4952,N_5121);
xor U7155 (N_7155,N_5615,N_4872);
nand U7156 (N_7156,N_5884,N_4943);
and U7157 (N_7157,N_5667,N_4832);
or U7158 (N_7158,N_5473,N_5136);
nand U7159 (N_7159,N_5021,N_5512);
nor U7160 (N_7160,N_5194,N_5080);
nand U7161 (N_7161,N_5757,N_5195);
nor U7162 (N_7162,N_5259,N_4996);
and U7163 (N_7163,N_5389,N_5365);
xor U7164 (N_7164,N_5259,N_5407);
and U7165 (N_7165,N_5164,N_5735);
xor U7166 (N_7166,N_5811,N_5627);
nand U7167 (N_7167,N_4934,N_5163);
and U7168 (N_7168,N_5387,N_5796);
and U7169 (N_7169,N_5910,N_5304);
and U7170 (N_7170,N_5391,N_5070);
xnor U7171 (N_7171,N_5744,N_5153);
or U7172 (N_7172,N_5630,N_4866);
or U7173 (N_7173,N_5893,N_5660);
xor U7174 (N_7174,N_5703,N_5301);
xnor U7175 (N_7175,N_4866,N_4833);
nand U7176 (N_7176,N_5809,N_4859);
nor U7177 (N_7177,N_5309,N_5686);
or U7178 (N_7178,N_4991,N_5357);
nand U7179 (N_7179,N_5549,N_5750);
xnor U7180 (N_7180,N_5397,N_5046);
xor U7181 (N_7181,N_5905,N_5782);
nor U7182 (N_7182,N_5107,N_5851);
and U7183 (N_7183,N_5823,N_5718);
or U7184 (N_7184,N_5404,N_5997);
nor U7185 (N_7185,N_5712,N_5561);
nor U7186 (N_7186,N_4958,N_5805);
and U7187 (N_7187,N_5988,N_4914);
or U7188 (N_7188,N_5526,N_4890);
nand U7189 (N_7189,N_5862,N_5710);
and U7190 (N_7190,N_5623,N_5283);
xor U7191 (N_7191,N_4963,N_5496);
nand U7192 (N_7192,N_5769,N_5007);
nor U7193 (N_7193,N_5562,N_5141);
xnor U7194 (N_7194,N_5905,N_5250);
and U7195 (N_7195,N_5464,N_5187);
and U7196 (N_7196,N_4812,N_4993);
nand U7197 (N_7197,N_5215,N_5222);
and U7198 (N_7198,N_5968,N_5445);
and U7199 (N_7199,N_4859,N_5689);
or U7200 (N_7200,N_6304,N_6144);
nor U7201 (N_7201,N_6604,N_7074);
and U7202 (N_7202,N_7149,N_6275);
nand U7203 (N_7203,N_6241,N_7086);
and U7204 (N_7204,N_6606,N_6184);
or U7205 (N_7205,N_6735,N_7189);
nor U7206 (N_7206,N_6871,N_6753);
and U7207 (N_7207,N_7010,N_7186);
or U7208 (N_7208,N_7005,N_6896);
and U7209 (N_7209,N_6398,N_6347);
nor U7210 (N_7210,N_6028,N_6808);
nand U7211 (N_7211,N_6927,N_7187);
xnor U7212 (N_7212,N_6107,N_7131);
xor U7213 (N_7213,N_6375,N_6907);
xnor U7214 (N_7214,N_6553,N_6024);
nor U7215 (N_7215,N_6039,N_6282);
or U7216 (N_7216,N_6548,N_6115);
and U7217 (N_7217,N_6605,N_6888);
nand U7218 (N_7218,N_6953,N_6861);
and U7219 (N_7219,N_6092,N_6578);
xor U7220 (N_7220,N_7178,N_6051);
xor U7221 (N_7221,N_6483,N_6038);
xor U7222 (N_7222,N_6854,N_6166);
nand U7223 (N_7223,N_7165,N_7160);
nand U7224 (N_7224,N_6392,N_6488);
xor U7225 (N_7225,N_6295,N_6732);
nor U7226 (N_7226,N_6614,N_7015);
and U7227 (N_7227,N_6187,N_6758);
and U7228 (N_7228,N_7112,N_6248);
or U7229 (N_7229,N_6318,N_6586);
nand U7230 (N_7230,N_6119,N_6780);
nand U7231 (N_7231,N_7142,N_6394);
and U7232 (N_7232,N_6105,N_7124);
and U7233 (N_7233,N_7105,N_6091);
xnor U7234 (N_7234,N_6499,N_7058);
or U7235 (N_7235,N_6078,N_7147);
nor U7236 (N_7236,N_6710,N_6910);
nor U7237 (N_7237,N_7044,N_6154);
nor U7238 (N_7238,N_6445,N_6147);
or U7239 (N_7239,N_6273,N_6243);
nand U7240 (N_7240,N_6058,N_6169);
and U7241 (N_7241,N_6164,N_6460);
or U7242 (N_7242,N_6934,N_6151);
nand U7243 (N_7243,N_6066,N_6879);
nor U7244 (N_7244,N_6146,N_6431);
or U7245 (N_7245,N_6903,N_6810);
nor U7246 (N_7246,N_7113,N_6638);
xnor U7247 (N_7247,N_6189,N_7175);
nand U7248 (N_7248,N_6603,N_7084);
nand U7249 (N_7249,N_6377,N_6359);
and U7250 (N_7250,N_7130,N_6938);
or U7251 (N_7251,N_6484,N_6966);
and U7252 (N_7252,N_6986,N_6426);
xnor U7253 (N_7253,N_6912,N_6079);
nand U7254 (N_7254,N_6517,N_6372);
and U7255 (N_7255,N_6579,N_6531);
or U7256 (N_7256,N_6805,N_6286);
xnor U7257 (N_7257,N_6178,N_6836);
nand U7258 (N_7258,N_6800,N_6556);
nand U7259 (N_7259,N_7034,N_6723);
xor U7260 (N_7260,N_7066,N_6618);
or U7261 (N_7261,N_6900,N_6947);
nor U7262 (N_7262,N_6891,N_6408);
nand U7263 (N_7263,N_6190,N_6328);
nand U7264 (N_7264,N_6923,N_6150);
or U7265 (N_7265,N_6961,N_6737);
xor U7266 (N_7266,N_6519,N_6686);
nor U7267 (N_7267,N_6003,N_6706);
nor U7268 (N_7268,N_6873,N_6155);
xnor U7269 (N_7269,N_6380,N_6617);
or U7270 (N_7270,N_6532,N_6515);
nor U7271 (N_7271,N_6012,N_6346);
and U7272 (N_7272,N_6186,N_6133);
and U7273 (N_7273,N_7199,N_6235);
and U7274 (N_7274,N_7038,N_7169);
xnor U7275 (N_7275,N_6340,N_6237);
xor U7276 (N_7276,N_6113,N_6486);
nor U7277 (N_7277,N_6283,N_6971);
nand U7278 (N_7278,N_6845,N_6229);
nand U7279 (N_7279,N_6453,N_6897);
nand U7280 (N_7280,N_6584,N_7181);
nor U7281 (N_7281,N_6569,N_6702);
or U7282 (N_7282,N_6314,N_6432);
nor U7283 (N_7283,N_6967,N_6238);
nor U7284 (N_7284,N_6552,N_7163);
nor U7285 (N_7285,N_6104,N_6547);
nor U7286 (N_7286,N_6396,N_6420);
nand U7287 (N_7287,N_6023,N_6355);
or U7288 (N_7288,N_6811,N_6371);
and U7289 (N_7289,N_6703,N_6998);
xnor U7290 (N_7290,N_6470,N_6352);
nand U7291 (N_7291,N_6819,N_6060);
nand U7292 (N_7292,N_6751,N_6650);
xor U7293 (N_7293,N_7123,N_6399);
or U7294 (N_7294,N_6919,N_6433);
or U7295 (N_7295,N_6884,N_6083);
nand U7296 (N_7296,N_6757,N_6441);
and U7297 (N_7297,N_6094,N_6628);
and U7298 (N_7298,N_6305,N_6715);
and U7299 (N_7299,N_6213,N_6833);
xnor U7300 (N_7300,N_7164,N_6320);
xnor U7301 (N_7301,N_6762,N_7013);
xnor U7302 (N_7302,N_6933,N_6937);
nand U7303 (N_7303,N_6110,N_6592);
or U7304 (N_7304,N_6661,N_6080);
and U7305 (N_7305,N_6463,N_6691);
and U7306 (N_7306,N_6921,N_6288);
or U7307 (N_7307,N_7056,N_6336);
or U7308 (N_7308,N_6990,N_6341);
or U7309 (N_7309,N_6536,N_6274);
and U7310 (N_7310,N_6177,N_7182);
and U7311 (N_7311,N_6088,N_6683);
nand U7312 (N_7312,N_7040,N_7051);
xnor U7313 (N_7313,N_7159,N_6600);
nand U7314 (N_7314,N_6830,N_6862);
nand U7315 (N_7315,N_6849,N_7155);
nor U7316 (N_7316,N_6450,N_6765);
nand U7317 (N_7317,N_6538,N_6973);
xnor U7318 (N_7318,N_6936,N_6682);
xor U7319 (N_7319,N_6595,N_6591);
nor U7320 (N_7320,N_6561,N_6803);
xnor U7321 (N_7321,N_6365,N_6882);
nor U7322 (N_7322,N_6989,N_6402);
nand U7323 (N_7323,N_6554,N_6053);
nand U7324 (N_7324,N_6458,N_6631);
nand U7325 (N_7325,N_7143,N_6145);
nand U7326 (N_7326,N_6315,N_6185);
nor U7327 (N_7327,N_6993,N_6050);
or U7328 (N_7328,N_6026,N_6120);
or U7329 (N_7329,N_6490,N_6768);
xor U7330 (N_7330,N_6639,N_7153);
nand U7331 (N_7331,N_6817,N_6807);
nor U7332 (N_7332,N_6156,N_7070);
xnor U7333 (N_7333,N_6256,N_6642);
and U7334 (N_7334,N_7104,N_6188);
nand U7335 (N_7335,N_6323,N_7102);
xor U7336 (N_7336,N_6027,N_6491);
or U7337 (N_7337,N_6322,N_6798);
nor U7338 (N_7338,N_6211,N_7185);
or U7339 (N_7339,N_6215,N_6766);
xor U7340 (N_7340,N_6730,N_6452);
or U7341 (N_7341,N_6364,N_6370);
or U7342 (N_7342,N_6793,N_6568);
nand U7343 (N_7343,N_6325,N_6302);
nor U7344 (N_7344,N_7110,N_6883);
nand U7345 (N_7345,N_6048,N_6387);
nor U7346 (N_7346,N_6977,N_6281);
xnor U7347 (N_7347,N_6137,N_6666);
or U7348 (N_7348,N_6485,N_6244);
xor U7349 (N_7349,N_6267,N_6017);
nand U7350 (N_7350,N_6307,N_7101);
xnor U7351 (N_7351,N_6056,N_6996);
and U7352 (N_7352,N_6222,N_6423);
nor U7353 (N_7353,N_7179,N_6257);
nand U7354 (N_7354,N_6597,N_6251);
nor U7355 (N_7355,N_6813,N_6799);
xor U7356 (N_7356,N_6559,N_6789);
or U7357 (N_7357,N_7018,N_6943);
nand U7358 (N_7358,N_6952,N_6941);
nor U7359 (N_7359,N_6928,N_6620);
nor U7360 (N_7360,N_6510,N_6680);
nand U7361 (N_7361,N_6195,N_6236);
and U7362 (N_7362,N_7145,N_6451);
or U7363 (N_7363,N_6863,N_6280);
nand U7364 (N_7364,N_7069,N_7111);
and U7365 (N_7365,N_6725,N_6250);
or U7366 (N_7366,N_7008,N_6640);
nor U7367 (N_7367,N_6974,N_6208);
xnor U7368 (N_7368,N_6129,N_6067);
and U7369 (N_7369,N_6696,N_6509);
xnor U7370 (N_7370,N_6095,N_6583);
or U7371 (N_7371,N_6424,N_6525);
and U7372 (N_7372,N_6914,N_6335);
nor U7373 (N_7373,N_6507,N_6034);
and U7374 (N_7374,N_6085,N_7127);
nor U7375 (N_7375,N_6774,N_6277);
nand U7376 (N_7376,N_7087,N_6664);
nand U7377 (N_7377,N_6763,N_6851);
nand U7378 (N_7378,N_6743,N_6988);
nand U7379 (N_7379,N_7037,N_6271);
nand U7380 (N_7380,N_6476,N_6261);
xnor U7381 (N_7381,N_6571,N_7139);
and U7382 (N_7382,N_6701,N_7036);
nand U7383 (N_7383,N_6268,N_6856);
nand U7384 (N_7384,N_6123,N_7117);
nand U7385 (N_7385,N_6376,N_6019);
nor U7386 (N_7386,N_7064,N_6407);
or U7387 (N_7387,N_7107,N_6464);
xnor U7388 (N_7388,N_6825,N_6815);
nand U7389 (N_7389,N_6136,N_6219);
or U7390 (N_7390,N_6869,N_6502);
nand U7391 (N_7391,N_6331,N_6125);
nand U7392 (N_7392,N_6514,N_6111);
or U7393 (N_7393,N_6511,N_6338);
and U7394 (N_7394,N_7126,N_6643);
and U7395 (N_7395,N_6127,N_6930);
and U7396 (N_7396,N_6073,N_6247);
xor U7397 (N_7397,N_7042,N_6090);
and U7398 (N_7398,N_6611,N_6995);
nor U7399 (N_7399,N_6724,N_7016);
nor U7400 (N_7400,N_6068,N_6658);
or U7401 (N_7401,N_6676,N_6632);
xor U7402 (N_7402,N_7055,N_7022);
nand U7403 (N_7403,N_6535,N_6626);
nand U7404 (N_7404,N_6349,N_7108);
and U7405 (N_7405,N_6874,N_7116);
or U7406 (N_7406,N_6116,N_6004);
or U7407 (N_7407,N_6563,N_6677);
and U7408 (N_7408,N_6908,N_6440);
or U7409 (N_7409,N_6594,N_6850);
and U7410 (N_7410,N_6773,N_6994);
and U7411 (N_7411,N_6522,N_6524);
nor U7412 (N_7412,N_6018,N_6567);
and U7413 (N_7413,N_6269,N_6599);
xor U7414 (N_7414,N_6161,N_7019);
nor U7415 (N_7415,N_6714,N_7148);
and U7416 (N_7416,N_6411,N_6985);
or U7417 (N_7417,N_6413,N_6081);
nand U7418 (N_7418,N_6368,N_6044);
nor U7419 (N_7419,N_6965,N_6802);
or U7420 (N_7420,N_6055,N_6881);
or U7421 (N_7421,N_6357,N_6103);
and U7422 (N_7422,N_6729,N_7043);
or U7423 (N_7423,N_6037,N_6152);
and U7424 (N_7424,N_6915,N_6687);
xor U7425 (N_7425,N_6386,N_6200);
and U7426 (N_7426,N_7188,N_6659);
and U7427 (N_7427,N_6596,N_6228);
nor U7428 (N_7428,N_6366,N_6459);
nor U7429 (N_7429,N_6876,N_6076);
nand U7430 (N_7430,N_6570,N_6976);
nand U7431 (N_7431,N_6446,N_6063);
nor U7432 (N_7432,N_6032,N_6647);
nor U7433 (N_7433,N_6875,N_6149);
or U7434 (N_7434,N_6447,N_6266);
nand U7435 (N_7435,N_6414,N_6218);
or U7436 (N_7436,N_6527,N_6254);
nand U7437 (N_7437,N_6400,N_7083);
xnor U7438 (N_7438,N_6521,N_6412);
or U7439 (N_7439,N_6427,N_6285);
and U7440 (N_7440,N_6086,N_6209);
nand U7441 (N_7441,N_6841,N_6645);
or U7442 (N_7442,N_6546,N_6652);
and U7443 (N_7443,N_6769,N_7026);
nor U7444 (N_7444,N_6886,N_6942);
nand U7445 (N_7445,N_6991,N_7002);
xnor U7446 (N_7446,N_7128,N_6679);
nor U7447 (N_7447,N_6795,N_6199);
nand U7448 (N_7448,N_6747,N_7196);
nor U7449 (N_7449,N_6287,N_6684);
and U7450 (N_7450,N_6010,N_6794);
xnor U7451 (N_7451,N_6972,N_6000);
nand U7452 (N_7452,N_6303,N_6772);
nor U7453 (N_7453,N_6621,N_6860);
and U7454 (N_7454,N_6496,N_6779);
or U7455 (N_7455,N_6675,N_7011);
xnor U7456 (N_7456,N_6098,N_7077);
nor U7457 (N_7457,N_6911,N_7052);
and U7458 (N_7458,N_7166,N_6405);
nor U7459 (N_7459,N_6818,N_6742);
nor U7460 (N_7460,N_6668,N_6651);
or U7461 (N_7461,N_6670,N_6240);
and U7462 (N_7462,N_6787,N_6958);
nor U7463 (N_7463,N_6940,N_6043);
nor U7464 (N_7464,N_6221,N_6252);
nor U7465 (N_7465,N_6395,N_6367);
nand U7466 (N_7466,N_6373,N_6859);
and U7467 (N_7467,N_6660,N_6135);
or U7468 (N_7468,N_6609,N_7191);
nor U7469 (N_7469,N_7053,N_6672);
or U7470 (N_7470,N_7158,N_6518);
and U7471 (N_7471,N_6528,N_6159);
nand U7472 (N_7472,N_6806,N_6950);
xnor U7473 (N_7473,N_6727,N_6170);
nand U7474 (N_7474,N_6138,N_6301);
nor U7475 (N_7475,N_6962,N_6025);
or U7476 (N_7476,N_6842,N_7020);
xor U7477 (N_7477,N_6868,N_6853);
and U7478 (N_7478,N_6984,N_6748);
nor U7479 (N_7479,N_6678,N_6981);
or U7480 (N_7480,N_6616,N_6540);
or U7481 (N_7481,N_7081,N_6719);
or U7482 (N_7482,N_6148,N_6316);
nand U7483 (N_7483,N_6122,N_6885);
xnor U7484 (N_7484,N_6009,N_6196);
and U7485 (N_7485,N_6663,N_6045);
nand U7486 (N_7486,N_6786,N_6270);
xnor U7487 (N_7487,N_6054,N_6619);
nand U7488 (N_7488,N_7039,N_6636);
xnor U7489 (N_7489,N_6179,N_6471);
nand U7490 (N_7490,N_6454,N_6646);
or U7491 (N_7491,N_6052,N_6635);
nand U7492 (N_7492,N_6410,N_6362);
nand U7493 (N_7493,N_6311,N_6158);
and U7494 (N_7494,N_6101,N_6733);
nor U7495 (N_7495,N_6877,N_6477);
nand U7496 (N_7496,N_7168,N_6382);
nand U7497 (N_7497,N_6838,N_7195);
nor U7498 (N_7498,N_6694,N_6968);
and U7499 (N_7499,N_6667,N_6982);
nand U7500 (N_7500,N_6770,N_6332);
and U7501 (N_7501,N_6143,N_6771);
and U7502 (N_7502,N_6342,N_6964);
nand U7503 (N_7503,N_6550,N_6530);
nor U7504 (N_7504,N_6214,N_6898);
xor U7505 (N_7505,N_6565,N_6734);
xor U7506 (N_7506,N_6746,N_6258);
and U7507 (N_7507,N_6627,N_6983);
or U7508 (N_7508,N_6172,N_6721);
nand U7509 (N_7509,N_6109,N_6601);
nand U7510 (N_7510,N_6587,N_7098);
and U7511 (N_7511,N_6064,N_6175);
and U7512 (N_7512,N_6681,N_6848);
and U7513 (N_7513,N_6566,N_6904);
nor U7514 (N_7514,N_6629,N_6126);
and U7515 (N_7515,N_6624,N_6397);
nor U7516 (N_7516,N_6654,N_6230);
nor U7517 (N_7517,N_6061,N_6865);
nor U7518 (N_7518,N_7093,N_6955);
or U7519 (N_7519,N_6893,N_6997);
xnor U7520 (N_7520,N_7017,N_6589);
or U7521 (N_7521,N_6558,N_7046);
or U7522 (N_7522,N_6245,N_6516);
nor U7523 (N_7523,N_6674,N_6226);
nor U7524 (N_7524,N_6478,N_6615);
and U7525 (N_7525,N_7106,N_6726);
xnor U7526 (N_7526,N_6935,N_7065);
nand U7527 (N_7527,N_6106,N_6761);
and U7528 (N_7528,N_6429,N_6070);
nor U7529 (N_7529,N_6598,N_6688);
xor U7530 (N_7530,N_6141,N_6231);
xnor U7531 (N_7531,N_6623,N_6383);
or U7532 (N_7532,N_6630,N_6253);
or U7533 (N_7533,N_6622,N_6449);
nand U7534 (N_7534,N_7041,N_6002);
nor U7535 (N_7535,N_7135,N_7192);
nor U7536 (N_7536,N_6404,N_6932);
nor U7537 (N_7537,N_6005,N_6954);
nor U7538 (N_7538,N_6291,N_6326);
xnor U7539 (N_7539,N_6916,N_6276);
or U7540 (N_7540,N_6889,N_6191);
xor U7541 (N_7541,N_6899,N_6831);
nor U7542 (N_7542,N_6262,N_6071);
and U7543 (N_7543,N_6969,N_6957);
and U7544 (N_7544,N_7027,N_6197);
nand U7545 (N_7545,N_6472,N_7177);
and U7546 (N_7546,N_6242,N_7047);
or U7547 (N_7547,N_6906,N_6168);
nor U7548 (N_7548,N_6448,N_6381);
and U7549 (N_7549,N_6379,N_6858);
and U7550 (N_7550,N_6369,N_6560);
xnor U7551 (N_7551,N_6298,N_7068);
nor U7552 (N_7552,N_6970,N_7067);
nand U7553 (N_7553,N_6909,N_6474);
nand U7554 (N_7554,N_6750,N_6712);
nand U7555 (N_7555,N_7174,N_6685);
xnor U7556 (N_7556,N_6887,N_6473);
nor U7557 (N_7557,N_6506,N_6093);
xor U7558 (N_7558,N_7035,N_6775);
xnor U7559 (N_7559,N_6541,N_6212);
nor U7560 (N_7560,N_6764,N_6931);
and U7561 (N_7561,N_7060,N_6492);
and U7562 (N_7562,N_6844,N_6839);
xnor U7563 (N_7563,N_7122,N_6812);
and U7564 (N_7564,N_6278,N_6832);
nand U7565 (N_7565,N_6895,N_6099);
or U7566 (N_7566,N_6574,N_6480);
xor U7567 (N_7567,N_7085,N_6279);
nor U7568 (N_7568,N_6422,N_6992);
xor U7569 (N_7569,N_6030,N_6011);
nor U7570 (N_7570,N_6926,N_6959);
nand U7571 (N_7571,N_6543,N_6007);
and U7572 (N_7572,N_6013,N_6084);
and U7573 (N_7573,N_6662,N_7021);
xnor U7574 (N_7574,N_6837,N_6198);
xor U7575 (N_7575,N_6755,N_6193);
or U7576 (N_7576,N_7152,N_6436);
or U7577 (N_7577,N_6108,N_7028);
nor U7578 (N_7578,N_6501,N_6358);
nor U7579 (N_7579,N_6948,N_6718);
xor U7580 (N_7580,N_6944,N_6872);
and U7581 (N_7581,N_7045,N_7198);
xnor U7582 (N_7582,N_6042,N_6612);
xor U7583 (N_7583,N_6533,N_6716);
nor U7584 (N_7584,N_6406,N_6206);
nor U7585 (N_7585,N_6393,N_6345);
nor U7586 (N_7586,N_6752,N_6022);
and U7587 (N_7587,N_7109,N_6713);
xnor U7588 (N_7588,N_7078,N_7009);
nand U7589 (N_7589,N_6929,N_7136);
xor U7590 (N_7590,N_7154,N_6846);
nand U7591 (N_7591,N_6334,N_7025);
nor U7592 (N_7592,N_6100,N_6390);
nor U7593 (N_7593,N_7133,N_7079);
nor U7594 (N_7594,N_6901,N_6739);
nand U7595 (N_7595,N_6754,N_6804);
xor U7596 (N_7596,N_6949,N_6537);
nand U7597 (N_7597,N_6163,N_6590);
nand U7598 (N_7598,N_6297,N_7063);
nor U7599 (N_7599,N_6319,N_6167);
or U7600 (N_7600,N_6657,N_6890);
xor U7601 (N_7601,N_6121,N_6731);
or U7602 (N_7602,N_6564,N_6649);
nor U7603 (N_7603,N_6210,N_7006);
xnor U7604 (N_7604,N_6756,N_6834);
and U7605 (N_7605,N_6435,N_6192);
or U7606 (N_7606,N_6749,N_6324);
nor U7607 (N_7607,N_6913,N_6634);
or U7608 (N_7608,N_6482,N_6788);
or U7609 (N_7609,N_7170,N_6920);
xor U7610 (N_7610,N_6892,N_6781);
nor U7611 (N_7611,N_6508,N_6465);
xnor U7612 (N_7612,N_6128,N_6783);
xor U7613 (N_7613,N_6264,N_6360);
and U7614 (N_7614,N_6625,N_7197);
nor U7615 (N_7615,N_7183,N_7033);
nand U7616 (N_7616,N_6728,N_6495);
xnor U7617 (N_7617,N_6759,N_6227);
nor U7618 (N_7618,N_7184,N_6239);
and U7619 (N_7619,N_6740,N_6489);
nor U7620 (N_7620,N_6343,N_6089);
nor U7621 (N_7621,N_6014,N_6956);
nand U7622 (N_7622,N_6717,N_6855);
nand U7623 (N_7623,N_6327,N_6827);
xor U7624 (N_7624,N_6284,N_6777);
and U7625 (N_7625,N_6689,N_6201);
nand U7626 (N_7626,N_6417,N_7141);
or U7627 (N_7627,N_7054,N_6031);
nor U7628 (N_7628,N_6401,N_6246);
and U7629 (N_7629,N_6437,N_6581);
and U7630 (N_7630,N_6207,N_6114);
xnor U7631 (N_7631,N_7125,N_6419);
or U7632 (N_7632,N_6461,N_7140);
and U7633 (N_7633,N_7115,N_6902);
nand U7634 (N_7634,N_6843,N_6608);
xnor U7635 (N_7635,N_7030,N_7171);
nor U7636 (N_7636,N_6194,N_6980);
or U7637 (N_7637,N_6035,N_6176);
nand U7638 (N_7638,N_6534,N_6745);
nand U7639 (N_7639,N_6880,N_6945);
xnor U7640 (N_7640,N_7144,N_6481);
nand U7641 (N_7641,N_6455,N_6385);
xnor U7642 (N_7642,N_6062,N_6263);
nand U7643 (N_7643,N_7029,N_7001);
and U7644 (N_7644,N_6015,N_6493);
xnor U7645 (N_7645,N_6337,N_6181);
or U7646 (N_7646,N_6487,N_6999);
or U7647 (N_7647,N_7118,N_7088);
nand U7648 (N_7648,N_6075,N_7012);
xor U7649 (N_7649,N_6102,N_7151);
and U7650 (N_7650,N_6310,N_6544);
and U7651 (N_7651,N_7096,N_6131);
nand U7652 (N_7652,N_7000,N_7076);
xnor U7653 (N_7653,N_7193,N_6697);
xor U7654 (N_7654,N_7146,N_6852);
or U7655 (N_7655,N_6542,N_6582);
nand U7656 (N_7656,N_6722,N_6700);
nand U7657 (N_7657,N_6409,N_6225);
and U7658 (N_7658,N_6479,N_6720);
xnor U7659 (N_7659,N_6699,N_6545);
nor U7660 (N_7660,N_6648,N_6939);
and U7661 (N_7661,N_7132,N_6006);
nor U7662 (N_7662,N_6669,N_6444);
and U7663 (N_7663,N_6290,N_7097);
and U7664 (N_7664,N_6814,N_6391);
or U7665 (N_7665,N_7080,N_6434);
xor U7666 (N_7666,N_6082,N_6421);
or U7667 (N_7667,N_6204,N_6607);
xor U7668 (N_7668,N_7003,N_6289);
xor U7669 (N_7669,N_6220,N_6785);
xnor U7670 (N_7670,N_6695,N_6828);
and U7671 (N_7671,N_6821,N_6403);
nor U7672 (N_7672,N_6801,N_6046);
or U7673 (N_7673,N_6555,N_6072);
nor U7674 (N_7674,N_7073,N_6124);
xnor U7675 (N_7675,N_6979,N_6260);
xor U7676 (N_7676,N_6760,N_6029);
or U7677 (N_7677,N_6351,N_6415);
or U7678 (N_7678,N_6653,N_6693);
and U7679 (N_7679,N_6498,N_6008);
nor U7680 (N_7680,N_6259,N_6174);
or U7681 (N_7681,N_6467,N_7014);
and U7682 (N_7682,N_6065,N_6462);
xnor U7683 (N_7683,N_6585,N_6216);
nor U7684 (N_7684,N_6905,N_6087);
nor U7685 (N_7685,N_6796,N_6791);
nor U7686 (N_7686,N_6790,N_6705);
or U7687 (N_7687,N_6497,N_6784);
and U7688 (N_7688,N_6665,N_6233);
nor U7689 (N_7689,N_6378,N_6171);
or U7690 (N_7690,N_6557,N_6249);
nand U7691 (N_7691,N_6438,N_6292);
nand U7692 (N_7692,N_6205,N_6057);
xor U7693 (N_7693,N_7049,N_6466);
nor U7694 (N_7694,N_6313,N_6265);
and U7695 (N_7695,N_7061,N_6878);
or U7696 (N_7696,N_6096,N_6097);
nor U7697 (N_7697,N_6822,N_6707);
and U7698 (N_7698,N_6308,N_6118);
nor U7699 (N_7699,N_6711,N_6041);
xnor U7700 (N_7700,N_6840,N_6580);
or U7701 (N_7701,N_6656,N_6293);
nor U7702 (N_7702,N_6140,N_6183);
xnor U7703 (N_7703,N_6312,N_6182);
and U7704 (N_7704,N_6112,N_6797);
or U7705 (N_7705,N_6778,N_7119);
and U7706 (N_7706,N_7090,N_6329);
or U7707 (N_7707,N_6576,N_6823);
xor U7708 (N_7708,N_6736,N_6468);
nor U7709 (N_7709,N_7114,N_7134);
xnor U7710 (N_7710,N_6457,N_7048);
xor U7711 (N_7711,N_6776,N_7050);
xnor U7712 (N_7712,N_6456,N_6077);
and U7713 (N_7713,N_6353,N_6987);
and U7714 (N_7714,N_6020,N_6069);
xnor U7715 (N_7715,N_7190,N_6049);
or U7716 (N_7716,N_6139,N_6520);
or U7717 (N_7717,N_6300,N_6356);
xnor U7718 (N_7718,N_6016,N_6512);
or U7719 (N_7719,N_6157,N_6165);
or U7720 (N_7720,N_6418,N_6782);
xnor U7721 (N_7721,N_6001,N_7057);
nand U7722 (N_7722,N_7082,N_6870);
nand U7723 (N_7723,N_6835,N_6153);
nand U7724 (N_7724,N_6575,N_6690);
nor U7725 (N_7725,N_7024,N_6917);
or U7726 (N_7726,N_6963,N_6299);
nand U7727 (N_7727,N_6443,N_6503);
nand U7728 (N_7728,N_6894,N_7071);
xor U7729 (N_7729,N_6255,N_6526);
and U7730 (N_7730,N_6350,N_6494);
nand U7731 (N_7731,N_6741,N_6272);
nand U7732 (N_7732,N_6610,N_7031);
or U7733 (N_7733,N_7150,N_6040);
or U7734 (N_7734,N_6602,N_6363);
nand U7735 (N_7735,N_6549,N_6074);
and U7736 (N_7736,N_6692,N_6033);
xnor U7737 (N_7737,N_7099,N_7059);
nand U7738 (N_7738,N_7180,N_6978);
or U7739 (N_7739,N_6866,N_7100);
xor U7740 (N_7740,N_6224,N_6132);
nand U7741 (N_7741,N_6330,N_7129);
and U7742 (N_7742,N_7137,N_7167);
nor U7743 (N_7743,N_6142,N_7121);
nor U7744 (N_7744,N_6036,N_6709);
or U7745 (N_7745,N_6162,N_6223);
nor U7746 (N_7746,N_7194,N_6294);
and U7747 (N_7747,N_6655,N_6348);
nor U7748 (N_7748,N_7094,N_6504);
nand U7749 (N_7749,N_6130,N_6809);
nor U7750 (N_7750,N_6975,N_6864);
and U7751 (N_7751,N_6924,N_6160);
xnor U7752 (N_7752,N_7162,N_6573);
nor U7753 (N_7753,N_7075,N_6059);
and U7754 (N_7754,N_6673,N_6384);
and U7755 (N_7755,N_6708,N_6562);
nand U7756 (N_7756,N_7157,N_6513);
or U7757 (N_7757,N_6234,N_7161);
and U7758 (N_7758,N_6816,N_6633);
nand U7759 (N_7759,N_6296,N_7091);
nor U7760 (N_7760,N_7173,N_6505);
nand U7761 (N_7761,N_6232,N_6439);
or U7762 (N_7762,N_6469,N_6173);
and U7763 (N_7763,N_6344,N_7138);
or U7764 (N_7764,N_6577,N_6321);
nor U7765 (N_7765,N_6361,N_6744);
nand U7766 (N_7766,N_7120,N_6572);
nand U7767 (N_7767,N_6047,N_6925);
nand U7768 (N_7768,N_7089,N_6767);
or U7769 (N_7769,N_7092,N_6339);
xnor U7770 (N_7770,N_6309,N_6824);
and U7771 (N_7771,N_6500,N_6704);
xor U7772 (N_7772,N_6551,N_6644);
and U7773 (N_7773,N_6922,N_6475);
nand U7774 (N_7774,N_6354,N_6428);
and U7775 (N_7775,N_6529,N_7072);
nor U7776 (N_7776,N_7095,N_6333);
nor U7777 (N_7777,N_6317,N_6134);
nor U7778 (N_7778,N_6374,N_6960);
or U7779 (N_7779,N_7004,N_6388);
nand U7780 (N_7780,N_6180,N_7176);
and U7781 (N_7781,N_6829,N_7172);
nor U7782 (N_7782,N_7062,N_6117);
or U7783 (N_7783,N_7156,N_6539);
xnor U7784 (N_7784,N_6857,N_6820);
xor U7785 (N_7785,N_6430,N_7032);
nand U7786 (N_7786,N_6523,N_6867);
nor U7787 (N_7787,N_6951,N_6637);
nor U7788 (N_7788,N_6416,N_7007);
and U7789 (N_7789,N_6021,N_6946);
xor U7790 (N_7790,N_7103,N_6918);
xnor U7791 (N_7791,N_6698,N_6593);
or U7792 (N_7792,N_6442,N_6217);
nand U7793 (N_7793,N_6389,N_6826);
or U7794 (N_7794,N_6671,N_6202);
nand U7795 (N_7795,N_6306,N_6738);
and U7796 (N_7796,N_6847,N_6613);
nor U7797 (N_7797,N_6425,N_7023);
nand U7798 (N_7798,N_6792,N_6641);
xnor U7799 (N_7799,N_6203,N_6588);
nor U7800 (N_7800,N_6464,N_6521);
nand U7801 (N_7801,N_6423,N_6001);
and U7802 (N_7802,N_7009,N_6255);
nor U7803 (N_7803,N_6216,N_7094);
and U7804 (N_7804,N_7159,N_6519);
nor U7805 (N_7805,N_7117,N_6645);
nor U7806 (N_7806,N_6517,N_6628);
xnor U7807 (N_7807,N_6911,N_6309);
nand U7808 (N_7808,N_7084,N_7071);
nor U7809 (N_7809,N_6121,N_6650);
or U7810 (N_7810,N_6642,N_6471);
or U7811 (N_7811,N_6148,N_6928);
nand U7812 (N_7812,N_6535,N_6016);
nor U7813 (N_7813,N_6733,N_6605);
xnor U7814 (N_7814,N_6150,N_6128);
nor U7815 (N_7815,N_6791,N_7153);
nand U7816 (N_7816,N_6563,N_6517);
nor U7817 (N_7817,N_6429,N_7050);
xor U7818 (N_7818,N_6973,N_6754);
and U7819 (N_7819,N_6115,N_6946);
nor U7820 (N_7820,N_7013,N_6429);
xnor U7821 (N_7821,N_6919,N_6904);
xnor U7822 (N_7822,N_6760,N_6405);
or U7823 (N_7823,N_6694,N_6255);
or U7824 (N_7824,N_6457,N_6543);
xnor U7825 (N_7825,N_6969,N_6139);
nor U7826 (N_7826,N_6732,N_6919);
and U7827 (N_7827,N_6341,N_6856);
xnor U7828 (N_7828,N_6689,N_6648);
nand U7829 (N_7829,N_6077,N_6372);
nor U7830 (N_7830,N_7028,N_6738);
and U7831 (N_7831,N_7141,N_6175);
or U7832 (N_7832,N_6003,N_6837);
or U7833 (N_7833,N_6693,N_6115);
and U7834 (N_7834,N_6282,N_6358);
or U7835 (N_7835,N_6416,N_6145);
nor U7836 (N_7836,N_6709,N_6747);
nor U7837 (N_7837,N_6770,N_6773);
xnor U7838 (N_7838,N_6221,N_6053);
nor U7839 (N_7839,N_6731,N_6565);
nor U7840 (N_7840,N_6691,N_6668);
xnor U7841 (N_7841,N_6495,N_6327);
nor U7842 (N_7842,N_6173,N_6360);
nand U7843 (N_7843,N_6135,N_7184);
and U7844 (N_7844,N_6715,N_6994);
nand U7845 (N_7845,N_6884,N_6380);
nand U7846 (N_7846,N_6277,N_6799);
nand U7847 (N_7847,N_6219,N_6144);
xor U7848 (N_7848,N_6059,N_6050);
nand U7849 (N_7849,N_7163,N_6067);
and U7850 (N_7850,N_7072,N_6997);
and U7851 (N_7851,N_6051,N_6433);
and U7852 (N_7852,N_6828,N_6722);
and U7853 (N_7853,N_6923,N_7178);
and U7854 (N_7854,N_6147,N_6157);
or U7855 (N_7855,N_6181,N_7060);
and U7856 (N_7856,N_6238,N_6787);
xor U7857 (N_7857,N_6044,N_6565);
and U7858 (N_7858,N_7194,N_6206);
nand U7859 (N_7859,N_6066,N_6045);
and U7860 (N_7860,N_6542,N_7139);
and U7861 (N_7861,N_6615,N_6257);
nor U7862 (N_7862,N_6472,N_6100);
and U7863 (N_7863,N_6093,N_6025);
xor U7864 (N_7864,N_7143,N_6233);
nand U7865 (N_7865,N_6533,N_6001);
nor U7866 (N_7866,N_6887,N_6336);
and U7867 (N_7867,N_6679,N_6664);
nor U7868 (N_7868,N_6940,N_6559);
xor U7869 (N_7869,N_6029,N_6971);
nand U7870 (N_7870,N_6019,N_6902);
nand U7871 (N_7871,N_6323,N_7075);
nor U7872 (N_7872,N_7086,N_6495);
or U7873 (N_7873,N_6046,N_6968);
nand U7874 (N_7874,N_6580,N_6690);
and U7875 (N_7875,N_6207,N_6563);
nor U7876 (N_7876,N_6322,N_6374);
xor U7877 (N_7877,N_6208,N_6395);
and U7878 (N_7878,N_6419,N_6212);
nand U7879 (N_7879,N_6427,N_7058);
nand U7880 (N_7880,N_6726,N_7031);
nor U7881 (N_7881,N_7116,N_6226);
and U7882 (N_7882,N_6851,N_6391);
or U7883 (N_7883,N_6493,N_6654);
nand U7884 (N_7884,N_6901,N_6462);
and U7885 (N_7885,N_6966,N_6299);
xnor U7886 (N_7886,N_6946,N_6224);
nor U7887 (N_7887,N_6933,N_6593);
nand U7888 (N_7888,N_6924,N_6134);
or U7889 (N_7889,N_6741,N_6784);
and U7890 (N_7890,N_6898,N_6729);
and U7891 (N_7891,N_6168,N_7131);
nor U7892 (N_7892,N_6745,N_6433);
and U7893 (N_7893,N_6453,N_6998);
and U7894 (N_7894,N_6999,N_6982);
xnor U7895 (N_7895,N_6034,N_6178);
nand U7896 (N_7896,N_6817,N_6355);
or U7897 (N_7897,N_6148,N_6196);
or U7898 (N_7898,N_6831,N_6957);
nor U7899 (N_7899,N_6520,N_7017);
xor U7900 (N_7900,N_6962,N_6374);
or U7901 (N_7901,N_6034,N_6156);
and U7902 (N_7902,N_6802,N_6420);
or U7903 (N_7903,N_7033,N_7124);
nand U7904 (N_7904,N_6768,N_6524);
xor U7905 (N_7905,N_6772,N_6853);
and U7906 (N_7906,N_6039,N_6219);
nand U7907 (N_7907,N_6949,N_6026);
or U7908 (N_7908,N_6450,N_6126);
or U7909 (N_7909,N_6302,N_6406);
and U7910 (N_7910,N_6479,N_6323);
nor U7911 (N_7911,N_6461,N_6675);
xor U7912 (N_7912,N_6174,N_6126);
and U7913 (N_7913,N_6923,N_6832);
nor U7914 (N_7914,N_6610,N_6328);
nor U7915 (N_7915,N_6188,N_7045);
xnor U7916 (N_7916,N_6878,N_6252);
nand U7917 (N_7917,N_7148,N_6626);
nor U7918 (N_7918,N_6709,N_6612);
xor U7919 (N_7919,N_7141,N_6675);
xnor U7920 (N_7920,N_6984,N_6598);
nand U7921 (N_7921,N_7130,N_6339);
nand U7922 (N_7922,N_6194,N_7049);
and U7923 (N_7923,N_6460,N_7183);
nor U7924 (N_7924,N_6636,N_6194);
and U7925 (N_7925,N_6134,N_6497);
nand U7926 (N_7926,N_7183,N_6885);
and U7927 (N_7927,N_6374,N_6815);
nor U7928 (N_7928,N_6562,N_6283);
nor U7929 (N_7929,N_7116,N_7155);
xnor U7930 (N_7930,N_6247,N_6610);
nand U7931 (N_7931,N_6999,N_6583);
and U7932 (N_7932,N_7088,N_6063);
xor U7933 (N_7933,N_6960,N_6514);
nor U7934 (N_7934,N_6440,N_6458);
and U7935 (N_7935,N_6549,N_7161);
nand U7936 (N_7936,N_6634,N_7133);
and U7937 (N_7937,N_6355,N_6204);
nor U7938 (N_7938,N_6264,N_6004);
and U7939 (N_7939,N_7180,N_7140);
nand U7940 (N_7940,N_7132,N_7037);
nor U7941 (N_7941,N_7004,N_7133);
xor U7942 (N_7942,N_6731,N_7180);
or U7943 (N_7943,N_6246,N_6639);
and U7944 (N_7944,N_6008,N_6525);
nand U7945 (N_7945,N_6972,N_6234);
and U7946 (N_7946,N_6487,N_6527);
nand U7947 (N_7947,N_6284,N_6694);
or U7948 (N_7948,N_6375,N_7032);
nor U7949 (N_7949,N_6653,N_6332);
nor U7950 (N_7950,N_6516,N_6199);
nand U7951 (N_7951,N_6154,N_6655);
and U7952 (N_7952,N_6092,N_7015);
nor U7953 (N_7953,N_7002,N_7176);
nand U7954 (N_7954,N_7110,N_6614);
nor U7955 (N_7955,N_6339,N_6083);
or U7956 (N_7956,N_6614,N_6572);
xor U7957 (N_7957,N_6123,N_6959);
nand U7958 (N_7958,N_6522,N_6378);
nor U7959 (N_7959,N_6264,N_6152);
nor U7960 (N_7960,N_7100,N_7103);
and U7961 (N_7961,N_6881,N_7059);
nor U7962 (N_7962,N_6341,N_6027);
nand U7963 (N_7963,N_6396,N_6833);
xnor U7964 (N_7964,N_6705,N_7130);
and U7965 (N_7965,N_6873,N_6781);
xnor U7966 (N_7966,N_6807,N_7184);
or U7967 (N_7967,N_7148,N_6206);
xnor U7968 (N_7968,N_6617,N_7157);
and U7969 (N_7969,N_6222,N_6598);
nand U7970 (N_7970,N_6491,N_6771);
nor U7971 (N_7971,N_6272,N_7026);
or U7972 (N_7972,N_6929,N_6253);
and U7973 (N_7973,N_6006,N_6119);
xor U7974 (N_7974,N_6196,N_6024);
nor U7975 (N_7975,N_6732,N_7119);
or U7976 (N_7976,N_6022,N_6664);
and U7977 (N_7977,N_6542,N_6981);
or U7978 (N_7978,N_6512,N_6391);
and U7979 (N_7979,N_6101,N_6611);
nor U7980 (N_7980,N_6739,N_6314);
or U7981 (N_7981,N_7021,N_7173);
nand U7982 (N_7982,N_6993,N_6815);
or U7983 (N_7983,N_6353,N_6288);
nand U7984 (N_7984,N_6527,N_6181);
xnor U7985 (N_7985,N_6313,N_6472);
xor U7986 (N_7986,N_7174,N_6699);
nand U7987 (N_7987,N_6441,N_6533);
and U7988 (N_7988,N_6072,N_6721);
nand U7989 (N_7989,N_7018,N_7019);
xor U7990 (N_7990,N_6711,N_7173);
nand U7991 (N_7991,N_6661,N_6307);
xor U7992 (N_7992,N_7098,N_7034);
or U7993 (N_7993,N_6077,N_6451);
xor U7994 (N_7994,N_6938,N_6563);
nand U7995 (N_7995,N_7030,N_6370);
and U7996 (N_7996,N_6289,N_6608);
or U7997 (N_7997,N_6836,N_6723);
xor U7998 (N_7998,N_7119,N_6746);
and U7999 (N_7999,N_6799,N_6814);
xor U8000 (N_8000,N_6873,N_7153);
and U8001 (N_8001,N_6675,N_6190);
nor U8002 (N_8002,N_6260,N_7016);
xnor U8003 (N_8003,N_6959,N_6103);
or U8004 (N_8004,N_6909,N_7156);
xnor U8005 (N_8005,N_6587,N_6950);
xnor U8006 (N_8006,N_6992,N_7099);
xor U8007 (N_8007,N_6142,N_6746);
xor U8008 (N_8008,N_6360,N_6866);
nor U8009 (N_8009,N_6617,N_6795);
and U8010 (N_8010,N_6342,N_6055);
and U8011 (N_8011,N_6804,N_6759);
xor U8012 (N_8012,N_7142,N_6637);
nand U8013 (N_8013,N_6599,N_7007);
xnor U8014 (N_8014,N_6887,N_6616);
xnor U8015 (N_8015,N_6453,N_6107);
nand U8016 (N_8016,N_6366,N_6535);
nor U8017 (N_8017,N_6076,N_6580);
and U8018 (N_8018,N_7076,N_6723);
xor U8019 (N_8019,N_6588,N_6002);
nor U8020 (N_8020,N_6537,N_6785);
or U8021 (N_8021,N_6128,N_6545);
nor U8022 (N_8022,N_7163,N_7021);
nor U8023 (N_8023,N_6635,N_6696);
nand U8024 (N_8024,N_7129,N_6643);
nor U8025 (N_8025,N_6386,N_6141);
or U8026 (N_8026,N_7155,N_7188);
or U8027 (N_8027,N_7115,N_6016);
or U8028 (N_8028,N_6276,N_6977);
or U8029 (N_8029,N_6831,N_6971);
nand U8030 (N_8030,N_7008,N_6107);
xor U8031 (N_8031,N_6332,N_6615);
nand U8032 (N_8032,N_6295,N_6140);
and U8033 (N_8033,N_7085,N_6687);
and U8034 (N_8034,N_6257,N_6105);
nor U8035 (N_8035,N_6754,N_6246);
nor U8036 (N_8036,N_7057,N_6719);
nor U8037 (N_8037,N_6682,N_6872);
and U8038 (N_8038,N_6818,N_6848);
xor U8039 (N_8039,N_6383,N_6960);
and U8040 (N_8040,N_6532,N_6992);
or U8041 (N_8041,N_6764,N_6490);
and U8042 (N_8042,N_6246,N_6555);
nor U8043 (N_8043,N_6398,N_6958);
xor U8044 (N_8044,N_6141,N_6145);
and U8045 (N_8045,N_6212,N_6977);
or U8046 (N_8046,N_6935,N_7062);
xor U8047 (N_8047,N_7120,N_7039);
xor U8048 (N_8048,N_7006,N_6922);
nor U8049 (N_8049,N_6755,N_6086);
and U8050 (N_8050,N_6470,N_7175);
xor U8051 (N_8051,N_6280,N_6552);
nand U8052 (N_8052,N_6119,N_6162);
or U8053 (N_8053,N_6934,N_6924);
nand U8054 (N_8054,N_6568,N_6868);
and U8055 (N_8055,N_7129,N_6115);
nand U8056 (N_8056,N_7083,N_6492);
and U8057 (N_8057,N_6569,N_6475);
and U8058 (N_8058,N_6787,N_6028);
and U8059 (N_8059,N_6580,N_7008);
and U8060 (N_8060,N_6994,N_6875);
nor U8061 (N_8061,N_6353,N_6180);
xor U8062 (N_8062,N_6724,N_6063);
or U8063 (N_8063,N_6577,N_6990);
or U8064 (N_8064,N_6557,N_6681);
or U8065 (N_8065,N_6282,N_6590);
nor U8066 (N_8066,N_6185,N_6223);
or U8067 (N_8067,N_6147,N_6001);
nor U8068 (N_8068,N_6257,N_6292);
xnor U8069 (N_8069,N_6603,N_7015);
nor U8070 (N_8070,N_6157,N_6438);
nand U8071 (N_8071,N_6654,N_6553);
and U8072 (N_8072,N_6784,N_6933);
nand U8073 (N_8073,N_6597,N_6724);
xor U8074 (N_8074,N_6595,N_6437);
nor U8075 (N_8075,N_6505,N_7027);
nand U8076 (N_8076,N_6426,N_6257);
xnor U8077 (N_8077,N_6693,N_6760);
nand U8078 (N_8078,N_6301,N_6081);
nand U8079 (N_8079,N_6878,N_6008);
and U8080 (N_8080,N_6011,N_6878);
or U8081 (N_8081,N_6310,N_6128);
or U8082 (N_8082,N_6625,N_6604);
or U8083 (N_8083,N_7176,N_6617);
xnor U8084 (N_8084,N_6989,N_6374);
nor U8085 (N_8085,N_6128,N_6509);
nand U8086 (N_8086,N_6344,N_6078);
nand U8087 (N_8087,N_6999,N_6091);
xor U8088 (N_8088,N_6928,N_7045);
or U8089 (N_8089,N_6880,N_6732);
nor U8090 (N_8090,N_6428,N_6331);
nor U8091 (N_8091,N_7179,N_6354);
xor U8092 (N_8092,N_6046,N_6581);
and U8093 (N_8093,N_6156,N_6681);
nor U8094 (N_8094,N_6981,N_6633);
nand U8095 (N_8095,N_7082,N_6163);
nand U8096 (N_8096,N_6740,N_6842);
nand U8097 (N_8097,N_7060,N_6184);
and U8098 (N_8098,N_7128,N_6557);
and U8099 (N_8099,N_6017,N_6373);
nand U8100 (N_8100,N_6488,N_7019);
xnor U8101 (N_8101,N_6406,N_6017);
or U8102 (N_8102,N_6864,N_6131);
nor U8103 (N_8103,N_6671,N_7130);
or U8104 (N_8104,N_6346,N_7134);
xor U8105 (N_8105,N_6387,N_6240);
or U8106 (N_8106,N_7157,N_6688);
nand U8107 (N_8107,N_7195,N_6234);
xor U8108 (N_8108,N_6083,N_6697);
or U8109 (N_8109,N_6264,N_6172);
nand U8110 (N_8110,N_7020,N_6196);
and U8111 (N_8111,N_6815,N_7038);
nor U8112 (N_8112,N_6530,N_6130);
nand U8113 (N_8113,N_6100,N_6414);
nor U8114 (N_8114,N_7095,N_6523);
or U8115 (N_8115,N_6539,N_6629);
nor U8116 (N_8116,N_6546,N_6246);
xor U8117 (N_8117,N_6303,N_7069);
or U8118 (N_8118,N_7173,N_6543);
and U8119 (N_8119,N_6842,N_7123);
and U8120 (N_8120,N_6252,N_6808);
or U8121 (N_8121,N_6100,N_6021);
nand U8122 (N_8122,N_6600,N_6590);
nor U8123 (N_8123,N_6295,N_7032);
or U8124 (N_8124,N_6434,N_6137);
or U8125 (N_8125,N_6857,N_6258);
nor U8126 (N_8126,N_6293,N_6171);
and U8127 (N_8127,N_6313,N_6744);
or U8128 (N_8128,N_6620,N_7051);
and U8129 (N_8129,N_6015,N_7101);
nor U8130 (N_8130,N_6592,N_7166);
nor U8131 (N_8131,N_6492,N_7066);
or U8132 (N_8132,N_6317,N_6138);
nor U8133 (N_8133,N_6307,N_6314);
nor U8134 (N_8134,N_6937,N_6335);
and U8135 (N_8135,N_6196,N_6039);
and U8136 (N_8136,N_6656,N_6010);
and U8137 (N_8137,N_6475,N_7084);
and U8138 (N_8138,N_6416,N_6975);
and U8139 (N_8139,N_6120,N_6331);
and U8140 (N_8140,N_6566,N_6898);
nor U8141 (N_8141,N_6931,N_7055);
nand U8142 (N_8142,N_6017,N_6558);
nand U8143 (N_8143,N_6440,N_7117);
nand U8144 (N_8144,N_7162,N_6277);
and U8145 (N_8145,N_6002,N_6756);
xnor U8146 (N_8146,N_7040,N_6823);
nand U8147 (N_8147,N_7106,N_6101);
nor U8148 (N_8148,N_6886,N_6227);
xnor U8149 (N_8149,N_6705,N_6853);
and U8150 (N_8150,N_7139,N_6187);
nor U8151 (N_8151,N_6688,N_6158);
nand U8152 (N_8152,N_6621,N_6922);
or U8153 (N_8153,N_7072,N_6544);
or U8154 (N_8154,N_6340,N_6335);
xor U8155 (N_8155,N_6546,N_6824);
and U8156 (N_8156,N_6280,N_6617);
xor U8157 (N_8157,N_6530,N_6201);
xor U8158 (N_8158,N_6530,N_6054);
xnor U8159 (N_8159,N_6716,N_6375);
nor U8160 (N_8160,N_6085,N_6225);
or U8161 (N_8161,N_6162,N_6192);
and U8162 (N_8162,N_6162,N_6149);
xnor U8163 (N_8163,N_6383,N_6335);
nand U8164 (N_8164,N_6426,N_6779);
nor U8165 (N_8165,N_6660,N_6126);
and U8166 (N_8166,N_6610,N_6671);
nor U8167 (N_8167,N_6677,N_6122);
xor U8168 (N_8168,N_6810,N_6761);
xnor U8169 (N_8169,N_6039,N_6152);
nand U8170 (N_8170,N_6758,N_6954);
and U8171 (N_8171,N_7071,N_6132);
xor U8172 (N_8172,N_6638,N_6071);
and U8173 (N_8173,N_6220,N_6852);
nor U8174 (N_8174,N_6309,N_7165);
and U8175 (N_8175,N_6329,N_6382);
nand U8176 (N_8176,N_6092,N_6986);
and U8177 (N_8177,N_6370,N_7115);
nand U8178 (N_8178,N_6527,N_6266);
and U8179 (N_8179,N_6398,N_6830);
and U8180 (N_8180,N_6351,N_6681);
or U8181 (N_8181,N_6429,N_6235);
nor U8182 (N_8182,N_6191,N_6060);
and U8183 (N_8183,N_7011,N_7042);
xor U8184 (N_8184,N_6772,N_6495);
or U8185 (N_8185,N_6415,N_6139);
nand U8186 (N_8186,N_6972,N_6454);
nor U8187 (N_8187,N_6970,N_6121);
nor U8188 (N_8188,N_6582,N_6731);
nand U8189 (N_8189,N_7091,N_6914);
nand U8190 (N_8190,N_6851,N_6720);
xnor U8191 (N_8191,N_6133,N_6953);
xnor U8192 (N_8192,N_6376,N_6121);
or U8193 (N_8193,N_6376,N_6176);
nor U8194 (N_8194,N_6730,N_6282);
and U8195 (N_8195,N_7069,N_6052);
nand U8196 (N_8196,N_6440,N_6939);
xnor U8197 (N_8197,N_6164,N_7069);
nor U8198 (N_8198,N_6801,N_6089);
or U8199 (N_8199,N_6321,N_6892);
nor U8200 (N_8200,N_6737,N_6124);
xnor U8201 (N_8201,N_7012,N_6455);
nand U8202 (N_8202,N_6788,N_6497);
xor U8203 (N_8203,N_6117,N_6473);
xnor U8204 (N_8204,N_6373,N_6064);
or U8205 (N_8205,N_6190,N_6237);
xnor U8206 (N_8206,N_6061,N_6300);
or U8207 (N_8207,N_6558,N_6981);
nand U8208 (N_8208,N_6891,N_6678);
or U8209 (N_8209,N_6506,N_6776);
and U8210 (N_8210,N_6423,N_7180);
nor U8211 (N_8211,N_6164,N_6592);
or U8212 (N_8212,N_6044,N_6250);
nor U8213 (N_8213,N_6189,N_6959);
or U8214 (N_8214,N_6869,N_6333);
nor U8215 (N_8215,N_6536,N_6400);
xnor U8216 (N_8216,N_6730,N_6062);
and U8217 (N_8217,N_6185,N_6623);
nor U8218 (N_8218,N_6701,N_6462);
nand U8219 (N_8219,N_7190,N_7111);
nor U8220 (N_8220,N_6497,N_6897);
nor U8221 (N_8221,N_6466,N_6791);
xnor U8222 (N_8222,N_6706,N_6958);
or U8223 (N_8223,N_6268,N_6935);
nand U8224 (N_8224,N_6658,N_6076);
or U8225 (N_8225,N_7138,N_6678);
nand U8226 (N_8226,N_6376,N_6746);
nand U8227 (N_8227,N_7131,N_6988);
nand U8228 (N_8228,N_6177,N_6292);
nor U8229 (N_8229,N_6267,N_6625);
nand U8230 (N_8230,N_6013,N_7056);
and U8231 (N_8231,N_6296,N_6128);
or U8232 (N_8232,N_6114,N_6827);
nand U8233 (N_8233,N_6888,N_6100);
or U8234 (N_8234,N_6061,N_6106);
nor U8235 (N_8235,N_6964,N_7163);
xor U8236 (N_8236,N_7199,N_6282);
or U8237 (N_8237,N_6679,N_7001);
and U8238 (N_8238,N_6509,N_6416);
nor U8239 (N_8239,N_6500,N_6285);
nor U8240 (N_8240,N_6923,N_7087);
nand U8241 (N_8241,N_6027,N_6105);
nor U8242 (N_8242,N_6412,N_6004);
xnor U8243 (N_8243,N_6634,N_6879);
or U8244 (N_8244,N_6022,N_6594);
or U8245 (N_8245,N_6057,N_6054);
and U8246 (N_8246,N_6914,N_6781);
nor U8247 (N_8247,N_6312,N_6876);
or U8248 (N_8248,N_6361,N_6278);
xor U8249 (N_8249,N_6388,N_6584);
or U8250 (N_8250,N_7103,N_6765);
nand U8251 (N_8251,N_6548,N_6906);
nand U8252 (N_8252,N_6694,N_6571);
nor U8253 (N_8253,N_6140,N_6040);
xor U8254 (N_8254,N_6070,N_6286);
xor U8255 (N_8255,N_6681,N_6529);
nand U8256 (N_8256,N_7188,N_6021);
xnor U8257 (N_8257,N_6316,N_6410);
nand U8258 (N_8258,N_6988,N_6422);
or U8259 (N_8259,N_6580,N_6593);
xor U8260 (N_8260,N_6919,N_6171);
nand U8261 (N_8261,N_6392,N_7042);
nor U8262 (N_8262,N_7036,N_7029);
nand U8263 (N_8263,N_6239,N_6946);
and U8264 (N_8264,N_7067,N_6468);
and U8265 (N_8265,N_7061,N_6249);
nand U8266 (N_8266,N_6909,N_6715);
and U8267 (N_8267,N_6424,N_7000);
nand U8268 (N_8268,N_6840,N_6283);
and U8269 (N_8269,N_6118,N_6044);
nand U8270 (N_8270,N_6343,N_6303);
xnor U8271 (N_8271,N_6613,N_6971);
nor U8272 (N_8272,N_6658,N_7006);
nand U8273 (N_8273,N_7109,N_7070);
xor U8274 (N_8274,N_6127,N_6943);
xnor U8275 (N_8275,N_6075,N_6369);
or U8276 (N_8276,N_6588,N_7112);
nor U8277 (N_8277,N_6303,N_6165);
xor U8278 (N_8278,N_6768,N_6462);
or U8279 (N_8279,N_6868,N_6646);
or U8280 (N_8280,N_6937,N_6984);
nor U8281 (N_8281,N_6672,N_6325);
and U8282 (N_8282,N_6248,N_7039);
xnor U8283 (N_8283,N_6179,N_6535);
xor U8284 (N_8284,N_6743,N_7109);
xnor U8285 (N_8285,N_6335,N_6124);
or U8286 (N_8286,N_6872,N_7173);
and U8287 (N_8287,N_6633,N_7008);
and U8288 (N_8288,N_6940,N_6378);
and U8289 (N_8289,N_6691,N_6506);
xor U8290 (N_8290,N_6913,N_6246);
nor U8291 (N_8291,N_6692,N_6070);
xor U8292 (N_8292,N_6696,N_6959);
xor U8293 (N_8293,N_6494,N_6022);
xor U8294 (N_8294,N_6924,N_6920);
xnor U8295 (N_8295,N_6020,N_6790);
nor U8296 (N_8296,N_6986,N_6070);
xnor U8297 (N_8297,N_6134,N_6243);
xnor U8298 (N_8298,N_6095,N_6963);
or U8299 (N_8299,N_6210,N_6839);
nand U8300 (N_8300,N_6702,N_6142);
xor U8301 (N_8301,N_6556,N_6448);
or U8302 (N_8302,N_6155,N_6655);
nor U8303 (N_8303,N_6815,N_6778);
or U8304 (N_8304,N_6506,N_6290);
xnor U8305 (N_8305,N_6084,N_6336);
nor U8306 (N_8306,N_6402,N_7111);
nand U8307 (N_8307,N_6640,N_6605);
xnor U8308 (N_8308,N_6683,N_6940);
xnor U8309 (N_8309,N_6415,N_6548);
nand U8310 (N_8310,N_6204,N_7193);
xor U8311 (N_8311,N_6226,N_7035);
nand U8312 (N_8312,N_6139,N_6375);
nor U8313 (N_8313,N_6797,N_7160);
nand U8314 (N_8314,N_6503,N_6007);
or U8315 (N_8315,N_6915,N_6766);
nor U8316 (N_8316,N_7058,N_6039);
nand U8317 (N_8317,N_6647,N_6519);
nand U8318 (N_8318,N_6375,N_6477);
nand U8319 (N_8319,N_6113,N_7152);
or U8320 (N_8320,N_6965,N_7150);
nor U8321 (N_8321,N_6905,N_6939);
nor U8322 (N_8322,N_6060,N_6220);
or U8323 (N_8323,N_6239,N_6446);
nor U8324 (N_8324,N_6372,N_6987);
nor U8325 (N_8325,N_7000,N_6054);
nor U8326 (N_8326,N_6647,N_6447);
nor U8327 (N_8327,N_6933,N_6643);
xor U8328 (N_8328,N_6258,N_7191);
nand U8329 (N_8329,N_6737,N_6188);
and U8330 (N_8330,N_6408,N_6750);
or U8331 (N_8331,N_6697,N_7106);
nor U8332 (N_8332,N_6901,N_6044);
nor U8333 (N_8333,N_6629,N_6203);
and U8334 (N_8334,N_7163,N_6992);
xnor U8335 (N_8335,N_6558,N_6722);
nand U8336 (N_8336,N_6024,N_6539);
nand U8337 (N_8337,N_6079,N_6030);
nor U8338 (N_8338,N_6285,N_6211);
nor U8339 (N_8339,N_6558,N_6332);
xor U8340 (N_8340,N_6143,N_6609);
and U8341 (N_8341,N_6253,N_6397);
and U8342 (N_8342,N_6128,N_6916);
and U8343 (N_8343,N_6071,N_6785);
xnor U8344 (N_8344,N_7123,N_6668);
nor U8345 (N_8345,N_6263,N_6707);
nand U8346 (N_8346,N_6735,N_6300);
xor U8347 (N_8347,N_7053,N_6626);
xor U8348 (N_8348,N_6404,N_6024);
or U8349 (N_8349,N_6374,N_6424);
xor U8350 (N_8350,N_6260,N_6810);
nor U8351 (N_8351,N_6069,N_6141);
nor U8352 (N_8352,N_6317,N_7153);
nand U8353 (N_8353,N_6236,N_6692);
xor U8354 (N_8354,N_6280,N_6103);
nand U8355 (N_8355,N_6685,N_6065);
and U8356 (N_8356,N_6005,N_6219);
or U8357 (N_8357,N_7192,N_6970);
nand U8358 (N_8358,N_6796,N_7131);
nor U8359 (N_8359,N_6957,N_6129);
nor U8360 (N_8360,N_6759,N_7037);
xor U8361 (N_8361,N_6610,N_6485);
or U8362 (N_8362,N_6556,N_7167);
and U8363 (N_8363,N_7105,N_6760);
nor U8364 (N_8364,N_6335,N_6128);
and U8365 (N_8365,N_6492,N_6304);
and U8366 (N_8366,N_6660,N_6634);
xnor U8367 (N_8367,N_7027,N_6599);
and U8368 (N_8368,N_6926,N_6462);
nand U8369 (N_8369,N_6542,N_6692);
xnor U8370 (N_8370,N_6794,N_6227);
or U8371 (N_8371,N_6110,N_6679);
nand U8372 (N_8372,N_7118,N_6817);
xor U8373 (N_8373,N_6421,N_7183);
xnor U8374 (N_8374,N_6865,N_6566);
nand U8375 (N_8375,N_6917,N_6110);
nand U8376 (N_8376,N_6048,N_6568);
and U8377 (N_8377,N_6312,N_6344);
nand U8378 (N_8378,N_6717,N_6311);
and U8379 (N_8379,N_7090,N_6585);
xor U8380 (N_8380,N_6906,N_7061);
xor U8381 (N_8381,N_7004,N_6240);
nand U8382 (N_8382,N_6570,N_6309);
nor U8383 (N_8383,N_6837,N_6124);
xnor U8384 (N_8384,N_6611,N_6676);
nor U8385 (N_8385,N_6666,N_6617);
nand U8386 (N_8386,N_6893,N_6815);
nand U8387 (N_8387,N_7044,N_6931);
xor U8388 (N_8388,N_6361,N_6919);
xor U8389 (N_8389,N_6503,N_6983);
nor U8390 (N_8390,N_6449,N_6490);
or U8391 (N_8391,N_6279,N_6493);
nand U8392 (N_8392,N_6549,N_6992);
nand U8393 (N_8393,N_6542,N_6757);
or U8394 (N_8394,N_6647,N_6225);
and U8395 (N_8395,N_6908,N_6281);
nand U8396 (N_8396,N_7034,N_6418);
nor U8397 (N_8397,N_6303,N_6158);
xnor U8398 (N_8398,N_6246,N_6078);
or U8399 (N_8399,N_6838,N_6912);
and U8400 (N_8400,N_8287,N_7411);
or U8401 (N_8401,N_7892,N_8104);
nor U8402 (N_8402,N_7498,N_7744);
and U8403 (N_8403,N_8351,N_8266);
nand U8404 (N_8404,N_7615,N_7624);
nor U8405 (N_8405,N_7972,N_7977);
nand U8406 (N_8406,N_7329,N_8067);
nor U8407 (N_8407,N_7726,N_7651);
or U8408 (N_8408,N_8007,N_7803);
or U8409 (N_8409,N_7525,N_8241);
nand U8410 (N_8410,N_7809,N_7682);
nand U8411 (N_8411,N_7938,N_7688);
nand U8412 (N_8412,N_8196,N_7221);
nor U8413 (N_8413,N_7420,N_7566);
nor U8414 (N_8414,N_7738,N_7272);
and U8415 (N_8415,N_7569,N_8210);
xor U8416 (N_8416,N_7655,N_8315);
or U8417 (N_8417,N_8192,N_8302);
and U8418 (N_8418,N_7294,N_7823);
or U8419 (N_8419,N_7259,N_7492);
nand U8420 (N_8420,N_7485,N_8329);
xor U8421 (N_8421,N_8167,N_8061);
xor U8422 (N_8422,N_7790,N_7969);
nand U8423 (N_8423,N_7465,N_7528);
nand U8424 (N_8424,N_8224,N_7399);
nor U8425 (N_8425,N_8347,N_7786);
xor U8426 (N_8426,N_7543,N_7880);
and U8427 (N_8427,N_7816,N_7585);
xnor U8428 (N_8428,N_8326,N_7451);
xnor U8429 (N_8429,N_8040,N_7495);
or U8430 (N_8430,N_7680,N_8060);
xor U8431 (N_8431,N_8166,N_7335);
nand U8432 (N_8432,N_7351,N_7521);
xnor U8433 (N_8433,N_7674,N_8298);
xor U8434 (N_8434,N_7642,N_7971);
nor U8435 (N_8435,N_8269,N_7445);
xnor U8436 (N_8436,N_7347,N_7519);
xnor U8437 (N_8437,N_7540,N_7866);
xor U8438 (N_8438,N_7441,N_8373);
xor U8439 (N_8439,N_7243,N_7960);
or U8440 (N_8440,N_7513,N_7340);
nand U8441 (N_8441,N_7722,N_7487);
and U8442 (N_8442,N_7978,N_7665);
and U8443 (N_8443,N_7862,N_8074);
and U8444 (N_8444,N_8297,N_8179);
nor U8445 (N_8445,N_8395,N_7620);
nor U8446 (N_8446,N_8130,N_8370);
or U8447 (N_8447,N_7906,N_7419);
nor U8448 (N_8448,N_8173,N_7743);
nand U8449 (N_8449,N_7919,N_8069);
xor U8450 (N_8450,N_8375,N_8139);
or U8451 (N_8451,N_7845,N_7872);
xor U8452 (N_8452,N_8125,N_7282);
and U8453 (N_8453,N_7962,N_7780);
or U8454 (N_8454,N_8265,N_8057);
nor U8455 (N_8455,N_7200,N_8378);
xnor U8456 (N_8456,N_8170,N_7380);
nand U8457 (N_8457,N_8252,N_7501);
or U8458 (N_8458,N_8384,N_8212);
and U8459 (N_8459,N_7493,N_7404);
nor U8460 (N_8460,N_7929,N_7580);
xnor U8461 (N_8461,N_7607,N_7240);
and U8462 (N_8462,N_7372,N_7371);
nand U8463 (N_8463,N_7810,N_7395);
nand U8464 (N_8464,N_7413,N_7705);
nor U8465 (N_8465,N_7770,N_7911);
and U8466 (N_8466,N_7409,N_7959);
nand U8467 (N_8467,N_7516,N_7853);
xor U8468 (N_8468,N_7625,N_7314);
nand U8469 (N_8469,N_7988,N_8320);
and U8470 (N_8470,N_8115,N_7251);
nand U8471 (N_8471,N_7937,N_7633);
nor U8472 (N_8472,N_8288,N_8133);
or U8473 (N_8473,N_8156,N_7337);
nor U8474 (N_8474,N_7366,N_8162);
nor U8475 (N_8475,N_7250,N_8394);
and U8476 (N_8476,N_7599,N_8289);
nor U8477 (N_8477,N_8312,N_8271);
nand U8478 (N_8478,N_7826,N_7631);
and U8479 (N_8479,N_7381,N_7812);
or U8480 (N_8480,N_7242,N_7747);
nor U8481 (N_8481,N_8286,N_7981);
nand U8482 (N_8482,N_7904,N_7632);
and U8483 (N_8483,N_7849,N_8092);
or U8484 (N_8484,N_7561,N_7795);
nand U8485 (N_8485,N_7568,N_7332);
and U8486 (N_8486,N_7547,N_7614);
and U8487 (N_8487,N_8119,N_8168);
or U8488 (N_8488,N_7634,N_8023);
xor U8489 (N_8489,N_7204,N_8025);
or U8490 (N_8490,N_7644,N_7458);
or U8491 (N_8491,N_8232,N_8377);
nand U8492 (N_8492,N_7377,N_8282);
nor U8493 (N_8493,N_7373,N_7753);
and U8494 (N_8494,N_7944,N_7742);
and U8495 (N_8495,N_7731,N_8042);
xnor U8496 (N_8496,N_7328,N_8111);
nor U8497 (N_8497,N_7920,N_7652);
and U8498 (N_8498,N_7418,N_7800);
or U8499 (N_8499,N_7414,N_8242);
and U8500 (N_8500,N_7980,N_7462);
or U8501 (N_8501,N_8360,N_7279);
xor U8502 (N_8502,N_8236,N_7496);
xor U8503 (N_8503,N_7215,N_7618);
xnor U8504 (N_8504,N_8274,N_7613);
nor U8505 (N_8505,N_8381,N_7439);
or U8506 (N_8506,N_7523,N_7338);
nor U8507 (N_8507,N_7581,N_7905);
nand U8508 (N_8508,N_7899,N_7252);
nor U8509 (N_8509,N_8197,N_7212);
and U8510 (N_8510,N_8134,N_7914);
nor U8511 (N_8511,N_7740,N_8002);
nand U8512 (N_8512,N_7942,N_8260);
xnor U8513 (N_8513,N_7352,N_8031);
nor U8514 (N_8514,N_8358,N_8335);
nor U8515 (N_8515,N_7604,N_8295);
and U8516 (N_8516,N_7894,N_7668);
nor U8517 (N_8517,N_8285,N_8026);
or U8518 (N_8518,N_7879,N_7921);
nor U8519 (N_8519,N_7497,N_7236);
or U8520 (N_8520,N_7284,N_7646);
and U8521 (N_8521,N_7684,N_7865);
nand U8522 (N_8522,N_8359,N_7428);
and U8523 (N_8523,N_7877,N_7951);
or U8524 (N_8524,N_7900,N_7400);
nor U8525 (N_8525,N_8293,N_7903);
xnor U8526 (N_8526,N_7341,N_7650);
nor U8527 (N_8527,N_8141,N_7510);
nand U8528 (N_8528,N_7601,N_8157);
or U8529 (N_8529,N_7720,N_8250);
nand U8530 (N_8530,N_7887,N_7896);
or U8531 (N_8531,N_7994,N_7602);
nand U8532 (N_8532,N_8207,N_7482);
nand U8533 (N_8533,N_7735,N_7793);
xnor U8534 (N_8534,N_7302,N_7410);
nand U8535 (N_8535,N_8277,N_7691);
xnor U8536 (N_8536,N_7608,N_7846);
and U8537 (N_8537,N_7721,N_8019);
nor U8538 (N_8538,N_8225,N_7966);
nor U8539 (N_8539,N_7574,N_7334);
nor U8540 (N_8540,N_7626,N_7955);
nor U8541 (N_8541,N_7368,N_7435);
nor U8542 (N_8542,N_7605,N_7756);
and U8543 (N_8543,N_7883,N_8055);
nand U8544 (N_8544,N_7564,N_7453);
xor U8545 (N_8545,N_7474,N_8175);
or U8546 (N_8546,N_7769,N_7713);
and U8547 (N_8547,N_7600,N_7692);
nor U8548 (N_8548,N_7354,N_7771);
and U8549 (N_8549,N_8107,N_7774);
nor U8550 (N_8550,N_7397,N_7822);
nand U8551 (N_8551,N_8362,N_7235);
nor U8552 (N_8552,N_7550,N_7270);
xnor U8553 (N_8553,N_8244,N_7830);
or U8554 (N_8554,N_7577,N_8331);
nor U8555 (N_8555,N_7464,N_7761);
nand U8556 (N_8556,N_7468,N_7289);
nor U8557 (N_8557,N_7255,N_8386);
nor U8558 (N_8558,N_7776,N_7385);
and U8559 (N_8559,N_8322,N_7998);
xor U8560 (N_8560,N_7670,N_7854);
and U8561 (N_8561,N_7583,N_8016);
xnor U8562 (N_8562,N_7783,N_7229);
xnor U8563 (N_8563,N_7333,N_7802);
xnor U8564 (N_8564,N_7737,N_7426);
nor U8565 (N_8565,N_7544,N_8138);
and U8566 (N_8566,N_7855,N_7820);
and U8567 (N_8567,N_7396,N_7842);
nor U8568 (N_8568,N_7836,N_8369);
and U8569 (N_8569,N_7787,N_8363);
nor U8570 (N_8570,N_7739,N_7637);
nand U8571 (N_8571,N_7517,N_7526);
nor U8572 (N_8572,N_7481,N_7751);
and U8573 (N_8573,N_8108,N_8233);
xnor U8574 (N_8574,N_7548,N_7835);
or U8575 (N_8575,N_8276,N_7433);
nand U8576 (N_8576,N_7384,N_8146);
xnor U8577 (N_8577,N_7870,N_8230);
nor U8578 (N_8578,N_8098,N_8171);
nor U8579 (N_8579,N_7365,N_7709);
nand U8580 (N_8580,N_7993,N_7764);
xor U8581 (N_8581,N_8261,N_8065);
or U8582 (N_8582,N_8063,N_8264);
xor U8583 (N_8583,N_7589,N_7362);
or U8584 (N_8584,N_7992,N_7344);
nand U8585 (N_8585,N_8334,N_8095);
or U8586 (N_8586,N_8313,N_7274);
xnor U8587 (N_8587,N_8050,N_7232);
nand U8588 (N_8588,N_7594,N_7443);
nor U8589 (N_8589,N_7330,N_8101);
or U8590 (N_8590,N_7719,N_7609);
and U8591 (N_8591,N_7661,N_7570);
and U8592 (N_8592,N_7687,N_8372);
or U8593 (N_8593,N_8137,N_8304);
xnor U8594 (N_8594,N_8237,N_7370);
xor U8595 (N_8595,N_7741,N_7407);
nand U8596 (N_8596,N_7991,N_8151);
or U8597 (N_8597,N_7582,N_7958);
or U8598 (N_8598,N_7961,N_7940);
nand U8599 (N_8599,N_7520,N_7898);
xor U8600 (N_8600,N_7246,N_7216);
nor U8601 (N_8601,N_8085,N_7832);
nand U8602 (N_8602,N_7275,N_8072);
and U8603 (N_8603,N_8239,N_8036);
xor U8604 (N_8604,N_7349,N_7767);
and U8605 (N_8605,N_7703,N_8164);
or U8606 (N_8606,N_7933,N_7621);
and U8607 (N_8607,N_7273,N_7488);
or U8608 (N_8608,N_7950,N_7657);
nand U8609 (N_8609,N_7533,N_7477);
nand U8610 (N_8610,N_7527,N_7659);
nand U8611 (N_8611,N_7936,N_7873);
and U8612 (N_8612,N_7374,N_7290);
xor U8613 (N_8613,N_8309,N_7808);
nand U8614 (N_8614,N_7825,N_8273);
nand U8615 (N_8615,N_7320,N_8317);
nor U8616 (N_8616,N_7804,N_7491);
and U8617 (N_8617,N_7454,N_7375);
and U8618 (N_8618,N_8314,N_8380);
xnor U8619 (N_8619,N_7319,N_7717);
nor U8620 (N_8620,N_7645,N_7857);
nand U8621 (N_8621,N_7871,N_8201);
nand U8622 (N_8622,N_8080,N_8012);
nor U8623 (N_8623,N_7518,N_8397);
xor U8624 (N_8624,N_7909,N_7502);
or U8625 (N_8625,N_7505,N_8299);
or U8626 (N_8626,N_7745,N_7405);
nand U8627 (N_8627,N_7326,N_7698);
nand U8628 (N_8628,N_7755,N_7442);
xor U8629 (N_8629,N_8364,N_8136);
nor U8630 (N_8630,N_7309,N_7423);
or U8631 (N_8631,N_7224,N_8020);
and U8632 (N_8632,N_8345,N_7785);
and U8633 (N_8633,N_8038,N_7323);
and U8634 (N_8634,N_8056,N_8033);
xnor U8635 (N_8635,N_7641,N_7847);
and U8636 (N_8636,N_7421,N_7922);
xor U8637 (N_8637,N_8300,N_7792);
xnor U8638 (N_8638,N_7943,N_7386);
nand U8639 (N_8639,N_8216,N_8219);
nor U8640 (N_8640,N_8118,N_7286);
nor U8641 (N_8641,N_8393,N_7974);
nand U8642 (N_8642,N_8017,N_8346);
xnor U8643 (N_8643,N_7534,N_7262);
nand U8644 (N_8644,N_7934,N_7918);
and U8645 (N_8645,N_7296,N_7401);
nor U8646 (N_8646,N_8245,N_7856);
nand U8647 (N_8647,N_8010,N_7440);
or U8648 (N_8648,N_8316,N_8319);
xor U8649 (N_8649,N_7554,N_7663);
or U8650 (N_8650,N_8218,N_8052);
xor U8651 (N_8651,N_7336,N_7575);
xnor U8652 (N_8652,N_7715,N_7844);
nor U8653 (N_8653,N_7701,N_8292);
nand U8654 (N_8654,N_7532,N_7990);
and U8655 (N_8655,N_7798,N_7382);
nand U8656 (N_8656,N_7486,N_7814);
and U8657 (N_8657,N_7983,N_8039);
nor U8658 (N_8658,N_7598,N_7559);
nor U8659 (N_8659,N_8024,N_7379);
xor U8660 (N_8660,N_8015,N_7287);
nor U8661 (N_8661,N_8140,N_8291);
and U8662 (N_8662,N_7402,N_7597);
and U8663 (N_8663,N_7310,N_8349);
nor U8664 (N_8664,N_7799,N_7868);
xnor U8665 (N_8665,N_7393,N_7447);
or U8666 (N_8666,N_8046,N_8235);
xor U8667 (N_8667,N_7712,N_7724);
nand U8668 (N_8668,N_7265,N_7245);
or U8669 (N_8669,N_8399,N_7834);
or U8670 (N_8670,N_7924,N_7263);
xnor U8671 (N_8671,N_8388,N_7662);
nor U8672 (N_8672,N_7324,N_7886);
nor U8673 (N_8673,N_7932,N_8228);
nand U8674 (N_8674,N_7711,N_7640);
or U8675 (N_8675,N_7696,N_8217);
or U8676 (N_8676,N_8160,N_8000);
xor U8677 (N_8677,N_7579,N_8323);
and U8678 (N_8678,N_7471,N_8051);
xnor U8679 (N_8679,N_8268,N_7925);
or U8680 (N_8680,N_8185,N_7506);
or U8681 (N_8681,N_7864,N_7733);
or U8682 (N_8682,N_8206,N_8357);
nor U8683 (N_8683,N_7444,N_7466);
and U8684 (N_8684,N_7541,N_7412);
nand U8685 (N_8685,N_7629,N_8145);
or U8686 (N_8686,N_7673,N_7233);
nor U8687 (N_8687,N_7995,N_8340);
nand U8688 (N_8688,N_7536,N_7630);
nor U8689 (N_8689,N_7389,N_8177);
nand U8690 (N_8690,N_7875,N_7360);
xnor U8691 (N_8691,N_7850,N_8041);
and U8692 (N_8692,N_7297,N_7638);
or U8693 (N_8693,N_8257,N_7611);
xnor U8694 (N_8694,N_8249,N_8120);
or U8695 (N_8695,N_7438,N_8066);
xnor U8696 (N_8696,N_8221,N_7285);
and U8697 (N_8697,N_7467,N_8321);
nor U8698 (N_8698,N_7965,N_7876);
and U8699 (N_8699,N_8213,N_7591);
nand U8700 (N_8700,N_8089,N_7267);
and U8701 (N_8701,N_8352,N_7860);
nand U8702 (N_8702,N_8090,N_7325);
nand U8703 (N_8703,N_8082,N_8374);
and U8704 (N_8704,N_8281,N_7472);
xor U8705 (N_8705,N_7238,N_7450);
nand U8706 (N_8706,N_7213,N_8009);
or U8707 (N_8707,N_8256,N_8021);
nand U8708 (N_8708,N_8011,N_7763);
or U8709 (N_8709,N_7895,N_7619);
nor U8710 (N_8710,N_7476,N_7693);
or U8711 (N_8711,N_8307,N_7503);
and U8712 (N_8712,N_7230,N_8032);
nand U8713 (N_8713,N_8106,N_8356);
nand U8714 (N_8714,N_8034,N_8076);
or U8715 (N_8715,N_7343,N_7913);
nor U8716 (N_8716,N_7346,N_7298);
nand U8717 (N_8717,N_7432,N_7313);
xnor U8718 (N_8718,N_7562,N_7775);
and U8719 (N_8719,N_7636,N_7801);
xor U8720 (N_8720,N_7507,N_8077);
or U8721 (N_8721,N_7436,N_8018);
and U8722 (N_8722,N_7654,N_7975);
nor U8723 (N_8723,N_7869,N_7345);
or U8724 (N_8724,N_7364,N_7478);
xor U8725 (N_8725,N_7839,N_8310);
and U8726 (N_8726,N_8113,N_8325);
and U8727 (N_8727,N_7817,N_7766);
and U8728 (N_8728,N_8172,N_7535);
and U8729 (N_8729,N_7963,N_7308);
or U8730 (N_8730,N_8396,N_7675);
xor U8731 (N_8731,N_7214,N_7578);
nand U8732 (N_8732,N_7928,N_7271);
or U8733 (N_8733,N_7268,N_7789);
or U8734 (N_8734,N_7653,N_8348);
xor U8735 (N_8735,N_7292,N_7734);
and U8736 (N_8736,N_7512,N_7976);
nand U8737 (N_8737,N_7264,N_7237);
and U8738 (N_8738,N_7768,N_7571);
and U8739 (N_8739,N_7821,N_7538);
or U8740 (N_8740,N_8391,N_7595);
nand U8741 (N_8741,N_8028,N_8267);
xor U8742 (N_8742,N_7218,N_8147);
nand U8743 (N_8743,N_7430,N_8301);
nor U8744 (N_8744,N_7730,N_7796);
xor U8745 (N_8745,N_7254,N_8376);
xor U8746 (N_8746,N_8182,N_7778);
or U8747 (N_8747,N_7228,N_7678);
nor U8748 (N_8748,N_7210,N_7996);
nand U8749 (N_8749,N_7446,N_7891);
nor U8750 (N_8750,N_7459,N_8068);
or U8751 (N_8751,N_7514,N_7773);
xor U8752 (N_8752,N_8103,N_7283);
xnor U8753 (N_8753,N_7448,N_7782);
and U8754 (N_8754,N_7457,N_8220);
nand U8755 (N_8755,N_8014,N_7939);
xor U8756 (N_8756,N_7952,N_7378);
nor U8757 (N_8757,N_7348,N_7838);
nor U8758 (N_8758,N_7217,N_7572);
or U8759 (N_8759,N_7322,N_8142);
or U8760 (N_8760,N_7556,N_7269);
nor U8761 (N_8761,N_7878,N_7388);
nand U8762 (N_8762,N_7718,N_8128);
nand U8763 (N_8763,N_8251,N_8193);
or U8764 (N_8764,N_8121,N_8129);
or U8765 (N_8765,N_7280,N_7278);
or U8766 (N_8766,N_8338,N_7261);
or U8767 (N_8767,N_8383,N_7777);
and U8768 (N_8768,N_8344,N_7356);
nand U8769 (N_8769,N_7431,N_7479);
xor U8770 (N_8770,N_7649,N_8081);
or U8771 (N_8771,N_7247,N_8027);
nand U8772 (N_8772,N_7707,N_8169);
and U8773 (N_8773,N_7949,N_7511);
xor U8774 (N_8774,N_7927,N_8342);
nand U8775 (N_8775,N_7954,N_7306);
nor U8776 (N_8776,N_7628,N_8385);
and U8777 (N_8777,N_7758,N_8387);
nor U8778 (N_8778,N_7957,N_7997);
or U8779 (N_8779,N_8200,N_8227);
xnor U8780 (N_8780,N_7484,N_7392);
xnor U8781 (N_8781,N_7676,N_7930);
or U8782 (N_8782,N_8231,N_7461);
xnor U8783 (N_8783,N_8006,N_8075);
or U8784 (N_8784,N_8222,N_7964);
and U8785 (N_8785,N_8116,N_7725);
xor U8786 (N_8786,N_7848,N_7987);
xnor U8787 (N_8787,N_8030,N_8270);
or U8788 (N_8788,N_7398,N_7425);
or U8789 (N_8789,N_7545,N_7858);
xor U8790 (N_8790,N_8091,N_7586);
and U8791 (N_8791,N_8202,N_8368);
xnor U8792 (N_8792,N_7353,N_7623);
nand U8793 (N_8793,N_7383,N_7647);
nor U8794 (N_8794,N_8094,N_7686);
nand U8795 (N_8795,N_7475,N_8070);
and U8796 (N_8796,N_8263,N_7304);
nand U8797 (N_8797,N_7391,N_8152);
nand U8798 (N_8798,N_7610,N_7449);
and U8799 (N_8799,N_7695,N_7480);
xnor U8800 (N_8800,N_8110,N_7982);
and U8801 (N_8801,N_8258,N_7403);
or U8802 (N_8802,N_7530,N_7815);
or U8803 (N_8803,N_7557,N_8238);
and U8804 (N_8804,N_8247,N_8045);
nor U8805 (N_8805,N_7897,N_8004);
and U8806 (N_8806,N_7437,N_7606);
xor U8807 (N_8807,N_8366,N_8187);
xor U8808 (N_8808,N_7300,N_7301);
and U8809 (N_8809,N_7794,N_7757);
xor U8810 (N_8810,N_8083,N_7408);
nand U8811 (N_8811,N_8163,N_7946);
or U8812 (N_8812,N_7361,N_8203);
nor U8813 (N_8813,N_7509,N_7874);
xor U8814 (N_8814,N_8022,N_8184);
xnor U8815 (N_8815,N_8336,N_8339);
nand U8816 (N_8816,N_8054,N_7881);
nor U8817 (N_8817,N_7728,N_7627);
or U8818 (N_8818,N_8390,N_7489);
nor U8819 (N_8819,N_7658,N_7683);
or U8820 (N_8820,N_8254,N_7941);
nand U8821 (N_8821,N_8341,N_7797);
nand U8822 (N_8822,N_7664,N_7256);
nand U8823 (N_8823,N_7754,N_8332);
xor U8824 (N_8824,N_7901,N_8240);
nor U8825 (N_8825,N_7549,N_7843);
xor U8826 (N_8826,N_7788,N_7394);
nor U8827 (N_8827,N_7318,N_7291);
xor U8828 (N_8828,N_8109,N_8333);
and U8829 (N_8829,N_7714,N_8096);
nor U8830 (N_8830,N_7205,N_8371);
xor U8831 (N_8831,N_7967,N_7916);
or U8832 (N_8832,N_8246,N_8278);
nand U8833 (N_8833,N_7910,N_7555);
nor U8834 (N_8834,N_7376,N_8029);
nor U8835 (N_8835,N_8234,N_7704);
xnor U8836 (N_8836,N_7305,N_8035);
nand U8837 (N_8837,N_8283,N_7303);
nand U8838 (N_8838,N_7494,N_7772);
nand U8839 (N_8839,N_7931,N_7827);
or U8840 (N_8840,N_8044,N_7603);
nand U8841 (N_8841,N_7546,N_7805);
xnor U8842 (N_8842,N_7915,N_7276);
and U8843 (N_8843,N_7833,N_8262);
or U8844 (N_8844,N_7463,N_8303);
xnor U8845 (N_8845,N_7429,N_7266);
or U8846 (N_8846,N_7884,N_8350);
and U8847 (N_8847,N_8229,N_7357);
or U8848 (N_8848,N_7945,N_7483);
nor U8849 (N_8849,N_7765,N_8208);
or U8850 (N_8850,N_7973,N_8191);
nor U8851 (N_8851,N_7784,N_8343);
nor U8852 (N_8852,N_7315,N_8355);
nand U8853 (N_8853,N_7708,N_7612);
xnor U8854 (N_8854,N_7202,N_7560);
and U8855 (N_8855,N_7588,N_7837);
nand U8856 (N_8856,N_7551,N_7907);
xor U8857 (N_8857,N_7359,N_8280);
and U8858 (N_8858,N_8209,N_8176);
xor U8859 (N_8859,N_7749,N_7706);
or U8860 (N_8860,N_8311,N_7355);
xnor U8861 (N_8861,N_7953,N_7750);
nand U8862 (N_8862,N_8155,N_7779);
nand U8863 (N_8863,N_8308,N_7417);
xor U8864 (N_8864,N_8058,N_8165);
or U8865 (N_8865,N_7327,N_8123);
or U8866 (N_8866,N_8306,N_7207);
or U8867 (N_8867,N_8389,N_8078);
or U8868 (N_8868,N_7867,N_7791);
or U8869 (N_8869,N_7748,N_8189);
and U8870 (N_8870,N_8154,N_7729);
nor U8871 (N_8871,N_7984,N_7656);
xor U8872 (N_8872,N_7852,N_7702);
nor U8873 (N_8873,N_8328,N_8088);
xor U8874 (N_8874,N_7759,N_8379);
and U8875 (N_8875,N_7917,N_7249);
or U8876 (N_8876,N_7912,N_7515);
and U8877 (N_8877,N_7316,N_7537);
or U8878 (N_8878,N_8354,N_8084);
xor U8879 (N_8879,N_7666,N_7222);
and U8880 (N_8880,N_8135,N_8178);
nand U8881 (N_8881,N_7893,N_8204);
nor U8882 (N_8882,N_8132,N_7989);
xor U8883 (N_8883,N_7746,N_7422);
or U8884 (N_8884,N_7452,N_8290);
or U8885 (N_8885,N_8284,N_8174);
and U8886 (N_8886,N_7293,N_8144);
xnor U8887 (N_8887,N_7225,N_7490);
nor U8888 (N_8888,N_8100,N_7312);
nor U8889 (N_8889,N_8102,N_8131);
and U8890 (N_8890,N_7552,N_8001);
or U8891 (N_8891,N_8272,N_7573);
xor U8892 (N_8892,N_7622,N_8398);
xnor U8893 (N_8893,N_8199,N_8073);
xnor U8894 (N_8894,N_8243,N_7470);
or U8895 (N_8895,N_8259,N_7635);
and U8896 (N_8896,N_7542,N_7358);
nand U8897 (N_8897,N_7339,N_7504);
or U8898 (N_8898,N_7576,N_7219);
nor U8899 (N_8899,N_7829,N_8127);
xor U8900 (N_8900,N_7567,N_7732);
xnor U8901 (N_8901,N_7807,N_7427);
nor U8902 (N_8902,N_7565,N_7669);
nor U8903 (N_8903,N_7828,N_7587);
nor U8904 (N_8904,N_7524,N_7956);
and U8905 (N_8905,N_7553,N_7277);
or U8906 (N_8906,N_7500,N_8105);
nand U8907 (N_8907,N_7239,N_7258);
xnor U8908 (N_8908,N_7762,N_7948);
xnor U8909 (N_8909,N_8124,N_7863);
xnor U8910 (N_8910,N_8086,N_8117);
xnor U8911 (N_8911,N_8305,N_8099);
nand U8912 (N_8912,N_7818,N_7689);
nor U8913 (N_8913,N_7434,N_7716);
nor U8914 (N_8914,N_8279,N_7947);
nor U8915 (N_8915,N_8255,N_8190);
xor U8916 (N_8916,N_7220,N_7985);
xor U8917 (N_8917,N_7529,N_8186);
nand U8918 (N_8918,N_8062,N_7616);
nand U8919 (N_8919,N_8097,N_7888);
nand U8920 (N_8920,N_7455,N_8226);
and U8921 (N_8921,N_8071,N_7596);
nand U8922 (N_8922,N_7979,N_8248);
nor U8923 (N_8923,N_8330,N_7889);
and U8924 (N_8924,N_7499,N_7813);
and U8925 (N_8925,N_7321,N_8382);
xnor U8926 (N_8926,N_8053,N_7257);
nor U8927 (N_8927,N_7968,N_7697);
and U8928 (N_8928,N_7643,N_7299);
nor U8929 (N_8929,N_7699,N_8059);
nand U8930 (N_8930,N_8214,N_8365);
and U8931 (N_8931,N_7908,N_8114);
and U8932 (N_8932,N_7592,N_8149);
or U8933 (N_8933,N_7752,N_8361);
and U8934 (N_8934,N_7760,N_8161);
nand U8935 (N_8935,N_8195,N_7208);
nor U8936 (N_8936,N_7781,N_7390);
nor U8937 (N_8937,N_7406,N_7201);
nand U8938 (N_8938,N_7456,N_7473);
nor U8939 (N_8939,N_7923,N_8126);
nand U8940 (N_8940,N_7679,N_7593);
and U8941 (N_8941,N_8064,N_7460);
xnor U8942 (N_8942,N_7648,N_8275);
xnor U8943 (N_8943,N_8367,N_7367);
nand U8944 (N_8944,N_8153,N_7671);
xnor U8945 (N_8945,N_7681,N_8198);
and U8946 (N_8946,N_8093,N_8013);
xor U8947 (N_8947,N_7253,N_7584);
and U8948 (N_8948,N_8087,N_7617);
nand U8949 (N_8949,N_8337,N_8223);
and U8950 (N_8950,N_7206,N_7415);
xor U8951 (N_8951,N_7824,N_7317);
or U8952 (N_8952,N_7539,N_7363);
and U8953 (N_8953,N_7986,N_7690);
xnor U8954 (N_8954,N_8183,N_8005);
or U8955 (N_8955,N_7639,N_7226);
xor U8956 (N_8956,N_7902,N_7311);
xnor U8957 (N_8957,N_8112,N_8215);
nor U8958 (N_8958,N_8194,N_8296);
or U8959 (N_8959,N_7244,N_8181);
xor U8960 (N_8960,N_7710,N_7342);
nor U8961 (N_8961,N_7522,N_7209);
xor U8962 (N_8962,N_8205,N_7369);
and U8963 (N_8963,N_7248,N_7727);
or U8964 (N_8964,N_7281,N_8148);
nor U8965 (N_8965,N_7882,N_7667);
nor U8966 (N_8966,N_7685,N_7260);
and U8967 (N_8967,N_7307,N_8188);
and U8968 (N_8968,N_7660,N_7231);
xnor U8969 (N_8969,N_7558,N_7387);
nor U8970 (N_8970,N_7859,N_7970);
and U8971 (N_8971,N_7531,N_8150);
xnor U8972 (N_8972,N_8327,N_7851);
nand U8973 (N_8973,N_7424,N_7295);
xor U8974 (N_8974,N_8353,N_7508);
nor U8975 (N_8975,N_8003,N_8180);
nand U8976 (N_8976,N_7831,N_7288);
nand U8977 (N_8977,N_7819,N_7840);
or U8978 (N_8978,N_8048,N_7203);
or U8979 (N_8979,N_8211,N_7736);
and U8980 (N_8980,N_8159,N_7234);
xnor U8981 (N_8981,N_8253,N_7885);
xor U8982 (N_8982,N_7811,N_7723);
and U8983 (N_8983,N_7926,N_8143);
nor U8984 (N_8984,N_7211,N_8324);
nand U8985 (N_8985,N_7677,N_7841);
or U8986 (N_8986,N_8318,N_8008);
xnor U8987 (N_8987,N_7999,N_8122);
xnor U8988 (N_8988,N_7241,N_7416);
and U8989 (N_8989,N_8158,N_8049);
and U8990 (N_8990,N_8294,N_7590);
nor U8991 (N_8991,N_7563,N_7331);
or U8992 (N_8992,N_7223,N_7890);
xnor U8993 (N_8993,N_8037,N_8079);
nor U8994 (N_8994,N_8047,N_7227);
or U8995 (N_8995,N_8043,N_7694);
nand U8996 (N_8996,N_8392,N_7672);
nand U8997 (N_8997,N_7700,N_7861);
nand U8998 (N_8998,N_7350,N_7806);
or U8999 (N_8999,N_7935,N_7469);
and U9000 (N_9000,N_7580,N_7788);
or U9001 (N_9001,N_8118,N_7626);
and U9002 (N_9002,N_8300,N_7610);
nand U9003 (N_9003,N_8138,N_7510);
xnor U9004 (N_9004,N_7834,N_7986);
or U9005 (N_9005,N_8144,N_7406);
nand U9006 (N_9006,N_7799,N_7918);
nor U9007 (N_9007,N_7942,N_7565);
and U9008 (N_9008,N_8351,N_7214);
and U9009 (N_9009,N_7355,N_8253);
nand U9010 (N_9010,N_8012,N_8382);
or U9011 (N_9011,N_8034,N_7407);
nor U9012 (N_9012,N_7775,N_7916);
nand U9013 (N_9013,N_7307,N_7592);
and U9014 (N_9014,N_7717,N_8387);
nor U9015 (N_9015,N_7306,N_8274);
xor U9016 (N_9016,N_8212,N_8103);
and U9017 (N_9017,N_8260,N_8268);
or U9018 (N_9018,N_7605,N_8133);
and U9019 (N_9019,N_8182,N_7996);
nor U9020 (N_9020,N_7964,N_7364);
and U9021 (N_9021,N_8091,N_7499);
and U9022 (N_9022,N_7212,N_7667);
nand U9023 (N_9023,N_7235,N_7801);
nor U9024 (N_9024,N_8353,N_7267);
or U9025 (N_9025,N_8124,N_7778);
and U9026 (N_9026,N_7758,N_7753);
and U9027 (N_9027,N_7652,N_8084);
xor U9028 (N_9028,N_7300,N_7765);
nor U9029 (N_9029,N_8366,N_7646);
nor U9030 (N_9030,N_8225,N_7869);
or U9031 (N_9031,N_8147,N_7485);
and U9032 (N_9032,N_8019,N_8277);
nand U9033 (N_9033,N_7252,N_7567);
xnor U9034 (N_9034,N_8254,N_7898);
nand U9035 (N_9035,N_7839,N_7452);
nor U9036 (N_9036,N_7207,N_7607);
nand U9037 (N_9037,N_8371,N_7239);
nand U9038 (N_9038,N_7523,N_7317);
and U9039 (N_9039,N_7516,N_7429);
nand U9040 (N_9040,N_7344,N_7967);
nand U9041 (N_9041,N_7215,N_7554);
and U9042 (N_9042,N_7952,N_7222);
and U9043 (N_9043,N_7305,N_8072);
xnor U9044 (N_9044,N_8161,N_7980);
or U9045 (N_9045,N_7375,N_8141);
xnor U9046 (N_9046,N_7902,N_7602);
nand U9047 (N_9047,N_7460,N_7704);
or U9048 (N_9048,N_7358,N_7319);
or U9049 (N_9049,N_8107,N_7482);
and U9050 (N_9050,N_7379,N_7955);
or U9051 (N_9051,N_7849,N_7453);
xnor U9052 (N_9052,N_7828,N_7578);
nor U9053 (N_9053,N_7335,N_8282);
nand U9054 (N_9054,N_7861,N_8092);
and U9055 (N_9055,N_7235,N_7777);
nor U9056 (N_9056,N_8253,N_7756);
or U9057 (N_9057,N_7574,N_7587);
nand U9058 (N_9058,N_7324,N_7770);
xor U9059 (N_9059,N_8322,N_7336);
nand U9060 (N_9060,N_7755,N_7745);
nor U9061 (N_9061,N_8350,N_7328);
nand U9062 (N_9062,N_7915,N_8168);
or U9063 (N_9063,N_7441,N_8122);
xor U9064 (N_9064,N_7922,N_7942);
nor U9065 (N_9065,N_7688,N_7979);
nand U9066 (N_9066,N_8320,N_7481);
nor U9067 (N_9067,N_8312,N_7936);
nor U9068 (N_9068,N_8088,N_7729);
xnor U9069 (N_9069,N_7987,N_7672);
and U9070 (N_9070,N_8276,N_7746);
xor U9071 (N_9071,N_8135,N_7310);
or U9072 (N_9072,N_7218,N_7838);
nor U9073 (N_9073,N_7242,N_7506);
nor U9074 (N_9074,N_7370,N_7606);
and U9075 (N_9075,N_7464,N_7402);
or U9076 (N_9076,N_7839,N_7628);
or U9077 (N_9077,N_7994,N_7203);
or U9078 (N_9078,N_8197,N_8325);
nand U9079 (N_9079,N_7354,N_7830);
nand U9080 (N_9080,N_7339,N_8399);
and U9081 (N_9081,N_8090,N_7702);
xor U9082 (N_9082,N_7347,N_7234);
or U9083 (N_9083,N_7601,N_7906);
xnor U9084 (N_9084,N_7622,N_7937);
nand U9085 (N_9085,N_7725,N_8137);
nand U9086 (N_9086,N_7480,N_7764);
and U9087 (N_9087,N_7431,N_7200);
and U9088 (N_9088,N_7399,N_7799);
xor U9089 (N_9089,N_7523,N_7450);
nor U9090 (N_9090,N_8237,N_7311);
xnor U9091 (N_9091,N_8227,N_8308);
and U9092 (N_9092,N_8010,N_7327);
and U9093 (N_9093,N_8157,N_7469);
xor U9094 (N_9094,N_7450,N_7411);
xnor U9095 (N_9095,N_8286,N_8201);
xnor U9096 (N_9096,N_7486,N_8044);
xor U9097 (N_9097,N_7573,N_7240);
and U9098 (N_9098,N_8020,N_8076);
nor U9099 (N_9099,N_8343,N_8152);
or U9100 (N_9100,N_7663,N_8135);
nor U9101 (N_9101,N_8055,N_7423);
and U9102 (N_9102,N_7844,N_7463);
and U9103 (N_9103,N_7830,N_7534);
and U9104 (N_9104,N_8045,N_7776);
nor U9105 (N_9105,N_7283,N_7919);
nor U9106 (N_9106,N_7746,N_7998);
or U9107 (N_9107,N_7899,N_8051);
and U9108 (N_9108,N_7622,N_7200);
nand U9109 (N_9109,N_7909,N_7253);
nand U9110 (N_9110,N_8364,N_7744);
nor U9111 (N_9111,N_8204,N_7881);
nor U9112 (N_9112,N_7684,N_7825);
xnor U9113 (N_9113,N_7441,N_8284);
nor U9114 (N_9114,N_8350,N_7829);
nor U9115 (N_9115,N_7642,N_7675);
nor U9116 (N_9116,N_7785,N_8241);
or U9117 (N_9117,N_8058,N_7840);
or U9118 (N_9118,N_7686,N_7799);
xor U9119 (N_9119,N_7394,N_7839);
nand U9120 (N_9120,N_7518,N_8172);
xnor U9121 (N_9121,N_7209,N_7989);
or U9122 (N_9122,N_7415,N_7277);
nor U9123 (N_9123,N_7608,N_8189);
and U9124 (N_9124,N_7551,N_8273);
and U9125 (N_9125,N_8169,N_8338);
or U9126 (N_9126,N_8117,N_8312);
nor U9127 (N_9127,N_8088,N_7270);
and U9128 (N_9128,N_7385,N_7948);
xnor U9129 (N_9129,N_7791,N_8378);
nand U9130 (N_9130,N_7234,N_8232);
or U9131 (N_9131,N_7656,N_7487);
and U9132 (N_9132,N_8109,N_8332);
nor U9133 (N_9133,N_7669,N_7854);
nor U9134 (N_9134,N_8392,N_7374);
nand U9135 (N_9135,N_7586,N_7881);
or U9136 (N_9136,N_7818,N_7232);
xor U9137 (N_9137,N_7524,N_7959);
or U9138 (N_9138,N_7718,N_8001);
nand U9139 (N_9139,N_8012,N_7919);
and U9140 (N_9140,N_7714,N_8090);
or U9141 (N_9141,N_7757,N_7905);
or U9142 (N_9142,N_7893,N_7643);
and U9143 (N_9143,N_8042,N_7730);
or U9144 (N_9144,N_7863,N_8380);
xor U9145 (N_9145,N_7961,N_8398);
nor U9146 (N_9146,N_8035,N_7584);
nor U9147 (N_9147,N_8038,N_8397);
nand U9148 (N_9148,N_8371,N_8355);
or U9149 (N_9149,N_7408,N_7433);
and U9150 (N_9150,N_7379,N_7334);
nand U9151 (N_9151,N_8379,N_8215);
or U9152 (N_9152,N_7478,N_7472);
nand U9153 (N_9153,N_7585,N_8353);
xnor U9154 (N_9154,N_8344,N_7501);
or U9155 (N_9155,N_8255,N_7621);
nor U9156 (N_9156,N_7996,N_7655);
and U9157 (N_9157,N_8107,N_8096);
and U9158 (N_9158,N_7701,N_8213);
or U9159 (N_9159,N_7483,N_7828);
nor U9160 (N_9160,N_7898,N_7999);
and U9161 (N_9161,N_7410,N_7249);
nand U9162 (N_9162,N_7731,N_7650);
nand U9163 (N_9163,N_7585,N_8099);
xor U9164 (N_9164,N_8088,N_8129);
and U9165 (N_9165,N_7304,N_7820);
or U9166 (N_9166,N_8125,N_7980);
xor U9167 (N_9167,N_7589,N_7746);
nor U9168 (N_9168,N_7432,N_8358);
and U9169 (N_9169,N_8285,N_7610);
nand U9170 (N_9170,N_7410,N_8034);
xnor U9171 (N_9171,N_8206,N_8316);
nand U9172 (N_9172,N_8303,N_7450);
nand U9173 (N_9173,N_8248,N_7499);
or U9174 (N_9174,N_7940,N_7454);
xnor U9175 (N_9175,N_8296,N_7600);
nor U9176 (N_9176,N_8313,N_7927);
or U9177 (N_9177,N_7550,N_7735);
nand U9178 (N_9178,N_7494,N_7657);
or U9179 (N_9179,N_7331,N_8023);
xnor U9180 (N_9180,N_8209,N_8041);
and U9181 (N_9181,N_7891,N_8281);
nand U9182 (N_9182,N_7289,N_7664);
xor U9183 (N_9183,N_8200,N_7549);
xor U9184 (N_9184,N_7413,N_7689);
or U9185 (N_9185,N_7670,N_8251);
or U9186 (N_9186,N_7535,N_8362);
nand U9187 (N_9187,N_7362,N_8061);
and U9188 (N_9188,N_8143,N_7561);
xnor U9189 (N_9189,N_7863,N_7365);
nor U9190 (N_9190,N_8037,N_8393);
nor U9191 (N_9191,N_7334,N_7864);
and U9192 (N_9192,N_7557,N_8263);
nand U9193 (N_9193,N_7240,N_8135);
nor U9194 (N_9194,N_7521,N_7846);
xnor U9195 (N_9195,N_7454,N_8295);
nand U9196 (N_9196,N_8368,N_7602);
nand U9197 (N_9197,N_8291,N_7671);
and U9198 (N_9198,N_7635,N_7295);
or U9199 (N_9199,N_8107,N_7264);
or U9200 (N_9200,N_7741,N_8073);
nor U9201 (N_9201,N_7512,N_7919);
nand U9202 (N_9202,N_7426,N_7273);
or U9203 (N_9203,N_8339,N_8149);
or U9204 (N_9204,N_8202,N_8347);
xor U9205 (N_9205,N_7631,N_7640);
or U9206 (N_9206,N_7225,N_8308);
nor U9207 (N_9207,N_7357,N_7424);
and U9208 (N_9208,N_7842,N_7697);
and U9209 (N_9209,N_8066,N_7242);
or U9210 (N_9210,N_7888,N_8140);
or U9211 (N_9211,N_7443,N_7807);
xnor U9212 (N_9212,N_7704,N_8032);
and U9213 (N_9213,N_8146,N_8203);
xor U9214 (N_9214,N_7536,N_7759);
or U9215 (N_9215,N_8263,N_7442);
or U9216 (N_9216,N_7469,N_8120);
and U9217 (N_9217,N_7401,N_8057);
nand U9218 (N_9218,N_7842,N_7572);
and U9219 (N_9219,N_7328,N_7204);
or U9220 (N_9220,N_8001,N_8289);
xnor U9221 (N_9221,N_7542,N_8389);
nor U9222 (N_9222,N_7874,N_7462);
nor U9223 (N_9223,N_8179,N_7665);
nor U9224 (N_9224,N_7779,N_7785);
and U9225 (N_9225,N_7816,N_7281);
nor U9226 (N_9226,N_7961,N_7284);
xnor U9227 (N_9227,N_7978,N_8317);
nor U9228 (N_9228,N_7847,N_8364);
nor U9229 (N_9229,N_8131,N_7380);
or U9230 (N_9230,N_8312,N_7240);
nor U9231 (N_9231,N_8097,N_8093);
nor U9232 (N_9232,N_7775,N_8122);
and U9233 (N_9233,N_7870,N_7293);
and U9234 (N_9234,N_7775,N_7245);
nor U9235 (N_9235,N_7361,N_7660);
and U9236 (N_9236,N_7622,N_7475);
or U9237 (N_9237,N_7372,N_7775);
and U9238 (N_9238,N_7250,N_8080);
and U9239 (N_9239,N_8216,N_8303);
xnor U9240 (N_9240,N_7505,N_7773);
xnor U9241 (N_9241,N_7975,N_7888);
xnor U9242 (N_9242,N_7346,N_7602);
and U9243 (N_9243,N_8270,N_8301);
and U9244 (N_9244,N_7709,N_8345);
nor U9245 (N_9245,N_7972,N_7925);
nor U9246 (N_9246,N_7873,N_8084);
nand U9247 (N_9247,N_8049,N_8179);
nor U9248 (N_9248,N_8296,N_7710);
nor U9249 (N_9249,N_7835,N_7910);
and U9250 (N_9250,N_7993,N_8104);
xor U9251 (N_9251,N_8196,N_7629);
or U9252 (N_9252,N_7394,N_8168);
nand U9253 (N_9253,N_7841,N_7350);
nor U9254 (N_9254,N_8307,N_7648);
or U9255 (N_9255,N_7976,N_7767);
or U9256 (N_9256,N_7853,N_7735);
xor U9257 (N_9257,N_8034,N_7408);
nand U9258 (N_9258,N_8351,N_8060);
nor U9259 (N_9259,N_7670,N_7343);
nor U9260 (N_9260,N_7417,N_7468);
and U9261 (N_9261,N_8174,N_7794);
xor U9262 (N_9262,N_8176,N_8092);
or U9263 (N_9263,N_7626,N_7218);
and U9264 (N_9264,N_7426,N_7332);
or U9265 (N_9265,N_7466,N_7551);
nor U9266 (N_9266,N_7701,N_8249);
nor U9267 (N_9267,N_8010,N_7686);
and U9268 (N_9268,N_8347,N_8180);
and U9269 (N_9269,N_7791,N_7591);
nor U9270 (N_9270,N_7400,N_7814);
xnor U9271 (N_9271,N_8210,N_8226);
or U9272 (N_9272,N_8032,N_7211);
or U9273 (N_9273,N_7413,N_8055);
or U9274 (N_9274,N_7402,N_8374);
xnor U9275 (N_9275,N_7878,N_8171);
nor U9276 (N_9276,N_7339,N_7768);
and U9277 (N_9277,N_7863,N_8167);
xor U9278 (N_9278,N_7928,N_8120);
nand U9279 (N_9279,N_7471,N_8085);
and U9280 (N_9280,N_7876,N_7992);
nand U9281 (N_9281,N_7494,N_7897);
and U9282 (N_9282,N_8279,N_8013);
and U9283 (N_9283,N_8313,N_7903);
nand U9284 (N_9284,N_7943,N_7548);
or U9285 (N_9285,N_7467,N_8247);
and U9286 (N_9286,N_8137,N_8328);
xor U9287 (N_9287,N_8220,N_7685);
or U9288 (N_9288,N_7344,N_7920);
or U9289 (N_9289,N_7729,N_8174);
xnor U9290 (N_9290,N_7853,N_8062);
or U9291 (N_9291,N_7335,N_8161);
nand U9292 (N_9292,N_7478,N_8335);
and U9293 (N_9293,N_7275,N_8027);
nand U9294 (N_9294,N_8127,N_7592);
or U9295 (N_9295,N_8209,N_8200);
nand U9296 (N_9296,N_7780,N_8390);
and U9297 (N_9297,N_7968,N_7613);
nor U9298 (N_9298,N_8381,N_7855);
nor U9299 (N_9299,N_7616,N_7661);
xor U9300 (N_9300,N_7277,N_7728);
and U9301 (N_9301,N_7795,N_8142);
nor U9302 (N_9302,N_7892,N_7809);
xor U9303 (N_9303,N_8035,N_8176);
xnor U9304 (N_9304,N_7767,N_8323);
xor U9305 (N_9305,N_7220,N_8159);
nor U9306 (N_9306,N_7433,N_8227);
nand U9307 (N_9307,N_7982,N_7678);
nor U9308 (N_9308,N_7559,N_8378);
nand U9309 (N_9309,N_7943,N_7634);
nand U9310 (N_9310,N_8247,N_7327);
or U9311 (N_9311,N_8292,N_8010);
nand U9312 (N_9312,N_7802,N_7300);
or U9313 (N_9313,N_7255,N_7729);
nand U9314 (N_9314,N_7966,N_7416);
nor U9315 (N_9315,N_7892,N_8208);
xor U9316 (N_9316,N_8064,N_7445);
nor U9317 (N_9317,N_7243,N_7548);
nand U9318 (N_9318,N_7695,N_7378);
nor U9319 (N_9319,N_7330,N_8134);
nand U9320 (N_9320,N_8333,N_7772);
or U9321 (N_9321,N_7677,N_7362);
and U9322 (N_9322,N_7205,N_8341);
nor U9323 (N_9323,N_8211,N_8192);
and U9324 (N_9324,N_8093,N_8115);
xnor U9325 (N_9325,N_8142,N_7510);
nor U9326 (N_9326,N_8038,N_8008);
and U9327 (N_9327,N_7881,N_7254);
nor U9328 (N_9328,N_8278,N_7717);
and U9329 (N_9329,N_7591,N_7672);
xor U9330 (N_9330,N_7354,N_7717);
or U9331 (N_9331,N_7255,N_7844);
and U9332 (N_9332,N_8093,N_8139);
xnor U9333 (N_9333,N_7879,N_7249);
nand U9334 (N_9334,N_8070,N_7354);
nand U9335 (N_9335,N_8176,N_8207);
or U9336 (N_9336,N_7989,N_8313);
nand U9337 (N_9337,N_7827,N_7221);
and U9338 (N_9338,N_7473,N_7598);
nor U9339 (N_9339,N_7579,N_7456);
nand U9340 (N_9340,N_7483,N_7497);
xor U9341 (N_9341,N_7268,N_7945);
and U9342 (N_9342,N_8299,N_7483);
and U9343 (N_9343,N_7616,N_8387);
or U9344 (N_9344,N_8010,N_7983);
nor U9345 (N_9345,N_8096,N_8010);
xor U9346 (N_9346,N_7710,N_7265);
nor U9347 (N_9347,N_7253,N_8343);
xor U9348 (N_9348,N_7904,N_8065);
and U9349 (N_9349,N_7837,N_7506);
nand U9350 (N_9350,N_8257,N_7952);
xnor U9351 (N_9351,N_7209,N_8151);
or U9352 (N_9352,N_7324,N_8125);
xnor U9353 (N_9353,N_7700,N_7216);
nand U9354 (N_9354,N_7359,N_7365);
xnor U9355 (N_9355,N_7965,N_7433);
nand U9356 (N_9356,N_7728,N_7982);
or U9357 (N_9357,N_8053,N_7880);
or U9358 (N_9358,N_8172,N_8137);
or U9359 (N_9359,N_7336,N_8034);
nand U9360 (N_9360,N_7416,N_7870);
or U9361 (N_9361,N_8216,N_8045);
nand U9362 (N_9362,N_8005,N_7756);
nor U9363 (N_9363,N_7931,N_7312);
or U9364 (N_9364,N_7364,N_7547);
xor U9365 (N_9365,N_8102,N_8026);
xnor U9366 (N_9366,N_7690,N_7645);
and U9367 (N_9367,N_7837,N_7623);
or U9368 (N_9368,N_8009,N_7849);
nor U9369 (N_9369,N_7479,N_7563);
and U9370 (N_9370,N_7465,N_8015);
or U9371 (N_9371,N_7730,N_7637);
nand U9372 (N_9372,N_8060,N_7409);
or U9373 (N_9373,N_8179,N_8339);
xnor U9374 (N_9374,N_7528,N_7260);
nor U9375 (N_9375,N_7354,N_8269);
nor U9376 (N_9376,N_7514,N_7946);
or U9377 (N_9377,N_7764,N_7487);
and U9378 (N_9378,N_7624,N_8269);
xnor U9379 (N_9379,N_8102,N_7630);
xor U9380 (N_9380,N_8007,N_7454);
or U9381 (N_9381,N_7414,N_7851);
and U9382 (N_9382,N_7375,N_7924);
and U9383 (N_9383,N_7579,N_7960);
nor U9384 (N_9384,N_8072,N_7350);
nor U9385 (N_9385,N_7555,N_7641);
or U9386 (N_9386,N_7763,N_7761);
nor U9387 (N_9387,N_7491,N_7885);
nand U9388 (N_9388,N_7871,N_8241);
and U9389 (N_9389,N_7609,N_8179);
xnor U9390 (N_9390,N_7733,N_8129);
and U9391 (N_9391,N_8092,N_7299);
xor U9392 (N_9392,N_7958,N_8238);
or U9393 (N_9393,N_8092,N_8065);
nor U9394 (N_9394,N_8320,N_8382);
nand U9395 (N_9395,N_7571,N_8171);
and U9396 (N_9396,N_8286,N_8059);
and U9397 (N_9397,N_8172,N_7675);
or U9398 (N_9398,N_7247,N_7881);
nand U9399 (N_9399,N_8339,N_8100);
nand U9400 (N_9400,N_8167,N_7818);
nor U9401 (N_9401,N_7646,N_7442);
and U9402 (N_9402,N_8344,N_8366);
and U9403 (N_9403,N_7703,N_8101);
xnor U9404 (N_9404,N_7279,N_7973);
and U9405 (N_9405,N_7375,N_7362);
and U9406 (N_9406,N_8088,N_8124);
xor U9407 (N_9407,N_8042,N_7372);
xnor U9408 (N_9408,N_7268,N_7624);
and U9409 (N_9409,N_7833,N_7445);
nor U9410 (N_9410,N_8300,N_8249);
nand U9411 (N_9411,N_7418,N_7472);
or U9412 (N_9412,N_7648,N_8057);
nand U9413 (N_9413,N_7644,N_7645);
xor U9414 (N_9414,N_8138,N_7771);
nand U9415 (N_9415,N_8332,N_7304);
nand U9416 (N_9416,N_8034,N_8107);
xnor U9417 (N_9417,N_7410,N_7403);
nor U9418 (N_9418,N_7387,N_8032);
nor U9419 (N_9419,N_7240,N_7220);
xor U9420 (N_9420,N_7914,N_7398);
nor U9421 (N_9421,N_8098,N_8256);
xnor U9422 (N_9422,N_7886,N_7685);
nor U9423 (N_9423,N_7499,N_7819);
and U9424 (N_9424,N_8203,N_7253);
or U9425 (N_9425,N_8397,N_7606);
xor U9426 (N_9426,N_7655,N_7443);
xnor U9427 (N_9427,N_8381,N_7968);
nor U9428 (N_9428,N_8300,N_7296);
or U9429 (N_9429,N_7481,N_7564);
xnor U9430 (N_9430,N_7410,N_7416);
xnor U9431 (N_9431,N_7759,N_7960);
or U9432 (N_9432,N_7631,N_7747);
nand U9433 (N_9433,N_8062,N_8149);
nand U9434 (N_9434,N_8027,N_7239);
or U9435 (N_9435,N_7245,N_7202);
and U9436 (N_9436,N_7979,N_8184);
nor U9437 (N_9437,N_7880,N_8106);
xnor U9438 (N_9438,N_8327,N_7638);
or U9439 (N_9439,N_7458,N_7615);
and U9440 (N_9440,N_8274,N_7837);
and U9441 (N_9441,N_7766,N_7600);
nor U9442 (N_9442,N_7729,N_7396);
or U9443 (N_9443,N_8307,N_8208);
and U9444 (N_9444,N_8072,N_7594);
nor U9445 (N_9445,N_7424,N_7990);
xor U9446 (N_9446,N_7378,N_7819);
xor U9447 (N_9447,N_7898,N_7888);
or U9448 (N_9448,N_7615,N_7611);
xnor U9449 (N_9449,N_8077,N_7577);
xor U9450 (N_9450,N_7296,N_7846);
or U9451 (N_9451,N_7517,N_7598);
xor U9452 (N_9452,N_7288,N_8129);
xor U9453 (N_9453,N_8129,N_8368);
or U9454 (N_9454,N_7346,N_8268);
nor U9455 (N_9455,N_8190,N_7299);
or U9456 (N_9456,N_7273,N_8186);
nor U9457 (N_9457,N_7467,N_8253);
or U9458 (N_9458,N_7755,N_7340);
and U9459 (N_9459,N_8372,N_7830);
and U9460 (N_9460,N_8121,N_7856);
or U9461 (N_9461,N_7901,N_7933);
xor U9462 (N_9462,N_8221,N_7292);
xor U9463 (N_9463,N_7810,N_7713);
and U9464 (N_9464,N_8187,N_7310);
and U9465 (N_9465,N_8283,N_8009);
or U9466 (N_9466,N_7490,N_7409);
xor U9467 (N_9467,N_8274,N_8100);
or U9468 (N_9468,N_7212,N_7898);
nor U9469 (N_9469,N_8238,N_8038);
and U9470 (N_9470,N_7667,N_7872);
or U9471 (N_9471,N_8193,N_7268);
xor U9472 (N_9472,N_7433,N_7766);
nor U9473 (N_9473,N_7500,N_8349);
and U9474 (N_9474,N_7394,N_7741);
xnor U9475 (N_9475,N_8366,N_8364);
and U9476 (N_9476,N_7816,N_7340);
and U9477 (N_9477,N_8319,N_8119);
nand U9478 (N_9478,N_7947,N_7644);
or U9479 (N_9479,N_7313,N_7743);
or U9480 (N_9480,N_8327,N_8236);
or U9481 (N_9481,N_8358,N_8148);
or U9482 (N_9482,N_8295,N_8171);
nor U9483 (N_9483,N_8346,N_7766);
or U9484 (N_9484,N_8037,N_7483);
or U9485 (N_9485,N_8045,N_7836);
nor U9486 (N_9486,N_8274,N_7229);
and U9487 (N_9487,N_7272,N_8097);
or U9488 (N_9488,N_7348,N_7455);
nand U9489 (N_9489,N_7931,N_7590);
nand U9490 (N_9490,N_7846,N_7350);
or U9491 (N_9491,N_7208,N_7650);
nand U9492 (N_9492,N_7500,N_8169);
nand U9493 (N_9493,N_8111,N_7758);
or U9494 (N_9494,N_7986,N_8258);
and U9495 (N_9495,N_7939,N_7750);
or U9496 (N_9496,N_8290,N_7242);
and U9497 (N_9497,N_7269,N_7732);
xnor U9498 (N_9498,N_7242,N_7342);
and U9499 (N_9499,N_7403,N_7977);
xor U9500 (N_9500,N_7493,N_8092);
xor U9501 (N_9501,N_7887,N_7722);
and U9502 (N_9502,N_8239,N_8124);
or U9503 (N_9503,N_7812,N_7392);
and U9504 (N_9504,N_7879,N_8181);
and U9505 (N_9505,N_7957,N_7419);
nor U9506 (N_9506,N_8154,N_7449);
nor U9507 (N_9507,N_8341,N_8296);
xor U9508 (N_9508,N_7478,N_8040);
nor U9509 (N_9509,N_8346,N_7452);
or U9510 (N_9510,N_7743,N_7573);
xor U9511 (N_9511,N_8145,N_7343);
nor U9512 (N_9512,N_8153,N_8382);
nor U9513 (N_9513,N_8281,N_8251);
or U9514 (N_9514,N_7520,N_7513);
and U9515 (N_9515,N_8393,N_7968);
xnor U9516 (N_9516,N_7517,N_7859);
or U9517 (N_9517,N_8133,N_8080);
and U9518 (N_9518,N_7763,N_7543);
or U9519 (N_9519,N_7855,N_7548);
xnor U9520 (N_9520,N_7934,N_7932);
nor U9521 (N_9521,N_8297,N_7238);
and U9522 (N_9522,N_8096,N_7597);
xor U9523 (N_9523,N_8148,N_7626);
xnor U9524 (N_9524,N_7996,N_7471);
nand U9525 (N_9525,N_7615,N_7440);
or U9526 (N_9526,N_8043,N_8243);
or U9527 (N_9527,N_7625,N_8209);
or U9528 (N_9528,N_7988,N_7447);
and U9529 (N_9529,N_7215,N_7684);
xor U9530 (N_9530,N_7719,N_7400);
and U9531 (N_9531,N_7654,N_7828);
nor U9532 (N_9532,N_7392,N_7279);
and U9533 (N_9533,N_7585,N_7857);
or U9534 (N_9534,N_7882,N_7874);
xor U9535 (N_9535,N_7240,N_7717);
or U9536 (N_9536,N_7772,N_7320);
xor U9537 (N_9537,N_8253,N_7938);
and U9538 (N_9538,N_7399,N_8384);
nand U9539 (N_9539,N_8294,N_8168);
or U9540 (N_9540,N_8304,N_7997);
or U9541 (N_9541,N_7327,N_7969);
and U9542 (N_9542,N_8332,N_7341);
nand U9543 (N_9543,N_8020,N_7670);
nand U9544 (N_9544,N_8162,N_8158);
and U9545 (N_9545,N_7769,N_7286);
or U9546 (N_9546,N_7618,N_8079);
nor U9547 (N_9547,N_7224,N_7825);
nand U9548 (N_9548,N_7904,N_7873);
nand U9549 (N_9549,N_7516,N_8367);
or U9550 (N_9550,N_7636,N_8018);
nand U9551 (N_9551,N_8099,N_7208);
nand U9552 (N_9552,N_8102,N_7848);
or U9553 (N_9553,N_8181,N_8324);
nand U9554 (N_9554,N_8298,N_8387);
and U9555 (N_9555,N_7891,N_8187);
or U9556 (N_9556,N_7972,N_7837);
and U9557 (N_9557,N_7783,N_7950);
xnor U9558 (N_9558,N_7389,N_7473);
and U9559 (N_9559,N_7308,N_8167);
xnor U9560 (N_9560,N_8104,N_8106);
xor U9561 (N_9561,N_8343,N_7270);
or U9562 (N_9562,N_7575,N_7329);
or U9563 (N_9563,N_7320,N_7994);
or U9564 (N_9564,N_8268,N_7466);
xor U9565 (N_9565,N_8081,N_7908);
or U9566 (N_9566,N_7506,N_7402);
nor U9567 (N_9567,N_8338,N_7951);
nand U9568 (N_9568,N_8007,N_8356);
or U9569 (N_9569,N_7899,N_8399);
nor U9570 (N_9570,N_7383,N_7693);
and U9571 (N_9571,N_7561,N_7997);
and U9572 (N_9572,N_8091,N_7306);
nor U9573 (N_9573,N_7282,N_7463);
and U9574 (N_9574,N_7536,N_7776);
or U9575 (N_9575,N_7500,N_7470);
nor U9576 (N_9576,N_8164,N_8162);
and U9577 (N_9577,N_7259,N_7707);
and U9578 (N_9578,N_8195,N_8222);
xor U9579 (N_9579,N_7848,N_8063);
or U9580 (N_9580,N_8296,N_7811);
nand U9581 (N_9581,N_8032,N_8163);
nand U9582 (N_9582,N_7533,N_7366);
xnor U9583 (N_9583,N_7486,N_8153);
xor U9584 (N_9584,N_7367,N_8188);
nand U9585 (N_9585,N_7558,N_8366);
and U9586 (N_9586,N_7388,N_8005);
and U9587 (N_9587,N_8026,N_7480);
or U9588 (N_9588,N_8013,N_7421);
nor U9589 (N_9589,N_8178,N_7702);
nor U9590 (N_9590,N_7597,N_8193);
or U9591 (N_9591,N_8119,N_7888);
xnor U9592 (N_9592,N_8069,N_7751);
or U9593 (N_9593,N_7494,N_7211);
xnor U9594 (N_9594,N_7431,N_7263);
nand U9595 (N_9595,N_8172,N_8310);
and U9596 (N_9596,N_7676,N_7493);
xor U9597 (N_9597,N_7903,N_7502);
and U9598 (N_9598,N_7510,N_8344);
nor U9599 (N_9599,N_7536,N_7689);
nor U9600 (N_9600,N_9251,N_8864);
and U9601 (N_9601,N_9390,N_8709);
or U9602 (N_9602,N_8693,N_8429);
xnor U9603 (N_9603,N_9269,N_9425);
xnor U9604 (N_9604,N_9054,N_9300);
xor U9605 (N_9605,N_9457,N_8951);
and U9606 (N_9606,N_8866,N_9452);
nand U9607 (N_9607,N_9286,N_8569);
nor U9608 (N_9608,N_9540,N_8753);
nand U9609 (N_9609,N_8938,N_8687);
nor U9610 (N_9610,N_8677,N_9239);
nor U9611 (N_9611,N_9258,N_9315);
xor U9612 (N_9612,N_8720,N_9422);
nor U9613 (N_9613,N_9584,N_8426);
or U9614 (N_9614,N_8921,N_8831);
and U9615 (N_9615,N_9108,N_8556);
xor U9616 (N_9616,N_9526,N_8694);
nand U9617 (N_9617,N_9417,N_9219);
and U9618 (N_9618,N_9277,N_9332);
nand U9619 (N_9619,N_8881,N_9103);
xnor U9620 (N_9620,N_9552,N_9056);
xnor U9621 (N_9621,N_8472,N_8581);
nand U9622 (N_9622,N_8447,N_8719);
nor U9623 (N_9623,N_8629,N_9205);
xor U9624 (N_9624,N_8946,N_8628);
or U9625 (N_9625,N_9194,N_8800);
or U9626 (N_9626,N_8684,N_9026);
nand U9627 (N_9627,N_8967,N_9267);
nand U9628 (N_9628,N_9558,N_9327);
and U9629 (N_9629,N_8869,N_8760);
nand U9630 (N_9630,N_8832,N_9066);
and U9631 (N_9631,N_9131,N_9582);
or U9632 (N_9632,N_8660,N_9069);
or U9633 (N_9633,N_9431,N_9491);
nor U9634 (N_9634,N_8873,N_9099);
and U9635 (N_9635,N_8579,N_9241);
nand U9636 (N_9636,N_9084,N_8773);
xor U9637 (N_9637,N_8667,N_9232);
and U9638 (N_9638,N_8476,N_9037);
xor U9639 (N_9639,N_9151,N_8735);
nor U9640 (N_9640,N_8595,N_8925);
or U9641 (N_9641,N_8699,N_8602);
nand U9642 (N_9642,N_8932,N_8734);
nor U9643 (N_9643,N_9342,N_9039);
nand U9644 (N_9644,N_9599,N_8910);
and U9645 (N_9645,N_9091,N_9531);
or U9646 (N_9646,N_9093,N_8902);
nor U9647 (N_9647,N_8570,N_8485);
nor U9648 (N_9648,N_8664,N_8525);
and U9649 (N_9649,N_9588,N_9271);
and U9650 (N_9650,N_8814,N_9578);
and U9651 (N_9651,N_9489,N_9338);
and U9652 (N_9652,N_8897,N_9587);
or U9653 (N_9653,N_8473,N_8515);
xnor U9654 (N_9654,N_8441,N_9055);
or U9655 (N_9655,N_9575,N_8909);
or U9656 (N_9656,N_8911,N_8731);
nor U9657 (N_9657,N_8463,N_8846);
nand U9658 (N_9658,N_9141,N_8914);
nor U9659 (N_9659,N_9238,N_9522);
or U9660 (N_9660,N_8712,N_9569);
and U9661 (N_9661,N_9157,N_9061);
xnor U9662 (N_9662,N_9573,N_9553);
and U9663 (N_9663,N_9323,N_8481);
or U9664 (N_9664,N_9303,N_9406);
nor U9665 (N_9665,N_8789,N_9351);
nor U9666 (N_9666,N_9427,N_8450);
and U9667 (N_9667,N_8561,N_9207);
nand U9668 (N_9668,N_9101,N_8844);
nand U9669 (N_9669,N_8875,N_9216);
nor U9670 (N_9670,N_8609,N_8793);
nor U9671 (N_9671,N_9096,N_8772);
xor U9672 (N_9672,N_8400,N_9571);
or U9673 (N_9673,N_9272,N_9397);
nand U9674 (N_9674,N_8586,N_9020);
nor U9675 (N_9675,N_9339,N_8531);
nand U9676 (N_9676,N_8536,N_9304);
xor U9677 (N_9677,N_8498,N_9004);
and U9678 (N_9678,N_8821,N_8607);
nand U9679 (N_9679,N_8795,N_9191);
nand U9680 (N_9680,N_9159,N_9509);
nor U9681 (N_9681,N_8484,N_9033);
nand U9682 (N_9682,N_9126,N_9129);
nor U9683 (N_9683,N_9329,N_9268);
or U9684 (N_9684,N_9192,N_9291);
nand U9685 (N_9685,N_8491,N_9376);
nand U9686 (N_9686,N_9551,N_8888);
and U9687 (N_9687,N_9403,N_9280);
and U9688 (N_9688,N_9174,N_9477);
and U9689 (N_9689,N_9369,N_8565);
or U9690 (N_9690,N_9316,N_9492);
nor U9691 (N_9691,N_9243,N_8679);
or U9692 (N_9692,N_8868,N_9279);
nor U9693 (N_9693,N_9097,N_8547);
nand U9694 (N_9694,N_9209,N_8992);
xor U9695 (N_9695,N_8872,N_8931);
xor U9696 (N_9696,N_8986,N_9325);
xnor U9697 (N_9697,N_8615,N_9168);
xnor U9698 (N_9698,N_9331,N_9005);
and U9699 (N_9699,N_9254,N_8727);
nor U9700 (N_9700,N_9319,N_9444);
or U9701 (N_9701,N_8907,N_9210);
nor U9702 (N_9702,N_8748,N_9125);
nand U9703 (N_9703,N_8955,N_9206);
nor U9704 (N_9704,N_8776,N_8895);
and U9705 (N_9705,N_8906,N_9434);
xnor U9706 (N_9706,N_9568,N_8940);
nand U9707 (N_9707,N_9514,N_8446);
or U9708 (N_9708,N_8436,N_8893);
nand U9709 (N_9709,N_9443,N_8454);
nor U9710 (N_9710,N_9340,N_8923);
xor U9711 (N_9711,N_9029,N_9428);
nor U9712 (N_9712,N_9357,N_8867);
or U9713 (N_9713,N_9440,N_8424);
or U9714 (N_9714,N_8670,N_9423);
or U9715 (N_9715,N_8422,N_8920);
nor U9716 (N_9716,N_9415,N_8585);
nor U9717 (N_9717,N_9077,N_9214);
nor U9718 (N_9718,N_9312,N_9455);
nand U9719 (N_9719,N_9062,N_8972);
nor U9720 (N_9720,N_8427,N_9374);
nand U9721 (N_9721,N_8702,N_9226);
nor U9722 (N_9722,N_9519,N_8738);
and U9723 (N_9723,N_9118,N_9565);
or U9724 (N_9724,N_8824,N_9336);
nor U9725 (N_9725,N_9405,N_9202);
nor U9726 (N_9726,N_9358,N_8656);
xnor U9727 (N_9727,N_8415,N_8421);
nor U9728 (N_9728,N_9309,N_8445);
or U9729 (N_9729,N_9187,N_9515);
or U9730 (N_9730,N_8448,N_8611);
nor U9731 (N_9731,N_8850,N_8665);
nand U9732 (N_9732,N_8730,N_8936);
and U9733 (N_9733,N_9524,N_8983);
or U9734 (N_9734,N_9433,N_8590);
nand U9735 (N_9735,N_9438,N_8937);
nand U9736 (N_9736,N_8577,N_8815);
and U9737 (N_9737,N_9314,N_9408);
xnor U9738 (N_9738,N_9242,N_9111);
or U9739 (N_9739,N_8811,N_9507);
xor U9740 (N_9740,N_8823,N_8542);
nand U9741 (N_9741,N_9143,N_8499);
nand U9742 (N_9742,N_8775,N_9577);
nand U9743 (N_9743,N_8874,N_9188);
and U9744 (N_9744,N_8971,N_8430);
xnor U9745 (N_9745,N_8588,N_9548);
nand U9746 (N_9746,N_9467,N_9412);
and U9747 (N_9747,N_9490,N_8742);
or U9748 (N_9748,N_8620,N_8442);
and U9749 (N_9749,N_8407,N_8903);
nand U9750 (N_9750,N_8507,N_8904);
or U9751 (N_9751,N_8543,N_9453);
or U9752 (N_9752,N_9025,N_8682);
nor U9753 (N_9753,N_9046,N_9088);
nand U9754 (N_9754,N_8489,N_8519);
xor U9755 (N_9755,N_9296,N_9245);
and U9756 (N_9756,N_8870,N_8638);
or U9757 (N_9757,N_8444,N_9119);
xor U9758 (N_9758,N_9154,N_8761);
or U9759 (N_9759,N_8653,N_9016);
nor U9760 (N_9760,N_8732,N_8750);
xor U9761 (N_9761,N_8996,N_8822);
nor U9762 (N_9762,N_8482,N_9089);
and U9763 (N_9763,N_8642,N_8845);
and U9764 (N_9764,N_9110,N_8755);
xor U9765 (N_9765,N_8621,N_9354);
or U9766 (N_9766,N_8458,N_8554);
xnor U9767 (N_9767,N_9419,N_8518);
nand U9768 (N_9768,N_8879,N_8568);
and U9769 (N_9769,N_8973,N_8840);
nand U9770 (N_9770,N_9495,N_8855);
nand U9771 (N_9771,N_9021,N_8401);
and U9772 (N_9772,N_9169,N_9480);
nand U9773 (N_9773,N_8540,N_8630);
nor U9774 (N_9774,N_8544,N_8759);
xor U9775 (N_9775,N_9372,N_8828);
nor U9776 (N_9776,N_9451,N_9344);
nand U9777 (N_9777,N_8898,N_9448);
nand U9778 (N_9778,N_8504,N_8598);
nor U9779 (N_9779,N_9474,N_8715);
and U9780 (N_9780,N_9090,N_8859);
or U9781 (N_9781,N_9442,N_8471);
nand U9782 (N_9782,N_8534,N_9416);
or U9783 (N_9783,N_8856,N_8989);
xnor U9784 (N_9784,N_8501,N_9098);
nand U9785 (N_9785,N_8756,N_8758);
nand U9786 (N_9786,N_9167,N_8669);
nor U9787 (N_9787,N_9537,N_9107);
or U9788 (N_9788,N_8635,N_9060);
nand U9789 (N_9789,N_8927,N_8562);
or U9790 (N_9790,N_8640,N_8995);
xnor U9791 (N_9791,N_9175,N_8580);
nor U9792 (N_9792,N_9384,N_9359);
or U9793 (N_9793,N_8456,N_9043);
or U9794 (N_9794,N_9032,N_9469);
nor U9795 (N_9795,N_9171,N_9117);
or U9796 (N_9796,N_8509,N_9550);
or U9797 (N_9797,N_9484,N_9064);
or U9798 (N_9798,N_9385,N_8626);
nand U9799 (N_9799,N_8794,N_8647);
and U9800 (N_9800,N_8985,N_9011);
nor U9801 (N_9801,N_9536,N_9498);
or U9802 (N_9802,N_9213,N_9204);
xor U9803 (N_9803,N_9549,N_8479);
xnor U9804 (N_9804,N_9186,N_9105);
nor U9805 (N_9805,N_8505,N_8560);
or U9806 (N_9806,N_9500,N_8807);
xnor U9807 (N_9807,N_9545,N_8691);
and U9808 (N_9808,N_8686,N_9306);
or U9809 (N_9809,N_9473,N_8723);
and U9810 (N_9810,N_8467,N_8412);
or U9811 (N_9811,N_8941,N_8876);
nand U9812 (N_9812,N_9466,N_9045);
or U9813 (N_9813,N_9356,N_9476);
or U9814 (N_9814,N_9247,N_8877);
xnor U9815 (N_9815,N_8468,N_8490);
or U9816 (N_9816,N_8729,N_8537);
nor U9817 (N_9817,N_9301,N_9257);
nand U9818 (N_9818,N_9420,N_8673);
or U9819 (N_9819,N_9225,N_9445);
or U9820 (N_9820,N_9389,N_9532);
xnor U9821 (N_9821,N_8680,N_9123);
xor U9822 (N_9822,N_9127,N_8563);
nand U9823 (N_9823,N_8644,N_8710);
or U9824 (N_9824,N_9023,N_9160);
xnor U9825 (N_9825,N_8606,N_9598);
nor U9826 (N_9826,N_8497,N_9449);
and U9827 (N_9827,N_9156,N_9377);
nor U9828 (N_9828,N_9246,N_9149);
nor U9829 (N_9829,N_9006,N_9557);
or U9830 (N_9830,N_8721,N_9485);
and U9831 (N_9831,N_9176,N_8934);
nor U9832 (N_9832,N_8403,N_8405);
or U9833 (N_9833,N_8672,N_8964);
xnor U9834 (N_9834,N_9145,N_9305);
and U9835 (N_9835,N_9392,N_8784);
and U9836 (N_9836,N_9590,N_8698);
and U9837 (N_9837,N_8806,N_8849);
or U9838 (N_9838,N_9220,N_8500);
nand U9839 (N_9839,N_8455,N_9136);
nand U9840 (N_9840,N_9177,N_8961);
nor U9841 (N_9841,N_9018,N_8880);
nor U9842 (N_9842,N_9413,N_9285);
nor U9843 (N_9843,N_8413,N_9193);
nor U9844 (N_9844,N_9065,N_9297);
nand U9845 (N_9845,N_8474,N_9439);
and U9846 (N_9846,N_9533,N_8438);
nand U9847 (N_9847,N_9530,N_9087);
xor U9848 (N_9848,N_9041,N_8551);
xnor U9849 (N_9849,N_8763,N_8997);
xnor U9850 (N_9850,N_8970,N_8512);
and U9851 (N_9851,N_9075,N_9402);
xor U9852 (N_9852,N_9040,N_9290);
nor U9853 (N_9853,N_8648,N_9208);
xnor U9854 (N_9854,N_9404,N_8549);
xor U9855 (N_9855,N_9252,N_8969);
nor U9856 (N_9856,N_8706,N_9592);
nand U9857 (N_9857,N_8674,N_9346);
xor U9858 (N_9858,N_8417,N_9371);
nand U9859 (N_9859,N_8817,N_8496);
nand U9860 (N_9860,N_9382,N_8954);
or U9861 (N_9861,N_8963,N_9106);
nor U9862 (N_9862,N_9036,N_8521);
nor U9863 (N_9863,N_9527,N_8882);
xor U9864 (N_9864,N_8764,N_9398);
and U9865 (N_9865,N_8567,N_8788);
nand U9866 (N_9866,N_8952,N_9094);
nand U9867 (N_9867,N_9487,N_9414);
nor U9868 (N_9868,N_8619,N_8947);
and U9869 (N_9869,N_8825,N_9203);
nor U9870 (N_9870,N_8975,N_9014);
or U9871 (N_9871,N_9463,N_9418);
and U9872 (N_9872,N_8812,N_9222);
nor U9873 (N_9873,N_9361,N_9072);
xor U9874 (N_9874,N_8885,N_8862);
nor U9875 (N_9875,N_9158,N_9295);
nor U9876 (N_9876,N_8443,N_8462);
and U9877 (N_9877,N_9421,N_9499);
or U9878 (N_9878,N_8836,N_8651);
and U9879 (N_9879,N_9092,N_9435);
and U9880 (N_9880,N_9504,N_8717);
or U9881 (N_9881,N_9053,N_9512);
nor U9882 (N_9882,N_9560,N_9050);
nand U9883 (N_9883,N_9049,N_9589);
and U9884 (N_9884,N_8613,N_8797);
and U9885 (N_9885,N_8899,N_8538);
or U9886 (N_9886,N_9270,N_8886);
or U9887 (N_9887,N_9283,N_9529);
nor U9888 (N_9888,N_9585,N_9259);
and U9889 (N_9889,N_9528,N_9482);
nand U9890 (N_9890,N_9429,N_8922);
or U9891 (N_9891,N_9027,N_8622);
nor U9892 (N_9892,N_9199,N_9395);
xnor U9893 (N_9893,N_8614,N_9113);
or U9894 (N_9894,N_8792,N_9124);
nand U9895 (N_9895,N_9458,N_8546);
and U9896 (N_9896,N_9535,N_8503);
nor U9897 (N_9897,N_9579,N_8819);
or U9898 (N_9898,N_9261,N_9566);
xnor U9899 (N_9899,N_8639,N_8736);
xor U9900 (N_9900,N_9365,N_8529);
nand U9901 (N_9901,N_9135,N_9211);
and U9902 (N_9902,N_9031,N_9424);
nand U9903 (N_9903,N_9063,N_8889);
nand U9904 (N_9904,N_9388,N_8786);
or U9905 (N_9905,N_8782,N_9275);
nor U9906 (N_9906,N_8998,N_9262);
and U9907 (N_9907,N_9355,N_9462);
xnor U9908 (N_9908,N_8659,N_8668);
nor U9909 (N_9909,N_8790,N_9068);
and U9910 (N_9910,N_8843,N_8692);
nor U9911 (N_9911,N_9003,N_8661);
xor U9912 (N_9912,N_9081,N_8666);
nor U9913 (N_9913,N_9007,N_9047);
nor U9914 (N_9914,N_8704,N_8420);
or U9915 (N_9915,N_8558,N_9576);
nand U9916 (N_9916,N_9539,N_8863);
xor U9917 (N_9917,N_9460,N_8655);
nand U9918 (N_9918,N_9360,N_9182);
xnor U9919 (N_9919,N_9180,N_8744);
or U9920 (N_9920,N_8978,N_8924);
nor U9921 (N_9921,N_9237,N_9379);
and U9922 (N_9922,N_9024,N_8528);
or U9923 (N_9923,N_9364,N_8584);
xor U9924 (N_9924,N_8627,N_8591);
nor U9925 (N_9925,N_8722,N_8587);
nand U9926 (N_9926,N_8487,N_9461);
and U9927 (N_9927,N_8728,N_8652);
xor U9928 (N_9928,N_9274,N_9085);
and U9929 (N_9929,N_8958,N_9030);
xnor U9930 (N_9930,N_8631,N_9562);
xnor U9931 (N_9931,N_8475,N_8557);
nor U9932 (N_9932,N_9133,N_9001);
nor U9933 (N_9933,N_8548,N_9185);
or U9934 (N_9934,N_8460,N_8532);
nor U9935 (N_9935,N_9475,N_8962);
nor U9936 (N_9936,N_8459,N_9307);
and U9937 (N_9937,N_9278,N_8827);
or U9938 (N_9938,N_8766,N_9407);
xor U9939 (N_9939,N_8469,N_8774);
or U9940 (N_9940,N_8610,N_8926);
xor U9941 (N_9941,N_9153,N_8625);
xor U9942 (N_9942,N_8726,N_9196);
nand U9943 (N_9943,N_9244,N_9010);
nand U9944 (N_9944,N_9543,N_8894);
xor U9945 (N_9945,N_8517,N_9074);
or U9946 (N_9946,N_9249,N_9446);
nand U9947 (N_9947,N_8948,N_8566);
and U9948 (N_9948,N_9464,N_8928);
or U9949 (N_9949,N_8861,N_8516);
or U9950 (N_9950,N_9481,N_9038);
or U9951 (N_9951,N_8833,N_9100);
nor U9952 (N_9952,N_9264,N_9044);
xnor U9953 (N_9953,N_8596,N_9015);
nand U9954 (N_9954,N_8705,N_8678);
nand U9955 (N_9955,N_8857,N_9510);
and U9956 (N_9956,N_9368,N_9596);
xor U9957 (N_9957,N_9200,N_8432);
or U9958 (N_9958,N_9282,N_9478);
and U9959 (N_9959,N_9459,N_9541);
or U9960 (N_9960,N_9104,N_8908);
xor U9961 (N_9961,N_9236,N_9181);
xor U9962 (N_9962,N_9265,N_8887);
nor U9963 (N_9963,N_9276,N_9559);
nor U9964 (N_9964,N_8465,N_8977);
xnor U9965 (N_9965,N_8520,N_8939);
or U9966 (N_9966,N_9542,N_8841);
nand U9967 (N_9967,N_8645,N_8739);
or U9968 (N_9968,N_9013,N_8681);
nor U9969 (N_9969,N_8419,N_8466);
nor U9970 (N_9970,N_8478,N_8690);
and U9971 (N_9971,N_9470,N_8771);
xnor U9972 (N_9972,N_8535,N_8539);
nand U9973 (N_9973,N_8810,N_8754);
and U9974 (N_9974,N_8671,N_8999);
or U9975 (N_9975,N_8829,N_8740);
or U9976 (N_9976,N_8935,N_9289);
or U9977 (N_9977,N_9447,N_8725);
xnor U9978 (N_9978,N_8891,N_8574);
nand U9979 (N_9979,N_8993,N_8597);
nand U9980 (N_9980,N_8960,N_8530);
and U9981 (N_9981,N_8650,N_8787);
and U9982 (N_9982,N_8675,N_9324);
nor U9983 (N_9983,N_9255,N_9347);
and U9984 (N_9984,N_8494,N_9353);
nor U9985 (N_9985,N_8733,N_8433);
nand U9986 (N_9986,N_8848,N_9224);
xnor U9987 (N_9987,N_8718,N_8777);
xor U9988 (N_9988,N_9130,N_9139);
nor U9989 (N_9989,N_8506,N_8492);
nor U9990 (N_9990,N_8979,N_8933);
nor U9991 (N_9991,N_9217,N_9563);
and U9992 (N_9992,N_8514,N_8765);
or U9993 (N_9993,N_9394,N_8747);
and U9994 (N_9994,N_9165,N_9002);
nor U9995 (N_9995,N_9233,N_8968);
nor U9996 (N_9996,N_9580,N_9586);
nor U9997 (N_9997,N_9116,N_8646);
xor U9998 (N_9998,N_8510,N_9378);
nand U9999 (N_9999,N_8953,N_8987);
xor U10000 (N_10000,N_9138,N_9163);
and U10001 (N_10001,N_8480,N_9076);
xor U10002 (N_10002,N_9366,N_8988);
nor U10003 (N_10003,N_8858,N_8526);
nor U10004 (N_10004,N_8663,N_8641);
xnor U10005 (N_10005,N_8594,N_9362);
xnor U10006 (N_10006,N_8428,N_8745);
or U10007 (N_10007,N_9052,N_8633);
nand U10008 (N_10008,N_9581,N_8802);
or U10009 (N_10009,N_8545,N_8783);
nor U10010 (N_10010,N_9253,N_8527);
nand U10011 (N_10011,N_9000,N_9070);
and U10012 (N_10012,N_9538,N_8483);
nor U10013 (N_10013,N_8418,N_8896);
and U10014 (N_10014,N_8623,N_8573);
xnor U10015 (N_10015,N_8683,N_8796);
or U10016 (N_10016,N_9079,N_9380);
nand U10017 (N_10017,N_9173,N_9078);
and U10018 (N_10018,N_9493,N_9393);
nor U10019 (N_10019,N_8883,N_9082);
and U10020 (N_10020,N_9299,N_8860);
nor U10021 (N_10021,N_9334,N_8779);
nand U10022 (N_10022,N_8617,N_8878);
nor U10023 (N_10023,N_8402,N_8950);
or U10024 (N_10024,N_9521,N_9067);
or U10025 (N_10025,N_9441,N_9383);
or U10026 (N_10026,N_9308,N_9561);
or U10027 (N_10027,N_8818,N_9137);
and U10028 (N_10028,N_9273,N_9333);
or U10029 (N_10029,N_8976,N_8834);
and U10030 (N_10030,N_9396,N_9172);
nand U10031 (N_10031,N_8711,N_8576);
and U10032 (N_10032,N_9281,N_9335);
or U10033 (N_10033,N_9349,N_8716);
nor U10034 (N_10034,N_9326,N_8533);
xnor U10035 (N_10035,N_9518,N_9432);
nor U10036 (N_10036,N_8847,N_9343);
xor U10037 (N_10037,N_9227,N_9472);
nor U10038 (N_10038,N_8612,N_9468);
nor U10039 (N_10039,N_9574,N_9221);
and U10040 (N_10040,N_8578,N_9302);
or U10041 (N_10041,N_8695,N_9164);
nand U10042 (N_10042,N_9230,N_8404);
nor U10043 (N_10043,N_8541,N_8616);
nand U10044 (N_10044,N_8632,N_9363);
xor U10045 (N_10045,N_8599,N_8945);
and U10046 (N_10046,N_8842,N_9086);
and U10047 (N_10047,N_9162,N_9328);
nor U10048 (N_10048,N_8464,N_9311);
and U10049 (N_10049,N_8416,N_9109);
and U10050 (N_10050,N_9148,N_8768);
or U10051 (N_10051,N_9313,N_8749);
or U10052 (N_10052,N_9042,N_9450);
and U10053 (N_10053,N_8780,N_8701);
nand U10054 (N_10054,N_9572,N_9348);
nand U10055 (N_10055,N_9583,N_8743);
xnor U10056 (N_10056,N_8658,N_8502);
or U10057 (N_10057,N_8707,N_9057);
and U10058 (N_10058,N_8488,N_9028);
or U10059 (N_10059,N_9525,N_8991);
nor U10060 (N_10060,N_8552,N_8820);
xnor U10061 (N_10061,N_9497,N_9112);
nand U10062 (N_10062,N_9375,N_8685);
and U10063 (N_10063,N_9352,N_8486);
and U10064 (N_10064,N_9494,N_8980);
or U10065 (N_10065,N_8522,N_9502);
or U10066 (N_10066,N_9409,N_9410);
nand U10067 (N_10067,N_9330,N_9523);
xnor U10068 (N_10068,N_9411,N_9229);
nor U10069 (N_10069,N_8643,N_9150);
or U10070 (N_10070,N_8511,N_8957);
nand U10071 (N_10071,N_8916,N_9059);
xnor U10072 (N_10072,N_8762,N_8959);
nor U10073 (N_10073,N_8697,N_8837);
nor U10074 (N_10074,N_8423,N_9310);
and U10075 (N_10075,N_8634,N_8930);
or U10076 (N_10076,N_8994,N_8654);
and U10077 (N_10077,N_8593,N_8984);
xnor U10078 (N_10078,N_9367,N_9190);
and U10079 (N_10079,N_8746,N_9546);
or U10080 (N_10080,N_8564,N_9430);
nand U10081 (N_10081,N_9520,N_9544);
xnor U10082 (N_10082,N_8791,N_9240);
and U10083 (N_10083,N_8477,N_9034);
nand U10084 (N_10084,N_9387,N_9386);
or U10085 (N_10085,N_9184,N_8890);
xor U10086 (N_10086,N_8804,N_8406);
or U10087 (N_10087,N_9121,N_9218);
and U10088 (N_10088,N_8461,N_9161);
nor U10089 (N_10089,N_9250,N_9556);
nor U10090 (N_10090,N_8440,N_8410);
xor U10091 (N_10091,N_9293,N_9166);
nor U10092 (N_10092,N_8605,N_9235);
or U10093 (N_10093,N_9051,N_8604);
nand U10094 (N_10094,N_9083,N_8495);
xor U10095 (N_10095,N_9009,N_8688);
nor U10096 (N_10096,N_9426,N_8751);
xnor U10097 (N_10097,N_9593,N_8676);
and U10098 (N_10098,N_8414,N_8965);
nor U10099 (N_10099,N_8425,N_9471);
nor U10100 (N_10100,N_8470,N_9058);
and U10101 (N_10101,N_9212,N_8905);
nand U10102 (N_10102,N_9201,N_9381);
nand U10103 (N_10103,N_8657,N_8919);
or U10104 (N_10104,N_9198,N_9144);
nand U10105 (N_10105,N_8550,N_8785);
xnor U10106 (N_10106,N_8603,N_8917);
xnor U10107 (N_10107,N_9505,N_8838);
nand U10108 (N_10108,N_9197,N_8508);
xor U10109 (N_10109,N_9292,N_8435);
nor U10110 (N_10110,N_9022,N_8411);
xor U10111 (N_10111,N_8452,N_8798);
xor U10112 (N_10112,N_9479,N_9132);
xor U10113 (N_10113,N_9234,N_9183);
nand U10114 (N_10114,N_9400,N_9178);
or U10115 (N_10115,N_8852,N_8408);
nor U10116 (N_10116,N_8805,N_9284);
nor U10117 (N_10117,N_9071,N_8724);
nor U10118 (N_10118,N_9555,N_8813);
xnor U10119 (N_10119,N_9223,N_8457);
and U10120 (N_10120,N_8524,N_9095);
nor U10121 (N_10121,N_9189,N_9288);
nor U10122 (N_10122,N_8708,N_9486);
or U10123 (N_10123,N_9215,N_9122);
or U10124 (N_10124,N_9102,N_8801);
xor U10125 (N_10125,N_9597,N_8409);
nor U10126 (N_10126,N_8649,N_9248);
or U10127 (N_10127,N_8689,N_9564);
and U10128 (N_10128,N_8929,N_8943);
and U10129 (N_10129,N_9437,N_9114);
nand U10130 (N_10130,N_8981,N_8575);
nor U10131 (N_10131,N_8600,N_9322);
xnor U10132 (N_10132,N_9146,N_9080);
nor U10133 (N_10133,N_8799,N_8966);
nor U10134 (N_10134,N_8637,N_9517);
nor U10135 (N_10135,N_8582,N_9341);
and U10136 (N_10136,N_9465,N_9595);
or U10137 (N_10137,N_8892,N_8990);
xnor U10138 (N_10138,N_8572,N_9152);
xor U10139 (N_10139,N_8830,N_8944);
nor U10140 (N_10140,N_8982,N_9155);
nand U10141 (N_10141,N_9513,N_9483);
xnor U10142 (N_10142,N_8592,N_8835);
xor U10143 (N_10143,N_9035,N_9260);
nor U10144 (N_10144,N_8559,N_9228);
and U10145 (N_10145,N_8513,N_9195);
xor U10146 (N_10146,N_9134,N_8781);
and U10147 (N_10147,N_8942,N_9140);
nor U10148 (N_10148,N_8451,N_9506);
or U10149 (N_10149,N_9454,N_8949);
or U10150 (N_10150,N_8839,N_9298);
or U10151 (N_10151,N_9401,N_9456);
and U10152 (N_10152,N_9256,N_8809);
and U10153 (N_10153,N_8871,N_9263);
and U10154 (N_10154,N_9128,N_9516);
nand U10155 (N_10155,N_8913,N_8714);
xor U10156 (N_10156,N_9503,N_8741);
nand U10157 (N_10157,N_8851,N_8912);
or U10158 (N_10158,N_9294,N_9534);
xor U10159 (N_10159,N_8608,N_9337);
or U10160 (N_10160,N_9570,N_8583);
or U10161 (N_10161,N_8778,N_8696);
nand U10162 (N_10162,N_8571,N_8915);
xor U10163 (N_10163,N_8618,N_8808);
xor U10164 (N_10164,N_8854,N_9501);
nor U10165 (N_10165,N_9373,N_8553);
nand U10166 (N_10166,N_8624,N_9488);
nand U10167 (N_10167,N_9170,N_9008);
xor U10168 (N_10168,N_8752,N_9567);
nor U10169 (N_10169,N_8816,N_8431);
xor U10170 (N_10170,N_8493,N_8449);
nor U10171 (N_10171,N_8434,N_8703);
nand U10172 (N_10172,N_8974,N_8662);
nor U10173 (N_10173,N_8453,N_9345);
or U10174 (N_10174,N_9399,N_9142);
or U10175 (N_10175,N_9594,N_9048);
nand U10176 (N_10176,N_9350,N_9147);
nand U10177 (N_10177,N_9436,N_9321);
and U10178 (N_10178,N_9511,N_9115);
or U10179 (N_10179,N_9508,N_8439);
nor U10180 (N_10180,N_8636,N_8601);
xnor U10181 (N_10181,N_9073,N_8767);
nor U10182 (N_10182,N_9370,N_8769);
or U10183 (N_10183,N_9179,N_9496);
xnor U10184 (N_10184,N_8956,N_9317);
and U10185 (N_10185,N_9019,N_9547);
nor U10186 (N_10186,N_8826,N_8803);
or U10187 (N_10187,N_9120,N_8770);
and U10188 (N_10188,N_8589,N_9554);
or U10189 (N_10189,N_9318,N_8918);
nand U10190 (N_10190,N_8865,N_9320);
xnor U10191 (N_10191,N_9266,N_8523);
nand U10192 (N_10192,N_8853,N_8757);
nand U10193 (N_10193,N_8437,N_9391);
or U10194 (N_10194,N_9231,N_9287);
nor U10195 (N_10195,N_8713,N_8884);
and U10196 (N_10196,N_8700,N_8555);
and U10197 (N_10197,N_9012,N_9591);
nand U10198 (N_10198,N_8737,N_8901);
nand U10199 (N_10199,N_9017,N_8900);
xor U10200 (N_10200,N_8930,N_8957);
or U10201 (N_10201,N_9107,N_8658);
xnor U10202 (N_10202,N_8453,N_8423);
or U10203 (N_10203,N_9105,N_9107);
nand U10204 (N_10204,N_8829,N_8617);
and U10205 (N_10205,N_8568,N_8991);
or U10206 (N_10206,N_8911,N_8521);
nor U10207 (N_10207,N_8651,N_8406);
nand U10208 (N_10208,N_8976,N_8941);
nor U10209 (N_10209,N_8739,N_8889);
nand U10210 (N_10210,N_9314,N_8489);
or U10211 (N_10211,N_9321,N_8640);
nor U10212 (N_10212,N_9228,N_9498);
nor U10213 (N_10213,N_8877,N_8690);
and U10214 (N_10214,N_8919,N_8616);
xor U10215 (N_10215,N_9032,N_9382);
nand U10216 (N_10216,N_9009,N_9384);
xnor U10217 (N_10217,N_8563,N_8990);
nor U10218 (N_10218,N_8433,N_9157);
xor U10219 (N_10219,N_8509,N_9520);
or U10220 (N_10220,N_8836,N_8881);
or U10221 (N_10221,N_9319,N_9410);
xnor U10222 (N_10222,N_9213,N_9425);
nor U10223 (N_10223,N_9039,N_9105);
xnor U10224 (N_10224,N_9167,N_8681);
nor U10225 (N_10225,N_8520,N_9056);
nand U10226 (N_10226,N_9345,N_9242);
xor U10227 (N_10227,N_8583,N_9518);
and U10228 (N_10228,N_8710,N_9254);
and U10229 (N_10229,N_9471,N_9268);
xor U10230 (N_10230,N_9167,N_8965);
nand U10231 (N_10231,N_8561,N_9170);
and U10232 (N_10232,N_9139,N_8792);
nand U10233 (N_10233,N_8485,N_8622);
xnor U10234 (N_10234,N_8763,N_8727);
nand U10235 (N_10235,N_8653,N_9380);
xnor U10236 (N_10236,N_8751,N_8718);
and U10237 (N_10237,N_8573,N_9144);
nand U10238 (N_10238,N_8491,N_8473);
xor U10239 (N_10239,N_8675,N_9145);
xor U10240 (N_10240,N_8653,N_9300);
or U10241 (N_10241,N_8855,N_9533);
nand U10242 (N_10242,N_8520,N_8669);
or U10243 (N_10243,N_9026,N_8998);
nand U10244 (N_10244,N_8780,N_9111);
or U10245 (N_10245,N_8502,N_8951);
xor U10246 (N_10246,N_8997,N_9097);
xor U10247 (N_10247,N_9276,N_9339);
xnor U10248 (N_10248,N_8773,N_9059);
and U10249 (N_10249,N_9060,N_9325);
or U10250 (N_10250,N_8736,N_8622);
nor U10251 (N_10251,N_8860,N_8500);
or U10252 (N_10252,N_8413,N_9347);
or U10253 (N_10253,N_9391,N_9026);
xor U10254 (N_10254,N_8803,N_9262);
and U10255 (N_10255,N_8773,N_9175);
and U10256 (N_10256,N_8813,N_9118);
xnor U10257 (N_10257,N_9039,N_9069);
nand U10258 (N_10258,N_9033,N_9589);
nor U10259 (N_10259,N_8877,N_9005);
xnor U10260 (N_10260,N_9454,N_8785);
or U10261 (N_10261,N_8571,N_8450);
nand U10262 (N_10262,N_8519,N_9009);
or U10263 (N_10263,N_9490,N_8743);
nand U10264 (N_10264,N_9043,N_9579);
nor U10265 (N_10265,N_9025,N_9033);
nor U10266 (N_10266,N_9397,N_8982);
nor U10267 (N_10267,N_9344,N_8869);
nand U10268 (N_10268,N_9029,N_9383);
nor U10269 (N_10269,N_8768,N_8937);
xor U10270 (N_10270,N_9491,N_9066);
nand U10271 (N_10271,N_8970,N_8961);
xor U10272 (N_10272,N_8528,N_9553);
nand U10273 (N_10273,N_9342,N_8676);
xor U10274 (N_10274,N_8645,N_8890);
and U10275 (N_10275,N_9275,N_9414);
nand U10276 (N_10276,N_8874,N_8811);
and U10277 (N_10277,N_8506,N_9347);
or U10278 (N_10278,N_8965,N_9484);
and U10279 (N_10279,N_8566,N_8694);
or U10280 (N_10280,N_8928,N_8794);
xnor U10281 (N_10281,N_8610,N_9100);
or U10282 (N_10282,N_8467,N_8458);
or U10283 (N_10283,N_9350,N_8961);
xor U10284 (N_10284,N_9366,N_8659);
xor U10285 (N_10285,N_9590,N_9016);
or U10286 (N_10286,N_8759,N_9243);
or U10287 (N_10287,N_8508,N_8927);
or U10288 (N_10288,N_8604,N_8443);
nor U10289 (N_10289,N_8771,N_8594);
or U10290 (N_10290,N_8847,N_8898);
nand U10291 (N_10291,N_9474,N_8677);
and U10292 (N_10292,N_9178,N_9512);
nand U10293 (N_10293,N_8656,N_8684);
nand U10294 (N_10294,N_8582,N_8792);
xor U10295 (N_10295,N_8594,N_9466);
nor U10296 (N_10296,N_8691,N_8941);
xnor U10297 (N_10297,N_9428,N_8762);
and U10298 (N_10298,N_8933,N_9125);
nand U10299 (N_10299,N_8697,N_8437);
or U10300 (N_10300,N_8925,N_9061);
and U10301 (N_10301,N_9230,N_9476);
and U10302 (N_10302,N_8954,N_9256);
or U10303 (N_10303,N_8794,N_8977);
or U10304 (N_10304,N_9487,N_9180);
nand U10305 (N_10305,N_9181,N_9160);
or U10306 (N_10306,N_9343,N_8638);
nand U10307 (N_10307,N_9282,N_8790);
or U10308 (N_10308,N_9286,N_9373);
xnor U10309 (N_10309,N_8578,N_9543);
xor U10310 (N_10310,N_8410,N_8852);
nor U10311 (N_10311,N_9265,N_8835);
xnor U10312 (N_10312,N_8685,N_8425);
xnor U10313 (N_10313,N_8584,N_9136);
or U10314 (N_10314,N_8567,N_9136);
or U10315 (N_10315,N_8579,N_8917);
xor U10316 (N_10316,N_8829,N_8814);
or U10317 (N_10317,N_9411,N_9572);
and U10318 (N_10318,N_9072,N_8832);
or U10319 (N_10319,N_9458,N_9140);
nand U10320 (N_10320,N_8987,N_8913);
nand U10321 (N_10321,N_9102,N_9134);
and U10322 (N_10322,N_8854,N_9266);
xnor U10323 (N_10323,N_8517,N_9313);
and U10324 (N_10324,N_9120,N_9055);
or U10325 (N_10325,N_8766,N_9405);
nand U10326 (N_10326,N_9031,N_8410);
nor U10327 (N_10327,N_9132,N_8685);
nor U10328 (N_10328,N_8467,N_8614);
or U10329 (N_10329,N_9302,N_8591);
and U10330 (N_10330,N_8616,N_9299);
xnor U10331 (N_10331,N_9026,N_9503);
nand U10332 (N_10332,N_8952,N_8478);
nor U10333 (N_10333,N_9197,N_8656);
xor U10334 (N_10334,N_8543,N_8985);
and U10335 (N_10335,N_8716,N_8478);
xor U10336 (N_10336,N_8831,N_9578);
nand U10337 (N_10337,N_8415,N_8616);
nand U10338 (N_10338,N_9035,N_8963);
and U10339 (N_10339,N_8701,N_8469);
xnor U10340 (N_10340,N_9520,N_8739);
or U10341 (N_10341,N_8426,N_9313);
nand U10342 (N_10342,N_9032,N_8704);
and U10343 (N_10343,N_9372,N_9016);
nand U10344 (N_10344,N_9093,N_8675);
and U10345 (N_10345,N_8616,N_9073);
or U10346 (N_10346,N_8525,N_9178);
nor U10347 (N_10347,N_9247,N_9442);
nor U10348 (N_10348,N_8442,N_9276);
xnor U10349 (N_10349,N_8780,N_8742);
nand U10350 (N_10350,N_8969,N_9061);
or U10351 (N_10351,N_9269,N_8790);
and U10352 (N_10352,N_8819,N_9563);
or U10353 (N_10353,N_8757,N_8558);
and U10354 (N_10354,N_9553,N_9517);
nand U10355 (N_10355,N_9240,N_8754);
nor U10356 (N_10356,N_8645,N_8656);
xnor U10357 (N_10357,N_8969,N_8707);
nand U10358 (N_10358,N_8485,N_8544);
and U10359 (N_10359,N_9086,N_8678);
and U10360 (N_10360,N_9300,N_9308);
or U10361 (N_10361,N_8517,N_8705);
and U10362 (N_10362,N_8625,N_9058);
nor U10363 (N_10363,N_8503,N_8402);
nor U10364 (N_10364,N_9302,N_8603);
nand U10365 (N_10365,N_8768,N_8979);
nand U10366 (N_10366,N_9096,N_8711);
xor U10367 (N_10367,N_8921,N_9259);
xnor U10368 (N_10368,N_8763,N_8410);
xnor U10369 (N_10369,N_8486,N_8445);
nand U10370 (N_10370,N_9511,N_9469);
or U10371 (N_10371,N_8649,N_9312);
and U10372 (N_10372,N_8636,N_9335);
nand U10373 (N_10373,N_8429,N_9246);
xnor U10374 (N_10374,N_8623,N_9533);
and U10375 (N_10375,N_9342,N_9466);
xor U10376 (N_10376,N_8836,N_8704);
xor U10377 (N_10377,N_8645,N_8910);
nand U10378 (N_10378,N_9448,N_8755);
nor U10379 (N_10379,N_8875,N_9561);
nor U10380 (N_10380,N_8772,N_8915);
xor U10381 (N_10381,N_8822,N_9185);
nand U10382 (N_10382,N_8886,N_9171);
and U10383 (N_10383,N_9275,N_8429);
xor U10384 (N_10384,N_9411,N_8942);
nor U10385 (N_10385,N_8719,N_9164);
or U10386 (N_10386,N_9266,N_9325);
nor U10387 (N_10387,N_9298,N_9322);
nand U10388 (N_10388,N_8752,N_9145);
nand U10389 (N_10389,N_9071,N_8767);
nor U10390 (N_10390,N_8499,N_9095);
or U10391 (N_10391,N_9289,N_9159);
nor U10392 (N_10392,N_8822,N_9264);
nand U10393 (N_10393,N_9480,N_9311);
nand U10394 (N_10394,N_9570,N_8958);
nor U10395 (N_10395,N_9500,N_9169);
and U10396 (N_10396,N_8627,N_8559);
nand U10397 (N_10397,N_9513,N_8849);
nand U10398 (N_10398,N_9194,N_8467);
nand U10399 (N_10399,N_8887,N_9188);
xor U10400 (N_10400,N_8531,N_8700);
and U10401 (N_10401,N_8785,N_9540);
nand U10402 (N_10402,N_9312,N_8888);
xor U10403 (N_10403,N_9220,N_8730);
nand U10404 (N_10404,N_8998,N_8533);
xnor U10405 (N_10405,N_8941,N_9206);
or U10406 (N_10406,N_9241,N_8457);
nand U10407 (N_10407,N_8548,N_8471);
and U10408 (N_10408,N_8646,N_9546);
xor U10409 (N_10409,N_8798,N_9570);
nor U10410 (N_10410,N_9347,N_9474);
nand U10411 (N_10411,N_9076,N_9520);
and U10412 (N_10412,N_8592,N_8922);
nand U10413 (N_10413,N_9546,N_9515);
and U10414 (N_10414,N_9460,N_8976);
and U10415 (N_10415,N_9544,N_9234);
nor U10416 (N_10416,N_8555,N_8747);
nand U10417 (N_10417,N_8875,N_8888);
nor U10418 (N_10418,N_8646,N_9374);
nand U10419 (N_10419,N_8554,N_8441);
nand U10420 (N_10420,N_8691,N_8786);
or U10421 (N_10421,N_8529,N_8450);
or U10422 (N_10422,N_8752,N_8951);
nand U10423 (N_10423,N_8503,N_8774);
nand U10424 (N_10424,N_8747,N_9284);
xnor U10425 (N_10425,N_9013,N_9285);
nand U10426 (N_10426,N_9122,N_8492);
nand U10427 (N_10427,N_8651,N_9009);
nor U10428 (N_10428,N_8432,N_9219);
and U10429 (N_10429,N_8408,N_8776);
and U10430 (N_10430,N_9285,N_9295);
nor U10431 (N_10431,N_8636,N_8982);
nor U10432 (N_10432,N_9323,N_9498);
xnor U10433 (N_10433,N_9594,N_8855);
nor U10434 (N_10434,N_9333,N_9032);
xor U10435 (N_10435,N_9562,N_8726);
nand U10436 (N_10436,N_8878,N_8708);
xor U10437 (N_10437,N_9490,N_9290);
nor U10438 (N_10438,N_8711,N_8597);
or U10439 (N_10439,N_9554,N_8419);
and U10440 (N_10440,N_9301,N_8700);
xor U10441 (N_10441,N_9367,N_8549);
and U10442 (N_10442,N_9268,N_9183);
nand U10443 (N_10443,N_8828,N_8844);
nor U10444 (N_10444,N_9443,N_8777);
nor U10445 (N_10445,N_9021,N_9569);
nand U10446 (N_10446,N_8931,N_9465);
and U10447 (N_10447,N_9119,N_8658);
and U10448 (N_10448,N_8819,N_9118);
nor U10449 (N_10449,N_8978,N_8554);
or U10450 (N_10450,N_9553,N_8814);
xor U10451 (N_10451,N_9330,N_8675);
nor U10452 (N_10452,N_8680,N_9151);
nor U10453 (N_10453,N_9426,N_9495);
or U10454 (N_10454,N_9303,N_9372);
nor U10455 (N_10455,N_9295,N_8468);
xnor U10456 (N_10456,N_9371,N_9398);
or U10457 (N_10457,N_8676,N_9328);
and U10458 (N_10458,N_9320,N_8828);
nor U10459 (N_10459,N_9317,N_9593);
nor U10460 (N_10460,N_9060,N_9121);
nor U10461 (N_10461,N_9044,N_8529);
xnor U10462 (N_10462,N_8797,N_9005);
and U10463 (N_10463,N_8969,N_9582);
xor U10464 (N_10464,N_8759,N_9238);
and U10465 (N_10465,N_9207,N_9595);
or U10466 (N_10466,N_8732,N_9399);
or U10467 (N_10467,N_9109,N_9477);
and U10468 (N_10468,N_8441,N_8794);
xor U10469 (N_10469,N_8524,N_8569);
and U10470 (N_10470,N_9556,N_9325);
nor U10471 (N_10471,N_9196,N_9195);
and U10472 (N_10472,N_8586,N_9383);
or U10473 (N_10473,N_8884,N_8801);
or U10474 (N_10474,N_8569,N_8532);
nor U10475 (N_10475,N_8571,N_9498);
and U10476 (N_10476,N_8404,N_8545);
or U10477 (N_10477,N_9324,N_8811);
or U10478 (N_10478,N_8802,N_8918);
nand U10479 (N_10479,N_9594,N_8885);
xnor U10480 (N_10480,N_8806,N_8404);
nand U10481 (N_10481,N_8596,N_8652);
xor U10482 (N_10482,N_8715,N_8680);
and U10483 (N_10483,N_8859,N_9391);
and U10484 (N_10484,N_8509,N_9580);
nor U10485 (N_10485,N_9460,N_9014);
and U10486 (N_10486,N_8642,N_9418);
nor U10487 (N_10487,N_9426,N_9382);
nor U10488 (N_10488,N_8828,N_9516);
or U10489 (N_10489,N_8841,N_8748);
xor U10490 (N_10490,N_8699,N_9168);
nand U10491 (N_10491,N_8514,N_8676);
xnor U10492 (N_10492,N_8430,N_8728);
and U10493 (N_10493,N_8633,N_8886);
and U10494 (N_10494,N_8424,N_9353);
xnor U10495 (N_10495,N_8897,N_9442);
nor U10496 (N_10496,N_8684,N_8421);
or U10497 (N_10497,N_9486,N_8672);
nor U10498 (N_10498,N_9458,N_8960);
xor U10499 (N_10499,N_8680,N_8622);
or U10500 (N_10500,N_9566,N_9557);
or U10501 (N_10501,N_8629,N_9075);
or U10502 (N_10502,N_9404,N_9577);
nand U10503 (N_10503,N_9092,N_8402);
nand U10504 (N_10504,N_9402,N_9172);
nor U10505 (N_10505,N_8890,N_9327);
xor U10506 (N_10506,N_9126,N_8752);
and U10507 (N_10507,N_8413,N_9543);
and U10508 (N_10508,N_9557,N_9568);
xnor U10509 (N_10509,N_9406,N_9093);
xnor U10510 (N_10510,N_9273,N_8939);
nor U10511 (N_10511,N_9284,N_8661);
nor U10512 (N_10512,N_8960,N_9595);
and U10513 (N_10513,N_8779,N_9388);
nor U10514 (N_10514,N_8682,N_9088);
and U10515 (N_10515,N_8732,N_8558);
nand U10516 (N_10516,N_9580,N_9487);
xnor U10517 (N_10517,N_9026,N_8627);
or U10518 (N_10518,N_8837,N_9505);
nor U10519 (N_10519,N_8820,N_9160);
xor U10520 (N_10520,N_9416,N_9212);
xnor U10521 (N_10521,N_8818,N_8491);
or U10522 (N_10522,N_9036,N_9150);
nor U10523 (N_10523,N_9552,N_8676);
or U10524 (N_10524,N_8879,N_8966);
or U10525 (N_10525,N_8413,N_8985);
nand U10526 (N_10526,N_8893,N_9433);
xnor U10527 (N_10527,N_9518,N_8430);
or U10528 (N_10528,N_8502,N_9301);
nand U10529 (N_10529,N_8982,N_8861);
and U10530 (N_10530,N_9212,N_9505);
nor U10531 (N_10531,N_8714,N_9174);
nor U10532 (N_10532,N_8416,N_8804);
nand U10533 (N_10533,N_8800,N_8789);
nand U10534 (N_10534,N_9572,N_9564);
nor U10535 (N_10535,N_9577,N_9271);
and U10536 (N_10536,N_9426,N_9419);
or U10537 (N_10537,N_8639,N_8606);
nand U10538 (N_10538,N_8652,N_8816);
xnor U10539 (N_10539,N_9590,N_8477);
xnor U10540 (N_10540,N_9328,N_8776);
or U10541 (N_10541,N_9285,N_9084);
nor U10542 (N_10542,N_9485,N_8464);
nor U10543 (N_10543,N_8751,N_9496);
nor U10544 (N_10544,N_9018,N_9195);
xnor U10545 (N_10545,N_8880,N_9475);
nor U10546 (N_10546,N_9551,N_8743);
nor U10547 (N_10547,N_9191,N_8473);
nand U10548 (N_10548,N_8449,N_9494);
or U10549 (N_10549,N_9125,N_8967);
nor U10550 (N_10550,N_8673,N_8815);
and U10551 (N_10551,N_8840,N_8846);
nor U10552 (N_10552,N_8557,N_8512);
or U10553 (N_10553,N_8478,N_9141);
xor U10554 (N_10554,N_9532,N_8514);
or U10555 (N_10555,N_8536,N_9282);
nand U10556 (N_10556,N_9475,N_8808);
nor U10557 (N_10557,N_8516,N_9118);
and U10558 (N_10558,N_9106,N_8446);
nor U10559 (N_10559,N_9451,N_9025);
and U10560 (N_10560,N_9567,N_9394);
nand U10561 (N_10561,N_8936,N_9525);
and U10562 (N_10562,N_9225,N_8653);
nor U10563 (N_10563,N_9499,N_8479);
or U10564 (N_10564,N_9484,N_8628);
nand U10565 (N_10565,N_8542,N_9278);
or U10566 (N_10566,N_8682,N_8855);
or U10567 (N_10567,N_8833,N_8431);
and U10568 (N_10568,N_8822,N_9105);
nand U10569 (N_10569,N_9085,N_8911);
nor U10570 (N_10570,N_8443,N_8650);
nor U10571 (N_10571,N_9210,N_8902);
nor U10572 (N_10572,N_8419,N_8819);
nand U10573 (N_10573,N_8933,N_9541);
and U10574 (N_10574,N_8590,N_8500);
or U10575 (N_10575,N_8742,N_8657);
xor U10576 (N_10576,N_8955,N_8765);
nand U10577 (N_10577,N_8634,N_9010);
nor U10578 (N_10578,N_9487,N_9469);
or U10579 (N_10579,N_9573,N_8871);
nand U10580 (N_10580,N_9062,N_8530);
or U10581 (N_10581,N_8595,N_8823);
nor U10582 (N_10582,N_9214,N_9467);
nand U10583 (N_10583,N_9265,N_9270);
or U10584 (N_10584,N_8515,N_8856);
nand U10585 (N_10585,N_9559,N_9442);
xor U10586 (N_10586,N_8554,N_9245);
xnor U10587 (N_10587,N_9538,N_8443);
and U10588 (N_10588,N_8998,N_9394);
or U10589 (N_10589,N_9456,N_8439);
and U10590 (N_10590,N_8849,N_8488);
nor U10591 (N_10591,N_8522,N_8407);
nand U10592 (N_10592,N_9573,N_9434);
nand U10593 (N_10593,N_9210,N_9358);
and U10594 (N_10594,N_9141,N_8726);
xor U10595 (N_10595,N_8953,N_8930);
or U10596 (N_10596,N_8684,N_9134);
and U10597 (N_10597,N_8937,N_9190);
nor U10598 (N_10598,N_8980,N_8457);
or U10599 (N_10599,N_8955,N_9537);
nand U10600 (N_10600,N_9119,N_9250);
nor U10601 (N_10601,N_9447,N_9332);
and U10602 (N_10602,N_8421,N_8896);
nor U10603 (N_10603,N_9507,N_9003);
nor U10604 (N_10604,N_9345,N_9059);
and U10605 (N_10605,N_8893,N_9095);
and U10606 (N_10606,N_9179,N_9512);
and U10607 (N_10607,N_9259,N_9337);
nor U10608 (N_10608,N_9221,N_8795);
nor U10609 (N_10609,N_9580,N_8786);
nand U10610 (N_10610,N_9177,N_8614);
and U10611 (N_10611,N_9481,N_9049);
or U10612 (N_10612,N_8707,N_8481);
and U10613 (N_10613,N_9022,N_8408);
and U10614 (N_10614,N_9239,N_8422);
or U10615 (N_10615,N_9441,N_9019);
or U10616 (N_10616,N_9271,N_8563);
nand U10617 (N_10617,N_8467,N_9428);
nand U10618 (N_10618,N_9272,N_8828);
and U10619 (N_10619,N_9213,N_8552);
xnor U10620 (N_10620,N_9233,N_9089);
nand U10621 (N_10621,N_9492,N_9554);
xnor U10622 (N_10622,N_9491,N_9300);
xnor U10623 (N_10623,N_9355,N_8826);
or U10624 (N_10624,N_8536,N_9128);
and U10625 (N_10625,N_9391,N_8927);
nand U10626 (N_10626,N_8644,N_9026);
xor U10627 (N_10627,N_8779,N_8855);
or U10628 (N_10628,N_8931,N_8669);
and U10629 (N_10629,N_8439,N_8483);
nor U10630 (N_10630,N_9488,N_8457);
xor U10631 (N_10631,N_9122,N_8584);
and U10632 (N_10632,N_9508,N_9217);
or U10633 (N_10633,N_9025,N_9591);
xor U10634 (N_10634,N_8959,N_9395);
nor U10635 (N_10635,N_8943,N_8779);
and U10636 (N_10636,N_8443,N_8774);
xnor U10637 (N_10637,N_8870,N_9514);
xor U10638 (N_10638,N_9451,N_9266);
xor U10639 (N_10639,N_9387,N_8777);
or U10640 (N_10640,N_8427,N_9541);
nand U10641 (N_10641,N_8558,N_8404);
nand U10642 (N_10642,N_8879,N_8931);
nand U10643 (N_10643,N_8718,N_9347);
xnor U10644 (N_10644,N_8636,N_9117);
nor U10645 (N_10645,N_9326,N_8591);
and U10646 (N_10646,N_9489,N_8430);
nand U10647 (N_10647,N_9570,N_9340);
and U10648 (N_10648,N_9279,N_8521);
nand U10649 (N_10649,N_9234,N_9490);
nor U10650 (N_10650,N_8755,N_9518);
and U10651 (N_10651,N_9145,N_8662);
and U10652 (N_10652,N_9152,N_9427);
xnor U10653 (N_10653,N_8993,N_8555);
nand U10654 (N_10654,N_9585,N_8614);
nor U10655 (N_10655,N_9245,N_8605);
nand U10656 (N_10656,N_9574,N_8457);
and U10657 (N_10657,N_9104,N_9343);
and U10658 (N_10658,N_9498,N_8708);
xnor U10659 (N_10659,N_8487,N_8654);
and U10660 (N_10660,N_8658,N_9341);
and U10661 (N_10661,N_9374,N_9120);
nand U10662 (N_10662,N_9338,N_8577);
xnor U10663 (N_10663,N_8927,N_8871);
nand U10664 (N_10664,N_8743,N_9237);
nand U10665 (N_10665,N_9429,N_8822);
and U10666 (N_10666,N_8588,N_8879);
nand U10667 (N_10667,N_9235,N_9115);
nor U10668 (N_10668,N_9398,N_9300);
nand U10669 (N_10669,N_9370,N_8919);
nand U10670 (N_10670,N_9156,N_8480);
nor U10671 (N_10671,N_9418,N_8771);
and U10672 (N_10672,N_8909,N_9225);
or U10673 (N_10673,N_9268,N_9014);
nor U10674 (N_10674,N_9085,N_9291);
xor U10675 (N_10675,N_8757,N_8473);
or U10676 (N_10676,N_9387,N_9002);
nand U10677 (N_10677,N_8704,N_9587);
nor U10678 (N_10678,N_8451,N_8523);
nor U10679 (N_10679,N_8506,N_8672);
and U10680 (N_10680,N_8639,N_9483);
xnor U10681 (N_10681,N_8790,N_9449);
xnor U10682 (N_10682,N_9536,N_9192);
or U10683 (N_10683,N_8728,N_8850);
and U10684 (N_10684,N_8883,N_9326);
nor U10685 (N_10685,N_9038,N_9518);
nor U10686 (N_10686,N_8576,N_9023);
nor U10687 (N_10687,N_8625,N_8575);
and U10688 (N_10688,N_9076,N_8899);
xnor U10689 (N_10689,N_9111,N_9268);
nor U10690 (N_10690,N_9336,N_8618);
xor U10691 (N_10691,N_8797,N_9588);
nand U10692 (N_10692,N_9504,N_9307);
nor U10693 (N_10693,N_8558,N_9479);
nor U10694 (N_10694,N_9233,N_8864);
and U10695 (N_10695,N_9178,N_8522);
or U10696 (N_10696,N_8589,N_8471);
and U10697 (N_10697,N_9007,N_9243);
and U10698 (N_10698,N_8615,N_8552);
or U10699 (N_10699,N_8474,N_8786);
or U10700 (N_10700,N_9394,N_8884);
nor U10701 (N_10701,N_8693,N_9496);
nor U10702 (N_10702,N_8503,N_8688);
nand U10703 (N_10703,N_8702,N_8696);
xor U10704 (N_10704,N_9441,N_8556);
nor U10705 (N_10705,N_9340,N_9327);
nand U10706 (N_10706,N_8957,N_8606);
nand U10707 (N_10707,N_9327,N_8897);
or U10708 (N_10708,N_8681,N_8768);
nor U10709 (N_10709,N_8894,N_8824);
and U10710 (N_10710,N_9563,N_9567);
nor U10711 (N_10711,N_9144,N_9299);
or U10712 (N_10712,N_9172,N_8641);
xor U10713 (N_10713,N_8843,N_8820);
or U10714 (N_10714,N_8513,N_8965);
nand U10715 (N_10715,N_8752,N_9543);
or U10716 (N_10716,N_9011,N_8813);
and U10717 (N_10717,N_9558,N_8400);
nand U10718 (N_10718,N_8429,N_8411);
xor U10719 (N_10719,N_8405,N_9490);
nor U10720 (N_10720,N_9116,N_8724);
nand U10721 (N_10721,N_8566,N_9105);
or U10722 (N_10722,N_8982,N_8710);
nor U10723 (N_10723,N_9446,N_9152);
and U10724 (N_10724,N_9436,N_8458);
xor U10725 (N_10725,N_9255,N_8760);
nand U10726 (N_10726,N_9089,N_8911);
nor U10727 (N_10727,N_8428,N_9426);
nand U10728 (N_10728,N_8757,N_9443);
nand U10729 (N_10729,N_9504,N_8619);
xor U10730 (N_10730,N_8454,N_8890);
nor U10731 (N_10731,N_9452,N_8924);
nand U10732 (N_10732,N_8874,N_8983);
nor U10733 (N_10733,N_8663,N_8993);
or U10734 (N_10734,N_9021,N_8584);
or U10735 (N_10735,N_9118,N_8989);
or U10736 (N_10736,N_9076,N_8470);
and U10737 (N_10737,N_8862,N_8478);
nor U10738 (N_10738,N_9312,N_8651);
xor U10739 (N_10739,N_8563,N_8895);
or U10740 (N_10740,N_8672,N_9592);
nand U10741 (N_10741,N_8813,N_9245);
and U10742 (N_10742,N_8610,N_8871);
or U10743 (N_10743,N_9113,N_8702);
xor U10744 (N_10744,N_9073,N_8750);
nor U10745 (N_10745,N_8564,N_9421);
xnor U10746 (N_10746,N_9065,N_9277);
nand U10747 (N_10747,N_9363,N_9051);
and U10748 (N_10748,N_9039,N_9538);
nand U10749 (N_10749,N_9118,N_9158);
xor U10750 (N_10750,N_9426,N_9225);
and U10751 (N_10751,N_8718,N_9491);
nand U10752 (N_10752,N_8856,N_9049);
nand U10753 (N_10753,N_9260,N_8791);
nor U10754 (N_10754,N_8499,N_9084);
xnor U10755 (N_10755,N_9273,N_9112);
nor U10756 (N_10756,N_8996,N_9078);
nor U10757 (N_10757,N_8488,N_9253);
xnor U10758 (N_10758,N_9571,N_9076);
and U10759 (N_10759,N_9366,N_8989);
xnor U10760 (N_10760,N_9025,N_8924);
nand U10761 (N_10761,N_9205,N_8892);
nor U10762 (N_10762,N_8660,N_8510);
and U10763 (N_10763,N_8605,N_9528);
nor U10764 (N_10764,N_9384,N_8906);
or U10765 (N_10765,N_8611,N_9095);
and U10766 (N_10766,N_9300,N_9081);
and U10767 (N_10767,N_8617,N_8766);
or U10768 (N_10768,N_9506,N_9486);
and U10769 (N_10769,N_8785,N_9291);
and U10770 (N_10770,N_9049,N_8631);
nand U10771 (N_10771,N_9506,N_8411);
and U10772 (N_10772,N_9346,N_8751);
nor U10773 (N_10773,N_9032,N_9192);
and U10774 (N_10774,N_8750,N_9113);
or U10775 (N_10775,N_9189,N_9524);
xnor U10776 (N_10776,N_9283,N_8471);
nor U10777 (N_10777,N_8946,N_8710);
nand U10778 (N_10778,N_8994,N_8805);
nand U10779 (N_10779,N_9175,N_8468);
nand U10780 (N_10780,N_9584,N_8976);
xnor U10781 (N_10781,N_9337,N_8915);
and U10782 (N_10782,N_9362,N_8462);
nor U10783 (N_10783,N_8994,N_9195);
nand U10784 (N_10784,N_9338,N_9000);
nor U10785 (N_10785,N_9174,N_8460);
nand U10786 (N_10786,N_8740,N_9417);
nor U10787 (N_10787,N_8951,N_8664);
and U10788 (N_10788,N_9008,N_9530);
xnor U10789 (N_10789,N_8802,N_8834);
or U10790 (N_10790,N_8611,N_8455);
xnor U10791 (N_10791,N_9153,N_9132);
or U10792 (N_10792,N_9232,N_8488);
xor U10793 (N_10793,N_8483,N_8930);
nor U10794 (N_10794,N_8833,N_8719);
xor U10795 (N_10795,N_8999,N_9168);
xor U10796 (N_10796,N_9067,N_9575);
xnor U10797 (N_10797,N_8706,N_9390);
xor U10798 (N_10798,N_8820,N_9343);
nand U10799 (N_10799,N_8881,N_8656);
nand U10800 (N_10800,N_10721,N_10372);
nor U10801 (N_10801,N_10131,N_10737);
and U10802 (N_10802,N_10300,N_10107);
and U10803 (N_10803,N_10215,N_9838);
nand U10804 (N_10804,N_10796,N_10074);
or U10805 (N_10805,N_10023,N_10393);
and U10806 (N_10806,N_10660,N_10236);
and U10807 (N_10807,N_9656,N_9957);
nand U10808 (N_10808,N_10744,N_10109);
and U10809 (N_10809,N_9954,N_9749);
or U10810 (N_10810,N_10212,N_9840);
nand U10811 (N_10811,N_10589,N_10592);
xnor U10812 (N_10812,N_10580,N_9972);
and U10813 (N_10813,N_9768,N_9779);
or U10814 (N_10814,N_10041,N_10134);
nor U10815 (N_10815,N_10062,N_10329);
and U10816 (N_10816,N_10351,N_10112);
nor U10817 (N_10817,N_10021,N_10797);
nand U10818 (N_10818,N_10216,N_9661);
and U10819 (N_10819,N_9645,N_9644);
xnor U10820 (N_10820,N_9652,N_9793);
nand U10821 (N_10821,N_10493,N_10222);
nor U10822 (N_10822,N_10475,N_10101);
nand U10823 (N_10823,N_9858,N_9654);
nand U10824 (N_10824,N_10069,N_10418);
xor U10825 (N_10825,N_10307,N_10358);
xnor U10826 (N_10826,N_10346,N_10297);
and U10827 (N_10827,N_10480,N_10534);
nor U10828 (N_10828,N_10170,N_10405);
nor U10829 (N_10829,N_10277,N_10442);
nand U10830 (N_10830,N_9717,N_10715);
and U10831 (N_10831,N_9657,N_9751);
nand U10832 (N_10832,N_9952,N_10410);
xnor U10833 (N_10833,N_9942,N_9807);
and U10834 (N_10834,N_10146,N_10298);
nand U10835 (N_10835,N_10100,N_10750);
or U10836 (N_10836,N_10164,N_9628);
and U10837 (N_10837,N_10070,N_9960);
nand U10838 (N_10838,N_10123,N_9669);
or U10839 (N_10839,N_10595,N_10273);
nand U10840 (N_10840,N_9785,N_9995);
xor U10841 (N_10841,N_10720,N_10621);
xor U10842 (N_10842,N_10600,N_10743);
nand U10843 (N_10843,N_9653,N_10427);
nand U10844 (N_10844,N_9755,N_9776);
and U10845 (N_10845,N_10508,N_10068);
and U10846 (N_10846,N_9873,N_9854);
nand U10847 (N_10847,N_10516,N_10067);
nand U10848 (N_10848,N_9701,N_9870);
nand U10849 (N_10849,N_10369,N_10723);
or U10850 (N_10850,N_10088,N_10285);
xor U10851 (N_10851,N_10455,N_10762);
xnor U10852 (N_10852,N_9745,N_10584);
nor U10853 (N_10853,N_10782,N_10717);
and U10854 (N_10854,N_10703,N_9765);
nand U10855 (N_10855,N_9947,N_10500);
nand U10856 (N_10856,N_10596,N_9912);
nor U10857 (N_10857,N_10634,N_10249);
or U10858 (N_10858,N_9961,N_9844);
nor U10859 (N_10859,N_10471,N_10624);
xnor U10860 (N_10860,N_9721,N_9875);
xnor U10861 (N_10861,N_10447,N_10356);
nor U10862 (N_10862,N_10226,N_9673);
and U10863 (N_10863,N_10323,N_9603);
or U10864 (N_10864,N_10110,N_10328);
xnor U10865 (N_10865,N_10566,N_10787);
xnor U10866 (N_10866,N_9898,N_9797);
and U10867 (N_10867,N_10177,N_10055);
or U10868 (N_10868,N_9635,N_9630);
nand U10869 (N_10869,N_10711,N_9773);
and U10870 (N_10870,N_10213,N_10675);
and U10871 (N_10871,N_9633,N_10003);
and U10872 (N_10872,N_10371,N_9623);
nor U10873 (N_10873,N_10160,N_10125);
nand U10874 (N_10874,N_9924,N_10748);
nand U10875 (N_10875,N_10487,N_10658);
nor U10876 (N_10876,N_9850,N_9762);
xnor U10877 (N_10877,N_9837,N_10609);
and U10878 (N_10878,N_9889,N_10384);
or U10879 (N_10879,N_9682,N_10034);
xor U10880 (N_10880,N_9909,N_10324);
or U10881 (N_10881,N_10257,N_9607);
nand U10882 (N_10882,N_10132,N_10504);
nand U10883 (N_10883,N_10666,N_10407);
and U10884 (N_10884,N_9910,N_10562);
nor U10885 (N_10885,N_9987,N_10630);
nand U10886 (N_10886,N_9977,N_10718);
nand U10887 (N_10887,N_9935,N_10684);
xnor U10888 (N_10888,N_10054,N_10518);
xnor U10889 (N_10889,N_10078,N_10312);
nor U10890 (N_10890,N_10081,N_9948);
and U10891 (N_10891,N_10044,N_10509);
xor U10892 (N_10892,N_10202,N_9710);
or U10893 (N_10893,N_10308,N_10191);
or U10894 (N_10894,N_10519,N_10671);
nor U10895 (N_10895,N_10408,N_10753);
nand U10896 (N_10896,N_9691,N_10036);
nor U10897 (N_10897,N_10238,N_10118);
xor U10898 (N_10898,N_9651,N_9887);
or U10899 (N_10899,N_10174,N_9930);
nor U10900 (N_10900,N_10449,N_10360);
nor U10901 (N_10901,N_10166,N_9668);
nand U10902 (N_10902,N_9696,N_10198);
xnor U10903 (N_10903,N_10057,N_10108);
xor U10904 (N_10904,N_10063,N_9883);
and U10905 (N_10905,N_10294,N_10138);
or U10906 (N_10906,N_10499,N_10714);
or U10907 (N_10907,N_10362,N_10367);
xnor U10908 (N_10908,N_9660,N_10223);
nor U10909 (N_10909,N_10093,N_10775);
and U10910 (N_10910,N_10565,N_9852);
nor U10911 (N_10911,N_10537,N_10317);
xnor U10912 (N_10912,N_9993,N_10029);
nand U10913 (N_10913,N_9687,N_10525);
nand U10914 (N_10914,N_10709,N_10186);
and U10915 (N_10915,N_10306,N_9800);
nand U10916 (N_10916,N_9980,N_10576);
xnor U10917 (N_10917,N_10610,N_9746);
nand U10918 (N_10918,N_10465,N_9845);
and U10919 (N_10919,N_9632,N_10413);
and U10920 (N_10920,N_10172,N_10645);
nand U10921 (N_10921,N_10183,N_10496);
or U10922 (N_10922,N_10698,N_10326);
or U10923 (N_10923,N_10615,N_10700);
nand U10924 (N_10924,N_10605,N_10613);
or U10925 (N_10925,N_10578,N_9784);
xor U10926 (N_10926,N_10339,N_9759);
nor U10927 (N_10927,N_9662,N_10373);
nand U10928 (N_10928,N_10084,N_10728);
nor U10929 (N_10929,N_10248,N_9692);
xor U10930 (N_10930,N_9629,N_10270);
or U10931 (N_10931,N_10757,N_9777);
or U10932 (N_10932,N_10602,N_10401);
nand U10933 (N_10933,N_9724,N_9842);
nand U10934 (N_10934,N_9833,N_10422);
nor U10935 (N_10935,N_9857,N_10338);
and U10936 (N_10936,N_10586,N_10106);
and U10937 (N_10937,N_10594,N_10667);
and U10938 (N_10938,N_10486,N_10451);
or U10939 (N_10939,N_10706,N_10195);
or U10940 (N_10940,N_9926,N_10309);
nor U10941 (N_10941,N_9665,N_10627);
or U10942 (N_10942,N_10391,N_10161);
and U10943 (N_10943,N_9631,N_10386);
nand U10944 (N_10944,N_10544,N_10253);
and U10945 (N_10945,N_10702,N_10217);
xor U10946 (N_10946,N_10090,N_10664);
or U10947 (N_10947,N_10210,N_10740);
nand U10948 (N_10948,N_9610,N_10235);
nand U10949 (N_10949,N_10739,N_9754);
xor U10950 (N_10950,N_9764,N_10563);
nand U10951 (N_10951,N_9973,N_10382);
or U10952 (N_10952,N_10794,N_10481);
and U10953 (N_10953,N_10561,N_9819);
and U10954 (N_10954,N_10431,N_9893);
xnor U10955 (N_10955,N_10414,N_9975);
nand U10956 (N_10956,N_10653,N_9982);
nand U10957 (N_10957,N_10406,N_10734);
and U10958 (N_10958,N_10502,N_10148);
and U10959 (N_10959,N_9684,N_10420);
nor U10960 (N_10960,N_9902,N_9802);
and U10961 (N_10961,N_10348,N_10587);
nor U10962 (N_10962,N_10548,N_10478);
nor U10963 (N_10963,N_10535,N_10683);
or U10964 (N_10964,N_9698,N_9625);
nand U10965 (N_10965,N_9864,N_10581);
nand U10966 (N_10966,N_9865,N_9695);
and U10967 (N_10967,N_9997,N_10488);
nor U10968 (N_10968,N_9674,N_10377);
nand U10969 (N_10969,N_10644,N_10462);
and U10970 (N_10970,N_10045,N_9822);
or U10971 (N_10971,N_10704,N_9782);
or U10972 (N_10972,N_10365,N_10189);
nor U10973 (N_10973,N_10521,N_9931);
or U10974 (N_10974,N_10343,N_9892);
nor U10975 (N_10975,N_10674,N_10010);
nor U10976 (N_10976,N_9938,N_10283);
nand U10977 (N_10977,N_10262,N_10553);
or U10978 (N_10978,N_10321,N_9795);
and U10979 (N_10979,N_9976,N_9703);
or U10980 (N_10980,N_10145,N_10231);
and U10981 (N_10981,N_10545,N_9693);
and U10982 (N_10982,N_10375,N_10278);
nand U10983 (N_10983,N_10559,N_10696);
nand U10984 (N_10984,N_10642,N_9820);
or U10985 (N_10985,N_10780,N_10685);
nand U10986 (N_10986,N_9715,N_9871);
or U10987 (N_10987,N_10479,N_10147);
xor U10988 (N_10988,N_10697,N_10793);
xor U10989 (N_10989,N_9805,N_9816);
nor U10990 (N_10990,N_10011,N_9879);
xnor U10991 (N_10991,N_9613,N_10228);
nand U10992 (N_10992,N_10736,N_9809);
nor U10993 (N_10993,N_9829,N_9915);
nor U10994 (N_10994,N_9876,N_10378);
nand U10995 (N_10995,N_10149,N_10532);
nand U10996 (N_10996,N_10175,N_10117);
and U10997 (N_10997,N_9786,N_10608);
or U10998 (N_10998,N_10423,N_10591);
or U10999 (N_10999,N_10686,N_10527);
xnor U11000 (N_11000,N_9944,N_10016);
nor U11001 (N_11001,N_10505,N_10182);
and U11002 (N_11002,N_9766,N_10681);
nor U11003 (N_11003,N_10390,N_10141);
and U11004 (N_11004,N_10655,N_10028);
or U11005 (N_11005,N_10180,N_10232);
nand U11006 (N_11006,N_10791,N_10256);
nor U11007 (N_11007,N_10176,N_9836);
nor U11008 (N_11008,N_10272,N_10344);
xor U11009 (N_11009,N_10370,N_10220);
or U11010 (N_11010,N_10547,N_10353);
nand U11011 (N_11011,N_9729,N_10243);
nor U11012 (N_11012,N_10233,N_10484);
nor U11013 (N_11013,N_9856,N_9831);
and U11014 (N_11014,N_10234,N_10474);
xor U11015 (N_11015,N_9801,N_10638);
xor U11016 (N_11016,N_10647,N_9906);
nand U11017 (N_11017,N_10281,N_10458);
xnor U11018 (N_11018,N_9641,N_10320);
xor U11019 (N_11019,N_9620,N_10741);
and U11020 (N_11020,N_10035,N_10713);
or U11021 (N_11021,N_10014,N_9925);
and U11022 (N_11022,N_10072,N_10207);
nor U11023 (N_11023,N_10032,N_10156);
nand U11024 (N_11024,N_10157,N_9771);
and U11025 (N_11025,N_10582,N_9895);
nand U11026 (N_11026,N_10204,N_10211);
xnor U11027 (N_11027,N_10064,N_10227);
xnor U11028 (N_11028,N_9677,N_9919);
xnor U11029 (N_11029,N_10473,N_9888);
or U11030 (N_11030,N_9953,N_10244);
xor U11031 (N_11031,N_9753,N_9928);
nand U11032 (N_11032,N_9742,N_9913);
nand U11033 (N_11033,N_9886,N_9604);
or U11034 (N_11034,N_9946,N_9705);
or U11035 (N_11035,N_9818,N_10389);
xor U11036 (N_11036,N_10461,N_10395);
xnor U11037 (N_11037,N_10575,N_10583);
nand U11038 (N_11038,N_10603,N_10517);
and U11039 (N_11039,N_10133,N_9951);
xor U11040 (N_11040,N_10073,N_10769);
nand U11041 (N_11041,N_10513,N_10716);
nand U11042 (N_11042,N_10366,N_10641);
nand U11043 (N_11043,N_10619,N_9861);
nand U11044 (N_11044,N_10319,N_9728);
nor U11045 (N_11045,N_9704,N_9659);
or U11046 (N_11046,N_10710,N_10444);
nor U11047 (N_11047,N_9646,N_10568);
nor U11048 (N_11048,N_10430,N_10026);
nand U11049 (N_11049,N_9970,N_10585);
nand U11050 (N_11050,N_9711,N_10543);
xor U11051 (N_11051,N_10295,N_9903);
or U11052 (N_11052,N_10733,N_9634);
nand U11053 (N_11053,N_9789,N_10038);
and U11054 (N_11054,N_9941,N_10047);
or U11055 (N_11055,N_10279,N_10002);
nand U11056 (N_11056,N_10662,N_10425);
or U11057 (N_11057,N_9647,N_10322);
or U11058 (N_11058,N_10424,N_10169);
or U11059 (N_11059,N_9823,N_10311);
and U11060 (N_11060,N_10103,N_9991);
xor U11061 (N_11061,N_10115,N_9914);
and U11062 (N_11062,N_10126,N_10538);
nand U11063 (N_11063,N_9979,N_10150);
or U11064 (N_11064,N_10102,N_10680);
nand U11065 (N_11065,N_9774,N_10622);
and U11066 (N_11066,N_10551,N_10552);
and U11067 (N_11067,N_10719,N_9978);
xor U11068 (N_11068,N_10007,N_10225);
or U11069 (N_11069,N_9923,N_9843);
xor U11070 (N_11070,N_10392,N_10795);
nor U11071 (N_11071,N_9621,N_10725);
nor U11072 (N_11072,N_10764,N_10554);
xnor U11073 (N_11073,N_10490,N_10053);
or U11074 (N_11074,N_10550,N_9694);
nor U11075 (N_11075,N_10492,N_10242);
xor U11076 (N_11076,N_9707,N_9996);
nand U11077 (N_11077,N_10699,N_10785);
xor U11078 (N_11078,N_9901,N_9963);
nand U11079 (N_11079,N_9758,N_10773);
xnor U11080 (N_11080,N_10152,N_10245);
nand U11081 (N_11081,N_9612,N_9968);
nor U11082 (N_11082,N_9722,N_9955);
nor U11083 (N_11083,N_10438,N_10334);
xor U11084 (N_11084,N_10193,N_10097);
nand U11085 (N_11085,N_10267,N_9747);
xor U11086 (N_11086,N_10315,N_9808);
xnor U11087 (N_11087,N_9832,N_10677);
nand U11088 (N_11088,N_10251,N_9943);
nor U11089 (N_11089,N_10436,N_10441);
and U11090 (N_11090,N_10403,N_10004);
and U11091 (N_11091,N_10105,N_10567);
xnor U11092 (N_11092,N_10087,N_10094);
nand U11093 (N_11093,N_9750,N_10031);
xnor U11094 (N_11094,N_10122,N_10464);
and U11095 (N_11095,N_10777,N_10650);
xnor U11096 (N_11096,N_10558,N_10676);
xnor U11097 (N_11097,N_10799,N_10264);
xor U11098 (N_11098,N_10665,N_10252);
or U11099 (N_11099,N_10142,N_10411);
xor U11100 (N_11100,N_9642,N_10625);
or U11101 (N_11101,N_10588,N_10540);
nor U11102 (N_11102,N_10357,N_9670);
nor U11103 (N_11103,N_10491,N_10203);
and U11104 (N_11104,N_10778,N_10679);
nor U11105 (N_11105,N_10310,N_10289);
or U11106 (N_11106,N_10798,N_9900);
or U11107 (N_11107,N_9846,N_10620);
nor U11108 (N_11108,N_10432,N_10687);
or U11109 (N_11109,N_9737,N_10606);
xor U11110 (N_11110,N_10765,N_9894);
nor U11111 (N_11111,N_10571,N_10789);
xor U11112 (N_11112,N_10639,N_10526);
or U11113 (N_11113,N_10507,N_10417);
and U11114 (N_11114,N_10305,N_10768);
nor U11115 (N_11115,N_10712,N_9853);
nor U11116 (N_11116,N_9908,N_10400);
or U11117 (N_11117,N_10098,N_10275);
xnor U11118 (N_11118,N_9981,N_9732);
nor U11119 (N_11119,N_9890,N_10165);
or U11120 (N_11120,N_10095,N_9839);
or U11121 (N_11121,N_10628,N_9663);
or U11122 (N_11122,N_9741,N_10426);
xor U11123 (N_11123,N_10668,N_10318);
xor U11124 (N_11124,N_10199,N_10776);
or U11125 (N_11125,N_9804,N_9932);
xor U11126 (N_11126,N_10524,N_9740);
nand U11127 (N_11127,N_10691,N_10135);
xnor U11128 (N_11128,N_10077,N_10397);
and U11129 (N_11129,N_10597,N_9880);
nand U11130 (N_11130,N_9867,N_10151);
nor U11131 (N_11131,N_10541,N_10396);
xnor U11132 (N_11132,N_10695,N_9866);
or U11133 (N_11133,N_10024,N_9618);
or U11134 (N_11134,N_10255,N_9803);
nand U11135 (N_11135,N_9811,N_9605);
and U11136 (N_11136,N_10607,N_10330);
nor U11137 (N_11137,N_10460,N_9859);
nand U11138 (N_11138,N_10271,N_10482);
nand U11139 (N_11139,N_10416,N_10246);
and U11140 (N_11140,N_10076,N_10494);
or U11141 (N_11141,N_10316,N_9974);
and U11142 (N_11142,N_9969,N_9984);
nand U11143 (N_11143,N_10746,N_10477);
or U11144 (N_11144,N_9769,N_10635);
nand U11145 (N_11145,N_9720,N_10497);
and U11146 (N_11146,N_10722,N_10197);
xor U11147 (N_11147,N_10506,N_9798);
nand U11148 (N_11148,N_10200,N_10448);
nor U11149 (N_11149,N_10332,N_9676);
and U11150 (N_11150,N_9992,N_10756);
and U11151 (N_11151,N_9950,N_9735);
and U11152 (N_11152,N_10171,N_10659);
xnor U11153 (N_11153,N_10701,N_10636);
nor U11154 (N_11154,N_10009,N_10124);
nor U11155 (N_11155,N_10618,N_9874);
nand U11156 (N_11156,N_9940,N_9649);
nor U11157 (N_11157,N_10304,N_9655);
or U11158 (N_11158,N_10091,N_10205);
or U11159 (N_11159,N_10688,N_10303);
or U11160 (N_11160,N_9916,N_10060);
nand U11161 (N_11161,N_9998,N_10219);
nor U11162 (N_11162,N_10089,N_10155);
nand U11163 (N_11163,N_10190,N_9706);
nor U11164 (N_11164,N_10669,N_9681);
nor U11165 (N_11165,N_9939,N_10292);
nand U11166 (N_11166,N_9964,N_9637);
or U11167 (N_11167,N_10459,N_10646);
xor U11168 (N_11168,N_10230,N_9855);
or U11169 (N_11169,N_10623,N_10086);
and U11170 (N_11170,N_9622,N_10663);
or U11171 (N_11171,N_10466,N_9882);
xnor U11172 (N_11172,N_10376,N_9686);
xor U11173 (N_11173,N_10269,N_10049);
and U11174 (N_11174,N_9849,N_10221);
nor U11175 (N_11175,N_10046,N_10654);
nand U11176 (N_11176,N_10616,N_10450);
and U11177 (N_11177,N_9863,N_10116);
xor U11178 (N_11178,N_10290,N_9799);
xor U11179 (N_11179,N_10192,N_10783);
xor U11180 (N_11180,N_9827,N_9937);
or U11181 (N_11181,N_9643,N_9884);
or U11182 (N_11182,N_9760,N_10162);
or U11183 (N_11183,N_10188,N_10005);
or U11184 (N_11184,N_10435,N_10560);
nand U11185 (N_11185,N_9985,N_10261);
and U11186 (N_11186,N_10542,N_10633);
xnor U11187 (N_11187,N_9949,N_9640);
and U11188 (N_11188,N_9962,N_10598);
nor U11189 (N_11189,N_9602,N_9601);
or U11190 (N_11190,N_10564,N_9986);
xnor U11191 (N_11191,N_9713,N_10179);
nand U11192 (N_11192,N_10184,N_9966);
or U11193 (N_11193,N_10331,N_10761);
or U11194 (N_11194,N_9787,N_10167);
xor U11195 (N_11195,N_10470,N_10579);
or U11196 (N_11196,N_10224,N_10286);
and U11197 (N_11197,N_9714,N_10130);
and U11198 (N_11198,N_10515,N_10453);
xnor U11199 (N_11199,N_10439,N_10614);
nand U11200 (N_11200,N_10394,N_10648);
nor U11201 (N_11201,N_9812,N_9817);
nor U11202 (N_11202,N_10388,N_10066);
nor U11203 (N_11203,N_10531,N_10240);
nor U11204 (N_11204,N_10751,N_9851);
nor U11205 (N_11205,N_9615,N_9790);
xor U11206 (N_11206,N_9835,N_10239);
nand U11207 (N_11207,N_10083,N_9617);
xnor U11208 (N_11208,N_9815,N_10314);
nor U11209 (N_11209,N_10380,N_10327);
nor U11210 (N_11210,N_9934,N_10682);
nor U11211 (N_11211,N_9756,N_10254);
nor U11212 (N_11212,N_9666,N_10387);
or U11213 (N_11213,N_10412,N_10409);
xor U11214 (N_11214,N_9994,N_10443);
or U11215 (N_11215,N_9783,N_9671);
or U11216 (N_11216,N_10335,N_10128);
and U11217 (N_11217,N_10043,N_10129);
and U11218 (N_11218,N_9614,N_10670);
nand U11219 (N_11219,N_10454,N_10693);
xor U11220 (N_11220,N_10570,N_10104);
xor U11221 (N_11221,N_10730,N_10689);
and U11222 (N_11222,N_10181,N_9794);
nor U11223 (N_11223,N_10065,N_9945);
nor U11224 (N_11224,N_10774,N_10139);
nand U11225 (N_11225,N_10381,N_10536);
xor U11226 (N_11226,N_9791,N_10355);
and U11227 (N_11227,N_10779,N_10738);
or U11228 (N_11228,N_9824,N_9796);
and U11229 (N_11229,N_9689,N_10079);
or U11230 (N_11230,N_9821,N_10260);
xor U11231 (N_11231,N_9697,N_9841);
nand U11232 (N_11232,N_10237,N_10732);
or U11233 (N_11233,N_10048,N_9936);
nor U11234 (N_11234,N_9770,N_10018);
xor U11235 (N_11235,N_9806,N_10333);
xnor U11236 (N_11236,N_10557,N_10555);
or U11237 (N_11237,N_9611,N_10434);
nand U11238 (N_11238,N_9626,N_10402);
or U11239 (N_11239,N_9716,N_10013);
xnor U11240 (N_11240,N_10452,N_9868);
nor U11241 (N_11241,N_10113,N_10061);
and U11242 (N_11242,N_9685,N_9619);
xnor U11243 (N_11243,N_10259,N_10569);
and U11244 (N_11244,N_10241,N_9727);
nor U11245 (N_11245,N_10040,N_10030);
xor U11246 (N_11246,N_10428,N_10052);
and U11247 (N_11247,N_9983,N_10092);
and U11248 (N_11248,N_9830,N_9744);
nor U11249 (N_11249,N_10533,N_9639);
and U11250 (N_11250,N_10185,N_10096);
xnor U11251 (N_11251,N_9967,N_10178);
nand U11252 (N_11252,N_9699,N_10291);
xor U11253 (N_11253,N_9638,N_10173);
or U11254 (N_11254,N_9965,N_10421);
nor U11255 (N_11255,N_9690,N_9897);
and U11256 (N_11256,N_10056,N_9679);
nor U11257 (N_11257,N_10604,N_10763);
and U11258 (N_11258,N_10398,N_9648);
nand U11259 (N_11259,N_10006,N_9726);
nand U11260 (N_11260,N_9907,N_10467);
nand U11261 (N_11261,N_10008,N_10349);
nor U11262 (N_11262,N_10530,N_9683);
and U11263 (N_11263,N_9872,N_10050);
and U11264 (N_11264,N_9667,N_10229);
and U11265 (N_11265,N_10788,N_10302);
or U11266 (N_11266,N_10293,N_10759);
nor U11267 (N_11267,N_10631,N_10726);
nand U11268 (N_11268,N_9825,N_10501);
nor U11269 (N_11269,N_10159,N_9920);
nand U11270 (N_11270,N_10752,N_9911);
xor U11271 (N_11271,N_10694,N_10483);
nand U11272 (N_11272,N_9725,N_9956);
nand U11273 (N_11273,N_10144,N_10637);
and U11274 (N_11274,N_9904,N_10601);
or U11275 (N_11275,N_9921,N_9734);
or U11276 (N_11276,N_10347,N_9989);
and U11277 (N_11277,N_9810,N_10656);
or U11278 (N_11278,N_10708,N_10282);
and U11279 (N_11279,N_9600,N_9761);
and U11280 (N_11280,N_9896,N_10770);
and U11281 (N_11281,N_10790,N_10114);
or U11282 (N_11282,N_10206,N_10280);
or U11283 (N_11283,N_9702,N_10218);
and U11284 (N_11284,N_10336,N_9828);
nor U11285 (N_11285,N_10556,N_10012);
and U11286 (N_11286,N_10617,N_10476);
xor U11287 (N_11287,N_10503,N_10258);
nand U11288 (N_11288,N_10341,N_10590);
or U11289 (N_11289,N_10051,N_10766);
or U11290 (N_11290,N_10154,N_10652);
nand U11291 (N_11291,N_10456,N_10364);
xnor U11292 (N_11292,N_10784,N_9636);
nor U11293 (N_11293,N_10099,N_9933);
nor U11294 (N_11294,N_9608,N_10692);
xnor U11295 (N_11295,N_10136,N_10284);
or U11296 (N_11296,N_10629,N_10379);
xnor U11297 (N_11297,N_10265,N_10127);
nand U11298 (N_11298,N_9834,N_9733);
nor U11299 (N_11299,N_10758,N_10071);
nor U11300 (N_11300,N_10368,N_10037);
xor U11301 (N_11301,N_10727,N_10268);
or U11302 (N_11302,N_10352,N_10001);
nor U11303 (N_11303,N_9606,N_10489);
xnor U11304 (N_11304,N_10022,N_10276);
nor U11305 (N_11305,N_10313,N_10153);
or U11306 (N_11306,N_10786,N_10196);
and U11307 (N_11307,N_10514,N_9877);
or U11308 (N_11308,N_10745,N_9738);
and U11309 (N_11309,N_10399,N_10288);
xor U11310 (N_11310,N_10523,N_10163);
xor U11311 (N_11311,N_10350,N_10760);
nand U11312 (N_11312,N_9748,N_10599);
nor U11313 (N_11313,N_10361,N_10143);
and U11314 (N_11314,N_10485,N_10299);
and U11315 (N_11315,N_9778,N_10168);
or U11316 (N_11316,N_9616,N_10643);
or U11317 (N_11317,N_9781,N_9767);
xor U11318 (N_11318,N_10781,N_9813);
or U11319 (N_11319,N_10137,N_9719);
or U11320 (N_11320,N_10075,N_10767);
nor U11321 (N_11321,N_10672,N_10301);
nand U11322 (N_11322,N_10121,N_10042);
nor U11323 (N_11323,N_10468,N_10082);
and U11324 (N_11324,N_10495,N_10574);
nand U11325 (N_11325,N_10015,N_10250);
nand U11326 (N_11326,N_10385,N_9917);
or U11327 (N_11327,N_9999,N_10632);
xnor U11328 (N_11328,N_10287,N_10498);
and U11329 (N_11329,N_10039,N_10457);
nand U11330 (N_11330,N_9709,N_10549);
nor U11331 (N_11331,N_9922,N_9990);
nor U11332 (N_11332,N_9775,N_9730);
nor U11333 (N_11333,N_9929,N_9678);
or U11334 (N_11334,N_10678,N_9988);
nor U11335 (N_11335,N_10440,N_10027);
xor U11336 (N_11336,N_9869,N_10263);
xor U11337 (N_11337,N_10187,N_10194);
nand U11338 (N_11338,N_10707,N_10437);
or U11339 (N_11339,N_9650,N_10345);
and U11340 (N_11340,N_10325,N_9757);
or U11341 (N_11341,N_10059,N_10747);
nor U11342 (N_11342,N_10419,N_10445);
nor U11343 (N_11343,N_10651,N_9848);
nand U11344 (N_11344,N_10019,N_10724);
and U11345 (N_11345,N_10731,N_10522);
nor U11346 (N_11346,N_10611,N_9885);
nor U11347 (N_11347,N_10539,N_10209);
xor U11348 (N_11348,N_9664,N_9927);
nor U11349 (N_11349,N_10749,N_10657);
nor U11350 (N_11350,N_10274,N_10577);
nand U11351 (N_11351,N_9763,N_10792);
nor U11352 (N_11352,N_10000,N_10742);
xnor U11353 (N_11353,N_10201,N_9905);
or U11354 (N_11354,N_9609,N_9743);
or U11355 (N_11355,N_10546,N_9708);
xor U11356 (N_11356,N_9739,N_10469);
nand U11357 (N_11357,N_9918,N_9891);
xor U11358 (N_11358,N_9718,N_10374);
xnor U11359 (N_11359,N_9731,N_9959);
nand U11360 (N_11360,N_10017,N_10772);
and U11361 (N_11361,N_10573,N_9624);
or U11362 (N_11362,N_9736,N_10446);
or U11363 (N_11363,N_10520,N_10771);
and U11364 (N_11364,N_10690,N_10080);
nand U11365 (N_11365,N_9672,N_10512);
or U11366 (N_11366,N_10529,N_10140);
and U11367 (N_11367,N_9826,N_9680);
or U11368 (N_11368,N_10119,N_10472);
or U11369 (N_11369,N_10593,N_9971);
or U11370 (N_11370,N_10020,N_9847);
xor U11371 (N_11371,N_10337,N_9881);
and U11372 (N_11372,N_9862,N_10266);
xnor U11373 (N_11373,N_10626,N_10340);
nand U11374 (N_11374,N_10612,N_10649);
or U11375 (N_11375,N_10433,N_10429);
xnor U11376 (N_11376,N_9792,N_10354);
or U11377 (N_11377,N_10025,N_9899);
or U11378 (N_11378,N_9772,N_10383);
nor U11379 (N_11379,N_10363,N_10640);
xnor U11380 (N_11380,N_10415,N_9780);
and U11381 (N_11381,N_10120,N_9958);
and U11382 (N_11382,N_10510,N_10208);
nor U11383 (N_11383,N_10058,N_10661);
xor U11384 (N_11384,N_9700,N_10085);
or U11385 (N_11385,N_10572,N_9878);
nor U11386 (N_11386,N_10296,N_10729);
xor U11387 (N_11387,N_9712,N_10214);
or U11388 (N_11388,N_10754,N_10342);
nand U11389 (N_11389,N_10735,N_10463);
nor U11390 (N_11390,N_10755,N_9627);
nor U11391 (N_11391,N_10673,N_9658);
xor U11392 (N_11392,N_9675,N_10247);
xnor U11393 (N_11393,N_9752,N_10158);
and U11394 (N_11394,N_9860,N_9814);
or U11395 (N_11395,N_10705,N_10528);
or U11396 (N_11396,N_10033,N_9688);
and U11397 (N_11397,N_10111,N_9788);
xor U11398 (N_11398,N_9723,N_10511);
nand U11399 (N_11399,N_10404,N_10359);
and U11400 (N_11400,N_10570,N_9839);
nand U11401 (N_11401,N_10087,N_9739);
nor U11402 (N_11402,N_10324,N_10053);
or U11403 (N_11403,N_10600,N_10259);
xor U11404 (N_11404,N_10491,N_9970);
and U11405 (N_11405,N_10312,N_9988);
and U11406 (N_11406,N_10384,N_9866);
or U11407 (N_11407,N_10404,N_9871);
nand U11408 (N_11408,N_9626,N_10336);
nand U11409 (N_11409,N_10078,N_9944);
xor U11410 (N_11410,N_10002,N_10297);
xor U11411 (N_11411,N_9945,N_10766);
and U11412 (N_11412,N_10331,N_10775);
nand U11413 (N_11413,N_9618,N_10580);
nor U11414 (N_11414,N_9782,N_9667);
nand U11415 (N_11415,N_9607,N_9700);
nand U11416 (N_11416,N_9603,N_9891);
and U11417 (N_11417,N_9660,N_9818);
or U11418 (N_11418,N_9681,N_10591);
and U11419 (N_11419,N_10575,N_10694);
and U11420 (N_11420,N_10786,N_10248);
nand U11421 (N_11421,N_9791,N_10471);
and U11422 (N_11422,N_9840,N_10194);
or U11423 (N_11423,N_10334,N_9660);
and U11424 (N_11424,N_10178,N_10037);
and U11425 (N_11425,N_10333,N_10346);
xor U11426 (N_11426,N_9660,N_10115);
or U11427 (N_11427,N_10246,N_10083);
or U11428 (N_11428,N_10491,N_10720);
nor U11429 (N_11429,N_10663,N_10381);
and U11430 (N_11430,N_9632,N_10048);
nand U11431 (N_11431,N_10127,N_10122);
or U11432 (N_11432,N_10514,N_10183);
nand U11433 (N_11433,N_10324,N_10082);
nand U11434 (N_11434,N_10265,N_10520);
xor U11435 (N_11435,N_10298,N_10153);
xor U11436 (N_11436,N_10682,N_10087);
or U11437 (N_11437,N_9967,N_9905);
xor U11438 (N_11438,N_10558,N_9741);
and U11439 (N_11439,N_10405,N_10239);
or U11440 (N_11440,N_10738,N_9791);
nand U11441 (N_11441,N_10483,N_10185);
or U11442 (N_11442,N_9697,N_10380);
nand U11443 (N_11443,N_10734,N_10667);
nand U11444 (N_11444,N_10267,N_9904);
xnor U11445 (N_11445,N_10345,N_10421);
xor U11446 (N_11446,N_9872,N_10143);
and U11447 (N_11447,N_10267,N_10306);
nand U11448 (N_11448,N_10107,N_10368);
xor U11449 (N_11449,N_10313,N_9754);
xnor U11450 (N_11450,N_10408,N_9770);
nand U11451 (N_11451,N_10378,N_9936);
or U11452 (N_11452,N_10377,N_10767);
xor U11453 (N_11453,N_9829,N_9959);
nor U11454 (N_11454,N_10647,N_10254);
and U11455 (N_11455,N_10117,N_9650);
or U11456 (N_11456,N_10377,N_10532);
xnor U11457 (N_11457,N_9634,N_9628);
nand U11458 (N_11458,N_10742,N_9929);
and U11459 (N_11459,N_10386,N_10130);
xnor U11460 (N_11460,N_10495,N_10470);
xnor U11461 (N_11461,N_9918,N_10089);
xor U11462 (N_11462,N_9835,N_10546);
nor U11463 (N_11463,N_10565,N_10177);
xnor U11464 (N_11464,N_10693,N_10635);
nand U11465 (N_11465,N_9985,N_10276);
or U11466 (N_11466,N_10203,N_10374);
and U11467 (N_11467,N_10328,N_10514);
nand U11468 (N_11468,N_10315,N_10708);
or U11469 (N_11469,N_9885,N_9621);
or U11470 (N_11470,N_10569,N_10428);
and U11471 (N_11471,N_9903,N_10511);
xnor U11472 (N_11472,N_10324,N_10274);
xnor U11473 (N_11473,N_10273,N_9949);
and U11474 (N_11474,N_10359,N_10612);
nor U11475 (N_11475,N_9807,N_10618);
nand U11476 (N_11476,N_10584,N_10555);
xnor U11477 (N_11477,N_10742,N_10412);
and U11478 (N_11478,N_10433,N_9806);
or U11479 (N_11479,N_9679,N_10588);
xnor U11480 (N_11480,N_9881,N_10612);
nand U11481 (N_11481,N_10575,N_10251);
and U11482 (N_11482,N_10026,N_9720);
or U11483 (N_11483,N_10122,N_10643);
nor U11484 (N_11484,N_9637,N_9718);
and U11485 (N_11485,N_9945,N_10602);
xnor U11486 (N_11486,N_9765,N_10623);
nor U11487 (N_11487,N_9696,N_9873);
or U11488 (N_11488,N_9733,N_9655);
nor U11489 (N_11489,N_10637,N_9986);
nor U11490 (N_11490,N_9697,N_10662);
or U11491 (N_11491,N_10344,N_10190);
nand U11492 (N_11492,N_10131,N_10777);
nand U11493 (N_11493,N_10185,N_10072);
nand U11494 (N_11494,N_9650,N_9670);
xnor U11495 (N_11495,N_10013,N_9637);
xnor U11496 (N_11496,N_10784,N_10298);
or U11497 (N_11497,N_10432,N_10178);
or U11498 (N_11498,N_9748,N_9930);
xor U11499 (N_11499,N_10759,N_10248);
or U11500 (N_11500,N_9742,N_10157);
or U11501 (N_11501,N_9827,N_9687);
and U11502 (N_11502,N_10126,N_10491);
xor U11503 (N_11503,N_10440,N_10093);
xnor U11504 (N_11504,N_10035,N_9804);
nand U11505 (N_11505,N_9774,N_10630);
nor U11506 (N_11506,N_10175,N_10235);
xor U11507 (N_11507,N_9734,N_10743);
or U11508 (N_11508,N_10668,N_10251);
or U11509 (N_11509,N_9636,N_9618);
nand U11510 (N_11510,N_9904,N_10284);
or U11511 (N_11511,N_10393,N_9686);
and U11512 (N_11512,N_10398,N_10430);
nand U11513 (N_11513,N_10292,N_10093);
or U11514 (N_11514,N_10352,N_10711);
nor U11515 (N_11515,N_9703,N_10514);
nand U11516 (N_11516,N_10123,N_9959);
xnor U11517 (N_11517,N_10427,N_10293);
or U11518 (N_11518,N_9789,N_9622);
nand U11519 (N_11519,N_9621,N_10363);
nand U11520 (N_11520,N_9998,N_9643);
or U11521 (N_11521,N_9634,N_9667);
and U11522 (N_11522,N_10095,N_10212);
nor U11523 (N_11523,N_9916,N_9815);
nor U11524 (N_11524,N_10287,N_9999);
or U11525 (N_11525,N_10626,N_9809);
or U11526 (N_11526,N_9842,N_9626);
and U11527 (N_11527,N_10498,N_10504);
nand U11528 (N_11528,N_10764,N_10261);
xnor U11529 (N_11529,N_10493,N_10138);
xnor U11530 (N_11530,N_10684,N_10032);
or U11531 (N_11531,N_10013,N_9992);
or U11532 (N_11532,N_10087,N_10508);
nor U11533 (N_11533,N_9677,N_10439);
nor U11534 (N_11534,N_9647,N_10406);
xnor U11535 (N_11535,N_10553,N_10533);
and U11536 (N_11536,N_10326,N_10592);
or U11537 (N_11537,N_10122,N_10315);
nor U11538 (N_11538,N_10034,N_9971);
nor U11539 (N_11539,N_10159,N_10212);
and U11540 (N_11540,N_10502,N_10385);
xor U11541 (N_11541,N_10751,N_10373);
nand U11542 (N_11542,N_9697,N_9960);
nor U11543 (N_11543,N_10578,N_10278);
nor U11544 (N_11544,N_9878,N_10492);
xnor U11545 (N_11545,N_10084,N_9985);
nand U11546 (N_11546,N_9706,N_10748);
and U11547 (N_11547,N_10057,N_10767);
nor U11548 (N_11548,N_10443,N_9893);
nand U11549 (N_11549,N_10110,N_9666);
xor U11550 (N_11550,N_10484,N_10732);
nor U11551 (N_11551,N_10197,N_9727);
nand U11552 (N_11552,N_9651,N_10037);
nor U11553 (N_11553,N_10480,N_10054);
nand U11554 (N_11554,N_10179,N_10730);
and U11555 (N_11555,N_9870,N_10555);
xnor U11556 (N_11556,N_10763,N_9779);
and U11557 (N_11557,N_9658,N_10266);
nand U11558 (N_11558,N_9905,N_9937);
and U11559 (N_11559,N_10188,N_10512);
nor U11560 (N_11560,N_9813,N_9853);
xor U11561 (N_11561,N_10089,N_10266);
and U11562 (N_11562,N_9917,N_10483);
or U11563 (N_11563,N_9943,N_9843);
nor U11564 (N_11564,N_9754,N_10752);
nand U11565 (N_11565,N_10698,N_10697);
nor U11566 (N_11566,N_10799,N_10518);
and U11567 (N_11567,N_9957,N_10588);
xnor U11568 (N_11568,N_10413,N_9996);
and U11569 (N_11569,N_9763,N_10715);
nor U11570 (N_11570,N_9684,N_9626);
or U11571 (N_11571,N_10405,N_10029);
and U11572 (N_11572,N_9788,N_9841);
or U11573 (N_11573,N_10383,N_9798);
and U11574 (N_11574,N_10495,N_10243);
nor U11575 (N_11575,N_10344,N_10269);
nand U11576 (N_11576,N_10569,N_10186);
or U11577 (N_11577,N_10181,N_9646);
nand U11578 (N_11578,N_9956,N_10322);
or U11579 (N_11579,N_10136,N_9860);
xnor U11580 (N_11580,N_10432,N_9779);
nand U11581 (N_11581,N_10726,N_9628);
xnor U11582 (N_11582,N_10385,N_10702);
nand U11583 (N_11583,N_10212,N_9746);
nand U11584 (N_11584,N_10496,N_10698);
or U11585 (N_11585,N_10619,N_10434);
or U11586 (N_11586,N_9974,N_10224);
xnor U11587 (N_11587,N_9860,N_10215);
or U11588 (N_11588,N_10301,N_10332);
xor U11589 (N_11589,N_9719,N_10622);
nor U11590 (N_11590,N_10490,N_10345);
nor U11591 (N_11591,N_10352,N_9761);
nand U11592 (N_11592,N_10140,N_10522);
and U11593 (N_11593,N_10068,N_10735);
nand U11594 (N_11594,N_9693,N_10134);
or U11595 (N_11595,N_9943,N_10765);
xnor U11596 (N_11596,N_10547,N_10332);
nor U11597 (N_11597,N_10172,N_10199);
nand U11598 (N_11598,N_10353,N_10683);
nand U11599 (N_11599,N_10590,N_10450);
and U11600 (N_11600,N_10698,N_10795);
or U11601 (N_11601,N_10485,N_10315);
xnor U11602 (N_11602,N_9840,N_10490);
or U11603 (N_11603,N_10454,N_10036);
and U11604 (N_11604,N_9778,N_9909);
nor U11605 (N_11605,N_9877,N_10413);
xor U11606 (N_11606,N_9737,N_10419);
nand U11607 (N_11607,N_10226,N_10760);
or U11608 (N_11608,N_9818,N_10762);
nand U11609 (N_11609,N_9909,N_10737);
or U11610 (N_11610,N_10178,N_10434);
xnor U11611 (N_11611,N_9782,N_10681);
and U11612 (N_11612,N_10002,N_9878);
and U11613 (N_11613,N_10047,N_9744);
nand U11614 (N_11614,N_10700,N_10282);
xor U11615 (N_11615,N_10786,N_10352);
or U11616 (N_11616,N_10123,N_10032);
and U11617 (N_11617,N_10174,N_9717);
nand U11618 (N_11618,N_10780,N_10405);
nand U11619 (N_11619,N_10321,N_9610);
and U11620 (N_11620,N_10053,N_10635);
and U11621 (N_11621,N_9872,N_9654);
nand U11622 (N_11622,N_9870,N_10469);
nor U11623 (N_11623,N_10684,N_9682);
nor U11624 (N_11624,N_10375,N_10527);
nor U11625 (N_11625,N_10125,N_10690);
and U11626 (N_11626,N_9710,N_10775);
or U11627 (N_11627,N_10229,N_10642);
or U11628 (N_11628,N_10404,N_9880);
or U11629 (N_11629,N_9709,N_9975);
xnor U11630 (N_11630,N_10086,N_10593);
nand U11631 (N_11631,N_9906,N_10571);
xor U11632 (N_11632,N_9747,N_9859);
or U11633 (N_11633,N_10431,N_10318);
and U11634 (N_11634,N_10618,N_9768);
and U11635 (N_11635,N_9665,N_10225);
xor U11636 (N_11636,N_10140,N_10051);
nor U11637 (N_11637,N_10430,N_10022);
and U11638 (N_11638,N_10272,N_9706);
nand U11639 (N_11639,N_10305,N_9950);
or U11640 (N_11640,N_10333,N_9814);
or U11641 (N_11641,N_9757,N_10095);
and U11642 (N_11642,N_9799,N_9975);
and U11643 (N_11643,N_10252,N_10141);
or U11644 (N_11644,N_10410,N_10478);
nor U11645 (N_11645,N_9857,N_9786);
nor U11646 (N_11646,N_9765,N_10385);
xor U11647 (N_11647,N_10769,N_10063);
nand U11648 (N_11648,N_10641,N_10034);
nand U11649 (N_11649,N_9924,N_10197);
nand U11650 (N_11650,N_9850,N_9753);
and U11651 (N_11651,N_10468,N_10091);
xor U11652 (N_11652,N_10589,N_9761);
or U11653 (N_11653,N_9920,N_9963);
xor U11654 (N_11654,N_10710,N_10524);
xnor U11655 (N_11655,N_9862,N_9658);
nand U11656 (N_11656,N_9702,N_9621);
xnor U11657 (N_11657,N_9881,N_10639);
nor U11658 (N_11658,N_9638,N_10288);
nand U11659 (N_11659,N_10176,N_10061);
and U11660 (N_11660,N_10514,N_10083);
nor U11661 (N_11661,N_10289,N_10428);
nor U11662 (N_11662,N_10259,N_10275);
or U11663 (N_11663,N_10656,N_10580);
nor U11664 (N_11664,N_9859,N_10463);
xor U11665 (N_11665,N_10695,N_10329);
or U11666 (N_11666,N_9997,N_9749);
and U11667 (N_11667,N_10044,N_9686);
xnor U11668 (N_11668,N_10690,N_10793);
and U11669 (N_11669,N_10190,N_10415);
nand U11670 (N_11670,N_10348,N_10607);
nand U11671 (N_11671,N_10053,N_10258);
and U11672 (N_11672,N_10077,N_9893);
nor U11673 (N_11673,N_9982,N_10425);
nor U11674 (N_11674,N_9667,N_10384);
nor U11675 (N_11675,N_10140,N_10167);
or U11676 (N_11676,N_9627,N_10785);
or U11677 (N_11677,N_9787,N_10373);
xnor U11678 (N_11678,N_9922,N_10686);
nand U11679 (N_11679,N_9636,N_10215);
and U11680 (N_11680,N_9709,N_9711);
nor U11681 (N_11681,N_10692,N_10182);
and U11682 (N_11682,N_10625,N_10226);
nand U11683 (N_11683,N_10522,N_9992);
or U11684 (N_11684,N_10570,N_9986);
nand U11685 (N_11685,N_10088,N_10682);
nor U11686 (N_11686,N_10676,N_9689);
and U11687 (N_11687,N_10377,N_10111);
and U11688 (N_11688,N_10355,N_10581);
nand U11689 (N_11689,N_10490,N_10274);
or U11690 (N_11690,N_10357,N_10307);
xnor U11691 (N_11691,N_10271,N_9790);
nor U11692 (N_11692,N_9984,N_9613);
and U11693 (N_11693,N_9717,N_10608);
nor U11694 (N_11694,N_10587,N_9826);
or U11695 (N_11695,N_9781,N_9757);
xnor U11696 (N_11696,N_10286,N_10703);
nor U11697 (N_11697,N_9936,N_10115);
xor U11698 (N_11698,N_9930,N_10200);
nand U11699 (N_11699,N_10023,N_10318);
nor U11700 (N_11700,N_9739,N_9951);
xnor U11701 (N_11701,N_10535,N_10040);
and U11702 (N_11702,N_9811,N_9993);
and U11703 (N_11703,N_9654,N_9607);
xor U11704 (N_11704,N_10757,N_10583);
and U11705 (N_11705,N_10694,N_10109);
xnor U11706 (N_11706,N_10071,N_10630);
and U11707 (N_11707,N_10534,N_10537);
nand U11708 (N_11708,N_10543,N_9893);
nand U11709 (N_11709,N_10078,N_10348);
nor U11710 (N_11710,N_10418,N_9895);
and U11711 (N_11711,N_10547,N_10266);
xor U11712 (N_11712,N_10071,N_10687);
or U11713 (N_11713,N_9646,N_10235);
nand U11714 (N_11714,N_10164,N_10609);
and U11715 (N_11715,N_10136,N_10624);
or U11716 (N_11716,N_10081,N_10414);
xnor U11717 (N_11717,N_10550,N_10652);
and U11718 (N_11718,N_9718,N_9623);
or U11719 (N_11719,N_10691,N_10494);
and U11720 (N_11720,N_9903,N_10574);
or U11721 (N_11721,N_9641,N_10713);
or U11722 (N_11722,N_10223,N_9930);
xnor U11723 (N_11723,N_9718,N_9716);
nand U11724 (N_11724,N_10654,N_10334);
or U11725 (N_11725,N_10259,N_10723);
and U11726 (N_11726,N_10402,N_10084);
and U11727 (N_11727,N_10178,N_10007);
nor U11728 (N_11728,N_9905,N_10446);
nand U11729 (N_11729,N_10667,N_10723);
and U11730 (N_11730,N_10364,N_10730);
nor U11731 (N_11731,N_9913,N_10200);
xor U11732 (N_11732,N_10252,N_10348);
xnor U11733 (N_11733,N_10313,N_10548);
nor U11734 (N_11734,N_10560,N_10024);
xnor U11735 (N_11735,N_10462,N_10017);
xor U11736 (N_11736,N_10033,N_10123);
nand U11737 (N_11737,N_10789,N_9675);
or U11738 (N_11738,N_10748,N_9662);
nand U11739 (N_11739,N_9848,N_10729);
nor U11740 (N_11740,N_10301,N_9850);
nand U11741 (N_11741,N_10217,N_10325);
xor U11742 (N_11742,N_10350,N_9652);
nand U11743 (N_11743,N_10329,N_10093);
or U11744 (N_11744,N_10302,N_10628);
and U11745 (N_11745,N_9758,N_9836);
xnor U11746 (N_11746,N_10243,N_10595);
or U11747 (N_11747,N_9619,N_9998);
and U11748 (N_11748,N_9767,N_10076);
nor U11749 (N_11749,N_10404,N_10018);
or U11750 (N_11750,N_10501,N_10693);
xnor U11751 (N_11751,N_9773,N_10754);
xnor U11752 (N_11752,N_9630,N_10471);
or U11753 (N_11753,N_10694,N_9877);
nand U11754 (N_11754,N_9696,N_9641);
xor U11755 (N_11755,N_10299,N_9812);
nand U11756 (N_11756,N_10257,N_10021);
xnor U11757 (N_11757,N_10107,N_10691);
nor U11758 (N_11758,N_9810,N_10574);
and U11759 (N_11759,N_10679,N_10329);
or U11760 (N_11760,N_10475,N_9981);
and U11761 (N_11761,N_10465,N_9635);
nor U11762 (N_11762,N_10794,N_10013);
nor U11763 (N_11763,N_10742,N_9617);
nor U11764 (N_11764,N_10276,N_10193);
and U11765 (N_11765,N_10721,N_10579);
nor U11766 (N_11766,N_10687,N_10465);
nor U11767 (N_11767,N_9934,N_10125);
nor U11768 (N_11768,N_10116,N_10289);
and U11769 (N_11769,N_10497,N_9610);
nand U11770 (N_11770,N_9878,N_10530);
and U11771 (N_11771,N_10222,N_10595);
nand U11772 (N_11772,N_9873,N_9876);
xor U11773 (N_11773,N_10773,N_10577);
nor U11774 (N_11774,N_10101,N_10718);
and U11775 (N_11775,N_10400,N_9624);
or U11776 (N_11776,N_10375,N_10123);
nor U11777 (N_11777,N_9935,N_9755);
nand U11778 (N_11778,N_10196,N_10093);
and U11779 (N_11779,N_9977,N_9855);
xor U11780 (N_11780,N_10391,N_10765);
nand U11781 (N_11781,N_10657,N_10086);
or U11782 (N_11782,N_10272,N_9799);
or U11783 (N_11783,N_10482,N_10452);
nor U11784 (N_11784,N_10709,N_10326);
nand U11785 (N_11785,N_9953,N_10582);
and U11786 (N_11786,N_9751,N_10736);
nor U11787 (N_11787,N_10267,N_10606);
nand U11788 (N_11788,N_10313,N_9618);
xnor U11789 (N_11789,N_10448,N_10462);
and U11790 (N_11790,N_9965,N_9970);
nor U11791 (N_11791,N_10343,N_10488);
xnor U11792 (N_11792,N_9785,N_9740);
nor U11793 (N_11793,N_10006,N_10202);
or U11794 (N_11794,N_10269,N_9966);
and U11795 (N_11795,N_10327,N_10259);
nor U11796 (N_11796,N_9743,N_9834);
xor U11797 (N_11797,N_9607,N_9980);
or U11798 (N_11798,N_9786,N_10387);
or U11799 (N_11799,N_9607,N_10458);
nor U11800 (N_11800,N_10436,N_10653);
xnor U11801 (N_11801,N_10540,N_10179);
and U11802 (N_11802,N_10633,N_10641);
and U11803 (N_11803,N_10415,N_10563);
and U11804 (N_11804,N_10048,N_10241);
xor U11805 (N_11805,N_10224,N_9791);
xnor U11806 (N_11806,N_9764,N_10058);
nor U11807 (N_11807,N_9949,N_10706);
nand U11808 (N_11808,N_10470,N_9887);
xor U11809 (N_11809,N_9882,N_10425);
and U11810 (N_11810,N_10274,N_10256);
nand U11811 (N_11811,N_9949,N_10290);
nand U11812 (N_11812,N_10390,N_10284);
or U11813 (N_11813,N_10201,N_10439);
or U11814 (N_11814,N_10084,N_10011);
nand U11815 (N_11815,N_10139,N_9877);
xor U11816 (N_11816,N_10423,N_9650);
nor U11817 (N_11817,N_10126,N_10679);
xnor U11818 (N_11818,N_10556,N_9931);
nand U11819 (N_11819,N_10158,N_9804);
nand U11820 (N_11820,N_10112,N_10781);
xnor U11821 (N_11821,N_10419,N_9674);
nor U11822 (N_11822,N_10322,N_10165);
nor U11823 (N_11823,N_10437,N_10688);
nor U11824 (N_11824,N_10472,N_9728);
xnor U11825 (N_11825,N_10621,N_10002);
and U11826 (N_11826,N_9857,N_10488);
nor U11827 (N_11827,N_9905,N_10500);
and U11828 (N_11828,N_9734,N_9883);
nand U11829 (N_11829,N_10783,N_9840);
nor U11830 (N_11830,N_10716,N_10011);
xnor U11831 (N_11831,N_9600,N_9615);
xor U11832 (N_11832,N_10306,N_10451);
and U11833 (N_11833,N_10082,N_10083);
nor U11834 (N_11834,N_10001,N_10002);
xor U11835 (N_11835,N_10785,N_9783);
xnor U11836 (N_11836,N_10165,N_9917);
nand U11837 (N_11837,N_10160,N_9726);
nor U11838 (N_11838,N_10392,N_10520);
xnor U11839 (N_11839,N_10079,N_9710);
and U11840 (N_11840,N_10661,N_10144);
nand U11841 (N_11841,N_9833,N_10499);
xor U11842 (N_11842,N_10550,N_9636);
or U11843 (N_11843,N_10496,N_10571);
xor U11844 (N_11844,N_9641,N_9965);
or U11845 (N_11845,N_9634,N_10559);
nor U11846 (N_11846,N_10726,N_10637);
nor U11847 (N_11847,N_10227,N_10154);
and U11848 (N_11848,N_10686,N_10169);
or U11849 (N_11849,N_10770,N_10173);
xor U11850 (N_11850,N_10538,N_10741);
xor U11851 (N_11851,N_10044,N_10653);
nand U11852 (N_11852,N_10122,N_9844);
or U11853 (N_11853,N_10361,N_9901);
or U11854 (N_11854,N_9796,N_9803);
nand U11855 (N_11855,N_10232,N_10394);
or U11856 (N_11856,N_10498,N_9846);
nor U11857 (N_11857,N_9816,N_9943);
nor U11858 (N_11858,N_10172,N_9992);
and U11859 (N_11859,N_10434,N_9748);
nor U11860 (N_11860,N_10571,N_10346);
and U11861 (N_11861,N_10596,N_10206);
xor U11862 (N_11862,N_10744,N_10593);
or U11863 (N_11863,N_9694,N_9806);
nor U11864 (N_11864,N_10550,N_10736);
nand U11865 (N_11865,N_10344,N_9926);
or U11866 (N_11866,N_10687,N_9793);
xor U11867 (N_11867,N_9698,N_10653);
nand U11868 (N_11868,N_9753,N_10327);
xnor U11869 (N_11869,N_10656,N_10629);
xor U11870 (N_11870,N_9925,N_10361);
nand U11871 (N_11871,N_10120,N_10545);
or U11872 (N_11872,N_10317,N_10255);
and U11873 (N_11873,N_10794,N_10014);
xnor U11874 (N_11874,N_9654,N_9957);
xor U11875 (N_11875,N_10496,N_10798);
or U11876 (N_11876,N_9774,N_10706);
xnor U11877 (N_11877,N_10774,N_10059);
nand U11878 (N_11878,N_10010,N_10452);
nor U11879 (N_11879,N_10459,N_10125);
and U11880 (N_11880,N_10312,N_9790);
nor U11881 (N_11881,N_10756,N_10336);
xor U11882 (N_11882,N_10742,N_9798);
or U11883 (N_11883,N_9678,N_9854);
and U11884 (N_11884,N_9907,N_9644);
nor U11885 (N_11885,N_10012,N_9743);
or U11886 (N_11886,N_10294,N_9806);
xor U11887 (N_11887,N_9827,N_10212);
nand U11888 (N_11888,N_10728,N_10185);
nand U11889 (N_11889,N_10221,N_10436);
and U11890 (N_11890,N_9774,N_10001);
or U11891 (N_11891,N_10273,N_10550);
or U11892 (N_11892,N_10332,N_10137);
nor U11893 (N_11893,N_10776,N_10054);
nand U11894 (N_11894,N_10283,N_9893);
xnor U11895 (N_11895,N_10406,N_9970);
or U11896 (N_11896,N_10730,N_10118);
nand U11897 (N_11897,N_9654,N_10575);
nand U11898 (N_11898,N_10030,N_10492);
xnor U11899 (N_11899,N_9848,N_9755);
xnor U11900 (N_11900,N_10630,N_10136);
nand U11901 (N_11901,N_9642,N_10761);
nand U11902 (N_11902,N_10508,N_9917);
or U11903 (N_11903,N_10025,N_10081);
xnor U11904 (N_11904,N_9919,N_10354);
nor U11905 (N_11905,N_10214,N_10596);
or U11906 (N_11906,N_9831,N_10458);
or U11907 (N_11907,N_10795,N_10427);
nor U11908 (N_11908,N_9812,N_10724);
nand U11909 (N_11909,N_10274,N_9600);
or U11910 (N_11910,N_10024,N_10309);
nor U11911 (N_11911,N_9985,N_9764);
xor U11912 (N_11912,N_10103,N_10543);
nor U11913 (N_11913,N_10774,N_10473);
xor U11914 (N_11914,N_10655,N_9772);
nor U11915 (N_11915,N_9952,N_10705);
and U11916 (N_11916,N_10491,N_10428);
xnor U11917 (N_11917,N_10266,N_10623);
nand U11918 (N_11918,N_10722,N_10472);
xor U11919 (N_11919,N_9807,N_10722);
nor U11920 (N_11920,N_9905,N_10448);
or U11921 (N_11921,N_10493,N_9649);
nor U11922 (N_11922,N_10368,N_9796);
xor U11923 (N_11923,N_10235,N_9988);
nor U11924 (N_11924,N_10175,N_9929);
or U11925 (N_11925,N_9875,N_9923);
nor U11926 (N_11926,N_10116,N_10566);
or U11927 (N_11927,N_10339,N_10709);
and U11928 (N_11928,N_10041,N_9824);
or U11929 (N_11929,N_10778,N_10594);
nor U11930 (N_11930,N_9880,N_10142);
and U11931 (N_11931,N_10328,N_10244);
and U11932 (N_11932,N_10416,N_10345);
xnor U11933 (N_11933,N_10144,N_9807);
or U11934 (N_11934,N_10287,N_10305);
nand U11935 (N_11935,N_10232,N_10357);
and U11936 (N_11936,N_10249,N_10489);
or U11937 (N_11937,N_9641,N_10419);
and U11938 (N_11938,N_10689,N_10764);
and U11939 (N_11939,N_10526,N_10002);
nand U11940 (N_11940,N_10188,N_10348);
xor U11941 (N_11941,N_10213,N_10226);
xnor U11942 (N_11942,N_9645,N_10302);
nor U11943 (N_11943,N_10533,N_10230);
or U11944 (N_11944,N_10452,N_10254);
nand U11945 (N_11945,N_9651,N_10793);
nor U11946 (N_11946,N_10181,N_9847);
or U11947 (N_11947,N_9665,N_9947);
nand U11948 (N_11948,N_10757,N_10436);
nand U11949 (N_11949,N_10381,N_10430);
xnor U11950 (N_11950,N_9940,N_10027);
nor U11951 (N_11951,N_9964,N_10741);
and U11952 (N_11952,N_10406,N_9807);
nand U11953 (N_11953,N_10351,N_9984);
nor U11954 (N_11954,N_10301,N_10564);
nand U11955 (N_11955,N_10516,N_10298);
xor U11956 (N_11956,N_10199,N_10462);
or U11957 (N_11957,N_9900,N_9774);
or U11958 (N_11958,N_10621,N_10579);
nand U11959 (N_11959,N_10707,N_10110);
nor U11960 (N_11960,N_10073,N_10117);
nor U11961 (N_11961,N_10575,N_10272);
and U11962 (N_11962,N_10672,N_10788);
xnor U11963 (N_11963,N_10715,N_10379);
xnor U11964 (N_11964,N_10258,N_10781);
nand U11965 (N_11965,N_10593,N_10307);
and U11966 (N_11966,N_10097,N_10525);
or U11967 (N_11967,N_10099,N_10776);
nor U11968 (N_11968,N_10346,N_10547);
or U11969 (N_11969,N_10153,N_10095);
nor U11970 (N_11970,N_10518,N_10449);
or U11971 (N_11971,N_9860,N_9726);
xnor U11972 (N_11972,N_9956,N_10693);
xnor U11973 (N_11973,N_10131,N_10281);
or U11974 (N_11974,N_10335,N_10138);
and U11975 (N_11975,N_10475,N_10679);
nor U11976 (N_11976,N_9822,N_9878);
xor U11977 (N_11977,N_10293,N_10666);
or U11978 (N_11978,N_10128,N_10002);
nor U11979 (N_11979,N_10624,N_9981);
or U11980 (N_11980,N_10645,N_10515);
nand U11981 (N_11981,N_9867,N_10437);
nand U11982 (N_11982,N_10585,N_10014);
nand U11983 (N_11983,N_10620,N_10512);
nor U11984 (N_11984,N_10246,N_9935);
nor U11985 (N_11985,N_10419,N_10193);
or U11986 (N_11986,N_9953,N_9812);
xnor U11987 (N_11987,N_10254,N_9986);
nor U11988 (N_11988,N_10566,N_10660);
nand U11989 (N_11989,N_10409,N_9889);
or U11990 (N_11990,N_10085,N_10459);
nor U11991 (N_11991,N_10467,N_9794);
nor U11992 (N_11992,N_10239,N_10573);
nand U11993 (N_11993,N_10478,N_10778);
nand U11994 (N_11994,N_9977,N_10058);
and U11995 (N_11995,N_10067,N_9717);
or U11996 (N_11996,N_10358,N_9682);
and U11997 (N_11997,N_10555,N_9663);
xor U11998 (N_11998,N_10002,N_9621);
xor U11999 (N_11999,N_10754,N_10176);
nand U12000 (N_12000,N_10957,N_11770);
nand U12001 (N_12001,N_10807,N_11384);
xor U12002 (N_12002,N_11662,N_11475);
or U12003 (N_12003,N_11661,N_10922);
nand U12004 (N_12004,N_11560,N_11516);
xor U12005 (N_12005,N_11272,N_10916);
xor U12006 (N_12006,N_11822,N_10900);
or U12007 (N_12007,N_11428,N_11613);
and U12008 (N_12008,N_11217,N_11978);
and U12009 (N_12009,N_11861,N_10869);
nor U12010 (N_12010,N_11216,N_11983);
xor U12011 (N_12011,N_11909,N_11769);
nand U12012 (N_12012,N_11860,N_11300);
nand U12013 (N_12013,N_10989,N_11830);
or U12014 (N_12014,N_10810,N_11468);
xnor U12015 (N_12015,N_10884,N_11893);
nand U12016 (N_12016,N_10819,N_11934);
nor U12017 (N_12017,N_11323,N_11365);
nor U12018 (N_12018,N_11891,N_11021);
xnor U12019 (N_12019,N_11695,N_11916);
nand U12020 (N_12020,N_11878,N_11454);
xor U12021 (N_12021,N_11673,N_11357);
nor U12022 (N_12022,N_11582,N_11678);
and U12023 (N_12023,N_11201,N_11172);
or U12024 (N_12024,N_11199,N_11832);
xnor U12025 (N_12025,N_11206,N_10947);
or U12026 (N_12026,N_11026,N_11815);
xnor U12027 (N_12027,N_11461,N_11786);
or U12028 (N_12028,N_11726,N_11898);
or U12029 (N_12029,N_11380,N_11858);
or U12030 (N_12030,N_11131,N_11594);
xnor U12031 (N_12031,N_11403,N_11095);
nor U12032 (N_12032,N_11553,N_11517);
nor U12033 (N_12033,N_10972,N_11449);
xor U12034 (N_12034,N_11746,N_11006);
nand U12035 (N_12035,N_10964,N_11321);
and U12036 (N_12036,N_11143,N_10962);
xor U12037 (N_12037,N_11163,N_11033);
nor U12038 (N_12038,N_11570,N_11540);
or U12039 (N_12039,N_11352,N_11165);
nor U12040 (N_12040,N_11686,N_11807);
nand U12041 (N_12041,N_10953,N_11839);
nand U12042 (N_12042,N_10968,N_11344);
or U12043 (N_12043,N_11486,N_11975);
and U12044 (N_12044,N_10805,N_10835);
and U12045 (N_12045,N_11181,N_11509);
or U12046 (N_12046,N_11631,N_11939);
xnor U12047 (N_12047,N_11132,N_11953);
or U12048 (N_12048,N_11342,N_11001);
nor U12049 (N_12049,N_11338,N_10847);
or U12050 (N_12050,N_10848,N_11957);
nand U12051 (N_12051,N_11521,N_11927);
or U12052 (N_12052,N_11652,N_10843);
nand U12053 (N_12053,N_11787,N_11680);
nand U12054 (N_12054,N_11888,N_10948);
xor U12055 (N_12055,N_11283,N_11932);
and U12056 (N_12056,N_11371,N_11489);
xor U12057 (N_12057,N_11402,N_11664);
xnor U12058 (N_12058,N_11361,N_10861);
and U12059 (N_12059,N_11298,N_11079);
nand U12060 (N_12060,N_11732,N_11801);
or U12061 (N_12061,N_11081,N_11471);
xor U12062 (N_12062,N_11022,N_11179);
nor U12063 (N_12063,N_11326,N_11968);
nand U12064 (N_12064,N_11353,N_11218);
or U12065 (N_12065,N_11847,N_11121);
and U12066 (N_12066,N_11423,N_11420);
xnor U12067 (N_12067,N_11134,N_11571);
or U12068 (N_12068,N_11077,N_10885);
xnor U12069 (N_12069,N_11349,N_11955);
or U12070 (N_12070,N_11929,N_11937);
nor U12071 (N_12071,N_11682,N_11679);
or U12072 (N_12072,N_11820,N_11119);
and U12073 (N_12073,N_11389,N_11914);
xor U12074 (N_12074,N_10841,N_10971);
and U12075 (N_12075,N_10886,N_11270);
or U12076 (N_12076,N_11392,N_11040);
nor U12077 (N_12077,N_11474,N_11854);
and U12078 (N_12078,N_10894,N_11938);
or U12079 (N_12079,N_11433,N_11487);
nand U12080 (N_12080,N_11379,N_11419);
and U12081 (N_12081,N_10907,N_10980);
nand U12082 (N_12082,N_11911,N_11717);
xnor U12083 (N_12083,N_11035,N_11176);
or U12084 (N_12084,N_11066,N_11778);
xnor U12085 (N_12085,N_11625,N_10936);
nand U12086 (N_12086,N_11166,N_11597);
and U12087 (N_12087,N_11834,N_11772);
or U12088 (N_12088,N_11109,N_11180);
xor U12089 (N_12089,N_10897,N_11824);
nand U12090 (N_12090,N_10902,N_10914);
nand U12091 (N_12091,N_10820,N_11354);
and U12092 (N_12092,N_10816,N_11332);
nor U12093 (N_12093,N_11325,N_11090);
xnor U12094 (N_12094,N_11434,N_11260);
nand U12095 (N_12095,N_11643,N_11826);
nand U12096 (N_12096,N_11532,N_10906);
or U12097 (N_12097,N_11991,N_11388);
and U12098 (N_12098,N_11562,N_11897);
or U12099 (N_12099,N_11480,N_11671);
xnor U12100 (N_12100,N_11313,N_11439);
nand U12101 (N_12101,N_11065,N_11093);
nand U12102 (N_12102,N_11627,N_11262);
nor U12103 (N_12103,N_10926,N_11641);
xnor U12104 (N_12104,N_11064,N_11327);
nand U12105 (N_12105,N_11687,N_10842);
nor U12106 (N_12106,N_11507,N_11405);
nor U12107 (N_12107,N_11398,N_11443);
nand U12108 (N_12108,N_11621,N_11092);
or U12109 (N_12109,N_11872,N_11237);
nor U12110 (N_12110,N_11923,N_11282);
nand U12111 (N_12111,N_11842,N_11039);
or U12112 (N_12112,N_11114,N_10988);
nor U12113 (N_12113,N_10998,N_11246);
nor U12114 (N_12114,N_10834,N_11568);
nor U12115 (N_12115,N_11611,N_11674);
nor U12116 (N_12116,N_11644,N_11779);
nand U12117 (N_12117,N_11817,N_11367);
and U12118 (N_12118,N_11551,N_10939);
nand U12119 (N_12119,N_11214,N_11950);
or U12120 (N_12120,N_11899,N_11989);
and U12121 (N_12121,N_11730,N_11299);
or U12122 (N_12122,N_11624,N_11152);
or U12123 (N_12123,N_11122,N_11783);
nor U12124 (N_12124,N_10875,N_11638);
nand U12125 (N_12125,N_11972,N_10977);
nand U12126 (N_12126,N_11045,N_11685);
xor U12127 (N_12127,N_11966,N_11767);
nor U12128 (N_12128,N_11233,N_11124);
xnor U12129 (N_12129,N_11426,N_11581);
nand U12130 (N_12130,N_11574,N_11034);
nor U12131 (N_12131,N_11104,N_11118);
nor U12132 (N_12132,N_11917,N_11951);
xnor U12133 (N_12133,N_11618,N_11210);
nor U12134 (N_12134,N_11054,N_11383);
or U12135 (N_12135,N_11413,N_11564);
nor U12136 (N_12136,N_10893,N_11969);
nor U12137 (N_12137,N_11016,N_11205);
nand U12138 (N_12138,N_11812,N_11762);
nand U12139 (N_12139,N_11760,N_10932);
and U12140 (N_12140,N_10942,N_11544);
and U12141 (N_12141,N_11608,N_10995);
nor U12142 (N_12142,N_11295,N_11215);
nand U12143 (N_12143,N_11761,N_11196);
and U12144 (N_12144,N_11515,N_11478);
xor U12145 (N_12145,N_11019,N_11345);
or U12146 (N_12146,N_11491,N_11438);
or U12147 (N_12147,N_11773,N_11514);
or U12148 (N_12148,N_11409,N_10908);
or U12149 (N_12149,N_11844,N_11575);
or U12150 (N_12150,N_11543,N_11069);
nor U12151 (N_12151,N_11788,N_11785);
nand U12152 (N_12152,N_11835,N_11829);
nor U12153 (N_12153,N_11460,N_10960);
nor U12154 (N_12154,N_11852,N_11241);
and U12155 (N_12155,N_11418,N_11235);
xor U12156 (N_12156,N_11038,N_11943);
xor U12157 (N_12157,N_11444,N_11137);
or U12158 (N_12158,N_11895,N_11286);
xnor U12159 (N_12159,N_10923,N_11138);
nor U12160 (N_12160,N_11536,N_11002);
xor U12161 (N_12161,N_11973,N_11942);
and U12162 (N_12162,N_11267,N_11567);
xnor U12163 (N_12163,N_11513,N_11111);
nor U12164 (N_12164,N_11525,N_11312);
and U12165 (N_12165,N_11187,N_11191);
nor U12166 (N_12166,N_11195,N_11289);
or U12167 (N_12167,N_11459,N_11322);
and U12168 (N_12168,N_11372,N_11947);
nand U12169 (N_12169,N_11646,N_11275);
xor U12170 (N_12170,N_11153,N_11430);
nand U12171 (N_12171,N_11976,N_11739);
xor U12172 (N_12172,N_11482,N_10825);
nor U12173 (N_12173,N_11078,N_11903);
and U12174 (N_12174,N_11936,N_11605);
and U12175 (N_12175,N_11068,N_11670);
and U12176 (N_12176,N_11333,N_11744);
xnor U12177 (N_12177,N_11424,N_11743);
and U12178 (N_12178,N_10991,N_11724);
nand U12179 (N_12179,N_11635,N_10876);
nor U12180 (N_12180,N_11971,N_10951);
and U12181 (N_12181,N_11960,N_11802);
nor U12182 (N_12182,N_11676,N_11098);
nor U12183 (N_12183,N_11590,N_11534);
nand U12184 (N_12184,N_11168,N_11223);
nor U12185 (N_12185,N_10822,N_11253);
nor U12186 (N_12186,N_11490,N_11974);
and U12187 (N_12187,N_11130,N_11264);
nand U12188 (N_12188,N_11320,N_11502);
or U12189 (N_12189,N_11127,N_11859);
and U12190 (N_12190,N_10896,N_11467);
xor U12191 (N_12191,N_11416,N_11873);
or U12192 (N_12192,N_11051,N_11711);
nand U12193 (N_12193,N_11539,N_10804);
nand U12194 (N_12194,N_10915,N_11626);
nor U12195 (N_12195,N_11297,N_10872);
xor U12196 (N_12196,N_11258,N_11811);
xnor U12197 (N_12197,N_11082,N_11393);
nand U12198 (N_12198,N_11836,N_11797);
or U12199 (N_12199,N_10992,N_11042);
nor U12200 (N_12200,N_10974,N_11465);
nor U12201 (N_12201,N_11658,N_10880);
or U12202 (N_12202,N_11378,N_11058);
nor U12203 (N_12203,N_11274,N_11287);
and U12204 (N_12204,N_11701,N_11579);
or U12205 (N_12205,N_11675,N_11554);
nand U12206 (N_12206,N_11410,N_11672);
and U12207 (N_12207,N_11018,N_11875);
nand U12208 (N_12208,N_11741,N_10878);
xnor U12209 (N_12209,N_11220,N_10899);
and U12210 (N_12210,N_10961,N_11339);
and U12211 (N_12211,N_11782,N_11310);
nand U12212 (N_12212,N_11883,N_11913);
nor U12213 (N_12213,N_11200,N_10818);
nand U12214 (N_12214,N_11504,N_11108);
and U12215 (N_12215,N_11905,N_11228);
nor U12216 (N_12216,N_11928,N_11716);
nand U12217 (N_12217,N_11466,N_10905);
xnor U12218 (N_12218,N_11161,N_11684);
and U12219 (N_12219,N_11318,N_11435);
nor U12220 (N_12220,N_11120,N_11995);
or U12221 (N_12221,N_11083,N_11585);
and U12222 (N_12222,N_11728,N_10823);
nor U12223 (N_12223,N_11655,N_11734);
nand U12224 (N_12224,N_11373,N_11303);
nor U12225 (N_12225,N_11473,N_11508);
and U12226 (N_12226,N_11007,N_11452);
xor U12227 (N_12227,N_11041,N_11128);
or U12228 (N_12228,N_11123,N_11902);
and U12229 (N_12229,N_10874,N_11948);
and U12230 (N_12230,N_11147,N_11248);
xnor U12231 (N_12231,N_11479,N_11804);
nand U12232 (N_12232,N_11979,N_11450);
nand U12233 (N_12233,N_11602,N_11369);
nor U12234 (N_12234,N_11714,N_11924);
or U12235 (N_12235,N_10803,N_11000);
nand U12236 (N_12236,N_10938,N_10853);
or U12237 (N_12237,N_10918,N_11962);
nand U12238 (N_12238,N_11387,N_11330);
xnor U12239 (N_12239,N_10845,N_11234);
nor U12240 (N_12240,N_11028,N_11591);
nor U12241 (N_12241,N_11394,N_10832);
nand U12242 (N_12242,N_10849,N_11053);
nand U12243 (N_12243,N_10935,N_11151);
and U12244 (N_12244,N_11988,N_11918);
or U12245 (N_12245,N_11453,N_11500);
or U12246 (N_12246,N_11697,N_10966);
and U12247 (N_12247,N_11926,N_11810);
and U12248 (N_12248,N_11250,N_11775);
xnor U12249 (N_12249,N_11864,N_11636);
nand U12250 (N_12250,N_11886,N_11876);
or U12251 (N_12251,N_11170,N_11519);
nor U12252 (N_12252,N_11062,N_11189);
and U12253 (N_12253,N_10913,N_11030);
xor U12254 (N_12254,N_11350,N_10865);
or U12255 (N_12255,N_10967,N_11319);
nor U12256 (N_12256,N_11238,N_11855);
nand U12257 (N_12257,N_11382,N_10944);
and U12258 (N_12258,N_11411,N_11277);
and U12259 (N_12259,N_10982,N_10840);
and U12260 (N_12260,N_10827,N_11550);
or U12261 (N_12261,N_11204,N_11110);
nand U12262 (N_12262,N_11495,N_11126);
and U12263 (N_12263,N_11073,N_11656);
and U12264 (N_12264,N_10930,N_11667);
xor U12265 (N_12265,N_11139,N_11930);
or U12266 (N_12266,N_10952,N_11055);
or U12267 (N_12267,N_11851,N_10917);
or U12268 (N_12268,N_11036,N_11247);
or U12269 (N_12269,N_11531,N_11072);
or U12270 (N_12270,N_11865,N_11524);
or U12271 (N_12271,N_11892,N_11004);
xor U12272 (N_12272,N_10839,N_11833);
and U12273 (N_12273,N_11542,N_11720);
nand U12274 (N_12274,N_11113,N_11156);
or U12275 (N_12275,N_11827,N_11399);
nor U12276 (N_12276,N_10850,N_11639);
xnor U12277 (N_12277,N_11445,N_11368);
nand U12278 (N_12278,N_11257,N_11884);
nand U12279 (N_12279,N_11376,N_11476);
nor U12280 (N_12280,N_11941,N_11010);
or U12281 (N_12281,N_10826,N_11381);
and U12282 (N_12282,N_11506,N_11406);
or U12283 (N_12283,N_11304,N_11584);
nor U12284 (N_12284,N_11343,N_11659);
or U12285 (N_12285,N_11483,N_11178);
nor U12286 (N_12286,N_11654,N_11601);
nand U12287 (N_12287,N_10950,N_11958);
nor U12288 (N_12288,N_11642,N_11651);
nor U12289 (N_12289,N_11771,N_11774);
or U12290 (N_12290,N_11900,N_10866);
nand U12291 (N_12291,N_11843,N_11186);
nand U12292 (N_12292,N_11169,N_11448);
nor U12293 (N_12293,N_11031,N_11634);
nand U12294 (N_12294,N_11512,N_11140);
nand U12295 (N_12295,N_11745,N_11391);
and U12296 (N_12296,N_11099,N_11202);
and U12297 (N_12297,N_11203,N_10846);
nor U12298 (N_12298,N_11401,N_11706);
xor U12299 (N_12299,N_11125,N_11014);
xnor U12300 (N_12300,N_11862,N_11965);
nor U12301 (N_12301,N_11457,N_11422);
xnor U12302 (N_12302,N_11451,N_10984);
xnor U12303 (N_12303,N_11414,N_11252);
and U12304 (N_12304,N_11725,N_11107);
and U12305 (N_12305,N_11084,N_11784);
or U12306 (N_12306,N_11141,N_11145);
nand U12307 (N_12307,N_10924,N_10931);
and U12308 (N_12308,N_11742,N_10859);
or U12309 (N_12309,N_10856,N_11647);
xnor U12310 (N_12310,N_10955,N_11425);
nand U12311 (N_12311,N_11650,N_11224);
or U12312 (N_12312,N_11341,N_11492);
xor U12313 (N_12313,N_11805,N_11155);
or U12314 (N_12314,N_11261,N_11528);
or U12315 (N_12315,N_11809,N_11185);
xor U12316 (N_12316,N_11046,N_11446);
nand U12317 (N_12317,N_11366,N_11669);
xor U12318 (N_12318,N_11870,N_11464);
nand U12319 (N_12319,N_11100,N_10892);
and U12320 (N_12320,N_11945,N_11329);
or U12321 (N_12321,N_11269,N_11292);
nand U12322 (N_12322,N_11691,N_11700);
nor U12323 (N_12323,N_10978,N_11211);
nor U12324 (N_12324,N_11593,N_10873);
xnor U12325 (N_12325,N_11059,N_11219);
and U12326 (N_12326,N_11091,N_11821);
xnor U12327 (N_12327,N_11102,N_11183);
nor U12328 (N_12328,N_11857,N_11793);
nand U12329 (N_12329,N_11708,N_11301);
and U12330 (N_12330,N_11094,N_11800);
nand U12331 (N_12331,N_11885,N_11290);
nand U12332 (N_12332,N_11458,N_11472);
and U12333 (N_12333,N_11236,N_10946);
and U12334 (N_12334,N_10813,N_11606);
nand U12335 (N_12335,N_11421,N_11400);
nor U12336 (N_12336,N_10986,N_11133);
xor U12337 (N_12337,N_11395,N_11044);
or U12338 (N_12338,N_11335,N_10985);
or U12339 (N_12339,N_10800,N_10976);
nand U12340 (N_12340,N_10860,N_11752);
and U12341 (N_12341,N_10844,N_11721);
nand U12342 (N_12342,N_11751,N_11047);
xnor U12343 (N_12343,N_11546,N_11037);
xnor U12344 (N_12344,N_11681,N_11566);
or U12345 (N_12345,N_11756,N_11755);
nor U12346 (N_12346,N_11148,N_11436);
or U12347 (N_12347,N_11221,N_11025);
or U12348 (N_12348,N_11154,N_11075);
or U12349 (N_12349,N_11008,N_10882);
xor U12350 (N_12350,N_10870,N_11529);
nand U12351 (N_12351,N_10994,N_10837);
nor U12352 (N_12352,N_11136,N_11177);
nor U12353 (N_12353,N_10997,N_11922);
nor U12354 (N_12354,N_11017,N_11629);
and U12355 (N_12355,N_11432,N_11694);
nand U12356 (N_12356,N_11919,N_10969);
or U12357 (N_12357,N_11986,N_11530);
nand U12358 (N_12358,N_11868,N_11085);
nand U12359 (N_12359,N_11408,N_11690);
or U12360 (N_12360,N_11526,N_11023);
or U12361 (N_12361,N_11846,N_11816);
and U12362 (N_12362,N_11912,N_11921);
or U12363 (N_12363,N_11496,N_11254);
or U12364 (N_12364,N_11729,N_10979);
or U12365 (N_12365,N_11276,N_10981);
and U12366 (N_12366,N_11780,N_11970);
xnor U12367 (N_12367,N_11964,N_10975);
xnor U12368 (N_12368,N_11493,N_11348);
xor U12369 (N_12369,N_11230,N_11867);
nor U12370 (N_12370,N_11285,N_10928);
xor U12371 (N_12371,N_11296,N_11803);
or U12372 (N_12372,N_11280,N_11523);
nor U12373 (N_12373,N_11628,N_11441);
or U12374 (N_12374,N_11781,N_11129);
xor U12375 (N_12375,N_11162,N_11887);
or U12376 (N_12376,N_11209,N_11731);
nand U12377 (N_12377,N_11555,N_11599);
nor U12378 (N_12378,N_11715,N_11190);
nand U12379 (N_12379,N_11198,N_10815);
or U12380 (N_12380,N_11896,N_11748);
nor U12381 (N_12381,N_10943,N_10817);
xor U12382 (N_12382,N_11710,N_11837);
or U12383 (N_12383,N_10887,N_11316);
xor U12384 (N_12384,N_10883,N_10811);
nand U12385 (N_12385,N_11407,N_11112);
or U12386 (N_12386,N_11841,N_11164);
nand U12387 (N_12387,N_11990,N_10831);
or U12388 (N_12388,N_11340,N_10927);
xnor U12389 (N_12389,N_10806,N_11719);
or U12390 (N_12390,N_11245,N_11749);
xor U12391 (N_12391,N_11279,N_11317);
and U12392 (N_12392,N_10921,N_11556);
xor U12393 (N_12393,N_11356,N_11825);
or U12394 (N_12394,N_11535,N_11364);
or U12395 (N_12395,N_11222,N_11309);
nor U12396 (N_12396,N_11533,N_10801);
nor U12397 (N_12397,N_11577,N_11753);
nand U12398 (N_12398,N_11565,N_10901);
or U12399 (N_12399,N_11935,N_11616);
and U12400 (N_12400,N_11984,N_11906);
xnor U12401 (N_12401,N_11231,N_11607);
or U12402 (N_12402,N_10836,N_11522);
or U12403 (N_12403,N_11548,N_11374);
and U12404 (N_12404,N_11076,N_11735);
or U12405 (N_12405,N_11754,N_11609);
nand U12406 (N_12406,N_11144,N_11703);
and U12407 (N_12407,N_11281,N_11808);
and U12408 (N_12408,N_11011,N_11657);
xor U12409 (N_12409,N_11184,N_11707);
and U12410 (N_12410,N_11889,N_11510);
or U12411 (N_12411,N_11175,N_11881);
nor U12412 (N_12412,N_11386,N_10934);
nor U12413 (N_12413,N_11256,N_11890);
xnor U12414 (N_12414,N_11346,N_10987);
xor U12415 (N_12415,N_11307,N_11712);
or U12416 (N_12416,N_11985,N_11996);
nor U12417 (N_12417,N_11167,N_11159);
and U12418 (N_12418,N_11484,N_11640);
and U12419 (N_12419,N_11397,N_11666);
or U12420 (N_12420,N_11576,N_11946);
xnor U12421 (N_12421,N_11265,N_11956);
nor U12422 (N_12422,N_11470,N_11765);
and U12423 (N_12423,N_11158,N_11251);
xor U12424 (N_12424,N_11561,N_11879);
nor U12425 (N_12425,N_11853,N_10937);
or U12426 (N_12426,N_10954,N_10833);
nor U12427 (N_12427,N_11440,N_11294);
or U12428 (N_12428,N_10895,N_11174);
and U12429 (N_12429,N_11901,N_11722);
or U12430 (N_12430,N_11595,N_10821);
nor U12431 (N_12431,N_11904,N_11305);
nand U12432 (N_12432,N_10996,N_11336);
nor U12433 (N_12433,N_11933,N_11370);
and U12434 (N_12434,N_11105,N_10881);
or U12435 (N_12435,N_11157,N_11437);
and U12436 (N_12436,N_11603,N_11067);
xor U12437 (N_12437,N_11630,N_11819);
and U12438 (N_12438,N_10808,N_11604);
or U12439 (N_12439,N_11663,N_10911);
nand U12440 (N_12440,N_11375,N_11363);
xnor U12441 (N_12441,N_11944,N_11677);
and U12442 (N_12442,N_11558,N_11963);
and U12443 (N_12443,N_11088,N_11359);
or U12444 (N_12444,N_11225,N_10862);
and U12445 (N_12445,N_11949,N_11520);
nor U12446 (N_12446,N_11337,N_11894);
or U12447 (N_12447,N_11981,N_11552);
or U12448 (N_12448,N_11024,N_10855);
or U12449 (N_12449,N_11665,N_10890);
nand U12450 (N_12450,N_11838,N_11763);
nor U12451 (N_12451,N_11226,N_11622);
or U12452 (N_12452,N_11813,N_11208);
and U12453 (N_12453,N_10912,N_10929);
nor U12454 (N_12454,N_11497,N_11463);
nand U12455 (N_12455,N_11699,N_11614);
and U12456 (N_12456,N_11135,N_11115);
or U12457 (N_12457,N_11266,N_11790);
nand U12458 (N_12458,N_11600,N_11877);
and U12459 (N_12459,N_11056,N_11334);
nor U12460 (N_12460,N_11511,N_11415);
and U12461 (N_12461,N_11920,N_11288);
and U12462 (N_12462,N_11547,N_11074);
xnor U12463 (N_12463,N_11498,N_11993);
nand U12464 (N_12464,N_10999,N_11740);
nor U12465 (N_12465,N_11660,N_11563);
nand U12466 (N_12466,N_10858,N_11572);
xor U12467 (N_12467,N_10983,N_11980);
nor U12468 (N_12468,N_11146,N_11057);
nor U12469 (N_12469,N_11586,N_11227);
nand U12470 (N_12470,N_11908,N_11188);
nand U12471 (N_12471,N_11689,N_11239);
or U12472 (N_12472,N_11431,N_11048);
nand U12473 (N_12473,N_11999,N_10802);
nor U12474 (N_12474,N_11462,N_11831);
and U12475 (N_12475,N_11106,N_10838);
nand U12476 (N_12476,N_10909,N_11610);
and U12477 (N_12477,N_11243,N_11845);
or U12478 (N_12478,N_11086,N_11538);
nor U12479 (N_12479,N_11587,N_11688);
or U12480 (N_12480,N_11750,N_11061);
nor U12481 (N_12481,N_11396,N_11173);
or U12482 (N_12482,N_11727,N_11961);
nand U12483 (N_12483,N_11747,N_10879);
nor U12484 (N_12484,N_11598,N_11043);
nand U12485 (N_12485,N_11032,N_11229);
nand U12486 (N_12486,N_11967,N_11615);
xnor U12487 (N_12487,N_11705,N_11080);
nor U12488 (N_12488,N_10877,N_11263);
nand U12489 (N_12489,N_11052,N_11799);
and U12490 (N_12490,N_11308,N_11549);
xor U12491 (N_12491,N_11977,N_11182);
or U12492 (N_12492,N_11557,N_11738);
nand U12493 (N_12493,N_11527,N_11823);
xor U12494 (N_12494,N_11702,N_10852);
and U12495 (N_12495,N_11160,N_11814);
xor U12496 (N_12496,N_11060,N_11736);
nor U12497 (N_12497,N_11583,N_11759);
and U12498 (N_12498,N_11481,N_11764);
nor U12499 (N_12499,N_11005,N_11013);
nand U12500 (N_12500,N_11915,N_11792);
and U12501 (N_12501,N_10888,N_11009);
xor U12502 (N_12502,N_10970,N_10965);
nor U12503 (N_12503,N_10973,N_11012);
or U12504 (N_12504,N_10871,N_11849);
or U12505 (N_12505,N_11244,N_11959);
nor U12506 (N_12506,N_11871,N_10940);
nor U12507 (N_12507,N_11632,N_10958);
nand U12508 (N_12508,N_11351,N_11347);
nor U12509 (N_12509,N_11869,N_11103);
nand U12510 (N_12510,N_11311,N_11417);
and U12511 (N_12511,N_11709,N_11580);
nor U12512 (N_12512,N_10851,N_11377);
and U12513 (N_12513,N_11171,N_11192);
nor U12514 (N_12514,N_11619,N_11070);
and U12515 (N_12515,N_11116,N_11668);
nand U12516 (N_12516,N_11207,N_11874);
or U12517 (N_12517,N_11952,N_10809);
xnor U12518 (N_12518,N_11050,N_11293);
nor U12519 (N_12519,N_11306,N_11455);
and U12520 (N_12520,N_11794,N_10891);
nand U12521 (N_12521,N_11150,N_11271);
or U12522 (N_12522,N_11477,N_10993);
nor U12523 (N_12523,N_11193,N_11940);
and U12524 (N_12524,N_11385,N_11617);
nand U12525 (N_12525,N_11789,N_10814);
nand U12526 (N_12526,N_11795,N_11798);
xnor U12527 (N_12527,N_10868,N_11278);
and U12528 (N_12528,N_11518,N_10959);
xor U12529 (N_12529,N_11994,N_10990);
and U12530 (N_12530,N_11291,N_11485);
nor U12531 (N_12531,N_11541,N_11362);
and U12532 (N_12532,N_11573,N_11331);
and U12533 (N_12533,N_11469,N_11404);
xor U12534 (N_12534,N_10903,N_11589);
nand U12535 (N_12535,N_11596,N_11427);
nor U12536 (N_12536,N_11796,N_11791);
or U12537 (N_12537,N_10830,N_11907);
xor U12538 (N_12538,N_11863,N_11197);
nand U12539 (N_12539,N_11494,N_11925);
xor U12540 (N_12540,N_11273,N_11649);
nand U12541 (N_12541,N_11213,N_11998);
nor U12542 (N_12542,N_11623,N_10867);
xnor U12543 (N_12543,N_11029,N_11015);
nand U12544 (N_12544,N_11806,N_11828);
nand U12545 (N_12545,N_11096,N_10963);
or U12546 (N_12546,N_11242,N_11488);
and U12547 (N_12547,N_11693,N_11848);
or U12548 (N_12548,N_11063,N_11982);
or U12549 (N_12549,N_10863,N_11776);
nor U12550 (N_12550,N_11360,N_11723);
nor U12551 (N_12551,N_11588,N_11003);
and U12552 (N_12552,N_11866,N_11733);
nand U12553 (N_12553,N_11442,N_11194);
or U12554 (N_12554,N_10941,N_11612);
and U12555 (N_12555,N_11818,N_11097);
nand U12556 (N_12556,N_11880,N_11324);
or U12557 (N_12557,N_10910,N_11954);
or U12558 (N_12558,N_11850,N_11089);
xnor U12559 (N_12559,N_10945,N_11569);
nand U12560 (N_12560,N_10854,N_11992);
xnor U12561 (N_12561,N_11259,N_11882);
nor U12562 (N_12562,N_11390,N_10812);
or U12563 (N_12563,N_11645,N_11302);
nand U12564 (N_12564,N_11758,N_11910);
xnor U12565 (N_12565,N_11718,N_11447);
nor U12566 (N_12566,N_11087,N_11505);
and U12567 (N_12567,N_11249,N_10925);
and U12568 (N_12568,N_11429,N_11559);
and U12569 (N_12569,N_11931,N_10889);
nand U12570 (N_12570,N_11149,N_10828);
or U12571 (N_12571,N_11328,N_10956);
xnor U12572 (N_12572,N_11620,N_11142);
and U12573 (N_12573,N_10898,N_11545);
and U12574 (N_12574,N_11737,N_11268);
or U12575 (N_12575,N_11537,N_11653);
xor U12576 (N_12576,N_11027,N_10824);
xnor U12577 (N_12577,N_11049,N_11240);
nor U12578 (N_12578,N_11358,N_11592);
and U12579 (N_12579,N_11997,N_11683);
xor U12580 (N_12580,N_11713,N_11777);
nand U12581 (N_12581,N_11456,N_11101);
nor U12582 (N_12582,N_11704,N_11412);
xor U12583 (N_12583,N_11698,N_11501);
nor U12584 (N_12584,N_11315,N_11648);
xnor U12585 (N_12585,N_10904,N_11212);
nand U12586 (N_12586,N_10933,N_10920);
and U12587 (N_12587,N_11503,N_11071);
nand U12588 (N_12588,N_11314,N_11766);
or U12589 (N_12589,N_11987,N_11633);
xor U12590 (N_12590,N_11355,N_11499);
xor U12591 (N_12591,N_11856,N_10857);
or U12592 (N_12592,N_11637,N_11020);
or U12593 (N_12593,N_10949,N_11284);
or U12594 (N_12594,N_10829,N_11255);
xnor U12595 (N_12595,N_11232,N_11757);
nor U12596 (N_12596,N_11840,N_11768);
nand U12597 (N_12597,N_10919,N_10864);
nand U12598 (N_12598,N_11117,N_11578);
nand U12599 (N_12599,N_11692,N_11696);
and U12600 (N_12600,N_11741,N_10983);
xor U12601 (N_12601,N_10820,N_11862);
nor U12602 (N_12602,N_11362,N_11755);
nor U12603 (N_12603,N_11328,N_11302);
nand U12604 (N_12604,N_11250,N_11882);
nand U12605 (N_12605,N_11953,N_10904);
nor U12606 (N_12606,N_11471,N_11476);
nand U12607 (N_12607,N_11422,N_11050);
xnor U12608 (N_12608,N_11899,N_10884);
and U12609 (N_12609,N_11275,N_11212);
xnor U12610 (N_12610,N_11557,N_11116);
and U12611 (N_12611,N_11731,N_11156);
xnor U12612 (N_12612,N_11449,N_11011);
and U12613 (N_12613,N_11353,N_11472);
or U12614 (N_12614,N_10942,N_11410);
nand U12615 (N_12615,N_11398,N_11240);
and U12616 (N_12616,N_11386,N_11125);
xnor U12617 (N_12617,N_11366,N_11644);
xor U12618 (N_12618,N_11001,N_11695);
xor U12619 (N_12619,N_11153,N_11025);
and U12620 (N_12620,N_11062,N_10813);
xnor U12621 (N_12621,N_11280,N_11473);
nor U12622 (N_12622,N_11093,N_10884);
nor U12623 (N_12623,N_11588,N_11454);
and U12624 (N_12624,N_11143,N_10934);
xor U12625 (N_12625,N_11732,N_11033);
or U12626 (N_12626,N_11337,N_11803);
xnor U12627 (N_12627,N_11468,N_11135);
nor U12628 (N_12628,N_11616,N_11230);
and U12629 (N_12629,N_11311,N_11025);
nor U12630 (N_12630,N_11468,N_11824);
nand U12631 (N_12631,N_11512,N_10921);
and U12632 (N_12632,N_10924,N_10966);
and U12633 (N_12633,N_11228,N_11618);
or U12634 (N_12634,N_11921,N_11364);
or U12635 (N_12635,N_11808,N_10926);
or U12636 (N_12636,N_10850,N_11679);
or U12637 (N_12637,N_11663,N_11946);
nand U12638 (N_12638,N_11648,N_10871);
nor U12639 (N_12639,N_11688,N_11631);
nand U12640 (N_12640,N_11250,N_11547);
or U12641 (N_12641,N_11635,N_10907);
xnor U12642 (N_12642,N_11544,N_11884);
xor U12643 (N_12643,N_11081,N_11860);
and U12644 (N_12644,N_11838,N_11132);
nor U12645 (N_12645,N_11380,N_11289);
xor U12646 (N_12646,N_11943,N_11340);
xnor U12647 (N_12647,N_11103,N_11562);
xnor U12648 (N_12648,N_10978,N_11459);
nor U12649 (N_12649,N_11371,N_11073);
xnor U12650 (N_12650,N_11439,N_11387);
and U12651 (N_12651,N_11332,N_10801);
xnor U12652 (N_12652,N_11937,N_11705);
or U12653 (N_12653,N_11081,N_11839);
nor U12654 (N_12654,N_11326,N_11641);
and U12655 (N_12655,N_11945,N_11377);
or U12656 (N_12656,N_11075,N_11329);
or U12657 (N_12657,N_11658,N_11227);
and U12658 (N_12658,N_11958,N_11702);
nand U12659 (N_12659,N_11303,N_11331);
and U12660 (N_12660,N_11167,N_11580);
or U12661 (N_12661,N_11879,N_11445);
or U12662 (N_12662,N_11863,N_11010);
or U12663 (N_12663,N_11065,N_11576);
and U12664 (N_12664,N_11487,N_11106);
xnor U12665 (N_12665,N_11980,N_11784);
xor U12666 (N_12666,N_11995,N_11287);
nand U12667 (N_12667,N_11340,N_11761);
nor U12668 (N_12668,N_11561,N_10963);
nand U12669 (N_12669,N_11998,N_11532);
and U12670 (N_12670,N_11467,N_11946);
and U12671 (N_12671,N_11560,N_11409);
xnor U12672 (N_12672,N_10890,N_11441);
nand U12673 (N_12673,N_11138,N_10864);
xnor U12674 (N_12674,N_11965,N_11527);
nand U12675 (N_12675,N_11751,N_11763);
nor U12676 (N_12676,N_11300,N_11001);
nand U12677 (N_12677,N_11838,N_11094);
xnor U12678 (N_12678,N_10803,N_11286);
or U12679 (N_12679,N_11511,N_11451);
xnor U12680 (N_12680,N_11157,N_11205);
or U12681 (N_12681,N_11583,N_11715);
nand U12682 (N_12682,N_11571,N_11389);
nor U12683 (N_12683,N_11923,N_11535);
xor U12684 (N_12684,N_11019,N_11038);
and U12685 (N_12685,N_11758,N_10889);
or U12686 (N_12686,N_11664,N_11427);
and U12687 (N_12687,N_11495,N_11461);
or U12688 (N_12688,N_11138,N_11818);
nand U12689 (N_12689,N_11721,N_11358);
nor U12690 (N_12690,N_11687,N_11278);
nand U12691 (N_12691,N_10979,N_11854);
nand U12692 (N_12692,N_11543,N_11447);
or U12693 (N_12693,N_11387,N_11107);
nor U12694 (N_12694,N_11182,N_11948);
and U12695 (N_12695,N_11424,N_11300);
xnor U12696 (N_12696,N_11915,N_11228);
nor U12697 (N_12697,N_10830,N_11151);
and U12698 (N_12698,N_11470,N_11301);
xor U12699 (N_12699,N_11075,N_11545);
nand U12700 (N_12700,N_10822,N_11407);
nor U12701 (N_12701,N_11827,N_11740);
and U12702 (N_12702,N_11108,N_11453);
and U12703 (N_12703,N_11380,N_11695);
nand U12704 (N_12704,N_11958,N_11667);
nor U12705 (N_12705,N_11494,N_11734);
and U12706 (N_12706,N_11826,N_11714);
and U12707 (N_12707,N_11774,N_11068);
or U12708 (N_12708,N_11808,N_11286);
xor U12709 (N_12709,N_11248,N_10962);
nand U12710 (N_12710,N_11051,N_11555);
xor U12711 (N_12711,N_11096,N_11213);
nand U12712 (N_12712,N_10830,N_11165);
nor U12713 (N_12713,N_11862,N_11610);
or U12714 (N_12714,N_11953,N_11375);
nand U12715 (N_12715,N_11253,N_11193);
and U12716 (N_12716,N_10882,N_11596);
and U12717 (N_12717,N_11955,N_10962);
or U12718 (N_12718,N_11517,N_10886);
and U12719 (N_12719,N_11754,N_11988);
or U12720 (N_12720,N_11534,N_11889);
nand U12721 (N_12721,N_11676,N_11010);
nand U12722 (N_12722,N_11099,N_11390);
nand U12723 (N_12723,N_11298,N_11677);
and U12724 (N_12724,N_11879,N_11272);
or U12725 (N_12725,N_11659,N_11446);
nor U12726 (N_12726,N_11460,N_11905);
and U12727 (N_12727,N_11684,N_11030);
or U12728 (N_12728,N_11085,N_10920);
and U12729 (N_12729,N_11771,N_11681);
or U12730 (N_12730,N_11736,N_11616);
or U12731 (N_12731,N_11649,N_11221);
xor U12732 (N_12732,N_11315,N_11077);
xor U12733 (N_12733,N_11269,N_11154);
nor U12734 (N_12734,N_11297,N_11270);
nor U12735 (N_12735,N_11368,N_11370);
and U12736 (N_12736,N_11201,N_11944);
xnor U12737 (N_12737,N_11589,N_11844);
xnor U12738 (N_12738,N_11197,N_11824);
nor U12739 (N_12739,N_11886,N_11644);
or U12740 (N_12740,N_11549,N_11647);
nand U12741 (N_12741,N_11604,N_10911);
and U12742 (N_12742,N_11255,N_11636);
and U12743 (N_12743,N_11457,N_11456);
or U12744 (N_12744,N_11853,N_11481);
nand U12745 (N_12745,N_11909,N_11076);
or U12746 (N_12746,N_11958,N_11545);
or U12747 (N_12747,N_11729,N_11825);
xnor U12748 (N_12748,N_10821,N_11562);
or U12749 (N_12749,N_10920,N_11887);
xor U12750 (N_12750,N_11876,N_11015);
nor U12751 (N_12751,N_11373,N_10980);
xnor U12752 (N_12752,N_10865,N_10957);
xnor U12753 (N_12753,N_10911,N_11739);
nor U12754 (N_12754,N_11212,N_11961);
nand U12755 (N_12755,N_11618,N_11844);
and U12756 (N_12756,N_11750,N_10862);
and U12757 (N_12757,N_11020,N_11372);
nor U12758 (N_12758,N_11326,N_11523);
nor U12759 (N_12759,N_11533,N_10892);
nand U12760 (N_12760,N_11395,N_11335);
nand U12761 (N_12761,N_11130,N_10809);
or U12762 (N_12762,N_11669,N_11943);
nand U12763 (N_12763,N_11982,N_11308);
xor U12764 (N_12764,N_11131,N_11443);
or U12765 (N_12765,N_11106,N_11747);
xnor U12766 (N_12766,N_11949,N_11049);
nand U12767 (N_12767,N_11056,N_11675);
or U12768 (N_12768,N_11306,N_11640);
xor U12769 (N_12769,N_11130,N_11506);
and U12770 (N_12770,N_11335,N_11547);
xor U12771 (N_12771,N_11316,N_11257);
xor U12772 (N_12772,N_11743,N_11772);
and U12773 (N_12773,N_11829,N_11630);
nand U12774 (N_12774,N_11457,N_11595);
nor U12775 (N_12775,N_11291,N_10918);
xnor U12776 (N_12776,N_11535,N_11747);
nor U12777 (N_12777,N_11897,N_11090);
nand U12778 (N_12778,N_11960,N_11930);
or U12779 (N_12779,N_11358,N_11500);
and U12780 (N_12780,N_11135,N_11881);
or U12781 (N_12781,N_11289,N_11738);
nand U12782 (N_12782,N_10853,N_10827);
xnor U12783 (N_12783,N_11007,N_10907);
or U12784 (N_12784,N_11941,N_11735);
nand U12785 (N_12785,N_11268,N_11931);
and U12786 (N_12786,N_11510,N_11433);
or U12787 (N_12787,N_11335,N_11076);
xnor U12788 (N_12788,N_11365,N_11888);
or U12789 (N_12789,N_11569,N_11089);
or U12790 (N_12790,N_11192,N_11949);
nor U12791 (N_12791,N_10814,N_11139);
and U12792 (N_12792,N_11939,N_11421);
nor U12793 (N_12793,N_11913,N_11231);
and U12794 (N_12794,N_11952,N_11237);
nor U12795 (N_12795,N_11031,N_11114);
and U12796 (N_12796,N_11707,N_11028);
and U12797 (N_12797,N_10872,N_11327);
or U12798 (N_12798,N_11308,N_10929);
nand U12799 (N_12799,N_11274,N_11966);
or U12800 (N_12800,N_11037,N_10966);
nor U12801 (N_12801,N_11649,N_11872);
nor U12802 (N_12802,N_11422,N_11673);
nor U12803 (N_12803,N_11253,N_10926);
xor U12804 (N_12804,N_11114,N_10856);
nor U12805 (N_12805,N_11650,N_11344);
nand U12806 (N_12806,N_11690,N_11748);
and U12807 (N_12807,N_11731,N_10808);
nand U12808 (N_12808,N_11768,N_11223);
and U12809 (N_12809,N_11438,N_11749);
and U12810 (N_12810,N_11353,N_11951);
xor U12811 (N_12811,N_11182,N_11215);
nor U12812 (N_12812,N_11862,N_11542);
and U12813 (N_12813,N_11760,N_11396);
nand U12814 (N_12814,N_11972,N_11507);
nor U12815 (N_12815,N_10890,N_11816);
xor U12816 (N_12816,N_11286,N_10939);
xor U12817 (N_12817,N_11022,N_11965);
nand U12818 (N_12818,N_11067,N_11833);
nand U12819 (N_12819,N_10902,N_11890);
or U12820 (N_12820,N_11600,N_11188);
xnor U12821 (N_12821,N_11493,N_11017);
xor U12822 (N_12822,N_11894,N_11373);
xnor U12823 (N_12823,N_11423,N_11510);
and U12824 (N_12824,N_11927,N_11682);
or U12825 (N_12825,N_11605,N_10996);
and U12826 (N_12826,N_10882,N_11056);
nor U12827 (N_12827,N_11623,N_10941);
nand U12828 (N_12828,N_11109,N_11631);
and U12829 (N_12829,N_11808,N_11748);
nand U12830 (N_12830,N_11604,N_11413);
and U12831 (N_12831,N_11310,N_10842);
or U12832 (N_12832,N_11471,N_10805);
nand U12833 (N_12833,N_11148,N_11179);
and U12834 (N_12834,N_11076,N_11468);
nand U12835 (N_12835,N_11412,N_11915);
and U12836 (N_12836,N_11707,N_11926);
and U12837 (N_12837,N_11424,N_11430);
and U12838 (N_12838,N_10881,N_11655);
and U12839 (N_12839,N_11006,N_11677);
nor U12840 (N_12840,N_11240,N_11715);
xor U12841 (N_12841,N_11285,N_11632);
or U12842 (N_12842,N_11380,N_11216);
or U12843 (N_12843,N_11453,N_11222);
or U12844 (N_12844,N_11820,N_10925);
and U12845 (N_12845,N_11370,N_10959);
nand U12846 (N_12846,N_10987,N_11176);
nor U12847 (N_12847,N_10909,N_11811);
or U12848 (N_12848,N_11525,N_11551);
nor U12849 (N_12849,N_10897,N_11764);
nor U12850 (N_12850,N_11901,N_11512);
and U12851 (N_12851,N_11761,N_11453);
nand U12852 (N_12852,N_10930,N_11391);
or U12853 (N_12853,N_11067,N_10866);
and U12854 (N_12854,N_11638,N_11774);
nor U12855 (N_12855,N_11819,N_11536);
nand U12856 (N_12856,N_11773,N_11166);
or U12857 (N_12857,N_10894,N_11726);
and U12858 (N_12858,N_11935,N_11408);
nand U12859 (N_12859,N_11415,N_11738);
and U12860 (N_12860,N_11335,N_11597);
nand U12861 (N_12861,N_11215,N_11367);
and U12862 (N_12862,N_10887,N_10826);
xnor U12863 (N_12863,N_11772,N_11139);
xnor U12864 (N_12864,N_11783,N_11483);
nor U12865 (N_12865,N_11223,N_11236);
nand U12866 (N_12866,N_11734,N_11341);
nand U12867 (N_12867,N_11562,N_11024);
nor U12868 (N_12868,N_10911,N_11060);
xnor U12869 (N_12869,N_10940,N_11342);
nor U12870 (N_12870,N_10882,N_11747);
nor U12871 (N_12871,N_11612,N_11803);
and U12872 (N_12872,N_11404,N_11494);
or U12873 (N_12873,N_11237,N_11464);
or U12874 (N_12874,N_11944,N_11207);
xor U12875 (N_12875,N_11356,N_10871);
and U12876 (N_12876,N_10882,N_11605);
nor U12877 (N_12877,N_10926,N_11432);
or U12878 (N_12878,N_11253,N_10829);
nand U12879 (N_12879,N_11462,N_11336);
and U12880 (N_12880,N_11809,N_11377);
nand U12881 (N_12881,N_11272,N_11475);
or U12882 (N_12882,N_11297,N_11198);
nand U12883 (N_12883,N_11341,N_11342);
nor U12884 (N_12884,N_11352,N_10986);
or U12885 (N_12885,N_11460,N_11017);
xnor U12886 (N_12886,N_11686,N_10944);
and U12887 (N_12887,N_11368,N_11910);
or U12888 (N_12888,N_11943,N_10838);
nand U12889 (N_12889,N_11735,N_11510);
nand U12890 (N_12890,N_11224,N_10803);
nor U12891 (N_12891,N_11911,N_11969);
xor U12892 (N_12892,N_11712,N_10949);
nor U12893 (N_12893,N_10914,N_11350);
xor U12894 (N_12894,N_11075,N_10886);
or U12895 (N_12895,N_10985,N_11424);
or U12896 (N_12896,N_11882,N_11792);
nor U12897 (N_12897,N_11323,N_10948);
xor U12898 (N_12898,N_10820,N_11735);
or U12899 (N_12899,N_10840,N_11873);
xnor U12900 (N_12900,N_11757,N_11988);
nor U12901 (N_12901,N_11369,N_11379);
xor U12902 (N_12902,N_11335,N_10844);
or U12903 (N_12903,N_11891,N_11001);
nand U12904 (N_12904,N_11312,N_11292);
or U12905 (N_12905,N_11395,N_11192);
nor U12906 (N_12906,N_10982,N_11088);
xor U12907 (N_12907,N_11584,N_11904);
or U12908 (N_12908,N_11647,N_11037);
nor U12909 (N_12909,N_11943,N_11649);
and U12910 (N_12910,N_11373,N_11289);
and U12911 (N_12911,N_11097,N_11540);
nand U12912 (N_12912,N_11477,N_11352);
nor U12913 (N_12913,N_10803,N_10907);
or U12914 (N_12914,N_11750,N_11074);
xor U12915 (N_12915,N_10857,N_11627);
and U12916 (N_12916,N_11566,N_11675);
nor U12917 (N_12917,N_11526,N_11940);
nand U12918 (N_12918,N_11967,N_11785);
and U12919 (N_12919,N_11906,N_11517);
nand U12920 (N_12920,N_10964,N_11446);
nor U12921 (N_12921,N_11315,N_11899);
xor U12922 (N_12922,N_11952,N_11410);
xnor U12923 (N_12923,N_11673,N_11059);
xnor U12924 (N_12924,N_11297,N_11336);
and U12925 (N_12925,N_10947,N_11200);
nand U12926 (N_12926,N_11836,N_11359);
or U12927 (N_12927,N_11177,N_11047);
xnor U12928 (N_12928,N_11275,N_11440);
xnor U12929 (N_12929,N_11951,N_11835);
xor U12930 (N_12930,N_11257,N_11037);
nand U12931 (N_12931,N_11664,N_10925);
xnor U12932 (N_12932,N_11474,N_11247);
and U12933 (N_12933,N_11960,N_10972);
xor U12934 (N_12934,N_10813,N_10997);
nor U12935 (N_12935,N_11426,N_11273);
or U12936 (N_12936,N_11400,N_10911);
nor U12937 (N_12937,N_11718,N_11397);
nand U12938 (N_12938,N_11291,N_11557);
and U12939 (N_12939,N_11082,N_11540);
or U12940 (N_12940,N_11759,N_11368);
nand U12941 (N_12941,N_11636,N_11416);
and U12942 (N_12942,N_11092,N_11757);
nor U12943 (N_12943,N_10852,N_11153);
nor U12944 (N_12944,N_11461,N_11348);
nor U12945 (N_12945,N_11706,N_10881);
nor U12946 (N_12946,N_11451,N_10843);
nand U12947 (N_12947,N_11258,N_10816);
xnor U12948 (N_12948,N_11126,N_11796);
or U12949 (N_12949,N_11592,N_11509);
nor U12950 (N_12950,N_10847,N_11748);
nor U12951 (N_12951,N_11399,N_11515);
or U12952 (N_12952,N_11437,N_10911);
nor U12953 (N_12953,N_11069,N_11881);
and U12954 (N_12954,N_11640,N_11744);
or U12955 (N_12955,N_10896,N_11457);
or U12956 (N_12956,N_11218,N_11408);
nor U12957 (N_12957,N_11566,N_11122);
xor U12958 (N_12958,N_11745,N_11561);
xor U12959 (N_12959,N_11822,N_11604);
nor U12960 (N_12960,N_11033,N_11232);
xor U12961 (N_12961,N_11626,N_10993);
and U12962 (N_12962,N_11695,N_11203);
nand U12963 (N_12963,N_11255,N_11813);
and U12964 (N_12964,N_11882,N_11863);
xnor U12965 (N_12965,N_11106,N_11462);
nor U12966 (N_12966,N_11335,N_11856);
nand U12967 (N_12967,N_11899,N_11319);
xnor U12968 (N_12968,N_11146,N_11703);
xnor U12969 (N_12969,N_11945,N_11361);
xnor U12970 (N_12970,N_11117,N_11554);
and U12971 (N_12971,N_11822,N_11323);
or U12972 (N_12972,N_11873,N_11467);
xnor U12973 (N_12973,N_11382,N_11964);
nor U12974 (N_12974,N_10935,N_11654);
nand U12975 (N_12975,N_11703,N_11562);
or U12976 (N_12976,N_11266,N_10923);
or U12977 (N_12977,N_11984,N_11249);
nand U12978 (N_12978,N_11776,N_11951);
nand U12979 (N_12979,N_11120,N_10962);
xor U12980 (N_12980,N_11809,N_11375);
xor U12981 (N_12981,N_11342,N_11695);
nand U12982 (N_12982,N_10953,N_10824);
and U12983 (N_12983,N_10922,N_11197);
nand U12984 (N_12984,N_10966,N_11003);
and U12985 (N_12985,N_11606,N_11062);
xnor U12986 (N_12986,N_11325,N_11201);
and U12987 (N_12987,N_11524,N_11624);
nand U12988 (N_12988,N_11828,N_11774);
nand U12989 (N_12989,N_11209,N_11673);
xnor U12990 (N_12990,N_11067,N_11088);
or U12991 (N_12991,N_11346,N_11126);
and U12992 (N_12992,N_11002,N_11026);
and U12993 (N_12993,N_10957,N_11064);
or U12994 (N_12994,N_11737,N_11777);
and U12995 (N_12995,N_10803,N_11998);
nand U12996 (N_12996,N_11049,N_11468);
and U12997 (N_12997,N_11041,N_11071);
xor U12998 (N_12998,N_11339,N_11588);
or U12999 (N_12999,N_11568,N_11593);
or U13000 (N_13000,N_11944,N_11560);
xor U13001 (N_13001,N_10921,N_11854);
and U13002 (N_13002,N_11583,N_11608);
nand U13003 (N_13003,N_11710,N_11762);
xnor U13004 (N_13004,N_11520,N_11856);
and U13005 (N_13005,N_11188,N_11259);
nand U13006 (N_13006,N_11798,N_11653);
nand U13007 (N_13007,N_11713,N_11812);
nand U13008 (N_13008,N_11378,N_11000);
nand U13009 (N_13009,N_11446,N_11647);
nand U13010 (N_13010,N_11315,N_11096);
nor U13011 (N_13011,N_11260,N_11997);
nand U13012 (N_13012,N_11616,N_11896);
or U13013 (N_13013,N_11976,N_11687);
xnor U13014 (N_13014,N_11461,N_10858);
nand U13015 (N_13015,N_11992,N_11469);
nor U13016 (N_13016,N_11747,N_10851);
xor U13017 (N_13017,N_11701,N_10801);
and U13018 (N_13018,N_10906,N_11117);
nand U13019 (N_13019,N_11747,N_11579);
nand U13020 (N_13020,N_11819,N_11439);
and U13021 (N_13021,N_11737,N_11346);
xnor U13022 (N_13022,N_11130,N_11003);
xnor U13023 (N_13023,N_11942,N_10841);
nand U13024 (N_13024,N_11249,N_10854);
or U13025 (N_13025,N_11051,N_10893);
nor U13026 (N_13026,N_11597,N_11257);
xnor U13027 (N_13027,N_11507,N_11054);
xor U13028 (N_13028,N_11437,N_10816);
and U13029 (N_13029,N_11153,N_11554);
or U13030 (N_13030,N_11750,N_10940);
and U13031 (N_13031,N_11180,N_11613);
xnor U13032 (N_13032,N_11585,N_11808);
and U13033 (N_13033,N_11831,N_11005);
and U13034 (N_13034,N_11042,N_11498);
and U13035 (N_13035,N_11334,N_10909);
xor U13036 (N_13036,N_11989,N_11884);
and U13037 (N_13037,N_10989,N_10819);
xor U13038 (N_13038,N_11369,N_10950);
and U13039 (N_13039,N_11246,N_11257);
nand U13040 (N_13040,N_11949,N_11529);
or U13041 (N_13041,N_11967,N_11529);
xor U13042 (N_13042,N_11808,N_11750);
nor U13043 (N_13043,N_11824,N_10827);
nor U13044 (N_13044,N_11057,N_11125);
or U13045 (N_13045,N_11443,N_11129);
nand U13046 (N_13046,N_11086,N_11066);
and U13047 (N_13047,N_11510,N_11141);
and U13048 (N_13048,N_11402,N_11681);
or U13049 (N_13049,N_11558,N_11922);
nor U13050 (N_13050,N_11210,N_11206);
or U13051 (N_13051,N_11737,N_11551);
nand U13052 (N_13052,N_11857,N_11767);
nor U13053 (N_13053,N_11218,N_10952);
and U13054 (N_13054,N_11773,N_11002);
or U13055 (N_13055,N_11624,N_11824);
nand U13056 (N_13056,N_11788,N_11136);
and U13057 (N_13057,N_11588,N_10932);
and U13058 (N_13058,N_11977,N_11455);
nand U13059 (N_13059,N_11939,N_11034);
xor U13060 (N_13060,N_11845,N_10931);
nor U13061 (N_13061,N_11112,N_11048);
xnor U13062 (N_13062,N_11436,N_11992);
nand U13063 (N_13063,N_11459,N_10886);
xnor U13064 (N_13064,N_11074,N_10893);
or U13065 (N_13065,N_11757,N_10975);
xnor U13066 (N_13066,N_11432,N_11904);
xnor U13067 (N_13067,N_11801,N_11809);
xnor U13068 (N_13068,N_11865,N_11213);
or U13069 (N_13069,N_10952,N_11829);
and U13070 (N_13070,N_11607,N_11527);
and U13071 (N_13071,N_11129,N_11351);
nand U13072 (N_13072,N_11756,N_11879);
xnor U13073 (N_13073,N_11072,N_11875);
xor U13074 (N_13074,N_11596,N_11586);
xnor U13075 (N_13075,N_11936,N_11090);
xor U13076 (N_13076,N_11579,N_10819);
nand U13077 (N_13077,N_11225,N_11865);
and U13078 (N_13078,N_10818,N_10948);
and U13079 (N_13079,N_11486,N_11003);
nor U13080 (N_13080,N_11114,N_11494);
and U13081 (N_13081,N_11641,N_11714);
xor U13082 (N_13082,N_11441,N_11468);
xnor U13083 (N_13083,N_10924,N_11744);
nand U13084 (N_13084,N_11582,N_11399);
and U13085 (N_13085,N_11152,N_11287);
nand U13086 (N_13086,N_11444,N_10996);
xor U13087 (N_13087,N_11248,N_11225);
xor U13088 (N_13088,N_11563,N_11889);
nor U13089 (N_13089,N_11783,N_11561);
xor U13090 (N_13090,N_11377,N_11051);
nor U13091 (N_13091,N_11468,N_10876);
xnor U13092 (N_13092,N_11126,N_11009);
nor U13093 (N_13093,N_11678,N_11234);
nor U13094 (N_13094,N_11513,N_11352);
or U13095 (N_13095,N_11006,N_11097);
nand U13096 (N_13096,N_11921,N_11714);
nor U13097 (N_13097,N_10985,N_11008);
nand U13098 (N_13098,N_11059,N_11101);
or U13099 (N_13099,N_11509,N_11585);
nand U13100 (N_13100,N_11821,N_11930);
nor U13101 (N_13101,N_11393,N_11214);
nand U13102 (N_13102,N_11994,N_11075);
or U13103 (N_13103,N_10823,N_10911);
and U13104 (N_13104,N_11240,N_11773);
xnor U13105 (N_13105,N_11616,N_11590);
and U13106 (N_13106,N_11160,N_11403);
or U13107 (N_13107,N_11904,N_11657);
and U13108 (N_13108,N_10939,N_11820);
nand U13109 (N_13109,N_11350,N_11663);
and U13110 (N_13110,N_10963,N_11081);
or U13111 (N_13111,N_11035,N_11091);
nand U13112 (N_13112,N_11101,N_11245);
nand U13113 (N_13113,N_11494,N_10854);
and U13114 (N_13114,N_11599,N_11320);
or U13115 (N_13115,N_11258,N_11430);
and U13116 (N_13116,N_11609,N_11732);
nand U13117 (N_13117,N_10957,N_11259);
or U13118 (N_13118,N_11517,N_10920);
nand U13119 (N_13119,N_11974,N_11721);
and U13120 (N_13120,N_11666,N_11392);
nand U13121 (N_13121,N_11691,N_10954);
nor U13122 (N_13122,N_11206,N_11380);
or U13123 (N_13123,N_11946,N_11033);
and U13124 (N_13124,N_11356,N_11817);
and U13125 (N_13125,N_10960,N_11694);
xnor U13126 (N_13126,N_10938,N_11326);
nand U13127 (N_13127,N_10983,N_11977);
and U13128 (N_13128,N_11462,N_11801);
and U13129 (N_13129,N_10883,N_11433);
and U13130 (N_13130,N_11524,N_11793);
xor U13131 (N_13131,N_11527,N_11092);
nor U13132 (N_13132,N_11140,N_11690);
xor U13133 (N_13133,N_11739,N_11614);
or U13134 (N_13134,N_10809,N_11909);
nor U13135 (N_13135,N_10895,N_11438);
or U13136 (N_13136,N_10907,N_11724);
nor U13137 (N_13137,N_11145,N_11019);
or U13138 (N_13138,N_11425,N_11151);
nand U13139 (N_13139,N_11318,N_11165);
or U13140 (N_13140,N_11986,N_10993);
nand U13141 (N_13141,N_11011,N_11175);
and U13142 (N_13142,N_11602,N_11368);
xnor U13143 (N_13143,N_11701,N_11480);
nor U13144 (N_13144,N_11149,N_11060);
nand U13145 (N_13145,N_11128,N_10811);
nand U13146 (N_13146,N_11081,N_11079);
or U13147 (N_13147,N_10924,N_11194);
and U13148 (N_13148,N_11572,N_10905);
nor U13149 (N_13149,N_11956,N_11555);
nor U13150 (N_13150,N_11057,N_11780);
or U13151 (N_13151,N_11754,N_11130);
and U13152 (N_13152,N_11650,N_10886);
or U13153 (N_13153,N_10999,N_11002);
or U13154 (N_13154,N_11586,N_11501);
or U13155 (N_13155,N_11520,N_10932);
xor U13156 (N_13156,N_11510,N_11760);
nor U13157 (N_13157,N_10911,N_11651);
nand U13158 (N_13158,N_11770,N_11895);
nand U13159 (N_13159,N_11518,N_11293);
xor U13160 (N_13160,N_11759,N_11896);
and U13161 (N_13161,N_11704,N_10969);
or U13162 (N_13162,N_11468,N_11306);
nor U13163 (N_13163,N_11125,N_11243);
or U13164 (N_13164,N_11147,N_10973);
or U13165 (N_13165,N_11240,N_10816);
nand U13166 (N_13166,N_11071,N_11922);
and U13167 (N_13167,N_11483,N_11107);
xnor U13168 (N_13168,N_11447,N_10981);
xor U13169 (N_13169,N_11145,N_11843);
or U13170 (N_13170,N_11846,N_11614);
xnor U13171 (N_13171,N_11177,N_11951);
xor U13172 (N_13172,N_11002,N_11781);
xnor U13173 (N_13173,N_11321,N_11557);
nor U13174 (N_13174,N_11493,N_11503);
nor U13175 (N_13175,N_10873,N_10847);
or U13176 (N_13176,N_11471,N_11649);
xor U13177 (N_13177,N_10986,N_10989);
and U13178 (N_13178,N_11414,N_10974);
and U13179 (N_13179,N_11051,N_11198);
xor U13180 (N_13180,N_11915,N_11196);
or U13181 (N_13181,N_11949,N_10943);
and U13182 (N_13182,N_11218,N_10854);
nor U13183 (N_13183,N_11095,N_10827);
nor U13184 (N_13184,N_10819,N_11299);
and U13185 (N_13185,N_11712,N_11843);
and U13186 (N_13186,N_11311,N_10829);
and U13187 (N_13187,N_11716,N_11847);
and U13188 (N_13188,N_11178,N_11068);
xnor U13189 (N_13189,N_11131,N_11351);
or U13190 (N_13190,N_11520,N_11765);
nand U13191 (N_13191,N_11892,N_10937);
nand U13192 (N_13192,N_11277,N_10936);
or U13193 (N_13193,N_11989,N_10873);
and U13194 (N_13194,N_11255,N_11696);
nand U13195 (N_13195,N_11063,N_11375);
xnor U13196 (N_13196,N_11825,N_11479);
nand U13197 (N_13197,N_11318,N_11561);
xnor U13198 (N_13198,N_11848,N_11025);
and U13199 (N_13199,N_11936,N_11708);
xnor U13200 (N_13200,N_13182,N_12338);
nand U13201 (N_13201,N_12989,N_12045);
and U13202 (N_13202,N_12099,N_12445);
xnor U13203 (N_13203,N_12805,N_13149);
xor U13204 (N_13204,N_12532,N_12649);
or U13205 (N_13205,N_12376,N_12325);
nand U13206 (N_13206,N_13188,N_12450);
xnor U13207 (N_13207,N_12051,N_12578);
nand U13208 (N_13208,N_13047,N_12977);
nor U13209 (N_13209,N_12144,N_12334);
nand U13210 (N_13210,N_12278,N_12226);
nor U13211 (N_13211,N_12545,N_12692);
and U13212 (N_13212,N_12435,N_13062);
or U13213 (N_13213,N_12710,N_13152);
nand U13214 (N_13214,N_12676,N_12975);
nand U13215 (N_13215,N_12414,N_13007);
nor U13216 (N_13216,N_12103,N_12017);
nand U13217 (N_13217,N_12912,N_12901);
or U13218 (N_13218,N_13115,N_12406);
xnor U13219 (N_13219,N_13135,N_12394);
and U13220 (N_13220,N_12238,N_12335);
or U13221 (N_13221,N_12909,N_12988);
nor U13222 (N_13222,N_13093,N_12429);
xnor U13223 (N_13223,N_12328,N_13076);
and U13224 (N_13224,N_12900,N_12834);
xnor U13225 (N_13225,N_12675,N_12930);
or U13226 (N_13226,N_12377,N_12397);
nor U13227 (N_13227,N_13069,N_12211);
nand U13228 (N_13228,N_12196,N_12519);
and U13229 (N_13229,N_12311,N_12498);
nor U13230 (N_13230,N_12958,N_12155);
xnor U13231 (N_13231,N_12422,N_12235);
nand U13232 (N_13232,N_12405,N_12974);
nor U13233 (N_13233,N_12143,N_12090);
or U13234 (N_13234,N_12077,N_12836);
and U13235 (N_13235,N_12247,N_12669);
and U13236 (N_13236,N_12789,N_13002);
and U13237 (N_13237,N_12526,N_12760);
xor U13238 (N_13238,N_12549,N_12221);
or U13239 (N_13239,N_12217,N_12704);
nor U13240 (N_13240,N_12633,N_13054);
xnor U13241 (N_13241,N_12352,N_12010);
nor U13242 (N_13242,N_12585,N_12448);
xnor U13243 (N_13243,N_12178,N_12112);
xor U13244 (N_13244,N_12971,N_12511);
or U13245 (N_13245,N_12348,N_12034);
and U13246 (N_13246,N_12561,N_13194);
nand U13247 (N_13247,N_12173,N_12798);
nor U13248 (N_13248,N_12772,N_12360);
nand U13249 (N_13249,N_12932,N_12058);
or U13250 (N_13250,N_12913,N_12269);
and U13251 (N_13251,N_12119,N_12992);
and U13252 (N_13252,N_12693,N_12088);
and U13253 (N_13253,N_12673,N_12479);
and U13254 (N_13254,N_12267,N_12597);
or U13255 (N_13255,N_12442,N_13013);
nor U13256 (N_13256,N_13190,N_12022);
and U13257 (N_13257,N_13014,N_13163);
and U13258 (N_13258,N_12408,N_12838);
nor U13259 (N_13259,N_12722,N_12052);
xor U13260 (N_13260,N_13070,N_12309);
nor U13261 (N_13261,N_12101,N_12691);
or U13262 (N_13262,N_12033,N_12850);
xor U13263 (N_13263,N_12421,N_12365);
or U13264 (N_13264,N_12940,N_12684);
or U13265 (N_13265,N_12830,N_13161);
xnor U13266 (N_13266,N_12128,N_12236);
nor U13267 (N_13267,N_12319,N_12094);
nor U13268 (N_13268,N_12391,N_12628);
or U13269 (N_13269,N_12194,N_12124);
xnor U13270 (N_13270,N_12493,N_12476);
nor U13271 (N_13271,N_12106,N_12835);
nor U13272 (N_13272,N_12813,N_12400);
and U13273 (N_13273,N_12314,N_12842);
nand U13274 (N_13274,N_12831,N_12025);
nor U13275 (N_13275,N_13109,N_13153);
nor U13276 (N_13276,N_12420,N_12794);
nor U13277 (N_13277,N_12199,N_13100);
nand U13278 (N_13278,N_12230,N_13063);
xor U13279 (N_13279,N_12753,N_12244);
nand U13280 (N_13280,N_12845,N_13136);
nand U13281 (N_13281,N_12412,N_12424);
nand U13282 (N_13282,N_12667,N_12959);
or U13283 (N_13283,N_12955,N_12113);
and U13284 (N_13284,N_12026,N_12573);
nor U13285 (N_13285,N_12541,N_12924);
nor U13286 (N_13286,N_12713,N_12733);
or U13287 (N_13287,N_13168,N_12741);
xor U13288 (N_13288,N_12287,N_12748);
nand U13289 (N_13289,N_12261,N_12492);
nor U13290 (N_13290,N_12617,N_12596);
xor U13291 (N_13291,N_13150,N_12851);
or U13292 (N_13292,N_13120,N_13140);
or U13293 (N_13293,N_12038,N_12188);
nand U13294 (N_13294,N_13199,N_13186);
nand U13295 (N_13295,N_12288,N_12891);
or U13296 (N_13296,N_12787,N_12849);
nor U13297 (N_13297,N_13071,N_12884);
or U13298 (N_13298,N_12824,N_12984);
xnor U13299 (N_13299,N_13009,N_12774);
nor U13300 (N_13300,N_13026,N_12192);
or U13301 (N_13301,N_12096,N_12019);
nor U13302 (N_13302,N_12207,N_12627);
and U13303 (N_13303,N_12461,N_12127);
nor U13304 (N_13304,N_12517,N_12591);
xor U13305 (N_13305,N_12757,N_13126);
xnor U13306 (N_13306,N_12042,N_13084);
nand U13307 (N_13307,N_12556,N_12462);
or U13308 (N_13308,N_13103,N_12393);
nor U13309 (N_13309,N_12949,N_12793);
nor U13310 (N_13310,N_12266,N_12866);
nor U13311 (N_13311,N_12255,N_13106);
and U13312 (N_13312,N_12159,N_12806);
nand U13313 (N_13313,N_12874,N_12666);
and U13314 (N_13314,N_12780,N_12623);
xnor U13315 (N_13315,N_12870,N_12060);
and U13316 (N_13316,N_12289,N_12799);
nor U13317 (N_13317,N_12146,N_12506);
nor U13318 (N_13318,N_12383,N_12725);
nor U13319 (N_13319,N_12833,N_12281);
or U13320 (N_13320,N_12547,N_12140);
xnor U13321 (N_13321,N_12726,N_12957);
or U13322 (N_13322,N_13086,N_12116);
nor U13323 (N_13323,N_12014,N_12037);
nand U13324 (N_13324,N_12009,N_12858);
and U13325 (N_13325,N_12998,N_12446);
xnor U13326 (N_13326,N_12951,N_13169);
nor U13327 (N_13327,N_12555,N_12470);
nand U13328 (N_13328,N_12847,N_12432);
or U13329 (N_13329,N_12624,N_12953);
nand U13330 (N_13330,N_12484,N_12568);
and U13331 (N_13331,N_12705,N_12657);
xnor U13332 (N_13332,N_12241,N_12650);
and U13333 (N_13333,N_13105,N_12061);
nand U13334 (N_13334,N_12018,N_12346);
nand U13335 (N_13335,N_13158,N_12183);
or U13336 (N_13336,N_12353,N_12911);
or U13337 (N_13337,N_12877,N_12648);
nand U13338 (N_13338,N_12210,N_12945);
and U13339 (N_13339,N_13024,N_12734);
xnor U13340 (N_13340,N_12730,N_12064);
or U13341 (N_13341,N_12301,N_12156);
nand U13342 (N_13342,N_12177,N_12347);
and U13343 (N_13343,N_12862,N_13176);
nand U13344 (N_13344,N_12469,N_12214);
xor U13345 (N_13345,N_12770,N_12482);
nand U13346 (N_13346,N_12980,N_12515);
nand U13347 (N_13347,N_12439,N_12990);
or U13348 (N_13348,N_12222,N_12187);
or U13349 (N_13349,N_13021,N_12619);
or U13350 (N_13350,N_12599,N_12375);
xor U13351 (N_13351,N_12665,N_12456);
and U13352 (N_13352,N_12563,N_12191);
and U13353 (N_13353,N_12812,N_13018);
nand U13354 (N_13354,N_13113,N_12349);
nor U13355 (N_13355,N_13000,N_12890);
xnor U13356 (N_13356,N_12296,N_12546);
nor U13357 (N_13357,N_12708,N_13088);
or U13358 (N_13358,N_12175,N_13080);
nand U13359 (N_13359,N_12759,N_13164);
or U13360 (N_13360,N_12618,N_12724);
nand U13361 (N_13361,N_12963,N_12495);
or U13362 (N_13362,N_12047,N_12571);
nand U13363 (N_13363,N_12290,N_13130);
and U13364 (N_13364,N_12853,N_12987);
nand U13365 (N_13365,N_13073,N_12950);
or U13366 (N_13366,N_12438,N_13079);
nand U13367 (N_13367,N_12031,N_12567);
or U13368 (N_13368,N_13145,N_12262);
or U13369 (N_13369,N_12897,N_12141);
xnor U13370 (N_13370,N_12712,N_13053);
or U13371 (N_13371,N_13144,N_12467);
or U13372 (N_13372,N_12473,N_12674);
and U13373 (N_13373,N_12586,N_13143);
and U13374 (N_13374,N_12065,N_12941);
nand U13375 (N_13375,N_12108,N_12006);
nor U13376 (N_13376,N_13022,N_13132);
or U13377 (N_13377,N_12100,N_12076);
or U13378 (N_13378,N_12778,N_12416);
nand U13379 (N_13379,N_12279,N_13028);
nor U13380 (N_13380,N_12982,N_12195);
nand U13381 (N_13381,N_12810,N_13008);
and U13382 (N_13382,N_13001,N_12149);
and U13383 (N_13383,N_12259,N_13032);
nand U13384 (N_13384,N_12749,N_12082);
nor U13385 (N_13385,N_12132,N_13174);
nor U13386 (N_13386,N_13065,N_12562);
or U13387 (N_13387,N_13020,N_12218);
nor U13388 (N_13388,N_12369,N_12703);
or U13389 (N_13389,N_13193,N_12661);
xor U13390 (N_13390,N_12978,N_12538);
and U13391 (N_13391,N_12709,N_12514);
nor U13392 (N_13392,N_13154,N_12443);
xor U13393 (N_13393,N_12933,N_12512);
or U13394 (N_13394,N_12433,N_12671);
nand U13395 (N_13395,N_12331,N_13035);
and U13396 (N_13396,N_12121,N_13127);
or U13397 (N_13397,N_13087,N_12613);
and U13398 (N_13398,N_13122,N_12804);
and U13399 (N_13399,N_12027,N_13061);
nand U13400 (N_13400,N_13139,N_12999);
or U13401 (N_13401,N_12735,N_12086);
or U13402 (N_13402,N_13175,N_12109);
xnor U13403 (N_13403,N_12659,N_12916);
xnor U13404 (N_13404,N_12727,N_12854);
or U13405 (N_13405,N_12316,N_12300);
xor U13406 (N_13406,N_12543,N_12679);
and U13407 (N_13407,N_12685,N_12865);
or U13408 (N_13408,N_12828,N_12323);
xor U13409 (N_13409,N_12773,N_13025);
xor U13410 (N_13410,N_12522,N_12537);
nand U13411 (N_13411,N_13082,N_12996);
nor U13412 (N_13412,N_12251,N_12176);
or U13413 (N_13413,N_12423,N_12308);
nor U13414 (N_13414,N_12658,N_12212);
xor U13415 (N_13415,N_12294,N_12044);
and U13416 (N_13416,N_12604,N_12872);
or U13417 (N_13417,N_12459,N_12914);
xnor U13418 (N_13418,N_12767,N_12036);
nand U13419 (N_13419,N_13090,N_12404);
or U13420 (N_13420,N_12181,N_13119);
xnor U13421 (N_13421,N_12788,N_12122);
xor U13422 (N_13422,N_13078,N_12956);
nand U13423 (N_13423,N_12926,N_12826);
nor U13424 (N_13424,N_13066,N_12465);
or U13425 (N_13425,N_12868,N_12057);
xor U13426 (N_13426,N_12732,N_12046);
nor U13427 (N_13427,N_12343,N_12286);
or U13428 (N_13428,N_12496,N_12431);
nor U13429 (N_13429,N_12464,N_12907);
and U13430 (N_13430,N_13006,N_12736);
nand U13431 (N_13431,N_12606,N_12592);
or U13432 (N_13432,N_12946,N_13151);
or U13433 (N_13433,N_12455,N_13166);
nand U13434 (N_13434,N_12477,N_12073);
nand U13435 (N_13435,N_13064,N_12695);
nand U13436 (N_13436,N_12209,N_13137);
nand U13437 (N_13437,N_13074,N_12552);
xnor U13438 (N_13438,N_12584,N_12312);
nand U13439 (N_13439,N_12983,N_12821);
or U13440 (N_13440,N_12066,N_12644);
nand U13441 (N_13441,N_12534,N_13015);
nand U13442 (N_13442,N_12997,N_12553);
or U13443 (N_13443,N_12361,N_13165);
xnor U13444 (N_13444,N_12960,N_12802);
nor U13445 (N_13445,N_12340,N_12254);
xor U13446 (N_13446,N_12848,N_12702);
xnor U13447 (N_13447,N_12837,N_12342);
and U13448 (N_13448,N_12973,N_12087);
nor U13449 (N_13449,N_12670,N_12224);
nand U13450 (N_13450,N_12668,N_12489);
and U13451 (N_13451,N_13179,N_12557);
and U13452 (N_13452,N_12133,N_13045);
nor U13453 (N_13453,N_12452,N_12878);
or U13454 (N_13454,N_12021,N_12663);
nor U13455 (N_13455,N_12728,N_12413);
nor U13456 (N_13456,N_13012,N_12513);
or U13457 (N_13457,N_12485,N_12655);
nand U13458 (N_13458,N_12822,N_12776);
or U13459 (N_13459,N_12751,N_13017);
xor U13460 (N_13460,N_12234,N_12969);
nand U13461 (N_13461,N_12341,N_13192);
xnor U13462 (N_13462,N_12024,N_12339);
and U13463 (N_13463,N_13030,N_12677);
xnor U13464 (N_13464,N_12203,N_12252);
or U13465 (N_13465,N_12929,N_13170);
or U13466 (N_13466,N_13075,N_12167);
or U13467 (N_13467,N_13048,N_12602);
and U13468 (N_13468,N_12682,N_13141);
xnor U13469 (N_13469,N_12250,N_12499);
xor U13470 (N_13470,N_12790,N_12783);
xnor U13471 (N_13471,N_12427,N_12204);
xnor U13472 (N_13472,N_12921,N_12239);
nand U13473 (N_13473,N_12115,N_12809);
xor U13474 (N_13474,N_12102,N_13029);
nand U13475 (N_13475,N_12059,N_12808);
nand U13476 (N_13476,N_12598,N_12453);
xnor U13477 (N_13477,N_12324,N_12638);
xnor U13478 (N_13478,N_12213,N_13038);
nand U13479 (N_13479,N_13129,N_12357);
nor U13480 (N_13480,N_12754,N_12993);
and U13481 (N_13481,N_12880,N_12601);
or U13482 (N_13482,N_12917,N_12871);
nand U13483 (N_13483,N_12220,N_12766);
xor U13484 (N_13484,N_12518,N_13184);
nor U13485 (N_13485,N_12320,N_12136);
xnor U13486 (N_13486,N_12707,N_12426);
nor U13487 (N_13487,N_12762,N_12777);
xor U13488 (N_13488,N_12994,N_12719);
and U13489 (N_13489,N_12931,N_13036);
nor U13490 (N_13490,N_13117,N_12005);
nor U13491 (N_13491,N_12040,N_13092);
or U13492 (N_13492,N_12886,N_13155);
xnor U13493 (N_13493,N_12329,N_12937);
nor U13494 (N_13494,N_12468,N_13104);
nand U13495 (N_13495,N_12322,N_13102);
xor U13496 (N_13496,N_12680,N_12899);
nor U13497 (N_13497,N_12852,N_12265);
and U13498 (N_13498,N_12402,N_12976);
xor U13499 (N_13499,N_12559,N_12827);
nand U13500 (N_13500,N_12646,N_12359);
nor U13501 (N_13501,N_12539,N_12151);
nand U13502 (N_13502,N_12080,N_12717);
nand U13503 (N_13503,N_12417,N_12313);
nand U13504 (N_13504,N_12407,N_12750);
or U13505 (N_13505,N_12030,N_12889);
and U13506 (N_13506,N_12344,N_13114);
nand U13507 (N_13507,N_12111,N_12867);
xnor U13508 (N_13508,N_12284,N_12345);
and U13509 (N_13509,N_12362,N_13031);
xnor U13510 (N_13510,N_12942,N_12282);
xnor U13511 (N_13511,N_13094,N_12160);
and U13512 (N_13512,N_13124,N_13187);
or U13513 (N_13513,N_12273,N_12007);
xor U13514 (N_13514,N_12049,N_13131);
nand U13515 (N_13515,N_12846,N_13148);
nand U13516 (N_13516,N_12274,N_12904);
nor U13517 (N_13517,N_12458,N_12825);
xnor U13518 (N_13518,N_12215,N_13003);
nor U13519 (N_13519,N_12268,N_12488);
xnor U13520 (N_13520,N_13058,N_12356);
nor U13521 (N_13521,N_12249,N_12185);
nand U13522 (N_13522,N_12330,N_12743);
and U13523 (N_13523,N_12283,N_12013);
nor U13524 (N_13524,N_12502,N_12321);
or U13525 (N_13525,N_12139,N_12678);
nand U13526 (N_13526,N_12130,N_12487);
nor U13527 (N_13527,N_12792,N_12480);
nand U13528 (N_13528,N_12686,N_12639);
nor U13529 (N_13529,N_13098,N_12118);
nand U13530 (N_13530,N_12965,N_12711);
xnor U13531 (N_13531,N_12164,N_12263);
or U13532 (N_13532,N_12656,N_12875);
and U13533 (N_13533,N_12197,N_12962);
or U13534 (N_13534,N_12841,N_13027);
nor U13535 (N_13535,N_12723,N_12003);
nand U13536 (N_13536,N_12739,N_12936);
and U13537 (N_13537,N_12554,N_12995);
nor U13538 (N_13538,N_13146,N_12582);
nand U13539 (N_13539,N_12530,N_12698);
nand U13540 (N_13540,N_12781,N_12257);
or U13541 (N_13541,N_12358,N_12523);
nor U13542 (N_13542,N_12070,N_13111);
xor U13543 (N_13543,N_12720,N_12944);
and U13544 (N_13544,N_13196,N_12075);
xor U13545 (N_13545,N_12947,N_12232);
and U13546 (N_13546,N_12486,N_12310);
and U13547 (N_13547,N_12908,N_12233);
or U13548 (N_13548,N_13178,N_12107);
and U13549 (N_13549,N_12071,N_12763);
nor U13550 (N_13550,N_12299,N_12228);
or U13551 (N_13551,N_12395,N_12169);
nand U13552 (N_13552,N_12903,N_12039);
or U13553 (N_13553,N_13142,N_13052);
nand U13554 (N_13554,N_12894,N_12954);
nor U13555 (N_13555,N_12008,N_12979);
nor U13556 (N_13556,N_13042,N_12654);
nor U13557 (N_13557,N_12634,N_12576);
and U13558 (N_13558,N_12385,N_12860);
or U13559 (N_13559,N_12387,N_12883);
and U13560 (N_13560,N_12147,N_12935);
or U13561 (N_13561,N_12608,N_12681);
or U13562 (N_13562,N_12418,N_12326);
nand U13563 (N_13563,N_12888,N_12869);
or U13564 (N_13564,N_12533,N_12202);
xnor U13565 (N_13565,N_12246,N_12354);
xnor U13566 (N_13566,N_12114,N_12784);
and U13567 (N_13567,N_12815,N_12105);
nand U13568 (N_13568,N_12505,N_12093);
nand U13569 (N_13569,N_13077,N_12803);
and U13570 (N_13570,N_12380,N_12531);
nand U13571 (N_13571,N_12264,N_12307);
nand U13572 (N_13572,N_12672,N_13044);
or U13573 (N_13573,N_12491,N_12068);
nor U13574 (N_13574,N_12165,N_12148);
and U13575 (N_13575,N_12647,N_12016);
nor U13576 (N_13576,N_12004,N_13167);
nor U13577 (N_13577,N_12398,N_12581);
nand U13578 (N_13578,N_13116,N_13040);
or U13579 (N_13579,N_13010,N_12260);
nand U13580 (N_13580,N_12516,N_12752);
nand U13581 (N_13581,N_12243,N_12721);
and U13582 (N_13582,N_12297,N_12829);
nor U13583 (N_13583,N_12524,N_12245);
nor U13584 (N_13584,N_12399,N_12182);
nand U13585 (N_13585,N_12688,N_12863);
nor U13586 (N_13586,N_12306,N_12508);
or U13587 (N_13587,N_12607,N_13060);
and U13588 (N_13588,N_12892,N_12174);
xor U13589 (N_13589,N_12621,N_12614);
nor U13590 (N_13590,N_12028,N_12928);
nand U13591 (N_13591,N_12740,N_12769);
nor U13592 (N_13592,N_12961,N_13096);
and U13593 (N_13593,N_12390,N_12536);
xor U13594 (N_13594,N_12304,N_12943);
and U13595 (N_13595,N_12079,N_12434);
or U13596 (N_13596,N_13110,N_12409);
nand U13597 (N_13597,N_12905,N_12653);
nor U13598 (N_13598,N_12474,N_12560);
xnor U13599 (N_13599,N_12460,N_12490);
or U13600 (N_13600,N_13059,N_13157);
or U13601 (N_13601,N_12305,N_12700);
xor U13602 (N_13602,N_13198,N_12651);
and U13603 (N_13603,N_12612,N_12163);
or U13604 (N_13604,N_12873,N_12095);
and U13605 (N_13605,N_12097,N_12231);
nand U13606 (N_13606,N_12336,N_13195);
and U13607 (N_13607,N_12504,N_12258);
nand U13608 (N_13608,N_12861,N_12225);
nand U13609 (N_13609,N_12415,N_12364);
and U13610 (N_13610,N_12817,N_12574);
nand U13611 (N_13611,N_12374,N_12823);
xnor U13612 (N_13612,N_12881,N_12782);
and U13613 (N_13613,N_12832,N_12367);
xor U13614 (N_13614,N_12200,N_12170);
xor U13615 (N_13615,N_12447,N_12451);
xor U13616 (N_13616,N_12089,N_12002);
xor U13617 (N_13617,N_12968,N_13081);
nand U13618 (N_13618,N_12967,N_12915);
xor U13619 (N_13619,N_12363,N_12755);
nor U13620 (N_13620,N_12270,N_13095);
xnor U13621 (N_13621,N_13123,N_13016);
and U13622 (N_13622,N_13050,N_12298);
and U13623 (N_13623,N_12172,N_12205);
nor U13624 (N_13624,N_12746,N_13067);
and U13625 (N_13625,N_12179,N_12229);
and U13626 (N_13626,N_12816,N_12419);
or U13627 (N_13627,N_12575,N_12050);
xor U13628 (N_13628,N_12758,N_12503);
or U13629 (N_13629,N_12664,N_12595);
xor U13630 (N_13630,N_12626,N_12069);
nor U13631 (N_13631,N_13162,N_12742);
or U13632 (N_13632,N_12548,N_12876);
and U13633 (N_13633,N_13134,N_13183);
nand U13634 (N_13634,N_12615,N_12227);
and U13635 (N_13635,N_13133,N_12198);
xnor U13636 (N_13636,N_12952,N_12764);
and U13637 (N_13637,N_12683,N_12193);
or U13638 (N_13638,N_13019,N_12898);
or U13639 (N_13639,N_12922,N_13101);
or U13640 (N_13640,N_12925,N_12466);
nand U13641 (N_13641,N_12551,N_12814);
nand U13642 (N_13642,N_12501,N_13121);
xnor U13643 (N_13643,N_12062,N_12237);
xnor U13644 (N_13644,N_13037,N_12129);
or U13645 (N_13645,N_12662,N_13189);
nand U13646 (N_13646,N_12392,N_12535);
and U13647 (N_13647,N_12544,N_13051);
nor U13648 (N_13648,N_12795,N_12223);
or U13649 (N_13649,N_12520,N_12565);
nor U13650 (N_13650,N_12622,N_12428);
or U13651 (N_13651,N_12893,N_12939);
or U13652 (N_13652,N_12403,N_12098);
nor U13653 (N_13653,N_12745,N_12190);
and U13654 (N_13654,N_12053,N_12839);
nand U13655 (N_13655,N_12441,N_12401);
or U13656 (N_13656,N_12189,N_12253);
and U13657 (N_13657,N_13068,N_12609);
or U13658 (N_13658,N_12509,N_12370);
xor U13659 (N_13659,N_12396,N_12389);
xnor U13660 (N_13660,N_12085,N_12012);
nor U13661 (N_13661,N_12463,N_13039);
and U13662 (N_13662,N_12964,N_13171);
nand U13663 (N_13663,N_12368,N_12475);
nand U13664 (N_13664,N_12775,N_12000);
or U13665 (N_13665,N_12919,N_12859);
and U13666 (N_13666,N_12840,N_12162);
and U13667 (N_13667,N_12593,N_12481);
and U13668 (N_13668,N_12055,N_12271);
or U13669 (N_13669,N_12272,N_12497);
and U13670 (N_13670,N_12818,N_12620);
nand U13671 (N_13671,N_13156,N_12280);
xnor U13672 (N_13672,N_12048,N_12587);
xor U13673 (N_13673,N_12152,N_12786);
and U13674 (N_13674,N_12910,N_12701);
nand U13675 (N_13675,N_12315,N_12590);
or U13676 (N_13676,N_13049,N_12570);
nand U13677 (N_13677,N_12337,N_12642);
or U13678 (N_13678,N_12494,N_13147);
xor U13679 (N_13679,N_12333,N_13083);
and U13680 (N_13680,N_12603,N_12275);
nor U13681 (N_13681,N_13191,N_12991);
or U13682 (N_13682,N_12938,N_13108);
nand U13683 (N_13683,N_12184,N_12366);
xor U13684 (N_13684,N_12747,N_12986);
nor U13685 (N_13685,N_12715,N_13125);
nand U13686 (N_13686,N_12110,N_12472);
and U13687 (N_13687,N_13160,N_12660);
and U13688 (N_13688,N_12011,N_12731);
or U13689 (N_13689,N_12457,N_12635);
xor U13690 (N_13690,N_12171,N_13185);
nand U13691 (N_13691,N_12043,N_12600);
nor U13692 (N_13692,N_12032,N_13112);
nand U13693 (N_13693,N_12437,N_12558);
or U13694 (N_13694,N_12694,N_12525);
nor U13695 (N_13695,N_12902,N_12120);
nor U13696 (N_13696,N_12706,N_12616);
and U13697 (N_13697,N_13138,N_12302);
nor U13698 (N_13698,N_12729,N_12765);
nand U13699 (N_13699,N_12153,N_12631);
and U13700 (N_13700,N_12918,N_12791);
xor U13701 (N_13701,N_12411,N_12293);
or U13702 (N_13702,N_12444,N_12500);
nor U13703 (N_13703,N_12410,N_12652);
nand U13704 (N_13704,N_12471,N_12081);
nor U13705 (N_13705,N_12083,N_12625);
and U13706 (N_13706,N_13099,N_13197);
and U13707 (N_13707,N_12569,N_12564);
nor U13708 (N_13708,N_12074,N_13057);
nand U13709 (N_13709,N_12425,N_12248);
or U13710 (N_13710,N_12478,N_13107);
nand U13711 (N_13711,N_12292,N_12796);
nor U13712 (N_13712,N_12528,N_12927);
and U13713 (N_13713,N_12295,N_12714);
and U13714 (N_13714,N_12355,N_12887);
xnor U13715 (N_13715,N_12150,N_12440);
or U13716 (N_13716,N_13173,N_12540);
nand U13717 (N_13717,N_12078,N_12882);
or U13718 (N_13718,N_12589,N_12201);
and U13719 (N_13719,N_12689,N_12158);
or U13720 (N_13720,N_13159,N_12072);
xnor U13721 (N_13721,N_12180,N_12744);
or U13722 (N_13722,N_13046,N_12843);
nand U13723 (N_13723,N_12327,N_12332);
or U13724 (N_13724,N_12168,N_13043);
nor U13725 (N_13725,N_12636,N_12800);
xor U13726 (N_13726,N_12242,N_12906);
or U13727 (N_13727,N_12588,N_12373);
nand U13728 (N_13728,N_12510,N_12449);
xor U13729 (N_13729,N_12696,N_12023);
nand U13730 (N_13730,N_13023,N_12125);
xnor U13731 (N_13731,N_12015,N_12436);
or U13732 (N_13732,N_13011,N_12161);
or U13733 (N_13733,N_13033,N_12208);
nor U13734 (N_13734,N_12923,N_12117);
nor U13735 (N_13735,N_12630,N_12126);
nor U13736 (N_13736,N_12864,N_12632);
nor U13737 (N_13737,N_12855,N_12041);
nand U13738 (N_13738,N_13089,N_13180);
and U13739 (N_13739,N_12020,N_12985);
nor U13740 (N_13740,N_12137,N_12084);
nor U13741 (N_13741,N_12388,N_12067);
or U13742 (N_13742,N_12583,N_13118);
nand U13743 (N_13743,N_12801,N_12697);
xnor U13744 (N_13744,N_12895,N_12579);
and U13745 (N_13745,N_12756,N_12157);
or U13746 (N_13746,N_12820,N_13091);
and U13747 (N_13747,N_12507,N_12029);
nand U13748 (N_13748,N_12219,N_12580);
and U13749 (N_13749,N_12610,N_12351);
nor U13750 (N_13750,N_12056,N_12372);
nand U13751 (N_13751,N_12629,N_12948);
nor U13752 (N_13752,N_12276,N_12145);
nand U13753 (N_13753,N_12811,N_12771);
xnor U13754 (N_13754,N_12885,N_12350);
or U13755 (N_13755,N_12142,N_12856);
nand U13756 (N_13756,N_12134,N_12206);
nand U13757 (N_13757,N_12371,N_12529);
or U13758 (N_13758,N_13005,N_12527);
xor U13759 (N_13759,N_12970,N_12761);
and U13760 (N_13760,N_12879,N_12896);
and U13761 (N_13761,N_13097,N_12386);
nor U13762 (N_13762,N_12285,N_12819);
nand U13763 (N_13763,N_12640,N_13041);
and U13764 (N_13764,N_12641,N_12779);
nand U13765 (N_13765,N_12857,N_12566);
nand U13766 (N_13766,N_12699,N_12291);
nor U13767 (N_13767,N_12138,N_12718);
xor U13768 (N_13768,N_12972,N_12382);
and U13769 (N_13769,N_12690,N_12154);
and U13770 (N_13770,N_12303,N_12797);
xnor U13771 (N_13771,N_13004,N_12381);
or U13772 (N_13772,N_12687,N_12123);
nor U13773 (N_13773,N_12785,N_12166);
and U13774 (N_13774,N_12384,N_12542);
and U13775 (N_13775,N_12605,N_13072);
and U13776 (N_13776,N_12550,N_13172);
xnor U13777 (N_13777,N_12317,N_12737);
nor U13778 (N_13778,N_12981,N_12637);
and U13779 (N_13779,N_12054,N_12643);
or U13780 (N_13780,N_12216,N_12934);
xnor U13781 (N_13781,N_12104,N_12483);
nor U13782 (N_13782,N_13128,N_13056);
nor U13783 (N_13783,N_12135,N_12379);
or U13784 (N_13784,N_12920,N_12454);
xnor U13785 (N_13785,N_13055,N_12277);
nor U13786 (N_13786,N_12577,N_12131);
or U13787 (N_13787,N_13034,N_12186);
nand U13788 (N_13788,N_12240,N_13177);
xnor U13789 (N_13789,N_12594,N_12378);
and U13790 (N_13790,N_12645,N_12572);
nand U13791 (N_13791,N_12966,N_13085);
nand U13792 (N_13792,N_12844,N_12091);
and U13793 (N_13793,N_12738,N_12035);
nor U13794 (N_13794,N_13181,N_12430);
and U13795 (N_13795,N_12256,N_12063);
xnor U13796 (N_13796,N_12807,N_12611);
or U13797 (N_13797,N_12001,N_12521);
nand U13798 (N_13798,N_12092,N_12318);
or U13799 (N_13799,N_12716,N_12768);
and U13800 (N_13800,N_12402,N_12547);
or U13801 (N_13801,N_12437,N_12955);
nand U13802 (N_13802,N_13104,N_12499);
and U13803 (N_13803,N_12605,N_12139);
xor U13804 (N_13804,N_12760,N_12813);
and U13805 (N_13805,N_12196,N_12484);
nor U13806 (N_13806,N_12080,N_12210);
xnor U13807 (N_13807,N_13183,N_12920);
or U13808 (N_13808,N_12307,N_13101);
nand U13809 (N_13809,N_13132,N_12556);
nor U13810 (N_13810,N_12407,N_12409);
xor U13811 (N_13811,N_12210,N_12620);
nor U13812 (N_13812,N_12976,N_12592);
xor U13813 (N_13813,N_12175,N_13014);
nor U13814 (N_13814,N_12289,N_12229);
xor U13815 (N_13815,N_12251,N_12778);
nor U13816 (N_13816,N_12558,N_12863);
or U13817 (N_13817,N_12589,N_12324);
nand U13818 (N_13818,N_12858,N_12945);
nand U13819 (N_13819,N_12377,N_12247);
nor U13820 (N_13820,N_12165,N_13139);
nand U13821 (N_13821,N_12554,N_12851);
nor U13822 (N_13822,N_12010,N_13188);
xnor U13823 (N_13823,N_12405,N_12945);
xnor U13824 (N_13824,N_12990,N_12602);
nand U13825 (N_13825,N_12881,N_12277);
nand U13826 (N_13826,N_13035,N_13067);
nand U13827 (N_13827,N_12474,N_12887);
xor U13828 (N_13828,N_12113,N_12248);
nor U13829 (N_13829,N_12529,N_12639);
xnor U13830 (N_13830,N_13174,N_12478);
and U13831 (N_13831,N_12651,N_12218);
or U13832 (N_13832,N_13036,N_12253);
nand U13833 (N_13833,N_12168,N_12381);
or U13834 (N_13834,N_12395,N_12742);
and U13835 (N_13835,N_13199,N_13033);
nand U13836 (N_13836,N_12576,N_13144);
and U13837 (N_13837,N_12349,N_12360);
nor U13838 (N_13838,N_12667,N_12110);
or U13839 (N_13839,N_12549,N_12141);
and U13840 (N_13840,N_12198,N_12720);
nor U13841 (N_13841,N_12817,N_12921);
nand U13842 (N_13842,N_12652,N_12544);
and U13843 (N_13843,N_12958,N_12784);
xnor U13844 (N_13844,N_12020,N_12612);
xnor U13845 (N_13845,N_13140,N_13190);
nand U13846 (N_13846,N_12598,N_13035);
nand U13847 (N_13847,N_12883,N_12603);
nand U13848 (N_13848,N_12659,N_12533);
xnor U13849 (N_13849,N_12545,N_13173);
nand U13850 (N_13850,N_12126,N_12148);
nand U13851 (N_13851,N_12185,N_12012);
and U13852 (N_13852,N_12496,N_12011);
or U13853 (N_13853,N_12082,N_12183);
xnor U13854 (N_13854,N_12735,N_12850);
and U13855 (N_13855,N_12365,N_12408);
and U13856 (N_13856,N_13033,N_12470);
nand U13857 (N_13857,N_12853,N_12526);
or U13858 (N_13858,N_13026,N_12101);
xor U13859 (N_13859,N_12620,N_13003);
nor U13860 (N_13860,N_12609,N_12582);
nand U13861 (N_13861,N_12859,N_12791);
or U13862 (N_13862,N_12405,N_12077);
or U13863 (N_13863,N_12234,N_12662);
and U13864 (N_13864,N_12708,N_12138);
nand U13865 (N_13865,N_12095,N_12914);
or U13866 (N_13866,N_12099,N_12264);
or U13867 (N_13867,N_12777,N_12948);
xnor U13868 (N_13868,N_12168,N_12829);
or U13869 (N_13869,N_12906,N_12487);
or U13870 (N_13870,N_12035,N_12781);
and U13871 (N_13871,N_13031,N_12666);
nand U13872 (N_13872,N_12936,N_12821);
xnor U13873 (N_13873,N_12788,N_12266);
nor U13874 (N_13874,N_13032,N_12016);
nand U13875 (N_13875,N_12320,N_13072);
or U13876 (N_13876,N_12776,N_12304);
or U13877 (N_13877,N_12425,N_13074);
nand U13878 (N_13878,N_12270,N_12862);
nor U13879 (N_13879,N_12152,N_12809);
and U13880 (N_13880,N_12909,N_12834);
nor U13881 (N_13881,N_12394,N_12462);
or U13882 (N_13882,N_12246,N_12881);
or U13883 (N_13883,N_12985,N_12061);
xnor U13884 (N_13884,N_12517,N_13091);
and U13885 (N_13885,N_12218,N_12366);
xnor U13886 (N_13886,N_12217,N_12677);
nand U13887 (N_13887,N_12452,N_12715);
nand U13888 (N_13888,N_13079,N_12050);
nor U13889 (N_13889,N_12596,N_12498);
and U13890 (N_13890,N_12328,N_12130);
nand U13891 (N_13891,N_12144,N_12614);
nor U13892 (N_13892,N_12307,N_12856);
or U13893 (N_13893,N_13064,N_12206);
xor U13894 (N_13894,N_13017,N_12383);
and U13895 (N_13895,N_12985,N_12439);
xnor U13896 (N_13896,N_12019,N_12476);
and U13897 (N_13897,N_12158,N_13119);
xor U13898 (N_13898,N_12678,N_12745);
or U13899 (N_13899,N_12590,N_12692);
xnor U13900 (N_13900,N_12283,N_12251);
and U13901 (N_13901,N_12233,N_12809);
xor U13902 (N_13902,N_13171,N_12180);
xor U13903 (N_13903,N_13134,N_12760);
nor U13904 (N_13904,N_12747,N_12490);
nor U13905 (N_13905,N_12628,N_13130);
or U13906 (N_13906,N_13061,N_12142);
or U13907 (N_13907,N_12963,N_13083);
nand U13908 (N_13908,N_13189,N_12673);
nor U13909 (N_13909,N_12305,N_12142);
or U13910 (N_13910,N_12901,N_12922);
or U13911 (N_13911,N_13191,N_12366);
or U13912 (N_13912,N_13185,N_12003);
or U13913 (N_13913,N_13099,N_12931);
xnor U13914 (N_13914,N_12100,N_12652);
and U13915 (N_13915,N_12953,N_12871);
or U13916 (N_13916,N_12151,N_12787);
and U13917 (N_13917,N_13039,N_12158);
nand U13918 (N_13918,N_12508,N_12105);
or U13919 (N_13919,N_12082,N_13169);
nor U13920 (N_13920,N_13092,N_13043);
and U13921 (N_13921,N_12494,N_12124);
nand U13922 (N_13922,N_12624,N_12231);
xnor U13923 (N_13923,N_12213,N_12240);
nand U13924 (N_13924,N_12651,N_12190);
or U13925 (N_13925,N_12993,N_12034);
nor U13926 (N_13926,N_13141,N_12015);
and U13927 (N_13927,N_12827,N_12370);
nand U13928 (N_13928,N_12592,N_12859);
or U13929 (N_13929,N_12319,N_12996);
nand U13930 (N_13930,N_12500,N_12971);
xnor U13931 (N_13931,N_12368,N_12572);
or U13932 (N_13932,N_12012,N_13048);
nand U13933 (N_13933,N_12865,N_13062);
and U13934 (N_13934,N_12727,N_12913);
or U13935 (N_13935,N_12697,N_12591);
and U13936 (N_13936,N_12148,N_12423);
nor U13937 (N_13937,N_12291,N_12165);
nand U13938 (N_13938,N_12618,N_12814);
or U13939 (N_13939,N_12792,N_12166);
nor U13940 (N_13940,N_12401,N_12506);
xor U13941 (N_13941,N_12598,N_12532);
or U13942 (N_13942,N_12510,N_12219);
or U13943 (N_13943,N_12805,N_13081);
and U13944 (N_13944,N_12444,N_12721);
xor U13945 (N_13945,N_12416,N_13061);
or U13946 (N_13946,N_12821,N_12041);
or U13947 (N_13947,N_12223,N_12030);
nor U13948 (N_13948,N_13137,N_12657);
nand U13949 (N_13949,N_13194,N_12810);
or U13950 (N_13950,N_13146,N_12527);
and U13951 (N_13951,N_12972,N_12664);
and U13952 (N_13952,N_12236,N_12071);
and U13953 (N_13953,N_12159,N_12360);
nand U13954 (N_13954,N_12574,N_12619);
nand U13955 (N_13955,N_12167,N_12044);
nor U13956 (N_13956,N_12867,N_12900);
xor U13957 (N_13957,N_12008,N_12974);
nor U13958 (N_13958,N_12361,N_12616);
and U13959 (N_13959,N_12257,N_12489);
or U13960 (N_13960,N_12881,N_12315);
and U13961 (N_13961,N_12778,N_12519);
xor U13962 (N_13962,N_12356,N_12573);
nand U13963 (N_13963,N_12177,N_12666);
and U13964 (N_13964,N_12076,N_13045);
or U13965 (N_13965,N_12504,N_13134);
xnor U13966 (N_13966,N_13101,N_13031);
xor U13967 (N_13967,N_13098,N_12428);
nand U13968 (N_13968,N_12142,N_13168);
nor U13969 (N_13969,N_12008,N_12273);
xnor U13970 (N_13970,N_12057,N_13124);
or U13971 (N_13971,N_13085,N_12695);
and U13972 (N_13972,N_12079,N_12923);
nand U13973 (N_13973,N_12528,N_12360);
nor U13974 (N_13974,N_13138,N_12376);
nor U13975 (N_13975,N_12782,N_12446);
nor U13976 (N_13976,N_12332,N_12046);
or U13977 (N_13977,N_12478,N_12324);
nand U13978 (N_13978,N_12080,N_12826);
or U13979 (N_13979,N_12521,N_12456);
nand U13980 (N_13980,N_12963,N_12481);
and U13981 (N_13981,N_12556,N_12073);
xor U13982 (N_13982,N_12714,N_12544);
nand U13983 (N_13983,N_12425,N_12671);
nor U13984 (N_13984,N_13145,N_12995);
and U13985 (N_13985,N_13135,N_12631);
and U13986 (N_13986,N_12187,N_12273);
nand U13987 (N_13987,N_12829,N_12096);
xor U13988 (N_13988,N_12140,N_12057);
nand U13989 (N_13989,N_13095,N_12019);
xnor U13990 (N_13990,N_12925,N_12364);
xor U13991 (N_13991,N_13181,N_12899);
nor U13992 (N_13992,N_12984,N_12393);
xnor U13993 (N_13993,N_12361,N_12352);
or U13994 (N_13994,N_12647,N_12433);
nand U13995 (N_13995,N_12325,N_12425);
xor U13996 (N_13996,N_12611,N_12613);
nor U13997 (N_13997,N_13082,N_12340);
nor U13998 (N_13998,N_12735,N_12621);
or U13999 (N_13999,N_12876,N_12798);
and U14000 (N_14000,N_13035,N_12654);
nor U14001 (N_14001,N_12496,N_12575);
nor U14002 (N_14002,N_12164,N_12313);
or U14003 (N_14003,N_12314,N_12397);
or U14004 (N_14004,N_12252,N_12330);
nand U14005 (N_14005,N_12809,N_12680);
or U14006 (N_14006,N_13164,N_12212);
and U14007 (N_14007,N_12188,N_12861);
and U14008 (N_14008,N_12174,N_12786);
xnor U14009 (N_14009,N_12733,N_12543);
xnor U14010 (N_14010,N_12296,N_12265);
and U14011 (N_14011,N_13048,N_12640);
and U14012 (N_14012,N_12150,N_13167);
xnor U14013 (N_14013,N_13138,N_12575);
xor U14014 (N_14014,N_13090,N_12643);
nor U14015 (N_14015,N_12929,N_12888);
nor U14016 (N_14016,N_12349,N_12576);
and U14017 (N_14017,N_13049,N_12668);
nor U14018 (N_14018,N_12019,N_12682);
nor U14019 (N_14019,N_12491,N_12634);
and U14020 (N_14020,N_12310,N_12510);
or U14021 (N_14021,N_12306,N_13062);
or U14022 (N_14022,N_12513,N_13144);
xnor U14023 (N_14023,N_12829,N_13181);
xor U14024 (N_14024,N_12347,N_13088);
xnor U14025 (N_14025,N_13046,N_12020);
and U14026 (N_14026,N_12159,N_12884);
or U14027 (N_14027,N_12099,N_12908);
or U14028 (N_14028,N_13122,N_12417);
and U14029 (N_14029,N_12309,N_12245);
and U14030 (N_14030,N_12777,N_12352);
xnor U14031 (N_14031,N_12566,N_13090);
or U14032 (N_14032,N_12444,N_12766);
nand U14033 (N_14033,N_12254,N_12371);
xnor U14034 (N_14034,N_12388,N_12521);
or U14035 (N_14035,N_12233,N_13057);
or U14036 (N_14036,N_12967,N_12210);
or U14037 (N_14037,N_12480,N_12623);
and U14038 (N_14038,N_12417,N_12539);
or U14039 (N_14039,N_12764,N_12820);
nor U14040 (N_14040,N_12817,N_13058);
xnor U14041 (N_14041,N_12945,N_12819);
nor U14042 (N_14042,N_12078,N_12218);
or U14043 (N_14043,N_13023,N_12780);
xnor U14044 (N_14044,N_12189,N_12305);
or U14045 (N_14045,N_12706,N_13098);
and U14046 (N_14046,N_12542,N_12706);
and U14047 (N_14047,N_13176,N_12643);
or U14048 (N_14048,N_12320,N_12680);
and U14049 (N_14049,N_12712,N_12798);
or U14050 (N_14050,N_13139,N_12665);
nand U14051 (N_14051,N_12826,N_12869);
nand U14052 (N_14052,N_12832,N_12064);
nor U14053 (N_14053,N_12921,N_12491);
nand U14054 (N_14054,N_12897,N_12472);
or U14055 (N_14055,N_12282,N_12434);
nand U14056 (N_14056,N_12478,N_12173);
and U14057 (N_14057,N_12823,N_12891);
xor U14058 (N_14058,N_12454,N_12447);
and U14059 (N_14059,N_12186,N_13096);
xnor U14060 (N_14060,N_13166,N_13187);
nand U14061 (N_14061,N_13128,N_13187);
nand U14062 (N_14062,N_12745,N_12442);
or U14063 (N_14063,N_13063,N_12553);
and U14064 (N_14064,N_12857,N_12590);
and U14065 (N_14065,N_12140,N_12286);
and U14066 (N_14066,N_12240,N_12457);
and U14067 (N_14067,N_13128,N_12154);
or U14068 (N_14068,N_13103,N_12054);
xnor U14069 (N_14069,N_12571,N_12587);
nor U14070 (N_14070,N_12128,N_12889);
and U14071 (N_14071,N_12887,N_13137);
and U14072 (N_14072,N_12466,N_12937);
and U14073 (N_14073,N_12321,N_12406);
or U14074 (N_14074,N_12409,N_12481);
nor U14075 (N_14075,N_13055,N_12475);
xnor U14076 (N_14076,N_12485,N_12519);
and U14077 (N_14077,N_12347,N_12521);
nand U14078 (N_14078,N_12023,N_12733);
and U14079 (N_14079,N_12896,N_12018);
or U14080 (N_14080,N_13159,N_13058);
or U14081 (N_14081,N_12315,N_13006);
xor U14082 (N_14082,N_13098,N_13137);
nand U14083 (N_14083,N_13107,N_12572);
or U14084 (N_14084,N_12900,N_12858);
nor U14085 (N_14085,N_13092,N_12993);
or U14086 (N_14086,N_12856,N_12287);
xnor U14087 (N_14087,N_12599,N_12318);
xnor U14088 (N_14088,N_13016,N_12438);
xor U14089 (N_14089,N_12193,N_12784);
xnor U14090 (N_14090,N_12384,N_12960);
nand U14091 (N_14091,N_12820,N_12248);
nor U14092 (N_14092,N_12744,N_12956);
or U14093 (N_14093,N_12323,N_12379);
or U14094 (N_14094,N_12209,N_12361);
and U14095 (N_14095,N_12144,N_12797);
xor U14096 (N_14096,N_12144,N_12840);
or U14097 (N_14097,N_12178,N_12737);
nor U14098 (N_14098,N_12154,N_12480);
nor U14099 (N_14099,N_12187,N_12161);
or U14100 (N_14100,N_12840,N_12146);
xor U14101 (N_14101,N_12117,N_12173);
xor U14102 (N_14102,N_12850,N_12209);
and U14103 (N_14103,N_12505,N_12348);
nor U14104 (N_14104,N_12823,N_13071);
nor U14105 (N_14105,N_12775,N_12433);
and U14106 (N_14106,N_12949,N_12265);
or U14107 (N_14107,N_12940,N_12954);
nand U14108 (N_14108,N_12517,N_12313);
nor U14109 (N_14109,N_12281,N_12748);
nor U14110 (N_14110,N_12722,N_12651);
xnor U14111 (N_14111,N_12652,N_12178);
and U14112 (N_14112,N_12737,N_13109);
or U14113 (N_14113,N_12208,N_13064);
xnor U14114 (N_14114,N_13099,N_12461);
and U14115 (N_14115,N_13028,N_13017);
or U14116 (N_14116,N_12175,N_12097);
and U14117 (N_14117,N_12709,N_12543);
or U14118 (N_14118,N_13164,N_12368);
nor U14119 (N_14119,N_12750,N_12217);
nor U14120 (N_14120,N_12233,N_12036);
or U14121 (N_14121,N_12808,N_12684);
nor U14122 (N_14122,N_12170,N_12156);
nand U14123 (N_14123,N_12656,N_12697);
nor U14124 (N_14124,N_12416,N_12548);
and U14125 (N_14125,N_12700,N_12916);
and U14126 (N_14126,N_12362,N_12575);
xor U14127 (N_14127,N_13114,N_12016);
xor U14128 (N_14128,N_13182,N_12408);
or U14129 (N_14129,N_12108,N_12201);
xnor U14130 (N_14130,N_13190,N_12800);
and U14131 (N_14131,N_12896,N_12602);
and U14132 (N_14132,N_13010,N_12915);
nand U14133 (N_14133,N_12017,N_12613);
nand U14134 (N_14134,N_12593,N_12873);
xor U14135 (N_14135,N_12540,N_13112);
and U14136 (N_14136,N_12544,N_12227);
or U14137 (N_14137,N_12440,N_13071);
nor U14138 (N_14138,N_12190,N_13092);
or U14139 (N_14139,N_12162,N_13154);
or U14140 (N_14140,N_12258,N_13103);
nand U14141 (N_14141,N_12425,N_12684);
and U14142 (N_14142,N_12919,N_13106);
nor U14143 (N_14143,N_12829,N_12478);
or U14144 (N_14144,N_12948,N_12224);
or U14145 (N_14145,N_12017,N_12992);
or U14146 (N_14146,N_12299,N_12041);
and U14147 (N_14147,N_12940,N_12056);
xor U14148 (N_14148,N_12469,N_12850);
and U14149 (N_14149,N_12747,N_12579);
and U14150 (N_14150,N_12902,N_13119);
xor U14151 (N_14151,N_12003,N_12653);
nand U14152 (N_14152,N_12263,N_12007);
or U14153 (N_14153,N_12101,N_12013);
nor U14154 (N_14154,N_12514,N_13072);
xnor U14155 (N_14155,N_12353,N_13112);
nor U14156 (N_14156,N_12345,N_12533);
and U14157 (N_14157,N_12707,N_12634);
xor U14158 (N_14158,N_12441,N_13159);
and U14159 (N_14159,N_12318,N_12498);
xor U14160 (N_14160,N_13162,N_13167);
nand U14161 (N_14161,N_12160,N_12755);
and U14162 (N_14162,N_12508,N_12753);
or U14163 (N_14163,N_12306,N_13131);
and U14164 (N_14164,N_12901,N_12771);
nor U14165 (N_14165,N_13137,N_12144);
and U14166 (N_14166,N_12861,N_12956);
and U14167 (N_14167,N_12802,N_13120);
nor U14168 (N_14168,N_12258,N_12392);
and U14169 (N_14169,N_12971,N_12781);
xnor U14170 (N_14170,N_12331,N_12191);
xor U14171 (N_14171,N_13005,N_12162);
and U14172 (N_14172,N_12018,N_12743);
and U14173 (N_14173,N_12577,N_12920);
nor U14174 (N_14174,N_12660,N_12362);
or U14175 (N_14175,N_12932,N_13146);
xor U14176 (N_14176,N_12585,N_12441);
nand U14177 (N_14177,N_12843,N_13080);
and U14178 (N_14178,N_12630,N_12381);
and U14179 (N_14179,N_12797,N_12706);
and U14180 (N_14180,N_12475,N_12051);
nor U14181 (N_14181,N_12753,N_12974);
and U14182 (N_14182,N_12318,N_12551);
nand U14183 (N_14183,N_13090,N_13052);
or U14184 (N_14184,N_12095,N_12915);
and U14185 (N_14185,N_12098,N_12670);
nor U14186 (N_14186,N_12370,N_12580);
xor U14187 (N_14187,N_12905,N_12387);
xnor U14188 (N_14188,N_12845,N_12696);
xor U14189 (N_14189,N_12470,N_12285);
and U14190 (N_14190,N_12119,N_13174);
nand U14191 (N_14191,N_13086,N_12701);
and U14192 (N_14192,N_12456,N_12676);
xor U14193 (N_14193,N_12634,N_12150);
nor U14194 (N_14194,N_13177,N_12936);
nand U14195 (N_14195,N_12349,N_12361);
nor U14196 (N_14196,N_13068,N_12750);
xor U14197 (N_14197,N_12567,N_12207);
nand U14198 (N_14198,N_12518,N_12993);
nand U14199 (N_14199,N_12168,N_12696);
or U14200 (N_14200,N_12308,N_13198);
or U14201 (N_14201,N_12341,N_12764);
nand U14202 (N_14202,N_12415,N_13045);
nor U14203 (N_14203,N_12199,N_12754);
and U14204 (N_14204,N_12217,N_13186);
or U14205 (N_14205,N_12565,N_12893);
xor U14206 (N_14206,N_12882,N_12968);
xnor U14207 (N_14207,N_12270,N_13110);
xor U14208 (N_14208,N_12273,N_13187);
or U14209 (N_14209,N_12306,N_12265);
nand U14210 (N_14210,N_13159,N_12650);
xor U14211 (N_14211,N_12548,N_12062);
nand U14212 (N_14212,N_12421,N_12048);
nand U14213 (N_14213,N_12930,N_12770);
nor U14214 (N_14214,N_12829,N_12635);
nor U14215 (N_14215,N_12863,N_13099);
and U14216 (N_14216,N_12114,N_12428);
nor U14217 (N_14217,N_12679,N_12407);
nand U14218 (N_14218,N_12722,N_12363);
and U14219 (N_14219,N_13021,N_12676);
nand U14220 (N_14220,N_12433,N_12370);
xnor U14221 (N_14221,N_12393,N_12999);
xor U14222 (N_14222,N_12391,N_12203);
or U14223 (N_14223,N_12396,N_12530);
nor U14224 (N_14224,N_13155,N_12552);
or U14225 (N_14225,N_13025,N_12948);
and U14226 (N_14226,N_13022,N_12158);
xor U14227 (N_14227,N_12159,N_13129);
and U14228 (N_14228,N_12019,N_12680);
and U14229 (N_14229,N_12630,N_12081);
or U14230 (N_14230,N_12906,N_12187);
nor U14231 (N_14231,N_12090,N_12341);
nand U14232 (N_14232,N_12136,N_12098);
nand U14233 (N_14233,N_12434,N_12307);
or U14234 (N_14234,N_13160,N_12891);
xor U14235 (N_14235,N_12392,N_12452);
and U14236 (N_14236,N_12250,N_12354);
nor U14237 (N_14237,N_12783,N_12901);
nand U14238 (N_14238,N_12161,N_12424);
nand U14239 (N_14239,N_12401,N_12305);
nand U14240 (N_14240,N_12168,N_12377);
xnor U14241 (N_14241,N_12336,N_12701);
and U14242 (N_14242,N_13124,N_12035);
nor U14243 (N_14243,N_12147,N_12237);
and U14244 (N_14244,N_13160,N_13128);
nor U14245 (N_14245,N_12801,N_12536);
and U14246 (N_14246,N_12265,N_12260);
nor U14247 (N_14247,N_13002,N_12785);
xnor U14248 (N_14248,N_12307,N_12139);
or U14249 (N_14249,N_12009,N_12860);
nor U14250 (N_14250,N_12202,N_12103);
nand U14251 (N_14251,N_12962,N_12589);
or U14252 (N_14252,N_12928,N_12192);
xor U14253 (N_14253,N_12518,N_12154);
nor U14254 (N_14254,N_12607,N_12981);
and U14255 (N_14255,N_12874,N_12169);
and U14256 (N_14256,N_13159,N_12409);
and U14257 (N_14257,N_12252,N_13017);
nand U14258 (N_14258,N_12013,N_12723);
xnor U14259 (N_14259,N_13066,N_13145);
and U14260 (N_14260,N_12885,N_12602);
or U14261 (N_14261,N_12930,N_12361);
and U14262 (N_14262,N_12538,N_12657);
xor U14263 (N_14263,N_13006,N_12810);
nand U14264 (N_14264,N_12840,N_12865);
xor U14265 (N_14265,N_13182,N_12017);
xor U14266 (N_14266,N_12758,N_13087);
xor U14267 (N_14267,N_12447,N_12561);
or U14268 (N_14268,N_12119,N_13063);
and U14269 (N_14269,N_12022,N_12373);
nand U14270 (N_14270,N_12920,N_12865);
and U14271 (N_14271,N_13051,N_12194);
nor U14272 (N_14272,N_12180,N_13153);
nor U14273 (N_14273,N_12602,N_12079);
nand U14274 (N_14274,N_12064,N_12327);
and U14275 (N_14275,N_13187,N_12625);
or U14276 (N_14276,N_13155,N_12880);
or U14277 (N_14277,N_12910,N_12297);
or U14278 (N_14278,N_12093,N_12928);
nand U14279 (N_14279,N_13199,N_12696);
nand U14280 (N_14280,N_12910,N_13131);
nand U14281 (N_14281,N_12711,N_12991);
xnor U14282 (N_14282,N_12457,N_12374);
xor U14283 (N_14283,N_12343,N_12847);
nor U14284 (N_14284,N_12888,N_12737);
or U14285 (N_14285,N_12828,N_12335);
and U14286 (N_14286,N_12277,N_13144);
nor U14287 (N_14287,N_12640,N_12853);
or U14288 (N_14288,N_12561,N_13165);
nand U14289 (N_14289,N_12073,N_12348);
xnor U14290 (N_14290,N_12398,N_12355);
nand U14291 (N_14291,N_12031,N_12082);
and U14292 (N_14292,N_12308,N_13190);
nand U14293 (N_14293,N_12364,N_12266);
xnor U14294 (N_14294,N_12982,N_12796);
nand U14295 (N_14295,N_12927,N_12300);
nand U14296 (N_14296,N_13106,N_12614);
or U14297 (N_14297,N_12097,N_12024);
and U14298 (N_14298,N_13109,N_13132);
and U14299 (N_14299,N_12221,N_12509);
nor U14300 (N_14300,N_12446,N_12120);
and U14301 (N_14301,N_12229,N_12730);
nand U14302 (N_14302,N_13074,N_12811);
and U14303 (N_14303,N_12386,N_12162);
nand U14304 (N_14304,N_12972,N_12865);
nor U14305 (N_14305,N_12587,N_12696);
nor U14306 (N_14306,N_12013,N_12326);
nand U14307 (N_14307,N_12045,N_12664);
xor U14308 (N_14308,N_12293,N_12870);
nor U14309 (N_14309,N_12858,N_12141);
or U14310 (N_14310,N_12626,N_12528);
nor U14311 (N_14311,N_12156,N_12594);
or U14312 (N_14312,N_12438,N_12533);
xnor U14313 (N_14313,N_13046,N_13086);
or U14314 (N_14314,N_12647,N_12872);
nor U14315 (N_14315,N_12808,N_13069);
nand U14316 (N_14316,N_12365,N_12223);
nor U14317 (N_14317,N_13006,N_12103);
and U14318 (N_14318,N_12040,N_13135);
nor U14319 (N_14319,N_13058,N_12140);
nor U14320 (N_14320,N_12979,N_12886);
nand U14321 (N_14321,N_12863,N_12199);
xnor U14322 (N_14322,N_12381,N_13073);
nor U14323 (N_14323,N_13046,N_12908);
xor U14324 (N_14324,N_12301,N_12334);
xnor U14325 (N_14325,N_12274,N_12683);
or U14326 (N_14326,N_12722,N_12846);
nand U14327 (N_14327,N_12757,N_12913);
and U14328 (N_14328,N_12639,N_12983);
nand U14329 (N_14329,N_12472,N_13140);
xnor U14330 (N_14330,N_12777,N_12587);
nor U14331 (N_14331,N_12475,N_13135);
or U14332 (N_14332,N_12782,N_13052);
and U14333 (N_14333,N_12230,N_12127);
xnor U14334 (N_14334,N_12981,N_12813);
nand U14335 (N_14335,N_13047,N_12881);
nand U14336 (N_14336,N_13029,N_12668);
xnor U14337 (N_14337,N_12201,N_12649);
or U14338 (N_14338,N_13016,N_13110);
xnor U14339 (N_14339,N_13078,N_13185);
nor U14340 (N_14340,N_12731,N_12318);
xnor U14341 (N_14341,N_13117,N_12812);
and U14342 (N_14342,N_13036,N_12262);
and U14343 (N_14343,N_12549,N_12091);
nor U14344 (N_14344,N_13185,N_13188);
nor U14345 (N_14345,N_12787,N_12102);
xnor U14346 (N_14346,N_12275,N_12918);
and U14347 (N_14347,N_12132,N_12075);
nor U14348 (N_14348,N_13102,N_12206);
and U14349 (N_14349,N_12497,N_12601);
nand U14350 (N_14350,N_12872,N_13177);
nor U14351 (N_14351,N_13090,N_12974);
nand U14352 (N_14352,N_12774,N_12297);
and U14353 (N_14353,N_12578,N_12175);
nor U14354 (N_14354,N_13147,N_12515);
or U14355 (N_14355,N_12712,N_12332);
nand U14356 (N_14356,N_13079,N_12007);
xnor U14357 (N_14357,N_13147,N_12653);
xor U14358 (N_14358,N_12056,N_12871);
nor U14359 (N_14359,N_12074,N_12603);
nand U14360 (N_14360,N_12660,N_12059);
xnor U14361 (N_14361,N_12465,N_12253);
or U14362 (N_14362,N_13197,N_12324);
and U14363 (N_14363,N_12804,N_12510);
nand U14364 (N_14364,N_12642,N_12958);
nand U14365 (N_14365,N_12502,N_12978);
and U14366 (N_14366,N_12489,N_12312);
nor U14367 (N_14367,N_12307,N_12517);
and U14368 (N_14368,N_12745,N_12104);
nand U14369 (N_14369,N_12167,N_12824);
and U14370 (N_14370,N_12600,N_12034);
nor U14371 (N_14371,N_13078,N_12572);
nor U14372 (N_14372,N_13030,N_13139);
nand U14373 (N_14373,N_12063,N_13007);
nand U14374 (N_14374,N_12226,N_12025);
and U14375 (N_14375,N_12299,N_12692);
nand U14376 (N_14376,N_12592,N_12862);
or U14377 (N_14377,N_12721,N_12309);
or U14378 (N_14378,N_12144,N_13004);
nor U14379 (N_14379,N_12399,N_12212);
nand U14380 (N_14380,N_12347,N_12746);
xnor U14381 (N_14381,N_12755,N_12548);
nand U14382 (N_14382,N_13088,N_12703);
nand U14383 (N_14383,N_12635,N_12426);
nand U14384 (N_14384,N_12599,N_12777);
nand U14385 (N_14385,N_13094,N_13004);
or U14386 (N_14386,N_12378,N_12671);
or U14387 (N_14387,N_12483,N_12539);
and U14388 (N_14388,N_12310,N_12053);
nand U14389 (N_14389,N_12241,N_12750);
nor U14390 (N_14390,N_13164,N_12082);
xnor U14391 (N_14391,N_12665,N_13041);
nand U14392 (N_14392,N_12132,N_13027);
and U14393 (N_14393,N_12902,N_13139);
and U14394 (N_14394,N_12032,N_12237);
nor U14395 (N_14395,N_12043,N_12852);
xnor U14396 (N_14396,N_12110,N_13186);
or U14397 (N_14397,N_12342,N_13140);
nand U14398 (N_14398,N_12870,N_12402);
and U14399 (N_14399,N_12371,N_12571);
nand U14400 (N_14400,N_13946,N_14244);
nand U14401 (N_14401,N_13875,N_13888);
nor U14402 (N_14402,N_13280,N_14075);
and U14403 (N_14403,N_13464,N_13955);
and U14404 (N_14404,N_13413,N_14373);
and U14405 (N_14405,N_14304,N_14045);
or U14406 (N_14406,N_14327,N_13659);
or U14407 (N_14407,N_13693,N_13795);
or U14408 (N_14408,N_13838,N_14203);
nand U14409 (N_14409,N_13764,N_13272);
nand U14410 (N_14410,N_13604,N_14156);
or U14411 (N_14411,N_13208,N_14054);
or U14412 (N_14412,N_13355,N_13590);
nor U14413 (N_14413,N_14112,N_14128);
or U14414 (N_14414,N_13293,N_13624);
and U14415 (N_14415,N_13341,N_13393);
or U14416 (N_14416,N_14052,N_13832);
nand U14417 (N_14417,N_13807,N_13645);
nor U14418 (N_14418,N_14238,N_13934);
and U14419 (N_14419,N_13559,N_14281);
and U14420 (N_14420,N_14387,N_13279);
xor U14421 (N_14421,N_14001,N_13502);
nor U14422 (N_14422,N_14019,N_13292);
nor U14423 (N_14423,N_14309,N_13840);
nand U14424 (N_14424,N_14114,N_13229);
and U14425 (N_14425,N_14258,N_13245);
and U14426 (N_14426,N_13906,N_14144);
or U14427 (N_14427,N_14395,N_13421);
xor U14428 (N_14428,N_13321,N_14053);
nor U14429 (N_14429,N_13535,N_13903);
nor U14430 (N_14430,N_13548,N_13568);
or U14431 (N_14431,N_13942,N_14357);
or U14432 (N_14432,N_13552,N_14242);
xor U14433 (N_14433,N_14367,N_13251);
and U14434 (N_14434,N_13597,N_13467);
xor U14435 (N_14435,N_13982,N_13486);
nor U14436 (N_14436,N_13753,N_13781);
nand U14437 (N_14437,N_13314,N_13687);
and U14438 (N_14438,N_14204,N_13473);
nor U14439 (N_14439,N_13556,N_14389);
and U14440 (N_14440,N_13519,N_14154);
nand U14441 (N_14441,N_14381,N_13423);
and U14442 (N_14442,N_13468,N_13709);
or U14443 (N_14443,N_14051,N_13299);
nor U14444 (N_14444,N_13787,N_14253);
and U14445 (N_14445,N_13793,N_13253);
or U14446 (N_14446,N_13534,N_13995);
nor U14447 (N_14447,N_13387,N_14352);
and U14448 (N_14448,N_13733,N_13352);
xnor U14449 (N_14449,N_13952,N_13738);
nand U14450 (N_14450,N_14050,N_13213);
or U14451 (N_14451,N_13480,N_14081);
nor U14452 (N_14452,N_13887,N_14089);
nand U14453 (N_14453,N_14251,N_13705);
or U14454 (N_14454,N_13349,N_13620);
xor U14455 (N_14455,N_13980,N_13586);
nand U14456 (N_14456,N_13471,N_14138);
nand U14457 (N_14457,N_14182,N_13858);
xnor U14458 (N_14458,N_13222,N_13905);
nand U14459 (N_14459,N_14032,N_13223);
nand U14460 (N_14460,N_14342,N_14007);
nor U14461 (N_14461,N_14266,N_14232);
xnor U14462 (N_14462,N_14091,N_14057);
and U14463 (N_14463,N_13895,N_13945);
xor U14464 (N_14464,N_14102,N_13667);
or U14465 (N_14465,N_13916,N_13706);
nand U14466 (N_14466,N_13907,N_13550);
or U14467 (N_14467,N_13288,N_14249);
or U14468 (N_14468,N_14212,N_14343);
or U14469 (N_14469,N_13329,N_14314);
or U14470 (N_14470,N_14196,N_13400);
nand U14471 (N_14471,N_13574,N_14298);
or U14472 (N_14472,N_14344,N_13405);
nor U14473 (N_14473,N_13318,N_13594);
nand U14474 (N_14474,N_13822,N_13201);
nor U14475 (N_14475,N_13869,N_13466);
nand U14476 (N_14476,N_13728,N_13827);
nor U14477 (N_14477,N_13252,N_13802);
xor U14478 (N_14478,N_13277,N_13569);
nand U14479 (N_14479,N_14390,N_14345);
or U14480 (N_14480,N_14276,N_13348);
and U14481 (N_14481,N_13500,N_14316);
xnor U14482 (N_14482,N_13211,N_13682);
nor U14483 (N_14483,N_13703,N_13830);
nor U14484 (N_14484,N_14312,N_13677);
nand U14485 (N_14485,N_13212,N_14347);
nand U14486 (N_14486,N_13224,N_13899);
nor U14487 (N_14487,N_13221,N_13570);
nor U14488 (N_14488,N_13607,N_13379);
nor U14489 (N_14489,N_13581,N_13459);
nor U14490 (N_14490,N_13704,N_14033);
or U14491 (N_14491,N_14093,N_13477);
nor U14492 (N_14492,N_13241,N_14169);
and U14493 (N_14493,N_14184,N_13302);
nor U14494 (N_14494,N_13300,N_14108);
and U14495 (N_14495,N_13449,N_13558);
or U14496 (N_14496,N_13600,N_13503);
or U14497 (N_14497,N_13488,N_13803);
and U14498 (N_14498,N_14025,N_13420);
xor U14499 (N_14499,N_13939,N_13725);
nand U14500 (N_14500,N_14132,N_14365);
xnor U14501 (N_14501,N_13937,N_13327);
nor U14502 (N_14502,N_13497,N_13894);
xor U14503 (N_14503,N_14077,N_14256);
nor U14504 (N_14504,N_14359,N_14239);
nand U14505 (N_14505,N_13542,N_13884);
nand U14506 (N_14506,N_13595,N_13819);
or U14507 (N_14507,N_14328,N_14146);
nand U14508 (N_14508,N_14267,N_13357);
nand U14509 (N_14509,N_13587,N_14178);
and U14510 (N_14510,N_13465,N_13317);
or U14511 (N_14511,N_14134,N_13755);
nand U14512 (N_14512,N_14264,N_14060);
and U14513 (N_14513,N_14125,N_14211);
and U14514 (N_14514,N_13472,N_14243);
or U14515 (N_14515,N_13271,N_13383);
xnor U14516 (N_14516,N_13306,N_13619);
nand U14517 (N_14517,N_13679,N_13825);
nand U14518 (N_14518,N_13561,N_13689);
and U14519 (N_14519,N_13790,N_14076);
and U14520 (N_14520,N_13384,N_13598);
xnor U14521 (N_14521,N_13707,N_14056);
and U14522 (N_14522,N_14164,N_13203);
or U14523 (N_14523,N_13653,N_14145);
xor U14524 (N_14524,N_13319,N_13397);
nor U14525 (N_14525,N_14029,N_14369);
or U14526 (N_14526,N_14319,N_13417);
and U14527 (N_14527,N_13258,N_14067);
and U14528 (N_14528,N_13774,N_13289);
and U14529 (N_14529,N_13647,N_13975);
or U14530 (N_14530,N_13315,N_13510);
nor U14531 (N_14531,N_13575,N_13901);
or U14532 (N_14532,N_14109,N_14168);
nand U14533 (N_14533,N_14170,N_14284);
and U14534 (N_14534,N_13640,N_13893);
nor U14535 (N_14535,N_14307,N_13308);
xor U14536 (N_14536,N_13275,N_13915);
or U14537 (N_14537,N_13770,N_13386);
and U14538 (N_14538,N_14136,N_14326);
nor U14539 (N_14539,N_13862,N_13381);
and U14540 (N_14540,N_13720,N_14382);
nor U14541 (N_14541,N_14008,N_13785);
or U14542 (N_14542,N_13515,N_13226);
nor U14543 (N_14543,N_14254,N_14252);
xor U14544 (N_14544,N_13833,N_14188);
xnor U14545 (N_14545,N_13429,N_14355);
or U14546 (N_14546,N_13750,N_13248);
nand U14547 (N_14547,N_13892,N_13380);
or U14548 (N_14548,N_14014,N_14377);
and U14549 (N_14549,N_13518,N_14257);
nor U14550 (N_14550,N_13873,N_13509);
nand U14551 (N_14551,N_13260,N_13451);
xnor U14552 (N_14552,N_13920,N_13722);
and U14553 (N_14553,N_13846,N_13741);
nor U14554 (N_14554,N_13369,N_13262);
xor U14555 (N_14555,N_13428,N_14227);
nand U14556 (N_14556,N_13419,N_13991);
and U14557 (N_14557,N_13462,N_13435);
nor U14558 (N_14558,N_14368,N_14152);
or U14559 (N_14559,N_14293,N_13736);
nand U14560 (N_14560,N_13220,N_13402);
xnor U14561 (N_14561,N_13266,N_13917);
nor U14562 (N_14562,N_14159,N_13636);
nor U14563 (N_14563,N_13896,N_13291);
or U14564 (N_14564,N_13748,N_14118);
nand U14565 (N_14565,N_14065,N_13931);
nand U14566 (N_14566,N_14058,N_13941);
xnor U14567 (N_14567,N_13611,N_13506);
xor U14568 (N_14568,N_13929,N_13806);
or U14569 (N_14569,N_14362,N_14062);
or U14570 (N_14570,N_14351,N_14139);
nand U14571 (N_14571,N_14332,N_13344);
nand U14572 (N_14572,N_13713,N_13727);
or U14573 (N_14573,N_13305,N_13239);
nor U14574 (N_14574,N_13623,N_13997);
nand U14575 (N_14575,N_14048,N_13734);
xnor U14576 (N_14576,N_13463,N_14094);
nand U14577 (N_14577,N_14215,N_14107);
or U14578 (N_14578,N_13921,N_13244);
and U14579 (N_14579,N_13246,N_13336);
and U14580 (N_14580,N_14099,N_13286);
nand U14581 (N_14581,N_14375,N_13643);
and U14582 (N_14582,N_14000,N_13673);
nor U14583 (N_14583,N_13670,N_13879);
or U14584 (N_14584,N_13566,N_14018);
and U14585 (N_14585,N_13525,N_13565);
nand U14586 (N_14586,N_14277,N_13439);
nor U14587 (N_14587,N_14294,N_13563);
nor U14588 (N_14588,N_13539,N_14040);
nand U14589 (N_14589,N_14106,N_13998);
nor U14590 (N_14590,N_13523,N_13885);
nor U14591 (N_14591,N_14208,N_14163);
or U14592 (N_14592,N_13639,N_13808);
or U14593 (N_14593,N_13256,N_13661);
or U14594 (N_14594,N_14031,N_14236);
or U14595 (N_14595,N_13278,N_14217);
xor U14596 (N_14596,N_13641,N_14071);
and U14597 (N_14597,N_13886,N_13541);
nand U14598 (N_14598,N_13814,N_13270);
or U14599 (N_14599,N_13672,N_13746);
nor U14600 (N_14600,N_14183,N_14246);
nor U14601 (N_14601,N_13767,N_13837);
nor U14602 (N_14602,N_14397,N_13865);
nand U14603 (N_14603,N_13403,N_13834);
nand U14604 (N_14604,N_13237,N_13512);
nand U14605 (N_14605,N_14041,N_14262);
and U14606 (N_14606,N_13216,N_13742);
and U14607 (N_14607,N_14047,N_14289);
and U14608 (N_14608,N_14228,N_13621);
nand U14609 (N_14609,N_13589,N_13333);
and U14610 (N_14610,N_13441,N_14147);
nor U14611 (N_14611,N_13322,N_13392);
xnor U14612 (N_14612,N_14366,N_13889);
xnor U14613 (N_14613,N_14015,N_14119);
xnor U14614 (N_14614,N_14069,N_13257);
and U14615 (N_14615,N_13789,N_14350);
and U14616 (N_14616,N_13655,N_13684);
nand U14617 (N_14617,N_14263,N_14330);
and U14618 (N_14618,N_13416,N_13868);
nand U14619 (N_14619,N_14167,N_14206);
nor U14620 (N_14620,N_13973,N_13508);
and U14621 (N_14621,N_13854,N_14165);
or U14622 (N_14622,N_13494,N_13591);
and U14623 (N_14623,N_13797,N_13533);
and U14624 (N_14624,N_13493,N_13880);
or U14625 (N_14625,N_13576,N_13855);
nor U14626 (N_14626,N_13301,N_13996);
or U14627 (N_14627,N_13207,N_14068);
xor U14628 (N_14628,N_13674,N_14175);
or U14629 (N_14629,N_13474,N_14292);
nand U14630 (N_14630,N_13630,N_13455);
or U14631 (N_14631,N_13671,N_13882);
nand U14632 (N_14632,N_14162,N_14197);
xor U14633 (N_14633,N_13702,N_14078);
nor U14634 (N_14634,N_13231,N_14143);
and U14635 (N_14635,N_14255,N_13695);
nor U14636 (N_14636,N_14198,N_13678);
xor U14637 (N_14637,N_13631,N_13475);
and U14638 (N_14638,N_13981,N_13448);
and U14639 (N_14639,N_14348,N_14038);
xor U14640 (N_14640,N_13759,N_13482);
or U14641 (N_14641,N_14288,N_14149);
nand U14642 (N_14642,N_13635,N_14354);
nand U14643 (N_14643,N_13902,N_13370);
xnor U14644 (N_14644,N_14226,N_14221);
nand U14645 (N_14645,N_14049,N_13577);
or U14646 (N_14646,N_14009,N_14231);
and U14647 (N_14647,N_13596,N_13382);
or U14648 (N_14648,N_13373,N_13994);
nor U14649 (N_14649,N_13544,N_13891);
or U14650 (N_14650,N_14092,N_14210);
nand U14651 (N_14651,N_14209,N_13656);
and U14652 (N_14652,N_13504,N_13514);
nand U14653 (N_14653,N_13965,N_13356);
xor U14654 (N_14654,N_14334,N_13276);
or U14655 (N_14655,N_13867,N_14336);
or U14656 (N_14656,N_13815,N_14115);
xor U14657 (N_14657,N_13911,N_13928);
nor U14658 (N_14658,N_14340,N_14237);
or U14659 (N_14659,N_13737,N_13217);
xor U14660 (N_14660,N_13951,N_14063);
or U14661 (N_14661,N_14085,N_13948);
or U14662 (N_14662,N_13681,N_14179);
nor U14663 (N_14663,N_14082,N_14270);
xnor U14664 (N_14664,N_14339,N_13985);
xnor U14665 (N_14665,N_13747,N_13940);
xor U14666 (N_14666,N_13859,N_13442);
nor U14667 (N_14667,N_14323,N_14005);
or U14668 (N_14668,N_13430,N_13849);
xor U14669 (N_14669,N_13233,N_13227);
and U14670 (N_14670,N_13206,N_13718);
xor U14671 (N_14671,N_13626,N_13404);
xor U14672 (N_14672,N_13492,N_13599);
and U14673 (N_14673,N_13912,N_13376);
and U14674 (N_14674,N_13805,N_14337);
or U14675 (N_14675,N_13527,N_13778);
xnor U14676 (N_14676,N_13218,N_14137);
and U14677 (N_14677,N_13295,N_14021);
and U14678 (N_14678,N_13555,N_14220);
xnor U14679 (N_14679,N_14308,N_14287);
nand U14680 (N_14680,N_13287,N_14177);
nand U14681 (N_14681,N_13378,N_13751);
nor U14682 (N_14682,N_13409,N_13766);
nand U14683 (N_14683,N_14153,N_13414);
nor U14684 (N_14684,N_13338,N_13826);
and U14685 (N_14685,N_14315,N_13371);
or U14686 (N_14686,N_14110,N_13777);
and U14687 (N_14687,N_14043,N_13490);
nand U14688 (N_14688,N_14207,N_13823);
and U14689 (N_14689,N_13769,N_13377);
xor U14690 (N_14690,N_13567,N_13717);
or U14691 (N_14691,N_13922,N_14121);
nand U14692 (N_14692,N_14130,N_13324);
and U14693 (N_14693,N_14361,N_13660);
and U14694 (N_14694,N_13507,N_14393);
or U14695 (N_14695,N_14202,N_13622);
nor U14696 (N_14696,N_14234,N_13909);
nand U14697 (N_14697,N_13969,N_14356);
nor U14698 (N_14698,N_13668,N_13365);
nand U14699 (N_14699,N_13296,N_13394);
or U14700 (N_14700,N_14218,N_13489);
nor U14701 (N_14701,N_14186,N_13938);
nand U14702 (N_14702,N_13263,N_13968);
nand U14703 (N_14703,N_13685,N_14034);
nand U14704 (N_14704,N_13723,N_13697);
xor U14705 (N_14705,N_13584,N_14370);
or U14706 (N_14706,N_13634,N_13786);
nor U14707 (N_14707,N_13583,N_13219);
nor U14708 (N_14708,N_13585,N_14012);
xnor U14709 (N_14709,N_13491,N_14072);
nor U14710 (N_14710,N_13234,N_13729);
nor U14711 (N_14711,N_13648,N_13551);
and U14712 (N_14712,N_13431,N_14300);
and U14713 (N_14713,N_13553,N_14098);
xnor U14714 (N_14714,N_13652,N_13651);
nor U14715 (N_14715,N_13664,N_13731);
or U14716 (N_14716,N_14297,N_13761);
nor U14717 (N_14717,N_14385,N_13358);
nand U14718 (N_14718,N_13714,N_13844);
and U14719 (N_14719,N_13970,N_13927);
xnor U14720 (N_14720,N_13616,N_13877);
and U14721 (N_14721,N_14245,N_14321);
or U14722 (N_14722,N_13269,N_13974);
or U14723 (N_14723,N_13521,N_13335);
or U14724 (N_14724,N_13399,N_14148);
nor U14725 (N_14725,N_13783,N_13863);
and U14726 (N_14726,N_13845,N_13547);
xnor U14727 (N_14727,N_13801,N_14299);
and U14728 (N_14728,N_14229,N_14037);
nand U14729 (N_14729,N_13476,N_14274);
and U14730 (N_14730,N_14087,N_13976);
nand U14731 (N_14731,N_13943,N_13285);
nand U14732 (N_14732,N_13540,N_14122);
nor U14733 (N_14733,N_13817,N_13613);
xor U14734 (N_14734,N_13243,N_14301);
nor U14735 (N_14735,N_13505,N_13726);
nor U14736 (N_14736,N_13366,N_13963);
or U14737 (N_14737,N_13593,N_13791);
nor U14738 (N_14738,N_14383,N_13739);
nand U14739 (N_14739,N_13949,N_14392);
nand U14740 (N_14740,N_14247,N_13560);
nand U14741 (N_14741,N_14026,N_13874);
nand U14742 (N_14742,N_13900,N_13440);
or U14743 (N_14743,N_13332,N_13388);
and U14744 (N_14744,N_13654,N_14088);
nand U14745 (N_14745,N_14261,N_13799);
nand U14746 (N_14746,N_14338,N_13612);
xnor U14747 (N_14747,N_13487,N_14142);
and U14748 (N_14748,N_14158,N_13989);
nor U14749 (N_14749,N_14320,N_13961);
or U14750 (N_14750,N_14272,N_13610);
or U14751 (N_14751,N_13484,N_13375);
nand U14752 (N_14752,N_13721,N_13368);
or U14753 (N_14753,N_13690,N_13944);
nor U14754 (N_14754,N_14317,N_13724);
and U14755 (N_14755,N_14113,N_13294);
nand U14756 (N_14756,N_13242,N_13427);
nand U14757 (N_14757,N_13663,N_14398);
nor U14758 (N_14758,N_14311,N_14331);
xor U14759 (N_14759,N_14013,N_14023);
or U14760 (N_14760,N_13537,N_13627);
and U14761 (N_14761,N_14278,N_13436);
xnor U14762 (N_14762,N_14187,N_14035);
nor U14763 (N_14763,N_14296,N_13214);
xor U14764 (N_14764,N_14101,N_13228);
nand U14765 (N_14765,N_14379,N_13346);
nand U14766 (N_14766,N_14039,N_13529);
and U14767 (N_14767,N_14283,N_13546);
xor U14768 (N_14768,N_14279,N_13323);
xor U14769 (N_14769,N_13520,N_13628);
or U14770 (N_14770,N_14141,N_13433);
xor U14771 (N_14771,N_13821,N_14268);
nor U14772 (N_14772,N_13408,N_14290);
or U14773 (N_14773,N_14027,N_14083);
nand U14774 (N_14774,N_14305,N_14192);
xor U14775 (N_14775,N_13342,N_13345);
nor U14776 (N_14776,N_13572,N_13878);
xor U14777 (N_14777,N_14002,N_13772);
and U14778 (N_14778,N_13259,N_13385);
nor U14779 (N_14779,N_14322,N_13364);
or U14780 (N_14780,N_13719,N_13637);
nand U14781 (N_14781,N_13710,N_14084);
and U14782 (N_14782,N_13735,N_13831);
or U14783 (N_14783,N_14346,N_13872);
xnor U14784 (N_14784,N_13812,N_13744);
nor U14785 (N_14785,N_13918,N_13617);
nand U14786 (N_14786,N_13924,N_13526);
nand U14787 (N_14787,N_13914,N_13443);
nor U14788 (N_14788,N_13304,N_13543);
nand U14789 (N_14789,N_13760,N_13794);
or U14790 (N_14790,N_14064,N_13910);
nor U14791 (N_14791,N_13530,N_13957);
xnor U14792 (N_14792,N_13438,N_13829);
nand U14793 (N_14793,N_13632,N_13501);
or U14794 (N_14794,N_14394,N_14017);
nor U14795 (N_14795,N_13273,N_13255);
nor U14796 (N_14796,N_13646,N_14195);
or U14797 (N_14797,N_13676,N_13768);
and U14798 (N_14798,N_14095,N_14117);
or U14799 (N_14799,N_13926,N_13424);
nor U14800 (N_14800,N_13485,N_14171);
nor U14801 (N_14801,N_13715,N_13771);
nand U14802 (N_14802,N_13665,N_14028);
xor U14803 (N_14803,N_14044,N_14105);
xnor U14804 (N_14804,N_14124,N_14024);
nand U14805 (N_14805,N_13391,N_14275);
or U14806 (N_14806,N_14127,N_14191);
xnor U14807 (N_14807,N_14310,N_13788);
or U14808 (N_14808,N_14172,N_13372);
and U14809 (N_14809,N_13412,N_13864);
and U14810 (N_14810,N_13784,N_14116);
and U14811 (N_14811,N_14399,N_14273);
or U14812 (N_14812,N_13337,N_14269);
xor U14813 (N_14813,N_14241,N_14248);
nand U14814 (N_14814,N_14120,N_13856);
or U14815 (N_14815,N_13692,N_13340);
xor U14816 (N_14816,N_13549,N_13396);
and U14817 (N_14817,N_13460,N_13669);
xor U14818 (N_14818,N_13694,N_13904);
xor U14819 (N_14819,N_13749,N_13511);
nor U14820 (N_14820,N_14066,N_13204);
or U14821 (N_14821,N_14123,N_13881);
or U14822 (N_14822,N_13608,N_13809);
or U14823 (N_14823,N_14129,N_14235);
or U14824 (N_14824,N_13516,N_13268);
nor U14825 (N_14825,N_13479,N_13615);
xor U14826 (N_14826,N_13618,N_13307);
or U14827 (N_14827,N_13601,N_14333);
xor U14828 (N_14828,N_14055,N_14073);
or U14829 (N_14829,N_13528,N_14157);
nor U14830 (N_14830,N_13842,N_14189);
or U14831 (N_14831,N_13432,N_13461);
nand U14832 (N_14832,N_14022,N_13913);
and U14833 (N_14833,N_13406,N_13389);
nand U14834 (N_14834,N_14216,N_14036);
and U14835 (N_14835,N_14160,N_13758);
xnor U14836 (N_14836,N_14097,N_13848);
nand U14837 (N_14837,N_13732,N_13495);
xor U14838 (N_14838,N_13499,N_14225);
nor U14839 (N_14839,N_13326,N_13363);
and U14840 (N_14840,N_13582,N_13283);
nand U14841 (N_14841,N_13452,N_13716);
nor U14842 (N_14842,N_13650,N_14004);
xnor U14843 (N_14843,N_13320,N_13792);
and U14844 (N_14844,N_14030,N_13267);
nand U14845 (N_14845,N_13513,N_13447);
or U14846 (N_14846,N_13847,N_13629);
nor U14847 (N_14847,N_14286,N_14161);
nor U14848 (N_14848,N_13853,N_13813);
or U14849 (N_14849,N_13290,N_13496);
nand U14850 (N_14850,N_13554,N_14271);
nor U14851 (N_14851,N_13779,N_13979);
xnor U14852 (N_14852,N_14302,N_13454);
or U14853 (N_14853,N_14010,N_14230);
or U14854 (N_14854,N_14003,N_13861);
nor U14855 (N_14855,N_13765,N_13798);
nor U14856 (N_14856,N_13850,N_14059);
or U14857 (N_14857,N_14046,N_14341);
nand U14858 (N_14858,N_14303,N_13686);
and U14859 (N_14859,N_13966,N_13298);
xor U14860 (N_14860,N_13411,N_13249);
and U14861 (N_14861,N_13757,N_13395);
xnor U14862 (N_14862,N_13457,N_13254);
or U14863 (N_14863,N_13312,N_13579);
xnor U14864 (N_14864,N_13274,N_13932);
xor U14865 (N_14865,N_14386,N_13410);
xnor U14866 (N_14866,N_14233,N_13811);
or U14867 (N_14867,N_13469,N_13841);
nor U14868 (N_14868,N_14155,N_13401);
and U14869 (N_14869,N_14166,N_14213);
xnor U14870 (N_14870,N_13418,N_13633);
nand U14871 (N_14871,N_14131,N_13870);
nand U14872 (N_14872,N_14086,N_14200);
xnor U14873 (N_14873,N_13964,N_14016);
nor U14874 (N_14874,N_13350,N_13782);
nand U14875 (N_14875,N_13481,N_14020);
and U14876 (N_14876,N_13522,N_14363);
nand U14877 (N_14877,N_13284,N_13680);
nor U14878 (N_14878,N_14080,N_13936);
nor U14879 (N_14879,N_13960,N_13343);
or U14880 (N_14880,N_13557,N_13580);
and U14881 (N_14881,N_14384,N_13588);
nor U14882 (N_14882,N_14173,N_13517);
xnor U14883 (N_14883,N_14176,N_13483);
nor U14884 (N_14884,N_14193,N_14295);
xnor U14885 (N_14885,N_13662,N_13609);
nand U14886 (N_14886,N_14259,N_14126);
xor U14887 (N_14887,N_13232,N_13642);
and U14888 (N_14888,N_13578,N_13605);
or U14889 (N_14889,N_13824,N_13238);
xnor U14890 (N_14890,N_14388,N_14201);
and U14891 (N_14891,N_13983,N_13247);
and U14892 (N_14892,N_13564,N_13776);
nand U14893 (N_14893,N_13407,N_13353);
and U14894 (N_14894,N_13754,N_14103);
xnor U14895 (N_14895,N_14151,N_13531);
or U14896 (N_14896,N_14180,N_13839);
or U14897 (N_14897,N_13860,N_13209);
or U14898 (N_14898,N_13956,N_13740);
nor U14899 (N_14899,N_13458,N_13804);
xnor U14900 (N_14900,N_13422,N_13993);
xnor U14901 (N_14901,N_13250,N_13532);
nand U14902 (N_14902,N_13359,N_14096);
or U14903 (N_14903,N_13282,N_13752);
xnor U14904 (N_14904,N_14325,N_13264);
nand U14905 (N_14905,N_13675,N_13959);
xor U14906 (N_14906,N_13743,N_13658);
or U14907 (N_14907,N_14396,N_13971);
or U14908 (N_14908,N_13967,N_14011);
and U14909 (N_14909,N_14260,N_14135);
or U14910 (N_14910,N_13202,N_13836);
nor U14911 (N_14911,N_13351,N_13745);
and U14912 (N_14912,N_13325,N_14358);
nor U14913 (N_14913,N_13657,N_13843);
nor U14914 (N_14914,N_13919,N_13456);
xor U14915 (N_14915,N_13711,N_13309);
nand U14916 (N_14916,N_13696,N_14223);
nand U14917 (N_14917,N_13361,N_14349);
nand U14918 (N_14918,N_13871,N_13898);
nor U14919 (N_14919,N_13450,N_13281);
nand U14920 (N_14920,N_14219,N_13478);
nor U14921 (N_14921,N_14104,N_13688);
or U14922 (N_14922,N_13992,N_14282);
xnor U14923 (N_14923,N_13691,N_13857);
or U14924 (N_14924,N_14214,N_13763);
nand U14925 (N_14925,N_13987,N_14199);
nor U14926 (N_14926,N_13331,N_13923);
nor U14927 (N_14927,N_13573,N_14090);
and U14928 (N_14928,N_13390,N_14194);
nand U14929 (N_14929,N_13313,N_13374);
and U14930 (N_14930,N_13930,N_14391);
xnor U14931 (N_14931,N_14374,N_13818);
nand U14932 (N_14932,N_13775,N_13666);
xnor U14933 (N_14933,N_13470,N_14079);
xnor U14934 (N_14934,N_13592,N_14291);
nand U14935 (N_14935,N_14285,N_14376);
and U14936 (N_14936,N_14372,N_13773);
or U14937 (N_14937,N_13614,N_14240);
and U14938 (N_14938,N_13712,N_14042);
and U14939 (N_14939,N_13852,N_13230);
nor U14940 (N_14940,N_13240,N_14265);
and U14941 (N_14941,N_13756,N_13730);
nand U14942 (N_14942,N_13235,N_13303);
and U14943 (N_14943,N_13215,N_14335);
nand U14944 (N_14944,N_14324,N_13972);
nor U14945 (N_14945,N_13780,N_13297);
nand U14946 (N_14946,N_13810,N_14250);
xor U14947 (N_14947,N_14006,N_13354);
or U14948 (N_14948,N_13708,N_14140);
xor U14949 (N_14949,N_13950,N_14380);
or U14950 (N_14950,N_14074,N_14111);
or U14951 (N_14951,N_13360,N_14306);
or U14952 (N_14952,N_13571,N_13434);
and U14953 (N_14953,N_13954,N_14190);
nand U14954 (N_14954,N_13426,N_13538);
nand U14955 (N_14955,N_14313,N_14070);
and U14956 (N_14956,N_13265,N_14364);
nand U14957 (N_14957,N_13334,N_13545);
or U14958 (N_14958,N_14222,N_13990);
nand U14959 (N_14959,N_13205,N_13683);
or U14960 (N_14960,N_13947,N_13953);
xnor U14961 (N_14961,N_13236,N_13316);
nor U14962 (N_14962,N_14318,N_13644);
or U14963 (N_14963,N_13890,N_13828);
and U14964 (N_14964,N_14185,N_13524);
nand U14965 (N_14965,N_13445,N_13958);
nand U14966 (N_14966,N_13649,N_13762);
xor U14967 (N_14967,N_14360,N_13698);
and U14968 (N_14968,N_13700,N_14329);
or U14969 (N_14969,N_13339,N_13328);
and U14970 (N_14970,N_13453,N_13796);
nand U14971 (N_14971,N_13978,N_13415);
nand U14972 (N_14972,N_13602,N_13925);
nand U14973 (N_14973,N_13225,N_13851);
or U14974 (N_14974,N_13367,N_13444);
nor U14975 (N_14975,N_13437,N_14378);
nor U14976 (N_14976,N_13835,N_13816);
nand U14977 (N_14977,N_14181,N_13800);
and U14978 (N_14978,N_13701,N_13962);
nand U14979 (N_14979,N_13200,N_13603);
or U14980 (N_14980,N_13933,N_14371);
or U14981 (N_14981,N_14174,N_13398);
nand U14982 (N_14982,N_13935,N_14224);
nand U14983 (N_14983,N_13425,N_13562);
nand U14984 (N_14984,N_14100,N_13977);
and U14985 (N_14985,N_13820,N_14353);
and U14986 (N_14986,N_13261,N_13984);
and U14987 (N_14987,N_13625,N_13908);
nor U14988 (N_14988,N_13311,N_13606);
and U14989 (N_14989,N_13876,N_13883);
nand U14990 (N_14990,N_13347,N_13986);
or U14991 (N_14991,N_13362,N_14205);
nand U14992 (N_14992,N_14061,N_13536);
xnor U14993 (N_14993,N_14150,N_13330);
and U14994 (N_14994,N_13999,N_13897);
xor U14995 (N_14995,N_13210,N_13638);
nor U14996 (N_14996,N_13866,N_13988);
xnor U14997 (N_14997,N_13310,N_13446);
xnor U14998 (N_14998,N_14280,N_13498);
nand U14999 (N_14999,N_13699,N_14133);
or U15000 (N_15000,N_13226,N_13529);
and U15001 (N_15001,N_13706,N_14321);
or U15002 (N_15002,N_13400,N_13500);
xor U15003 (N_15003,N_13814,N_13691);
and U15004 (N_15004,N_13220,N_13548);
and U15005 (N_15005,N_14268,N_14328);
xnor U15006 (N_15006,N_13868,N_14379);
nand U15007 (N_15007,N_13995,N_13611);
nor U15008 (N_15008,N_14371,N_14226);
nor U15009 (N_15009,N_13649,N_14123);
nor U15010 (N_15010,N_14040,N_13901);
xnor U15011 (N_15011,N_13455,N_13315);
xnor U15012 (N_15012,N_14047,N_13303);
and U15013 (N_15013,N_13829,N_13306);
and U15014 (N_15014,N_13259,N_14378);
and U15015 (N_15015,N_14184,N_13478);
nor U15016 (N_15016,N_14350,N_14202);
or U15017 (N_15017,N_14083,N_14118);
xor U15018 (N_15018,N_13374,N_13822);
nor U15019 (N_15019,N_14176,N_13991);
and U15020 (N_15020,N_14053,N_14213);
and U15021 (N_15021,N_14142,N_13565);
or U15022 (N_15022,N_13844,N_13759);
and U15023 (N_15023,N_14284,N_13847);
xor U15024 (N_15024,N_14147,N_13602);
xor U15025 (N_15025,N_13811,N_13893);
or U15026 (N_15026,N_13552,N_13997);
nand U15027 (N_15027,N_13800,N_14156);
xor U15028 (N_15028,N_14319,N_13599);
nand U15029 (N_15029,N_13773,N_13937);
nor U15030 (N_15030,N_14309,N_14295);
or U15031 (N_15031,N_14153,N_14363);
or U15032 (N_15032,N_13423,N_13827);
xor U15033 (N_15033,N_13375,N_13784);
nand U15034 (N_15034,N_14136,N_14116);
and U15035 (N_15035,N_13683,N_13719);
nor U15036 (N_15036,N_13494,N_13767);
xnor U15037 (N_15037,N_13685,N_14135);
or U15038 (N_15038,N_13994,N_13885);
and U15039 (N_15039,N_14075,N_13330);
xnor U15040 (N_15040,N_14097,N_14363);
xor U15041 (N_15041,N_13990,N_13651);
nand U15042 (N_15042,N_14382,N_14218);
or U15043 (N_15043,N_13231,N_14002);
xor U15044 (N_15044,N_13250,N_13702);
or U15045 (N_15045,N_13796,N_13501);
nor U15046 (N_15046,N_14014,N_14239);
nand U15047 (N_15047,N_13588,N_13291);
and U15048 (N_15048,N_14372,N_13800);
nor U15049 (N_15049,N_13502,N_13509);
nor U15050 (N_15050,N_14143,N_14328);
xor U15051 (N_15051,N_13755,N_13851);
nand U15052 (N_15052,N_13992,N_13823);
nand U15053 (N_15053,N_13528,N_13996);
nor U15054 (N_15054,N_13942,N_13317);
xor U15055 (N_15055,N_13936,N_14163);
and U15056 (N_15056,N_14381,N_14181);
nand U15057 (N_15057,N_13769,N_13821);
nand U15058 (N_15058,N_13247,N_13939);
and U15059 (N_15059,N_13256,N_13272);
xor U15060 (N_15060,N_14198,N_13659);
and U15061 (N_15061,N_14375,N_14090);
nand U15062 (N_15062,N_13463,N_13709);
nor U15063 (N_15063,N_13572,N_13257);
nand U15064 (N_15064,N_14343,N_13664);
and U15065 (N_15065,N_13990,N_13742);
nor U15066 (N_15066,N_14321,N_14282);
and U15067 (N_15067,N_14348,N_13902);
or U15068 (N_15068,N_13376,N_13360);
or U15069 (N_15069,N_13605,N_13304);
and U15070 (N_15070,N_13850,N_14351);
and U15071 (N_15071,N_14326,N_13808);
or U15072 (N_15072,N_13998,N_13633);
and U15073 (N_15073,N_13603,N_14106);
nand U15074 (N_15074,N_13876,N_13223);
nand U15075 (N_15075,N_14224,N_14180);
nor U15076 (N_15076,N_13876,N_13727);
nor U15077 (N_15077,N_13406,N_14376);
nor U15078 (N_15078,N_13288,N_13200);
xnor U15079 (N_15079,N_13480,N_13451);
xnor U15080 (N_15080,N_13349,N_13721);
nand U15081 (N_15081,N_13544,N_13578);
nor U15082 (N_15082,N_13273,N_13752);
and U15083 (N_15083,N_13554,N_13617);
nand U15084 (N_15084,N_13728,N_13752);
nand U15085 (N_15085,N_13388,N_13515);
nand U15086 (N_15086,N_14068,N_13792);
xnor U15087 (N_15087,N_13454,N_13674);
nand U15088 (N_15088,N_13807,N_14181);
or U15089 (N_15089,N_13508,N_13637);
nand U15090 (N_15090,N_13828,N_13449);
nor U15091 (N_15091,N_13469,N_14380);
xor U15092 (N_15092,N_13460,N_13650);
nor U15093 (N_15093,N_13979,N_13215);
and U15094 (N_15094,N_13752,N_14234);
and U15095 (N_15095,N_13691,N_13884);
or U15096 (N_15096,N_13500,N_13636);
and U15097 (N_15097,N_13964,N_13843);
nand U15098 (N_15098,N_13544,N_13535);
and U15099 (N_15099,N_13751,N_13920);
and U15100 (N_15100,N_13975,N_13995);
nand U15101 (N_15101,N_13982,N_14332);
nand U15102 (N_15102,N_13856,N_14370);
or U15103 (N_15103,N_13399,N_13734);
and U15104 (N_15104,N_13297,N_14077);
and U15105 (N_15105,N_13332,N_13712);
or U15106 (N_15106,N_13268,N_13513);
nand U15107 (N_15107,N_13361,N_14363);
nor U15108 (N_15108,N_13697,N_13715);
and U15109 (N_15109,N_14372,N_13553);
xnor U15110 (N_15110,N_14154,N_13878);
xnor U15111 (N_15111,N_13298,N_13799);
nand U15112 (N_15112,N_13539,N_13771);
nand U15113 (N_15113,N_14352,N_14102);
nand U15114 (N_15114,N_13487,N_14238);
xor U15115 (N_15115,N_13529,N_14190);
nor U15116 (N_15116,N_13787,N_13838);
or U15117 (N_15117,N_14155,N_13966);
and U15118 (N_15118,N_13539,N_13892);
xnor U15119 (N_15119,N_14058,N_13336);
xor U15120 (N_15120,N_13765,N_13852);
nand U15121 (N_15121,N_13582,N_14390);
nand U15122 (N_15122,N_13641,N_13394);
xor U15123 (N_15123,N_14115,N_13721);
xnor U15124 (N_15124,N_14286,N_13690);
xnor U15125 (N_15125,N_13212,N_13685);
nor U15126 (N_15126,N_13308,N_13567);
nor U15127 (N_15127,N_13372,N_14091);
nand U15128 (N_15128,N_14333,N_14245);
or U15129 (N_15129,N_13660,N_14008);
and U15130 (N_15130,N_13690,N_13226);
xor U15131 (N_15131,N_14169,N_13932);
or U15132 (N_15132,N_14090,N_13254);
or U15133 (N_15133,N_13700,N_13806);
xor U15134 (N_15134,N_13531,N_13429);
and U15135 (N_15135,N_13315,N_13344);
xor U15136 (N_15136,N_13625,N_13564);
nand U15137 (N_15137,N_13591,N_13781);
or U15138 (N_15138,N_14112,N_13423);
nor U15139 (N_15139,N_13217,N_14079);
xnor U15140 (N_15140,N_13625,N_13877);
xor U15141 (N_15141,N_13428,N_13385);
nor U15142 (N_15142,N_13326,N_14349);
or U15143 (N_15143,N_13636,N_13810);
or U15144 (N_15144,N_13620,N_13200);
or U15145 (N_15145,N_13823,N_14072);
nor U15146 (N_15146,N_14372,N_13814);
and U15147 (N_15147,N_13294,N_13556);
and U15148 (N_15148,N_14390,N_13929);
and U15149 (N_15149,N_14160,N_14066);
nor U15150 (N_15150,N_13474,N_13525);
and U15151 (N_15151,N_13714,N_13832);
or U15152 (N_15152,N_14086,N_14103);
xnor U15153 (N_15153,N_13964,N_13687);
xnor U15154 (N_15154,N_13906,N_13998);
nand U15155 (N_15155,N_13281,N_13276);
and U15156 (N_15156,N_13516,N_13207);
nor U15157 (N_15157,N_13262,N_13700);
nand U15158 (N_15158,N_13671,N_14193);
nor U15159 (N_15159,N_13500,N_14267);
xnor U15160 (N_15160,N_14311,N_13907);
nand U15161 (N_15161,N_14124,N_13841);
or U15162 (N_15162,N_13277,N_13671);
nand U15163 (N_15163,N_13721,N_13660);
xor U15164 (N_15164,N_13366,N_13924);
and U15165 (N_15165,N_14097,N_13538);
xor U15166 (N_15166,N_14381,N_14326);
and U15167 (N_15167,N_13250,N_13522);
or U15168 (N_15168,N_13741,N_14145);
xnor U15169 (N_15169,N_13397,N_13676);
nor U15170 (N_15170,N_14326,N_13399);
xnor U15171 (N_15171,N_14187,N_13290);
nand U15172 (N_15172,N_14348,N_13374);
nand U15173 (N_15173,N_13759,N_13870);
and U15174 (N_15174,N_13242,N_13876);
xor U15175 (N_15175,N_13223,N_13348);
and U15176 (N_15176,N_13262,N_13417);
or U15177 (N_15177,N_13520,N_13537);
and U15178 (N_15178,N_13398,N_13247);
nand U15179 (N_15179,N_14350,N_13773);
xnor U15180 (N_15180,N_14135,N_13312);
or U15181 (N_15181,N_13375,N_14068);
nand U15182 (N_15182,N_13651,N_13692);
nand U15183 (N_15183,N_14030,N_13509);
nor U15184 (N_15184,N_13208,N_13280);
nor U15185 (N_15185,N_13353,N_14395);
nor U15186 (N_15186,N_13301,N_13984);
xnor U15187 (N_15187,N_13833,N_14266);
xor U15188 (N_15188,N_13900,N_13976);
nand U15189 (N_15189,N_14208,N_14331);
nor U15190 (N_15190,N_13827,N_13816);
and U15191 (N_15191,N_13505,N_14316);
xnor U15192 (N_15192,N_13599,N_13538);
and U15193 (N_15193,N_14146,N_13542);
nand U15194 (N_15194,N_13864,N_13392);
nand U15195 (N_15195,N_13464,N_13200);
nand U15196 (N_15196,N_13295,N_13868);
nor U15197 (N_15197,N_13619,N_13706);
nand U15198 (N_15198,N_13655,N_14319);
and U15199 (N_15199,N_13909,N_14107);
xor U15200 (N_15200,N_13330,N_14155);
nand U15201 (N_15201,N_13896,N_13925);
nand U15202 (N_15202,N_14175,N_13469);
xor U15203 (N_15203,N_13883,N_13679);
or U15204 (N_15204,N_13237,N_14211);
xnor U15205 (N_15205,N_13568,N_13398);
nand U15206 (N_15206,N_14219,N_13497);
and U15207 (N_15207,N_14332,N_13451);
nor U15208 (N_15208,N_13372,N_13963);
and U15209 (N_15209,N_13292,N_14190);
and U15210 (N_15210,N_13240,N_13512);
nand U15211 (N_15211,N_13581,N_13314);
or U15212 (N_15212,N_13859,N_13269);
xnor U15213 (N_15213,N_14179,N_14139);
xor U15214 (N_15214,N_14092,N_13857);
and U15215 (N_15215,N_13375,N_13534);
xor U15216 (N_15216,N_14075,N_13694);
xnor U15217 (N_15217,N_14326,N_14146);
nor U15218 (N_15218,N_14301,N_13265);
or U15219 (N_15219,N_13224,N_13852);
nand U15220 (N_15220,N_13548,N_14084);
xnor U15221 (N_15221,N_13917,N_13761);
xor U15222 (N_15222,N_13589,N_13532);
and U15223 (N_15223,N_14291,N_13990);
or U15224 (N_15224,N_13310,N_13580);
nor U15225 (N_15225,N_13483,N_13452);
xnor U15226 (N_15226,N_13747,N_14227);
and U15227 (N_15227,N_13225,N_13417);
nand U15228 (N_15228,N_14182,N_14356);
nor U15229 (N_15229,N_14379,N_13226);
or U15230 (N_15230,N_13235,N_14344);
and U15231 (N_15231,N_13854,N_14188);
or U15232 (N_15232,N_13357,N_14321);
or U15233 (N_15233,N_13890,N_14055);
nand U15234 (N_15234,N_13677,N_14191);
nand U15235 (N_15235,N_13757,N_13740);
xor U15236 (N_15236,N_13594,N_13454);
xor U15237 (N_15237,N_14357,N_14107);
nor U15238 (N_15238,N_14000,N_14342);
xnor U15239 (N_15239,N_13900,N_14241);
and U15240 (N_15240,N_13270,N_14174);
or U15241 (N_15241,N_14113,N_13808);
nand U15242 (N_15242,N_13281,N_14222);
nor U15243 (N_15243,N_13910,N_14261);
nor U15244 (N_15244,N_14231,N_13561);
or U15245 (N_15245,N_13771,N_14288);
xor U15246 (N_15246,N_13733,N_14137);
and U15247 (N_15247,N_13528,N_14091);
and U15248 (N_15248,N_13324,N_14240);
nand U15249 (N_15249,N_13226,N_13686);
or U15250 (N_15250,N_13964,N_14121);
xor U15251 (N_15251,N_14138,N_13625);
or U15252 (N_15252,N_13475,N_13252);
nand U15253 (N_15253,N_14079,N_13214);
or U15254 (N_15254,N_13507,N_13735);
xor U15255 (N_15255,N_13401,N_13531);
or U15256 (N_15256,N_13823,N_14117);
and U15257 (N_15257,N_13742,N_13741);
nand U15258 (N_15258,N_13242,N_13222);
nand U15259 (N_15259,N_13308,N_14047);
and U15260 (N_15260,N_13799,N_13450);
nor U15261 (N_15261,N_13418,N_14004);
and U15262 (N_15262,N_14316,N_14129);
xnor U15263 (N_15263,N_13265,N_14127);
nand U15264 (N_15264,N_14095,N_14340);
xnor U15265 (N_15265,N_14178,N_13259);
xor U15266 (N_15266,N_13767,N_13954);
and U15267 (N_15267,N_14251,N_13373);
or U15268 (N_15268,N_14175,N_13273);
and U15269 (N_15269,N_13624,N_13549);
or U15270 (N_15270,N_14281,N_14237);
or U15271 (N_15271,N_14199,N_13837);
nand U15272 (N_15272,N_13968,N_14334);
or U15273 (N_15273,N_14363,N_13203);
and U15274 (N_15274,N_13568,N_13207);
or U15275 (N_15275,N_14103,N_13881);
nand U15276 (N_15276,N_13616,N_14003);
xor U15277 (N_15277,N_13864,N_14373);
nand U15278 (N_15278,N_13544,N_13824);
or U15279 (N_15279,N_13416,N_14187);
or U15280 (N_15280,N_14304,N_13445);
and U15281 (N_15281,N_13893,N_13310);
xnor U15282 (N_15282,N_14110,N_13406);
or U15283 (N_15283,N_13815,N_13942);
or U15284 (N_15284,N_13459,N_13582);
and U15285 (N_15285,N_13490,N_13202);
or U15286 (N_15286,N_14154,N_13574);
nor U15287 (N_15287,N_14108,N_13490);
nand U15288 (N_15288,N_13643,N_13780);
xnor U15289 (N_15289,N_13426,N_14205);
and U15290 (N_15290,N_14265,N_13925);
and U15291 (N_15291,N_13966,N_13326);
xor U15292 (N_15292,N_13383,N_13288);
nor U15293 (N_15293,N_14330,N_13243);
xor U15294 (N_15294,N_14269,N_13232);
or U15295 (N_15295,N_13699,N_13329);
xor U15296 (N_15296,N_14322,N_14135);
nor U15297 (N_15297,N_14310,N_13828);
nor U15298 (N_15298,N_13633,N_13829);
or U15299 (N_15299,N_13535,N_13395);
nand U15300 (N_15300,N_14070,N_13465);
or U15301 (N_15301,N_13499,N_13518);
nor U15302 (N_15302,N_13242,N_13482);
nor U15303 (N_15303,N_13880,N_13591);
or U15304 (N_15304,N_13472,N_13457);
nand U15305 (N_15305,N_14261,N_13602);
xor U15306 (N_15306,N_13464,N_13336);
or U15307 (N_15307,N_13262,N_13430);
nand U15308 (N_15308,N_13371,N_13326);
or U15309 (N_15309,N_13707,N_13623);
or U15310 (N_15310,N_13403,N_14095);
nand U15311 (N_15311,N_13881,N_13316);
or U15312 (N_15312,N_13789,N_13903);
xor U15313 (N_15313,N_13698,N_13444);
nor U15314 (N_15314,N_13783,N_13486);
nor U15315 (N_15315,N_13967,N_14331);
or U15316 (N_15316,N_13483,N_14369);
xnor U15317 (N_15317,N_14037,N_14291);
or U15318 (N_15318,N_13979,N_13924);
nor U15319 (N_15319,N_13280,N_13249);
or U15320 (N_15320,N_14278,N_13455);
or U15321 (N_15321,N_13454,N_14100);
xnor U15322 (N_15322,N_13468,N_14347);
or U15323 (N_15323,N_14268,N_14136);
nor U15324 (N_15324,N_13353,N_13791);
xnor U15325 (N_15325,N_13676,N_13470);
nor U15326 (N_15326,N_13254,N_13249);
nand U15327 (N_15327,N_13646,N_13506);
xor U15328 (N_15328,N_13793,N_13901);
xor U15329 (N_15329,N_14227,N_13515);
nand U15330 (N_15330,N_13368,N_13728);
nor U15331 (N_15331,N_13807,N_14281);
xnor U15332 (N_15332,N_14175,N_13832);
xnor U15333 (N_15333,N_13874,N_13245);
or U15334 (N_15334,N_13490,N_14194);
and U15335 (N_15335,N_13984,N_13643);
nand U15336 (N_15336,N_14142,N_14076);
xor U15337 (N_15337,N_13662,N_13377);
or U15338 (N_15338,N_14224,N_13335);
nor U15339 (N_15339,N_13277,N_13565);
nand U15340 (N_15340,N_13710,N_13902);
nand U15341 (N_15341,N_14192,N_13587);
nor U15342 (N_15342,N_13746,N_13442);
and U15343 (N_15343,N_13314,N_13507);
and U15344 (N_15344,N_13694,N_13555);
and U15345 (N_15345,N_13290,N_13352);
nand U15346 (N_15346,N_14024,N_13321);
nor U15347 (N_15347,N_13501,N_13898);
nand U15348 (N_15348,N_14081,N_13974);
nor U15349 (N_15349,N_13826,N_14014);
nand U15350 (N_15350,N_13765,N_14326);
and U15351 (N_15351,N_13683,N_14018);
nor U15352 (N_15352,N_14332,N_13729);
and U15353 (N_15353,N_13855,N_13200);
and U15354 (N_15354,N_13516,N_13360);
or U15355 (N_15355,N_13267,N_13399);
nor U15356 (N_15356,N_13511,N_13329);
nand U15357 (N_15357,N_13635,N_14207);
xor U15358 (N_15358,N_13335,N_13696);
nand U15359 (N_15359,N_13336,N_13890);
and U15360 (N_15360,N_13864,N_13950);
xnor U15361 (N_15361,N_14031,N_14337);
nor U15362 (N_15362,N_14211,N_14078);
nor U15363 (N_15363,N_14318,N_13473);
xnor U15364 (N_15364,N_14228,N_13587);
and U15365 (N_15365,N_13638,N_13797);
nor U15366 (N_15366,N_13304,N_13918);
or U15367 (N_15367,N_13426,N_14166);
xor U15368 (N_15368,N_14168,N_14336);
nor U15369 (N_15369,N_13467,N_13203);
xnor U15370 (N_15370,N_13866,N_13422);
and U15371 (N_15371,N_14140,N_13940);
nand U15372 (N_15372,N_13729,N_14310);
xnor U15373 (N_15373,N_13992,N_14265);
or U15374 (N_15374,N_14111,N_13924);
xnor U15375 (N_15375,N_13674,N_13503);
or U15376 (N_15376,N_14185,N_13337);
nor U15377 (N_15377,N_14365,N_13853);
nor U15378 (N_15378,N_14191,N_13368);
nor U15379 (N_15379,N_14169,N_13714);
or U15380 (N_15380,N_14245,N_13914);
and U15381 (N_15381,N_13226,N_13398);
and U15382 (N_15382,N_14120,N_13201);
nor U15383 (N_15383,N_13962,N_13623);
nor U15384 (N_15384,N_13985,N_13520);
and U15385 (N_15385,N_13500,N_14296);
and U15386 (N_15386,N_13531,N_13595);
and U15387 (N_15387,N_13707,N_13636);
and U15388 (N_15388,N_13395,N_13903);
nor U15389 (N_15389,N_14300,N_14376);
nand U15390 (N_15390,N_13724,N_13938);
nand U15391 (N_15391,N_13818,N_13977);
and U15392 (N_15392,N_13657,N_13461);
or U15393 (N_15393,N_14305,N_13621);
or U15394 (N_15394,N_14022,N_13814);
nor U15395 (N_15395,N_13499,N_13983);
nor U15396 (N_15396,N_13925,N_13480);
nand U15397 (N_15397,N_13594,N_13239);
nand U15398 (N_15398,N_13269,N_13217);
and U15399 (N_15399,N_14230,N_13401);
or U15400 (N_15400,N_13456,N_14128);
nor U15401 (N_15401,N_13367,N_13845);
xnor U15402 (N_15402,N_14038,N_13793);
and U15403 (N_15403,N_13910,N_13414);
nor U15404 (N_15404,N_13805,N_14085);
xnor U15405 (N_15405,N_13977,N_13674);
nor U15406 (N_15406,N_13764,N_13973);
xor U15407 (N_15407,N_14298,N_13745);
xor U15408 (N_15408,N_13722,N_13813);
xnor U15409 (N_15409,N_13961,N_13570);
nand U15410 (N_15410,N_14215,N_14100);
or U15411 (N_15411,N_14327,N_13966);
or U15412 (N_15412,N_13576,N_13940);
and U15413 (N_15413,N_14375,N_14001);
or U15414 (N_15414,N_14362,N_13545);
or U15415 (N_15415,N_14031,N_14280);
nor U15416 (N_15416,N_13804,N_13557);
or U15417 (N_15417,N_13973,N_14180);
nor U15418 (N_15418,N_13620,N_13420);
xor U15419 (N_15419,N_13654,N_13692);
xor U15420 (N_15420,N_13591,N_13496);
xor U15421 (N_15421,N_14120,N_13503);
nor U15422 (N_15422,N_14300,N_14081);
or U15423 (N_15423,N_13359,N_13337);
xor U15424 (N_15424,N_14109,N_13846);
or U15425 (N_15425,N_13722,N_13670);
and U15426 (N_15426,N_13561,N_14313);
and U15427 (N_15427,N_13257,N_14118);
nor U15428 (N_15428,N_13481,N_14114);
nand U15429 (N_15429,N_13497,N_14117);
or U15430 (N_15430,N_13424,N_14375);
and U15431 (N_15431,N_13607,N_13394);
nor U15432 (N_15432,N_14285,N_13364);
nor U15433 (N_15433,N_13761,N_13875);
or U15434 (N_15434,N_13852,N_14003);
or U15435 (N_15435,N_13938,N_13497);
nand U15436 (N_15436,N_14312,N_14316);
nand U15437 (N_15437,N_14280,N_14032);
or U15438 (N_15438,N_13314,N_14187);
nand U15439 (N_15439,N_14398,N_14066);
nor U15440 (N_15440,N_14385,N_14163);
and U15441 (N_15441,N_14319,N_14221);
or U15442 (N_15442,N_13453,N_13897);
or U15443 (N_15443,N_13629,N_13526);
xnor U15444 (N_15444,N_14108,N_13871);
nand U15445 (N_15445,N_13892,N_13846);
or U15446 (N_15446,N_13808,N_13857);
nor U15447 (N_15447,N_14197,N_13600);
and U15448 (N_15448,N_14091,N_13788);
xor U15449 (N_15449,N_14006,N_13812);
nand U15450 (N_15450,N_13617,N_13956);
or U15451 (N_15451,N_13255,N_14348);
or U15452 (N_15452,N_14206,N_13658);
or U15453 (N_15453,N_14332,N_14156);
or U15454 (N_15454,N_13897,N_14151);
xnor U15455 (N_15455,N_13994,N_13608);
and U15456 (N_15456,N_13394,N_14067);
or U15457 (N_15457,N_14289,N_14315);
nand U15458 (N_15458,N_13666,N_13448);
nor U15459 (N_15459,N_13742,N_13488);
nor U15460 (N_15460,N_13438,N_13668);
and U15461 (N_15461,N_14398,N_13215);
xnor U15462 (N_15462,N_14200,N_14373);
and U15463 (N_15463,N_13535,N_13922);
and U15464 (N_15464,N_13926,N_13287);
nor U15465 (N_15465,N_13713,N_14172);
nand U15466 (N_15466,N_13226,N_13415);
xor U15467 (N_15467,N_13231,N_13744);
xnor U15468 (N_15468,N_13790,N_14364);
nand U15469 (N_15469,N_13354,N_13942);
nor U15470 (N_15470,N_13998,N_13454);
and U15471 (N_15471,N_13548,N_13697);
nand U15472 (N_15472,N_14160,N_13900);
nor U15473 (N_15473,N_13360,N_13397);
nor U15474 (N_15474,N_14121,N_14194);
nor U15475 (N_15475,N_13841,N_13969);
nor U15476 (N_15476,N_13889,N_13877);
and U15477 (N_15477,N_14011,N_13919);
nand U15478 (N_15478,N_13757,N_13726);
xnor U15479 (N_15479,N_13381,N_13321);
xnor U15480 (N_15480,N_14197,N_13493);
xor U15481 (N_15481,N_14191,N_13933);
nand U15482 (N_15482,N_14336,N_14398);
nand U15483 (N_15483,N_14201,N_13632);
nand U15484 (N_15484,N_14232,N_13933);
or U15485 (N_15485,N_14264,N_14224);
nor U15486 (N_15486,N_13250,N_13958);
nand U15487 (N_15487,N_14019,N_13563);
xnor U15488 (N_15488,N_13418,N_13897);
xor U15489 (N_15489,N_13383,N_14370);
xor U15490 (N_15490,N_14307,N_14229);
nor U15491 (N_15491,N_13698,N_13962);
xor U15492 (N_15492,N_14239,N_13891);
and U15493 (N_15493,N_13853,N_14027);
xnor U15494 (N_15494,N_13418,N_13645);
or U15495 (N_15495,N_13588,N_14190);
nor U15496 (N_15496,N_13630,N_14066);
and U15497 (N_15497,N_13770,N_14006);
xor U15498 (N_15498,N_14147,N_13752);
or U15499 (N_15499,N_14384,N_14377);
and U15500 (N_15500,N_13490,N_13246);
and U15501 (N_15501,N_13904,N_13423);
and U15502 (N_15502,N_14217,N_14032);
or U15503 (N_15503,N_14347,N_13280);
nand U15504 (N_15504,N_13443,N_13271);
and U15505 (N_15505,N_14396,N_13625);
and U15506 (N_15506,N_13889,N_13281);
and U15507 (N_15507,N_14268,N_13913);
xor U15508 (N_15508,N_13355,N_14243);
or U15509 (N_15509,N_14269,N_14078);
nor U15510 (N_15510,N_14361,N_13956);
nand U15511 (N_15511,N_14102,N_13218);
xnor U15512 (N_15512,N_14295,N_14334);
nand U15513 (N_15513,N_13628,N_13673);
nand U15514 (N_15514,N_14005,N_13291);
xnor U15515 (N_15515,N_14321,N_13742);
nand U15516 (N_15516,N_14192,N_13803);
nand U15517 (N_15517,N_13981,N_13918);
and U15518 (N_15518,N_13331,N_13745);
nor U15519 (N_15519,N_14105,N_13945);
xnor U15520 (N_15520,N_14067,N_13604);
and U15521 (N_15521,N_14014,N_14223);
nor U15522 (N_15522,N_13200,N_13954);
nand U15523 (N_15523,N_14216,N_13468);
or U15524 (N_15524,N_14361,N_13594);
or U15525 (N_15525,N_14094,N_13962);
nor U15526 (N_15526,N_13240,N_13392);
nand U15527 (N_15527,N_13229,N_14278);
xor U15528 (N_15528,N_14162,N_13275);
nand U15529 (N_15529,N_14210,N_13956);
or U15530 (N_15530,N_14227,N_14099);
xor U15531 (N_15531,N_13328,N_13482);
nor U15532 (N_15532,N_14333,N_13407);
xor U15533 (N_15533,N_14304,N_13971);
and U15534 (N_15534,N_13881,N_13956);
and U15535 (N_15535,N_13751,N_13668);
nand U15536 (N_15536,N_14094,N_14102);
or U15537 (N_15537,N_13400,N_13816);
and U15538 (N_15538,N_14365,N_13254);
nor U15539 (N_15539,N_13488,N_13466);
xor U15540 (N_15540,N_13843,N_13954);
nand U15541 (N_15541,N_13984,N_13612);
or U15542 (N_15542,N_14281,N_14151);
nor U15543 (N_15543,N_14198,N_14108);
and U15544 (N_15544,N_14166,N_13678);
xor U15545 (N_15545,N_14081,N_14289);
nand U15546 (N_15546,N_13545,N_14118);
xnor U15547 (N_15547,N_13990,N_13714);
or U15548 (N_15548,N_13517,N_13337);
nand U15549 (N_15549,N_13258,N_13530);
nand U15550 (N_15550,N_13954,N_13408);
or U15551 (N_15551,N_13801,N_14341);
xor U15552 (N_15552,N_14045,N_13462);
or U15553 (N_15553,N_13745,N_14047);
and U15554 (N_15554,N_13261,N_13726);
and U15555 (N_15555,N_13773,N_13594);
xnor U15556 (N_15556,N_13476,N_14266);
or U15557 (N_15557,N_14295,N_14202);
nor U15558 (N_15558,N_13320,N_13348);
and U15559 (N_15559,N_13761,N_13869);
nand U15560 (N_15560,N_13486,N_13235);
nor U15561 (N_15561,N_14214,N_13667);
and U15562 (N_15562,N_13780,N_13745);
and U15563 (N_15563,N_13612,N_14341);
nor U15564 (N_15564,N_14305,N_13970);
nor U15565 (N_15565,N_14188,N_13939);
or U15566 (N_15566,N_13339,N_13717);
xnor U15567 (N_15567,N_14197,N_13693);
xor U15568 (N_15568,N_13315,N_14087);
and U15569 (N_15569,N_13639,N_13671);
or U15570 (N_15570,N_13616,N_13621);
and U15571 (N_15571,N_13362,N_14227);
xnor U15572 (N_15572,N_14029,N_13833);
nand U15573 (N_15573,N_14179,N_13651);
and U15574 (N_15574,N_14367,N_13696);
xnor U15575 (N_15575,N_13963,N_14235);
nand U15576 (N_15576,N_14365,N_13403);
or U15577 (N_15577,N_14273,N_13674);
or U15578 (N_15578,N_14325,N_13457);
or U15579 (N_15579,N_13669,N_13658);
nand U15580 (N_15580,N_13704,N_13749);
nand U15581 (N_15581,N_14038,N_13677);
or U15582 (N_15582,N_13668,N_13270);
nor U15583 (N_15583,N_14226,N_13363);
xor U15584 (N_15584,N_13654,N_13388);
nor U15585 (N_15585,N_14150,N_13894);
or U15586 (N_15586,N_14285,N_14030);
xnor U15587 (N_15587,N_14222,N_14335);
nor U15588 (N_15588,N_14090,N_14106);
xnor U15589 (N_15589,N_14083,N_13329);
or U15590 (N_15590,N_13848,N_13412);
xnor U15591 (N_15591,N_14154,N_13738);
nand U15592 (N_15592,N_13259,N_13616);
nor U15593 (N_15593,N_14100,N_13930);
and U15594 (N_15594,N_13640,N_14385);
nor U15595 (N_15595,N_13992,N_14064);
nor U15596 (N_15596,N_14380,N_13530);
xor U15597 (N_15597,N_13267,N_13647);
and U15598 (N_15598,N_13346,N_13577);
nand U15599 (N_15599,N_13804,N_14275);
xnor U15600 (N_15600,N_14554,N_14960);
nand U15601 (N_15601,N_15398,N_14463);
and U15602 (N_15602,N_14908,N_15538);
nand U15603 (N_15603,N_14706,N_14905);
xor U15604 (N_15604,N_15566,N_14431);
nand U15605 (N_15605,N_15010,N_14473);
and U15606 (N_15606,N_14883,N_15114);
nand U15607 (N_15607,N_15453,N_15514);
xnor U15608 (N_15608,N_15599,N_15009);
nor U15609 (N_15609,N_14612,N_15157);
xor U15610 (N_15610,N_15493,N_15390);
or U15611 (N_15611,N_15097,N_15221);
xnor U15612 (N_15612,N_14848,N_15048);
nor U15613 (N_15613,N_14722,N_15203);
xor U15614 (N_15614,N_14646,N_15594);
and U15615 (N_15615,N_14520,N_14618);
nor U15616 (N_15616,N_15196,N_14629);
xnor U15617 (N_15617,N_15422,N_15581);
and U15618 (N_15618,N_14928,N_15050);
nor U15619 (N_15619,N_14776,N_14506);
nor U15620 (N_15620,N_15132,N_15045);
or U15621 (N_15621,N_14593,N_15273);
nand U15622 (N_15622,N_15477,N_15076);
or U15623 (N_15623,N_15144,N_15558);
nand U15624 (N_15624,N_15393,N_15253);
nand U15625 (N_15625,N_14620,N_14790);
or U15626 (N_15626,N_15201,N_15420);
or U15627 (N_15627,N_14862,N_14433);
xnor U15628 (N_15628,N_15371,N_15384);
nor U15629 (N_15629,N_15129,N_14560);
nor U15630 (N_15630,N_15254,N_15309);
nor U15631 (N_15631,N_14673,N_15532);
nand U15632 (N_15632,N_15434,N_15507);
and U15633 (N_15633,N_14505,N_14992);
or U15634 (N_15634,N_14421,N_14887);
nand U15635 (N_15635,N_15155,N_15184);
or U15636 (N_15636,N_15524,N_15106);
xor U15637 (N_15637,N_14746,N_14546);
xor U15638 (N_15638,N_14884,N_14654);
xnor U15639 (N_15639,N_14532,N_14570);
xnor U15640 (N_15640,N_14951,N_15510);
nand U15641 (N_15641,N_15481,N_14780);
or U15642 (N_15642,N_14692,N_15505);
and U15643 (N_15643,N_15211,N_15570);
or U15644 (N_15644,N_15437,N_15412);
and U15645 (N_15645,N_15576,N_15466);
nor U15646 (N_15646,N_14541,N_14796);
or U15647 (N_15647,N_15128,N_15082);
or U15648 (N_15648,N_15270,N_14828);
and U15649 (N_15649,N_15386,N_15419);
nand U15650 (N_15650,N_15153,N_14902);
xor U15651 (N_15651,N_14488,N_14669);
xor U15652 (N_15652,N_14551,N_14571);
xor U15653 (N_15653,N_15158,N_15498);
or U15654 (N_15654,N_14415,N_15376);
and U15655 (N_15655,N_15069,N_14925);
nor U15656 (N_15656,N_14765,N_15455);
xor U15657 (N_15657,N_15164,N_15206);
and U15658 (N_15658,N_15468,N_14726);
nor U15659 (N_15659,N_15587,N_14753);
and U15660 (N_15660,N_15573,N_14601);
nor U15661 (N_15661,N_14875,N_14708);
nor U15662 (N_15662,N_15344,N_15315);
nor U15663 (N_15663,N_14589,N_15336);
and U15664 (N_15664,N_14536,N_15145);
nand U15665 (N_15665,N_14988,N_15277);
xnor U15666 (N_15666,N_15127,N_14579);
xnor U15667 (N_15667,N_14482,N_15290);
nand U15668 (N_15668,N_15259,N_15428);
and U15669 (N_15669,N_15197,N_15240);
nand U15670 (N_15670,N_14958,N_15559);
nand U15671 (N_15671,N_14975,N_15204);
xnor U15672 (N_15672,N_14794,N_14610);
and U15673 (N_15673,N_14762,N_15202);
and U15674 (N_15674,N_14870,N_15301);
nand U15675 (N_15675,N_14854,N_14721);
and U15676 (N_15676,N_14631,N_14922);
and U15677 (N_15677,N_14662,N_15054);
and U15678 (N_15678,N_14542,N_15289);
or U15679 (N_15679,N_14868,N_14619);
nand U15680 (N_15680,N_14758,N_15073);
and U15681 (N_15681,N_14627,N_15094);
and U15682 (N_15682,N_14643,N_15355);
or U15683 (N_15683,N_14731,N_15295);
xnor U15684 (N_15684,N_14413,N_15503);
or U15685 (N_15685,N_15396,N_15552);
or U15686 (N_15686,N_15354,N_15190);
or U15687 (N_15687,N_14760,N_15572);
nor U15688 (N_15688,N_15228,N_14537);
or U15689 (N_15689,N_14750,N_15193);
or U15690 (N_15690,N_14489,N_14691);
nand U15691 (N_15691,N_15349,N_15238);
and U15692 (N_15692,N_15329,N_14432);
or U15693 (N_15693,N_15018,N_14989);
or U15694 (N_15694,N_14914,N_14947);
or U15695 (N_15695,N_14526,N_14448);
nor U15696 (N_15696,N_14769,N_15230);
and U15697 (N_15697,N_14650,N_15124);
and U15698 (N_15698,N_14476,N_15011);
and U15699 (N_15699,N_15095,N_14671);
xor U15700 (N_15700,N_15316,N_14604);
xor U15701 (N_15701,N_14569,N_15084);
nor U15702 (N_15702,N_15154,N_14451);
or U15703 (N_15703,N_15087,N_14584);
nor U15704 (N_15704,N_15348,N_14998);
nor U15705 (N_15705,N_14982,N_15590);
nor U15706 (N_15706,N_14971,N_14785);
or U15707 (N_15707,N_15163,N_15125);
or U15708 (N_15708,N_14996,N_15431);
nand U15709 (N_15709,N_15026,N_14934);
and U15710 (N_15710,N_14458,N_15509);
and U15711 (N_15711,N_15310,N_14402);
and U15712 (N_15712,N_14830,N_14430);
xor U15713 (N_15713,N_14952,N_14889);
and U15714 (N_15714,N_14798,N_15225);
xnor U15715 (N_15715,N_15183,N_15533);
nor U15716 (N_15716,N_14876,N_15502);
xnor U15717 (N_15717,N_15229,N_15460);
nand U15718 (N_15718,N_15022,N_14895);
xnor U15719 (N_15719,N_15584,N_14841);
nor U15720 (N_15720,N_14857,N_15194);
xor U15721 (N_15721,N_15529,N_15372);
and U15722 (N_15722,N_14441,N_14446);
nor U15723 (N_15723,N_14937,N_14549);
or U15724 (N_15724,N_14616,N_15334);
xor U15725 (N_15725,N_14575,N_15023);
nand U15726 (N_15726,N_15318,N_14617);
nor U15727 (N_15727,N_14797,N_14578);
and U15728 (N_15728,N_15062,N_14930);
or U15729 (N_15729,N_15521,N_15282);
nand U15730 (N_15730,N_15494,N_14401);
nor U15731 (N_15731,N_14877,N_14698);
and U15732 (N_15732,N_14553,N_14603);
xnor U15733 (N_15733,N_15130,N_15464);
and U15734 (N_15734,N_15089,N_14519);
or U15735 (N_15735,N_15473,N_14525);
nor U15736 (N_15736,N_14995,N_14703);
nand U15737 (N_15737,N_15199,N_15262);
nand U15738 (N_15738,N_15359,N_14932);
nor U15739 (N_15739,N_15569,N_14545);
nor U15740 (N_15740,N_15265,N_14592);
and U15741 (N_15741,N_14510,N_14831);
nand U15742 (N_15742,N_14814,N_15066);
xnor U15743 (N_15743,N_15088,N_15450);
xor U15744 (N_15744,N_15403,N_15239);
xnor U15745 (N_15745,N_14727,N_15563);
xor U15746 (N_15746,N_14832,N_14948);
or U15747 (N_15747,N_15519,N_15245);
and U15748 (N_15748,N_14602,N_14943);
nand U15749 (N_15749,N_14422,N_15352);
or U15750 (N_15750,N_14550,N_14836);
or U15751 (N_15751,N_15070,N_14909);
nor U15752 (N_15752,N_14994,N_15139);
and U15753 (N_15753,N_14968,N_14405);
nand U15754 (N_15754,N_15171,N_14504);
xnor U15755 (N_15755,N_14702,N_15243);
nand U15756 (N_15756,N_14880,N_14480);
and U15757 (N_15757,N_15444,N_15058);
nand U15758 (N_15758,N_15074,N_15340);
xor U15759 (N_15759,N_15525,N_15374);
xor U15760 (N_15760,N_15233,N_14719);
nor U15761 (N_15761,N_14900,N_15452);
xnor U15762 (N_15762,N_14795,N_14573);
or U15763 (N_15763,N_14462,N_15491);
nor U15764 (N_15764,N_15476,N_15469);
xor U15765 (N_15765,N_15006,N_14660);
xor U15766 (N_15766,N_14508,N_15261);
nand U15767 (N_15767,N_14490,N_14632);
and U15768 (N_15768,N_15005,N_14756);
or U15769 (N_15769,N_14655,N_15085);
xor U15770 (N_15770,N_14978,N_15571);
nand U15771 (N_15771,N_14891,N_15195);
nand U15772 (N_15772,N_15350,N_15322);
xnor U15773 (N_15773,N_14853,N_15513);
nand U15774 (N_15774,N_14899,N_14675);
xor U15775 (N_15775,N_14443,N_15160);
nor U15776 (N_15776,N_14511,N_15362);
xnor U15777 (N_15777,N_14543,N_14723);
or U15778 (N_15778,N_14946,N_15442);
xor U15779 (N_15779,N_14621,N_14626);
nor U15780 (N_15780,N_15380,N_15086);
nor U15781 (N_15781,N_15459,N_15330);
nor U15782 (N_15782,N_15119,N_15165);
or U15783 (N_15783,N_15326,N_14921);
and U15784 (N_15784,N_14640,N_14893);
nand U15785 (N_15785,N_14533,N_14582);
or U15786 (N_15786,N_14624,N_14426);
nor U15787 (N_15787,N_14827,N_14897);
xor U15788 (N_15788,N_15304,N_15418);
nor U15789 (N_15789,N_14858,N_15036);
and U15790 (N_15790,N_14474,N_15294);
and U15791 (N_15791,N_15044,N_15592);
xnor U15792 (N_15792,N_15324,N_15472);
nor U15793 (N_15793,N_15223,N_14724);
and U15794 (N_15794,N_14491,N_15241);
nor U15795 (N_15795,N_15451,N_15042);
and U15796 (N_15796,N_15131,N_15121);
and U15797 (N_15797,N_15497,N_14436);
xnor U15798 (N_15798,N_15341,N_15575);
nand U15799 (N_15799,N_15339,N_15067);
or U15800 (N_15800,N_14926,N_15365);
or U15801 (N_15801,N_15504,N_14901);
nand U15802 (N_15802,N_14407,N_15439);
and U15803 (N_15803,N_14962,N_14613);
and U15804 (N_15804,N_15387,N_14514);
nand U15805 (N_15805,N_14561,N_14645);
nand U15806 (N_15806,N_14745,N_15142);
nor U15807 (N_15807,N_15205,N_14665);
or U15808 (N_15808,N_14406,N_14498);
nor U15809 (N_15809,N_15098,N_15520);
xnor U15810 (N_15810,N_15499,N_14826);
or U15811 (N_15811,N_15079,N_14772);
and U15812 (N_15812,N_15480,N_14714);
and U15813 (N_15813,N_15385,N_15053);
nor U15814 (N_15814,N_14412,N_15120);
nor U15815 (N_15815,N_15101,N_15425);
and U15816 (N_15816,N_14434,N_14641);
xor U15817 (N_15817,N_15443,N_15293);
or U15818 (N_15818,N_15134,N_14588);
nor U15819 (N_15819,N_15256,N_15413);
nand U15820 (N_15820,N_14997,N_15394);
xor U15821 (N_15821,N_15207,N_15056);
nor U15822 (N_15822,N_15028,N_15361);
xnor U15823 (N_15823,N_15284,N_14786);
and U15824 (N_15824,N_15537,N_14587);
nor U15825 (N_15825,N_14615,N_14972);
nor U15826 (N_15826,N_14453,N_15091);
xnor U15827 (N_15827,N_15250,N_15260);
nor U15828 (N_15828,N_14779,N_15008);
nor U15829 (N_15829,N_14580,N_15217);
nor U15830 (N_15830,N_14591,N_15181);
nor U15831 (N_15831,N_15030,N_14559);
nand U15832 (N_15832,N_15501,N_15589);
nor U15833 (N_15833,N_15059,N_15429);
nand U15834 (N_15834,N_14509,N_15447);
or U15835 (N_15835,N_14981,N_15432);
or U15836 (N_15836,N_14802,N_14608);
xor U15837 (N_15837,N_15231,N_15515);
and U15838 (N_15838,N_15483,N_15252);
nand U15839 (N_15839,N_15567,N_14682);
nor U15840 (N_15840,N_15105,N_15280);
nor U15841 (N_15841,N_14459,N_15297);
or U15842 (N_15842,N_14622,N_14651);
and U15843 (N_15843,N_14737,N_14529);
nor U15844 (N_15844,N_15313,N_14452);
nor U15845 (N_15845,N_14888,N_14685);
or U15846 (N_15846,N_14961,N_15535);
nand U15847 (N_15847,N_14563,N_15470);
or U15848 (N_15848,N_14865,N_15555);
or U15849 (N_15849,N_14479,N_15189);
nor U15850 (N_15850,N_14470,N_15072);
nor U15851 (N_15851,N_14892,N_14885);
nand U15852 (N_15852,N_15077,N_14941);
xor U15853 (N_15853,N_15090,N_14985);
nand U15854 (N_15854,N_14823,N_14771);
or U15855 (N_15855,N_15423,N_15540);
nor U15856 (N_15856,N_14789,N_15441);
and U15857 (N_15857,N_15518,N_15291);
nand U15858 (N_15858,N_14486,N_15402);
nand U15859 (N_15859,N_15577,N_14761);
and U15860 (N_15860,N_14528,N_15320);
nand U15861 (N_15861,N_15063,N_15288);
xor U15862 (N_15862,N_14548,N_15110);
nor U15863 (N_15863,N_15414,N_14423);
nor U15864 (N_15864,N_14648,N_15246);
or U15865 (N_15865,N_14538,N_14863);
and U15866 (N_15866,N_14799,N_14792);
xor U15867 (N_15867,N_15364,N_15568);
nor U15868 (N_15868,N_14524,N_14572);
xnor U15869 (N_15869,N_15415,N_15038);
or U15870 (N_15870,N_14477,N_14979);
xnor U15871 (N_15871,N_14429,N_14449);
and U15872 (N_15872,N_15550,N_15172);
or U15873 (N_15873,N_15191,N_15484);
and U15874 (N_15874,N_15025,N_15029);
or U15875 (N_15875,N_15174,N_14967);
xor U15876 (N_15876,N_15440,N_15149);
xnor U15877 (N_15877,N_14805,N_14754);
xnor U15878 (N_15878,N_15312,N_14609);
and U15879 (N_15879,N_15546,N_14577);
xnor U15880 (N_15880,N_14438,N_15511);
nor U15881 (N_15881,N_14690,N_15399);
nor U15882 (N_15882,N_14628,N_15554);
xor U15883 (N_15883,N_14447,N_14864);
nor U15884 (N_15884,N_14787,N_14534);
or U15885 (N_15885,N_14784,N_14636);
xnor U15886 (N_15886,N_15317,N_15162);
xor U15887 (N_15887,N_14567,N_15266);
or U15888 (N_15888,N_15526,N_14903);
nor U15889 (N_15889,N_14400,N_15248);
or U15890 (N_15890,N_14878,N_14833);
or U15891 (N_15891,N_14715,N_15357);
nor U15892 (N_15892,N_15338,N_15186);
nand U15893 (N_15893,N_15283,N_14816);
and U15894 (N_15894,N_15015,N_15118);
nand U15895 (N_15895,N_15219,N_14896);
and U15896 (N_15896,N_15557,N_14849);
or U15897 (N_15897,N_15421,N_15553);
and U15898 (N_15898,N_15411,N_15113);
or U15899 (N_15899,N_15373,N_14801);
or U15900 (N_15900,N_15180,N_15115);
xor U15901 (N_15901,N_15031,N_14800);
or U15902 (N_15902,N_15595,N_15182);
xor U15903 (N_15903,N_14770,N_14658);
nor U15904 (N_15904,N_14700,N_14838);
nor U15905 (N_15905,N_15369,N_15222);
nor U15906 (N_15906,N_15075,N_15343);
nor U15907 (N_15907,N_15331,N_14991);
and U15908 (N_15908,N_15517,N_15578);
and U15909 (N_15909,N_14667,N_14741);
or U15910 (N_15910,N_14974,N_15523);
xnor U15911 (N_15911,N_15522,N_14803);
nand U15912 (N_15912,N_14475,N_14859);
nor U15913 (N_15913,N_15337,N_14817);
nand U15914 (N_15914,N_15156,N_15016);
and U15915 (N_15915,N_15408,N_14681);
nor U15916 (N_15916,N_15167,N_14950);
xor U15917 (N_15917,N_15548,N_15588);
xnor U15918 (N_15918,N_14683,N_14873);
xor U15919 (N_15919,N_15416,N_15170);
nor U15920 (N_15920,N_15148,N_14425);
xor U15921 (N_15921,N_14906,N_15133);
or U15922 (N_15922,N_14720,N_15549);
nor U15923 (N_15923,N_14953,N_15478);
nand U15924 (N_15924,N_14813,N_14711);
and U15925 (N_15925,N_15208,N_15582);
and U15926 (N_15926,N_15212,N_15560);
nand U15927 (N_15927,N_14512,N_14846);
xor U15928 (N_15928,N_15116,N_15328);
nor U15929 (N_15929,N_14562,N_14469);
or U15930 (N_15930,N_15351,N_14924);
nor U15931 (N_15931,N_15534,N_15389);
xnor U15932 (N_15932,N_14842,N_15068);
nand U15933 (N_15933,N_14844,N_15489);
and U15934 (N_15934,N_15020,N_14420);
nor U15935 (N_15935,N_15307,N_15475);
and U15936 (N_15936,N_14728,N_14501);
and U15937 (N_15937,N_15500,N_15490);
nand U15938 (N_15938,N_14736,N_15407);
or U15939 (N_15939,N_15308,N_15556);
nor U15940 (N_15940,N_15378,N_14850);
nor U15941 (N_15941,N_15302,N_15319);
nor U15942 (N_15942,N_14494,N_14478);
nand U15943 (N_15943,N_14574,N_15287);
nand U15944 (N_15944,N_15479,N_14917);
nor U15945 (N_15945,N_14938,N_14912);
or U15946 (N_15946,N_15001,N_14749);
nand U15947 (N_15947,N_14598,N_14484);
and U15948 (N_15948,N_15409,N_15081);
xnor U15949 (N_15949,N_14808,N_15014);
or U15950 (N_15950,N_15579,N_14515);
or U15951 (N_15951,N_14485,N_14596);
and U15952 (N_15952,N_15435,N_15449);
or U15953 (N_15953,N_14481,N_14642);
nor U15954 (N_15954,N_14625,N_14834);
nor U15955 (N_15955,N_15227,N_15391);
nor U15956 (N_15956,N_15092,N_14516);
nor U15957 (N_15957,N_15257,N_14806);
and U15958 (N_15958,N_14471,N_15152);
xnor U15959 (N_15959,N_15039,N_15258);
nor U15960 (N_15960,N_15188,N_14732);
xor U15961 (N_15961,N_14751,N_15143);
xnor U15962 (N_15962,N_14819,N_15383);
xor U15963 (N_15963,N_15392,N_14913);
and U15964 (N_15964,N_15104,N_15057);
xnor U15965 (N_15965,N_14839,N_14969);
xnor U15966 (N_15966,N_14963,N_15333);
and U15967 (N_15967,N_14791,N_14623);
xor U15968 (N_15968,N_14513,N_14686);
nand U15969 (N_15969,N_14860,N_14442);
and U15970 (N_15970,N_14716,N_15405);
nor U15971 (N_15971,N_15137,N_15064);
nand U15972 (N_15972,N_14977,N_15544);
or U15973 (N_15973,N_15198,N_15345);
xor U15974 (N_15974,N_15462,N_14633);
xnor U15975 (N_15975,N_14767,N_14630);
and U15976 (N_15976,N_14777,N_14748);
xnor U15977 (N_15977,N_14717,N_15551);
xor U15978 (N_15978,N_15249,N_14499);
nor U15979 (N_15979,N_14467,N_15168);
xnor U15980 (N_15980,N_14581,N_15296);
nor U15981 (N_15981,N_15096,N_15235);
xnor U15982 (N_15982,N_15013,N_15236);
xor U15983 (N_15983,N_14807,N_14676);
and U15984 (N_15984,N_14911,N_15400);
or U15985 (N_15985,N_14500,N_15485);
nand U15986 (N_15986,N_14644,N_14647);
nor U15987 (N_15987,N_14866,N_14531);
nand U15988 (N_15988,N_14468,N_14666);
and U15989 (N_15989,N_14530,N_15281);
xnor U15990 (N_15990,N_15046,N_14689);
or U15991 (N_15991,N_14409,N_15303);
and U15992 (N_15992,N_15580,N_14544);
or U15993 (N_15993,N_15574,N_15210);
xor U15994 (N_15994,N_14855,N_14466);
or U15995 (N_15995,N_15264,N_15360);
or U15996 (N_15996,N_14403,N_15173);
or U15997 (N_15997,N_14916,N_15179);
nand U15998 (N_15998,N_14915,N_15424);
or U15999 (N_15999,N_14634,N_14718);
or U16000 (N_16000,N_14812,N_15187);
or U16001 (N_16001,N_15033,N_15456);
nand U16002 (N_16002,N_14547,N_14931);
nand U16003 (N_16003,N_14557,N_14585);
and U16004 (N_16004,N_15112,N_15040);
nand U16005 (N_16005,N_14444,N_15109);
nand U16006 (N_16006,N_14495,N_15080);
nand U16007 (N_16007,N_14918,N_14735);
xor U16008 (N_16008,N_15213,N_14611);
nor U16009 (N_16009,N_14417,N_14653);
or U16010 (N_16010,N_15516,N_15035);
and U16011 (N_16011,N_14699,N_14450);
nor U16012 (N_16012,N_14954,N_15426);
xnor U16013 (N_16013,N_15508,N_14688);
xnor U16014 (N_16014,N_14697,N_15314);
xnor U16015 (N_16015,N_15275,N_14566);
and U16016 (N_16016,N_14704,N_15108);
or U16017 (N_16017,N_14440,N_14740);
or U16018 (N_16018,N_14811,N_14957);
or U16019 (N_16019,N_14733,N_15463);
nand U16020 (N_16020,N_14773,N_15461);
or U16021 (N_16021,N_15458,N_14738);
xnor U16022 (N_16022,N_15327,N_14496);
and U16023 (N_16023,N_15123,N_14465);
nor U16024 (N_16024,N_14861,N_14419);
nand U16025 (N_16025,N_15285,N_14986);
and U16026 (N_16026,N_15306,N_15545);
nand U16027 (N_16027,N_14874,N_14517);
nand U16028 (N_16028,N_14492,N_14781);
xnor U16029 (N_16029,N_14672,N_14695);
nor U16030 (N_16030,N_14639,N_14818);
nand U16031 (N_16031,N_15276,N_14674);
or U16032 (N_16032,N_15024,N_15430);
nand U16033 (N_16033,N_15126,N_14710);
nor U16034 (N_16034,N_15366,N_14539);
xor U16035 (N_16035,N_15596,N_15438);
nand U16036 (N_16036,N_14693,N_14680);
and U16037 (N_16037,N_14904,N_14411);
nand U16038 (N_16038,N_15216,N_15486);
nor U16039 (N_16039,N_15093,N_14990);
nor U16040 (N_16040,N_15536,N_14763);
nor U16041 (N_16041,N_15177,N_14929);
and U16042 (N_16042,N_15278,N_14744);
or U16043 (N_16043,N_14678,N_14872);
nand U16044 (N_16044,N_15274,N_15032);
xnor U16045 (N_16045,N_15325,N_15585);
or U16046 (N_16046,N_15017,N_14568);
nand U16047 (N_16047,N_15003,N_14663);
nor U16048 (N_16048,N_15543,N_15103);
xnor U16049 (N_16049,N_14701,N_15159);
nand U16050 (N_16050,N_15247,N_14821);
nand U16051 (N_16051,N_15279,N_15332);
and U16052 (N_16052,N_15083,N_15530);
and U16053 (N_16053,N_14775,N_14757);
and U16054 (N_16054,N_14856,N_14600);
and U16055 (N_16055,N_15427,N_15012);
xnor U16056 (N_16056,N_15021,N_15433);
xnor U16057 (N_16057,N_14461,N_14435);
xor U16058 (N_16058,N_15226,N_14942);
or U16059 (N_16059,N_14661,N_15528);
xor U16060 (N_16060,N_14964,N_14822);
nand U16061 (N_16061,N_15542,N_14927);
nand U16062 (N_16062,N_14472,N_14656);
and U16063 (N_16063,N_14712,N_14679);
nand U16064 (N_16064,N_15060,N_15541);
nor U16065 (N_16065,N_14556,N_14910);
and U16066 (N_16066,N_14483,N_15410);
nor U16067 (N_16067,N_14595,N_15446);
and U16068 (N_16068,N_15487,N_15271);
xnor U16069 (N_16069,N_15251,N_14424);
and U16070 (N_16070,N_14768,N_15111);
xnor U16071 (N_16071,N_15467,N_14793);
nand U16072 (N_16072,N_15146,N_14752);
or U16073 (N_16073,N_15356,N_15272);
or U16074 (N_16074,N_15591,N_14670);
nor U16075 (N_16075,N_14976,N_14898);
nand U16076 (N_16076,N_15300,N_14778);
xor U16077 (N_16077,N_14843,N_14677);
and U16078 (N_16078,N_14586,N_14696);
nand U16079 (N_16079,N_15368,N_14414);
xor U16080 (N_16080,N_15051,N_14583);
nor U16081 (N_16081,N_14933,N_15061);
nand U16082 (N_16082,N_14936,N_14966);
nand U16083 (N_16083,N_15448,N_14637);
and U16084 (N_16084,N_14923,N_15457);
and U16085 (N_16085,N_15454,N_15482);
xnor U16086 (N_16086,N_14457,N_14920);
nand U16087 (N_16087,N_14907,N_15506);
or U16088 (N_16088,N_15564,N_14919);
or U16089 (N_16089,N_14521,N_15353);
xnor U16090 (N_16090,N_15381,N_14455);
nor U16091 (N_16091,N_14945,N_15004);
nor U16092 (N_16092,N_15027,N_15214);
xnor U16093 (N_16093,N_14871,N_14829);
nand U16094 (N_16094,N_14522,N_15047);
and U16095 (N_16095,N_14555,N_15140);
and U16096 (N_16096,N_15000,N_14523);
nand U16097 (N_16097,N_15237,N_15007);
or U16098 (N_16098,N_14788,N_15185);
xnor U16099 (N_16099,N_14493,N_15220);
nor U16100 (N_16100,N_14652,N_14747);
or U16101 (N_16101,N_15263,N_15397);
or U16102 (N_16102,N_15200,N_15147);
xor U16103 (N_16103,N_14886,N_15292);
xnor U16104 (N_16104,N_14694,N_14687);
and U16105 (N_16105,N_15102,N_14851);
nor U16106 (N_16106,N_14867,N_15122);
nor U16107 (N_16107,N_15417,N_14774);
xnor U16108 (N_16108,N_14766,N_15586);
xor U16109 (N_16109,N_15107,N_14879);
nor U16110 (N_16110,N_14664,N_15268);
nor U16111 (N_16111,N_15565,N_14894);
nor U16112 (N_16112,N_15512,N_14742);
nor U16113 (N_16113,N_14999,N_14955);
nor U16114 (N_16114,N_14764,N_14940);
and U16115 (N_16115,N_15166,N_14881);
or U16116 (N_16116,N_14558,N_15150);
nor U16117 (N_16117,N_14820,N_14428);
or U16118 (N_16118,N_14410,N_15065);
xnor U16119 (N_16119,N_15136,N_15347);
and U16120 (N_16120,N_15041,N_15436);
and U16121 (N_16121,N_15161,N_15311);
or U16122 (N_16122,N_14576,N_15547);
and U16123 (N_16123,N_15178,N_15404);
nand U16124 (N_16124,N_15593,N_15232);
and U16125 (N_16125,N_15342,N_15401);
xor U16126 (N_16126,N_14730,N_14815);
and U16127 (N_16127,N_15135,N_15176);
or U16128 (N_16128,N_14606,N_15055);
and U16129 (N_16129,N_14605,N_14668);
xor U16130 (N_16130,N_14707,N_14404);
and U16131 (N_16131,N_14439,N_14684);
or U16132 (N_16132,N_14502,N_15234);
or U16133 (N_16133,N_15286,N_15242);
nand U16134 (N_16134,N_14837,N_15244);
or U16135 (N_16135,N_15192,N_14810);
and U16136 (N_16136,N_14959,N_14965);
nor U16137 (N_16137,N_15363,N_15465);
or U16138 (N_16138,N_14993,N_15305);
and U16139 (N_16139,N_15474,N_15335);
or U16140 (N_16140,N_14824,N_14882);
and U16141 (N_16141,N_15099,N_14734);
xor U16142 (N_16142,N_15488,N_14845);
xor U16143 (N_16143,N_15527,N_14607);
xnor U16144 (N_16144,N_15492,N_14594);
xor U16145 (N_16145,N_15406,N_15471);
and U16146 (N_16146,N_15395,N_14987);
nor U16147 (N_16147,N_14939,N_15019);
nor U16148 (N_16148,N_15377,N_14739);
nand U16149 (N_16149,N_14507,N_15367);
and U16150 (N_16150,N_15370,N_14729);
xnor U16151 (N_16151,N_14649,N_14638);
nor U16152 (N_16152,N_14599,N_15034);
nor U16153 (N_16153,N_15002,N_15496);
nor U16154 (N_16154,N_14956,N_15255);
nor U16155 (N_16155,N_14835,N_15495);
and U16156 (N_16156,N_14427,N_14935);
xnor U16157 (N_16157,N_14725,N_14755);
nor U16158 (N_16158,N_15445,N_14503);
nor U16159 (N_16159,N_14809,N_14464);
xnor U16160 (N_16160,N_14840,N_15531);
and U16161 (N_16161,N_15382,N_14659);
and U16162 (N_16162,N_14949,N_15215);
nand U16163 (N_16163,N_14705,N_14454);
and U16164 (N_16164,N_15138,N_14890);
xnor U16165 (N_16165,N_15269,N_15375);
or U16166 (N_16166,N_14709,N_14847);
xor U16167 (N_16167,N_15583,N_15379);
or U16168 (N_16168,N_14825,N_14869);
nor U16169 (N_16169,N_15218,N_15562);
and U16170 (N_16170,N_15043,N_15358);
xor U16171 (N_16171,N_14635,N_15078);
or U16172 (N_16172,N_15561,N_15169);
xor U16173 (N_16173,N_14497,N_15071);
nor U16174 (N_16174,N_14456,N_14540);
nand U16175 (N_16175,N_15539,N_15346);
xnor U16176 (N_16176,N_14984,N_15298);
nand U16177 (N_16177,N_15388,N_14614);
nand U16178 (N_16178,N_14597,N_14804);
and U16179 (N_16179,N_14743,N_14445);
xnor U16180 (N_16180,N_14552,N_14487);
nor U16181 (N_16181,N_14564,N_15117);
and U16182 (N_16182,N_15141,N_15100);
nand U16183 (N_16183,N_14970,N_14418);
xnor U16184 (N_16184,N_15267,N_14527);
xor U16185 (N_16185,N_14565,N_15052);
and U16186 (N_16186,N_14657,N_15224);
xor U16187 (N_16187,N_15299,N_14437);
nor U16188 (N_16188,N_15597,N_14944);
nand U16189 (N_16189,N_15598,N_15037);
and U16190 (N_16190,N_14460,N_15151);
and U16191 (N_16191,N_14983,N_15321);
nand U16192 (N_16192,N_14782,N_14416);
nor U16193 (N_16193,N_15049,N_14783);
nand U16194 (N_16194,N_15175,N_14535);
xor U16195 (N_16195,N_14590,N_14980);
xnor U16196 (N_16196,N_14518,N_14973);
xor U16197 (N_16197,N_15323,N_15209);
and U16198 (N_16198,N_14408,N_14759);
nand U16199 (N_16199,N_14713,N_14852);
or U16200 (N_16200,N_15078,N_15353);
xnor U16201 (N_16201,N_15261,N_14848);
xnor U16202 (N_16202,N_15299,N_15174);
xnor U16203 (N_16203,N_14445,N_15079);
nor U16204 (N_16204,N_14477,N_15583);
or U16205 (N_16205,N_15020,N_14456);
nor U16206 (N_16206,N_14914,N_14797);
nand U16207 (N_16207,N_14998,N_14770);
xor U16208 (N_16208,N_14962,N_15406);
or U16209 (N_16209,N_14975,N_15568);
or U16210 (N_16210,N_15343,N_15333);
nand U16211 (N_16211,N_15049,N_14991);
nand U16212 (N_16212,N_15595,N_15153);
nor U16213 (N_16213,N_15297,N_15073);
and U16214 (N_16214,N_15233,N_15150);
or U16215 (N_16215,N_14587,N_14424);
or U16216 (N_16216,N_14605,N_14732);
xor U16217 (N_16217,N_14637,N_15138);
nand U16218 (N_16218,N_15153,N_14706);
nor U16219 (N_16219,N_14472,N_14854);
nor U16220 (N_16220,N_14978,N_15171);
and U16221 (N_16221,N_14531,N_15111);
and U16222 (N_16222,N_14955,N_15155);
nor U16223 (N_16223,N_14514,N_14682);
and U16224 (N_16224,N_14438,N_15428);
xor U16225 (N_16225,N_15168,N_14603);
and U16226 (N_16226,N_14967,N_14509);
or U16227 (N_16227,N_14679,N_14787);
nand U16228 (N_16228,N_15480,N_14914);
and U16229 (N_16229,N_15056,N_15381);
xnor U16230 (N_16230,N_14416,N_15115);
nand U16231 (N_16231,N_14967,N_14920);
and U16232 (N_16232,N_15175,N_14732);
xor U16233 (N_16233,N_15089,N_14826);
and U16234 (N_16234,N_15582,N_15204);
xor U16235 (N_16235,N_14957,N_15312);
xor U16236 (N_16236,N_14732,N_15311);
or U16237 (N_16237,N_14558,N_14824);
nand U16238 (N_16238,N_15434,N_14483);
or U16239 (N_16239,N_14783,N_14409);
or U16240 (N_16240,N_15133,N_15520);
xnor U16241 (N_16241,N_14616,N_14488);
and U16242 (N_16242,N_14770,N_14827);
nor U16243 (N_16243,N_14847,N_14920);
xnor U16244 (N_16244,N_14553,N_15459);
and U16245 (N_16245,N_14505,N_15125);
nor U16246 (N_16246,N_15210,N_14918);
and U16247 (N_16247,N_14600,N_14403);
nor U16248 (N_16248,N_14829,N_14697);
or U16249 (N_16249,N_15056,N_15169);
nand U16250 (N_16250,N_15559,N_14615);
and U16251 (N_16251,N_14664,N_15061);
nor U16252 (N_16252,N_15225,N_14468);
or U16253 (N_16253,N_14991,N_15568);
and U16254 (N_16254,N_15366,N_14455);
xnor U16255 (N_16255,N_15320,N_14435);
nand U16256 (N_16256,N_14591,N_15049);
or U16257 (N_16257,N_15343,N_15160);
nor U16258 (N_16258,N_15426,N_15033);
or U16259 (N_16259,N_14808,N_15360);
or U16260 (N_16260,N_15114,N_15315);
and U16261 (N_16261,N_15235,N_14788);
or U16262 (N_16262,N_15055,N_14647);
xor U16263 (N_16263,N_14699,N_14443);
xor U16264 (N_16264,N_15051,N_14613);
xor U16265 (N_16265,N_15442,N_15208);
and U16266 (N_16266,N_15258,N_14550);
nor U16267 (N_16267,N_15230,N_14970);
nor U16268 (N_16268,N_14830,N_14551);
xnor U16269 (N_16269,N_14860,N_14595);
nor U16270 (N_16270,N_14446,N_15016);
xor U16271 (N_16271,N_14707,N_15199);
nand U16272 (N_16272,N_15280,N_14668);
and U16273 (N_16273,N_15592,N_14564);
xnor U16274 (N_16274,N_15553,N_15496);
xor U16275 (N_16275,N_14483,N_15542);
nand U16276 (N_16276,N_15208,N_14991);
or U16277 (N_16277,N_15297,N_14500);
xor U16278 (N_16278,N_14894,N_15196);
xor U16279 (N_16279,N_15350,N_15383);
xor U16280 (N_16280,N_15122,N_15011);
or U16281 (N_16281,N_14436,N_14746);
nand U16282 (N_16282,N_15108,N_14470);
nand U16283 (N_16283,N_15386,N_15550);
nor U16284 (N_16284,N_15462,N_15198);
nand U16285 (N_16285,N_14507,N_15590);
nor U16286 (N_16286,N_15205,N_15500);
nand U16287 (N_16287,N_14995,N_14408);
nand U16288 (N_16288,N_15409,N_15088);
xnor U16289 (N_16289,N_14680,N_15094);
or U16290 (N_16290,N_14619,N_15431);
nand U16291 (N_16291,N_14850,N_14848);
and U16292 (N_16292,N_15244,N_15525);
and U16293 (N_16293,N_14491,N_14626);
and U16294 (N_16294,N_15375,N_15319);
nand U16295 (N_16295,N_15078,N_14576);
and U16296 (N_16296,N_15398,N_15017);
xnor U16297 (N_16297,N_14989,N_14574);
or U16298 (N_16298,N_15109,N_15463);
and U16299 (N_16299,N_15333,N_15582);
or U16300 (N_16300,N_15385,N_15411);
nand U16301 (N_16301,N_14883,N_14727);
xnor U16302 (N_16302,N_15070,N_15072);
nand U16303 (N_16303,N_14625,N_14849);
or U16304 (N_16304,N_15554,N_14760);
nor U16305 (N_16305,N_15420,N_14842);
xnor U16306 (N_16306,N_15104,N_14971);
nor U16307 (N_16307,N_14519,N_15080);
nor U16308 (N_16308,N_15454,N_14515);
or U16309 (N_16309,N_15332,N_14903);
xor U16310 (N_16310,N_15110,N_15138);
and U16311 (N_16311,N_15451,N_14835);
or U16312 (N_16312,N_15172,N_15315);
nand U16313 (N_16313,N_14647,N_14962);
nand U16314 (N_16314,N_14560,N_14874);
nor U16315 (N_16315,N_14580,N_15091);
xnor U16316 (N_16316,N_15062,N_14983);
and U16317 (N_16317,N_14963,N_14700);
or U16318 (N_16318,N_15460,N_15377);
nor U16319 (N_16319,N_15457,N_14976);
or U16320 (N_16320,N_14485,N_15415);
xor U16321 (N_16321,N_14650,N_14930);
xnor U16322 (N_16322,N_15443,N_14506);
or U16323 (N_16323,N_14678,N_14910);
nor U16324 (N_16324,N_14546,N_14544);
nor U16325 (N_16325,N_14675,N_15310);
or U16326 (N_16326,N_15087,N_14719);
xnor U16327 (N_16327,N_14858,N_14897);
and U16328 (N_16328,N_15451,N_15355);
xnor U16329 (N_16329,N_15044,N_15339);
xnor U16330 (N_16330,N_14422,N_14676);
xnor U16331 (N_16331,N_14766,N_15218);
and U16332 (N_16332,N_14684,N_14508);
nand U16333 (N_16333,N_15136,N_15483);
nand U16334 (N_16334,N_15445,N_14453);
nand U16335 (N_16335,N_15242,N_15366);
and U16336 (N_16336,N_15007,N_15419);
and U16337 (N_16337,N_15468,N_15104);
xor U16338 (N_16338,N_15031,N_15008);
nand U16339 (N_16339,N_14812,N_15203);
or U16340 (N_16340,N_15568,N_15491);
nand U16341 (N_16341,N_14862,N_14679);
and U16342 (N_16342,N_14965,N_15540);
nor U16343 (N_16343,N_14689,N_14467);
nor U16344 (N_16344,N_15417,N_14721);
nand U16345 (N_16345,N_14518,N_14783);
nand U16346 (N_16346,N_15529,N_14691);
nand U16347 (N_16347,N_15426,N_14691);
xor U16348 (N_16348,N_15084,N_15392);
nor U16349 (N_16349,N_14477,N_14573);
xnor U16350 (N_16350,N_15203,N_15242);
xor U16351 (N_16351,N_14670,N_14898);
nor U16352 (N_16352,N_15435,N_14470);
xor U16353 (N_16353,N_15315,N_14891);
xnor U16354 (N_16354,N_15145,N_15367);
nor U16355 (N_16355,N_14585,N_14786);
and U16356 (N_16356,N_15530,N_14674);
and U16357 (N_16357,N_14648,N_15345);
xnor U16358 (N_16358,N_15150,N_15141);
or U16359 (N_16359,N_14742,N_15299);
xor U16360 (N_16360,N_15216,N_14601);
nand U16361 (N_16361,N_15503,N_15058);
or U16362 (N_16362,N_14455,N_14916);
nor U16363 (N_16363,N_14711,N_15089);
and U16364 (N_16364,N_14671,N_14619);
xor U16365 (N_16365,N_15563,N_14893);
or U16366 (N_16366,N_15270,N_14674);
nand U16367 (N_16367,N_14873,N_14851);
nand U16368 (N_16368,N_14787,N_14995);
nand U16369 (N_16369,N_14861,N_14539);
nand U16370 (N_16370,N_15342,N_14634);
xnor U16371 (N_16371,N_15236,N_14955);
nor U16372 (N_16372,N_14977,N_14856);
nand U16373 (N_16373,N_14630,N_14761);
nor U16374 (N_16374,N_14601,N_15100);
and U16375 (N_16375,N_14516,N_14701);
nor U16376 (N_16376,N_14439,N_14677);
nor U16377 (N_16377,N_15363,N_14647);
xor U16378 (N_16378,N_15583,N_14967);
nand U16379 (N_16379,N_15460,N_14912);
or U16380 (N_16380,N_15572,N_15035);
nor U16381 (N_16381,N_14951,N_14606);
xor U16382 (N_16382,N_15181,N_14529);
and U16383 (N_16383,N_14896,N_14956);
nand U16384 (N_16384,N_15332,N_15084);
and U16385 (N_16385,N_14414,N_15459);
nand U16386 (N_16386,N_14802,N_15174);
xnor U16387 (N_16387,N_14733,N_15032);
nand U16388 (N_16388,N_14936,N_14988);
or U16389 (N_16389,N_15498,N_15599);
nand U16390 (N_16390,N_15075,N_15164);
nand U16391 (N_16391,N_15459,N_15107);
xnor U16392 (N_16392,N_14979,N_14941);
xor U16393 (N_16393,N_14555,N_15199);
xor U16394 (N_16394,N_15360,N_14498);
and U16395 (N_16395,N_15305,N_14592);
or U16396 (N_16396,N_14404,N_14683);
or U16397 (N_16397,N_15133,N_14789);
nand U16398 (N_16398,N_14414,N_15086);
xnor U16399 (N_16399,N_14810,N_15200);
or U16400 (N_16400,N_15404,N_14469);
xor U16401 (N_16401,N_15156,N_14783);
and U16402 (N_16402,N_15044,N_14514);
nand U16403 (N_16403,N_15262,N_15269);
nor U16404 (N_16404,N_14838,N_15596);
xor U16405 (N_16405,N_14682,N_15394);
and U16406 (N_16406,N_14674,N_14682);
and U16407 (N_16407,N_14928,N_15003);
or U16408 (N_16408,N_14652,N_14984);
nor U16409 (N_16409,N_14563,N_14725);
nand U16410 (N_16410,N_14957,N_14949);
nor U16411 (N_16411,N_14513,N_15452);
nand U16412 (N_16412,N_15123,N_14478);
nand U16413 (N_16413,N_15317,N_14928);
nand U16414 (N_16414,N_15195,N_15555);
and U16415 (N_16415,N_14638,N_15343);
xnor U16416 (N_16416,N_14763,N_14998);
nor U16417 (N_16417,N_14703,N_14686);
and U16418 (N_16418,N_15209,N_15066);
or U16419 (N_16419,N_14847,N_14785);
xor U16420 (N_16420,N_15593,N_15145);
nor U16421 (N_16421,N_15155,N_14560);
and U16422 (N_16422,N_15086,N_15068);
nand U16423 (N_16423,N_15051,N_15581);
nor U16424 (N_16424,N_14500,N_14584);
nor U16425 (N_16425,N_15230,N_15059);
xnor U16426 (N_16426,N_15395,N_15424);
xnor U16427 (N_16427,N_15576,N_15231);
and U16428 (N_16428,N_15233,N_14763);
xor U16429 (N_16429,N_15060,N_15495);
or U16430 (N_16430,N_14717,N_14849);
nor U16431 (N_16431,N_14728,N_14946);
and U16432 (N_16432,N_15168,N_15573);
and U16433 (N_16433,N_14815,N_14597);
and U16434 (N_16434,N_14526,N_14596);
nor U16435 (N_16435,N_15343,N_14460);
nor U16436 (N_16436,N_15255,N_14782);
nor U16437 (N_16437,N_14580,N_15278);
or U16438 (N_16438,N_14582,N_14425);
xnor U16439 (N_16439,N_14737,N_15101);
nor U16440 (N_16440,N_15259,N_14820);
and U16441 (N_16441,N_14499,N_14615);
nand U16442 (N_16442,N_14651,N_14669);
or U16443 (N_16443,N_15131,N_14511);
and U16444 (N_16444,N_15339,N_14938);
or U16445 (N_16445,N_14857,N_15477);
or U16446 (N_16446,N_14520,N_15253);
nand U16447 (N_16447,N_15295,N_14458);
xnor U16448 (N_16448,N_15555,N_15244);
xnor U16449 (N_16449,N_14433,N_14493);
nor U16450 (N_16450,N_15484,N_14562);
and U16451 (N_16451,N_15367,N_14453);
and U16452 (N_16452,N_15140,N_15126);
and U16453 (N_16453,N_15596,N_14709);
xnor U16454 (N_16454,N_15349,N_14652);
and U16455 (N_16455,N_14994,N_14551);
and U16456 (N_16456,N_15161,N_15557);
or U16457 (N_16457,N_15187,N_15146);
or U16458 (N_16458,N_14977,N_14649);
nand U16459 (N_16459,N_14602,N_15174);
xnor U16460 (N_16460,N_14792,N_15482);
and U16461 (N_16461,N_15438,N_14944);
or U16462 (N_16462,N_15594,N_14706);
nor U16463 (N_16463,N_15529,N_15395);
and U16464 (N_16464,N_15157,N_15586);
or U16465 (N_16465,N_15340,N_14437);
or U16466 (N_16466,N_15330,N_14430);
xor U16467 (N_16467,N_15156,N_14435);
nor U16468 (N_16468,N_14960,N_14754);
and U16469 (N_16469,N_14877,N_15382);
and U16470 (N_16470,N_15284,N_14756);
xor U16471 (N_16471,N_15182,N_15567);
or U16472 (N_16472,N_15387,N_15262);
or U16473 (N_16473,N_14786,N_14957);
and U16474 (N_16474,N_14814,N_14428);
nor U16475 (N_16475,N_14503,N_15070);
xor U16476 (N_16476,N_15051,N_15515);
and U16477 (N_16477,N_14780,N_14574);
nor U16478 (N_16478,N_14401,N_15407);
xor U16479 (N_16479,N_14889,N_14976);
nand U16480 (N_16480,N_15372,N_15592);
nand U16481 (N_16481,N_14763,N_14988);
nor U16482 (N_16482,N_14811,N_14964);
nand U16483 (N_16483,N_14895,N_15095);
and U16484 (N_16484,N_15459,N_14523);
and U16485 (N_16485,N_14608,N_15379);
nand U16486 (N_16486,N_15469,N_15490);
xor U16487 (N_16487,N_14805,N_14556);
or U16488 (N_16488,N_15511,N_14434);
or U16489 (N_16489,N_15562,N_14666);
nand U16490 (N_16490,N_14599,N_14845);
xnor U16491 (N_16491,N_15457,N_15182);
or U16492 (N_16492,N_14728,N_14766);
xor U16493 (N_16493,N_15301,N_15055);
nand U16494 (N_16494,N_15057,N_15008);
and U16495 (N_16495,N_15072,N_15448);
and U16496 (N_16496,N_15529,N_15194);
nand U16497 (N_16497,N_15172,N_14513);
nor U16498 (N_16498,N_14487,N_15483);
and U16499 (N_16499,N_14524,N_14588);
xnor U16500 (N_16500,N_14491,N_15074);
nand U16501 (N_16501,N_15465,N_14852);
and U16502 (N_16502,N_15275,N_14907);
and U16503 (N_16503,N_14949,N_15226);
xor U16504 (N_16504,N_15411,N_15329);
and U16505 (N_16505,N_15475,N_14761);
or U16506 (N_16506,N_15113,N_15330);
and U16507 (N_16507,N_14826,N_14509);
nand U16508 (N_16508,N_14798,N_14442);
nand U16509 (N_16509,N_14636,N_15021);
and U16510 (N_16510,N_14853,N_14668);
xor U16511 (N_16511,N_14803,N_15080);
or U16512 (N_16512,N_14915,N_14997);
nand U16513 (N_16513,N_15218,N_14484);
and U16514 (N_16514,N_14948,N_14723);
or U16515 (N_16515,N_15539,N_14836);
nor U16516 (N_16516,N_15059,N_14753);
nand U16517 (N_16517,N_14790,N_15442);
or U16518 (N_16518,N_15354,N_14641);
or U16519 (N_16519,N_15007,N_14539);
nand U16520 (N_16520,N_15322,N_15407);
nand U16521 (N_16521,N_15536,N_14710);
or U16522 (N_16522,N_14841,N_15144);
nor U16523 (N_16523,N_14972,N_15512);
and U16524 (N_16524,N_14617,N_14993);
and U16525 (N_16525,N_14862,N_14411);
or U16526 (N_16526,N_14691,N_14499);
xnor U16527 (N_16527,N_14474,N_14436);
and U16528 (N_16528,N_14583,N_15089);
nor U16529 (N_16529,N_15194,N_14422);
nor U16530 (N_16530,N_14880,N_14730);
nand U16531 (N_16531,N_15146,N_14865);
and U16532 (N_16532,N_14527,N_15108);
nand U16533 (N_16533,N_15163,N_14656);
nor U16534 (N_16534,N_15406,N_14696);
nand U16535 (N_16535,N_14814,N_14503);
and U16536 (N_16536,N_14961,N_15468);
nand U16537 (N_16537,N_14789,N_14788);
nor U16538 (N_16538,N_14497,N_15154);
nor U16539 (N_16539,N_14457,N_15329);
and U16540 (N_16540,N_14529,N_15500);
nor U16541 (N_16541,N_14819,N_14638);
nor U16542 (N_16542,N_14549,N_15560);
xnor U16543 (N_16543,N_14698,N_14958);
and U16544 (N_16544,N_14538,N_14541);
nand U16545 (N_16545,N_15474,N_14993);
nand U16546 (N_16546,N_14419,N_15233);
and U16547 (N_16547,N_15307,N_14840);
xor U16548 (N_16548,N_14538,N_15421);
xor U16549 (N_16549,N_15515,N_14712);
or U16550 (N_16550,N_15417,N_15355);
and U16551 (N_16551,N_15548,N_15324);
nor U16552 (N_16552,N_15378,N_14823);
and U16553 (N_16553,N_14907,N_15564);
nand U16554 (N_16554,N_15045,N_15208);
xor U16555 (N_16555,N_14426,N_15403);
and U16556 (N_16556,N_14763,N_14633);
or U16557 (N_16557,N_15477,N_14687);
xnor U16558 (N_16558,N_14763,N_15400);
and U16559 (N_16559,N_14591,N_14877);
nor U16560 (N_16560,N_15285,N_15204);
nor U16561 (N_16561,N_15438,N_15281);
and U16562 (N_16562,N_15057,N_15534);
nor U16563 (N_16563,N_15477,N_14722);
nor U16564 (N_16564,N_14559,N_14560);
xor U16565 (N_16565,N_14945,N_15254);
and U16566 (N_16566,N_14686,N_14769);
nand U16567 (N_16567,N_15539,N_15341);
and U16568 (N_16568,N_15007,N_14971);
and U16569 (N_16569,N_15192,N_14829);
nand U16570 (N_16570,N_15275,N_14582);
nand U16571 (N_16571,N_15551,N_15087);
or U16572 (N_16572,N_14709,N_15529);
nand U16573 (N_16573,N_14675,N_14472);
nand U16574 (N_16574,N_15231,N_15390);
nor U16575 (N_16575,N_14633,N_15020);
or U16576 (N_16576,N_15292,N_15459);
nor U16577 (N_16577,N_14454,N_15473);
nor U16578 (N_16578,N_14931,N_15123);
nand U16579 (N_16579,N_14932,N_14676);
or U16580 (N_16580,N_14618,N_14621);
or U16581 (N_16581,N_14706,N_15051);
or U16582 (N_16582,N_14584,N_14402);
and U16583 (N_16583,N_14930,N_14444);
nand U16584 (N_16584,N_14556,N_14866);
and U16585 (N_16585,N_14668,N_15529);
xnor U16586 (N_16586,N_15034,N_14416);
or U16587 (N_16587,N_14934,N_14896);
xnor U16588 (N_16588,N_15204,N_14406);
and U16589 (N_16589,N_14747,N_14951);
xnor U16590 (N_16590,N_14567,N_14716);
nand U16591 (N_16591,N_14479,N_15182);
or U16592 (N_16592,N_15591,N_14568);
xor U16593 (N_16593,N_14740,N_14976);
nor U16594 (N_16594,N_14574,N_14490);
and U16595 (N_16595,N_15148,N_15180);
nand U16596 (N_16596,N_14638,N_15320);
nand U16597 (N_16597,N_14720,N_14934);
nand U16598 (N_16598,N_15479,N_15397);
nand U16599 (N_16599,N_14696,N_14437);
nand U16600 (N_16600,N_14541,N_14639);
and U16601 (N_16601,N_15497,N_14776);
nand U16602 (N_16602,N_15240,N_15477);
xor U16603 (N_16603,N_15052,N_14965);
nand U16604 (N_16604,N_14796,N_14562);
and U16605 (N_16605,N_14993,N_15086);
or U16606 (N_16606,N_15426,N_15122);
nand U16607 (N_16607,N_15039,N_14651);
nand U16608 (N_16608,N_15146,N_15064);
nor U16609 (N_16609,N_15196,N_15378);
xor U16610 (N_16610,N_14455,N_14940);
or U16611 (N_16611,N_15503,N_15018);
nand U16612 (N_16612,N_15576,N_15134);
and U16613 (N_16613,N_14636,N_14423);
and U16614 (N_16614,N_15046,N_14996);
nor U16615 (N_16615,N_15106,N_14843);
xnor U16616 (N_16616,N_14809,N_14482);
or U16617 (N_16617,N_14872,N_14851);
nor U16618 (N_16618,N_15114,N_15158);
nand U16619 (N_16619,N_14555,N_15550);
nor U16620 (N_16620,N_14509,N_14733);
xnor U16621 (N_16621,N_15306,N_15556);
and U16622 (N_16622,N_14771,N_14402);
xnor U16623 (N_16623,N_15215,N_14948);
or U16624 (N_16624,N_15503,N_15597);
nor U16625 (N_16625,N_15540,N_14723);
or U16626 (N_16626,N_15296,N_14713);
xor U16627 (N_16627,N_14509,N_15502);
xnor U16628 (N_16628,N_15392,N_15351);
and U16629 (N_16629,N_14676,N_15132);
xnor U16630 (N_16630,N_15289,N_15131);
nor U16631 (N_16631,N_14991,N_14564);
and U16632 (N_16632,N_15455,N_14585);
and U16633 (N_16633,N_15372,N_14857);
xor U16634 (N_16634,N_15119,N_14616);
nor U16635 (N_16635,N_15037,N_15395);
nor U16636 (N_16636,N_15182,N_14731);
nand U16637 (N_16637,N_14704,N_15423);
or U16638 (N_16638,N_15383,N_14569);
xor U16639 (N_16639,N_14419,N_14859);
xor U16640 (N_16640,N_15356,N_14517);
nand U16641 (N_16641,N_14476,N_14536);
nand U16642 (N_16642,N_15044,N_15544);
nor U16643 (N_16643,N_15473,N_14847);
nand U16644 (N_16644,N_14731,N_14559);
xnor U16645 (N_16645,N_15048,N_15530);
nand U16646 (N_16646,N_15266,N_14490);
xor U16647 (N_16647,N_14686,N_15287);
xnor U16648 (N_16648,N_15193,N_15336);
nand U16649 (N_16649,N_14979,N_14878);
nor U16650 (N_16650,N_15426,N_15068);
nand U16651 (N_16651,N_14821,N_15365);
or U16652 (N_16652,N_15290,N_14877);
nand U16653 (N_16653,N_14414,N_14925);
nand U16654 (N_16654,N_14550,N_14784);
or U16655 (N_16655,N_15306,N_14649);
xor U16656 (N_16656,N_15132,N_15205);
nor U16657 (N_16657,N_14712,N_15258);
or U16658 (N_16658,N_14743,N_15388);
nand U16659 (N_16659,N_15116,N_14698);
and U16660 (N_16660,N_14673,N_14641);
xnor U16661 (N_16661,N_15365,N_15239);
nand U16662 (N_16662,N_14923,N_15396);
and U16663 (N_16663,N_14806,N_14695);
nor U16664 (N_16664,N_14628,N_15490);
or U16665 (N_16665,N_15044,N_14819);
xnor U16666 (N_16666,N_15073,N_15380);
and U16667 (N_16667,N_15410,N_14853);
or U16668 (N_16668,N_15160,N_14992);
nand U16669 (N_16669,N_15559,N_14973);
or U16670 (N_16670,N_14975,N_14525);
and U16671 (N_16671,N_15565,N_14481);
xnor U16672 (N_16672,N_14426,N_15222);
nand U16673 (N_16673,N_15408,N_15446);
or U16674 (N_16674,N_15179,N_14740);
nand U16675 (N_16675,N_14414,N_14729);
nand U16676 (N_16676,N_15162,N_14871);
nor U16677 (N_16677,N_15361,N_14448);
nand U16678 (N_16678,N_14708,N_14780);
nor U16679 (N_16679,N_15458,N_15233);
and U16680 (N_16680,N_15338,N_15468);
nand U16681 (N_16681,N_14659,N_14588);
nor U16682 (N_16682,N_15594,N_14513);
and U16683 (N_16683,N_14450,N_15024);
nor U16684 (N_16684,N_15331,N_15452);
xnor U16685 (N_16685,N_14777,N_14821);
and U16686 (N_16686,N_14463,N_14555);
nand U16687 (N_16687,N_14621,N_14608);
xor U16688 (N_16688,N_14420,N_14614);
or U16689 (N_16689,N_14650,N_14595);
nor U16690 (N_16690,N_15482,N_14638);
nand U16691 (N_16691,N_15449,N_14458);
nand U16692 (N_16692,N_15302,N_15028);
or U16693 (N_16693,N_15396,N_15541);
and U16694 (N_16694,N_15193,N_15460);
or U16695 (N_16695,N_15454,N_14783);
nand U16696 (N_16696,N_14716,N_14734);
nor U16697 (N_16697,N_14823,N_15285);
nand U16698 (N_16698,N_15238,N_14409);
nor U16699 (N_16699,N_14646,N_15357);
and U16700 (N_16700,N_15147,N_14600);
or U16701 (N_16701,N_15424,N_14850);
nor U16702 (N_16702,N_14861,N_14740);
and U16703 (N_16703,N_14496,N_15131);
nor U16704 (N_16704,N_15430,N_15350);
and U16705 (N_16705,N_15320,N_15139);
nor U16706 (N_16706,N_14876,N_15338);
xnor U16707 (N_16707,N_14928,N_15472);
nand U16708 (N_16708,N_14857,N_14714);
xnor U16709 (N_16709,N_14406,N_15484);
and U16710 (N_16710,N_14849,N_15246);
or U16711 (N_16711,N_14435,N_15410);
and U16712 (N_16712,N_14436,N_15576);
and U16713 (N_16713,N_15500,N_14873);
xnor U16714 (N_16714,N_14931,N_14422);
or U16715 (N_16715,N_14988,N_15527);
and U16716 (N_16716,N_15561,N_14916);
nand U16717 (N_16717,N_15546,N_14546);
xnor U16718 (N_16718,N_15361,N_15171);
and U16719 (N_16719,N_15473,N_15354);
or U16720 (N_16720,N_15559,N_15532);
nor U16721 (N_16721,N_14983,N_14939);
xnor U16722 (N_16722,N_15162,N_14585);
or U16723 (N_16723,N_14612,N_14404);
nand U16724 (N_16724,N_14404,N_14489);
nand U16725 (N_16725,N_14760,N_14814);
and U16726 (N_16726,N_14657,N_15439);
xor U16727 (N_16727,N_15061,N_14862);
nor U16728 (N_16728,N_15098,N_14658);
nand U16729 (N_16729,N_15019,N_15403);
or U16730 (N_16730,N_15186,N_14820);
xnor U16731 (N_16731,N_14758,N_14817);
xor U16732 (N_16732,N_14486,N_14865);
or U16733 (N_16733,N_15212,N_15404);
or U16734 (N_16734,N_15419,N_15097);
nor U16735 (N_16735,N_15066,N_15249);
xor U16736 (N_16736,N_14864,N_15181);
and U16737 (N_16737,N_14535,N_14969);
or U16738 (N_16738,N_15149,N_15578);
and U16739 (N_16739,N_15323,N_15152);
or U16740 (N_16740,N_15039,N_14665);
nand U16741 (N_16741,N_14401,N_15077);
nand U16742 (N_16742,N_14524,N_14754);
nor U16743 (N_16743,N_14805,N_15220);
or U16744 (N_16744,N_15184,N_15207);
nor U16745 (N_16745,N_14718,N_15434);
xor U16746 (N_16746,N_14455,N_14970);
nor U16747 (N_16747,N_14425,N_15452);
and U16748 (N_16748,N_14405,N_14794);
or U16749 (N_16749,N_14713,N_15176);
xor U16750 (N_16750,N_14769,N_15330);
xnor U16751 (N_16751,N_14441,N_15465);
xor U16752 (N_16752,N_15067,N_14814);
and U16753 (N_16753,N_14748,N_14586);
or U16754 (N_16754,N_15247,N_14809);
xor U16755 (N_16755,N_14887,N_14460);
nand U16756 (N_16756,N_14783,N_15126);
nor U16757 (N_16757,N_15486,N_14569);
nand U16758 (N_16758,N_15144,N_14527);
nor U16759 (N_16759,N_14438,N_14792);
xor U16760 (N_16760,N_15305,N_14430);
nand U16761 (N_16761,N_15303,N_15164);
or U16762 (N_16762,N_15516,N_15381);
xnor U16763 (N_16763,N_14497,N_14438);
xnor U16764 (N_16764,N_14696,N_14655);
and U16765 (N_16765,N_14528,N_14436);
and U16766 (N_16766,N_14452,N_15009);
nand U16767 (N_16767,N_14514,N_14951);
xnor U16768 (N_16768,N_14687,N_15270);
nor U16769 (N_16769,N_15011,N_14818);
xor U16770 (N_16770,N_14851,N_14508);
and U16771 (N_16771,N_14936,N_14534);
and U16772 (N_16772,N_14957,N_14862);
xnor U16773 (N_16773,N_15001,N_14491);
xor U16774 (N_16774,N_14979,N_14830);
nor U16775 (N_16775,N_14649,N_15207);
xor U16776 (N_16776,N_15311,N_14459);
nor U16777 (N_16777,N_14866,N_14525);
xor U16778 (N_16778,N_14810,N_14519);
xnor U16779 (N_16779,N_15132,N_15186);
nor U16780 (N_16780,N_14986,N_15175);
and U16781 (N_16781,N_14558,N_14748);
xnor U16782 (N_16782,N_14782,N_14632);
or U16783 (N_16783,N_15287,N_14679);
and U16784 (N_16784,N_15207,N_14754);
nand U16785 (N_16785,N_14795,N_15107);
xor U16786 (N_16786,N_15571,N_15453);
and U16787 (N_16787,N_15420,N_15599);
nand U16788 (N_16788,N_15369,N_15392);
and U16789 (N_16789,N_14471,N_14938);
nand U16790 (N_16790,N_14863,N_14748);
nand U16791 (N_16791,N_15486,N_14702);
nor U16792 (N_16792,N_15160,N_14723);
or U16793 (N_16793,N_14670,N_15380);
and U16794 (N_16794,N_14853,N_15444);
or U16795 (N_16795,N_14753,N_14587);
nor U16796 (N_16796,N_14886,N_15084);
or U16797 (N_16797,N_15033,N_14722);
xnor U16798 (N_16798,N_14804,N_14922);
nand U16799 (N_16799,N_15335,N_14746);
and U16800 (N_16800,N_15817,N_15789);
or U16801 (N_16801,N_15685,N_16554);
nand U16802 (N_16802,N_15998,N_15719);
xor U16803 (N_16803,N_15938,N_15637);
nand U16804 (N_16804,N_16207,N_15921);
or U16805 (N_16805,N_15820,N_15754);
and U16806 (N_16806,N_15923,N_16672);
nand U16807 (N_16807,N_16665,N_16799);
and U16808 (N_16808,N_16736,N_15623);
nand U16809 (N_16809,N_15641,N_15629);
nor U16810 (N_16810,N_16788,N_15744);
nand U16811 (N_16811,N_15759,N_16668);
xnor U16812 (N_16812,N_16352,N_16447);
nand U16813 (N_16813,N_16408,N_16413);
or U16814 (N_16814,N_16473,N_15811);
xor U16815 (N_16815,N_16085,N_15720);
nor U16816 (N_16816,N_16164,N_16055);
nand U16817 (N_16817,N_16224,N_15781);
xnor U16818 (N_16818,N_16083,N_16195);
and U16819 (N_16819,N_16200,N_15922);
and U16820 (N_16820,N_16300,N_16429);
nand U16821 (N_16821,N_16093,N_16574);
and U16822 (N_16822,N_16534,N_15813);
nand U16823 (N_16823,N_15612,N_16040);
and U16824 (N_16824,N_16761,N_15855);
nor U16825 (N_16825,N_16231,N_15653);
xor U16826 (N_16826,N_16734,N_16148);
nand U16827 (N_16827,N_15925,N_16637);
or U16828 (N_16828,N_15770,N_16094);
and U16829 (N_16829,N_15906,N_15687);
and U16830 (N_16830,N_16233,N_15694);
xor U16831 (N_16831,N_16054,N_15668);
nor U16832 (N_16832,N_15859,N_15965);
nand U16833 (N_16833,N_16732,N_15627);
or U16834 (N_16834,N_16489,N_16517);
or U16835 (N_16835,N_15725,N_16620);
or U16836 (N_16836,N_15871,N_16718);
or U16837 (N_16837,N_15600,N_16425);
nand U16838 (N_16838,N_16560,N_15778);
nand U16839 (N_16839,N_16267,N_16174);
xor U16840 (N_16840,N_16452,N_16492);
and U16841 (N_16841,N_16405,N_16333);
nor U16842 (N_16842,N_16623,N_16027);
or U16843 (N_16843,N_16307,N_16302);
xnor U16844 (N_16844,N_16442,N_15702);
nor U16845 (N_16845,N_16234,N_15904);
xor U16846 (N_16846,N_16343,N_16645);
nor U16847 (N_16847,N_16721,N_15837);
and U16848 (N_16848,N_16244,N_16380);
nor U16849 (N_16849,N_15706,N_15800);
or U16850 (N_16850,N_16357,N_15870);
nor U16851 (N_16851,N_16003,N_15776);
and U16852 (N_16852,N_16203,N_16256);
nor U16853 (N_16853,N_15667,N_16689);
or U16854 (N_16854,N_16419,N_16169);
nand U16855 (N_16855,N_16043,N_15948);
xor U16856 (N_16856,N_15967,N_16258);
nand U16857 (N_16857,N_15768,N_16015);
nor U16858 (N_16858,N_16118,N_16313);
or U16859 (N_16859,N_16596,N_16061);
nor U16860 (N_16860,N_16626,N_16284);
nand U16861 (N_16861,N_16296,N_16058);
and U16862 (N_16862,N_16167,N_16650);
xor U16863 (N_16863,N_15609,N_16124);
nand U16864 (N_16864,N_15951,N_16250);
xor U16865 (N_16865,N_16056,N_16099);
xnor U16866 (N_16866,N_16774,N_16475);
or U16867 (N_16867,N_16340,N_15635);
and U16868 (N_16868,N_16392,N_15894);
or U16869 (N_16869,N_15712,N_16023);
nor U16870 (N_16870,N_16433,N_16444);
nand U16871 (N_16871,N_16342,N_15836);
nand U16872 (N_16872,N_15830,N_16711);
xor U16873 (N_16873,N_16611,N_15735);
or U16874 (N_16874,N_16314,N_15815);
nor U16875 (N_16875,N_16485,N_16230);
nand U16876 (N_16876,N_16019,N_15673);
and U16877 (N_16877,N_16555,N_16745);
or U16878 (N_16878,N_16441,N_16563);
or U16879 (N_16879,N_16630,N_16335);
and U16880 (N_16880,N_16037,N_16079);
nor U16881 (N_16881,N_15850,N_16614);
nor U16882 (N_16882,N_15677,N_16101);
or U16883 (N_16883,N_15785,N_15994);
and U16884 (N_16884,N_16599,N_15752);
or U16885 (N_16885,N_16683,N_15821);
xor U16886 (N_16886,N_16483,N_16422);
or U16887 (N_16887,N_15734,N_15606);
or U16888 (N_16888,N_16190,N_15617);
and U16889 (N_16889,N_15903,N_16038);
nor U16890 (N_16890,N_16400,N_16225);
and U16891 (N_16891,N_16321,N_16359);
xor U16892 (N_16892,N_16798,N_16782);
or U16893 (N_16893,N_16382,N_16308);
xnor U16894 (N_16894,N_16778,N_16561);
xor U16895 (N_16895,N_16468,N_16522);
or U16896 (N_16896,N_16281,N_16744);
nor U16897 (N_16897,N_16295,N_16748);
nand U16898 (N_16898,N_16715,N_15795);
nor U16899 (N_16899,N_15611,N_16185);
or U16900 (N_16900,N_16417,N_16770);
xor U16901 (N_16901,N_15895,N_16679);
and U16902 (N_16902,N_16292,N_16609);
nor U16903 (N_16903,N_16202,N_16116);
or U16904 (N_16904,N_15805,N_16605);
or U16905 (N_16905,N_16445,N_15680);
xor U16906 (N_16906,N_15711,N_16407);
xnor U16907 (N_16907,N_16133,N_16552);
nand U16908 (N_16908,N_16199,N_16198);
and U16909 (N_16909,N_16348,N_16228);
and U16910 (N_16910,N_15783,N_16414);
and U16911 (N_16911,N_15639,N_16653);
and U16912 (N_16912,N_16384,N_16182);
or U16913 (N_16913,N_15981,N_16050);
xnor U16914 (N_16914,N_16081,N_16304);
xor U16915 (N_16915,N_15970,N_15832);
or U16916 (N_16916,N_16006,N_15630);
nand U16917 (N_16917,N_16379,N_16676);
and U16918 (N_16918,N_16151,N_15898);
and U16919 (N_16919,N_16719,N_16480);
or U16920 (N_16920,N_16510,N_15896);
and U16921 (N_16921,N_16593,N_16428);
nor U16922 (N_16922,N_16353,N_16360);
and U16923 (N_16923,N_15890,N_15780);
nand U16924 (N_16924,N_16212,N_16642);
nor U16925 (N_16925,N_15900,N_16471);
xnor U16926 (N_16926,N_16502,N_16113);
and U16927 (N_16927,N_16294,N_16288);
xnor U16928 (N_16928,N_15941,N_16712);
nand U16929 (N_16929,N_16699,N_16354);
xnor U16930 (N_16930,N_15721,N_15853);
xnor U16931 (N_16931,N_15714,N_15621);
xor U16932 (N_16932,N_16646,N_15717);
and U16933 (N_16933,N_16029,N_15848);
nor U16934 (N_16934,N_15866,N_16771);
xnor U16935 (N_16935,N_15786,N_16196);
and U16936 (N_16936,N_15672,N_16588);
nand U16937 (N_16937,N_16365,N_16532);
nor U16938 (N_16938,N_15634,N_15675);
nand U16939 (N_16939,N_15899,N_16168);
nand U16940 (N_16940,N_16063,N_16070);
and U16941 (N_16941,N_16001,N_16479);
xnor U16942 (N_16942,N_15852,N_16240);
or U16943 (N_16943,N_16418,N_16613);
or U16944 (N_16944,N_15885,N_16740);
xor U16945 (N_16945,N_16498,N_15860);
nor U16946 (N_16946,N_16166,N_16438);
or U16947 (N_16947,N_16410,N_16443);
xnor U16948 (N_16948,N_16172,N_16355);
nor U16949 (N_16949,N_16252,N_15701);
xnor U16950 (N_16950,N_16635,N_16406);
nand U16951 (N_16951,N_16536,N_15681);
nor U16952 (N_16952,N_15933,N_16533);
nand U16953 (N_16953,N_16135,N_16312);
nor U16954 (N_16954,N_16482,N_16493);
xor U16955 (N_16955,N_15788,N_15695);
xnor U16956 (N_16956,N_15757,N_16477);
nand U16957 (N_16957,N_16173,N_16681);
and U16958 (N_16958,N_16104,N_15937);
nand U16959 (N_16959,N_16797,N_15690);
and U16960 (N_16960,N_15882,N_16045);
or U16961 (N_16961,N_15908,N_16499);
xnor U16962 (N_16962,N_15716,N_15819);
xor U16963 (N_16963,N_15743,N_16092);
nor U16964 (N_16964,N_16161,N_16470);
nor U16965 (N_16965,N_16076,N_16235);
nor U16966 (N_16966,N_16602,N_16159);
xnor U16967 (N_16967,N_15935,N_15699);
nand U16968 (N_16968,N_15608,N_16507);
nand U16969 (N_16969,N_16634,N_16690);
xnor U16970 (N_16970,N_16729,N_15990);
nor U16971 (N_16971,N_16165,N_15912);
or U16972 (N_16972,N_16180,N_15614);
nor U16973 (N_16973,N_15671,N_16263);
or U16974 (N_16974,N_16520,N_16000);
nand U16975 (N_16975,N_16759,N_16286);
and U16976 (N_16976,N_15825,N_16097);
nand U16977 (N_16977,N_15814,N_15909);
nand U16978 (N_16978,N_15968,N_15652);
nand U16979 (N_16979,N_16285,N_16440);
nand U16980 (N_16980,N_16649,N_16559);
xnor U16981 (N_16981,N_16432,N_15802);
xnor U16982 (N_16982,N_15983,N_15979);
nor U16983 (N_16983,N_15644,N_16578);
xor U16984 (N_16984,N_16030,N_15794);
nor U16985 (N_16985,N_16059,N_15982);
nor U16986 (N_16986,N_16463,N_15868);
nand U16987 (N_16987,N_16330,N_16108);
nor U16988 (N_16988,N_16742,N_16792);
nand U16989 (N_16989,N_16717,N_15897);
or U16990 (N_16990,N_15741,N_15834);
xor U16991 (N_16991,N_15625,N_15801);
nor U16992 (N_16992,N_16261,N_16455);
nor U16993 (N_16993,N_16299,N_16666);
or U16994 (N_16994,N_16075,N_15881);
and U16995 (N_16995,N_16171,N_16550);
xnor U16996 (N_16996,N_16591,N_15707);
nand U16997 (N_16997,N_15700,N_15989);
or U16998 (N_16998,N_16458,N_16476);
nand U16999 (N_16999,N_15993,N_15964);
and U17000 (N_17000,N_16631,N_16089);
and U17001 (N_17001,N_15915,N_16389);
nand U17002 (N_17002,N_16052,N_16727);
xor U17003 (N_17003,N_16607,N_16095);
nor U17004 (N_17004,N_16325,N_15732);
and U17005 (N_17005,N_16277,N_15656);
and U17006 (N_17006,N_16763,N_16098);
xnor U17007 (N_17007,N_15976,N_15650);
xor U17008 (N_17008,N_16714,N_15618);
nor U17009 (N_17009,N_16018,N_16724);
nor U17010 (N_17010,N_16518,N_16786);
or U17011 (N_17011,N_15746,N_15664);
xnor U17012 (N_17012,N_15958,N_15854);
xor U17013 (N_17013,N_16460,N_15601);
xor U17014 (N_17014,N_15946,N_16112);
nand U17015 (N_17015,N_15874,N_15875);
nor U17016 (N_17016,N_15843,N_16746);
nand U17017 (N_17017,N_15987,N_15683);
and U17018 (N_17018,N_16011,N_16377);
or U17019 (N_17019,N_15772,N_16239);
nand U17020 (N_17020,N_15957,N_15791);
and U17021 (N_17021,N_15808,N_16680);
nand U17022 (N_17022,N_16741,N_16752);
nor U17023 (N_17023,N_16287,N_15978);
or U17024 (N_17024,N_16396,N_15771);
xnor U17025 (N_17025,N_16695,N_15901);
xor U17026 (N_17026,N_16504,N_16386);
xnor U17027 (N_17027,N_16765,N_16109);
xor U17028 (N_17028,N_16531,N_15709);
and U17029 (N_17029,N_16696,N_15997);
xor U17030 (N_17030,N_16328,N_15610);
nand U17031 (N_17031,N_15659,N_16192);
nand U17032 (N_17032,N_16662,N_16211);
nand U17033 (N_17033,N_16659,N_16539);
and U17034 (N_17034,N_15844,N_16339);
nand U17035 (N_17035,N_16290,N_15628);
nor U17036 (N_17036,N_16158,N_16776);
nand U17037 (N_17037,N_16508,N_16412);
nor U17038 (N_17038,N_16437,N_16065);
and U17039 (N_17039,N_16457,N_15750);
nand U17040 (N_17040,N_16692,N_16454);
nand U17041 (N_17041,N_16615,N_16436);
nor U17042 (N_17042,N_16720,N_16257);
nor U17043 (N_17043,N_16698,N_16487);
xor U17044 (N_17044,N_15742,N_16512);
and U17045 (N_17045,N_16223,N_16600);
xnor U17046 (N_17046,N_16048,N_16506);
xor U17047 (N_17047,N_16152,N_16024);
or U17048 (N_17048,N_16769,N_16648);
xor U17049 (N_17049,N_15995,N_16035);
and U17050 (N_17050,N_16728,N_16704);
nand U17051 (N_17051,N_16162,N_16570);
and U17052 (N_17052,N_16254,N_15774);
xnor U17053 (N_17053,N_16766,N_15674);
or U17054 (N_17054,N_16237,N_15991);
or U17055 (N_17055,N_16028,N_16523);
or U17056 (N_17056,N_15764,N_16515);
or U17057 (N_17057,N_16276,N_15929);
nor U17058 (N_17058,N_15782,N_16067);
and U17059 (N_17059,N_16556,N_16047);
nand U17060 (N_17060,N_15838,N_16176);
xnor U17061 (N_17061,N_16633,N_15986);
and U17062 (N_17062,N_16126,N_16305);
and U17063 (N_17063,N_16044,N_16332);
nand U17064 (N_17064,N_16669,N_16186);
nor U17065 (N_17065,N_15739,N_16383);
and U17066 (N_17066,N_16586,N_15822);
nand U17067 (N_17067,N_16587,N_15684);
or U17068 (N_17068,N_16416,N_16575);
and U17069 (N_17069,N_16639,N_16795);
and U17070 (N_17070,N_16545,N_15867);
or U17071 (N_17071,N_15797,N_15698);
or U17072 (N_17072,N_15841,N_16465);
and U17073 (N_17073,N_15691,N_16751);
and U17074 (N_17074,N_15793,N_16255);
nand U17075 (N_17075,N_15930,N_16638);
nor U17076 (N_17076,N_16145,N_16005);
xor U17077 (N_17077,N_16528,N_15977);
or U17078 (N_17078,N_16137,N_16686);
and U17079 (N_17079,N_16731,N_16282);
and U17080 (N_17080,N_16459,N_16421);
nor U17081 (N_17081,N_16178,N_16260);
nor U17082 (N_17082,N_16664,N_16289);
xor U17083 (N_17083,N_15773,N_16007);
nand U17084 (N_17084,N_15931,N_16147);
nand U17085 (N_17085,N_15758,N_15862);
or U17086 (N_17086,N_16341,N_16146);
xnor U17087 (N_17087,N_16114,N_16391);
nor U17088 (N_17088,N_16326,N_16411);
and U17089 (N_17089,N_16709,N_16086);
or U17090 (N_17090,N_16657,N_16371);
xnor U17091 (N_17091,N_15718,N_16791);
or U17092 (N_17092,N_15737,N_15902);
xnor U17093 (N_17093,N_16706,N_16567);
nor U17094 (N_17094,N_15810,N_15613);
and U17095 (N_17095,N_15662,N_16363);
or U17096 (N_17096,N_16478,N_16245);
nand U17097 (N_17097,N_15665,N_16356);
and U17098 (N_17098,N_16395,N_16042);
nor U17099 (N_17099,N_16119,N_16236);
nor U17100 (N_17100,N_16549,N_15682);
nor U17101 (N_17101,N_16541,N_16542);
nor U17102 (N_17102,N_15777,N_16625);
xor U17103 (N_17103,N_15956,N_15666);
xnor U17104 (N_17104,N_15911,N_16214);
and U17105 (N_17105,N_15910,N_15869);
nand U17106 (N_17106,N_16129,N_15858);
xnor U17107 (N_17107,N_16793,N_16265);
xnor U17108 (N_17108,N_15705,N_16713);
xnor U17109 (N_17109,N_16311,N_16163);
nor U17110 (N_17110,N_16381,N_16540);
nand U17111 (N_17111,N_16322,N_15926);
and U17112 (N_17112,N_16025,N_16547);
nand U17113 (N_17113,N_15604,N_16138);
and U17114 (N_17114,N_15944,N_16481);
xor U17115 (N_17115,N_16450,N_16553);
xnor U17116 (N_17116,N_16544,N_16346);
nor U17117 (N_17117,N_15887,N_16582);
nor U17118 (N_17118,N_16057,N_16269);
or U17119 (N_17119,N_15745,N_16122);
xnor U17120 (N_17120,N_15864,N_15823);
or U17121 (N_17121,N_16082,N_16026);
and U17122 (N_17122,N_16039,N_15607);
nand U17123 (N_17123,N_16601,N_16010);
nand U17124 (N_17124,N_16674,N_16175);
and U17125 (N_17125,N_16197,N_16394);
nor U17126 (N_17126,N_15729,N_15704);
nand U17127 (N_17127,N_16643,N_16273);
or U17128 (N_17128,N_15829,N_16621);
and U17129 (N_17129,N_16297,N_16426);
and U17130 (N_17130,N_15715,N_15688);
xor U17131 (N_17131,N_16521,N_16703);
or U17132 (N_17132,N_16682,N_16446);
nand U17133 (N_17133,N_16364,N_16266);
and U17134 (N_17134,N_16397,N_16415);
nor U17135 (N_17135,N_16678,N_16758);
or U17136 (N_17136,N_15605,N_16608);
xor U17137 (N_17137,N_16739,N_16590);
nand U17138 (N_17138,N_15846,N_15703);
nand U17139 (N_17139,N_15723,N_16527);
nor U17140 (N_17140,N_16157,N_16191);
and U17141 (N_17141,N_16624,N_16110);
nor U17142 (N_17142,N_15766,N_15886);
or U17143 (N_17143,N_16456,N_16577);
nand U17144 (N_17144,N_16697,N_16738);
and U17145 (N_17145,N_16153,N_16249);
xor U17146 (N_17146,N_16217,N_16209);
nor U17147 (N_17147,N_15996,N_16309);
and U17148 (N_17148,N_16768,N_15818);
and U17149 (N_17149,N_16338,N_15943);
xor U17150 (N_17150,N_15863,N_16501);
or U17151 (N_17151,N_16324,N_16336);
nand U17152 (N_17152,N_15924,N_16494);
nor U17153 (N_17153,N_15660,N_16262);
nor U17154 (N_17154,N_16500,N_15812);
xnor U17155 (N_17155,N_16726,N_15733);
or U17156 (N_17156,N_15669,N_15927);
xor U17157 (N_17157,N_15692,N_16617);
nand U17158 (N_17158,N_16275,N_16107);
or U17159 (N_17159,N_15952,N_15816);
xnor U17160 (N_17160,N_16194,N_16131);
nand U17161 (N_17161,N_16790,N_15615);
nand U17162 (N_17162,N_16671,N_15809);
or U17163 (N_17163,N_16663,N_16378);
and U17164 (N_17164,N_16072,N_16767);
xnor U17165 (N_17165,N_16573,N_15792);
and U17166 (N_17166,N_16210,N_16078);
and U17167 (N_17167,N_16090,N_15796);
and U17168 (N_17168,N_16017,N_15747);
nand U17169 (N_17169,N_16616,N_16700);
and U17170 (N_17170,N_16051,N_16448);
or U17171 (N_17171,N_15697,N_16362);
nor U17172 (N_17172,N_16760,N_16337);
xnor U17173 (N_17173,N_16246,N_16369);
nor U17174 (N_17174,N_16451,N_15616);
or U17175 (N_17175,N_16497,N_15648);
and U17176 (N_17176,N_16347,N_16772);
nand U17177 (N_17177,N_15765,N_15972);
and U17178 (N_17178,N_16431,N_15831);
and U17179 (N_17179,N_16495,N_16142);
and U17180 (N_17180,N_16598,N_16318);
and U17181 (N_17181,N_15955,N_16543);
xnor U17182 (N_17182,N_15636,N_16677);
or U17183 (N_17183,N_15973,N_16002);
nand U17184 (N_17184,N_15678,N_16610);
xnor U17185 (N_17185,N_15856,N_16647);
nand U17186 (N_17186,N_15646,N_16096);
nand U17187 (N_17187,N_15798,N_16794);
xnor U17188 (N_17188,N_16319,N_16579);
nand U17189 (N_17189,N_16773,N_16566);
xnor U17190 (N_17190,N_16514,N_16215);
xnor U17191 (N_17191,N_16221,N_15932);
xor U17192 (N_17192,N_16144,N_16705);
or U17193 (N_17193,N_15693,N_16537);
xnor U17194 (N_17194,N_16399,N_15872);
nor U17195 (N_17195,N_16509,N_16062);
xor U17196 (N_17196,N_16466,N_16141);
nand U17197 (N_17197,N_15649,N_16177);
nand U17198 (N_17198,N_16667,N_16316);
and U17199 (N_17199,N_16461,N_16701);
and U17200 (N_17200,N_15827,N_16708);
nor U17201 (N_17201,N_15961,N_16184);
nor U17202 (N_17202,N_16564,N_16125);
or U17203 (N_17203,N_16551,N_16684);
or U17204 (N_17204,N_15824,N_16583);
and U17205 (N_17205,N_15845,N_16021);
and U17206 (N_17206,N_16012,N_15661);
nor U17207 (N_17207,N_15891,N_16427);
nand U17208 (N_17208,N_16375,N_15857);
nor U17209 (N_17209,N_15738,N_16117);
and U17210 (N_17210,N_16688,N_16320);
nor U17211 (N_17211,N_16423,N_16462);
nor U17212 (N_17212,N_15945,N_16120);
nor U17213 (N_17213,N_16503,N_16298);
and U17214 (N_17214,N_16796,N_16248);
nor U17215 (N_17215,N_16034,N_15751);
nand U17216 (N_17216,N_16376,N_15727);
xor U17217 (N_17217,N_16612,N_15835);
nand U17218 (N_17218,N_16439,N_16361);
nor U17219 (N_17219,N_16247,N_15631);
nor U17220 (N_17220,N_15876,N_16603);
nor U17221 (N_17221,N_15960,N_16123);
or U17222 (N_17222,N_16130,N_15992);
and U17223 (N_17223,N_16291,N_16519);
or U17224 (N_17224,N_16513,N_16474);
nor U17225 (N_17225,N_16764,N_16754);
or U17226 (N_17226,N_16747,N_16218);
nor U17227 (N_17227,N_15626,N_16576);
nor U17228 (N_17228,N_15740,N_16505);
xor U17229 (N_17229,N_15971,N_15767);
and U17230 (N_17230,N_16393,N_16031);
nor U17231 (N_17231,N_16403,N_16208);
xor U17232 (N_17232,N_15663,N_16486);
nor U17233 (N_17233,N_16229,N_16716);
xnor U17234 (N_17234,N_15839,N_16750);
xnor U17235 (N_17235,N_16660,N_16402);
xnor U17236 (N_17236,N_15645,N_16735);
nor U17237 (N_17237,N_16449,N_16629);
or U17238 (N_17238,N_15748,N_16074);
and U17239 (N_17239,N_15934,N_16004);
and U17240 (N_17240,N_15713,N_15784);
nand U17241 (N_17241,N_16160,N_15710);
or U17242 (N_17242,N_16488,N_15657);
nor U17243 (N_17243,N_16526,N_15947);
nor U17244 (N_17244,N_16193,N_16585);
and U17245 (N_17245,N_16226,N_15679);
and U17246 (N_17246,N_16032,N_16756);
xnor U17247 (N_17247,N_16641,N_16222);
nor U17248 (N_17248,N_15884,N_15787);
and U17249 (N_17249,N_16757,N_16087);
nand U17250 (N_17250,N_16737,N_16604);
nand U17251 (N_17251,N_16775,N_16580);
and U17252 (N_17252,N_16344,N_16187);
or U17253 (N_17253,N_16565,N_16132);
xor U17254 (N_17254,N_15879,N_15651);
or U17255 (N_17255,N_16420,N_15779);
nor U17256 (N_17256,N_16385,N_16350);
nand U17257 (N_17257,N_16524,N_16189);
nor U17258 (N_17258,N_16306,N_15883);
xnor U17259 (N_17259,N_15936,N_15962);
and U17260 (N_17260,N_16636,N_16430);
and U17261 (N_17261,N_16644,N_16278);
nand U17262 (N_17262,N_15756,N_16069);
nand U17263 (N_17263,N_16216,N_16068);
nand U17264 (N_17264,N_16219,N_16315);
nor U17265 (N_17265,N_16435,N_15963);
nand U17266 (N_17266,N_16009,N_16694);
nor U17267 (N_17267,N_16049,N_15975);
nor U17268 (N_17268,N_15755,N_16743);
nor U17269 (N_17269,N_15966,N_15919);
or U17270 (N_17270,N_16755,N_15833);
nor U17271 (N_17271,N_16388,N_16651);
or U17272 (N_17272,N_15893,N_16722);
or U17273 (N_17273,N_15762,N_16789);
nor U17274 (N_17274,N_15670,N_16253);
xor U17275 (N_17275,N_16139,N_16584);
or U17276 (N_17276,N_15622,N_16293);
xor U17277 (N_17277,N_15953,N_15775);
nand U17278 (N_17278,N_15799,N_16673);
and U17279 (N_17279,N_16149,N_16241);
or U17280 (N_17280,N_16170,N_15658);
and U17281 (N_17281,N_15632,N_16100);
nand U17282 (N_17282,N_16535,N_16453);
or U17283 (N_17283,N_15696,N_15847);
or U17284 (N_17284,N_15760,N_15803);
xor U17285 (N_17285,N_15728,N_15840);
or U17286 (N_17286,N_16374,N_15914);
xnor U17287 (N_17287,N_16490,N_16205);
and U17288 (N_17288,N_16548,N_16053);
and U17289 (N_17289,N_16781,N_16546);
xor U17290 (N_17290,N_15731,N_15918);
nand U17291 (N_17291,N_16730,N_15726);
nor U17292 (N_17292,N_16390,N_16589);
nand U17293 (N_17293,N_16538,N_16370);
or U17294 (N_17294,N_16401,N_15655);
nor U17295 (N_17295,N_16105,N_16264);
nor U17296 (N_17296,N_16329,N_16283);
nand U17297 (N_17297,N_16143,N_16317);
nor U17298 (N_17298,N_16127,N_15753);
nand U17299 (N_17299,N_15638,N_16301);
and U17300 (N_17300,N_15602,N_16484);
and U17301 (N_17301,N_16310,N_15877);
nor U17302 (N_17302,N_16594,N_16562);
nand U17303 (N_17303,N_16424,N_15603);
nor U17304 (N_17304,N_16749,N_16622);
or U17305 (N_17305,N_15769,N_15880);
nand U17306 (N_17306,N_16372,N_16206);
or U17307 (N_17307,N_16787,N_15633);
and U17308 (N_17308,N_15969,N_16077);
or U17309 (N_17309,N_16592,N_15790);
nor U17310 (N_17310,N_16345,N_15878);
and U17311 (N_17311,N_16785,N_16060);
xnor U17312 (N_17312,N_16777,N_16183);
and U17313 (N_17313,N_16073,N_15942);
xnor U17314 (N_17314,N_16707,N_16103);
xor U17315 (N_17315,N_15804,N_16762);
xnor U17316 (N_17316,N_16046,N_16387);
or U17317 (N_17317,N_16581,N_16274);
or U17318 (N_17318,N_16628,N_15730);
nor U17319 (N_17319,N_15959,N_16111);
xnor U17320 (N_17320,N_15928,N_15892);
nand U17321 (N_17321,N_15954,N_16213);
and U17322 (N_17322,N_15676,N_16136);
or U17323 (N_17323,N_16597,N_15722);
nand U17324 (N_17324,N_15939,N_16702);
xor U17325 (N_17325,N_15807,N_15985);
nor U17326 (N_17326,N_16268,N_15916);
and U17327 (N_17327,N_16102,N_16154);
nor U17328 (N_17328,N_16618,N_16572);
xor U17329 (N_17329,N_15624,N_16525);
nor U17330 (N_17330,N_16693,N_16238);
nand U17331 (N_17331,N_16367,N_16529);
xor U17332 (N_17332,N_16279,N_15888);
or U17333 (N_17333,N_16179,N_16656);
nand U17334 (N_17334,N_15724,N_15749);
nor U17335 (N_17335,N_16733,N_16409);
xor U17336 (N_17336,N_16654,N_16008);
and U17337 (N_17337,N_16632,N_15920);
nand U17338 (N_17338,N_15984,N_16084);
nand U17339 (N_17339,N_16155,N_15907);
or U17340 (N_17340,N_16349,N_16464);
and U17341 (N_17341,N_16569,N_16251);
nand U17342 (N_17342,N_16134,N_16036);
nor U17343 (N_17343,N_16516,N_16181);
and U17344 (N_17344,N_16652,N_16472);
and U17345 (N_17345,N_15736,N_15686);
xnor U17346 (N_17346,N_16398,N_16627);
nor U17347 (N_17347,N_16150,N_15826);
nand U17348 (N_17348,N_16270,N_15974);
nor U17349 (N_17349,N_16220,N_16691);
and U17350 (N_17350,N_16753,N_15949);
or U17351 (N_17351,N_16358,N_16725);
and U17352 (N_17352,N_16280,N_15763);
xor U17353 (N_17353,N_15654,N_15849);
and U17354 (N_17354,N_15828,N_16779);
or U17355 (N_17355,N_16303,N_15913);
xor U17356 (N_17356,N_16723,N_16351);
nor U17357 (N_17357,N_16373,N_15917);
and U17358 (N_17358,N_16571,N_16115);
and U17359 (N_17359,N_16156,N_16121);
nand U17360 (N_17360,N_16404,N_16511);
xnor U17361 (N_17361,N_16467,N_16366);
and U17362 (N_17362,N_16655,N_15865);
and U17363 (N_17363,N_16064,N_16658);
nand U17364 (N_17364,N_16201,N_16323);
nor U17365 (N_17365,N_16368,N_16661);
or U17366 (N_17366,N_16595,N_15988);
and U17367 (N_17367,N_16242,N_16232);
and U17368 (N_17368,N_16619,N_16071);
or U17369 (N_17369,N_16685,N_16227);
nand U17370 (N_17370,N_15940,N_16013);
and U17371 (N_17371,N_16530,N_16334);
xnor U17372 (N_17372,N_15689,N_16080);
and U17373 (N_17373,N_15620,N_16491);
and U17374 (N_17374,N_16020,N_16033);
and U17375 (N_17375,N_16243,N_15861);
xor U17376 (N_17376,N_15980,N_16204);
nand U17377 (N_17377,N_16557,N_15950);
xor U17378 (N_17378,N_16188,N_15761);
and U17379 (N_17379,N_16106,N_16568);
and U17380 (N_17380,N_16558,N_15889);
nand U17381 (N_17381,N_15640,N_15806);
xnor U17382 (N_17382,N_16469,N_16606);
xor U17383 (N_17383,N_16088,N_16014);
or U17384 (N_17384,N_15851,N_15647);
nand U17385 (N_17385,N_16272,N_16259);
xnor U17386 (N_17386,N_16783,N_16041);
xor U17387 (N_17387,N_15619,N_16687);
nand U17388 (N_17388,N_16710,N_16327);
nand U17389 (N_17389,N_15708,N_16675);
or U17390 (N_17390,N_16331,N_16780);
xor U17391 (N_17391,N_16128,N_15873);
nand U17392 (N_17392,N_15999,N_15842);
xor U17393 (N_17393,N_16016,N_15905);
nand U17394 (N_17394,N_16784,N_16271);
nand U17395 (N_17395,N_16022,N_16091);
or U17396 (N_17396,N_16496,N_15643);
xnor U17397 (N_17397,N_16434,N_16066);
xor U17398 (N_17398,N_16640,N_16140);
xor U17399 (N_17399,N_15642,N_16670);
or U17400 (N_17400,N_16534,N_16008);
and U17401 (N_17401,N_16759,N_16294);
xnor U17402 (N_17402,N_15801,N_16071);
xnor U17403 (N_17403,N_16746,N_16620);
and U17404 (N_17404,N_16444,N_16251);
and U17405 (N_17405,N_16098,N_16342);
nand U17406 (N_17406,N_15933,N_16746);
nand U17407 (N_17407,N_15902,N_16050);
or U17408 (N_17408,N_15897,N_16447);
nor U17409 (N_17409,N_15736,N_15657);
and U17410 (N_17410,N_16653,N_16487);
xnor U17411 (N_17411,N_16654,N_15794);
and U17412 (N_17412,N_16176,N_16458);
and U17413 (N_17413,N_16308,N_16273);
xnor U17414 (N_17414,N_15827,N_16535);
or U17415 (N_17415,N_15829,N_15778);
or U17416 (N_17416,N_16471,N_16698);
or U17417 (N_17417,N_16199,N_16390);
and U17418 (N_17418,N_16478,N_16343);
xnor U17419 (N_17419,N_15880,N_15801);
and U17420 (N_17420,N_16523,N_16632);
and U17421 (N_17421,N_16124,N_16324);
nand U17422 (N_17422,N_16235,N_16068);
nand U17423 (N_17423,N_15849,N_15791);
xor U17424 (N_17424,N_16019,N_15668);
nand U17425 (N_17425,N_15652,N_15708);
nand U17426 (N_17426,N_16135,N_16516);
and U17427 (N_17427,N_16588,N_15825);
nand U17428 (N_17428,N_15756,N_15728);
nand U17429 (N_17429,N_15780,N_16597);
or U17430 (N_17430,N_16560,N_15728);
nor U17431 (N_17431,N_15782,N_16060);
or U17432 (N_17432,N_15868,N_16507);
nor U17433 (N_17433,N_16380,N_16522);
xnor U17434 (N_17434,N_16099,N_15871);
xor U17435 (N_17435,N_16407,N_15757);
nor U17436 (N_17436,N_15775,N_16280);
nand U17437 (N_17437,N_15885,N_16634);
or U17438 (N_17438,N_16723,N_16763);
nand U17439 (N_17439,N_16209,N_16749);
and U17440 (N_17440,N_15932,N_15988);
and U17441 (N_17441,N_16708,N_16427);
xor U17442 (N_17442,N_16629,N_16038);
xor U17443 (N_17443,N_16001,N_16252);
nand U17444 (N_17444,N_16062,N_15797);
and U17445 (N_17445,N_16652,N_15615);
nor U17446 (N_17446,N_16611,N_15974);
nand U17447 (N_17447,N_15772,N_15899);
nand U17448 (N_17448,N_16628,N_16541);
and U17449 (N_17449,N_15922,N_16736);
nand U17450 (N_17450,N_15685,N_16255);
and U17451 (N_17451,N_16246,N_16531);
and U17452 (N_17452,N_15704,N_16635);
xor U17453 (N_17453,N_15961,N_15851);
or U17454 (N_17454,N_16535,N_16011);
or U17455 (N_17455,N_16561,N_16777);
xnor U17456 (N_17456,N_16426,N_16474);
and U17457 (N_17457,N_16751,N_15793);
nand U17458 (N_17458,N_16132,N_16131);
or U17459 (N_17459,N_15841,N_15699);
and U17460 (N_17460,N_15994,N_16074);
nand U17461 (N_17461,N_16502,N_16435);
and U17462 (N_17462,N_16793,N_15788);
and U17463 (N_17463,N_16630,N_15794);
nor U17464 (N_17464,N_15657,N_16116);
and U17465 (N_17465,N_16223,N_15922);
xor U17466 (N_17466,N_16166,N_15931);
nand U17467 (N_17467,N_15858,N_16449);
and U17468 (N_17468,N_15692,N_15908);
and U17469 (N_17469,N_16063,N_16749);
nand U17470 (N_17470,N_15793,N_16001);
nor U17471 (N_17471,N_16467,N_15612);
xnor U17472 (N_17472,N_15820,N_16044);
or U17473 (N_17473,N_16797,N_15616);
or U17474 (N_17474,N_16186,N_16194);
or U17475 (N_17475,N_15610,N_16005);
or U17476 (N_17476,N_16574,N_15978);
nand U17477 (N_17477,N_16219,N_15660);
or U17478 (N_17478,N_16610,N_15679);
or U17479 (N_17479,N_16394,N_16258);
nand U17480 (N_17480,N_15759,N_16302);
or U17481 (N_17481,N_15876,N_16272);
nand U17482 (N_17482,N_15904,N_16479);
nor U17483 (N_17483,N_16793,N_16778);
nor U17484 (N_17484,N_16023,N_16542);
or U17485 (N_17485,N_16610,N_16614);
xor U17486 (N_17486,N_16542,N_15935);
xor U17487 (N_17487,N_15667,N_16024);
xor U17488 (N_17488,N_15824,N_15902);
nand U17489 (N_17489,N_16335,N_16689);
and U17490 (N_17490,N_16313,N_16511);
or U17491 (N_17491,N_15838,N_16111);
xnor U17492 (N_17492,N_15617,N_15988);
nand U17493 (N_17493,N_15606,N_16361);
xor U17494 (N_17494,N_16420,N_16479);
nand U17495 (N_17495,N_15988,N_16307);
or U17496 (N_17496,N_15760,N_16786);
or U17497 (N_17497,N_16600,N_15710);
xor U17498 (N_17498,N_16402,N_15611);
or U17499 (N_17499,N_15811,N_16438);
xnor U17500 (N_17500,N_16113,N_16576);
and U17501 (N_17501,N_16409,N_15741);
nor U17502 (N_17502,N_16561,N_16596);
xor U17503 (N_17503,N_16580,N_15901);
or U17504 (N_17504,N_16088,N_15991);
nand U17505 (N_17505,N_16259,N_16049);
nor U17506 (N_17506,N_16419,N_16027);
nor U17507 (N_17507,N_16499,N_16175);
and U17508 (N_17508,N_15794,N_16615);
nand U17509 (N_17509,N_16314,N_15630);
nand U17510 (N_17510,N_16440,N_16493);
nor U17511 (N_17511,N_16404,N_16044);
nand U17512 (N_17512,N_16454,N_16428);
nor U17513 (N_17513,N_16311,N_15920);
or U17514 (N_17514,N_16174,N_16145);
or U17515 (N_17515,N_16773,N_16253);
and U17516 (N_17516,N_16654,N_16333);
nor U17517 (N_17517,N_15809,N_16042);
or U17518 (N_17518,N_15913,N_16297);
and U17519 (N_17519,N_15855,N_16334);
and U17520 (N_17520,N_16290,N_16044);
and U17521 (N_17521,N_15781,N_15856);
and U17522 (N_17522,N_15602,N_16643);
nor U17523 (N_17523,N_16463,N_16498);
nor U17524 (N_17524,N_16394,N_16410);
xor U17525 (N_17525,N_16540,N_16731);
xor U17526 (N_17526,N_15682,N_15612);
xnor U17527 (N_17527,N_15969,N_16212);
nand U17528 (N_17528,N_16529,N_16123);
and U17529 (N_17529,N_15651,N_15690);
or U17530 (N_17530,N_15762,N_16731);
nor U17531 (N_17531,N_16376,N_16124);
xor U17532 (N_17532,N_16124,N_16023);
and U17533 (N_17533,N_16053,N_15703);
xnor U17534 (N_17534,N_16718,N_16172);
or U17535 (N_17535,N_15994,N_16324);
or U17536 (N_17536,N_16147,N_15929);
nand U17537 (N_17537,N_16162,N_16522);
nand U17538 (N_17538,N_16496,N_16610);
and U17539 (N_17539,N_16429,N_16725);
or U17540 (N_17540,N_15967,N_16425);
xnor U17541 (N_17541,N_16769,N_16370);
xnor U17542 (N_17542,N_16607,N_16614);
or U17543 (N_17543,N_16518,N_16387);
xnor U17544 (N_17544,N_15754,N_16459);
nor U17545 (N_17545,N_16736,N_15821);
nor U17546 (N_17546,N_15957,N_15720);
xnor U17547 (N_17547,N_16130,N_16328);
or U17548 (N_17548,N_15829,N_16563);
and U17549 (N_17549,N_16138,N_16688);
xor U17550 (N_17550,N_16214,N_15791);
xnor U17551 (N_17551,N_16792,N_16451);
nor U17552 (N_17552,N_15994,N_16073);
nand U17553 (N_17553,N_16328,N_15818);
xor U17554 (N_17554,N_16480,N_16598);
nor U17555 (N_17555,N_16483,N_16271);
nor U17556 (N_17556,N_15648,N_16128);
nand U17557 (N_17557,N_16266,N_15638);
nor U17558 (N_17558,N_15621,N_15986);
or U17559 (N_17559,N_16663,N_16760);
nor U17560 (N_17560,N_16554,N_16253);
xnor U17561 (N_17561,N_16539,N_16301);
nand U17562 (N_17562,N_15727,N_16779);
and U17563 (N_17563,N_15769,N_16103);
or U17564 (N_17564,N_15665,N_16101);
xnor U17565 (N_17565,N_16406,N_16229);
or U17566 (N_17566,N_16287,N_15629);
and U17567 (N_17567,N_16100,N_16020);
or U17568 (N_17568,N_16676,N_15998);
or U17569 (N_17569,N_15904,N_16398);
or U17570 (N_17570,N_15895,N_16762);
or U17571 (N_17571,N_16756,N_16630);
nand U17572 (N_17572,N_16704,N_15844);
nand U17573 (N_17573,N_15863,N_15794);
or U17574 (N_17574,N_16661,N_15842);
xnor U17575 (N_17575,N_16482,N_16478);
and U17576 (N_17576,N_16601,N_16025);
xnor U17577 (N_17577,N_16297,N_16632);
and U17578 (N_17578,N_15871,N_15629);
or U17579 (N_17579,N_15871,N_16232);
nor U17580 (N_17580,N_16754,N_15961);
or U17581 (N_17581,N_16726,N_16380);
and U17582 (N_17582,N_15813,N_16599);
or U17583 (N_17583,N_15745,N_16562);
or U17584 (N_17584,N_15814,N_16367);
or U17585 (N_17585,N_15933,N_15874);
xnor U17586 (N_17586,N_15991,N_16155);
xor U17587 (N_17587,N_16090,N_16478);
and U17588 (N_17588,N_16603,N_15989);
nand U17589 (N_17589,N_15628,N_15998);
and U17590 (N_17590,N_16714,N_16320);
nand U17591 (N_17591,N_16195,N_15936);
xor U17592 (N_17592,N_15948,N_16113);
nand U17593 (N_17593,N_16091,N_16228);
or U17594 (N_17594,N_15913,N_16622);
xor U17595 (N_17595,N_15787,N_15692);
and U17596 (N_17596,N_16107,N_16128);
nand U17597 (N_17597,N_16032,N_15790);
xnor U17598 (N_17598,N_15890,N_15624);
or U17599 (N_17599,N_16683,N_16577);
and U17600 (N_17600,N_16678,N_16368);
nand U17601 (N_17601,N_16474,N_16467);
or U17602 (N_17602,N_15893,N_16255);
and U17603 (N_17603,N_16656,N_16264);
nand U17604 (N_17604,N_15833,N_16046);
nor U17605 (N_17605,N_16762,N_16211);
xor U17606 (N_17606,N_16579,N_15662);
nor U17607 (N_17607,N_16367,N_16791);
xor U17608 (N_17608,N_16410,N_15943);
xnor U17609 (N_17609,N_16643,N_16272);
xor U17610 (N_17610,N_16796,N_16461);
xor U17611 (N_17611,N_16238,N_15953);
nor U17612 (N_17612,N_16615,N_15661);
nor U17613 (N_17613,N_16670,N_16761);
nor U17614 (N_17614,N_16053,N_15942);
nor U17615 (N_17615,N_15691,N_16448);
and U17616 (N_17616,N_16111,N_16349);
nor U17617 (N_17617,N_16659,N_16483);
nand U17618 (N_17618,N_16599,N_16647);
or U17619 (N_17619,N_16354,N_16183);
nor U17620 (N_17620,N_16308,N_15819);
or U17621 (N_17621,N_16564,N_16094);
and U17622 (N_17622,N_15820,N_16182);
nor U17623 (N_17623,N_16382,N_15763);
nor U17624 (N_17624,N_16024,N_16063);
or U17625 (N_17625,N_16316,N_16431);
nor U17626 (N_17626,N_16405,N_15695);
nand U17627 (N_17627,N_15736,N_16148);
and U17628 (N_17628,N_16172,N_15758);
and U17629 (N_17629,N_15833,N_16588);
xor U17630 (N_17630,N_16268,N_15607);
or U17631 (N_17631,N_16025,N_16663);
xnor U17632 (N_17632,N_16651,N_15904);
and U17633 (N_17633,N_16303,N_16568);
nand U17634 (N_17634,N_15799,N_15724);
or U17635 (N_17635,N_16517,N_16327);
nor U17636 (N_17636,N_16174,N_15699);
nor U17637 (N_17637,N_16688,N_16501);
nor U17638 (N_17638,N_16758,N_16277);
xnor U17639 (N_17639,N_16357,N_15972);
xnor U17640 (N_17640,N_16157,N_15615);
xor U17641 (N_17641,N_15941,N_16525);
and U17642 (N_17642,N_16166,N_16383);
nand U17643 (N_17643,N_16175,N_16643);
or U17644 (N_17644,N_16612,N_16494);
nor U17645 (N_17645,N_16621,N_15676);
nor U17646 (N_17646,N_15858,N_15803);
or U17647 (N_17647,N_16518,N_16733);
or U17648 (N_17648,N_16739,N_16791);
or U17649 (N_17649,N_15706,N_15906);
nand U17650 (N_17650,N_15993,N_16347);
or U17651 (N_17651,N_16561,N_16094);
and U17652 (N_17652,N_16745,N_16516);
xor U17653 (N_17653,N_15740,N_16223);
or U17654 (N_17654,N_16493,N_16048);
nand U17655 (N_17655,N_16060,N_16754);
nor U17656 (N_17656,N_16029,N_16407);
and U17657 (N_17657,N_15778,N_16017);
nand U17658 (N_17658,N_15776,N_16603);
or U17659 (N_17659,N_16350,N_16792);
nand U17660 (N_17660,N_16415,N_15767);
and U17661 (N_17661,N_16049,N_16716);
and U17662 (N_17662,N_16448,N_16233);
xnor U17663 (N_17663,N_15960,N_16593);
or U17664 (N_17664,N_16342,N_15895);
or U17665 (N_17665,N_16577,N_15880);
xor U17666 (N_17666,N_16796,N_15981);
and U17667 (N_17667,N_16549,N_16338);
or U17668 (N_17668,N_16481,N_15617);
xor U17669 (N_17669,N_16133,N_15931);
and U17670 (N_17670,N_16090,N_16252);
and U17671 (N_17671,N_16116,N_16147);
nand U17672 (N_17672,N_16722,N_15881);
nand U17673 (N_17673,N_15755,N_15689);
nand U17674 (N_17674,N_15756,N_15650);
nand U17675 (N_17675,N_16663,N_16276);
nand U17676 (N_17676,N_15732,N_15774);
nor U17677 (N_17677,N_15799,N_15875);
and U17678 (N_17678,N_16021,N_16396);
nand U17679 (N_17679,N_16664,N_16629);
nand U17680 (N_17680,N_15858,N_16650);
nor U17681 (N_17681,N_16661,N_15647);
nand U17682 (N_17682,N_16720,N_16639);
and U17683 (N_17683,N_16677,N_15627);
or U17684 (N_17684,N_16782,N_16155);
or U17685 (N_17685,N_15667,N_15752);
nand U17686 (N_17686,N_16076,N_16174);
nor U17687 (N_17687,N_15612,N_16448);
xor U17688 (N_17688,N_16009,N_16171);
and U17689 (N_17689,N_16122,N_15947);
nand U17690 (N_17690,N_16115,N_16486);
xnor U17691 (N_17691,N_16629,N_15808);
and U17692 (N_17692,N_15718,N_16765);
xnor U17693 (N_17693,N_15867,N_16372);
and U17694 (N_17694,N_15968,N_16462);
xor U17695 (N_17695,N_16367,N_16133);
xnor U17696 (N_17696,N_16258,N_16371);
nor U17697 (N_17697,N_16303,N_15911);
nor U17698 (N_17698,N_15648,N_16392);
xor U17699 (N_17699,N_16760,N_15926);
nor U17700 (N_17700,N_16542,N_16772);
nor U17701 (N_17701,N_16796,N_16452);
and U17702 (N_17702,N_16355,N_15715);
nand U17703 (N_17703,N_15742,N_15710);
nand U17704 (N_17704,N_16194,N_16018);
and U17705 (N_17705,N_15695,N_16655);
or U17706 (N_17706,N_16054,N_16150);
xnor U17707 (N_17707,N_15701,N_16692);
nand U17708 (N_17708,N_15785,N_15955);
xnor U17709 (N_17709,N_16053,N_16021);
nand U17710 (N_17710,N_16163,N_16753);
or U17711 (N_17711,N_16262,N_15961);
xnor U17712 (N_17712,N_16524,N_16668);
and U17713 (N_17713,N_16262,N_16515);
nand U17714 (N_17714,N_16341,N_16726);
nand U17715 (N_17715,N_15883,N_15605);
nand U17716 (N_17716,N_16250,N_16079);
nand U17717 (N_17717,N_15933,N_16298);
nor U17718 (N_17718,N_16142,N_16587);
nand U17719 (N_17719,N_16684,N_16288);
nand U17720 (N_17720,N_16535,N_15880);
and U17721 (N_17721,N_16034,N_16734);
nand U17722 (N_17722,N_16372,N_16586);
and U17723 (N_17723,N_16408,N_15864);
or U17724 (N_17724,N_15894,N_16022);
and U17725 (N_17725,N_16446,N_16245);
and U17726 (N_17726,N_16051,N_16506);
nor U17727 (N_17727,N_15872,N_15893);
xnor U17728 (N_17728,N_15725,N_16027);
nor U17729 (N_17729,N_15706,N_15981);
and U17730 (N_17730,N_16412,N_16019);
xor U17731 (N_17731,N_16474,N_16011);
or U17732 (N_17732,N_15875,N_16398);
and U17733 (N_17733,N_16348,N_16256);
or U17734 (N_17734,N_15755,N_16510);
and U17735 (N_17735,N_16624,N_16743);
or U17736 (N_17736,N_15602,N_15607);
xnor U17737 (N_17737,N_16194,N_15853);
nor U17738 (N_17738,N_15698,N_16390);
or U17739 (N_17739,N_15706,N_16444);
nor U17740 (N_17740,N_16547,N_16526);
nor U17741 (N_17741,N_16393,N_16009);
nor U17742 (N_17742,N_16384,N_15646);
nor U17743 (N_17743,N_16474,N_16036);
nor U17744 (N_17744,N_16402,N_16453);
nor U17745 (N_17745,N_16092,N_16324);
nand U17746 (N_17746,N_15640,N_16236);
and U17747 (N_17747,N_15861,N_16158);
or U17748 (N_17748,N_15982,N_16362);
xor U17749 (N_17749,N_15799,N_16247);
xor U17750 (N_17750,N_15747,N_16545);
or U17751 (N_17751,N_16357,N_16033);
xor U17752 (N_17752,N_16257,N_16217);
nor U17753 (N_17753,N_16101,N_15792);
nand U17754 (N_17754,N_16454,N_16689);
nor U17755 (N_17755,N_16401,N_16459);
xnor U17756 (N_17756,N_16564,N_16329);
and U17757 (N_17757,N_16286,N_16549);
nor U17758 (N_17758,N_16335,N_16041);
nor U17759 (N_17759,N_16037,N_16628);
and U17760 (N_17760,N_16487,N_16675);
nor U17761 (N_17761,N_16134,N_16375);
nor U17762 (N_17762,N_15893,N_16726);
nand U17763 (N_17763,N_15923,N_16474);
nor U17764 (N_17764,N_16612,N_16600);
or U17765 (N_17765,N_15688,N_15689);
and U17766 (N_17766,N_16706,N_16480);
nand U17767 (N_17767,N_16685,N_15760);
nand U17768 (N_17768,N_16119,N_16408);
and U17769 (N_17769,N_15850,N_15959);
xor U17770 (N_17770,N_16129,N_16594);
or U17771 (N_17771,N_16607,N_16146);
nor U17772 (N_17772,N_15620,N_16158);
nor U17773 (N_17773,N_16667,N_15630);
xnor U17774 (N_17774,N_15934,N_16797);
nand U17775 (N_17775,N_15838,N_16284);
or U17776 (N_17776,N_16109,N_15609);
or U17777 (N_17777,N_15658,N_16627);
and U17778 (N_17778,N_15705,N_16780);
or U17779 (N_17779,N_15685,N_16031);
and U17780 (N_17780,N_16377,N_15786);
nand U17781 (N_17781,N_15817,N_16346);
nand U17782 (N_17782,N_16448,N_15759);
nand U17783 (N_17783,N_16641,N_16749);
xor U17784 (N_17784,N_15846,N_16257);
nand U17785 (N_17785,N_15783,N_16010);
and U17786 (N_17786,N_16598,N_16653);
and U17787 (N_17787,N_15813,N_16043);
and U17788 (N_17788,N_15614,N_15963);
nand U17789 (N_17789,N_16032,N_16170);
or U17790 (N_17790,N_16305,N_16508);
nand U17791 (N_17791,N_16412,N_16223);
nand U17792 (N_17792,N_16342,N_16676);
and U17793 (N_17793,N_15833,N_15744);
and U17794 (N_17794,N_15854,N_16525);
or U17795 (N_17795,N_15827,N_16133);
nor U17796 (N_17796,N_15835,N_15634);
nand U17797 (N_17797,N_15670,N_16591);
nand U17798 (N_17798,N_16663,N_15635);
or U17799 (N_17799,N_16042,N_16335);
or U17800 (N_17800,N_15602,N_15672);
and U17801 (N_17801,N_15784,N_16397);
and U17802 (N_17802,N_15937,N_16691);
and U17803 (N_17803,N_16217,N_16353);
or U17804 (N_17804,N_16271,N_16108);
nor U17805 (N_17805,N_16530,N_16711);
xnor U17806 (N_17806,N_15618,N_15601);
and U17807 (N_17807,N_15612,N_16585);
xor U17808 (N_17808,N_16256,N_16027);
or U17809 (N_17809,N_16446,N_16550);
xnor U17810 (N_17810,N_15758,N_16799);
and U17811 (N_17811,N_16713,N_16001);
nor U17812 (N_17812,N_16187,N_16163);
and U17813 (N_17813,N_15874,N_16500);
or U17814 (N_17814,N_16590,N_16570);
nand U17815 (N_17815,N_15923,N_16148);
and U17816 (N_17816,N_15608,N_16615);
or U17817 (N_17817,N_16551,N_15955);
nor U17818 (N_17818,N_16123,N_16164);
and U17819 (N_17819,N_16616,N_16233);
or U17820 (N_17820,N_15919,N_16059);
or U17821 (N_17821,N_16515,N_16481);
nand U17822 (N_17822,N_16106,N_16370);
nor U17823 (N_17823,N_15920,N_16347);
nand U17824 (N_17824,N_15662,N_15738);
or U17825 (N_17825,N_15616,N_16226);
nand U17826 (N_17826,N_16440,N_16165);
and U17827 (N_17827,N_16537,N_15765);
xor U17828 (N_17828,N_16280,N_16070);
nand U17829 (N_17829,N_16737,N_16105);
nand U17830 (N_17830,N_16278,N_15753);
nor U17831 (N_17831,N_16382,N_16204);
nand U17832 (N_17832,N_15998,N_16660);
and U17833 (N_17833,N_16761,N_16135);
nor U17834 (N_17834,N_15647,N_15631);
and U17835 (N_17835,N_16060,N_16562);
nor U17836 (N_17836,N_15951,N_16190);
or U17837 (N_17837,N_15739,N_15953);
or U17838 (N_17838,N_15790,N_16745);
xnor U17839 (N_17839,N_16442,N_15705);
or U17840 (N_17840,N_16761,N_16587);
nand U17841 (N_17841,N_16768,N_16552);
nand U17842 (N_17842,N_15769,N_16429);
nand U17843 (N_17843,N_15678,N_16513);
and U17844 (N_17844,N_16653,N_16226);
and U17845 (N_17845,N_16435,N_16674);
nand U17846 (N_17846,N_16612,N_16330);
and U17847 (N_17847,N_15806,N_15614);
xor U17848 (N_17848,N_15828,N_15653);
xnor U17849 (N_17849,N_16598,N_16699);
and U17850 (N_17850,N_15979,N_15762);
xnor U17851 (N_17851,N_16713,N_16736);
nand U17852 (N_17852,N_16654,N_15748);
xor U17853 (N_17853,N_16364,N_16153);
nor U17854 (N_17854,N_16251,N_15887);
nand U17855 (N_17855,N_15911,N_16543);
or U17856 (N_17856,N_16332,N_15613);
or U17857 (N_17857,N_16351,N_16255);
nand U17858 (N_17858,N_15905,N_15624);
or U17859 (N_17859,N_16636,N_16793);
and U17860 (N_17860,N_15993,N_15992);
nor U17861 (N_17861,N_16486,N_16084);
and U17862 (N_17862,N_16156,N_16644);
xnor U17863 (N_17863,N_16618,N_16357);
nor U17864 (N_17864,N_16717,N_16408);
xnor U17865 (N_17865,N_16785,N_16503);
or U17866 (N_17866,N_16547,N_16456);
or U17867 (N_17867,N_16211,N_15609);
and U17868 (N_17868,N_15829,N_16156);
and U17869 (N_17869,N_15777,N_16294);
xnor U17870 (N_17870,N_15956,N_15781);
nor U17871 (N_17871,N_15861,N_16789);
or U17872 (N_17872,N_16378,N_16700);
or U17873 (N_17873,N_15651,N_15799);
xor U17874 (N_17874,N_16177,N_16679);
nor U17875 (N_17875,N_16514,N_16712);
and U17876 (N_17876,N_16364,N_16246);
or U17877 (N_17877,N_16597,N_15670);
nand U17878 (N_17878,N_15897,N_16555);
nand U17879 (N_17879,N_15999,N_16386);
nand U17880 (N_17880,N_16723,N_15702);
xnor U17881 (N_17881,N_16196,N_15782);
and U17882 (N_17882,N_16467,N_16730);
nor U17883 (N_17883,N_16371,N_16004);
nand U17884 (N_17884,N_15977,N_15739);
and U17885 (N_17885,N_16208,N_16059);
nor U17886 (N_17886,N_16507,N_16149);
nand U17887 (N_17887,N_15617,N_16729);
nor U17888 (N_17888,N_16099,N_15921);
nor U17889 (N_17889,N_16596,N_16438);
nand U17890 (N_17890,N_16508,N_15716);
xor U17891 (N_17891,N_16579,N_16191);
nand U17892 (N_17892,N_16678,N_16608);
and U17893 (N_17893,N_15964,N_15955);
nand U17894 (N_17894,N_15954,N_16015);
nand U17895 (N_17895,N_15686,N_15677);
xnor U17896 (N_17896,N_16694,N_15930);
and U17897 (N_17897,N_16655,N_16355);
xor U17898 (N_17898,N_16154,N_16520);
and U17899 (N_17899,N_16249,N_16290);
nand U17900 (N_17900,N_16153,N_15772);
or U17901 (N_17901,N_15628,N_16752);
or U17902 (N_17902,N_15702,N_16079);
and U17903 (N_17903,N_15900,N_16081);
or U17904 (N_17904,N_16063,N_16450);
or U17905 (N_17905,N_15826,N_16798);
nand U17906 (N_17906,N_15730,N_16018);
nand U17907 (N_17907,N_16099,N_15986);
or U17908 (N_17908,N_16679,N_15714);
or U17909 (N_17909,N_16569,N_16539);
and U17910 (N_17910,N_16656,N_16558);
and U17911 (N_17911,N_15870,N_15672);
xnor U17912 (N_17912,N_16158,N_16787);
and U17913 (N_17913,N_15803,N_16038);
or U17914 (N_17914,N_16482,N_16602);
nor U17915 (N_17915,N_16366,N_16334);
and U17916 (N_17916,N_16799,N_16296);
or U17917 (N_17917,N_16665,N_15953);
nand U17918 (N_17918,N_15765,N_16601);
nand U17919 (N_17919,N_16355,N_16714);
or U17920 (N_17920,N_16075,N_16270);
xnor U17921 (N_17921,N_16515,N_16020);
nand U17922 (N_17922,N_16446,N_16004);
nand U17923 (N_17923,N_16107,N_16782);
and U17924 (N_17924,N_15904,N_15941);
and U17925 (N_17925,N_16026,N_16737);
nor U17926 (N_17926,N_16220,N_16776);
nand U17927 (N_17927,N_16395,N_15803);
nand U17928 (N_17928,N_16303,N_16204);
xor U17929 (N_17929,N_16267,N_15793);
xnor U17930 (N_17930,N_16076,N_16495);
xor U17931 (N_17931,N_16453,N_16240);
or U17932 (N_17932,N_16249,N_15996);
or U17933 (N_17933,N_15956,N_16575);
nor U17934 (N_17934,N_15701,N_15730);
nor U17935 (N_17935,N_16786,N_15874);
or U17936 (N_17936,N_16177,N_16221);
nand U17937 (N_17937,N_16512,N_15625);
or U17938 (N_17938,N_16582,N_15776);
nor U17939 (N_17939,N_16521,N_15845);
nand U17940 (N_17940,N_16304,N_15852);
nand U17941 (N_17941,N_16247,N_16356);
nor U17942 (N_17942,N_16094,N_16123);
nand U17943 (N_17943,N_16404,N_16712);
and U17944 (N_17944,N_16289,N_16288);
nor U17945 (N_17945,N_16268,N_15817);
nand U17946 (N_17946,N_15627,N_16216);
nand U17947 (N_17947,N_16212,N_15801);
and U17948 (N_17948,N_15724,N_15706);
or U17949 (N_17949,N_16023,N_15671);
nor U17950 (N_17950,N_15868,N_16514);
nand U17951 (N_17951,N_16615,N_16051);
nor U17952 (N_17952,N_16416,N_16043);
xor U17953 (N_17953,N_16214,N_16759);
or U17954 (N_17954,N_16545,N_16444);
and U17955 (N_17955,N_16258,N_16706);
xor U17956 (N_17956,N_15748,N_16500);
nor U17957 (N_17957,N_16353,N_16623);
and U17958 (N_17958,N_16372,N_16782);
nor U17959 (N_17959,N_16783,N_16101);
nor U17960 (N_17960,N_16433,N_16412);
nor U17961 (N_17961,N_16544,N_16644);
nor U17962 (N_17962,N_16007,N_16791);
and U17963 (N_17963,N_15811,N_16028);
nand U17964 (N_17964,N_16433,N_16508);
xnor U17965 (N_17965,N_15870,N_16509);
xnor U17966 (N_17966,N_15788,N_16125);
nor U17967 (N_17967,N_16237,N_16792);
or U17968 (N_17968,N_15866,N_16048);
nor U17969 (N_17969,N_15913,N_15984);
nand U17970 (N_17970,N_16528,N_16669);
xnor U17971 (N_17971,N_16423,N_16092);
xor U17972 (N_17972,N_16272,N_16468);
nand U17973 (N_17973,N_16398,N_15720);
and U17974 (N_17974,N_16242,N_16279);
or U17975 (N_17975,N_16549,N_15952);
and U17976 (N_17976,N_15996,N_16569);
xor U17977 (N_17977,N_16755,N_15948);
nand U17978 (N_17978,N_16434,N_16353);
nand U17979 (N_17979,N_16567,N_16748);
or U17980 (N_17980,N_16265,N_16616);
and U17981 (N_17981,N_15726,N_15628);
and U17982 (N_17982,N_16319,N_16711);
and U17983 (N_17983,N_16005,N_16788);
xnor U17984 (N_17984,N_16299,N_16210);
or U17985 (N_17985,N_15858,N_16388);
and U17986 (N_17986,N_16133,N_16095);
xor U17987 (N_17987,N_16151,N_16765);
xnor U17988 (N_17988,N_16237,N_16227);
nor U17989 (N_17989,N_15646,N_16238);
or U17990 (N_17990,N_16728,N_16451);
and U17991 (N_17991,N_16326,N_16601);
and U17992 (N_17992,N_15653,N_15996);
xnor U17993 (N_17993,N_16027,N_16442);
or U17994 (N_17994,N_16786,N_15947);
nor U17995 (N_17995,N_16130,N_15690);
and U17996 (N_17996,N_16175,N_16184);
or U17997 (N_17997,N_16343,N_16120);
or U17998 (N_17998,N_15810,N_15779);
or U17999 (N_17999,N_16572,N_16759);
and U18000 (N_18000,N_17364,N_17240);
nand U18001 (N_18001,N_16841,N_17348);
or U18002 (N_18002,N_17310,N_17816);
nor U18003 (N_18003,N_17641,N_17646);
and U18004 (N_18004,N_16907,N_17077);
nor U18005 (N_18005,N_17629,N_17184);
or U18006 (N_18006,N_17623,N_17100);
and U18007 (N_18007,N_17192,N_17758);
nor U18008 (N_18008,N_17849,N_17377);
nand U18009 (N_18009,N_16962,N_17673);
and U18010 (N_18010,N_17877,N_17667);
nand U18011 (N_18011,N_17954,N_17945);
or U18012 (N_18012,N_17859,N_17135);
and U18013 (N_18013,N_16982,N_17122);
or U18014 (N_18014,N_17761,N_17888);
or U18015 (N_18015,N_16884,N_17148);
or U18016 (N_18016,N_16826,N_17496);
or U18017 (N_18017,N_16993,N_17666);
nor U18018 (N_18018,N_17055,N_17004);
nand U18019 (N_18019,N_17752,N_17337);
nor U18020 (N_18020,N_17225,N_16895);
or U18021 (N_18021,N_17080,N_17290);
nand U18022 (N_18022,N_16900,N_17716);
and U18023 (N_18023,N_17145,N_17901);
or U18024 (N_18024,N_17951,N_16913);
nand U18025 (N_18025,N_17132,N_17168);
or U18026 (N_18026,N_17340,N_17410);
nand U18027 (N_18027,N_16911,N_17297);
nor U18028 (N_18028,N_17490,N_16844);
nor U18029 (N_18029,N_16818,N_17081);
nor U18030 (N_18030,N_17579,N_16978);
nor U18031 (N_18031,N_16922,N_17458);
nor U18032 (N_18032,N_17737,N_17210);
nand U18033 (N_18033,N_17228,N_17281);
and U18034 (N_18034,N_17968,N_16874);
or U18035 (N_18035,N_17024,N_17986);
xnor U18036 (N_18036,N_17503,N_17621);
nand U18037 (N_18037,N_17524,N_17067);
or U18038 (N_18038,N_17618,N_16887);
or U18039 (N_18039,N_17078,N_16921);
xor U18040 (N_18040,N_17560,N_17513);
or U18041 (N_18041,N_16869,N_17108);
nor U18042 (N_18042,N_17685,N_16805);
and U18043 (N_18043,N_16981,N_17878);
nor U18044 (N_18044,N_17101,N_17527);
and U18045 (N_18045,N_17402,N_17703);
or U18046 (N_18046,N_17766,N_16945);
nor U18047 (N_18047,N_16901,N_17076);
and U18048 (N_18048,N_17091,N_16850);
nand U18049 (N_18049,N_17537,N_17043);
or U18050 (N_18050,N_17614,N_17701);
and U18051 (N_18051,N_17834,N_17116);
xnor U18052 (N_18052,N_17987,N_17421);
xor U18053 (N_18053,N_17399,N_17050);
xnor U18054 (N_18054,N_17429,N_16822);
nand U18055 (N_18055,N_17449,N_17584);
nand U18056 (N_18056,N_17327,N_17261);
nand U18057 (N_18057,N_17869,N_17131);
xnor U18058 (N_18058,N_16983,N_16906);
xor U18059 (N_18059,N_17475,N_17670);
nor U18060 (N_18060,N_17709,N_17549);
and U18061 (N_18061,N_16834,N_17936);
xnor U18062 (N_18062,N_17523,N_17127);
nor U18063 (N_18063,N_17124,N_17249);
nand U18064 (N_18064,N_16836,N_16927);
and U18065 (N_18065,N_17084,N_17931);
nand U18066 (N_18066,N_17302,N_17823);
and U18067 (N_18067,N_16828,N_17982);
or U18068 (N_18068,N_17197,N_17052);
and U18069 (N_18069,N_17495,N_17895);
nor U18070 (N_18070,N_17640,N_17587);
and U18071 (N_18071,N_17468,N_17238);
and U18072 (N_18072,N_17740,N_17346);
and U18073 (N_18073,N_17999,N_17072);
and U18074 (N_18074,N_17710,N_17383);
or U18075 (N_18075,N_17892,N_17543);
and U18076 (N_18076,N_17242,N_17967);
xnor U18077 (N_18077,N_17023,N_17368);
nor U18078 (N_18078,N_17218,N_17862);
nor U18079 (N_18079,N_17566,N_17095);
xnor U18080 (N_18080,N_17934,N_16827);
nand U18081 (N_18081,N_17759,N_17071);
or U18082 (N_18082,N_17564,N_17381);
and U18083 (N_18083,N_17448,N_17734);
nand U18084 (N_18084,N_17409,N_17048);
nand U18085 (N_18085,N_17502,N_17695);
nand U18086 (N_18086,N_17167,N_17994);
or U18087 (N_18087,N_17263,N_17802);
and U18088 (N_18088,N_17217,N_17749);
and U18089 (N_18089,N_16871,N_16939);
and U18090 (N_18090,N_16882,N_17099);
xor U18091 (N_18091,N_17785,N_17721);
xor U18092 (N_18092,N_17158,N_17470);
and U18093 (N_18093,N_17864,N_17649);
nand U18094 (N_18094,N_17684,N_17571);
or U18095 (N_18095,N_17898,N_17538);
nand U18096 (N_18096,N_17041,N_17234);
xor U18097 (N_18097,N_17021,N_17746);
or U18098 (N_18098,N_17034,N_17014);
nor U18099 (N_18099,N_16925,N_17985);
and U18100 (N_18100,N_17176,N_17501);
and U18101 (N_18101,N_17635,N_17844);
xnor U18102 (N_18102,N_17057,N_17175);
nor U18103 (N_18103,N_17605,N_16876);
or U18104 (N_18104,N_17883,N_17322);
or U18105 (N_18105,N_17194,N_17277);
and U18106 (N_18106,N_17965,N_16917);
or U18107 (N_18107,N_17296,N_16999);
nand U18108 (N_18108,N_17966,N_17569);
or U18109 (N_18109,N_17442,N_17731);
nand U18110 (N_18110,N_17704,N_17254);
and U18111 (N_18111,N_17995,N_17642);
and U18112 (N_18112,N_17585,N_17222);
and U18113 (N_18113,N_17972,N_17239);
and U18114 (N_18114,N_17483,N_17195);
xor U18115 (N_18115,N_17547,N_16992);
or U18116 (N_18116,N_17265,N_17284);
xnor U18117 (N_18117,N_17374,N_17891);
nor U18118 (N_18118,N_17899,N_17671);
and U18119 (N_18119,N_17434,N_17793);
xor U18120 (N_18120,N_16944,N_17732);
xnor U18121 (N_18121,N_17681,N_17988);
nor U18122 (N_18122,N_17427,N_17253);
nand U18123 (N_18123,N_17736,N_17541);
nand U18124 (N_18124,N_17404,N_17847);
and U18125 (N_18125,N_17181,N_17497);
nand U18126 (N_18126,N_16909,N_17329);
and U18127 (N_18127,N_17193,N_17748);
and U18128 (N_18128,N_17262,N_17879);
nand U18129 (N_18129,N_17609,N_17688);
xnor U18130 (N_18130,N_17622,N_17713);
and U18131 (N_18131,N_17797,N_16879);
nand U18132 (N_18132,N_17143,N_17663);
xor U18133 (N_18133,N_17515,N_16984);
nand U18134 (N_18134,N_17930,N_17370);
xor U18135 (N_18135,N_16866,N_17976);
xnor U18136 (N_18136,N_17577,N_17744);
and U18137 (N_18137,N_17516,N_17717);
nor U18138 (N_18138,N_17038,N_17506);
or U18139 (N_18139,N_17856,N_17973);
nor U18140 (N_18140,N_17173,N_17300);
nor U18141 (N_18141,N_17546,N_17820);
xnor U18142 (N_18142,N_16891,N_17144);
nand U18143 (N_18143,N_16898,N_17489);
or U18144 (N_18144,N_16812,N_17147);
and U18145 (N_18145,N_17590,N_16801);
nand U18146 (N_18146,N_17104,N_17119);
and U18147 (N_18147,N_17990,N_17697);
and U18148 (N_18148,N_17806,N_17553);
nand U18149 (N_18149,N_17243,N_17433);
xnor U18150 (N_18150,N_17159,N_17803);
nor U18151 (N_18151,N_16936,N_17616);
and U18152 (N_18152,N_17015,N_17380);
and U18153 (N_18153,N_17397,N_17728);
nor U18154 (N_18154,N_16859,N_16855);
or U18155 (N_18155,N_17114,N_16896);
nor U18156 (N_18156,N_17037,N_17852);
nand U18157 (N_18157,N_17298,N_17267);
or U18158 (N_18158,N_17059,N_17929);
or U18159 (N_18159,N_17186,N_17794);
and U18160 (N_18160,N_17418,N_17657);
or U18161 (N_18161,N_17873,N_17705);
or U18162 (N_18162,N_17465,N_16967);
or U18163 (N_18163,N_16905,N_16990);
and U18164 (N_18164,N_16964,N_17808);
xor U18165 (N_18165,N_17536,N_17739);
xor U18166 (N_18166,N_17610,N_17010);
and U18167 (N_18167,N_17426,N_17318);
nor U18168 (N_18168,N_17919,N_17304);
xor U18169 (N_18169,N_17113,N_17435);
xnor U18170 (N_18170,N_17837,N_17578);
or U18171 (N_18171,N_17157,N_17530);
nand U18172 (N_18172,N_17089,N_17109);
or U18173 (N_18173,N_17593,N_17488);
or U18174 (N_18174,N_17164,N_17648);
or U18175 (N_18175,N_17805,N_17678);
xnor U18176 (N_18176,N_17958,N_17884);
xor U18177 (N_18177,N_17767,N_17013);
xor U18178 (N_18178,N_16889,N_17920);
xor U18179 (N_18179,N_17248,N_17970);
and U18180 (N_18180,N_17338,N_16833);
nor U18181 (N_18181,N_17754,N_17692);
xor U18182 (N_18182,N_17473,N_17063);
xnor U18183 (N_18183,N_17851,N_17129);
xor U18184 (N_18184,N_17075,N_17796);
nand U18185 (N_18185,N_17682,N_17382);
nand U18186 (N_18186,N_17742,N_17664);
or U18187 (N_18187,N_17366,N_16975);
or U18188 (N_18188,N_16814,N_17983);
or U18189 (N_18189,N_17904,N_17362);
nor U18190 (N_18190,N_17231,N_16858);
nor U18191 (N_18191,N_17843,N_17001);
and U18192 (N_18192,N_17392,N_17699);
nor U18193 (N_18193,N_17624,N_17203);
or U18194 (N_18194,N_17450,N_17079);
nand U18195 (N_18195,N_17092,N_16877);
xnor U18196 (N_18196,N_17950,N_17464);
xor U18197 (N_18197,N_17961,N_17532);
nand U18198 (N_18198,N_16809,N_17662);
or U18199 (N_18199,N_16848,N_17997);
and U18200 (N_18200,N_17319,N_17125);
or U18201 (N_18201,N_17839,N_17485);
or U18202 (N_18202,N_17918,N_17902);
and U18203 (N_18203,N_17923,N_17581);
nor U18204 (N_18204,N_17514,N_17783);
xor U18205 (N_18205,N_17006,N_17601);
and U18206 (N_18206,N_17446,N_17595);
and U18207 (N_18207,N_17447,N_17051);
nor U18208 (N_18208,N_17555,N_17224);
nor U18209 (N_18209,N_17712,N_17706);
or U18210 (N_18210,N_17860,N_17762);
and U18211 (N_18211,N_16968,N_17975);
and U18212 (N_18212,N_16838,N_17198);
nor U18213 (N_18213,N_17894,N_17280);
xnor U18214 (N_18214,N_17611,N_17285);
or U18215 (N_18215,N_17227,N_17669);
and U18216 (N_18216,N_17617,N_17299);
xor U18217 (N_18217,N_16943,N_16923);
nand U18218 (N_18218,N_17525,N_17686);
or U18219 (N_18219,N_17369,N_17720);
xor U18220 (N_18220,N_17508,N_17065);
nor U18221 (N_18221,N_17343,N_17871);
nand U18222 (N_18222,N_17171,N_17137);
or U18223 (N_18223,N_17729,N_17628);
xor U18224 (N_18224,N_16952,N_17246);
xor U18225 (N_18225,N_16947,N_17947);
or U18226 (N_18226,N_17120,N_17565);
or U18227 (N_18227,N_17942,N_17411);
and U18228 (N_18228,N_17341,N_17317);
and U18229 (N_18229,N_17308,N_17066);
or U18230 (N_18230,N_17551,N_17260);
or U18231 (N_18231,N_17866,N_17165);
xor U18232 (N_18232,N_17268,N_17439);
nand U18233 (N_18233,N_17801,N_17756);
and U18234 (N_18234,N_16807,N_17251);
nor U18235 (N_18235,N_17028,N_17134);
nor U18236 (N_18236,N_17870,N_17890);
nand U18237 (N_18237,N_17645,N_17840);
nand U18238 (N_18238,N_17303,N_17707);
nor U18239 (N_18239,N_17539,N_17149);
and U18240 (N_18240,N_17906,N_17196);
or U18241 (N_18241,N_16878,N_17278);
xnor U18242 (N_18242,N_17389,N_16926);
and U18243 (N_18243,N_17693,N_17757);
and U18244 (N_18244,N_17674,N_17575);
or U18245 (N_18245,N_17255,N_17353);
or U18246 (N_18246,N_16919,N_17054);
and U18247 (N_18247,N_16846,N_17781);
nand U18248 (N_18248,N_17221,N_17305);
nand U18249 (N_18249,N_16890,N_16932);
and U18250 (N_18250,N_17123,N_17924);
xor U18251 (N_18251,N_17107,N_17270);
nor U18252 (N_18252,N_16847,N_17312);
or U18253 (N_18253,N_16872,N_17311);
and U18254 (N_18254,N_17003,N_17455);
xnor U18255 (N_18255,N_17774,N_17580);
and U18256 (N_18256,N_17651,N_17033);
xnor U18257 (N_18257,N_17215,N_17384);
xor U18258 (N_18258,N_17454,N_17842);
or U18259 (N_18259,N_17955,N_16934);
or U18260 (N_18260,N_17128,N_17658);
and U18261 (N_18261,N_17599,N_17292);
xnor U18262 (N_18262,N_17561,N_17600);
or U18263 (N_18263,N_17183,N_17726);
or U18264 (N_18264,N_17769,N_17563);
nor U18265 (N_18265,N_17428,N_17828);
and U18266 (N_18266,N_17582,N_17387);
and U18267 (N_18267,N_17675,N_17882);
or U18268 (N_18268,N_17815,N_17250);
and U18269 (N_18269,N_17174,N_17462);
nor U18270 (N_18270,N_17804,N_16885);
or U18271 (N_18271,N_17719,N_17938);
nand U18272 (N_18272,N_17160,N_17235);
xor U18273 (N_18273,N_17474,N_17336);
and U18274 (N_18274,N_16970,N_17944);
and U18275 (N_18275,N_17914,N_17504);
or U18276 (N_18276,N_17291,N_16963);
xor U18277 (N_18277,N_17625,N_16986);
nand U18278 (N_18278,N_17472,N_17591);
or U18279 (N_18279,N_17588,N_17596);
nor U18280 (N_18280,N_17136,N_17032);
or U18281 (N_18281,N_17069,N_16953);
or U18282 (N_18282,N_17214,N_17492);
nand U18283 (N_18283,N_16980,N_17589);
xnor U18284 (N_18284,N_16816,N_17948);
nand U18285 (N_18285,N_17416,N_17632);
nand U18286 (N_18286,N_17391,N_17654);
nor U18287 (N_18287,N_16957,N_17204);
nor U18288 (N_18288,N_17026,N_17896);
or U18289 (N_18289,N_17324,N_17573);
xor U18290 (N_18290,N_17367,N_17825);
and U18291 (N_18291,N_17469,N_17090);
and U18292 (N_18292,N_17019,N_17049);
or U18293 (N_18293,N_17979,N_17403);
nand U18294 (N_18294,N_16966,N_17738);
nand U18295 (N_18295,N_17521,N_17724);
xor U18296 (N_18296,N_17045,N_17396);
or U18297 (N_18297,N_17482,N_17103);
xor U18298 (N_18298,N_16883,N_17245);
xor U18299 (N_18299,N_17112,N_16832);
nor U18300 (N_18300,N_17208,N_16976);
nand U18301 (N_18301,N_17638,N_17971);
and U18302 (N_18302,N_17111,N_17598);
or U18303 (N_18303,N_17633,N_17205);
nand U18304 (N_18304,N_17486,N_16802);
nand U18305 (N_18305,N_16950,N_17544);
xor U18306 (N_18306,N_17799,N_17309);
xor U18307 (N_18307,N_17574,N_17620);
and U18308 (N_18308,N_17375,N_17874);
and U18309 (N_18309,N_17928,N_17730);
xor U18310 (N_18310,N_16820,N_17957);
nor U18311 (N_18311,N_17548,N_17060);
or U18312 (N_18312,N_17778,N_16830);
or U18313 (N_18313,N_16839,N_17567);
xnor U18314 (N_18314,N_16835,N_16861);
nand U18315 (N_18315,N_17977,N_17349);
or U18316 (N_18316,N_17008,N_17679);
or U18317 (N_18317,N_17354,N_17334);
or U18318 (N_18318,N_17660,N_16849);
xnor U18319 (N_18319,N_16920,N_17035);
nor U18320 (N_18320,N_17018,N_17911);
or U18321 (N_18321,N_17763,N_17542);
and U18322 (N_18322,N_17202,N_17594);
nor U18323 (N_18323,N_17405,N_17022);
nor U18324 (N_18324,N_17325,N_17875);
nand U18325 (N_18325,N_17016,N_17518);
nand U18326 (N_18326,N_17096,N_17313);
or U18327 (N_18327,N_17845,N_17833);
or U18328 (N_18328,N_17652,N_17810);
and U18329 (N_18329,N_17187,N_17415);
or U18330 (N_18330,N_17727,N_17020);
or U18331 (N_18331,N_16902,N_16823);
and U18332 (N_18332,N_17420,N_17247);
and U18333 (N_18333,N_17180,N_17953);
or U18334 (N_18334,N_17230,N_17419);
or U18335 (N_18335,N_17074,N_17959);
and U18336 (N_18336,N_17960,N_17848);
nor U18337 (N_18337,N_17602,N_17216);
xnor U18338 (N_18338,N_17283,N_17913);
nand U18339 (N_18339,N_16880,N_17690);
nor U18340 (N_18340,N_17150,N_17784);
and U18341 (N_18341,N_17282,N_17212);
nor U18342 (N_18342,N_16935,N_17677);
nor U18343 (N_18343,N_17656,N_17443);
nor U18344 (N_18344,N_17597,N_17499);
nand U18345 (N_18345,N_17698,N_17639);
and U18346 (N_18346,N_17105,N_17494);
or U18347 (N_18347,N_17572,N_17330);
and U18348 (N_18348,N_17926,N_16863);
nor U18349 (N_18349,N_17694,N_16965);
nor U18350 (N_18350,N_16806,N_17715);
and U18351 (N_18351,N_17522,N_17829);
nor U18352 (N_18352,N_17743,N_17082);
or U18353 (N_18353,N_16867,N_16951);
and U18354 (N_18354,N_17306,N_17029);
nor U18355 (N_18355,N_16933,N_17142);
and U18356 (N_18356,N_17272,N_17903);
nor U18357 (N_18357,N_17155,N_17770);
xor U18358 (N_18358,N_16930,N_17819);
xnor U18359 (N_18359,N_17991,N_17407);
or U18360 (N_18360,N_17937,N_17735);
nor U18361 (N_18361,N_17812,N_16973);
nor U18362 (N_18362,N_17307,N_17011);
nand U18363 (N_18363,N_16987,N_16995);
nor U18364 (N_18364,N_17627,N_16804);
and U18365 (N_18365,N_17252,N_17905);
nand U18366 (N_18366,N_16937,N_17568);
and U18367 (N_18367,N_16958,N_16940);
nor U18368 (N_18368,N_17718,N_17725);
or U18369 (N_18369,N_17047,N_17027);
nor U18370 (N_18370,N_17347,N_17413);
and U18371 (N_18371,N_17378,N_17333);
xnor U18372 (N_18372,N_17294,N_17151);
xor U18373 (N_18373,N_17529,N_17887);
or U18374 (N_18374,N_17432,N_17753);
or U18375 (N_18375,N_16994,N_17807);
or U18376 (N_18376,N_17691,N_16843);
or U18377 (N_18377,N_17244,N_17655);
or U18378 (N_18378,N_17213,N_17273);
nor U18379 (N_18379,N_17335,N_17363);
xor U18380 (N_18380,N_17741,N_17643);
nor U18381 (N_18381,N_16854,N_17339);
nand U18382 (N_18382,N_16931,N_17189);
nor U18383 (N_18383,N_17241,N_17821);
nand U18384 (N_18384,N_17751,N_17814);
or U18385 (N_18385,N_17838,N_17893);
or U18386 (N_18386,N_17800,N_17361);
nor U18387 (N_18387,N_17876,N_17780);
nand U18388 (N_18388,N_16893,N_17962);
nand U18389 (N_18389,N_17162,N_17714);
nor U18390 (N_18390,N_16831,N_17417);
or U18391 (N_18391,N_17626,N_17236);
or U18392 (N_18392,N_17747,N_17453);
xor U18393 (N_18393,N_17659,N_16998);
nand U18394 (N_18394,N_16969,N_17786);
or U18395 (N_18395,N_16904,N_17009);
nor U18396 (N_18396,N_17535,N_17394);
or U18397 (N_18397,N_17776,N_17723);
xnor U18398 (N_18398,N_17030,N_17696);
and U18399 (N_18399,N_17156,N_16948);
xor U18400 (N_18400,N_16860,N_17811);
nor U18401 (N_18401,N_17771,N_17117);
xor U18402 (N_18402,N_16903,N_17907);
nor U18403 (N_18403,N_17813,N_17817);
xnor U18404 (N_18404,N_17445,N_17088);
nor U18405 (N_18405,N_16821,N_17841);
xnor U18406 (N_18406,N_17355,N_17326);
xor U18407 (N_18407,N_17855,N_17676);
nand U18408 (N_18408,N_17526,N_16870);
nand U18409 (N_18409,N_17031,N_17083);
xnor U18410 (N_18410,N_17315,N_16955);
xor U18411 (N_18411,N_17398,N_17507);
xnor U18412 (N_18412,N_17393,N_17467);
nor U18413 (N_18413,N_17201,N_17604);
nor U18414 (N_18414,N_16808,N_16989);
xor U18415 (N_18415,N_17005,N_17379);
nand U18416 (N_18416,N_17352,N_17058);
and U18417 (N_18417,N_17471,N_17256);
nand U18418 (N_18418,N_16815,N_17064);
nand U18419 (N_18419,N_17661,N_17012);
xnor U18420 (N_18420,N_17386,N_17138);
and U18421 (N_18421,N_17765,N_16840);
or U18422 (N_18422,N_17927,N_17457);
nor U18423 (N_18423,N_17650,N_17170);
nand U18424 (N_18424,N_17395,N_16856);
nand U18425 (N_18425,N_16864,N_17512);
nor U18426 (N_18426,N_17606,N_16888);
xnor U18427 (N_18427,N_17460,N_17153);
nand U18428 (N_18428,N_16916,N_17680);
nand U18429 (N_18429,N_17764,N_17872);
and U18430 (N_18430,N_17371,N_17557);
or U18431 (N_18431,N_16915,N_17653);
or U18432 (N_18432,N_16972,N_17424);
nand U18433 (N_18433,N_17933,N_17053);
nand U18434 (N_18434,N_16941,N_17868);
and U18435 (N_18435,N_17607,N_17044);
nor U18436 (N_18436,N_17269,N_17487);
and U18437 (N_18437,N_17832,N_16914);
or U18438 (N_18438,N_16918,N_17790);
or U18439 (N_18439,N_17068,N_17480);
xor U18440 (N_18440,N_17912,N_16912);
or U18441 (N_18441,N_17613,N_17826);
nor U18442 (N_18442,N_16829,N_17073);
and U18443 (N_18443,N_17351,N_16881);
and U18444 (N_18444,N_17552,N_17233);
and U18445 (N_18445,N_17830,N_17232);
nand U18446 (N_18446,N_17408,N_16929);
xor U18447 (N_18447,N_17969,N_17087);
and U18448 (N_18448,N_16865,N_16897);
or U18449 (N_18449,N_17191,N_17981);
or U18450 (N_18450,N_17939,N_17388);
and U18451 (N_18451,N_17209,N_17425);
nand U18452 (N_18452,N_17850,N_17372);
or U18453 (N_18453,N_17700,N_17788);
nand U18454 (N_18454,N_17154,N_16988);
xnor U18455 (N_18455,N_17925,N_17711);
and U18456 (N_18456,N_17644,N_17295);
xnor U18457 (N_18457,N_17978,N_17782);
and U18458 (N_18458,N_17358,N_17288);
nor U18459 (N_18459,N_17963,N_17886);
nor U18460 (N_18460,N_16837,N_17097);
and U18461 (N_18461,N_17360,N_16862);
nand U18462 (N_18462,N_17559,N_17356);
and U18463 (N_18463,N_17836,N_17775);
or U18464 (N_18464,N_16886,N_17373);
or U18465 (N_18465,N_16985,N_17062);
or U18466 (N_18466,N_17199,N_17534);
or U18467 (N_18467,N_17853,N_17858);
xnor U18468 (N_18468,N_16961,N_16825);
nor U18469 (N_18469,N_16857,N_17528);
xor U18470 (N_18470,N_17921,N_17226);
and U18471 (N_18471,N_17085,N_17478);
nand U18472 (N_18472,N_17094,N_16824);
nand U18473 (N_18473,N_17406,N_17275);
nand U18474 (N_18474,N_17121,N_17390);
or U18475 (N_18475,N_17177,N_17854);
or U18476 (N_18476,N_17046,N_17636);
nor U18477 (N_18477,N_17025,N_17570);
nand U18478 (N_18478,N_17110,N_17412);
or U18479 (N_18479,N_17056,N_16971);
nor U18480 (N_18480,N_17172,N_16938);
nor U18481 (N_18481,N_16974,N_17932);
and U18482 (N_18482,N_17683,N_17206);
and U18483 (N_18483,N_17665,N_17211);
and U18484 (N_18484,N_17964,N_17061);
or U18485 (N_18485,N_17900,N_17550);
nor U18486 (N_18486,N_17867,N_17444);
and U18487 (N_18487,N_16817,N_17795);
or U18488 (N_18488,N_17274,N_16813);
nand U18489 (N_18489,N_17586,N_17332);
nand U18490 (N_18490,N_17889,N_17493);
and U18491 (N_18491,N_17000,N_17603);
xnor U18492 (N_18492,N_17702,N_17342);
or U18493 (N_18493,N_17608,N_17376);
nor U18494 (N_18494,N_17491,N_17505);
nor U18495 (N_18495,N_17185,N_16811);
or U18496 (N_18496,N_16873,N_17321);
and U18497 (N_18497,N_17481,N_17440);
or U18498 (N_18498,N_17276,N_17791);
nor U18499 (N_18499,N_17431,N_17558);
or U18500 (N_18500,N_16842,N_17102);
nand U18501 (N_18501,N_17520,N_17792);
nor U18502 (N_18502,N_16977,N_17946);
and U18503 (N_18503,N_17466,N_17498);
nor U18504 (N_18504,N_17831,N_17554);
xor U18505 (N_18505,N_17477,N_16851);
xnor U18506 (N_18506,N_17880,N_17093);
nand U18507 (N_18507,N_17190,N_17863);
xnor U18508 (N_18508,N_17974,N_17809);
or U18509 (N_18509,N_17998,N_17846);
xnor U18510 (N_18510,N_17456,N_17822);
xor U18511 (N_18511,N_17941,N_17940);
xor U18512 (N_18512,N_17178,N_17865);
and U18513 (N_18513,N_17989,N_17229);
and U18514 (N_18514,N_17519,N_16942);
xor U18515 (N_18515,N_17002,N_17509);
xnor U18516 (N_18516,N_17824,N_17344);
and U18517 (N_18517,N_17264,N_17949);
nand U18518 (N_18518,N_17007,N_17583);
nor U18519 (N_18519,N_17689,N_17357);
and U18520 (N_18520,N_17106,N_17461);
or U18521 (N_18521,N_17414,N_16910);
xnor U18522 (N_18522,N_17637,N_17182);
nor U18523 (N_18523,N_17017,N_17086);
xor U18524 (N_18524,N_17163,N_17992);
nand U18525 (N_18525,N_17188,N_16853);
nand U18526 (N_18526,N_17286,N_16868);
nand U18527 (N_18527,N_17293,N_17237);
nand U18528 (N_18528,N_17687,N_17672);
nand U18529 (N_18529,N_17993,N_17301);
and U18530 (N_18530,N_17562,N_17984);
nor U18531 (N_18531,N_17320,N_17885);
nor U18532 (N_18532,N_17750,N_17220);
nor U18533 (N_18533,N_17287,N_17768);
nand U18534 (N_18534,N_17039,N_16810);
nand U18535 (N_18535,N_17271,N_17722);
and U18536 (N_18536,N_16908,N_17040);
xnor U18537 (N_18537,N_17909,N_17556);
nor U18538 (N_18538,N_17818,N_17479);
nand U18539 (N_18539,N_17630,N_17861);
or U18540 (N_18540,N_17359,N_17459);
or U18541 (N_18541,N_17070,N_16892);
and U18542 (N_18542,N_17935,N_17331);
and U18543 (N_18543,N_17152,N_17612);
xor U18544 (N_18544,N_17772,N_17798);
xor U18545 (N_18545,N_16852,N_16996);
or U18546 (N_18546,N_16960,N_16899);
or U18547 (N_18547,N_17279,N_17787);
and U18548 (N_18548,N_17634,N_17436);
xnor U18549 (N_18549,N_16959,N_17511);
or U18550 (N_18550,N_17219,N_17365);
nor U18551 (N_18551,N_17166,N_17323);
and U18552 (N_18552,N_17316,N_16956);
xnor U18553 (N_18553,N_17897,N_17345);
nor U18554 (N_18554,N_17259,N_17140);
xnor U18555 (N_18555,N_17956,N_17141);
and U18556 (N_18556,N_17733,N_17223);
nor U18557 (N_18557,N_17118,N_17708);
nand U18558 (N_18558,N_17881,N_17827);
nand U18559 (N_18559,N_17668,N_17036);
and U18560 (N_18560,N_17910,N_17042);
or U18561 (N_18561,N_17517,N_17476);
nor U18562 (N_18562,N_17576,N_17615);
xnor U18563 (N_18563,N_17200,N_16954);
and U18564 (N_18564,N_17533,N_17328);
or U18565 (N_18565,N_17789,N_17161);
xor U18566 (N_18566,N_16997,N_16924);
and U18567 (N_18567,N_17314,N_17463);
and U18568 (N_18568,N_17400,N_17115);
nand U18569 (N_18569,N_17510,N_16845);
nand U18570 (N_18570,N_17451,N_16946);
and U18571 (N_18571,N_17773,N_17835);
xnor U18572 (N_18572,N_16819,N_17441);
or U18573 (N_18573,N_17133,N_16800);
nand U18574 (N_18574,N_16949,N_17916);
or U18575 (N_18575,N_17258,N_17619);
and U18576 (N_18576,N_17452,N_17760);
nor U18577 (N_18577,N_17169,N_16803);
and U18578 (N_18578,N_16894,N_17540);
or U18579 (N_18579,N_17755,N_17130);
nand U18580 (N_18580,N_17857,N_17179);
or U18581 (N_18581,N_17908,N_17266);
nand U18582 (N_18582,N_17545,N_17980);
and U18583 (N_18583,N_16875,N_17943);
and U18584 (N_18584,N_17917,N_17422);
or U18585 (N_18585,N_16979,N_17139);
nor U18586 (N_18586,N_17423,N_17647);
and U18587 (N_18587,N_17146,N_17401);
xor U18588 (N_18588,N_17385,N_17631);
xnor U18589 (N_18589,N_17952,N_17531);
nor U18590 (N_18590,N_17350,N_17592);
or U18591 (N_18591,N_17745,N_17098);
nand U18592 (N_18592,N_16991,N_17777);
and U18593 (N_18593,N_17437,N_17996);
nand U18594 (N_18594,N_17438,N_17207);
or U18595 (N_18595,N_17126,N_17257);
nand U18596 (N_18596,N_17500,N_17779);
xnor U18597 (N_18597,N_17915,N_17484);
or U18598 (N_18598,N_17430,N_17922);
nand U18599 (N_18599,N_17289,N_16928);
and U18600 (N_18600,N_17672,N_17511);
nor U18601 (N_18601,N_16901,N_17906);
xor U18602 (N_18602,N_17206,N_17667);
or U18603 (N_18603,N_17579,N_17355);
and U18604 (N_18604,N_17825,N_17063);
and U18605 (N_18605,N_17967,N_17535);
and U18606 (N_18606,N_17678,N_17777);
or U18607 (N_18607,N_17919,N_17041);
xnor U18608 (N_18608,N_17545,N_17216);
nor U18609 (N_18609,N_17586,N_17036);
or U18610 (N_18610,N_17910,N_17007);
or U18611 (N_18611,N_17534,N_17834);
xor U18612 (N_18612,N_17258,N_17503);
or U18613 (N_18613,N_17707,N_17176);
xnor U18614 (N_18614,N_17985,N_16852);
nand U18615 (N_18615,N_16857,N_17467);
nor U18616 (N_18616,N_16983,N_17191);
nand U18617 (N_18617,N_17977,N_17643);
xor U18618 (N_18618,N_17859,N_17867);
nor U18619 (N_18619,N_17932,N_17988);
or U18620 (N_18620,N_17622,N_16823);
nor U18621 (N_18621,N_17634,N_17060);
xor U18622 (N_18622,N_16999,N_16844);
nand U18623 (N_18623,N_17240,N_17326);
nor U18624 (N_18624,N_17365,N_17103);
nand U18625 (N_18625,N_16861,N_17484);
nand U18626 (N_18626,N_17947,N_17106);
or U18627 (N_18627,N_17783,N_17811);
or U18628 (N_18628,N_17089,N_17674);
nor U18629 (N_18629,N_17599,N_17284);
nor U18630 (N_18630,N_16827,N_16955);
xnor U18631 (N_18631,N_17452,N_17698);
and U18632 (N_18632,N_16861,N_17089);
and U18633 (N_18633,N_17397,N_17990);
xnor U18634 (N_18634,N_17019,N_16918);
or U18635 (N_18635,N_17700,N_17961);
nand U18636 (N_18636,N_17341,N_17381);
xor U18637 (N_18637,N_17779,N_17525);
or U18638 (N_18638,N_17219,N_16850);
nor U18639 (N_18639,N_17060,N_16863);
xnor U18640 (N_18640,N_17911,N_17661);
xnor U18641 (N_18641,N_17994,N_17762);
nand U18642 (N_18642,N_17234,N_17921);
or U18643 (N_18643,N_17979,N_17374);
xnor U18644 (N_18644,N_17832,N_16858);
nor U18645 (N_18645,N_17208,N_17889);
or U18646 (N_18646,N_17079,N_17768);
or U18647 (N_18647,N_17684,N_16915);
nand U18648 (N_18648,N_17874,N_16930);
or U18649 (N_18649,N_17369,N_17750);
xor U18650 (N_18650,N_16894,N_17759);
or U18651 (N_18651,N_17126,N_17727);
and U18652 (N_18652,N_17950,N_17560);
or U18653 (N_18653,N_17206,N_17125);
and U18654 (N_18654,N_17382,N_17793);
nand U18655 (N_18655,N_17251,N_17677);
xor U18656 (N_18656,N_16893,N_17253);
nor U18657 (N_18657,N_17515,N_17901);
or U18658 (N_18658,N_17555,N_17795);
nor U18659 (N_18659,N_16894,N_17133);
xor U18660 (N_18660,N_16836,N_17941);
or U18661 (N_18661,N_17226,N_17521);
nor U18662 (N_18662,N_17739,N_17492);
or U18663 (N_18663,N_17405,N_17926);
xnor U18664 (N_18664,N_17431,N_17078);
or U18665 (N_18665,N_17922,N_17711);
and U18666 (N_18666,N_17684,N_16996);
xor U18667 (N_18667,N_17237,N_17605);
nor U18668 (N_18668,N_17133,N_16900);
nor U18669 (N_18669,N_17788,N_17777);
nor U18670 (N_18670,N_17103,N_17994);
or U18671 (N_18671,N_17847,N_17874);
or U18672 (N_18672,N_17298,N_17820);
xor U18673 (N_18673,N_17205,N_17668);
or U18674 (N_18674,N_17622,N_17077);
xnor U18675 (N_18675,N_17648,N_17623);
nor U18676 (N_18676,N_17823,N_17445);
nand U18677 (N_18677,N_17102,N_17216);
xnor U18678 (N_18678,N_17916,N_17732);
nand U18679 (N_18679,N_17572,N_17419);
xor U18680 (N_18680,N_16904,N_17455);
xnor U18681 (N_18681,N_17673,N_17143);
nand U18682 (N_18682,N_17023,N_17319);
xnor U18683 (N_18683,N_17148,N_17988);
and U18684 (N_18684,N_16904,N_17792);
xor U18685 (N_18685,N_17743,N_17138);
and U18686 (N_18686,N_16871,N_16953);
nor U18687 (N_18687,N_17419,N_17092);
or U18688 (N_18688,N_17545,N_17776);
or U18689 (N_18689,N_17149,N_17674);
and U18690 (N_18690,N_17305,N_17820);
nand U18691 (N_18691,N_16916,N_17562);
xor U18692 (N_18692,N_17416,N_17780);
nor U18693 (N_18693,N_16825,N_17107);
xnor U18694 (N_18694,N_17797,N_17863);
and U18695 (N_18695,N_17493,N_16923);
nor U18696 (N_18696,N_16902,N_17114);
nand U18697 (N_18697,N_17164,N_17566);
xnor U18698 (N_18698,N_17708,N_17310);
nor U18699 (N_18699,N_17399,N_16981);
nand U18700 (N_18700,N_17403,N_17351);
nor U18701 (N_18701,N_16930,N_17815);
nand U18702 (N_18702,N_16893,N_17745);
xnor U18703 (N_18703,N_17791,N_17831);
nor U18704 (N_18704,N_16845,N_16968);
or U18705 (N_18705,N_17170,N_17557);
xnor U18706 (N_18706,N_16938,N_17677);
or U18707 (N_18707,N_16849,N_17276);
xnor U18708 (N_18708,N_17775,N_17179);
xor U18709 (N_18709,N_17378,N_17486);
or U18710 (N_18710,N_16907,N_17099);
xor U18711 (N_18711,N_17979,N_17265);
xor U18712 (N_18712,N_16927,N_17222);
nand U18713 (N_18713,N_17997,N_17343);
xnor U18714 (N_18714,N_17830,N_17835);
nor U18715 (N_18715,N_16919,N_17673);
or U18716 (N_18716,N_17735,N_17251);
nor U18717 (N_18717,N_17595,N_16977);
and U18718 (N_18718,N_17949,N_17394);
xnor U18719 (N_18719,N_17520,N_17744);
and U18720 (N_18720,N_17459,N_17457);
xor U18721 (N_18721,N_16948,N_17985);
nor U18722 (N_18722,N_17235,N_17955);
nand U18723 (N_18723,N_16914,N_17195);
nor U18724 (N_18724,N_17201,N_17811);
and U18725 (N_18725,N_17449,N_17719);
nor U18726 (N_18726,N_17936,N_16879);
xor U18727 (N_18727,N_16904,N_17039);
nand U18728 (N_18728,N_16863,N_17172);
or U18729 (N_18729,N_17617,N_16807);
nand U18730 (N_18730,N_17021,N_16851);
nand U18731 (N_18731,N_17962,N_16840);
or U18732 (N_18732,N_17392,N_17069);
and U18733 (N_18733,N_17931,N_17412);
and U18734 (N_18734,N_17652,N_16955);
xnor U18735 (N_18735,N_17031,N_17514);
nand U18736 (N_18736,N_17680,N_17193);
nand U18737 (N_18737,N_17304,N_17623);
and U18738 (N_18738,N_17080,N_17981);
and U18739 (N_18739,N_17934,N_17335);
xor U18740 (N_18740,N_17660,N_17591);
or U18741 (N_18741,N_17792,N_17238);
nor U18742 (N_18742,N_17606,N_17192);
xnor U18743 (N_18743,N_17558,N_16844);
nor U18744 (N_18744,N_17961,N_17325);
nand U18745 (N_18745,N_17982,N_16970);
xnor U18746 (N_18746,N_17705,N_17405);
or U18747 (N_18747,N_17127,N_17557);
xnor U18748 (N_18748,N_17110,N_17055);
nand U18749 (N_18749,N_17941,N_17401);
nor U18750 (N_18750,N_17163,N_16992);
xnor U18751 (N_18751,N_17169,N_17948);
and U18752 (N_18752,N_17466,N_17360);
nor U18753 (N_18753,N_16838,N_17177);
or U18754 (N_18754,N_17381,N_17511);
or U18755 (N_18755,N_17916,N_17657);
or U18756 (N_18756,N_17386,N_17793);
and U18757 (N_18757,N_16939,N_17436);
nand U18758 (N_18758,N_17177,N_17289);
or U18759 (N_18759,N_17976,N_17301);
nand U18760 (N_18760,N_17949,N_17363);
nor U18761 (N_18761,N_17429,N_17672);
and U18762 (N_18762,N_17826,N_17416);
or U18763 (N_18763,N_17494,N_17719);
nor U18764 (N_18764,N_16876,N_17057);
nand U18765 (N_18765,N_16836,N_17756);
nand U18766 (N_18766,N_17127,N_17462);
xor U18767 (N_18767,N_17239,N_17579);
and U18768 (N_18768,N_17836,N_17690);
and U18769 (N_18769,N_17284,N_17514);
and U18770 (N_18770,N_17268,N_17064);
or U18771 (N_18771,N_17149,N_17320);
nor U18772 (N_18772,N_16969,N_17114);
xnor U18773 (N_18773,N_17368,N_17272);
nor U18774 (N_18774,N_17378,N_17386);
or U18775 (N_18775,N_17885,N_17626);
nand U18776 (N_18776,N_17568,N_17194);
and U18777 (N_18777,N_16984,N_17469);
or U18778 (N_18778,N_17487,N_17809);
nand U18779 (N_18779,N_17462,N_17748);
or U18780 (N_18780,N_16832,N_17771);
and U18781 (N_18781,N_17220,N_17678);
xnor U18782 (N_18782,N_17041,N_16835);
xnor U18783 (N_18783,N_17080,N_17609);
and U18784 (N_18784,N_17378,N_16840);
and U18785 (N_18785,N_17952,N_17007);
or U18786 (N_18786,N_17365,N_17778);
or U18787 (N_18787,N_17607,N_17728);
xor U18788 (N_18788,N_17764,N_17226);
nor U18789 (N_18789,N_17198,N_17044);
and U18790 (N_18790,N_17543,N_17610);
or U18791 (N_18791,N_17517,N_17157);
and U18792 (N_18792,N_16892,N_17347);
xnor U18793 (N_18793,N_16906,N_17494);
or U18794 (N_18794,N_17757,N_17241);
xor U18795 (N_18795,N_17833,N_17742);
or U18796 (N_18796,N_17877,N_16876);
or U18797 (N_18797,N_16859,N_17323);
and U18798 (N_18798,N_17649,N_16958);
nor U18799 (N_18799,N_17375,N_16983);
or U18800 (N_18800,N_16933,N_17444);
or U18801 (N_18801,N_17219,N_17311);
nand U18802 (N_18802,N_17117,N_17737);
or U18803 (N_18803,N_16910,N_17984);
and U18804 (N_18804,N_17441,N_17993);
nor U18805 (N_18805,N_17216,N_17609);
and U18806 (N_18806,N_17828,N_17124);
nor U18807 (N_18807,N_17429,N_16970);
nor U18808 (N_18808,N_17848,N_17592);
xor U18809 (N_18809,N_16985,N_17833);
and U18810 (N_18810,N_17713,N_17442);
nand U18811 (N_18811,N_16871,N_17298);
xnor U18812 (N_18812,N_16835,N_17155);
nand U18813 (N_18813,N_16886,N_17461);
nor U18814 (N_18814,N_17831,N_17030);
xor U18815 (N_18815,N_17293,N_17365);
and U18816 (N_18816,N_17133,N_17539);
or U18817 (N_18817,N_17725,N_16808);
nand U18818 (N_18818,N_17894,N_17649);
nor U18819 (N_18819,N_17101,N_17653);
or U18820 (N_18820,N_17599,N_17557);
and U18821 (N_18821,N_17667,N_16929);
xor U18822 (N_18822,N_17720,N_17114);
and U18823 (N_18823,N_17290,N_17293);
and U18824 (N_18824,N_17860,N_17137);
nand U18825 (N_18825,N_17557,N_17662);
xnor U18826 (N_18826,N_17996,N_17245);
nand U18827 (N_18827,N_16938,N_17407);
nor U18828 (N_18828,N_16997,N_16996);
and U18829 (N_18829,N_17555,N_16852);
xnor U18830 (N_18830,N_16974,N_17170);
and U18831 (N_18831,N_17043,N_17737);
nor U18832 (N_18832,N_17873,N_17377);
or U18833 (N_18833,N_17122,N_16997);
xor U18834 (N_18834,N_16990,N_17020);
nor U18835 (N_18835,N_17493,N_17345);
nand U18836 (N_18836,N_17635,N_17060);
and U18837 (N_18837,N_17142,N_17077);
and U18838 (N_18838,N_16906,N_17091);
or U18839 (N_18839,N_17209,N_17990);
and U18840 (N_18840,N_16828,N_17947);
or U18841 (N_18841,N_17048,N_17674);
nor U18842 (N_18842,N_17022,N_16861);
nor U18843 (N_18843,N_17511,N_16845);
or U18844 (N_18844,N_17178,N_17037);
nor U18845 (N_18845,N_17097,N_17540);
nand U18846 (N_18846,N_17044,N_17867);
xnor U18847 (N_18847,N_17288,N_17499);
xor U18848 (N_18848,N_16887,N_17998);
xor U18849 (N_18849,N_17529,N_17802);
or U18850 (N_18850,N_17789,N_16866);
or U18851 (N_18851,N_16852,N_17197);
nor U18852 (N_18852,N_16883,N_16993);
nand U18853 (N_18853,N_17038,N_16880);
nor U18854 (N_18854,N_17524,N_16887);
and U18855 (N_18855,N_17951,N_17630);
and U18856 (N_18856,N_17361,N_17606);
and U18857 (N_18857,N_17244,N_17033);
and U18858 (N_18858,N_17076,N_17769);
or U18859 (N_18859,N_17789,N_17838);
nand U18860 (N_18860,N_16961,N_16804);
and U18861 (N_18861,N_16982,N_17801);
nor U18862 (N_18862,N_17058,N_17563);
xor U18863 (N_18863,N_17530,N_17502);
nand U18864 (N_18864,N_16959,N_17410);
nand U18865 (N_18865,N_17349,N_17418);
or U18866 (N_18866,N_17841,N_17313);
or U18867 (N_18867,N_17127,N_17248);
and U18868 (N_18868,N_17550,N_17977);
nand U18869 (N_18869,N_17791,N_16845);
xnor U18870 (N_18870,N_17837,N_17876);
nand U18871 (N_18871,N_17480,N_17327);
nand U18872 (N_18872,N_17489,N_17066);
xnor U18873 (N_18873,N_17554,N_17736);
xnor U18874 (N_18874,N_17514,N_17636);
xnor U18875 (N_18875,N_17053,N_16888);
nor U18876 (N_18876,N_16939,N_17315);
or U18877 (N_18877,N_17332,N_17947);
nand U18878 (N_18878,N_17195,N_17776);
nand U18879 (N_18879,N_16988,N_17577);
nand U18880 (N_18880,N_17570,N_17981);
or U18881 (N_18881,N_17623,N_17381);
nand U18882 (N_18882,N_17055,N_17596);
or U18883 (N_18883,N_17059,N_17867);
and U18884 (N_18884,N_17571,N_17671);
nand U18885 (N_18885,N_17332,N_16836);
nor U18886 (N_18886,N_17311,N_17251);
xor U18887 (N_18887,N_17542,N_17377);
or U18888 (N_18888,N_17323,N_17295);
or U18889 (N_18889,N_17138,N_17689);
or U18890 (N_18890,N_16882,N_17055);
and U18891 (N_18891,N_17074,N_17266);
nor U18892 (N_18892,N_17403,N_17017);
nand U18893 (N_18893,N_17299,N_17776);
nor U18894 (N_18894,N_17861,N_17689);
nor U18895 (N_18895,N_16845,N_17515);
and U18896 (N_18896,N_17779,N_16880);
xor U18897 (N_18897,N_17332,N_17191);
or U18898 (N_18898,N_17365,N_17180);
nand U18899 (N_18899,N_17013,N_16848);
or U18900 (N_18900,N_17380,N_17991);
xor U18901 (N_18901,N_17565,N_17100);
or U18902 (N_18902,N_17066,N_17098);
xor U18903 (N_18903,N_17183,N_17506);
xor U18904 (N_18904,N_16873,N_17865);
nor U18905 (N_18905,N_16811,N_17301);
or U18906 (N_18906,N_17080,N_17488);
xnor U18907 (N_18907,N_17501,N_16817);
nor U18908 (N_18908,N_17322,N_17979);
nand U18909 (N_18909,N_17211,N_17097);
xor U18910 (N_18910,N_17061,N_17439);
nand U18911 (N_18911,N_17626,N_17599);
nand U18912 (N_18912,N_17359,N_17887);
and U18913 (N_18913,N_17335,N_17195);
xnor U18914 (N_18914,N_17901,N_17191);
or U18915 (N_18915,N_17620,N_17570);
or U18916 (N_18916,N_17032,N_17589);
or U18917 (N_18917,N_17598,N_17635);
nand U18918 (N_18918,N_16823,N_16854);
xor U18919 (N_18919,N_17569,N_17313);
or U18920 (N_18920,N_16928,N_17950);
and U18921 (N_18921,N_17780,N_17044);
nor U18922 (N_18922,N_17417,N_17491);
xnor U18923 (N_18923,N_17193,N_17771);
nor U18924 (N_18924,N_17732,N_17183);
nor U18925 (N_18925,N_17169,N_17138);
and U18926 (N_18926,N_17746,N_16839);
and U18927 (N_18927,N_16857,N_17164);
or U18928 (N_18928,N_17938,N_16952);
and U18929 (N_18929,N_17662,N_17571);
or U18930 (N_18930,N_16969,N_17540);
xor U18931 (N_18931,N_17422,N_17454);
and U18932 (N_18932,N_17918,N_17016);
and U18933 (N_18933,N_17135,N_17307);
nor U18934 (N_18934,N_17339,N_17906);
nand U18935 (N_18935,N_17662,N_17750);
nand U18936 (N_18936,N_16983,N_17554);
xor U18937 (N_18937,N_17231,N_17257);
nand U18938 (N_18938,N_17602,N_17221);
nand U18939 (N_18939,N_17041,N_17938);
or U18940 (N_18940,N_17539,N_17733);
nor U18941 (N_18941,N_17834,N_17582);
or U18942 (N_18942,N_17104,N_17432);
and U18943 (N_18943,N_17940,N_17620);
nand U18944 (N_18944,N_17756,N_17262);
nand U18945 (N_18945,N_16916,N_17494);
xor U18946 (N_18946,N_17352,N_17908);
nand U18947 (N_18947,N_17579,N_17893);
and U18948 (N_18948,N_17235,N_17602);
xor U18949 (N_18949,N_16856,N_17133);
xnor U18950 (N_18950,N_17110,N_17807);
nor U18951 (N_18951,N_17745,N_16902);
or U18952 (N_18952,N_17680,N_17868);
nand U18953 (N_18953,N_17069,N_17766);
nor U18954 (N_18954,N_17031,N_17851);
xor U18955 (N_18955,N_17641,N_17244);
and U18956 (N_18956,N_17528,N_16820);
or U18957 (N_18957,N_16805,N_17433);
xnor U18958 (N_18958,N_16871,N_16897);
nor U18959 (N_18959,N_17103,N_17216);
xnor U18960 (N_18960,N_16817,N_17414);
nor U18961 (N_18961,N_17687,N_16897);
nor U18962 (N_18962,N_17516,N_16910);
nor U18963 (N_18963,N_17466,N_16971);
or U18964 (N_18964,N_17054,N_17603);
nor U18965 (N_18965,N_17799,N_17562);
xor U18966 (N_18966,N_17208,N_16946);
or U18967 (N_18967,N_17641,N_17288);
nor U18968 (N_18968,N_16875,N_17751);
nand U18969 (N_18969,N_17461,N_17783);
nand U18970 (N_18970,N_17739,N_17828);
and U18971 (N_18971,N_17927,N_17374);
xor U18972 (N_18972,N_17968,N_17003);
nand U18973 (N_18973,N_17214,N_17923);
xor U18974 (N_18974,N_17156,N_17422);
nand U18975 (N_18975,N_17544,N_17423);
xnor U18976 (N_18976,N_16845,N_17570);
nor U18977 (N_18977,N_17220,N_17394);
and U18978 (N_18978,N_16886,N_17951);
nor U18979 (N_18979,N_17537,N_17476);
or U18980 (N_18980,N_16810,N_17825);
nand U18981 (N_18981,N_16824,N_16899);
nor U18982 (N_18982,N_17130,N_17391);
xor U18983 (N_18983,N_17661,N_17486);
or U18984 (N_18984,N_17079,N_16813);
or U18985 (N_18985,N_16878,N_17131);
and U18986 (N_18986,N_17518,N_17306);
or U18987 (N_18987,N_16885,N_17019);
nor U18988 (N_18988,N_16922,N_17456);
and U18989 (N_18989,N_17919,N_17990);
nand U18990 (N_18990,N_17830,N_17361);
xor U18991 (N_18991,N_16937,N_17893);
nand U18992 (N_18992,N_16900,N_17283);
or U18993 (N_18993,N_17156,N_17201);
or U18994 (N_18994,N_17318,N_17916);
and U18995 (N_18995,N_17023,N_17892);
xnor U18996 (N_18996,N_17468,N_17360);
nor U18997 (N_18997,N_16907,N_16892);
or U18998 (N_18998,N_16842,N_17728);
xnor U18999 (N_18999,N_17909,N_17207);
nand U19000 (N_19000,N_17325,N_17104);
nor U19001 (N_19001,N_17933,N_17722);
nand U19002 (N_19002,N_17209,N_17450);
and U19003 (N_19003,N_17259,N_17981);
and U19004 (N_19004,N_17535,N_17653);
or U19005 (N_19005,N_17693,N_17701);
xnor U19006 (N_19006,N_17859,N_17561);
nand U19007 (N_19007,N_17533,N_17183);
nor U19008 (N_19008,N_17056,N_17077);
xor U19009 (N_19009,N_17203,N_17149);
and U19010 (N_19010,N_17713,N_17716);
xor U19011 (N_19011,N_17241,N_16982);
and U19012 (N_19012,N_17292,N_17661);
nor U19013 (N_19013,N_17236,N_17512);
or U19014 (N_19014,N_17066,N_17688);
and U19015 (N_19015,N_17166,N_17637);
and U19016 (N_19016,N_17623,N_17457);
nand U19017 (N_19017,N_17899,N_17314);
xnor U19018 (N_19018,N_17965,N_17446);
nand U19019 (N_19019,N_17587,N_17881);
and U19020 (N_19020,N_16928,N_17270);
or U19021 (N_19021,N_17755,N_17464);
nor U19022 (N_19022,N_17557,N_17916);
xor U19023 (N_19023,N_17647,N_17418);
and U19024 (N_19024,N_17595,N_17339);
xnor U19025 (N_19025,N_17274,N_17198);
xnor U19026 (N_19026,N_17881,N_17753);
nand U19027 (N_19027,N_17420,N_17007);
nand U19028 (N_19028,N_17211,N_17463);
xnor U19029 (N_19029,N_16997,N_17370);
xnor U19030 (N_19030,N_17626,N_17847);
nor U19031 (N_19031,N_17169,N_16981);
xor U19032 (N_19032,N_17372,N_17414);
and U19033 (N_19033,N_16904,N_17390);
and U19034 (N_19034,N_17569,N_17862);
nor U19035 (N_19035,N_17158,N_17079);
xnor U19036 (N_19036,N_17659,N_16905);
or U19037 (N_19037,N_17396,N_17319);
or U19038 (N_19038,N_17865,N_16899);
and U19039 (N_19039,N_17080,N_17942);
nand U19040 (N_19040,N_16999,N_17182);
or U19041 (N_19041,N_17607,N_17434);
nor U19042 (N_19042,N_17288,N_17636);
nand U19043 (N_19043,N_17398,N_17537);
nand U19044 (N_19044,N_17768,N_17369);
nand U19045 (N_19045,N_17679,N_17597);
xnor U19046 (N_19046,N_17795,N_17510);
and U19047 (N_19047,N_17272,N_17168);
nor U19048 (N_19048,N_17454,N_17546);
nor U19049 (N_19049,N_16886,N_16949);
xor U19050 (N_19050,N_17448,N_16995);
nor U19051 (N_19051,N_16908,N_16967);
and U19052 (N_19052,N_17058,N_17822);
nor U19053 (N_19053,N_16966,N_16975);
xnor U19054 (N_19054,N_17704,N_17239);
xnor U19055 (N_19055,N_17077,N_17073);
nand U19056 (N_19056,N_17000,N_17562);
or U19057 (N_19057,N_17245,N_17929);
nor U19058 (N_19058,N_17658,N_17232);
nand U19059 (N_19059,N_17271,N_17578);
or U19060 (N_19060,N_16991,N_16894);
xnor U19061 (N_19061,N_16986,N_17127);
nand U19062 (N_19062,N_17973,N_17371);
xor U19063 (N_19063,N_17833,N_17439);
or U19064 (N_19064,N_17144,N_17507);
or U19065 (N_19065,N_17246,N_17316);
and U19066 (N_19066,N_17224,N_17758);
or U19067 (N_19067,N_17554,N_17613);
and U19068 (N_19068,N_16956,N_17371);
xor U19069 (N_19069,N_17768,N_17040);
nor U19070 (N_19070,N_17602,N_17062);
or U19071 (N_19071,N_17060,N_17002);
xor U19072 (N_19072,N_17124,N_17585);
or U19073 (N_19073,N_17160,N_17580);
nor U19074 (N_19074,N_17355,N_17746);
nand U19075 (N_19075,N_17439,N_17484);
or U19076 (N_19076,N_17496,N_17559);
nor U19077 (N_19077,N_17821,N_16946);
or U19078 (N_19078,N_17218,N_17247);
nor U19079 (N_19079,N_16829,N_17643);
and U19080 (N_19080,N_17235,N_16875);
nor U19081 (N_19081,N_17437,N_17815);
and U19082 (N_19082,N_16960,N_17158);
and U19083 (N_19083,N_16868,N_17964);
nand U19084 (N_19084,N_17157,N_17978);
and U19085 (N_19085,N_17297,N_17202);
nand U19086 (N_19086,N_17968,N_17296);
nand U19087 (N_19087,N_16929,N_16826);
xnor U19088 (N_19088,N_17409,N_17189);
or U19089 (N_19089,N_17913,N_17946);
nand U19090 (N_19090,N_17937,N_17393);
xnor U19091 (N_19091,N_17588,N_17834);
nor U19092 (N_19092,N_16961,N_17592);
and U19093 (N_19093,N_17718,N_17289);
xor U19094 (N_19094,N_17509,N_16872);
nor U19095 (N_19095,N_17099,N_17753);
and U19096 (N_19096,N_17076,N_17383);
nor U19097 (N_19097,N_17744,N_17150);
and U19098 (N_19098,N_17663,N_17664);
xor U19099 (N_19099,N_16804,N_17400);
nor U19100 (N_19100,N_17897,N_17001);
nor U19101 (N_19101,N_17061,N_17875);
or U19102 (N_19102,N_17882,N_17072);
xnor U19103 (N_19103,N_17478,N_17166);
nand U19104 (N_19104,N_17715,N_17679);
or U19105 (N_19105,N_17252,N_17630);
nand U19106 (N_19106,N_17765,N_17303);
or U19107 (N_19107,N_17555,N_17712);
or U19108 (N_19108,N_17666,N_17172);
and U19109 (N_19109,N_16857,N_17935);
nand U19110 (N_19110,N_17184,N_17202);
or U19111 (N_19111,N_17208,N_17295);
nor U19112 (N_19112,N_17055,N_17371);
or U19113 (N_19113,N_17499,N_17581);
nand U19114 (N_19114,N_17525,N_17377);
and U19115 (N_19115,N_17746,N_16869);
xor U19116 (N_19116,N_16816,N_17312);
nand U19117 (N_19117,N_17702,N_17663);
and U19118 (N_19118,N_17939,N_17004);
or U19119 (N_19119,N_17177,N_17407);
nand U19120 (N_19120,N_16950,N_17000);
nor U19121 (N_19121,N_17698,N_17336);
nor U19122 (N_19122,N_17356,N_17499);
xor U19123 (N_19123,N_16924,N_17904);
nor U19124 (N_19124,N_17381,N_17039);
nand U19125 (N_19125,N_17544,N_17621);
or U19126 (N_19126,N_16835,N_17344);
and U19127 (N_19127,N_17266,N_17793);
and U19128 (N_19128,N_17969,N_17771);
nand U19129 (N_19129,N_17567,N_17485);
or U19130 (N_19130,N_17873,N_17020);
or U19131 (N_19131,N_16901,N_17180);
or U19132 (N_19132,N_17576,N_17727);
and U19133 (N_19133,N_17471,N_17873);
or U19134 (N_19134,N_17915,N_16964);
or U19135 (N_19135,N_16968,N_17958);
or U19136 (N_19136,N_17903,N_17152);
or U19137 (N_19137,N_17178,N_17882);
xor U19138 (N_19138,N_17850,N_17933);
xnor U19139 (N_19139,N_16839,N_17652);
nand U19140 (N_19140,N_17843,N_17753);
and U19141 (N_19141,N_17263,N_17654);
nor U19142 (N_19142,N_16815,N_17301);
nor U19143 (N_19143,N_16866,N_17354);
or U19144 (N_19144,N_17942,N_16916);
nor U19145 (N_19145,N_17308,N_17001);
nand U19146 (N_19146,N_17119,N_17444);
or U19147 (N_19147,N_17021,N_17039);
and U19148 (N_19148,N_17464,N_17484);
nor U19149 (N_19149,N_17332,N_17673);
nand U19150 (N_19150,N_17623,N_17214);
xor U19151 (N_19151,N_17396,N_17184);
nor U19152 (N_19152,N_17951,N_17609);
and U19153 (N_19153,N_17713,N_17968);
or U19154 (N_19154,N_17921,N_16820);
nand U19155 (N_19155,N_16980,N_17197);
or U19156 (N_19156,N_17969,N_17857);
and U19157 (N_19157,N_17835,N_16808);
or U19158 (N_19158,N_17325,N_17607);
nor U19159 (N_19159,N_17020,N_17926);
or U19160 (N_19160,N_16977,N_17996);
nor U19161 (N_19161,N_16860,N_17759);
nor U19162 (N_19162,N_17379,N_17629);
nor U19163 (N_19163,N_16957,N_17493);
nand U19164 (N_19164,N_17321,N_17946);
or U19165 (N_19165,N_17296,N_16993);
xor U19166 (N_19166,N_17413,N_17834);
or U19167 (N_19167,N_17036,N_17795);
xor U19168 (N_19168,N_17498,N_17636);
nor U19169 (N_19169,N_17677,N_17227);
nand U19170 (N_19170,N_17862,N_17489);
and U19171 (N_19171,N_16993,N_16945);
and U19172 (N_19172,N_17477,N_17502);
and U19173 (N_19173,N_17741,N_17589);
xnor U19174 (N_19174,N_16864,N_17449);
xor U19175 (N_19175,N_17285,N_17006);
nand U19176 (N_19176,N_17251,N_17724);
nor U19177 (N_19177,N_17945,N_17770);
xnor U19178 (N_19178,N_17512,N_17994);
or U19179 (N_19179,N_16864,N_17813);
nand U19180 (N_19180,N_17297,N_17073);
xnor U19181 (N_19181,N_16934,N_16850);
or U19182 (N_19182,N_17019,N_17491);
or U19183 (N_19183,N_17222,N_17987);
nand U19184 (N_19184,N_17249,N_17292);
nor U19185 (N_19185,N_17652,N_17298);
and U19186 (N_19186,N_17303,N_17822);
xor U19187 (N_19187,N_17048,N_17741);
xnor U19188 (N_19188,N_17506,N_17682);
or U19189 (N_19189,N_17296,N_17978);
or U19190 (N_19190,N_16926,N_17946);
nand U19191 (N_19191,N_17616,N_17787);
xnor U19192 (N_19192,N_17092,N_17410);
xor U19193 (N_19193,N_17759,N_17480);
or U19194 (N_19194,N_16871,N_17003);
nand U19195 (N_19195,N_17495,N_17317);
nor U19196 (N_19196,N_17203,N_16935);
nor U19197 (N_19197,N_17876,N_17593);
or U19198 (N_19198,N_17009,N_17856);
xor U19199 (N_19199,N_17913,N_17774);
nand U19200 (N_19200,N_18307,N_18272);
xnor U19201 (N_19201,N_18814,N_18070);
or U19202 (N_19202,N_18024,N_18815);
nor U19203 (N_19203,N_18335,N_18473);
or U19204 (N_19204,N_18046,N_19027);
xor U19205 (N_19205,N_18373,N_18397);
nor U19206 (N_19206,N_18975,N_18792);
nand U19207 (N_19207,N_18704,N_18953);
or U19208 (N_19208,N_18169,N_18677);
xor U19209 (N_19209,N_18230,N_18366);
nand U19210 (N_19210,N_19047,N_18336);
nor U19211 (N_19211,N_18858,N_18487);
nand U19212 (N_19212,N_18508,N_18263);
or U19213 (N_19213,N_18740,N_18493);
and U19214 (N_19214,N_18591,N_18637);
or U19215 (N_19215,N_18352,N_19020);
nor U19216 (N_19216,N_19181,N_18795);
xnor U19217 (N_19217,N_19143,N_18678);
or U19218 (N_19218,N_18729,N_18048);
and U19219 (N_19219,N_18101,N_18471);
nor U19220 (N_19220,N_18089,N_18497);
nor U19221 (N_19221,N_18383,N_18350);
and U19222 (N_19222,N_18519,N_19040);
or U19223 (N_19223,N_18482,N_19116);
nor U19224 (N_19224,N_18430,N_18710);
nor U19225 (N_19225,N_19009,N_18153);
xnor U19226 (N_19226,N_19042,N_18833);
xnor U19227 (N_19227,N_18088,N_18159);
xor U19228 (N_19228,N_18650,N_18440);
and U19229 (N_19229,N_18539,N_18458);
and U19230 (N_19230,N_19097,N_18062);
or U19231 (N_19231,N_18364,N_19140);
and U19232 (N_19232,N_18511,N_18767);
xor U19233 (N_19233,N_18593,N_18249);
nand U19234 (N_19234,N_18402,N_18906);
or U19235 (N_19235,N_19115,N_18813);
nand U19236 (N_19236,N_18055,N_19048);
xnor U19237 (N_19237,N_19018,N_18550);
xor U19238 (N_19238,N_18128,N_18888);
nand U19239 (N_19239,N_18097,N_18433);
nor U19240 (N_19240,N_19099,N_18042);
or U19241 (N_19241,N_18047,N_18285);
nor U19242 (N_19242,N_18106,N_18974);
nand U19243 (N_19243,N_19026,N_18531);
nor U19244 (N_19244,N_18093,N_18890);
xor U19245 (N_19245,N_18573,N_18067);
or U19246 (N_19246,N_18465,N_18312);
nor U19247 (N_19247,N_18468,N_18532);
or U19248 (N_19248,N_18641,N_18713);
nand U19249 (N_19249,N_18948,N_18492);
or U19250 (N_19250,N_18469,N_18254);
nor U19251 (N_19251,N_18051,N_18321);
nand U19252 (N_19252,N_18059,N_18269);
or U19253 (N_19253,N_18859,N_19112);
nand U19254 (N_19254,N_18624,N_18739);
and U19255 (N_19255,N_18178,N_18297);
nand U19256 (N_19256,N_19182,N_18568);
and U19257 (N_19257,N_18026,N_18078);
nand U19258 (N_19258,N_18698,N_18738);
nor U19259 (N_19259,N_18001,N_18464);
xor U19260 (N_19260,N_18140,N_19141);
nor U19261 (N_19261,N_18123,N_18134);
and U19262 (N_19262,N_18775,N_18883);
nand U19263 (N_19263,N_18937,N_18176);
nor U19264 (N_19264,N_18198,N_18310);
or U19265 (N_19265,N_18594,N_19194);
nor U19266 (N_19266,N_18561,N_18645);
and U19267 (N_19267,N_19089,N_18356);
nor U19268 (N_19268,N_18011,N_18894);
nor U19269 (N_19269,N_19006,N_18248);
nand U19270 (N_19270,N_18914,N_18368);
and U19271 (N_19271,N_18590,N_18582);
or U19272 (N_19272,N_18571,N_18537);
and U19273 (N_19273,N_18455,N_18797);
and U19274 (N_19274,N_19168,N_18835);
nor U19275 (N_19275,N_18982,N_18708);
and U19276 (N_19276,N_19073,N_18292);
nor U19277 (N_19277,N_18586,N_18023);
nand U19278 (N_19278,N_18535,N_18118);
nand U19279 (N_19279,N_18395,N_18856);
nor U19280 (N_19280,N_18040,N_18862);
and U19281 (N_19281,N_18298,N_18563);
and U19282 (N_19282,N_18750,N_18077);
xor U19283 (N_19283,N_18965,N_19050);
nand U19284 (N_19284,N_18824,N_18617);
xor U19285 (N_19285,N_18060,N_18640);
nor U19286 (N_19286,N_18081,N_18562);
nand U19287 (N_19287,N_19060,N_18257);
or U19288 (N_19288,N_18278,N_18161);
and U19289 (N_19289,N_18821,N_19051);
nor U19290 (N_19290,N_18706,N_18091);
and U19291 (N_19291,N_18545,N_18449);
and U19292 (N_19292,N_18991,N_19142);
or U19293 (N_19293,N_18012,N_18733);
xnor U19294 (N_19294,N_18960,N_18502);
nor U19295 (N_19295,N_18300,N_18111);
or U19296 (N_19296,N_18661,N_19176);
nor U19297 (N_19297,N_18786,N_18341);
nand U19298 (N_19298,N_18942,N_18480);
and U19299 (N_19299,N_18674,N_18790);
xor U19300 (N_19300,N_19123,N_18208);
xnor U19301 (N_19301,N_18877,N_19064);
or U19302 (N_19302,N_18185,N_18226);
xor U19303 (N_19303,N_19052,N_19049);
and U19304 (N_19304,N_18680,N_18512);
xnor U19305 (N_19305,N_18370,N_19175);
xnor U19306 (N_19306,N_18816,N_18037);
nor U19307 (N_19307,N_18660,N_18553);
nand U19308 (N_19308,N_18918,N_18063);
nand U19309 (N_19309,N_18578,N_19127);
and U19310 (N_19310,N_18145,N_18524);
nor U19311 (N_19311,N_18486,N_18781);
or U19312 (N_19312,N_18201,N_18256);
or U19313 (N_19313,N_19013,N_18827);
xnor U19314 (N_19314,N_18453,N_18533);
or U19315 (N_19315,N_19122,N_18941);
nand U19316 (N_19316,N_18391,N_19139);
xor U19317 (N_19317,N_18907,N_18478);
xnor U19318 (N_19318,N_18901,N_18522);
xnor U19319 (N_19319,N_18569,N_18308);
xnor U19320 (N_19320,N_19164,N_18837);
or U19321 (N_19321,N_18233,N_18283);
xnor U19322 (N_19322,N_18013,N_18261);
nor U19323 (N_19323,N_18135,N_18270);
nor U19324 (N_19324,N_18943,N_18105);
nand U19325 (N_19325,N_18673,N_19184);
xnor U19326 (N_19326,N_18629,N_18425);
nor U19327 (N_19327,N_18043,N_18966);
and U19328 (N_19328,N_19120,N_18481);
xor U19329 (N_19329,N_19104,N_18782);
nand U19330 (N_19330,N_18769,N_18228);
and U19331 (N_19331,N_18005,N_18252);
and U19332 (N_19332,N_18080,N_18071);
xnor U19333 (N_19333,N_18268,N_18324);
xor U19334 (N_19334,N_18304,N_18855);
or U19335 (N_19335,N_18699,N_19171);
xnor U19336 (N_19336,N_18957,N_18371);
xor U19337 (N_19337,N_18068,N_18009);
or U19338 (N_19338,N_18191,N_19069);
and U19339 (N_19339,N_18848,N_19147);
nor U19340 (N_19340,N_19111,N_18452);
xor U19341 (N_19341,N_18838,N_18860);
or U19342 (N_19342,N_18034,N_18603);
or U19343 (N_19343,N_18404,N_18021);
or U19344 (N_19344,N_19102,N_19028);
and U19345 (N_19345,N_18853,N_18638);
or U19346 (N_19346,N_18791,N_18812);
and U19347 (N_19347,N_18273,N_18830);
xnor U19348 (N_19348,N_18551,N_18843);
and U19349 (N_19349,N_18499,N_18483);
nor U19350 (N_19350,N_18203,N_18496);
xor U19351 (N_19351,N_19088,N_18032);
xnor U19352 (N_19352,N_18224,N_18946);
or U19353 (N_19353,N_18155,N_18355);
nand U19354 (N_19354,N_18179,N_18820);
nand U19355 (N_19355,N_18672,N_18983);
or U19356 (N_19356,N_18229,N_18700);
or U19357 (N_19357,N_18994,N_19080);
nand U19358 (N_19358,N_18314,N_18489);
xnor U19359 (N_19359,N_18380,N_18065);
nand U19360 (N_19360,N_18902,N_18676);
nand U19361 (N_19361,N_18899,N_18625);
nand U19362 (N_19362,N_18150,N_18470);
and U19363 (N_19363,N_18615,N_18703);
nor U19364 (N_19364,N_18151,N_18963);
or U19365 (N_19365,N_18354,N_18845);
or U19366 (N_19366,N_19094,N_18527);
nor U19367 (N_19367,N_18258,N_19197);
and U19368 (N_19368,N_18961,N_18655);
or U19369 (N_19369,N_19173,N_18094);
nor U19370 (N_19370,N_18611,N_18969);
xor U19371 (N_19371,N_18358,N_19129);
or U19372 (N_19372,N_18851,N_18175);
nor U19373 (N_19373,N_18113,N_18944);
nand U19374 (N_19374,N_18104,N_18437);
nor U19375 (N_19375,N_19025,N_18765);
and U19376 (N_19376,N_19023,N_18211);
or U19377 (N_19377,N_18320,N_19119);
nor U19378 (N_19378,N_18474,N_18755);
xnor U19379 (N_19379,N_18548,N_19046);
and U19380 (N_19380,N_19074,N_18056);
or U19381 (N_19381,N_19004,N_19044);
xor U19382 (N_19382,N_18940,N_18751);
nor U19383 (N_19383,N_18073,N_18540);
nor U19384 (N_19384,N_18659,N_18932);
nand U19385 (N_19385,N_18521,N_18656);
or U19386 (N_19386,N_18993,N_19126);
and U19387 (N_19387,N_18086,N_18122);
nand U19388 (N_19388,N_18217,N_19188);
or U19389 (N_19389,N_18980,N_18085);
and U19390 (N_19390,N_18072,N_18694);
nor U19391 (N_19391,N_18552,N_18149);
xor U19392 (N_19392,N_18276,N_18016);
or U19393 (N_19393,N_19106,N_18780);
and U19394 (N_19394,N_19059,N_18579);
xnor U19395 (N_19395,N_18887,N_18313);
nand U19396 (N_19396,N_19014,N_18507);
nor U19397 (N_19397,N_19062,N_18014);
xnor U19398 (N_19398,N_18714,N_18082);
nor U19399 (N_19399,N_18435,N_18628);
and U19400 (N_19400,N_18744,N_18187);
and U19401 (N_19401,N_18162,N_18008);
nand U19402 (N_19402,N_18183,N_18083);
xnor U19403 (N_19403,N_18917,N_19057);
nand U19404 (N_19404,N_18018,N_18290);
and U19405 (N_19405,N_18800,N_19160);
or U19406 (N_19406,N_18280,N_18662);
nor U19407 (N_19407,N_18538,N_18536);
nor U19408 (N_19408,N_19151,N_18971);
xor U19409 (N_19409,N_18558,N_19153);
xor U19410 (N_19410,N_19183,N_18265);
or U19411 (N_19411,N_18959,N_18927);
or U19412 (N_19412,N_19086,N_18761);
nor U19413 (N_19413,N_18523,N_18041);
nand U19414 (N_19414,N_18626,N_18117);
nor U19415 (N_19415,N_18630,N_18115);
nand U19416 (N_19416,N_18984,N_18951);
nand U19417 (N_19417,N_18216,N_18864);
or U19418 (N_19418,N_18243,N_18379);
nand U19419 (N_19419,N_18096,N_19136);
or U19420 (N_19420,N_18757,N_18319);
and U19421 (N_19421,N_18362,N_18061);
or U19422 (N_19422,N_18163,N_18448);
or U19423 (N_19423,N_18172,N_18842);
nor U19424 (N_19424,N_18635,N_18876);
and U19425 (N_19425,N_18412,N_18770);
nor U19426 (N_19426,N_18495,N_19072);
and U19427 (N_19427,N_18620,N_19092);
and U19428 (N_19428,N_18367,N_18653);
nand U19429 (N_19429,N_18614,N_18107);
or U19430 (N_19430,N_18777,N_19007);
or U19431 (N_19431,N_18510,N_18166);
or U19432 (N_19432,N_18543,N_18390);
or U19433 (N_19433,N_19003,N_18618);
nand U19434 (N_19434,N_18743,N_18422);
nand U19435 (N_19435,N_18142,N_18879);
xor U19436 (N_19436,N_18409,N_18095);
or U19437 (N_19437,N_19081,N_18730);
nand U19438 (N_19438,N_19128,N_19021);
xnor U19439 (N_19439,N_18418,N_18649);
and U19440 (N_19440,N_19082,N_18520);
and U19441 (N_19441,N_18050,N_18663);
nand U19442 (N_19442,N_18337,N_18922);
nand U19443 (N_19443,N_19162,N_18567);
xnor U19444 (N_19444,N_18693,N_18330);
xor U19445 (N_19445,N_18441,N_18718);
or U19446 (N_19446,N_18587,N_18723);
nor U19447 (N_19447,N_18627,N_18873);
and U19448 (N_19448,N_19019,N_18173);
nand U19449 (N_19449,N_18881,N_18462);
nand U19450 (N_19450,N_18702,N_18664);
nand U19451 (N_19451,N_18245,N_18189);
nor U19452 (N_19452,N_18875,N_18950);
or U19453 (N_19453,N_18774,N_19087);
and U19454 (N_19454,N_19083,N_19022);
or U19455 (N_19455,N_18834,N_18803);
nand U19456 (N_19456,N_18808,N_18177);
xnor U19457 (N_19457,N_18847,N_18472);
or U19458 (N_19458,N_18728,N_18504);
and U19459 (N_19459,N_18002,N_18930);
nand U19460 (N_19460,N_18075,N_18736);
and U19461 (N_19461,N_18817,N_18326);
nand U19462 (N_19462,N_18505,N_18793);
nor U19463 (N_19463,N_18406,N_18109);
or U19464 (N_19464,N_18636,N_18724);
xor U19465 (N_19465,N_19103,N_19187);
xnor U19466 (N_19466,N_18910,N_18498);
nor U19467 (N_19467,N_18271,N_18707);
or U19468 (N_19468,N_18926,N_18799);
xnor U19469 (N_19469,N_18939,N_18976);
or U19470 (N_19470,N_18642,N_18444);
nor U19471 (N_19471,N_19002,N_18184);
xnor U19472 (N_19472,N_18334,N_19193);
nor U19473 (N_19473,N_18995,N_18160);
or U19474 (N_19474,N_18839,N_18340);
nor U19475 (N_19475,N_18732,N_18125);
nor U19476 (N_19476,N_19066,N_18076);
nor U19477 (N_19477,N_19117,N_18238);
or U19478 (N_19478,N_19031,N_18035);
or U19479 (N_19479,N_19055,N_18343);
nor U19480 (N_19480,N_18205,N_18908);
and U19481 (N_19481,N_18589,N_19156);
or U19482 (N_19482,N_18031,N_19096);
nor U19483 (N_19483,N_19155,N_18410);
nor U19484 (N_19484,N_18003,N_18281);
nand U19485 (N_19485,N_18844,N_19146);
and U19486 (N_19486,N_18675,N_18385);
or U19487 (N_19487,N_18992,N_18260);
nor U19488 (N_19488,N_18439,N_19110);
and U19489 (N_19489,N_18819,N_18904);
nor U19490 (N_19490,N_19163,N_18365);
or U19491 (N_19491,N_18981,N_18069);
nand U19492 (N_19492,N_18494,N_18116);
xor U19493 (N_19493,N_18697,N_18857);
nand U19494 (N_19494,N_18696,N_19093);
or U19495 (N_19495,N_19078,N_18180);
or U19496 (N_19496,N_18999,N_18490);
nor U19497 (N_19497,N_18604,N_18361);
xor U19498 (N_19498,N_18760,N_18333);
nand U19499 (N_19499,N_18526,N_18802);
nand U19500 (N_19500,N_18606,N_18588);
xnor U19501 (N_19501,N_19172,N_18121);
and U19502 (N_19502,N_18152,N_18949);
or U19503 (N_19503,N_18424,N_18053);
xnor U19504 (N_19504,N_19125,N_18933);
nand U19505 (N_19505,N_18514,N_19035);
nand U19506 (N_19506,N_18921,N_18779);
nand U19507 (N_19507,N_18120,N_18554);
nor U19508 (N_19508,N_18202,N_18010);
and U19509 (N_19509,N_18220,N_18204);
and U19510 (N_19510,N_18690,N_18924);
xor U19511 (N_19511,N_18099,N_19121);
and U19512 (N_19512,N_19090,N_18954);
or U19513 (N_19513,N_18234,N_18773);
and U19514 (N_19514,N_18004,N_18349);
xor U19515 (N_19515,N_18872,N_18477);
and U19516 (N_19516,N_18282,N_19012);
nor U19517 (N_19517,N_18832,N_18978);
xor U19518 (N_19518,N_18293,N_18039);
nand U19519 (N_19519,N_18616,N_18098);
nor U19520 (N_19520,N_18893,N_19079);
and U19521 (N_19521,N_18546,N_18669);
nor U19522 (N_19522,N_18193,N_18989);
or U19523 (N_19523,N_18393,N_18878);
xnor U19524 (N_19524,N_18416,N_18237);
and U19525 (N_19525,N_19076,N_18500);
and U19526 (N_19526,N_18164,N_18771);
or U19527 (N_19527,N_19058,N_18445);
or U19528 (N_19528,N_19054,N_19095);
nor U19529 (N_19529,N_18199,N_18753);
xnor U19530 (N_19530,N_18442,N_19185);
or U19531 (N_19531,N_18979,N_18219);
nor U19532 (N_19532,N_18689,N_18168);
or U19533 (N_19533,N_18811,N_18936);
nor U19534 (N_19534,N_18413,N_18749);
and U19535 (N_19535,N_18928,N_18398);
nand U19536 (N_19536,N_18619,N_18691);
nor U19537 (N_19537,N_18622,N_18846);
xor U19538 (N_19538,N_19135,N_18828);
or U19539 (N_19539,N_18905,N_19016);
nor U19540 (N_19540,N_18381,N_18332);
nor U19541 (N_19541,N_18900,N_18581);
nand U19542 (N_19542,N_18403,N_18671);
or U19543 (N_19543,N_18885,N_18264);
nand U19544 (N_19544,N_18633,N_18998);
and U19545 (N_19545,N_18392,N_18598);
or U19546 (N_19546,N_18209,N_18214);
xnor U19547 (N_19547,N_18737,N_18870);
and U19548 (N_19548,N_19170,N_19138);
or U19549 (N_19549,N_18102,N_19177);
nand U19550 (N_19550,N_18850,N_18192);
nand U19551 (N_19551,N_18267,N_18654);
or U19552 (N_19552,N_18665,N_18717);
and U19553 (N_19553,N_18131,N_18419);
and U19554 (N_19554,N_18952,N_18019);
and U19555 (N_19555,N_18207,N_18955);
or U19556 (N_19556,N_18388,N_18716);
nor U19557 (N_19557,N_18488,N_18849);
nand U19558 (N_19558,N_18503,N_18911);
and U19559 (N_19559,N_19061,N_18129);
xor U19560 (N_19560,N_18359,N_19137);
and U19561 (N_19561,N_19033,N_18171);
or U19562 (N_19562,N_18566,N_18556);
and U19563 (N_19563,N_18146,N_19100);
xnor U19564 (N_19564,N_18612,N_18124);
xnor U19565 (N_19565,N_18597,N_18829);
nand U19566 (N_19566,N_19065,N_18977);
or U19567 (N_19567,N_18913,N_18789);
and U19568 (N_19568,N_18363,N_18372);
or U19569 (N_19569,N_18734,N_18657);
nand U19570 (N_19570,N_18241,N_18181);
and U19571 (N_19571,N_18338,N_18547);
nand U19572 (N_19572,N_18647,N_19145);
or U19573 (N_19573,N_18174,N_18644);
and U19574 (N_19574,N_18938,N_18242);
nand U19575 (N_19575,N_18295,N_18064);
nand U19576 (N_19576,N_18621,N_18897);
nor U19577 (N_19577,N_18188,N_18138);
nor U19578 (N_19578,N_18294,N_18592);
and U19579 (N_19579,N_18025,N_18580);
nor U19580 (N_19580,N_18762,N_18868);
nand U19581 (N_19581,N_18218,N_18253);
and U19582 (N_19582,N_18309,N_18331);
or U19583 (N_19583,N_19154,N_18528);
xor U19584 (N_19584,N_18684,N_18892);
nor U19585 (N_19585,N_18867,N_19113);
and U19586 (N_19586,N_19053,N_18132);
nand U19587 (N_19587,N_18577,N_19008);
or U19588 (N_19588,N_18090,N_19161);
nor U19589 (N_19589,N_18206,N_18387);
xor U19590 (N_19590,N_18456,N_19131);
or U19591 (N_19591,N_19000,N_18222);
and U19592 (N_19592,N_18608,N_18414);
nand U19593 (N_19593,N_18317,N_18555);
nor U19594 (N_19594,N_18934,N_19190);
and U19595 (N_19595,N_19024,N_18017);
nand U19596 (N_19596,N_18686,N_18475);
xor U19597 (N_19597,N_18215,N_18167);
and U19598 (N_19598,N_18854,N_18079);
and U19599 (N_19599,N_19041,N_18726);
and U19600 (N_19600,N_18240,N_18599);
xor U19601 (N_19601,N_18796,N_18727);
xnor U19602 (N_19602,N_18623,N_18920);
nor U19603 (N_19603,N_18764,N_19034);
nor U19604 (N_19604,N_19075,N_18250);
and U19605 (N_19605,N_18299,N_18049);
or U19606 (N_19606,N_18666,N_18027);
and U19607 (N_19607,N_18709,N_18148);
or U19608 (N_19608,N_18668,N_18756);
nand U19609 (N_19609,N_19152,N_18156);
nor U19610 (N_19610,N_18197,N_18557);
and U19611 (N_19611,N_18423,N_18194);
nor U19612 (N_19612,N_18236,N_18329);
nor U19613 (N_19613,N_18720,N_18513);
and U19614 (N_19614,N_19108,N_18605);
or U19615 (N_19615,N_18692,N_18182);
nand U19616 (N_19616,N_18719,N_18565);
xor U19617 (N_19617,N_18251,N_18100);
nand U19618 (N_19618,N_18570,N_18575);
nand U19619 (N_19619,N_18898,N_18766);
nand U19620 (N_19620,N_19105,N_18758);
and U19621 (N_19621,N_19101,N_19144);
or U19622 (N_19622,N_18057,N_18157);
xnor U19623 (N_19623,N_18962,N_19070);
or U19624 (N_19624,N_18119,N_18327);
xnor U19625 (N_19625,N_18970,N_19077);
and U19626 (N_19626,N_18288,N_18852);
nand U19627 (N_19627,N_18609,N_19030);
and U19628 (N_19628,N_18741,N_18509);
or U19629 (N_19629,N_18103,N_18378);
nand U19630 (N_19630,N_18996,N_18136);
nand U19631 (N_19631,N_19174,N_18092);
nor U19632 (N_19632,N_19010,N_18648);
xnor U19633 (N_19633,N_18126,N_19191);
or U19634 (N_19634,N_18432,N_18600);
and U19635 (N_19635,N_18420,N_18376);
nand U19636 (N_19636,N_18431,N_18542);
or U19637 (N_19637,N_18227,N_18840);
xor U19638 (N_19638,N_18798,N_19029);
xor U19639 (N_19639,N_18342,N_19001);
and U19640 (N_19640,N_18231,N_18190);
xnor U19641 (N_19641,N_19038,N_18195);
nand U19642 (N_19642,N_18006,N_18357);
and U19643 (N_19643,N_18255,N_18968);
xnor U19644 (N_19644,N_18244,N_18772);
nand U19645 (N_19645,N_18742,N_18262);
nor U19646 (N_19646,N_18454,N_18754);
or U19647 (N_19647,N_18303,N_19039);
xnor U19648 (N_19648,N_18447,N_18515);
and U19649 (N_19649,N_19067,N_19189);
nor U19650 (N_19650,N_19037,N_18682);
nor U19651 (N_19651,N_19159,N_18595);
nand U19652 (N_19652,N_18748,N_18466);
and U19653 (N_19653,N_18054,N_18705);
nor U19654 (N_19654,N_18446,N_18344);
or U19655 (N_19655,N_18863,N_18541);
xnor U19656 (N_19656,N_18108,N_18822);
or U19657 (N_19657,N_19107,N_18912);
nor U19658 (N_19658,N_18602,N_18831);
nor U19659 (N_19659,N_18711,N_18210);
nor U19660 (N_19660,N_18158,N_18396);
and U19661 (N_19661,N_18417,N_18316);
nand U19662 (N_19662,N_18683,N_18639);
and U19663 (N_19663,N_18374,N_18200);
and U19664 (N_19664,N_18015,N_18658);
nor U19665 (N_19665,N_18865,N_19005);
and U19666 (N_19666,N_18722,N_18836);
xor U19667 (N_19667,N_18339,N_18929);
nand U19668 (N_19668,N_18916,N_18945);
nand U19669 (N_19669,N_18318,N_18052);
nor U19670 (N_19670,N_18776,N_18646);
or U19671 (N_19671,N_18461,N_18348);
nand U19672 (N_19672,N_18484,N_18323);
and U19673 (N_19673,N_18346,N_18246);
and U19674 (N_19674,N_18935,N_18130);
nor U19675 (N_19675,N_18925,N_18479);
xnor U19676 (N_19676,N_19068,N_18964);
or U19677 (N_19677,N_19158,N_18903);
xnor U19678 (N_19678,N_18020,N_18287);
nand U19679 (N_19679,N_19017,N_18634);
xor U19680 (N_19680,N_18874,N_18225);
or U19681 (N_19681,N_19045,N_19071);
nand U19682 (N_19682,N_18389,N_18601);
nor U19683 (N_19683,N_18408,N_19150);
and U19684 (N_19684,N_18377,N_18560);
and U19685 (N_19685,N_18884,N_18947);
and U19686 (N_19686,N_18576,N_18411);
xnor U19687 (N_19687,N_18029,N_18747);
and U19688 (N_19688,N_19124,N_18745);
or U19689 (N_19689,N_18559,N_18967);
nor U19690 (N_19690,N_18752,N_18141);
nor U19691 (N_19691,N_18289,N_18328);
and U19692 (N_19692,N_18405,N_18544);
and U19693 (N_19693,N_18033,N_18574);
or U19694 (N_19694,N_18667,N_18186);
and U19695 (N_19695,N_18144,N_18154);
xnor U19696 (N_19696,N_19114,N_18746);
nand U19697 (N_19697,N_19085,N_18306);
nor U19698 (N_19698,N_18074,N_18235);
nor U19699 (N_19699,N_18139,N_18030);
or U19700 (N_19700,N_19063,N_18460);
nand U19701 (N_19701,N_18768,N_18170);
xnor U19702 (N_19702,N_19056,N_19098);
or U19703 (N_19703,N_19133,N_18805);
nor U19704 (N_19704,N_19166,N_18375);
xnor U19705 (N_19705,N_18322,N_19032);
xnor U19706 (N_19706,N_18286,N_18823);
or U19707 (N_19707,N_19165,N_18818);
nand U19708 (N_19708,N_18436,N_18259);
nor U19709 (N_19709,N_18007,N_18931);
or U19710 (N_19710,N_18681,N_18221);
nor U19711 (N_19711,N_18985,N_18997);
nor U19712 (N_19712,N_18421,N_18632);
nor U19713 (N_19713,N_18787,N_19091);
nor U19714 (N_19714,N_18651,N_19148);
and U19715 (N_19715,N_19192,N_19015);
nor U19716 (N_19716,N_19157,N_18147);
and U19717 (N_19717,N_18889,N_18266);
xnor U19718 (N_19718,N_18399,N_18987);
nor U19719 (N_19719,N_18919,N_18807);
nor U19720 (N_19720,N_18973,N_18763);
or U19721 (N_19721,N_18880,N_18386);
nor U19722 (N_19722,N_18463,N_18712);
and U19723 (N_19723,N_19130,N_18806);
nand U19724 (N_19724,N_18809,N_18501);
and U19725 (N_19725,N_18701,N_19084);
or U19726 (N_19726,N_18585,N_18534);
nor U19727 (N_19727,N_19199,N_19011);
nor U19728 (N_19728,N_18296,N_18685);
nor U19729 (N_19729,N_18457,N_18516);
nor U19730 (N_19730,N_19169,N_18427);
and U19731 (N_19731,N_18794,N_18382);
and U19732 (N_19732,N_18045,N_19118);
nand U19733 (N_19733,N_18058,N_18400);
and U19734 (N_19734,N_18347,N_18788);
or U19735 (N_19735,N_19134,N_18165);
nor U19736 (N_19736,N_18459,N_18044);
and U19737 (N_19737,N_18572,N_18284);
or U19738 (N_19738,N_18429,N_18583);
or U19739 (N_19739,N_18353,N_18518);
xnor U19740 (N_19740,N_18247,N_18886);
nor U19741 (N_19741,N_18394,N_18022);
and U19742 (N_19742,N_19149,N_18909);
or U19743 (N_19743,N_18112,N_18785);
or U19744 (N_19744,N_18735,N_19198);
and U19745 (N_19745,N_18415,N_18279);
nor U19746 (N_19746,N_18360,N_19178);
nand U19747 (N_19747,N_18426,N_18110);
and U19748 (N_19748,N_18066,N_18384);
xor U19749 (N_19749,N_18613,N_18972);
and U19750 (N_19750,N_18467,N_18212);
xnor U19751 (N_19751,N_18564,N_18000);
and U19752 (N_19752,N_18784,N_18990);
nand U19753 (N_19753,N_18315,N_18407);
nor U19754 (N_19754,N_18721,N_18596);
xor U19755 (N_19755,N_18491,N_18895);
xnor U19756 (N_19756,N_19195,N_18731);
xnor U19757 (N_19757,N_19167,N_18783);
xnor U19758 (N_19758,N_19132,N_18958);
xnor U19759 (N_19759,N_18305,N_18028);
nor U19760 (N_19760,N_18778,N_18670);
nand U19761 (N_19761,N_18369,N_18438);
and U19762 (N_19762,N_18351,N_18915);
and U19763 (N_19763,N_18239,N_18825);
or U19764 (N_19764,N_19109,N_18196);
nor U19765 (N_19765,N_19036,N_18631);
xnor U19766 (N_19766,N_18274,N_19180);
xnor U19767 (N_19767,N_18302,N_18826);
nor U19768 (N_19768,N_18451,N_18804);
nor U19769 (N_19769,N_18549,N_18450);
or U19770 (N_19770,N_18127,N_18810);
and U19771 (N_19771,N_18275,N_19043);
nor U19772 (N_19772,N_18988,N_18896);
nor U19773 (N_19773,N_18143,N_18301);
and U19774 (N_19774,N_18137,N_18869);
and U19775 (N_19775,N_18801,N_18087);
xor U19776 (N_19776,N_18679,N_18506);
xor U19777 (N_19777,N_18866,N_18443);
xnor U19778 (N_19778,N_19196,N_18325);
nor U19779 (N_19779,N_18882,N_18525);
or U19780 (N_19780,N_18841,N_18476);
nand U19781 (N_19781,N_18610,N_18428);
and U19782 (N_19782,N_18725,N_18133);
or U19783 (N_19783,N_18345,N_18923);
nor U19784 (N_19784,N_18114,N_18891);
xnor U19785 (N_19785,N_18861,N_18584);
nor U19786 (N_19786,N_19179,N_18291);
nor U19787 (N_19787,N_18607,N_18232);
xnor U19788 (N_19788,N_18434,N_18277);
xnor U19789 (N_19789,N_18652,N_18643);
xnor U19790 (N_19790,N_18084,N_18986);
xor U19791 (N_19791,N_18687,N_18956);
and U19792 (N_19792,N_18213,N_18485);
xnor U19793 (N_19793,N_18517,N_18223);
or U19794 (N_19794,N_18688,N_18871);
nor U19795 (N_19795,N_18759,N_18311);
nor U19796 (N_19796,N_18036,N_18401);
and U19797 (N_19797,N_18038,N_18529);
xnor U19798 (N_19798,N_19186,N_18715);
xor U19799 (N_19799,N_18530,N_18695);
and U19800 (N_19800,N_19034,N_18314);
xor U19801 (N_19801,N_18197,N_18175);
nor U19802 (N_19802,N_19072,N_18050);
or U19803 (N_19803,N_18583,N_18815);
nand U19804 (N_19804,N_18240,N_18879);
nand U19805 (N_19805,N_18889,N_18831);
xnor U19806 (N_19806,N_18328,N_18178);
and U19807 (N_19807,N_18856,N_19022);
or U19808 (N_19808,N_18864,N_18464);
or U19809 (N_19809,N_18631,N_18352);
nor U19810 (N_19810,N_18266,N_18600);
or U19811 (N_19811,N_18559,N_18481);
xnor U19812 (N_19812,N_18411,N_19095);
and U19813 (N_19813,N_18075,N_18276);
or U19814 (N_19814,N_18627,N_18764);
and U19815 (N_19815,N_18466,N_18541);
and U19816 (N_19816,N_18849,N_18602);
and U19817 (N_19817,N_18294,N_18831);
and U19818 (N_19818,N_18284,N_18776);
nor U19819 (N_19819,N_18191,N_18441);
xor U19820 (N_19820,N_18726,N_18499);
or U19821 (N_19821,N_18992,N_18876);
and U19822 (N_19822,N_19106,N_18524);
nor U19823 (N_19823,N_18992,N_18770);
nor U19824 (N_19824,N_18353,N_18810);
or U19825 (N_19825,N_18628,N_18720);
nor U19826 (N_19826,N_18392,N_18913);
or U19827 (N_19827,N_18368,N_18174);
xor U19828 (N_19828,N_18629,N_18370);
nor U19829 (N_19829,N_19011,N_18737);
xor U19830 (N_19830,N_18541,N_18066);
xor U19831 (N_19831,N_18878,N_19096);
xnor U19832 (N_19832,N_18537,N_18457);
nand U19833 (N_19833,N_18101,N_18855);
or U19834 (N_19834,N_18573,N_18532);
nand U19835 (N_19835,N_18625,N_18130);
or U19836 (N_19836,N_19009,N_18027);
nor U19837 (N_19837,N_18029,N_18944);
xnor U19838 (N_19838,N_18489,N_18850);
or U19839 (N_19839,N_18507,N_18344);
or U19840 (N_19840,N_18921,N_18186);
or U19841 (N_19841,N_18941,N_18486);
or U19842 (N_19842,N_18211,N_18746);
nor U19843 (N_19843,N_19040,N_18564);
xor U19844 (N_19844,N_18912,N_18108);
nand U19845 (N_19845,N_18334,N_18477);
and U19846 (N_19846,N_18328,N_19139);
nand U19847 (N_19847,N_18109,N_18644);
xor U19848 (N_19848,N_18243,N_19156);
xor U19849 (N_19849,N_18211,N_18440);
xnor U19850 (N_19850,N_18899,N_18365);
or U19851 (N_19851,N_18429,N_18674);
xnor U19852 (N_19852,N_18978,N_19063);
nand U19853 (N_19853,N_18499,N_18948);
or U19854 (N_19854,N_19036,N_18683);
nand U19855 (N_19855,N_18566,N_18416);
xor U19856 (N_19856,N_19187,N_18621);
and U19857 (N_19857,N_18232,N_18703);
and U19858 (N_19858,N_19082,N_18153);
and U19859 (N_19859,N_18392,N_18544);
nor U19860 (N_19860,N_18788,N_18196);
nor U19861 (N_19861,N_18675,N_19079);
nand U19862 (N_19862,N_18554,N_19160);
or U19863 (N_19863,N_18799,N_19184);
and U19864 (N_19864,N_18347,N_18785);
nand U19865 (N_19865,N_19056,N_18319);
xor U19866 (N_19866,N_18684,N_18543);
or U19867 (N_19867,N_18670,N_18575);
xor U19868 (N_19868,N_18399,N_18247);
xnor U19869 (N_19869,N_18673,N_19196);
nand U19870 (N_19870,N_18117,N_18666);
and U19871 (N_19871,N_18774,N_18875);
and U19872 (N_19872,N_18135,N_18525);
and U19873 (N_19873,N_18390,N_18978);
and U19874 (N_19874,N_18403,N_18416);
nor U19875 (N_19875,N_18521,N_19082);
or U19876 (N_19876,N_18019,N_18824);
nand U19877 (N_19877,N_18848,N_19039);
and U19878 (N_19878,N_18154,N_19156);
nor U19879 (N_19879,N_18349,N_18214);
nor U19880 (N_19880,N_18272,N_18850);
nand U19881 (N_19881,N_18923,N_18506);
and U19882 (N_19882,N_19185,N_18150);
nor U19883 (N_19883,N_18101,N_19069);
nor U19884 (N_19884,N_18731,N_19124);
or U19885 (N_19885,N_19184,N_18642);
nand U19886 (N_19886,N_18837,N_19191);
nor U19887 (N_19887,N_18435,N_18103);
nor U19888 (N_19888,N_18479,N_18650);
nor U19889 (N_19889,N_18394,N_18424);
and U19890 (N_19890,N_19150,N_18032);
and U19891 (N_19891,N_18733,N_19168);
and U19892 (N_19892,N_18141,N_18200);
and U19893 (N_19893,N_18087,N_18188);
or U19894 (N_19894,N_18360,N_18657);
or U19895 (N_19895,N_18503,N_19199);
or U19896 (N_19896,N_18634,N_18439);
nand U19897 (N_19897,N_18420,N_18123);
and U19898 (N_19898,N_18712,N_18420);
nor U19899 (N_19899,N_18788,N_18581);
nor U19900 (N_19900,N_18071,N_18615);
nor U19901 (N_19901,N_18995,N_18475);
or U19902 (N_19902,N_18237,N_18271);
nand U19903 (N_19903,N_18077,N_18813);
nand U19904 (N_19904,N_19185,N_18206);
nand U19905 (N_19905,N_18335,N_18656);
nand U19906 (N_19906,N_19150,N_19167);
nor U19907 (N_19907,N_18611,N_18002);
nand U19908 (N_19908,N_18872,N_19121);
and U19909 (N_19909,N_18003,N_18489);
and U19910 (N_19910,N_18397,N_18161);
xor U19911 (N_19911,N_18928,N_18951);
or U19912 (N_19912,N_18408,N_18335);
nor U19913 (N_19913,N_18464,N_19001);
and U19914 (N_19914,N_18390,N_18051);
and U19915 (N_19915,N_18062,N_19089);
and U19916 (N_19916,N_18622,N_18063);
and U19917 (N_19917,N_18869,N_18854);
nor U19918 (N_19918,N_18271,N_18776);
and U19919 (N_19919,N_19150,N_18066);
and U19920 (N_19920,N_19108,N_18081);
xor U19921 (N_19921,N_18352,N_18681);
xnor U19922 (N_19922,N_18125,N_19040);
and U19923 (N_19923,N_19199,N_18542);
or U19924 (N_19924,N_18081,N_18393);
nor U19925 (N_19925,N_18545,N_19158);
xnor U19926 (N_19926,N_18394,N_19191);
and U19927 (N_19927,N_18942,N_18517);
and U19928 (N_19928,N_18079,N_19107);
xor U19929 (N_19929,N_18195,N_18770);
or U19930 (N_19930,N_18170,N_18543);
nand U19931 (N_19931,N_18327,N_18061);
nor U19932 (N_19932,N_18717,N_18224);
or U19933 (N_19933,N_18023,N_18308);
nor U19934 (N_19934,N_18048,N_18209);
nand U19935 (N_19935,N_18023,N_18941);
nand U19936 (N_19936,N_18913,N_18490);
nand U19937 (N_19937,N_19130,N_18654);
and U19938 (N_19938,N_19108,N_19001);
and U19939 (N_19939,N_18317,N_18795);
or U19940 (N_19940,N_18755,N_19143);
nand U19941 (N_19941,N_18607,N_18731);
or U19942 (N_19942,N_18384,N_19086);
or U19943 (N_19943,N_18702,N_18754);
xnor U19944 (N_19944,N_18453,N_18732);
nor U19945 (N_19945,N_18921,N_18241);
nand U19946 (N_19946,N_18737,N_18817);
and U19947 (N_19947,N_18462,N_18972);
xnor U19948 (N_19948,N_18058,N_18220);
nor U19949 (N_19949,N_18838,N_18713);
or U19950 (N_19950,N_18028,N_18580);
xor U19951 (N_19951,N_18988,N_18916);
or U19952 (N_19952,N_19037,N_18959);
xor U19953 (N_19953,N_18649,N_18992);
or U19954 (N_19954,N_18839,N_18112);
and U19955 (N_19955,N_19103,N_18178);
nor U19956 (N_19956,N_18744,N_18839);
or U19957 (N_19957,N_18878,N_18654);
nor U19958 (N_19958,N_18702,N_18629);
or U19959 (N_19959,N_18298,N_18078);
or U19960 (N_19960,N_18650,N_19157);
xnor U19961 (N_19961,N_19014,N_18945);
or U19962 (N_19962,N_18328,N_18194);
nand U19963 (N_19963,N_18626,N_18993);
nand U19964 (N_19964,N_18850,N_18152);
or U19965 (N_19965,N_18473,N_19079);
xor U19966 (N_19966,N_18342,N_18226);
or U19967 (N_19967,N_18752,N_18646);
nor U19968 (N_19968,N_18896,N_19027);
nor U19969 (N_19969,N_18939,N_19103);
or U19970 (N_19970,N_18047,N_18999);
nand U19971 (N_19971,N_18766,N_18288);
nor U19972 (N_19972,N_18536,N_18891);
xnor U19973 (N_19973,N_18096,N_18712);
nor U19974 (N_19974,N_18299,N_18082);
xnor U19975 (N_19975,N_18420,N_18071);
nor U19976 (N_19976,N_19038,N_19093);
or U19977 (N_19977,N_18827,N_18851);
and U19978 (N_19978,N_18696,N_19006);
nand U19979 (N_19979,N_18583,N_18618);
xor U19980 (N_19980,N_18290,N_18109);
nor U19981 (N_19981,N_18833,N_18154);
or U19982 (N_19982,N_19025,N_18525);
xor U19983 (N_19983,N_18205,N_19196);
xor U19984 (N_19984,N_18544,N_18782);
nand U19985 (N_19985,N_19172,N_18247);
or U19986 (N_19986,N_18424,N_18203);
or U19987 (N_19987,N_18712,N_18898);
nor U19988 (N_19988,N_18859,N_19069);
and U19989 (N_19989,N_18878,N_18193);
xnor U19990 (N_19990,N_18239,N_18103);
and U19991 (N_19991,N_18542,N_19145);
or U19992 (N_19992,N_19027,N_18336);
or U19993 (N_19993,N_18132,N_18164);
or U19994 (N_19994,N_18488,N_18266);
nand U19995 (N_19995,N_18422,N_18343);
and U19996 (N_19996,N_18778,N_18027);
or U19997 (N_19997,N_18428,N_18582);
nand U19998 (N_19998,N_19198,N_18564);
xnor U19999 (N_19999,N_18238,N_18185);
or U20000 (N_20000,N_18583,N_18238);
and U20001 (N_20001,N_19173,N_18210);
nand U20002 (N_20002,N_18231,N_18775);
nor U20003 (N_20003,N_18564,N_18603);
nand U20004 (N_20004,N_18668,N_18504);
and U20005 (N_20005,N_18201,N_18274);
xor U20006 (N_20006,N_18303,N_18345);
and U20007 (N_20007,N_18516,N_18123);
and U20008 (N_20008,N_19007,N_18403);
or U20009 (N_20009,N_18610,N_19143);
xnor U20010 (N_20010,N_18503,N_18763);
or U20011 (N_20011,N_18331,N_18250);
and U20012 (N_20012,N_18945,N_19010);
and U20013 (N_20013,N_18874,N_18905);
nor U20014 (N_20014,N_18671,N_18068);
nor U20015 (N_20015,N_18872,N_18819);
nor U20016 (N_20016,N_18402,N_18761);
xor U20017 (N_20017,N_18515,N_18092);
or U20018 (N_20018,N_18472,N_18594);
and U20019 (N_20019,N_18604,N_18028);
nor U20020 (N_20020,N_19157,N_18799);
xnor U20021 (N_20021,N_18419,N_18647);
or U20022 (N_20022,N_19098,N_18371);
xnor U20023 (N_20023,N_18975,N_18339);
nor U20024 (N_20024,N_18214,N_18660);
nor U20025 (N_20025,N_18163,N_18634);
and U20026 (N_20026,N_18536,N_18478);
nand U20027 (N_20027,N_18065,N_18492);
xnor U20028 (N_20028,N_19189,N_18375);
nand U20029 (N_20029,N_18368,N_18133);
or U20030 (N_20030,N_18924,N_18051);
xnor U20031 (N_20031,N_19079,N_18678);
nor U20032 (N_20032,N_18723,N_18222);
xnor U20033 (N_20033,N_18222,N_18233);
xor U20034 (N_20034,N_18714,N_18232);
xnor U20035 (N_20035,N_18055,N_19122);
nand U20036 (N_20036,N_18097,N_18736);
xnor U20037 (N_20037,N_18753,N_19147);
and U20038 (N_20038,N_18816,N_18168);
nand U20039 (N_20039,N_18761,N_19196);
nand U20040 (N_20040,N_18807,N_18626);
nand U20041 (N_20041,N_18173,N_18436);
and U20042 (N_20042,N_18802,N_19079);
nand U20043 (N_20043,N_18677,N_18031);
and U20044 (N_20044,N_18853,N_18630);
nand U20045 (N_20045,N_18935,N_18366);
and U20046 (N_20046,N_18044,N_18620);
and U20047 (N_20047,N_19022,N_18661);
and U20048 (N_20048,N_18402,N_18180);
and U20049 (N_20049,N_18752,N_18948);
or U20050 (N_20050,N_18164,N_19047);
xor U20051 (N_20051,N_18955,N_19036);
and U20052 (N_20052,N_18639,N_18446);
or U20053 (N_20053,N_19043,N_18542);
or U20054 (N_20054,N_19076,N_19054);
or U20055 (N_20055,N_18397,N_18492);
or U20056 (N_20056,N_18308,N_18862);
nor U20057 (N_20057,N_19091,N_18040);
and U20058 (N_20058,N_18996,N_18641);
and U20059 (N_20059,N_18665,N_18534);
and U20060 (N_20060,N_18517,N_18602);
or U20061 (N_20061,N_18435,N_18163);
nor U20062 (N_20062,N_18942,N_18345);
nand U20063 (N_20063,N_18928,N_18711);
nand U20064 (N_20064,N_18413,N_19167);
xnor U20065 (N_20065,N_19038,N_18496);
xnor U20066 (N_20066,N_18126,N_18957);
and U20067 (N_20067,N_18931,N_18728);
xnor U20068 (N_20068,N_19020,N_18367);
nor U20069 (N_20069,N_18757,N_18398);
or U20070 (N_20070,N_18850,N_18446);
or U20071 (N_20071,N_18074,N_18436);
or U20072 (N_20072,N_19046,N_19195);
xnor U20073 (N_20073,N_19106,N_18642);
nand U20074 (N_20074,N_18739,N_18009);
xnor U20075 (N_20075,N_18813,N_18526);
nand U20076 (N_20076,N_18160,N_18165);
and U20077 (N_20077,N_18346,N_18687);
nor U20078 (N_20078,N_18442,N_18567);
nand U20079 (N_20079,N_18110,N_18189);
or U20080 (N_20080,N_18077,N_18654);
nand U20081 (N_20081,N_19021,N_18610);
xor U20082 (N_20082,N_18221,N_19198);
nor U20083 (N_20083,N_18813,N_18844);
or U20084 (N_20084,N_18482,N_18371);
and U20085 (N_20085,N_18258,N_19020);
nand U20086 (N_20086,N_19036,N_18959);
xor U20087 (N_20087,N_18261,N_19120);
or U20088 (N_20088,N_18281,N_18425);
nand U20089 (N_20089,N_18070,N_18722);
nand U20090 (N_20090,N_18879,N_18288);
or U20091 (N_20091,N_18681,N_19138);
xor U20092 (N_20092,N_18797,N_18547);
and U20093 (N_20093,N_18614,N_18544);
nand U20094 (N_20094,N_18097,N_19036);
xnor U20095 (N_20095,N_18845,N_18404);
nand U20096 (N_20096,N_18673,N_19174);
nand U20097 (N_20097,N_18904,N_18845);
and U20098 (N_20098,N_18641,N_18544);
xnor U20099 (N_20099,N_18623,N_18017);
and U20100 (N_20100,N_19005,N_18516);
xnor U20101 (N_20101,N_18657,N_18153);
xnor U20102 (N_20102,N_19008,N_18985);
or U20103 (N_20103,N_18867,N_19137);
nor U20104 (N_20104,N_18399,N_18697);
nor U20105 (N_20105,N_18365,N_18787);
xnor U20106 (N_20106,N_18183,N_18136);
or U20107 (N_20107,N_18140,N_18753);
and U20108 (N_20108,N_18522,N_19180);
nor U20109 (N_20109,N_18308,N_18117);
or U20110 (N_20110,N_18195,N_18083);
nor U20111 (N_20111,N_18221,N_18380);
xnor U20112 (N_20112,N_19023,N_18632);
and U20113 (N_20113,N_18882,N_18686);
nand U20114 (N_20114,N_18075,N_18109);
nor U20115 (N_20115,N_19004,N_19038);
and U20116 (N_20116,N_18789,N_18427);
nor U20117 (N_20117,N_18904,N_18579);
nand U20118 (N_20118,N_18723,N_18449);
nand U20119 (N_20119,N_18708,N_18610);
nand U20120 (N_20120,N_18403,N_18818);
or U20121 (N_20121,N_18056,N_18222);
xor U20122 (N_20122,N_18734,N_19051);
nand U20123 (N_20123,N_18767,N_18309);
or U20124 (N_20124,N_18742,N_19149);
xor U20125 (N_20125,N_18478,N_18654);
xnor U20126 (N_20126,N_18420,N_18011);
or U20127 (N_20127,N_18064,N_18220);
and U20128 (N_20128,N_18787,N_18280);
nor U20129 (N_20129,N_18897,N_18617);
nor U20130 (N_20130,N_19192,N_18931);
and U20131 (N_20131,N_18261,N_18192);
nor U20132 (N_20132,N_19026,N_18979);
nor U20133 (N_20133,N_18065,N_18201);
xor U20134 (N_20134,N_18110,N_18248);
and U20135 (N_20135,N_19185,N_18263);
nor U20136 (N_20136,N_18724,N_18964);
nand U20137 (N_20137,N_19143,N_19053);
nor U20138 (N_20138,N_19075,N_18328);
nor U20139 (N_20139,N_18280,N_19187);
xnor U20140 (N_20140,N_18117,N_18842);
and U20141 (N_20141,N_18892,N_18569);
or U20142 (N_20142,N_18834,N_19067);
xnor U20143 (N_20143,N_19092,N_18240);
and U20144 (N_20144,N_18762,N_18382);
or U20145 (N_20145,N_19142,N_18834);
nor U20146 (N_20146,N_18672,N_19062);
nor U20147 (N_20147,N_18643,N_18488);
nor U20148 (N_20148,N_18299,N_19094);
xnor U20149 (N_20149,N_18180,N_18319);
and U20150 (N_20150,N_18727,N_19106);
or U20151 (N_20151,N_19184,N_18165);
nor U20152 (N_20152,N_18522,N_18575);
or U20153 (N_20153,N_18910,N_18475);
nor U20154 (N_20154,N_18908,N_18185);
xor U20155 (N_20155,N_18297,N_18057);
xnor U20156 (N_20156,N_18363,N_18703);
xnor U20157 (N_20157,N_18482,N_19141);
nand U20158 (N_20158,N_18066,N_18538);
or U20159 (N_20159,N_19180,N_18024);
and U20160 (N_20160,N_18547,N_19163);
nand U20161 (N_20161,N_18140,N_19058);
xnor U20162 (N_20162,N_18261,N_19074);
or U20163 (N_20163,N_19109,N_19151);
nand U20164 (N_20164,N_18405,N_18740);
and U20165 (N_20165,N_18060,N_18964);
or U20166 (N_20166,N_18034,N_19070);
or U20167 (N_20167,N_18486,N_19185);
nor U20168 (N_20168,N_18755,N_18533);
nor U20169 (N_20169,N_18016,N_18996);
nand U20170 (N_20170,N_18812,N_18796);
nand U20171 (N_20171,N_18501,N_18329);
and U20172 (N_20172,N_18632,N_18377);
and U20173 (N_20173,N_18593,N_18868);
nor U20174 (N_20174,N_18579,N_18525);
nand U20175 (N_20175,N_18074,N_18524);
nor U20176 (N_20176,N_18969,N_18143);
and U20177 (N_20177,N_18276,N_18137);
nand U20178 (N_20178,N_18202,N_18332);
xnor U20179 (N_20179,N_18151,N_18208);
nand U20180 (N_20180,N_18428,N_18832);
nand U20181 (N_20181,N_18849,N_18503);
or U20182 (N_20182,N_19103,N_18520);
or U20183 (N_20183,N_18227,N_18631);
or U20184 (N_20184,N_18619,N_18402);
nor U20185 (N_20185,N_18747,N_18713);
nor U20186 (N_20186,N_18569,N_18826);
or U20187 (N_20187,N_19070,N_18526);
and U20188 (N_20188,N_18428,N_19148);
and U20189 (N_20189,N_18491,N_18358);
nor U20190 (N_20190,N_18663,N_18960);
xor U20191 (N_20191,N_19103,N_18245);
nor U20192 (N_20192,N_18456,N_18748);
and U20193 (N_20193,N_19183,N_18500);
xnor U20194 (N_20194,N_18299,N_18690);
xnor U20195 (N_20195,N_18411,N_19157);
or U20196 (N_20196,N_18779,N_18951);
and U20197 (N_20197,N_18914,N_18929);
nand U20198 (N_20198,N_18137,N_18802);
xnor U20199 (N_20199,N_19074,N_19096);
nand U20200 (N_20200,N_18623,N_19075);
or U20201 (N_20201,N_18680,N_19140);
xor U20202 (N_20202,N_18669,N_18018);
nand U20203 (N_20203,N_18475,N_19179);
nor U20204 (N_20204,N_18452,N_18423);
and U20205 (N_20205,N_19084,N_18388);
nand U20206 (N_20206,N_18841,N_18690);
or U20207 (N_20207,N_18655,N_18306);
nor U20208 (N_20208,N_18005,N_18433);
or U20209 (N_20209,N_18465,N_18345);
xor U20210 (N_20210,N_18335,N_18162);
or U20211 (N_20211,N_18188,N_18144);
or U20212 (N_20212,N_18727,N_18296);
or U20213 (N_20213,N_18125,N_18971);
or U20214 (N_20214,N_18148,N_18934);
and U20215 (N_20215,N_18005,N_19101);
nor U20216 (N_20216,N_18731,N_18071);
xnor U20217 (N_20217,N_18891,N_19116);
xnor U20218 (N_20218,N_18071,N_18911);
nor U20219 (N_20219,N_18357,N_18700);
nor U20220 (N_20220,N_18266,N_18758);
nand U20221 (N_20221,N_18234,N_18845);
nand U20222 (N_20222,N_19084,N_18510);
or U20223 (N_20223,N_18085,N_18104);
nand U20224 (N_20224,N_18259,N_18988);
nand U20225 (N_20225,N_18725,N_18510);
xnor U20226 (N_20226,N_18182,N_18714);
and U20227 (N_20227,N_18892,N_18447);
or U20228 (N_20228,N_19007,N_19066);
xnor U20229 (N_20229,N_18134,N_18957);
xnor U20230 (N_20230,N_18218,N_18041);
nor U20231 (N_20231,N_19028,N_18121);
or U20232 (N_20232,N_19189,N_19196);
or U20233 (N_20233,N_19131,N_18883);
xnor U20234 (N_20234,N_18739,N_18207);
nor U20235 (N_20235,N_18945,N_18585);
or U20236 (N_20236,N_18123,N_19034);
nand U20237 (N_20237,N_18235,N_19015);
nor U20238 (N_20238,N_18483,N_18004);
nor U20239 (N_20239,N_18277,N_18581);
xor U20240 (N_20240,N_18660,N_18374);
and U20241 (N_20241,N_18125,N_18145);
and U20242 (N_20242,N_19045,N_18920);
nor U20243 (N_20243,N_18635,N_18309);
xnor U20244 (N_20244,N_18070,N_18011);
nor U20245 (N_20245,N_18392,N_18878);
and U20246 (N_20246,N_18444,N_18736);
nand U20247 (N_20247,N_18173,N_18314);
xnor U20248 (N_20248,N_18809,N_19150);
xnor U20249 (N_20249,N_18834,N_18963);
and U20250 (N_20250,N_18727,N_18622);
or U20251 (N_20251,N_18386,N_18115);
xnor U20252 (N_20252,N_19101,N_18255);
or U20253 (N_20253,N_18532,N_18403);
nand U20254 (N_20254,N_18328,N_19156);
xor U20255 (N_20255,N_18256,N_18143);
nand U20256 (N_20256,N_18502,N_18881);
nor U20257 (N_20257,N_18441,N_18479);
nor U20258 (N_20258,N_19157,N_18833);
and U20259 (N_20259,N_18407,N_18111);
nor U20260 (N_20260,N_18009,N_18221);
xnor U20261 (N_20261,N_18856,N_19178);
nand U20262 (N_20262,N_18709,N_18311);
nor U20263 (N_20263,N_18198,N_18616);
nor U20264 (N_20264,N_18460,N_18934);
xnor U20265 (N_20265,N_18832,N_18065);
nand U20266 (N_20266,N_18387,N_18011);
nand U20267 (N_20267,N_19021,N_18167);
nor U20268 (N_20268,N_19033,N_18900);
nor U20269 (N_20269,N_19180,N_18568);
and U20270 (N_20270,N_19135,N_19005);
nand U20271 (N_20271,N_19029,N_18927);
and U20272 (N_20272,N_18417,N_18287);
nor U20273 (N_20273,N_19131,N_18815);
nor U20274 (N_20274,N_18354,N_18343);
xor U20275 (N_20275,N_18094,N_18337);
xnor U20276 (N_20276,N_18124,N_18996);
or U20277 (N_20277,N_18544,N_18359);
and U20278 (N_20278,N_18094,N_18778);
or U20279 (N_20279,N_18238,N_18827);
and U20280 (N_20280,N_18314,N_18804);
xor U20281 (N_20281,N_18633,N_18205);
nor U20282 (N_20282,N_18362,N_18731);
xor U20283 (N_20283,N_19011,N_18541);
or U20284 (N_20284,N_18691,N_18347);
nand U20285 (N_20285,N_19008,N_18131);
nand U20286 (N_20286,N_18094,N_19069);
and U20287 (N_20287,N_18669,N_18713);
xor U20288 (N_20288,N_18454,N_18514);
nand U20289 (N_20289,N_18894,N_19193);
nand U20290 (N_20290,N_19138,N_18155);
or U20291 (N_20291,N_18321,N_19093);
or U20292 (N_20292,N_18230,N_18289);
nor U20293 (N_20293,N_18098,N_18726);
xnor U20294 (N_20294,N_19154,N_18868);
xnor U20295 (N_20295,N_18204,N_18275);
or U20296 (N_20296,N_18873,N_18058);
and U20297 (N_20297,N_19088,N_18390);
nand U20298 (N_20298,N_18552,N_18266);
nand U20299 (N_20299,N_18714,N_18535);
xor U20300 (N_20300,N_18364,N_18817);
xor U20301 (N_20301,N_18676,N_18492);
nand U20302 (N_20302,N_18823,N_19162);
nor U20303 (N_20303,N_18172,N_18337);
or U20304 (N_20304,N_19140,N_18218);
nand U20305 (N_20305,N_18907,N_18666);
xor U20306 (N_20306,N_18059,N_19111);
and U20307 (N_20307,N_18555,N_18554);
and U20308 (N_20308,N_18604,N_18896);
nand U20309 (N_20309,N_18282,N_18771);
xor U20310 (N_20310,N_18748,N_18408);
xor U20311 (N_20311,N_18976,N_18812);
nand U20312 (N_20312,N_18760,N_18521);
or U20313 (N_20313,N_18401,N_19124);
nor U20314 (N_20314,N_19168,N_18145);
nand U20315 (N_20315,N_18203,N_18228);
and U20316 (N_20316,N_18267,N_18726);
xnor U20317 (N_20317,N_18999,N_18462);
nand U20318 (N_20318,N_18944,N_18399);
nor U20319 (N_20319,N_18369,N_18312);
xor U20320 (N_20320,N_18960,N_19163);
nor U20321 (N_20321,N_18595,N_18902);
nor U20322 (N_20322,N_18660,N_18129);
nand U20323 (N_20323,N_18530,N_19059);
nor U20324 (N_20324,N_18461,N_18669);
nand U20325 (N_20325,N_18582,N_18627);
and U20326 (N_20326,N_18328,N_18657);
xor U20327 (N_20327,N_18263,N_18309);
and U20328 (N_20328,N_18547,N_18321);
nand U20329 (N_20329,N_18217,N_19111);
xor U20330 (N_20330,N_18728,N_18700);
nand U20331 (N_20331,N_18284,N_19026);
nand U20332 (N_20332,N_18202,N_18108);
and U20333 (N_20333,N_18738,N_18214);
or U20334 (N_20334,N_18061,N_19092);
or U20335 (N_20335,N_18368,N_18665);
nand U20336 (N_20336,N_18132,N_18294);
or U20337 (N_20337,N_18267,N_18731);
nand U20338 (N_20338,N_18454,N_19168);
or U20339 (N_20339,N_19176,N_18723);
nor U20340 (N_20340,N_19072,N_18906);
and U20341 (N_20341,N_18751,N_18083);
xnor U20342 (N_20342,N_18721,N_18088);
nand U20343 (N_20343,N_18847,N_18409);
and U20344 (N_20344,N_18475,N_18274);
and U20345 (N_20345,N_18348,N_19071);
nor U20346 (N_20346,N_19082,N_18196);
nor U20347 (N_20347,N_18783,N_18145);
or U20348 (N_20348,N_18451,N_18929);
xor U20349 (N_20349,N_18147,N_18171);
or U20350 (N_20350,N_18779,N_18461);
and U20351 (N_20351,N_18420,N_18135);
nand U20352 (N_20352,N_18478,N_19130);
xor U20353 (N_20353,N_19085,N_18159);
nor U20354 (N_20354,N_18895,N_18102);
xnor U20355 (N_20355,N_18097,N_18809);
and U20356 (N_20356,N_18597,N_19035);
or U20357 (N_20357,N_18788,N_18208);
nand U20358 (N_20358,N_18388,N_19069);
nand U20359 (N_20359,N_18393,N_18552);
xnor U20360 (N_20360,N_18709,N_19035);
nand U20361 (N_20361,N_19024,N_18471);
xor U20362 (N_20362,N_18558,N_18050);
and U20363 (N_20363,N_19003,N_18543);
and U20364 (N_20364,N_18424,N_18381);
and U20365 (N_20365,N_19073,N_18005);
or U20366 (N_20366,N_19168,N_18560);
nor U20367 (N_20367,N_18993,N_18938);
xor U20368 (N_20368,N_18299,N_18588);
xnor U20369 (N_20369,N_18723,N_18314);
nand U20370 (N_20370,N_18451,N_18877);
xor U20371 (N_20371,N_18485,N_18416);
or U20372 (N_20372,N_18446,N_18995);
nand U20373 (N_20373,N_19086,N_18991);
and U20374 (N_20374,N_18227,N_18914);
nor U20375 (N_20375,N_18044,N_18809);
and U20376 (N_20376,N_19195,N_18974);
nand U20377 (N_20377,N_19147,N_19035);
and U20378 (N_20378,N_18282,N_18328);
and U20379 (N_20379,N_18707,N_18302);
and U20380 (N_20380,N_19139,N_19030);
nand U20381 (N_20381,N_18729,N_18488);
nand U20382 (N_20382,N_18504,N_18872);
or U20383 (N_20383,N_18660,N_18125);
xnor U20384 (N_20384,N_18195,N_19082);
xnor U20385 (N_20385,N_18370,N_19187);
nand U20386 (N_20386,N_18820,N_19141);
nand U20387 (N_20387,N_18793,N_19068);
nand U20388 (N_20388,N_18247,N_18185);
xnor U20389 (N_20389,N_18676,N_18087);
xor U20390 (N_20390,N_18440,N_18046);
and U20391 (N_20391,N_18625,N_18960);
nand U20392 (N_20392,N_18613,N_18158);
and U20393 (N_20393,N_18411,N_18338);
nand U20394 (N_20394,N_18938,N_18059);
xor U20395 (N_20395,N_18488,N_18454);
nor U20396 (N_20396,N_19100,N_18984);
or U20397 (N_20397,N_18389,N_18241);
and U20398 (N_20398,N_18656,N_18734);
xnor U20399 (N_20399,N_18056,N_18345);
or U20400 (N_20400,N_19363,N_20069);
xor U20401 (N_20401,N_19616,N_19640);
nand U20402 (N_20402,N_20231,N_20386);
nand U20403 (N_20403,N_20011,N_19409);
nand U20404 (N_20404,N_20132,N_20047);
xnor U20405 (N_20405,N_19232,N_19690);
and U20406 (N_20406,N_19367,N_19334);
nand U20407 (N_20407,N_19327,N_19303);
or U20408 (N_20408,N_19242,N_20381);
or U20409 (N_20409,N_20064,N_19301);
and U20410 (N_20410,N_20026,N_20012);
or U20411 (N_20411,N_19673,N_19472);
xor U20412 (N_20412,N_19308,N_19651);
or U20413 (N_20413,N_20030,N_19588);
and U20414 (N_20414,N_19755,N_19699);
nand U20415 (N_20415,N_20344,N_19740);
nor U20416 (N_20416,N_20315,N_20355);
or U20417 (N_20417,N_20086,N_20188);
xor U20418 (N_20418,N_19785,N_19638);
or U20419 (N_20419,N_20345,N_20314);
nor U20420 (N_20420,N_19473,N_19375);
nand U20421 (N_20421,N_19520,N_19676);
or U20422 (N_20422,N_19280,N_20158);
and U20423 (N_20423,N_19576,N_19790);
or U20424 (N_20424,N_19979,N_20334);
xor U20425 (N_20425,N_19340,N_19641);
nand U20426 (N_20426,N_19617,N_19621);
nor U20427 (N_20427,N_19282,N_20361);
nand U20428 (N_20428,N_19749,N_19867);
xor U20429 (N_20429,N_19969,N_19729);
xor U20430 (N_20430,N_20117,N_19670);
or U20431 (N_20431,N_19335,N_19239);
nor U20432 (N_20432,N_19618,N_20294);
nor U20433 (N_20433,N_19578,N_19836);
or U20434 (N_20434,N_19201,N_19241);
xnor U20435 (N_20435,N_19684,N_19840);
or U20436 (N_20436,N_20002,N_20271);
xnor U20437 (N_20437,N_19493,N_19961);
nand U20438 (N_20438,N_19654,N_19792);
and U20439 (N_20439,N_19438,N_19696);
and U20440 (N_20440,N_19607,N_19681);
nor U20441 (N_20441,N_20096,N_19389);
or U20442 (N_20442,N_19765,N_20202);
nor U20443 (N_20443,N_20050,N_19336);
and U20444 (N_20444,N_20240,N_19310);
nor U20445 (N_20445,N_20254,N_20384);
xnor U20446 (N_20446,N_19508,N_19882);
nor U20447 (N_20447,N_20126,N_20343);
nor U20448 (N_20448,N_19933,N_20159);
nand U20449 (N_20449,N_20098,N_19397);
xnor U20450 (N_20450,N_19543,N_19581);
nor U20451 (N_20451,N_19223,N_19796);
nor U20452 (N_20452,N_20018,N_19999);
and U20453 (N_20453,N_20360,N_19539);
or U20454 (N_20454,N_20037,N_19844);
xnor U20455 (N_20455,N_20211,N_19881);
nor U20456 (N_20456,N_19260,N_19548);
xor U20457 (N_20457,N_19847,N_20264);
nor U20458 (N_20458,N_19551,N_19828);
or U20459 (N_20459,N_20010,N_20189);
xnor U20460 (N_20460,N_19626,N_19970);
nor U20461 (N_20461,N_20329,N_19276);
nand U20462 (N_20462,N_19871,N_20341);
nand U20463 (N_20463,N_19243,N_20387);
xor U20464 (N_20464,N_19876,N_19518);
nand U20465 (N_20465,N_19379,N_19939);
nor U20466 (N_20466,N_19853,N_19500);
and U20467 (N_20467,N_20125,N_20080);
and U20468 (N_20468,N_20149,N_20145);
or U20469 (N_20469,N_19787,N_20127);
or U20470 (N_20470,N_19893,N_19810);
nor U20471 (N_20471,N_20019,N_20089);
nor U20472 (N_20472,N_19622,N_20169);
or U20473 (N_20473,N_19487,N_19281);
and U20474 (N_20474,N_19982,N_19212);
nand U20475 (N_20475,N_19989,N_19325);
xor U20476 (N_20476,N_19675,N_19770);
xor U20477 (N_20477,N_19935,N_20319);
xor U20478 (N_20478,N_19877,N_19665);
nor U20479 (N_20479,N_19978,N_19800);
and U20480 (N_20480,N_20272,N_19501);
xor U20481 (N_20481,N_19863,N_19403);
nand U20482 (N_20482,N_19822,N_19304);
xnor U20483 (N_20483,N_20155,N_19658);
and U20484 (N_20484,N_19577,N_19421);
or U20485 (N_20485,N_20181,N_19407);
or U20486 (N_20486,N_19402,N_19388);
xor U20487 (N_20487,N_19290,N_19394);
nor U20488 (N_20488,N_19324,N_19595);
and U20489 (N_20489,N_19597,N_19778);
and U20490 (N_20490,N_19573,N_19716);
and U20491 (N_20491,N_19246,N_19943);
nor U20492 (N_20492,N_19783,N_20092);
or U20493 (N_20493,N_19483,N_19383);
nor U20494 (N_20494,N_19846,N_20348);
nand U20495 (N_20495,N_19444,N_20061);
nor U20496 (N_20496,N_19495,N_19488);
nor U20497 (N_20497,N_19779,N_20239);
and U20498 (N_20498,N_19255,N_20168);
xnor U20499 (N_20499,N_19951,N_19371);
xnor U20500 (N_20500,N_20337,N_19489);
and U20501 (N_20501,N_19851,N_19730);
nand U20502 (N_20502,N_19378,N_20303);
nand U20503 (N_20503,N_19464,N_20393);
nand U20504 (N_20504,N_19359,N_20325);
xnor U20505 (N_20505,N_20242,N_19479);
xnor U20506 (N_20506,N_19208,N_19793);
xor U20507 (N_20507,N_20099,N_19313);
nand U20508 (N_20508,N_20156,N_19656);
or U20509 (N_20509,N_19580,N_19429);
nor U20510 (N_20510,N_19899,N_20249);
nand U20511 (N_20511,N_19385,N_20114);
nand U20512 (N_20512,N_20213,N_19680);
nand U20513 (N_20513,N_19975,N_20015);
or U20514 (N_20514,N_19249,N_19467);
or U20515 (N_20515,N_19251,N_19774);
nand U20516 (N_20516,N_19902,N_20200);
and U20517 (N_20517,N_20196,N_19226);
nand U20518 (N_20518,N_20038,N_20235);
or U20519 (N_20519,N_19620,N_19210);
nand U20520 (N_20520,N_20215,N_19672);
and U20521 (N_20521,N_20136,N_19372);
xnor U20522 (N_20522,N_19806,N_19235);
xnor U20523 (N_20523,N_19669,N_19504);
xor U20524 (N_20524,N_19914,N_19315);
and U20525 (N_20525,N_19756,N_19752);
xnor U20526 (N_20526,N_20265,N_19590);
nor U20527 (N_20527,N_20005,N_20372);
and U20528 (N_20528,N_20287,N_20142);
and U20529 (N_20529,N_19406,N_19530);
and U20530 (N_20530,N_19491,N_19405);
xnor U20531 (N_20531,N_20238,N_19203);
or U20532 (N_20532,N_19744,N_19652);
and U20533 (N_20533,N_19305,N_19995);
and U20534 (N_20534,N_20317,N_19717);
nor U20535 (N_20535,N_19627,N_19857);
and U20536 (N_20536,N_20116,N_19370);
nor U20537 (N_20537,N_20301,N_20305);
nand U20538 (N_20538,N_20129,N_19206);
xnor U20539 (N_20539,N_19554,N_19459);
and U20540 (N_20540,N_19237,N_19984);
xor U20541 (N_20541,N_19994,N_19368);
xor U20542 (N_20542,N_19601,N_20346);
and U20543 (N_20543,N_19482,N_20109);
and U20544 (N_20544,N_19814,N_20100);
nor U20545 (N_20545,N_20173,N_20003);
nor U20546 (N_20546,N_19811,N_19525);
nor U20547 (N_20547,N_20042,N_19695);
or U20548 (N_20548,N_19916,N_20212);
or U20549 (N_20549,N_20302,N_20163);
nand U20550 (N_20550,N_20363,N_19683);
nor U20551 (N_20551,N_19529,N_20322);
nand U20552 (N_20552,N_20201,N_19706);
and U20553 (N_20553,N_20152,N_20359);
xor U20554 (N_20554,N_20261,N_19874);
nor U20555 (N_20555,N_19436,N_20347);
or U20556 (N_20556,N_19326,N_19927);
xnor U20557 (N_20557,N_20021,N_20110);
nor U20558 (N_20558,N_20377,N_19637);
and U20559 (N_20559,N_19231,N_19538);
or U20560 (N_20560,N_20093,N_19748);
nor U20561 (N_20561,N_20247,N_19718);
or U20562 (N_20562,N_20192,N_19751);
xnor U20563 (N_20563,N_19789,N_20321);
and U20564 (N_20564,N_19647,N_19702);
xnor U20565 (N_20565,N_19870,N_19498);
and U20566 (N_20566,N_20318,N_19380);
nand U20567 (N_20567,N_20139,N_19445);
and U20568 (N_20568,N_19583,N_19587);
or U20569 (N_20569,N_19950,N_19250);
and U20570 (N_20570,N_19945,N_19600);
nand U20571 (N_20571,N_20198,N_19780);
and U20572 (N_20572,N_19991,N_19289);
xor U20573 (N_20573,N_20107,N_19968);
xor U20574 (N_20574,N_19760,N_20310);
nor U20575 (N_20575,N_19211,N_19434);
nor U20576 (N_20576,N_20079,N_19430);
nand U20577 (N_20577,N_20216,N_20101);
nor U20578 (N_20578,N_20282,N_20224);
and U20579 (N_20579,N_19906,N_19485);
and U20580 (N_20580,N_19817,N_19492);
and U20581 (N_20581,N_20326,N_19966);
xnor U20582 (N_20582,N_20180,N_19563);
or U20583 (N_20583,N_20274,N_19410);
or U20584 (N_20584,N_19514,N_19294);
and U20585 (N_20585,N_19727,N_19602);
nand U20586 (N_20586,N_20394,N_19471);
or U20587 (N_20587,N_19350,N_19738);
xor U20588 (N_20588,N_19511,N_19609);
nand U20589 (N_20589,N_19781,N_20095);
nor U20590 (N_20590,N_20185,N_19664);
nand U20591 (N_20591,N_20000,N_19688);
nand U20592 (N_20592,N_20046,N_20122);
or U20593 (N_20593,N_19455,N_20245);
nor U20594 (N_20594,N_19366,N_19777);
nor U20595 (N_20595,N_20225,N_19446);
and U20596 (N_20596,N_19798,N_19413);
and U20597 (N_20597,N_19465,N_19424);
or U20598 (N_20598,N_19582,N_20327);
nand U20599 (N_20599,N_20278,N_19234);
nand U20600 (N_20600,N_19428,N_19829);
and U20601 (N_20601,N_19293,N_20074);
or U20602 (N_20602,N_19956,N_20062);
or U20603 (N_20603,N_19229,N_20285);
and U20604 (N_20604,N_20141,N_20124);
xnor U20605 (N_20605,N_19432,N_20164);
and U20606 (N_20606,N_19894,N_19924);
nor U20607 (N_20607,N_19506,N_19571);
and U20608 (N_20608,N_19599,N_20260);
and U20609 (N_20609,N_19905,N_19722);
nor U20610 (N_20610,N_19624,N_19767);
xnor U20611 (N_20611,N_20090,N_20277);
or U20612 (N_20612,N_19457,N_19929);
and U20613 (N_20613,N_20056,N_19476);
and U20614 (N_20614,N_19864,N_19946);
or U20615 (N_20615,N_20320,N_19723);
or U20616 (N_20616,N_19395,N_19821);
or U20617 (N_20617,N_19425,N_19784);
or U20618 (N_20618,N_19944,N_19998);
or U20619 (N_20619,N_20053,N_19941);
xnor U20620 (N_20620,N_19655,N_19630);
xnor U20621 (N_20621,N_20258,N_20121);
nor U20622 (N_20622,N_19295,N_19805);
nand U20623 (N_20623,N_20082,N_19981);
nand U20624 (N_20624,N_19328,N_19861);
nand U20625 (N_20625,N_19236,N_19297);
nand U20626 (N_20626,N_19570,N_20177);
and U20627 (N_20627,N_20267,N_19856);
xor U20628 (N_20628,N_20025,N_19801);
or U20629 (N_20629,N_19608,N_19419);
xor U20630 (N_20630,N_20256,N_19463);
or U20631 (N_20631,N_19919,N_19558);
xnor U20632 (N_20632,N_20352,N_19412);
and U20633 (N_20633,N_19568,N_19386);
and U20634 (N_20634,N_20076,N_20383);
and U20635 (N_20635,N_19537,N_19947);
xnor U20636 (N_20636,N_20229,N_19786);
nor U20637 (N_20637,N_20299,N_19224);
xor U20638 (N_20638,N_19408,N_19967);
nand U20639 (N_20639,N_19272,N_20203);
nand U20640 (N_20640,N_19948,N_19362);
xor U20641 (N_20641,N_19593,N_19973);
nand U20642 (N_20642,N_20246,N_19866);
nand U20643 (N_20643,N_19341,N_19753);
nor U20644 (N_20644,N_19598,N_19709);
nand U20645 (N_20645,N_19938,N_20108);
xor U20646 (N_20646,N_19625,N_19277);
nand U20647 (N_20647,N_19648,N_19585);
nor U20648 (N_20648,N_20342,N_19332);
nand U20649 (N_20649,N_19400,N_19261);
nand U20650 (N_20650,N_19339,N_19816);
nor U20651 (N_20651,N_20051,N_19725);
xor U20652 (N_20652,N_20307,N_19831);
or U20653 (N_20653,N_19567,N_20378);
or U20654 (N_20654,N_20392,N_20066);
and U20655 (N_20655,N_20388,N_20028);
nor U20656 (N_20656,N_20123,N_19536);
xor U20657 (N_20657,N_19468,N_19960);
nor U20658 (N_20658,N_19992,N_19497);
or U20659 (N_20659,N_19420,N_19505);
xnor U20660 (N_20660,N_19639,N_19515);
or U20661 (N_20661,N_20281,N_19976);
and U20662 (N_20662,N_19782,N_19565);
nand U20663 (N_20663,N_20205,N_19264);
nand U20664 (N_20664,N_19480,N_19912);
or U20665 (N_20665,N_20370,N_19374);
and U20666 (N_20666,N_19643,N_19671);
nor U20667 (N_20667,N_20134,N_19592);
xnor U20668 (N_20668,N_19214,N_19746);
nand U20669 (N_20669,N_20353,N_19742);
nor U20670 (N_20670,N_19823,N_19309);
xnor U20671 (N_20671,N_19762,N_19605);
and U20672 (N_20672,N_19202,N_19757);
nor U20673 (N_20673,N_19776,N_19841);
and U20674 (N_20674,N_19584,N_19298);
xnor U20675 (N_20675,N_19721,N_20362);
or U20676 (N_20676,N_19963,N_20244);
nand U20677 (N_20677,N_19908,N_19330);
and U20678 (N_20678,N_19815,N_19833);
or U20679 (N_20679,N_20286,N_20255);
xor U20680 (N_20680,N_20014,N_19606);
nor U20681 (N_20681,N_19628,N_20350);
xnor U20682 (N_20682,N_19553,N_19878);
nor U20683 (N_20683,N_19311,N_19443);
and U20684 (N_20684,N_19775,N_19830);
xnor U20685 (N_20685,N_19707,N_19435);
and U20686 (N_20686,N_20029,N_19353);
xnor U20687 (N_20687,N_20300,N_20036);
or U20688 (N_20688,N_19270,N_19342);
nand U20689 (N_20689,N_20374,N_19766);
nor U20690 (N_20690,N_20330,N_20219);
and U20691 (N_20691,N_19256,N_19314);
nor U20692 (N_20692,N_20041,N_19418);
xor U20693 (N_20693,N_19439,N_19238);
and U20694 (N_20694,N_19347,N_20222);
or U20695 (N_20695,N_19644,N_20071);
xnor U20696 (N_20696,N_19306,N_19209);
nand U20697 (N_20697,N_19269,N_20087);
nor U20698 (N_20698,N_20351,N_20376);
or U20699 (N_20699,N_19322,N_20073);
xnor U20700 (N_20700,N_20338,N_19254);
xnor U20701 (N_20701,N_20221,N_19678);
xor U20702 (N_20702,N_19897,N_20223);
and U20703 (N_20703,N_19858,N_19736);
and U20704 (N_20704,N_19855,N_19391);
nor U20705 (N_20705,N_20228,N_19426);
xnor U20706 (N_20706,N_19512,N_20335);
nand U20707 (N_20707,N_19804,N_19885);
or U20708 (N_20708,N_19319,N_19977);
nand U20709 (N_20709,N_19411,N_20054);
xnor U20710 (N_20710,N_20251,N_19358);
xor U20711 (N_20711,N_19575,N_19503);
or U20712 (N_20712,N_20369,N_19631);
nand U20713 (N_20713,N_19926,N_20263);
and U20714 (N_20714,N_19925,N_19453);
or U20715 (N_20715,N_19845,N_19292);
xor U20716 (N_20716,N_19523,N_20072);
xor U20717 (N_20717,N_20308,N_20398);
and U20718 (N_20718,N_20140,N_19594);
nand U20719 (N_20719,N_19441,N_20232);
xnor U20720 (N_20720,N_19741,N_19527);
or U20721 (N_20721,N_19259,N_20133);
or U20722 (N_20722,N_19552,N_19803);
xnor U20723 (N_20723,N_19771,N_20153);
and U20724 (N_20724,N_19531,N_19974);
and U20725 (N_20725,N_19824,N_19450);
or U20726 (N_20726,N_19291,N_20027);
nand U20727 (N_20727,N_20316,N_20375);
and U20728 (N_20728,N_20128,N_20312);
and U20729 (N_20729,N_19909,N_20234);
xnor U20730 (N_20730,N_20217,N_20328);
nand U20731 (N_20731,N_20382,N_19940);
or U20732 (N_20732,N_20389,N_20017);
nand U20733 (N_20733,N_19398,N_19275);
nand U20734 (N_20734,N_19884,N_19228);
nor U20735 (N_20735,N_19603,N_19839);
and U20736 (N_20736,N_20022,N_19623);
xnor U20737 (N_20737,N_20118,N_19686);
and U20738 (N_20738,N_20333,N_20016);
nor U20739 (N_20739,N_20137,N_19392);
nor U20740 (N_20740,N_19888,N_20004);
nor U20741 (N_20741,N_19710,N_20236);
or U20742 (N_20742,N_19509,N_19456);
and U20743 (N_20743,N_19393,N_19333);
and U20744 (N_20744,N_19555,N_20008);
and U20745 (N_20745,N_20191,N_20237);
and U20746 (N_20746,N_20077,N_20395);
nor U20747 (N_20747,N_20120,N_19891);
nor U20748 (N_20748,N_19962,N_19859);
nand U20749 (N_20749,N_20357,N_19703);
and U20750 (N_20750,N_19448,N_19896);
xor U20751 (N_20751,N_20257,N_19376);
and U20752 (N_20752,N_19691,N_19221);
nand U20753 (N_20753,N_19451,N_19542);
nand U20754 (N_20754,N_19461,N_19470);
nand U20755 (N_20755,N_19460,N_19474);
or U20756 (N_20756,N_20060,N_20033);
and U20757 (N_20757,N_19615,N_19835);
xnor U20758 (N_20758,N_19533,N_19910);
nand U20759 (N_20759,N_19307,N_19838);
and U20760 (N_20760,N_19633,N_19317);
nor U20761 (N_20761,N_19701,N_19343);
nand U20762 (N_20762,N_19337,N_19355);
xnor U20763 (N_20763,N_19452,N_19484);
xor U20764 (N_20764,N_19708,N_20035);
xnor U20765 (N_20765,N_20144,N_19613);
or U20766 (N_20766,N_19666,N_19930);
xnor U20767 (N_20767,N_19879,N_19954);
xnor U20768 (N_20768,N_20193,N_19204);
or U20769 (N_20769,N_20354,N_20070);
xor U20770 (N_20770,N_19502,N_19689);
or U20771 (N_20771,N_19271,N_19399);
nor U20772 (N_20772,N_19218,N_20266);
and U20773 (N_20773,N_19850,N_19352);
or U20774 (N_20774,N_20009,N_20323);
xor U20775 (N_20775,N_19528,N_19566);
xor U20776 (N_20776,N_19257,N_20206);
and U20777 (N_20777,N_19387,N_19612);
and U20778 (N_20778,N_19714,N_19918);
or U20779 (N_20779,N_20289,N_20367);
xor U20780 (N_20780,N_20218,N_19478);
or U20781 (N_20781,N_19754,N_19263);
nor U20782 (N_20782,N_19667,N_19225);
or U20783 (N_20783,N_20296,N_19219);
xor U20784 (N_20784,N_19813,N_19917);
or U20785 (N_20785,N_19384,N_20262);
nand U20786 (N_20786,N_20045,N_20365);
nand U20787 (N_20787,N_20088,N_19296);
and U20788 (N_20788,N_20293,N_19579);
or U20789 (N_20789,N_19915,N_19959);
and U20790 (N_20790,N_20270,N_19732);
and U20791 (N_20791,N_19820,N_19610);
or U20792 (N_20792,N_20063,N_19807);
and U20793 (N_20793,N_19494,N_19556);
xor U20794 (N_20794,N_19344,N_20055);
xnor U20795 (N_20795,N_19284,N_19769);
nor U20796 (N_20796,N_19526,N_19901);
or U20797 (N_20797,N_19300,N_19278);
nand U20798 (N_20798,N_19283,N_20368);
and U20799 (N_20799,N_19390,N_19247);
nand U20800 (N_20800,N_19705,N_20052);
and U20801 (N_20801,N_19205,N_19517);
or U20802 (N_20802,N_19636,N_20176);
nand U20803 (N_20803,N_19988,N_20150);
nor U20804 (N_20804,N_19745,N_19869);
and U20805 (N_20805,N_20194,N_19739);
nor U20806 (N_20806,N_19589,N_20085);
and U20807 (N_20807,N_19466,N_20184);
or U20808 (N_20808,N_20166,N_19507);
and U20809 (N_20809,N_20183,N_19832);
xor U20810 (N_20810,N_20208,N_20143);
xnor U20811 (N_20811,N_19791,N_19713);
or U20812 (N_20812,N_19734,N_19351);
nand U20813 (N_20813,N_19662,N_20044);
nor U20814 (N_20814,N_19697,N_20031);
or U20815 (N_20815,N_20336,N_20001);
xor U20816 (N_20816,N_19416,N_20364);
or U20817 (N_20817,N_20146,N_19299);
nand U20818 (N_20818,N_19726,N_19724);
nor U20819 (N_20819,N_19486,N_19320);
and U20820 (N_20820,N_19475,N_19852);
or U20821 (N_20821,N_19213,N_20112);
nor U20822 (N_20822,N_19516,N_19875);
xnor U20823 (N_20823,N_20174,N_19848);
nand U20824 (N_20824,N_19761,N_19377);
nand U20825 (N_20825,N_19922,N_19904);
or U20826 (N_20826,N_20324,N_19733);
nor U20827 (N_20827,N_19937,N_19913);
nor U20828 (N_20828,N_19818,N_20160);
or U20829 (N_20829,N_20340,N_19728);
nor U20830 (N_20830,N_19715,N_19510);
or U20831 (N_20831,N_19381,N_19653);
nor U20832 (N_20832,N_20298,N_19427);
and U20833 (N_20833,N_20253,N_19442);
nor U20834 (N_20834,N_20280,N_19361);
and U20835 (N_20835,N_20131,N_19996);
nand U20836 (N_20836,N_20304,N_19849);
and U20837 (N_20837,N_19862,N_20356);
and U20838 (N_20838,N_19712,N_19354);
nor U20839 (N_20839,N_20250,N_19700);
and U20840 (N_20840,N_20040,N_19302);
and U20841 (N_20841,N_19704,N_19980);
nor U20842 (N_20842,N_20175,N_20306);
and U20843 (N_20843,N_20339,N_20048);
and U20844 (N_20844,N_19860,N_20102);
or U20845 (N_20845,N_20162,N_20391);
or U20846 (N_20846,N_19266,N_19809);
nor U20847 (N_20847,N_20259,N_19596);
and U20848 (N_20848,N_19288,N_19635);
nor U20849 (N_20849,N_19279,N_20268);
nand U20850 (N_20850,N_19329,N_20113);
nand U20851 (N_20851,N_20366,N_19604);
and U20852 (N_20852,N_20248,N_20288);
nand U20853 (N_20853,N_19216,N_20199);
or U20854 (N_20854,N_20275,N_19997);
nand U20855 (N_20855,N_19663,N_19356);
nand U20856 (N_20856,N_20013,N_20230);
xnor U20857 (N_20857,N_19253,N_20243);
or U20858 (N_20858,N_20078,N_19668);
nor U20859 (N_20859,N_20309,N_19903);
and U20860 (N_20860,N_19369,N_19660);
nand U20861 (N_20861,N_19462,N_20097);
nand U20862 (N_20862,N_20380,N_19719);
nor U20863 (N_20863,N_19795,N_19481);
nand U20864 (N_20864,N_20034,N_19346);
or U20865 (N_20865,N_19957,N_20103);
nand U20866 (N_20866,N_19768,N_19634);
or U20867 (N_20867,N_20130,N_19540);
and U20868 (N_20868,N_19262,N_19572);
nor U20869 (N_20869,N_19422,N_19569);
or U20870 (N_20870,N_19447,N_20138);
xnor U20871 (N_20871,N_19928,N_19687);
xor U20872 (N_20872,N_19611,N_19711);
nand U20873 (N_20873,N_20178,N_20220);
nor U20874 (N_20874,N_19348,N_19985);
xnor U20875 (N_20875,N_19972,N_20279);
or U20876 (N_20876,N_20195,N_19971);
or U20877 (N_20877,N_19396,N_19797);
nor U20878 (N_20878,N_20227,N_19345);
nand U20879 (N_20879,N_19477,N_20115);
nand U20880 (N_20880,N_20241,N_20332);
nand U20881 (N_20881,N_20081,N_19258);
xnor U20882 (N_20882,N_19230,N_19524);
and U20883 (N_20883,N_19513,N_19758);
xnor U20884 (N_20884,N_19574,N_19535);
and U20885 (N_20885,N_20358,N_19887);
or U20886 (N_20886,N_19731,N_20371);
nand U20887 (N_20887,N_19316,N_19215);
or U20888 (N_20888,N_19349,N_20399);
or U20889 (N_20889,N_20154,N_19331);
nor U20890 (N_20890,N_20059,N_19222);
or U20891 (N_20891,N_19240,N_19321);
nor U20892 (N_20892,N_20067,N_19949);
xnor U20893 (N_20893,N_19433,N_19562);
xnor U20894 (N_20894,N_19401,N_19458);
or U20895 (N_20895,N_20204,N_20390);
nand U20896 (N_20896,N_19287,N_19440);
and U20897 (N_20897,N_19469,N_19936);
or U20898 (N_20898,N_20167,N_19872);
and U20899 (N_20899,N_19990,N_19759);
xnor U20900 (N_20900,N_19534,N_19364);
nor U20901 (N_20901,N_19265,N_19496);
xnor U20902 (N_20902,N_19747,N_19318);
and U20903 (N_20903,N_20058,N_19642);
nor U20904 (N_20904,N_19490,N_20106);
nand U20905 (N_20905,N_19245,N_19646);
and U20906 (N_20906,N_20084,N_19737);
xor U20907 (N_20907,N_19920,N_19983);
or U20908 (N_20908,N_20083,N_19557);
or U20909 (N_20909,N_19559,N_20373);
nand U20910 (N_20910,N_19549,N_20276);
or U20911 (N_20911,N_19923,N_19886);
nor U20912 (N_20912,N_19252,N_20379);
nor U20913 (N_20913,N_19499,N_20151);
xor U20914 (N_20914,N_19772,N_19248);
and U20915 (N_20915,N_20068,N_19679);
xor U20916 (N_20916,N_20385,N_19865);
xor U20917 (N_20917,N_20187,N_20283);
xor U20918 (N_20918,N_19244,N_19217);
xnor U20919 (N_20919,N_20396,N_20297);
nand U20920 (N_20920,N_19547,N_20207);
nor U20921 (N_20921,N_20023,N_19907);
or U20922 (N_20922,N_20111,N_20157);
xor U20923 (N_20923,N_19286,N_19892);
or U20924 (N_20924,N_19645,N_20172);
and U20925 (N_20925,N_20313,N_19550);
nor U20926 (N_20926,N_20075,N_19677);
xor U20927 (N_20927,N_19285,N_20226);
or U20928 (N_20928,N_20190,N_20214);
and U20929 (N_20929,N_19373,N_19227);
nand U20930 (N_20930,N_19357,N_20147);
nand U20931 (N_20931,N_19545,N_20209);
nor U20932 (N_20932,N_20182,N_19743);
nand U20933 (N_20933,N_19764,N_19532);
nor U20934 (N_20934,N_19932,N_20269);
nand U20935 (N_20935,N_19763,N_20020);
xor U20936 (N_20936,N_19694,N_20197);
xor U20937 (N_20937,N_19808,N_19895);
or U20938 (N_20938,N_20233,N_19799);
nand U20939 (N_20939,N_19873,N_19953);
or U20940 (N_20940,N_19773,N_20331);
nand U20941 (N_20941,N_20032,N_19843);
and U20942 (N_20942,N_19586,N_20165);
and U20943 (N_20943,N_19890,N_19685);
or U20944 (N_20944,N_19360,N_19819);
and U20945 (N_20945,N_19274,N_19521);
xnor U20946 (N_20946,N_20170,N_19735);
nor U20947 (N_20947,N_20273,N_19564);
nor U20948 (N_20948,N_20290,N_19207);
nand U20949 (N_20949,N_19889,N_19323);
or U20950 (N_20950,N_20119,N_19883);
and U20951 (N_20951,N_19682,N_19720);
or U20952 (N_20952,N_19788,N_19868);
xor U20953 (N_20953,N_19415,N_19544);
xor U20954 (N_20954,N_19591,N_19423);
nand U20955 (N_20955,N_19561,N_19921);
and U20956 (N_20956,N_19431,N_19365);
nor U20957 (N_20957,N_19842,N_19546);
xor U20958 (N_20958,N_19417,N_20065);
xnor U20959 (N_20959,N_19200,N_19812);
or U20960 (N_20960,N_19854,N_19965);
xnor U20961 (N_20961,N_19692,N_19657);
nand U20962 (N_20962,N_19834,N_19449);
nor U20963 (N_20963,N_19942,N_19220);
xnor U20964 (N_20964,N_19273,N_20292);
or U20965 (N_20965,N_20043,N_20105);
nor U20966 (N_20966,N_19382,N_20161);
nor U20967 (N_20967,N_19898,N_19827);
or U20968 (N_20968,N_20039,N_19987);
or U20969 (N_20969,N_20091,N_19649);
and U20970 (N_20970,N_19312,N_20057);
or U20971 (N_20971,N_20135,N_19268);
or U20972 (N_20972,N_20006,N_20186);
or U20973 (N_20973,N_19964,N_19880);
nor U20974 (N_20974,N_20295,N_19825);
nor U20975 (N_20975,N_19650,N_20311);
or U20976 (N_20976,N_20397,N_19661);
nand U20977 (N_20977,N_20024,N_19750);
nand U20978 (N_20978,N_19693,N_19802);
and U20979 (N_20979,N_19437,N_19522);
nand U20980 (N_20980,N_19560,N_20291);
nor U20981 (N_20981,N_20094,N_20007);
nor U20982 (N_20982,N_19404,N_19837);
or U20983 (N_20983,N_19826,N_19414);
nor U20984 (N_20984,N_20179,N_19698);
nand U20985 (N_20985,N_19614,N_19338);
nor U20986 (N_20986,N_19900,N_20349);
nand U20987 (N_20987,N_19619,N_19629);
xor U20988 (N_20988,N_19541,N_20252);
and U20989 (N_20989,N_19233,N_19952);
xor U20990 (N_20990,N_19659,N_20104);
xor U20991 (N_20991,N_19267,N_19632);
nor U20992 (N_20992,N_19934,N_20210);
nand U20993 (N_20993,N_19794,N_20148);
nand U20994 (N_20994,N_19931,N_19674);
xnor U20995 (N_20995,N_19955,N_19958);
nand U20996 (N_20996,N_20049,N_20171);
nand U20997 (N_20997,N_19911,N_20284);
or U20998 (N_20998,N_19454,N_19993);
xor U20999 (N_20999,N_19519,N_19986);
nor U21000 (N_21000,N_19281,N_20239);
nor U21001 (N_21001,N_19263,N_19446);
nor U21002 (N_21002,N_20362,N_19297);
nand U21003 (N_21003,N_19397,N_20038);
nor U21004 (N_21004,N_19995,N_20194);
xnor U21005 (N_21005,N_19243,N_19549);
and U21006 (N_21006,N_19696,N_20392);
and U21007 (N_21007,N_19791,N_19477);
and U21008 (N_21008,N_20000,N_19901);
xor U21009 (N_21009,N_19894,N_20017);
nand U21010 (N_21010,N_19650,N_20116);
or U21011 (N_21011,N_19748,N_19408);
or U21012 (N_21012,N_20013,N_20047);
xor U21013 (N_21013,N_20340,N_20329);
xnor U21014 (N_21014,N_20291,N_19574);
and U21015 (N_21015,N_19824,N_19249);
nor U21016 (N_21016,N_20176,N_19475);
and U21017 (N_21017,N_20087,N_20287);
and U21018 (N_21018,N_19453,N_19236);
nor U21019 (N_21019,N_19778,N_19983);
or U21020 (N_21020,N_19334,N_19771);
and U21021 (N_21021,N_19942,N_19852);
xnor U21022 (N_21022,N_19435,N_19905);
xor U21023 (N_21023,N_19594,N_20296);
or U21024 (N_21024,N_20223,N_19961);
xor U21025 (N_21025,N_19243,N_20056);
or U21026 (N_21026,N_20321,N_19919);
nor U21027 (N_21027,N_20295,N_19375);
xor U21028 (N_21028,N_19967,N_20105);
or U21029 (N_21029,N_19446,N_19929);
nand U21030 (N_21030,N_20185,N_19225);
nand U21031 (N_21031,N_20099,N_19618);
and U21032 (N_21032,N_19464,N_20351);
xor U21033 (N_21033,N_19831,N_19979);
nand U21034 (N_21034,N_20020,N_19702);
or U21035 (N_21035,N_19580,N_19234);
nand U21036 (N_21036,N_19689,N_20063);
nand U21037 (N_21037,N_19614,N_19909);
and U21038 (N_21038,N_20227,N_19983);
and U21039 (N_21039,N_20177,N_19821);
nor U21040 (N_21040,N_20208,N_20271);
and U21041 (N_21041,N_20387,N_19596);
nand U21042 (N_21042,N_19604,N_19319);
nand U21043 (N_21043,N_19281,N_19944);
or U21044 (N_21044,N_19671,N_19677);
xnor U21045 (N_21045,N_19611,N_19809);
or U21046 (N_21046,N_19437,N_20044);
nor U21047 (N_21047,N_19516,N_19380);
nand U21048 (N_21048,N_20213,N_19645);
or U21049 (N_21049,N_19566,N_19879);
and U21050 (N_21050,N_19216,N_19730);
nand U21051 (N_21051,N_20347,N_19710);
xor U21052 (N_21052,N_19687,N_19845);
nor U21053 (N_21053,N_19214,N_19833);
nand U21054 (N_21054,N_19286,N_20362);
or U21055 (N_21055,N_19362,N_20107);
and U21056 (N_21056,N_19906,N_20108);
or U21057 (N_21057,N_19270,N_19969);
and U21058 (N_21058,N_20324,N_19979);
nand U21059 (N_21059,N_19520,N_20031);
xnor U21060 (N_21060,N_20081,N_20105);
or U21061 (N_21061,N_20043,N_19957);
nor U21062 (N_21062,N_19247,N_19433);
or U21063 (N_21063,N_19698,N_19785);
and U21064 (N_21064,N_20021,N_19893);
xnor U21065 (N_21065,N_19934,N_20294);
nand U21066 (N_21066,N_20271,N_19975);
or U21067 (N_21067,N_19346,N_19771);
nand U21068 (N_21068,N_19644,N_20204);
and U21069 (N_21069,N_19918,N_19886);
xnor U21070 (N_21070,N_19996,N_20137);
or U21071 (N_21071,N_19647,N_19999);
xnor U21072 (N_21072,N_19836,N_20184);
nand U21073 (N_21073,N_19710,N_19339);
nand U21074 (N_21074,N_19765,N_19310);
nor U21075 (N_21075,N_19889,N_19920);
or U21076 (N_21076,N_19224,N_19998);
nor U21077 (N_21077,N_20208,N_19800);
and U21078 (N_21078,N_20383,N_19567);
xnor U21079 (N_21079,N_19694,N_20083);
xnor U21080 (N_21080,N_20074,N_20325);
and U21081 (N_21081,N_20112,N_19625);
nand U21082 (N_21082,N_19495,N_19390);
xnor U21083 (N_21083,N_19838,N_19986);
xnor U21084 (N_21084,N_19384,N_20205);
nand U21085 (N_21085,N_20232,N_19522);
xnor U21086 (N_21086,N_19607,N_20140);
xnor U21087 (N_21087,N_20150,N_20163);
nand U21088 (N_21088,N_19513,N_19789);
nor U21089 (N_21089,N_19987,N_20197);
nor U21090 (N_21090,N_20218,N_19821);
nor U21091 (N_21091,N_20088,N_19651);
nor U21092 (N_21092,N_19995,N_20216);
and U21093 (N_21093,N_20380,N_20204);
xnor U21094 (N_21094,N_19288,N_20337);
nand U21095 (N_21095,N_19485,N_19838);
nor U21096 (N_21096,N_19665,N_19453);
nor U21097 (N_21097,N_19318,N_19368);
xor U21098 (N_21098,N_20141,N_19905);
nor U21099 (N_21099,N_19917,N_19581);
or U21100 (N_21100,N_19783,N_20090);
and U21101 (N_21101,N_20158,N_19607);
nor U21102 (N_21102,N_19971,N_20128);
nor U21103 (N_21103,N_20111,N_20044);
xor U21104 (N_21104,N_19417,N_20376);
and U21105 (N_21105,N_19250,N_20108);
xor U21106 (N_21106,N_19499,N_19560);
xor U21107 (N_21107,N_20035,N_19307);
and U21108 (N_21108,N_20181,N_20049);
xnor U21109 (N_21109,N_19735,N_20142);
nand U21110 (N_21110,N_19877,N_19619);
or U21111 (N_21111,N_19366,N_19265);
or U21112 (N_21112,N_19588,N_20237);
nand U21113 (N_21113,N_20263,N_19778);
nor U21114 (N_21114,N_19238,N_19662);
nand U21115 (N_21115,N_20067,N_19517);
or U21116 (N_21116,N_19945,N_20275);
and U21117 (N_21117,N_19794,N_19901);
or U21118 (N_21118,N_19620,N_19822);
or U21119 (N_21119,N_20110,N_20162);
xor U21120 (N_21120,N_20335,N_19863);
and U21121 (N_21121,N_19883,N_19760);
or U21122 (N_21122,N_19608,N_20373);
nor U21123 (N_21123,N_19396,N_19380);
or U21124 (N_21124,N_20036,N_19670);
nand U21125 (N_21125,N_19490,N_20170);
and U21126 (N_21126,N_19643,N_19246);
nor U21127 (N_21127,N_20173,N_19296);
and U21128 (N_21128,N_20313,N_19880);
xnor U21129 (N_21129,N_19296,N_20227);
and U21130 (N_21130,N_19838,N_19321);
nand U21131 (N_21131,N_19398,N_19941);
xor U21132 (N_21132,N_20165,N_19653);
nand U21133 (N_21133,N_20179,N_19248);
nand U21134 (N_21134,N_20005,N_19671);
nand U21135 (N_21135,N_19627,N_20268);
xnor U21136 (N_21136,N_19810,N_19459);
nand U21137 (N_21137,N_20145,N_19693);
nor U21138 (N_21138,N_19506,N_19342);
nand U21139 (N_21139,N_19506,N_20131);
nand U21140 (N_21140,N_20060,N_20144);
and U21141 (N_21141,N_20255,N_19783);
and U21142 (N_21142,N_19284,N_20104);
and U21143 (N_21143,N_19220,N_19256);
xor U21144 (N_21144,N_20388,N_19205);
xor U21145 (N_21145,N_19784,N_19689);
xnor U21146 (N_21146,N_20195,N_20388);
or U21147 (N_21147,N_19419,N_19257);
and U21148 (N_21148,N_20088,N_20377);
nand U21149 (N_21149,N_19667,N_19528);
nor U21150 (N_21150,N_19412,N_19516);
and U21151 (N_21151,N_20251,N_20082);
nand U21152 (N_21152,N_19593,N_20066);
nand U21153 (N_21153,N_20255,N_19354);
nor U21154 (N_21154,N_19619,N_20082);
xor U21155 (N_21155,N_20134,N_19703);
xor U21156 (N_21156,N_20289,N_19678);
and U21157 (N_21157,N_20319,N_20253);
nand U21158 (N_21158,N_19636,N_19979);
or U21159 (N_21159,N_19289,N_19834);
or U21160 (N_21160,N_19267,N_19516);
nand U21161 (N_21161,N_20127,N_19449);
xor U21162 (N_21162,N_19883,N_19250);
xnor U21163 (N_21163,N_19559,N_19400);
xor U21164 (N_21164,N_20170,N_19770);
xor U21165 (N_21165,N_19513,N_19339);
xor U21166 (N_21166,N_20105,N_19856);
or U21167 (N_21167,N_19343,N_20230);
or U21168 (N_21168,N_19584,N_19448);
nand U21169 (N_21169,N_20300,N_19661);
or U21170 (N_21170,N_19977,N_19633);
and U21171 (N_21171,N_19805,N_19746);
or U21172 (N_21172,N_19632,N_19254);
and U21173 (N_21173,N_20281,N_19699);
nand U21174 (N_21174,N_20065,N_20022);
nand U21175 (N_21175,N_19379,N_19617);
xor U21176 (N_21176,N_19724,N_19747);
nor U21177 (N_21177,N_19898,N_20009);
nor U21178 (N_21178,N_19676,N_19683);
xor U21179 (N_21179,N_19301,N_20223);
or U21180 (N_21180,N_19206,N_19758);
xnor U21181 (N_21181,N_19471,N_20159);
and U21182 (N_21182,N_19232,N_20004);
or U21183 (N_21183,N_19378,N_20380);
and U21184 (N_21184,N_19357,N_19682);
and U21185 (N_21185,N_20091,N_19557);
nand U21186 (N_21186,N_19253,N_19782);
and U21187 (N_21187,N_19822,N_19389);
xnor U21188 (N_21188,N_20143,N_19357);
xnor U21189 (N_21189,N_20190,N_20015);
xor U21190 (N_21190,N_19697,N_19350);
and U21191 (N_21191,N_20117,N_19520);
nand U21192 (N_21192,N_19570,N_19237);
nor U21193 (N_21193,N_19985,N_19461);
nand U21194 (N_21194,N_19507,N_20185);
nor U21195 (N_21195,N_19480,N_20087);
xor U21196 (N_21196,N_19827,N_19311);
nor U21197 (N_21197,N_19326,N_19485);
and U21198 (N_21198,N_20339,N_20094);
xnor U21199 (N_21199,N_19723,N_19775);
and U21200 (N_21200,N_19983,N_19352);
xnor U21201 (N_21201,N_20124,N_19469);
or U21202 (N_21202,N_19264,N_20107);
xnor U21203 (N_21203,N_20325,N_19260);
or U21204 (N_21204,N_19427,N_19787);
nand U21205 (N_21205,N_19912,N_19567);
and U21206 (N_21206,N_19516,N_19868);
xnor U21207 (N_21207,N_19351,N_19246);
or U21208 (N_21208,N_20128,N_20213);
nor U21209 (N_21209,N_20341,N_20151);
and U21210 (N_21210,N_20094,N_19447);
nand U21211 (N_21211,N_20364,N_20202);
xnor U21212 (N_21212,N_19380,N_20109);
xnor U21213 (N_21213,N_19243,N_20252);
and U21214 (N_21214,N_19326,N_19309);
nor U21215 (N_21215,N_19710,N_19715);
xor U21216 (N_21216,N_19603,N_20160);
and U21217 (N_21217,N_20273,N_20347);
nand U21218 (N_21218,N_19236,N_20376);
and U21219 (N_21219,N_20038,N_19963);
xor U21220 (N_21220,N_19303,N_19283);
nand U21221 (N_21221,N_20007,N_20013);
nor U21222 (N_21222,N_19944,N_19733);
or U21223 (N_21223,N_20016,N_19362);
or U21224 (N_21224,N_19923,N_19450);
or U21225 (N_21225,N_19200,N_19659);
nor U21226 (N_21226,N_19200,N_19619);
nor U21227 (N_21227,N_19769,N_20123);
xor U21228 (N_21228,N_19454,N_19302);
nand U21229 (N_21229,N_19447,N_20319);
and U21230 (N_21230,N_20115,N_20344);
xnor U21231 (N_21231,N_19503,N_20010);
nor U21232 (N_21232,N_19697,N_19978);
nor U21233 (N_21233,N_19850,N_20163);
nor U21234 (N_21234,N_19587,N_19446);
nand U21235 (N_21235,N_19869,N_20086);
nand U21236 (N_21236,N_19864,N_19688);
or U21237 (N_21237,N_20330,N_19468);
or U21238 (N_21238,N_19445,N_19870);
xor U21239 (N_21239,N_20063,N_19939);
or U21240 (N_21240,N_20168,N_19302);
nor U21241 (N_21241,N_19639,N_20293);
nor U21242 (N_21242,N_19202,N_20365);
or U21243 (N_21243,N_19684,N_19457);
nor U21244 (N_21244,N_19661,N_19236);
nand U21245 (N_21245,N_20058,N_19946);
nor U21246 (N_21246,N_19542,N_19607);
and U21247 (N_21247,N_20230,N_19300);
and U21248 (N_21248,N_19802,N_19815);
or U21249 (N_21249,N_19373,N_19916);
xor U21250 (N_21250,N_20053,N_19519);
or U21251 (N_21251,N_20004,N_20363);
nor U21252 (N_21252,N_19967,N_19827);
nor U21253 (N_21253,N_19591,N_19854);
nor U21254 (N_21254,N_19971,N_19894);
nand U21255 (N_21255,N_19977,N_20108);
nor U21256 (N_21256,N_19950,N_20393);
nor U21257 (N_21257,N_19580,N_19370);
xor U21258 (N_21258,N_19382,N_19981);
xnor U21259 (N_21259,N_20269,N_19217);
nor U21260 (N_21260,N_19802,N_19877);
nand U21261 (N_21261,N_19492,N_19626);
nor U21262 (N_21262,N_20024,N_20296);
nor U21263 (N_21263,N_19627,N_20178);
or U21264 (N_21264,N_19307,N_19958);
nor U21265 (N_21265,N_20223,N_20324);
and U21266 (N_21266,N_20152,N_19929);
and U21267 (N_21267,N_19370,N_19441);
nor U21268 (N_21268,N_20230,N_19971);
nand U21269 (N_21269,N_19735,N_19723);
xnor U21270 (N_21270,N_19597,N_19531);
or U21271 (N_21271,N_19775,N_19760);
nor U21272 (N_21272,N_19224,N_19663);
nand U21273 (N_21273,N_20031,N_19669);
xor U21274 (N_21274,N_20348,N_20335);
nand U21275 (N_21275,N_19698,N_20058);
nor U21276 (N_21276,N_19403,N_20203);
nand U21277 (N_21277,N_19709,N_19544);
nand U21278 (N_21278,N_19319,N_19941);
nor U21279 (N_21279,N_19734,N_19684);
nand U21280 (N_21280,N_19714,N_20148);
or U21281 (N_21281,N_19614,N_19734);
nor U21282 (N_21282,N_19597,N_20202);
nor U21283 (N_21283,N_19957,N_19583);
or U21284 (N_21284,N_20027,N_20157);
nand U21285 (N_21285,N_19793,N_20387);
or U21286 (N_21286,N_19649,N_19374);
nor U21287 (N_21287,N_20366,N_19939);
xnor U21288 (N_21288,N_19525,N_19733);
nand U21289 (N_21289,N_19427,N_19445);
nor U21290 (N_21290,N_19610,N_20150);
and U21291 (N_21291,N_19225,N_20387);
nand U21292 (N_21292,N_19252,N_19983);
and U21293 (N_21293,N_20164,N_19822);
nand U21294 (N_21294,N_19345,N_20230);
and U21295 (N_21295,N_20112,N_20189);
nor U21296 (N_21296,N_20011,N_20352);
or U21297 (N_21297,N_19234,N_20170);
and U21298 (N_21298,N_19520,N_19511);
nand U21299 (N_21299,N_19552,N_20266);
nand U21300 (N_21300,N_19537,N_20075);
nand U21301 (N_21301,N_19419,N_19219);
xnor U21302 (N_21302,N_19948,N_19835);
and U21303 (N_21303,N_19847,N_19943);
or U21304 (N_21304,N_20104,N_20179);
nor U21305 (N_21305,N_19567,N_19502);
nand U21306 (N_21306,N_19532,N_20030);
nand U21307 (N_21307,N_19423,N_20268);
nand U21308 (N_21308,N_19939,N_20282);
nand U21309 (N_21309,N_19498,N_19975);
or U21310 (N_21310,N_19684,N_20022);
and U21311 (N_21311,N_19221,N_19770);
nand U21312 (N_21312,N_19654,N_19274);
or U21313 (N_21313,N_20236,N_19951);
and U21314 (N_21314,N_19403,N_20274);
nor U21315 (N_21315,N_20372,N_19527);
or U21316 (N_21316,N_19544,N_19854);
and U21317 (N_21317,N_19789,N_19214);
xor U21318 (N_21318,N_20254,N_19219);
and U21319 (N_21319,N_20261,N_20164);
nand U21320 (N_21320,N_19320,N_19602);
nor U21321 (N_21321,N_19969,N_19399);
xnor U21322 (N_21322,N_20386,N_19578);
and U21323 (N_21323,N_19892,N_20136);
nor U21324 (N_21324,N_20263,N_20190);
or U21325 (N_21325,N_20291,N_19895);
nand U21326 (N_21326,N_19684,N_19377);
xor U21327 (N_21327,N_20075,N_19248);
nor U21328 (N_21328,N_19818,N_19685);
xor U21329 (N_21329,N_19529,N_19933);
or U21330 (N_21330,N_20099,N_19234);
and U21331 (N_21331,N_19731,N_19924);
nor U21332 (N_21332,N_19334,N_19361);
nand U21333 (N_21333,N_20223,N_19300);
nand U21334 (N_21334,N_19367,N_19799);
nor U21335 (N_21335,N_20219,N_20161);
nor U21336 (N_21336,N_19308,N_20097);
nand U21337 (N_21337,N_19504,N_19923);
nor U21338 (N_21338,N_20253,N_19310);
nand U21339 (N_21339,N_19732,N_19522);
nand U21340 (N_21340,N_20133,N_19489);
or U21341 (N_21341,N_20094,N_19318);
nor U21342 (N_21342,N_19967,N_19450);
xnor U21343 (N_21343,N_19444,N_20378);
and U21344 (N_21344,N_20118,N_20397);
or U21345 (N_21345,N_19483,N_20193);
nand U21346 (N_21346,N_19290,N_19980);
xnor U21347 (N_21347,N_19601,N_19972);
and U21348 (N_21348,N_19747,N_20019);
and U21349 (N_21349,N_19691,N_19296);
and U21350 (N_21350,N_20241,N_20000);
nor U21351 (N_21351,N_20352,N_19725);
nor U21352 (N_21352,N_19500,N_19729);
nand U21353 (N_21353,N_19505,N_19376);
and U21354 (N_21354,N_20008,N_19588);
nand U21355 (N_21355,N_19338,N_20334);
and U21356 (N_21356,N_19371,N_20014);
nand U21357 (N_21357,N_19242,N_19458);
and U21358 (N_21358,N_19821,N_20075);
and U21359 (N_21359,N_19843,N_20111);
and U21360 (N_21360,N_19768,N_19836);
nand U21361 (N_21361,N_20007,N_20099);
or U21362 (N_21362,N_19613,N_19518);
nand U21363 (N_21363,N_19567,N_19501);
nand U21364 (N_21364,N_19838,N_19845);
nand U21365 (N_21365,N_20271,N_19295);
and U21366 (N_21366,N_19215,N_20320);
and U21367 (N_21367,N_19252,N_19626);
or U21368 (N_21368,N_19853,N_19999);
and U21369 (N_21369,N_20254,N_20238);
or U21370 (N_21370,N_19692,N_20022);
nand U21371 (N_21371,N_20182,N_20160);
nor U21372 (N_21372,N_20067,N_20137);
nand U21373 (N_21373,N_19754,N_19314);
xnor U21374 (N_21374,N_20399,N_20145);
and U21375 (N_21375,N_19364,N_20032);
and U21376 (N_21376,N_19350,N_19801);
nor U21377 (N_21377,N_19501,N_19638);
and U21378 (N_21378,N_19684,N_20201);
nand U21379 (N_21379,N_19697,N_20195);
and U21380 (N_21380,N_20061,N_20144);
or U21381 (N_21381,N_20165,N_19583);
or U21382 (N_21382,N_20230,N_20362);
xnor U21383 (N_21383,N_19510,N_19428);
nor U21384 (N_21384,N_19706,N_20232);
xor U21385 (N_21385,N_19515,N_20224);
nor U21386 (N_21386,N_19960,N_19474);
nor U21387 (N_21387,N_19454,N_19459);
and U21388 (N_21388,N_20089,N_20184);
and U21389 (N_21389,N_19506,N_19914);
nor U21390 (N_21390,N_19996,N_19358);
nor U21391 (N_21391,N_20054,N_20291);
or U21392 (N_21392,N_20080,N_20204);
nor U21393 (N_21393,N_19364,N_19603);
or U21394 (N_21394,N_19913,N_19206);
nor U21395 (N_21395,N_19723,N_19504);
and U21396 (N_21396,N_20224,N_19773);
and U21397 (N_21397,N_19485,N_19236);
nand U21398 (N_21398,N_19996,N_19804);
or U21399 (N_21399,N_20194,N_19684);
or U21400 (N_21400,N_20272,N_19552);
nor U21401 (N_21401,N_20179,N_19326);
nor U21402 (N_21402,N_19319,N_19638);
and U21403 (N_21403,N_19792,N_20346);
and U21404 (N_21404,N_20167,N_20173);
xnor U21405 (N_21405,N_19617,N_19354);
and U21406 (N_21406,N_20075,N_20270);
nor U21407 (N_21407,N_20280,N_20191);
nand U21408 (N_21408,N_19520,N_19377);
nor U21409 (N_21409,N_20070,N_19430);
or U21410 (N_21410,N_19644,N_19767);
xnor U21411 (N_21411,N_20123,N_19748);
nand U21412 (N_21412,N_19513,N_19738);
or U21413 (N_21413,N_19627,N_19974);
nor U21414 (N_21414,N_20065,N_19562);
nand U21415 (N_21415,N_19835,N_19403);
xor U21416 (N_21416,N_20109,N_19660);
or U21417 (N_21417,N_19236,N_19712);
nand U21418 (N_21418,N_19804,N_19911);
xor U21419 (N_21419,N_19835,N_20109);
xor U21420 (N_21420,N_19550,N_19930);
nor U21421 (N_21421,N_19710,N_20094);
nor U21422 (N_21422,N_19536,N_19585);
nor U21423 (N_21423,N_19436,N_20226);
or U21424 (N_21424,N_19274,N_19850);
xnor U21425 (N_21425,N_19902,N_19584);
and U21426 (N_21426,N_19975,N_19918);
xnor U21427 (N_21427,N_20246,N_19626);
nor U21428 (N_21428,N_20195,N_19515);
nor U21429 (N_21429,N_19226,N_20296);
xor U21430 (N_21430,N_19722,N_19887);
nand U21431 (N_21431,N_19958,N_19308);
xor U21432 (N_21432,N_20092,N_20334);
or U21433 (N_21433,N_20185,N_20360);
nand U21434 (N_21434,N_19409,N_19341);
or U21435 (N_21435,N_19316,N_20053);
nand U21436 (N_21436,N_19661,N_20264);
or U21437 (N_21437,N_19647,N_19576);
and U21438 (N_21438,N_20195,N_20001);
or U21439 (N_21439,N_19259,N_19766);
nand U21440 (N_21440,N_19778,N_20225);
nand U21441 (N_21441,N_19313,N_20308);
nor U21442 (N_21442,N_19559,N_20229);
xnor U21443 (N_21443,N_19369,N_19266);
nor U21444 (N_21444,N_20152,N_20086);
or U21445 (N_21445,N_20044,N_19692);
nand U21446 (N_21446,N_19478,N_19925);
nand U21447 (N_21447,N_19363,N_19572);
nor U21448 (N_21448,N_19813,N_20388);
or U21449 (N_21449,N_19371,N_19258);
and U21450 (N_21450,N_19734,N_20317);
nand U21451 (N_21451,N_19950,N_20391);
and U21452 (N_21452,N_19367,N_19240);
nor U21453 (N_21453,N_19257,N_20296);
xor U21454 (N_21454,N_20137,N_19672);
and U21455 (N_21455,N_19649,N_19335);
or U21456 (N_21456,N_19355,N_20388);
xnor U21457 (N_21457,N_19995,N_19716);
nand U21458 (N_21458,N_19932,N_19332);
or U21459 (N_21459,N_19804,N_19825);
and U21460 (N_21460,N_19275,N_19477);
or U21461 (N_21461,N_19527,N_19614);
or U21462 (N_21462,N_19928,N_19584);
nor U21463 (N_21463,N_19620,N_20151);
and U21464 (N_21464,N_19804,N_19450);
xnor U21465 (N_21465,N_19284,N_20239);
nor U21466 (N_21466,N_19972,N_19331);
and U21467 (N_21467,N_19341,N_19328);
and U21468 (N_21468,N_20399,N_19654);
nor U21469 (N_21469,N_20182,N_19441);
and U21470 (N_21470,N_20116,N_19290);
nor U21471 (N_21471,N_19287,N_20198);
xnor U21472 (N_21472,N_20049,N_19957);
xnor U21473 (N_21473,N_19707,N_19956);
xnor U21474 (N_21474,N_20319,N_20356);
nand U21475 (N_21475,N_19969,N_19245);
nand U21476 (N_21476,N_20079,N_19972);
nor U21477 (N_21477,N_19407,N_19282);
or U21478 (N_21478,N_20089,N_20384);
xnor U21479 (N_21479,N_20176,N_19665);
and U21480 (N_21480,N_19537,N_19581);
nand U21481 (N_21481,N_19484,N_20220);
xor U21482 (N_21482,N_19509,N_20312);
and U21483 (N_21483,N_20249,N_19693);
and U21484 (N_21484,N_19854,N_19667);
nor U21485 (N_21485,N_19255,N_19337);
xor U21486 (N_21486,N_20091,N_19592);
and U21487 (N_21487,N_19797,N_19475);
nor U21488 (N_21488,N_20005,N_20057);
xor U21489 (N_21489,N_19249,N_19208);
and U21490 (N_21490,N_20004,N_19747);
and U21491 (N_21491,N_19711,N_19529);
nor U21492 (N_21492,N_20363,N_19351);
or U21493 (N_21493,N_19783,N_19547);
xnor U21494 (N_21494,N_19490,N_19814);
xnor U21495 (N_21495,N_20376,N_20281);
and U21496 (N_21496,N_20218,N_20322);
and U21497 (N_21497,N_19374,N_20066);
xor U21498 (N_21498,N_19847,N_20084);
nand U21499 (N_21499,N_20007,N_19987);
nor U21500 (N_21500,N_19389,N_19636);
and U21501 (N_21501,N_20093,N_19683);
and U21502 (N_21502,N_20244,N_19397);
or U21503 (N_21503,N_19750,N_20371);
or U21504 (N_21504,N_19297,N_20005);
xnor U21505 (N_21505,N_19835,N_19794);
nor U21506 (N_21506,N_19791,N_19267);
nand U21507 (N_21507,N_19650,N_19844);
nor U21508 (N_21508,N_20302,N_19968);
or U21509 (N_21509,N_19836,N_19358);
or U21510 (N_21510,N_19888,N_19486);
or U21511 (N_21511,N_19875,N_20190);
nor U21512 (N_21512,N_19488,N_20100);
xnor U21513 (N_21513,N_19231,N_19956);
and U21514 (N_21514,N_20254,N_19698);
nor U21515 (N_21515,N_20141,N_19793);
and U21516 (N_21516,N_20058,N_19209);
or U21517 (N_21517,N_20243,N_19704);
nor U21518 (N_21518,N_19406,N_20099);
xnor U21519 (N_21519,N_20300,N_19327);
xor U21520 (N_21520,N_19688,N_19647);
nand U21521 (N_21521,N_19739,N_19774);
xnor U21522 (N_21522,N_19678,N_19748);
nor U21523 (N_21523,N_19963,N_19292);
nand U21524 (N_21524,N_19687,N_19756);
or U21525 (N_21525,N_19901,N_19881);
and U21526 (N_21526,N_19882,N_20231);
or U21527 (N_21527,N_19629,N_19833);
nand U21528 (N_21528,N_19871,N_19578);
and U21529 (N_21529,N_20120,N_20330);
xnor U21530 (N_21530,N_20183,N_19772);
xnor U21531 (N_21531,N_19853,N_19721);
and U21532 (N_21532,N_19471,N_19660);
nand U21533 (N_21533,N_20166,N_19704);
nor U21534 (N_21534,N_19282,N_19517);
xnor U21535 (N_21535,N_19398,N_19911);
or U21536 (N_21536,N_20220,N_19803);
and U21537 (N_21537,N_19596,N_19584);
xnor U21538 (N_21538,N_19865,N_19499);
nor U21539 (N_21539,N_20326,N_19953);
nor U21540 (N_21540,N_19286,N_19983);
nor U21541 (N_21541,N_20122,N_19867);
and U21542 (N_21542,N_19425,N_19225);
nand U21543 (N_21543,N_20318,N_19719);
xor U21544 (N_21544,N_19863,N_19218);
nand U21545 (N_21545,N_19524,N_19461);
nand U21546 (N_21546,N_19677,N_19808);
nor U21547 (N_21547,N_19249,N_19510);
or U21548 (N_21548,N_19451,N_19742);
nand U21549 (N_21549,N_19442,N_19219);
and U21550 (N_21550,N_19987,N_20362);
or U21551 (N_21551,N_19831,N_19332);
nand U21552 (N_21552,N_19910,N_20229);
xnor U21553 (N_21553,N_19510,N_19745);
nand U21554 (N_21554,N_19320,N_19697);
nor U21555 (N_21555,N_19807,N_19784);
and U21556 (N_21556,N_20257,N_20033);
and U21557 (N_21557,N_20299,N_19637);
xor U21558 (N_21558,N_19491,N_20195);
nor U21559 (N_21559,N_19362,N_20209);
nor U21560 (N_21560,N_19973,N_19888);
nor U21561 (N_21561,N_20304,N_19331);
nand U21562 (N_21562,N_19268,N_19750);
nor U21563 (N_21563,N_19216,N_19742);
xor U21564 (N_21564,N_19901,N_19891);
xor U21565 (N_21565,N_20187,N_19344);
nor U21566 (N_21566,N_19648,N_19875);
nor U21567 (N_21567,N_19347,N_20374);
or U21568 (N_21568,N_20276,N_19618);
and U21569 (N_21569,N_19204,N_20263);
or U21570 (N_21570,N_20064,N_20009);
xnor U21571 (N_21571,N_19489,N_19765);
xor U21572 (N_21572,N_19849,N_19378);
or U21573 (N_21573,N_20276,N_20030);
nor U21574 (N_21574,N_19306,N_19660);
nor U21575 (N_21575,N_19712,N_20164);
nand U21576 (N_21576,N_19290,N_19316);
xor U21577 (N_21577,N_20043,N_19794);
or U21578 (N_21578,N_19490,N_20064);
and U21579 (N_21579,N_20069,N_19449);
nor U21580 (N_21580,N_20036,N_19904);
nor U21581 (N_21581,N_20241,N_19631);
nand U21582 (N_21582,N_19526,N_19765);
and U21583 (N_21583,N_20259,N_20157);
nand U21584 (N_21584,N_20292,N_20111);
and U21585 (N_21585,N_19961,N_20315);
nand U21586 (N_21586,N_19408,N_19241);
xnor U21587 (N_21587,N_20166,N_19347);
nand U21588 (N_21588,N_19441,N_19202);
and U21589 (N_21589,N_19986,N_20392);
or U21590 (N_21590,N_20205,N_20095);
nor U21591 (N_21591,N_19357,N_20292);
and U21592 (N_21592,N_19642,N_19576);
nand U21593 (N_21593,N_19426,N_20174);
xnor U21594 (N_21594,N_20310,N_19521);
nor U21595 (N_21595,N_20136,N_19742);
and U21596 (N_21596,N_19931,N_20120);
and U21597 (N_21597,N_20357,N_19601);
and U21598 (N_21598,N_19834,N_19415);
nor U21599 (N_21599,N_19581,N_19490);
and U21600 (N_21600,N_20436,N_21561);
nor U21601 (N_21601,N_20488,N_20551);
xnor U21602 (N_21602,N_20697,N_21302);
nand U21603 (N_21603,N_21495,N_21291);
xnor U21604 (N_21604,N_20520,N_21278);
nor U21605 (N_21605,N_20595,N_20861);
xor U21606 (N_21606,N_21140,N_20995);
or U21607 (N_21607,N_21457,N_21388);
nand U21608 (N_21608,N_21306,N_21204);
or U21609 (N_21609,N_21368,N_20678);
and U21610 (N_21610,N_20826,N_20792);
nor U21611 (N_21611,N_20926,N_21118);
and U21612 (N_21612,N_20968,N_21122);
xor U21613 (N_21613,N_21314,N_21079);
nand U21614 (N_21614,N_21395,N_20870);
nor U21615 (N_21615,N_21459,N_21530);
nand U21616 (N_21616,N_21003,N_21198);
nor U21617 (N_21617,N_21045,N_20925);
and U21618 (N_21618,N_20529,N_20539);
and U21619 (N_21619,N_21563,N_21564);
or U21620 (N_21620,N_20450,N_21181);
nor U21621 (N_21621,N_21013,N_20898);
or U21622 (N_21622,N_20648,N_21018);
nor U21623 (N_21623,N_20901,N_21266);
or U21624 (N_21624,N_20430,N_20515);
nor U21625 (N_21625,N_20560,N_20542);
xor U21626 (N_21626,N_20512,N_20670);
xnor U21627 (N_21627,N_21133,N_21321);
and U21628 (N_21628,N_20504,N_20969);
or U21629 (N_21629,N_21475,N_21543);
nand U21630 (N_21630,N_20781,N_21059);
nand U21631 (N_21631,N_20526,N_20786);
nor U21632 (N_21632,N_21505,N_21086);
nor U21633 (N_21633,N_20958,N_20837);
xor U21634 (N_21634,N_20650,N_21139);
nor U21635 (N_21635,N_21248,N_21216);
nor U21636 (N_21636,N_21332,N_21579);
nor U21637 (N_21637,N_20710,N_20664);
xor U21638 (N_21638,N_21326,N_20846);
and U21639 (N_21639,N_21386,N_20772);
xnor U21640 (N_21640,N_21218,N_20506);
or U21641 (N_21641,N_21017,N_20745);
or U21642 (N_21642,N_21214,N_21051);
nand U21643 (N_21643,N_20936,N_21322);
nand U21644 (N_21644,N_21485,N_20696);
and U21645 (N_21645,N_20619,N_20530);
nor U21646 (N_21646,N_21043,N_20695);
nor U21647 (N_21647,N_20991,N_21477);
nor U21648 (N_21648,N_20419,N_20495);
xnor U21649 (N_21649,N_20460,N_21022);
or U21650 (N_21650,N_21330,N_20623);
xor U21651 (N_21651,N_21424,N_20747);
and U21652 (N_21652,N_20730,N_20802);
and U21653 (N_21653,N_21279,N_21262);
nand U21654 (N_21654,N_20957,N_21597);
and U21655 (N_21655,N_20765,N_20501);
nand U21656 (N_21656,N_21200,N_21098);
nand U21657 (N_21657,N_20513,N_21483);
and U21658 (N_21658,N_20559,N_21168);
xnor U21659 (N_21659,N_21491,N_20514);
nand U21660 (N_21660,N_21587,N_21565);
and U21661 (N_21661,N_21039,N_21105);
and U21662 (N_21662,N_21557,N_21578);
xnor U21663 (N_21663,N_20585,N_20437);
nand U21664 (N_21664,N_20653,N_21504);
nand U21665 (N_21665,N_20531,N_21351);
xor U21666 (N_21666,N_20828,N_20647);
nand U21667 (N_21667,N_21244,N_20796);
or U21668 (N_21668,N_21325,N_20609);
nor U21669 (N_21669,N_20541,N_20694);
and U21670 (N_21670,N_20836,N_21206);
or U21671 (N_21671,N_21531,N_21427);
xnor U21672 (N_21672,N_20987,N_21331);
or U21673 (N_21673,N_21113,N_21099);
xnor U21674 (N_21674,N_20610,N_20919);
and U21675 (N_21675,N_20645,N_21102);
xor U21676 (N_21676,N_21342,N_21169);
nand U21677 (N_21677,N_20461,N_21519);
or U21678 (N_21678,N_21375,N_21577);
or U21679 (N_21679,N_20438,N_20472);
nand U21680 (N_21680,N_20762,N_21154);
nor U21681 (N_21681,N_21152,N_20895);
or U21682 (N_21682,N_20462,N_21467);
and U21683 (N_21683,N_20689,N_21445);
and U21684 (N_21684,N_21145,N_21123);
nand U21685 (N_21685,N_20743,N_21219);
or U21686 (N_21686,N_20660,N_21560);
and U21687 (N_21687,N_21398,N_20739);
nor U21688 (N_21688,N_20459,N_20847);
xor U21689 (N_21689,N_21469,N_21106);
or U21690 (N_21690,N_20833,N_20582);
and U21691 (N_21691,N_20661,N_20722);
xor U21692 (N_21692,N_21307,N_21525);
or U21693 (N_21693,N_20517,N_20476);
or U21694 (N_21694,N_20561,N_21005);
nor U21695 (N_21695,N_20606,N_21015);
nand U21696 (N_21696,N_21054,N_21409);
nand U21697 (N_21697,N_21383,N_21456);
nand U21698 (N_21698,N_20983,N_21189);
nor U21699 (N_21699,N_20852,N_21134);
and U21700 (N_21700,N_20814,N_21496);
and U21701 (N_21701,N_20916,N_20713);
and U21702 (N_21702,N_21261,N_20753);
xnor U21703 (N_21703,N_20912,N_20931);
and U21704 (N_21704,N_20558,N_20600);
xor U21705 (N_21705,N_21430,N_20475);
xor U21706 (N_21706,N_21372,N_21008);
and U21707 (N_21707,N_20598,N_20769);
nand U21708 (N_21708,N_21156,N_20776);
nor U21709 (N_21709,N_20599,N_21444);
and U21710 (N_21710,N_21173,N_21364);
and U21711 (N_21711,N_21570,N_20808);
or U21712 (N_21712,N_20857,N_20646);
or U21713 (N_21713,N_21545,N_21104);
nor U21714 (N_21714,N_20627,N_21425);
xor U21715 (N_21715,N_20589,N_21362);
or U21716 (N_21716,N_20620,N_21247);
nand U21717 (N_21717,N_21510,N_20679);
xnor U21718 (N_21718,N_21144,N_21275);
nor U21719 (N_21719,N_21452,N_20939);
nor U21720 (N_21720,N_20920,N_21205);
xnor U21721 (N_21721,N_20990,N_20942);
or U21722 (N_21722,N_21340,N_21396);
nor U21723 (N_21723,N_21230,N_20644);
nor U21724 (N_21724,N_21356,N_20911);
xor U21725 (N_21725,N_21111,N_21517);
xor U21726 (N_21726,N_21448,N_21450);
xor U21727 (N_21727,N_21366,N_20510);
nand U21728 (N_21728,N_20789,N_20402);
xor U21729 (N_21729,N_20737,N_20825);
xor U21730 (N_21730,N_20928,N_20963);
nor U21731 (N_21731,N_20625,N_20701);
nor U21732 (N_21732,N_20929,N_20955);
and U21733 (N_21733,N_20863,N_20432);
xnor U21734 (N_21734,N_20824,N_21064);
xnor U21735 (N_21735,N_21527,N_20470);
xor U21736 (N_21736,N_20817,N_20856);
or U21737 (N_21737,N_21470,N_21514);
xnor U21738 (N_21738,N_21007,N_21049);
or U21739 (N_21739,N_21567,N_21107);
nand U21740 (N_21740,N_20552,N_20652);
xnor U21741 (N_21741,N_20700,N_21374);
nor U21742 (N_21742,N_21016,N_21373);
and U21743 (N_21743,N_21103,N_21112);
nor U21744 (N_21744,N_21135,N_20649);
nand U21745 (N_21745,N_21593,N_20575);
nand U21746 (N_21746,N_21025,N_21050);
or U21747 (N_21747,N_20499,N_21091);
nand U21748 (N_21748,N_21087,N_20704);
nor U21749 (N_21749,N_20937,N_20671);
or U21750 (N_21750,N_21419,N_21500);
or U21751 (N_21751,N_21382,N_20994);
nand U21752 (N_21752,N_20715,N_21129);
xor U21753 (N_21753,N_21063,N_21384);
nand U21754 (N_21754,N_21207,N_20758);
or U21755 (N_21755,N_21153,N_20434);
nand U21756 (N_21756,N_21175,N_21131);
xor U21757 (N_21757,N_21268,N_20793);
or U21758 (N_21758,N_21329,N_20917);
nand U21759 (N_21759,N_21060,N_21237);
or U21760 (N_21760,N_20413,N_20643);
xor U21761 (N_21761,N_21088,N_21595);
and U21762 (N_21762,N_21501,N_20570);
or U21763 (N_21763,N_21355,N_20822);
nor U21764 (N_21764,N_20734,N_21455);
and U21765 (N_21765,N_20489,N_21480);
and U21766 (N_21766,N_20746,N_21413);
nand U21767 (N_21767,N_20617,N_20707);
nand U21768 (N_21768,N_20741,N_20744);
nor U21769 (N_21769,N_21257,N_21432);
nand U21770 (N_21770,N_20611,N_21164);
nand U21771 (N_21771,N_21594,N_20634);
xor U21772 (N_21772,N_21172,N_20540);
xnor U21773 (N_21773,N_20950,N_21232);
and U21774 (N_21774,N_20618,N_20806);
and U21775 (N_21775,N_20705,N_20468);
nand U21776 (N_21776,N_21271,N_20799);
and U21777 (N_21777,N_20457,N_21532);
or U21778 (N_21778,N_20684,N_21488);
and U21779 (N_21779,N_21334,N_20573);
nor U21780 (N_21780,N_20960,N_21202);
nand U21781 (N_21781,N_21192,N_21072);
nor U21782 (N_21782,N_20401,N_20621);
or U21783 (N_21783,N_21160,N_20777);
nand U21784 (N_21784,N_21370,N_20778);
nor U21785 (N_21785,N_21223,N_21288);
or U21786 (N_21786,N_21150,N_21171);
nor U21787 (N_21787,N_21414,N_21367);
and U21788 (N_21788,N_21224,N_20435);
and U21789 (N_21789,N_21081,N_21379);
or U21790 (N_21790,N_20732,N_21085);
or U21791 (N_21791,N_21341,N_20569);
nand U21792 (N_21792,N_21141,N_21109);
xnor U21793 (N_21793,N_21253,N_20673);
or U21794 (N_21794,N_20426,N_21599);
or U21795 (N_21795,N_21494,N_21255);
or U21796 (N_21796,N_20924,N_21451);
xnor U21797 (N_21797,N_20997,N_20736);
nand U21798 (N_21798,N_21231,N_21337);
and U21799 (N_21799,N_21260,N_20632);
nor U21800 (N_21800,N_21211,N_20980);
nor U21801 (N_21801,N_21352,N_20742);
or U21802 (N_21802,N_21497,N_21296);
xor U21803 (N_21803,N_21486,N_20502);
and U21804 (N_21804,N_20760,N_21209);
nor U21805 (N_21805,N_21110,N_21363);
or U21806 (N_21806,N_20505,N_20400);
nor U21807 (N_21807,N_20784,N_20441);
xnor U21808 (N_21808,N_21250,N_21267);
nand U21809 (N_21809,N_20731,N_20654);
or U21810 (N_21810,N_21127,N_20616);
xor U21811 (N_21811,N_21286,N_21083);
xnor U21812 (N_21812,N_20768,N_20718);
nor U21813 (N_21813,N_20479,N_21507);
nand U21814 (N_21814,N_21259,N_21070);
nor U21815 (N_21815,N_20500,N_21242);
xor U21816 (N_21816,N_20840,N_20439);
or U21817 (N_21817,N_21193,N_20940);
or U21818 (N_21818,N_21299,N_21512);
nor U21819 (N_21819,N_20448,N_20951);
xnor U21820 (N_21820,N_20961,N_20424);
nor U21821 (N_21821,N_20574,N_20615);
or U21822 (N_21822,N_21024,N_21534);
and U21823 (N_21823,N_20887,N_20474);
and U21824 (N_21824,N_20491,N_21023);
xor U21825 (N_21825,N_21442,N_21208);
and U21826 (N_21826,N_20528,N_20959);
nor U21827 (N_21827,N_21499,N_21138);
or U21828 (N_21828,N_21040,N_21201);
nor U21829 (N_21829,N_20578,N_20985);
xor U21830 (N_21830,N_21069,N_20442);
or U21831 (N_21831,N_20603,N_20412);
or U21832 (N_21832,N_21041,N_21526);
xnor U21833 (N_21833,N_21392,N_21163);
and U21834 (N_21834,N_21184,N_20555);
nor U21835 (N_21835,N_20922,N_21055);
nor U21836 (N_21836,N_20761,N_20456);
nor U21837 (N_21837,N_21280,N_20706);
and U21838 (N_21838,N_21272,N_20878);
nor U21839 (N_21839,N_20804,N_20910);
nor U21840 (N_21840,N_20674,N_20563);
xnor U21841 (N_21841,N_20899,N_20659);
nand U21842 (N_21842,N_21136,N_21101);
xor U21843 (N_21843,N_21227,N_21585);
nor U21844 (N_21844,N_21137,N_20818);
nand U21845 (N_21845,N_20536,N_21581);
xnor U21846 (N_21846,N_20820,N_20841);
nor U21847 (N_21847,N_20717,N_21550);
xor U21848 (N_21848,N_21197,N_20642);
nand U21849 (N_21849,N_20680,N_21402);
nor U21850 (N_21850,N_20867,N_21580);
nand U21851 (N_21851,N_21044,N_20974);
xnor U21852 (N_21852,N_20699,N_21555);
xor U21853 (N_21853,N_21377,N_20411);
nor U21854 (N_21854,N_20809,N_20735);
nor U21855 (N_21855,N_20449,N_20755);
and U21856 (N_21856,N_20440,N_21057);
and U21857 (N_21857,N_21026,N_21598);
nor U21858 (N_21858,N_20879,N_20467);
and U21859 (N_21859,N_21312,N_20473);
and U21860 (N_21860,N_21174,N_20894);
nand U21861 (N_21861,N_20834,N_20947);
or U21862 (N_21862,N_20945,N_20794);
nor U21863 (N_21863,N_21343,N_20738);
xnor U21864 (N_21864,N_21407,N_21001);
nand U21865 (N_21865,N_21421,N_20759);
or U21866 (N_21866,N_21270,N_21317);
xnor U21867 (N_21867,N_20481,N_21084);
xnor U21868 (N_21868,N_21394,N_21339);
or U21869 (N_21869,N_20444,N_20798);
nand U21870 (N_21870,N_20909,N_21359);
nand U21871 (N_21871,N_21195,N_21465);
nor U21872 (N_21872,N_20408,N_20535);
nand U21873 (N_21873,N_20845,N_21096);
or U21874 (N_21874,N_21126,N_21498);
or U21875 (N_21875,N_20884,N_21361);
nor U21876 (N_21876,N_20830,N_20921);
nor U21877 (N_21877,N_21116,N_20729);
nor U21878 (N_21878,N_21019,N_20638);
xnor U21879 (N_21879,N_21516,N_20976);
nand U21880 (N_21880,N_20810,N_20771);
or U21881 (N_21881,N_20888,N_20483);
nand U21882 (N_21882,N_21385,N_20405);
or U21883 (N_21883,N_21588,N_20604);
xnor U21884 (N_21884,N_20409,N_21241);
xor U21885 (N_21885,N_20859,N_21165);
xnor U21886 (N_21886,N_20767,N_20494);
xor U21887 (N_21887,N_21380,N_21426);
nand U21888 (N_21888,N_21324,N_20900);
or U21889 (N_21889,N_21575,N_20832);
nor U21890 (N_21890,N_21090,N_20544);
nor U21891 (N_21891,N_21428,N_21574);
xor U21892 (N_21892,N_21011,N_21401);
or U21893 (N_21893,N_21590,N_21520);
or U21894 (N_21894,N_20865,N_20429);
nor U21895 (N_21895,N_20905,N_21474);
nor U21896 (N_21896,N_20593,N_21252);
and U21897 (N_21897,N_21052,N_20756);
or U21898 (N_21898,N_20629,N_20724);
nand U21899 (N_21899,N_21433,N_21410);
and U21900 (N_21900,N_20795,N_20787);
nor U21901 (N_21901,N_20581,N_20537);
nand U21902 (N_21902,N_20877,N_21573);
and U21903 (N_21903,N_20675,N_21082);
xor U21904 (N_21904,N_20893,N_20658);
and U21905 (N_21905,N_20605,N_20907);
or U21906 (N_21906,N_20757,N_20883);
nand U21907 (N_21907,N_20667,N_20485);
nand U21908 (N_21908,N_20404,N_20607);
or U21909 (N_21909,N_20886,N_20972);
nor U21910 (N_21910,N_20524,N_20676);
and U21911 (N_21911,N_21400,N_21157);
and U21912 (N_21912,N_20518,N_21158);
xnor U21913 (N_21913,N_20709,N_21269);
nand U21914 (N_21914,N_21535,N_20498);
xnor U21915 (N_21915,N_21404,N_21481);
and U21916 (N_21916,N_20588,N_20783);
nand U21917 (N_21917,N_20596,N_21177);
nor U21918 (N_21918,N_20406,N_20641);
or U21919 (N_21919,N_21490,N_20612);
nor U21920 (N_21920,N_20933,N_20601);
or U21921 (N_21921,N_20967,N_21586);
xnor U21922 (N_21922,N_21417,N_21552);
nor U21923 (N_21923,N_20938,N_21547);
and U21924 (N_21924,N_21142,N_20511);
and U21925 (N_21925,N_21066,N_21021);
xnor U21926 (N_21926,N_20516,N_20428);
nand U21927 (N_21927,N_20477,N_21371);
and U21928 (N_21928,N_20547,N_21249);
nand U21929 (N_21929,N_20666,N_21551);
xnor U21930 (N_21930,N_21418,N_20949);
or U21931 (N_21931,N_20527,N_21309);
xnor U21932 (N_21932,N_20848,N_20977);
and U21933 (N_21933,N_21596,N_20764);
nor U21934 (N_21934,N_20838,N_21243);
xnor U21935 (N_21935,N_20779,N_20628);
xnor U21936 (N_21936,N_21524,N_21365);
nand U21937 (N_21937,N_20443,N_20640);
or U21938 (N_21938,N_20656,N_20876);
nand U21939 (N_21939,N_21254,N_20571);
nor U21940 (N_21940,N_20948,N_20874);
or U21941 (N_21941,N_21592,N_21540);
or U21942 (N_21942,N_21196,N_21221);
xor U21943 (N_21943,N_20851,N_21391);
nand U21944 (N_21944,N_20813,N_21493);
nand U21945 (N_21945,N_20835,N_21313);
or U21946 (N_21946,N_20932,N_21478);
nor U21947 (N_21947,N_20478,N_21285);
or U21948 (N_21948,N_20631,N_21037);
nor U21949 (N_21949,N_20608,N_20885);
xnor U21950 (N_21950,N_20725,N_21360);
or U21951 (N_21951,N_20698,N_21548);
xnor U21952 (N_21952,N_21075,N_21074);
or U21953 (N_21953,N_21130,N_21303);
and U21954 (N_21954,N_21294,N_20637);
xnor U21955 (N_21955,N_20831,N_20984);
xnor U21956 (N_21956,N_20770,N_21284);
xnor U21957 (N_21957,N_20418,N_20891);
and U21958 (N_21958,N_21357,N_20850);
and U21959 (N_21959,N_21420,N_21287);
and U21960 (N_21960,N_20594,N_20780);
nor U21961 (N_21961,N_20855,N_21148);
nand U21962 (N_21962,N_21440,N_21030);
or U21963 (N_21963,N_20962,N_21187);
and U21964 (N_21964,N_20869,N_21194);
nor U21965 (N_21965,N_21539,N_20415);
nor U21966 (N_21966,N_21029,N_20538);
and U21967 (N_21967,N_21036,N_20882);
or U21968 (N_21968,N_20935,N_20819);
xnor U21969 (N_21969,N_20812,N_21034);
xnor U21970 (N_21970,N_21387,N_21397);
or U21971 (N_21971,N_20720,N_20897);
xor U21972 (N_21972,N_20989,N_21210);
nand U21973 (N_21973,N_21487,N_21310);
xor U21974 (N_21974,N_20493,N_21229);
or U21975 (N_21975,N_21178,N_21078);
nand U21976 (N_21976,N_20453,N_20733);
and U21977 (N_21977,N_20534,N_21390);
nand U21978 (N_21978,N_20971,N_20892);
nor U21979 (N_21979,N_21089,N_20790);
nand U21980 (N_21980,N_21128,N_21553);
nor U21981 (N_21981,N_21191,N_20827);
xor U21982 (N_21982,N_20486,N_20844);
xnor U21983 (N_21983,N_21233,N_20714);
or U21984 (N_21984,N_20702,N_20711);
xnor U21985 (N_21985,N_21453,N_21061);
nand U21986 (N_21986,N_21238,N_20480);
nand U21987 (N_21987,N_21589,N_21258);
or U21988 (N_21988,N_21518,N_21071);
xnor U21989 (N_21989,N_21320,N_20451);
and U21990 (N_21990,N_20657,N_21542);
and U21991 (N_21991,N_21028,N_20577);
nand U21992 (N_21992,N_21464,N_20803);
or U21993 (N_21993,N_21020,N_20525);
nand U21994 (N_21994,N_21529,N_20941);
xor U21995 (N_21995,N_20956,N_21335);
xnor U21996 (N_21996,N_21185,N_20889);
xnor U21997 (N_21997,N_21429,N_20993);
xnor U21998 (N_21998,N_21117,N_20626);
nor U21999 (N_21999,N_20455,N_21014);
nand U22000 (N_22000,N_21319,N_21276);
nand U22001 (N_22001,N_21115,N_21159);
or U22002 (N_22002,N_21436,N_20952);
nand U22003 (N_22003,N_21047,N_21067);
or U22004 (N_22004,N_20965,N_20782);
nand U22005 (N_22005,N_20665,N_21423);
nand U22006 (N_22006,N_20583,N_21166);
or U22007 (N_22007,N_21073,N_20496);
and U22008 (N_22008,N_21220,N_21549);
xnor U22009 (N_22009,N_20677,N_21240);
or U22010 (N_22010,N_20797,N_21348);
and U22011 (N_22011,N_20447,N_20903);
xor U22012 (N_22012,N_21068,N_21333);
nand U22013 (N_22013,N_20556,N_20853);
and U22014 (N_22014,N_21095,N_20981);
nand U22015 (N_22015,N_21076,N_20785);
nor U22016 (N_22016,N_21473,N_21308);
nor U22017 (N_22017,N_21591,N_21544);
nand U22018 (N_22018,N_20403,N_20427);
or U22019 (N_22019,N_20622,N_20508);
nand U22020 (N_22020,N_21032,N_21472);
or U22021 (N_22021,N_21146,N_20821);
or U22022 (N_22022,N_21293,N_21234);
or U22023 (N_22023,N_20548,N_21225);
and U22024 (N_22024,N_21461,N_21358);
or U22025 (N_22025,N_21449,N_21318);
or U22026 (N_22026,N_20452,N_21522);
or U22027 (N_22027,N_21186,N_21264);
nand U22028 (N_22028,N_21323,N_21002);
and U22029 (N_22029,N_21511,N_21304);
or U22030 (N_22030,N_20549,N_21566);
nand U22031 (N_22031,N_21378,N_20996);
nor U22032 (N_22032,N_21031,N_21119);
xor U22033 (N_22033,N_20954,N_20823);
nor U22034 (N_22034,N_20807,N_20687);
and U22035 (N_22035,N_21062,N_21537);
nor U22036 (N_22036,N_20572,N_20862);
nor U22037 (N_22037,N_21155,N_21056);
nand U22038 (N_22038,N_21143,N_21554);
xor U22039 (N_22039,N_20550,N_20872);
nand U22040 (N_22040,N_20918,N_21283);
nor U22041 (N_22041,N_20988,N_20721);
or U22042 (N_22042,N_20975,N_20964);
and U22043 (N_22043,N_21506,N_20446);
nand U22044 (N_22044,N_20692,N_21289);
or U22045 (N_22045,N_20519,N_20766);
or U22046 (N_22046,N_20639,N_21167);
nor U22047 (N_22047,N_20849,N_20579);
xor U22048 (N_22048,N_21503,N_21513);
nor U22049 (N_22049,N_20586,N_20636);
or U22050 (N_22050,N_21212,N_20973);
or U22051 (N_22051,N_21058,N_20597);
nor U22052 (N_22052,N_20564,N_20816);
nor U22053 (N_22053,N_20842,N_20946);
xor U22054 (N_22054,N_21263,N_21301);
and U22055 (N_22055,N_21471,N_20682);
nor U22056 (N_22056,N_21046,N_20425);
or U22057 (N_22057,N_20592,N_21298);
nor U22058 (N_22058,N_21097,N_20576);
nand U22059 (N_22059,N_21179,N_21559);
and U22060 (N_22060,N_20748,N_21369);
and U22061 (N_22061,N_20690,N_21479);
nand U22062 (N_22062,N_20423,N_21033);
xnor U22063 (N_22063,N_21149,N_21010);
nand U22064 (N_22064,N_21038,N_21523);
or U22065 (N_22065,N_21381,N_20811);
xor U22066 (N_22066,N_20999,N_21441);
xor U22067 (N_22067,N_21093,N_20584);
and U22068 (N_22068,N_20466,N_20407);
nor U22069 (N_22069,N_21239,N_21415);
xnor U22070 (N_22070,N_20708,N_20986);
and U22071 (N_22071,N_20465,N_21411);
nor U22072 (N_22072,N_20979,N_21576);
and U22073 (N_22073,N_21403,N_20871);
nand U22074 (N_22074,N_20740,N_20906);
nand U22075 (N_22075,N_20915,N_20908);
nor U22076 (N_22076,N_20587,N_21203);
nor U22077 (N_22077,N_20410,N_20873);
xor U22078 (N_22078,N_20775,N_21538);
nor U22079 (N_22079,N_21408,N_21476);
nor U22080 (N_22080,N_21406,N_20716);
nor U22081 (N_22081,N_21108,N_21226);
xor U22082 (N_22082,N_21431,N_20633);
nor U22083 (N_22083,N_21416,N_20902);
nor U22084 (N_22084,N_21468,N_20417);
or U22085 (N_22085,N_21161,N_21434);
and U22086 (N_22086,N_20864,N_21274);
or U22087 (N_22087,N_21170,N_21295);
and U22088 (N_22088,N_21399,N_20805);
nor U22089 (N_22089,N_20728,N_20463);
nand U22090 (N_22090,N_21281,N_20727);
nand U22091 (N_22091,N_20751,N_21114);
nor U22092 (N_22092,N_20523,N_20655);
nor U22093 (N_22093,N_21053,N_21292);
nor U22094 (N_22094,N_21245,N_21151);
and U22095 (N_22095,N_20422,N_20507);
nand U22096 (N_22096,N_20568,N_20854);
or U22097 (N_22097,N_21336,N_20913);
xor U22098 (N_22098,N_20445,N_21251);
nor U22099 (N_22099,N_20693,N_20492);
nand U22100 (N_22100,N_20591,N_21572);
and U22101 (N_22101,N_20509,N_21222);
or U22102 (N_22102,N_20943,N_21277);
nand U22103 (N_22103,N_20454,N_21327);
nand U22104 (N_22104,N_21094,N_20482);
nand U22105 (N_22105,N_20567,N_21290);
and U22106 (N_22106,N_21443,N_21147);
and U22107 (N_22107,N_20866,N_20992);
xor U22108 (N_22108,N_21124,N_21546);
nor U22109 (N_22109,N_20839,N_20553);
or U22110 (N_22110,N_21346,N_20546);
xor U22111 (N_22111,N_20414,N_20686);
xnor U22112 (N_22112,N_21315,N_20497);
nand U22113 (N_22113,N_21120,N_21035);
xor U22114 (N_22114,N_21092,N_20557);
nor U22115 (N_22115,N_21347,N_21482);
nand U22116 (N_22116,N_20890,N_21042);
xnor U22117 (N_22117,N_21508,N_20613);
xor U22118 (N_22118,N_20433,N_21080);
xnor U22119 (N_22119,N_21182,N_21435);
nand U22120 (N_22120,N_20416,N_20774);
nor U22121 (N_22121,N_20602,N_21492);
nand U22122 (N_22122,N_21405,N_21305);
nand U22123 (N_22123,N_20420,N_20914);
nand U22124 (N_22124,N_20858,N_21509);
nand U22125 (N_22125,N_21533,N_20934);
and U22126 (N_22126,N_20763,N_20503);
nor U22127 (N_22127,N_20614,N_21583);
nand U22128 (N_22128,N_20554,N_21183);
xnor U22129 (N_22129,N_20712,N_20953);
xnor U22130 (N_22130,N_20545,N_20881);
nor U22131 (N_22131,N_20944,N_21462);
or U22132 (N_22132,N_21000,N_21256);
xnor U22133 (N_22133,N_21353,N_20800);
nand U22134 (N_22134,N_20624,N_20484);
xnor U22135 (N_22135,N_21562,N_20801);
xnor U22136 (N_22136,N_20860,N_20978);
and U22137 (N_22137,N_21228,N_20726);
nor U22138 (N_22138,N_20685,N_21100);
or U22139 (N_22139,N_21521,N_21012);
nor U22140 (N_22140,N_21376,N_21460);
and U22141 (N_22141,N_20875,N_20923);
nor U22142 (N_22142,N_20843,N_20896);
nand U22143 (N_22143,N_21125,N_21300);
xor U22144 (N_22144,N_21077,N_20998);
and U22145 (N_22145,N_21199,N_21217);
or U22146 (N_22146,N_21393,N_20719);
xor U22147 (N_22147,N_21344,N_21282);
or U22148 (N_22148,N_21350,N_21265);
nor U22149 (N_22149,N_20815,N_21180);
or U22150 (N_22150,N_21489,N_20683);
nand U22151 (N_22151,N_21458,N_20752);
xor U22152 (N_22152,N_20562,N_21190);
nand U22153 (N_22153,N_21484,N_20469);
or U22154 (N_22154,N_20672,N_20691);
nand U22155 (N_22155,N_20788,N_20565);
xnor U22156 (N_22156,N_21515,N_20904);
or U22157 (N_22157,N_20723,N_21528);
nand U22158 (N_22158,N_21006,N_21132);
nor U22159 (N_22159,N_20773,N_20533);
or U22160 (N_22160,N_21454,N_21389);
xor U22161 (N_22161,N_21541,N_20750);
nand U22162 (N_22162,N_20471,N_21446);
nor U22163 (N_22163,N_20590,N_20580);
nor U22164 (N_22164,N_21438,N_20522);
xor U22165 (N_22165,N_20543,N_21558);
and U22166 (N_22166,N_21354,N_20458);
or U22167 (N_22167,N_21536,N_20490);
or U22168 (N_22168,N_20754,N_21162);
and U22169 (N_22169,N_21009,N_20703);
nor U22170 (N_22170,N_21311,N_21235);
nor U22171 (N_22171,N_20688,N_21236);
xnor U22172 (N_22172,N_21571,N_21338);
nand U22173 (N_22173,N_20927,N_21316);
nor U22174 (N_22174,N_20868,N_20791);
nor U22175 (N_22175,N_21065,N_20681);
and U22176 (N_22176,N_21349,N_21447);
nor U22177 (N_22177,N_20669,N_20668);
and U22178 (N_22178,N_21213,N_21556);
xnor U22179 (N_22179,N_20532,N_20880);
nand U22180 (N_22180,N_20651,N_20749);
and U22181 (N_22181,N_20464,N_21568);
nand U22182 (N_22182,N_21437,N_21273);
nand U22183 (N_22183,N_20566,N_21027);
or U22184 (N_22184,N_20521,N_21582);
nand U22185 (N_22185,N_21176,N_21569);
or U22186 (N_22186,N_20421,N_20662);
nor U22187 (N_22187,N_21466,N_20663);
xnor U22188 (N_22188,N_21188,N_21502);
nand U22189 (N_22189,N_20431,N_21328);
nor U22190 (N_22190,N_20635,N_20966);
nor U22191 (N_22191,N_21412,N_20930);
xor U22192 (N_22192,N_21345,N_21422);
nand U22193 (N_22193,N_21004,N_21439);
xor U22194 (N_22194,N_21215,N_20970);
nand U22195 (N_22195,N_21048,N_21246);
nor U22196 (N_22196,N_20829,N_20982);
or U22197 (N_22197,N_21584,N_21463);
or U22198 (N_22198,N_20630,N_20487);
xor U22199 (N_22199,N_21121,N_21297);
nand U22200 (N_22200,N_21060,N_20538);
or U22201 (N_22201,N_21328,N_21448);
or U22202 (N_22202,N_20711,N_21583);
or U22203 (N_22203,N_20874,N_20715);
or U22204 (N_22204,N_20824,N_20717);
and U22205 (N_22205,N_20553,N_20938);
nand U22206 (N_22206,N_20907,N_20942);
nand U22207 (N_22207,N_20751,N_21350);
xnor U22208 (N_22208,N_21087,N_20620);
nand U22209 (N_22209,N_21476,N_20957);
or U22210 (N_22210,N_21556,N_21074);
xor U22211 (N_22211,N_20945,N_20974);
and U22212 (N_22212,N_21454,N_21034);
or U22213 (N_22213,N_21369,N_21221);
and U22214 (N_22214,N_20660,N_21384);
nand U22215 (N_22215,N_20641,N_21251);
and U22216 (N_22216,N_20601,N_21286);
nand U22217 (N_22217,N_21057,N_21322);
nand U22218 (N_22218,N_20628,N_20638);
nor U22219 (N_22219,N_21469,N_21586);
nand U22220 (N_22220,N_21212,N_21185);
nand U22221 (N_22221,N_21028,N_21239);
nor U22222 (N_22222,N_21452,N_21507);
nor U22223 (N_22223,N_20906,N_21307);
nand U22224 (N_22224,N_21520,N_21140);
nor U22225 (N_22225,N_21521,N_20765);
xor U22226 (N_22226,N_20887,N_20968);
nand U22227 (N_22227,N_20964,N_20791);
or U22228 (N_22228,N_21146,N_21488);
and U22229 (N_22229,N_20609,N_20892);
and U22230 (N_22230,N_21576,N_21434);
and U22231 (N_22231,N_20413,N_20594);
nand U22232 (N_22232,N_21303,N_20560);
xnor U22233 (N_22233,N_20739,N_21176);
xor U22234 (N_22234,N_21204,N_20455);
nor U22235 (N_22235,N_21043,N_20440);
and U22236 (N_22236,N_20905,N_21088);
nand U22237 (N_22237,N_21382,N_21012);
or U22238 (N_22238,N_21578,N_20893);
or U22239 (N_22239,N_20425,N_21585);
nand U22240 (N_22240,N_20620,N_20523);
or U22241 (N_22241,N_21480,N_20404);
nand U22242 (N_22242,N_20856,N_20706);
or U22243 (N_22243,N_21309,N_20865);
xnor U22244 (N_22244,N_21362,N_20824);
or U22245 (N_22245,N_21548,N_20540);
nand U22246 (N_22246,N_21475,N_20511);
xnor U22247 (N_22247,N_20791,N_20464);
and U22248 (N_22248,N_21319,N_20504);
and U22249 (N_22249,N_21369,N_20497);
nand U22250 (N_22250,N_20745,N_21546);
xor U22251 (N_22251,N_20871,N_20993);
nand U22252 (N_22252,N_20569,N_20652);
nand U22253 (N_22253,N_20812,N_21025);
nand U22254 (N_22254,N_21368,N_20850);
or U22255 (N_22255,N_20754,N_21415);
xor U22256 (N_22256,N_20645,N_20594);
or U22257 (N_22257,N_21128,N_21201);
or U22258 (N_22258,N_21366,N_20421);
xnor U22259 (N_22259,N_20696,N_21121);
or U22260 (N_22260,N_20510,N_20459);
nand U22261 (N_22261,N_20936,N_20785);
and U22262 (N_22262,N_21070,N_21533);
or U22263 (N_22263,N_21156,N_20730);
nand U22264 (N_22264,N_21040,N_20589);
nand U22265 (N_22265,N_20630,N_21462);
nor U22266 (N_22266,N_20600,N_20826);
and U22267 (N_22267,N_20992,N_20547);
nor U22268 (N_22268,N_21505,N_20821);
and U22269 (N_22269,N_21395,N_21101);
nand U22270 (N_22270,N_21364,N_20803);
nor U22271 (N_22271,N_20631,N_20663);
or U22272 (N_22272,N_21469,N_20987);
nand U22273 (N_22273,N_21381,N_21177);
nor U22274 (N_22274,N_21262,N_21348);
nor U22275 (N_22275,N_21460,N_21375);
or U22276 (N_22276,N_20979,N_21190);
or U22277 (N_22277,N_21394,N_20879);
or U22278 (N_22278,N_21085,N_20922);
and U22279 (N_22279,N_21419,N_20908);
nand U22280 (N_22280,N_21009,N_21177);
and U22281 (N_22281,N_20464,N_20750);
and U22282 (N_22282,N_21105,N_20980);
nand U22283 (N_22283,N_21435,N_21533);
nand U22284 (N_22284,N_20747,N_20509);
or U22285 (N_22285,N_21128,N_20534);
and U22286 (N_22286,N_21043,N_20714);
or U22287 (N_22287,N_21020,N_21562);
or U22288 (N_22288,N_20974,N_20441);
xor U22289 (N_22289,N_20443,N_21196);
xnor U22290 (N_22290,N_21306,N_20537);
xor U22291 (N_22291,N_21161,N_20882);
nor U22292 (N_22292,N_20929,N_20902);
and U22293 (N_22293,N_21055,N_21490);
nor U22294 (N_22294,N_20857,N_21497);
xor U22295 (N_22295,N_21140,N_21493);
or U22296 (N_22296,N_21094,N_20839);
nand U22297 (N_22297,N_20807,N_21436);
or U22298 (N_22298,N_20832,N_20752);
and U22299 (N_22299,N_21058,N_21208);
and U22300 (N_22300,N_21428,N_21595);
or U22301 (N_22301,N_20434,N_20875);
and U22302 (N_22302,N_21145,N_20565);
and U22303 (N_22303,N_20549,N_20820);
or U22304 (N_22304,N_21203,N_20936);
and U22305 (N_22305,N_21236,N_20958);
or U22306 (N_22306,N_20684,N_21172);
or U22307 (N_22307,N_20651,N_21155);
and U22308 (N_22308,N_21576,N_21518);
nand U22309 (N_22309,N_21298,N_21426);
nor U22310 (N_22310,N_20869,N_21085);
or U22311 (N_22311,N_21355,N_21467);
xor U22312 (N_22312,N_20524,N_21017);
xnor U22313 (N_22313,N_20972,N_20434);
and U22314 (N_22314,N_21091,N_20775);
xnor U22315 (N_22315,N_20648,N_20621);
nand U22316 (N_22316,N_20766,N_20564);
nand U22317 (N_22317,N_20453,N_21334);
nand U22318 (N_22318,N_20792,N_21083);
nor U22319 (N_22319,N_20897,N_20732);
or U22320 (N_22320,N_20766,N_21242);
xnor U22321 (N_22321,N_20558,N_21009);
and U22322 (N_22322,N_20948,N_21287);
xor U22323 (N_22323,N_21373,N_21432);
nand U22324 (N_22324,N_20610,N_21264);
or U22325 (N_22325,N_21230,N_20517);
nor U22326 (N_22326,N_20607,N_21290);
and U22327 (N_22327,N_20661,N_21076);
and U22328 (N_22328,N_20962,N_20853);
nand U22329 (N_22329,N_20569,N_20590);
nor U22330 (N_22330,N_20447,N_20503);
xor U22331 (N_22331,N_21347,N_20755);
nor U22332 (N_22332,N_20947,N_21089);
nand U22333 (N_22333,N_20644,N_20820);
and U22334 (N_22334,N_20521,N_20763);
nand U22335 (N_22335,N_20791,N_20857);
or U22336 (N_22336,N_20630,N_20564);
xnor U22337 (N_22337,N_20671,N_20504);
xor U22338 (N_22338,N_21172,N_20655);
nor U22339 (N_22339,N_20472,N_20545);
or U22340 (N_22340,N_20868,N_21184);
nand U22341 (N_22341,N_20788,N_20887);
or U22342 (N_22342,N_21219,N_21417);
nand U22343 (N_22343,N_21293,N_20518);
nor U22344 (N_22344,N_21205,N_20596);
nor U22345 (N_22345,N_20412,N_21146);
xnor U22346 (N_22346,N_21048,N_20421);
xnor U22347 (N_22347,N_21127,N_21328);
and U22348 (N_22348,N_21213,N_20889);
nand U22349 (N_22349,N_21054,N_21533);
nor U22350 (N_22350,N_20766,N_21410);
and U22351 (N_22351,N_20610,N_21177);
nor U22352 (N_22352,N_20649,N_21025);
nor U22353 (N_22353,N_21090,N_20502);
or U22354 (N_22354,N_21388,N_20733);
nor U22355 (N_22355,N_20685,N_20984);
or U22356 (N_22356,N_21322,N_21344);
or U22357 (N_22357,N_20844,N_20892);
nor U22358 (N_22358,N_20706,N_20629);
nor U22359 (N_22359,N_21473,N_21544);
xor U22360 (N_22360,N_21386,N_20547);
nor U22361 (N_22361,N_20823,N_21587);
and U22362 (N_22362,N_20698,N_21330);
and U22363 (N_22363,N_20684,N_21227);
or U22364 (N_22364,N_20994,N_20638);
and U22365 (N_22365,N_21178,N_21195);
nand U22366 (N_22366,N_20777,N_20804);
xor U22367 (N_22367,N_20649,N_21003);
nor U22368 (N_22368,N_21545,N_21056);
xor U22369 (N_22369,N_20439,N_20956);
nor U22370 (N_22370,N_20953,N_20453);
nand U22371 (N_22371,N_21582,N_21473);
nand U22372 (N_22372,N_21445,N_21067);
xnor U22373 (N_22373,N_21050,N_20571);
xor U22374 (N_22374,N_20501,N_20464);
nand U22375 (N_22375,N_21496,N_20455);
nor U22376 (N_22376,N_20843,N_21465);
and U22377 (N_22377,N_20877,N_20864);
xnor U22378 (N_22378,N_21108,N_21507);
nand U22379 (N_22379,N_21128,N_20940);
xnor U22380 (N_22380,N_20510,N_20432);
nand U22381 (N_22381,N_20707,N_20594);
and U22382 (N_22382,N_21004,N_21218);
nand U22383 (N_22383,N_20903,N_21474);
or U22384 (N_22384,N_21111,N_21088);
xor U22385 (N_22385,N_21043,N_21590);
and U22386 (N_22386,N_20903,N_21059);
nand U22387 (N_22387,N_20463,N_20676);
nor U22388 (N_22388,N_20890,N_21517);
nand U22389 (N_22389,N_21485,N_21342);
or U22390 (N_22390,N_21294,N_20474);
nand U22391 (N_22391,N_20871,N_21120);
nor U22392 (N_22392,N_20603,N_21557);
and U22393 (N_22393,N_21069,N_20710);
nor U22394 (N_22394,N_20490,N_20503);
nand U22395 (N_22395,N_20616,N_20593);
xnor U22396 (N_22396,N_21306,N_21465);
nor U22397 (N_22397,N_20885,N_21538);
nor U22398 (N_22398,N_20966,N_21318);
or U22399 (N_22399,N_21540,N_20549);
xor U22400 (N_22400,N_20754,N_21485);
or U22401 (N_22401,N_20421,N_21418);
xnor U22402 (N_22402,N_21486,N_20734);
nand U22403 (N_22403,N_21004,N_21253);
nor U22404 (N_22404,N_20897,N_20746);
xor U22405 (N_22405,N_20628,N_21268);
or U22406 (N_22406,N_20593,N_20524);
and U22407 (N_22407,N_21111,N_21131);
nand U22408 (N_22408,N_20877,N_20656);
and U22409 (N_22409,N_21597,N_21346);
xor U22410 (N_22410,N_21454,N_20664);
nor U22411 (N_22411,N_21316,N_21145);
and U22412 (N_22412,N_20962,N_20473);
xnor U22413 (N_22413,N_21492,N_20521);
and U22414 (N_22414,N_20635,N_20510);
nand U22415 (N_22415,N_20435,N_20523);
and U22416 (N_22416,N_20665,N_21550);
nor U22417 (N_22417,N_21294,N_21087);
nand U22418 (N_22418,N_21561,N_20873);
nor U22419 (N_22419,N_21376,N_20530);
and U22420 (N_22420,N_20531,N_20863);
and U22421 (N_22421,N_21400,N_20630);
xnor U22422 (N_22422,N_21351,N_21288);
or U22423 (N_22423,N_20521,N_21309);
or U22424 (N_22424,N_21015,N_20997);
xor U22425 (N_22425,N_20465,N_20428);
and U22426 (N_22426,N_20474,N_20746);
nor U22427 (N_22427,N_20751,N_21475);
nor U22428 (N_22428,N_21282,N_21356);
nand U22429 (N_22429,N_21206,N_20882);
and U22430 (N_22430,N_20502,N_20761);
nand U22431 (N_22431,N_21408,N_20834);
nor U22432 (N_22432,N_20493,N_21195);
or U22433 (N_22433,N_20530,N_20724);
and U22434 (N_22434,N_20758,N_20441);
xnor U22435 (N_22435,N_20873,N_21514);
nor U22436 (N_22436,N_21398,N_21342);
or U22437 (N_22437,N_20725,N_20744);
and U22438 (N_22438,N_21586,N_20902);
nor U22439 (N_22439,N_20746,N_21066);
or U22440 (N_22440,N_20848,N_20670);
nor U22441 (N_22441,N_20859,N_20704);
or U22442 (N_22442,N_20573,N_20945);
xor U22443 (N_22443,N_21551,N_21307);
nand U22444 (N_22444,N_20677,N_21307);
nor U22445 (N_22445,N_20563,N_20661);
xor U22446 (N_22446,N_21585,N_21446);
and U22447 (N_22447,N_21439,N_21280);
or U22448 (N_22448,N_20993,N_20818);
and U22449 (N_22449,N_21190,N_21557);
and U22450 (N_22450,N_20489,N_21285);
xnor U22451 (N_22451,N_20501,N_21364);
xnor U22452 (N_22452,N_20565,N_20753);
and U22453 (N_22453,N_20898,N_21210);
and U22454 (N_22454,N_21000,N_20409);
and U22455 (N_22455,N_21179,N_21294);
xor U22456 (N_22456,N_21540,N_21320);
nand U22457 (N_22457,N_21217,N_20804);
nor U22458 (N_22458,N_21464,N_20860);
xor U22459 (N_22459,N_21463,N_20884);
or U22460 (N_22460,N_21262,N_20539);
nor U22461 (N_22461,N_20435,N_21388);
nor U22462 (N_22462,N_20450,N_21051);
xnor U22463 (N_22463,N_20758,N_21575);
nand U22464 (N_22464,N_21371,N_21475);
nor U22465 (N_22465,N_21014,N_20807);
and U22466 (N_22466,N_21327,N_21207);
and U22467 (N_22467,N_20824,N_20435);
or U22468 (N_22468,N_20609,N_21214);
xor U22469 (N_22469,N_20477,N_20820);
nand U22470 (N_22470,N_20878,N_21428);
xor U22471 (N_22471,N_20914,N_20521);
and U22472 (N_22472,N_21326,N_20794);
nand U22473 (N_22473,N_20587,N_20542);
nand U22474 (N_22474,N_21241,N_21472);
nor U22475 (N_22475,N_20523,N_21441);
or U22476 (N_22476,N_21497,N_21147);
and U22477 (N_22477,N_21378,N_20908);
and U22478 (N_22478,N_20535,N_20874);
xnor U22479 (N_22479,N_20736,N_21471);
xor U22480 (N_22480,N_20999,N_20696);
or U22481 (N_22481,N_21379,N_21215);
and U22482 (N_22482,N_21523,N_20493);
nand U22483 (N_22483,N_20641,N_21435);
nand U22484 (N_22484,N_20448,N_21064);
xor U22485 (N_22485,N_20486,N_20744);
or U22486 (N_22486,N_20584,N_20777);
xnor U22487 (N_22487,N_20813,N_20593);
and U22488 (N_22488,N_21080,N_20847);
and U22489 (N_22489,N_21427,N_21015);
and U22490 (N_22490,N_21578,N_20864);
or U22491 (N_22491,N_20647,N_21158);
nand U22492 (N_22492,N_21358,N_20552);
nand U22493 (N_22493,N_20818,N_21542);
nor U22494 (N_22494,N_20690,N_21460);
nor U22495 (N_22495,N_21390,N_20714);
or U22496 (N_22496,N_20612,N_20442);
xor U22497 (N_22497,N_20991,N_20541);
and U22498 (N_22498,N_20504,N_20708);
or U22499 (N_22499,N_20471,N_21164);
and U22500 (N_22500,N_21460,N_21513);
and U22501 (N_22501,N_21008,N_20551);
and U22502 (N_22502,N_20769,N_20705);
nor U22503 (N_22503,N_21270,N_21462);
xnor U22504 (N_22504,N_21293,N_20839);
xnor U22505 (N_22505,N_20998,N_21397);
or U22506 (N_22506,N_20781,N_20738);
xnor U22507 (N_22507,N_21339,N_21080);
or U22508 (N_22508,N_21362,N_20751);
and U22509 (N_22509,N_21082,N_20957);
and U22510 (N_22510,N_20414,N_20775);
nor U22511 (N_22511,N_21477,N_20783);
nand U22512 (N_22512,N_20545,N_20846);
nor U22513 (N_22513,N_21185,N_21391);
and U22514 (N_22514,N_20793,N_21491);
or U22515 (N_22515,N_21217,N_21096);
nor U22516 (N_22516,N_20543,N_20924);
and U22517 (N_22517,N_21361,N_21565);
and U22518 (N_22518,N_20655,N_21063);
nor U22519 (N_22519,N_20457,N_20931);
xnor U22520 (N_22520,N_21176,N_21071);
xor U22521 (N_22521,N_21375,N_20858);
and U22522 (N_22522,N_20542,N_21153);
xor U22523 (N_22523,N_21289,N_20966);
or U22524 (N_22524,N_21567,N_20855);
nand U22525 (N_22525,N_21580,N_21508);
and U22526 (N_22526,N_20472,N_20905);
nand U22527 (N_22527,N_20672,N_21115);
nor U22528 (N_22528,N_20866,N_20898);
nand U22529 (N_22529,N_20848,N_20711);
or U22530 (N_22530,N_21084,N_20629);
or U22531 (N_22531,N_20678,N_21161);
and U22532 (N_22532,N_21442,N_21488);
xor U22533 (N_22533,N_20831,N_21499);
nor U22534 (N_22534,N_21534,N_21591);
or U22535 (N_22535,N_21154,N_21238);
nand U22536 (N_22536,N_20420,N_21096);
or U22537 (N_22537,N_20523,N_20680);
or U22538 (N_22538,N_21597,N_20558);
and U22539 (N_22539,N_21484,N_20491);
xor U22540 (N_22540,N_21340,N_20696);
xnor U22541 (N_22541,N_21213,N_20691);
nand U22542 (N_22542,N_20491,N_20721);
nor U22543 (N_22543,N_21474,N_20559);
or U22544 (N_22544,N_20400,N_20659);
or U22545 (N_22545,N_20694,N_21352);
nor U22546 (N_22546,N_21280,N_20781);
nand U22547 (N_22547,N_20694,N_20858);
and U22548 (N_22548,N_21354,N_21321);
xor U22549 (N_22549,N_21492,N_20618);
nor U22550 (N_22550,N_21508,N_20930);
nand U22551 (N_22551,N_20756,N_21087);
and U22552 (N_22552,N_20449,N_20531);
or U22553 (N_22553,N_21498,N_20822);
and U22554 (N_22554,N_20508,N_20869);
nor U22555 (N_22555,N_20464,N_21494);
xnor U22556 (N_22556,N_20807,N_21006);
nor U22557 (N_22557,N_20782,N_20728);
or U22558 (N_22558,N_21245,N_20768);
nor U22559 (N_22559,N_21407,N_20688);
and U22560 (N_22560,N_21366,N_20780);
or U22561 (N_22561,N_20424,N_20806);
nand U22562 (N_22562,N_21039,N_20789);
and U22563 (N_22563,N_20980,N_20505);
and U22564 (N_22564,N_20847,N_20920);
and U22565 (N_22565,N_20731,N_20644);
nor U22566 (N_22566,N_20617,N_20952);
nor U22567 (N_22567,N_20463,N_20610);
nor U22568 (N_22568,N_20847,N_21102);
nand U22569 (N_22569,N_20567,N_21557);
nand U22570 (N_22570,N_20665,N_21125);
nand U22571 (N_22571,N_21205,N_21181);
xor U22572 (N_22572,N_20783,N_21461);
nor U22573 (N_22573,N_21301,N_21078);
nand U22574 (N_22574,N_20616,N_21331);
nand U22575 (N_22575,N_21279,N_20690);
nor U22576 (N_22576,N_20687,N_20835);
and U22577 (N_22577,N_21546,N_20844);
nor U22578 (N_22578,N_20552,N_21137);
xor U22579 (N_22579,N_20867,N_21092);
xnor U22580 (N_22580,N_20604,N_20880);
nor U22581 (N_22581,N_20602,N_21275);
nand U22582 (N_22582,N_21255,N_21318);
and U22583 (N_22583,N_20663,N_20699);
or U22584 (N_22584,N_21385,N_21190);
or U22585 (N_22585,N_21487,N_20666);
nand U22586 (N_22586,N_21068,N_20556);
nand U22587 (N_22587,N_20898,N_21074);
nor U22588 (N_22588,N_20951,N_21263);
nand U22589 (N_22589,N_20539,N_20501);
or U22590 (N_22590,N_21432,N_21597);
and U22591 (N_22591,N_21108,N_21207);
and U22592 (N_22592,N_21431,N_21229);
or U22593 (N_22593,N_20567,N_21034);
or U22594 (N_22594,N_20933,N_20599);
xnor U22595 (N_22595,N_20498,N_20662);
or U22596 (N_22596,N_21432,N_21288);
and U22597 (N_22597,N_21325,N_20755);
or U22598 (N_22598,N_20776,N_20729);
xnor U22599 (N_22599,N_21295,N_20576);
nand U22600 (N_22600,N_20599,N_20943);
nand U22601 (N_22601,N_21427,N_20920);
or U22602 (N_22602,N_21489,N_21519);
nor U22603 (N_22603,N_20940,N_20587);
nor U22604 (N_22604,N_20786,N_21011);
nor U22605 (N_22605,N_21522,N_21211);
nor U22606 (N_22606,N_21072,N_20706);
nor U22607 (N_22607,N_20751,N_21082);
nand U22608 (N_22608,N_20872,N_21152);
and U22609 (N_22609,N_20453,N_21215);
nand U22610 (N_22610,N_21442,N_21436);
and U22611 (N_22611,N_20738,N_20720);
and U22612 (N_22612,N_21173,N_21567);
and U22613 (N_22613,N_21006,N_20747);
nand U22614 (N_22614,N_21198,N_20412);
nor U22615 (N_22615,N_20494,N_21022);
nand U22616 (N_22616,N_20545,N_21201);
nand U22617 (N_22617,N_20464,N_20638);
nand U22618 (N_22618,N_21159,N_20718);
nor U22619 (N_22619,N_20846,N_20543);
xnor U22620 (N_22620,N_20421,N_21358);
xor U22621 (N_22621,N_21147,N_21032);
xor U22622 (N_22622,N_21512,N_21078);
xnor U22623 (N_22623,N_20822,N_21472);
or U22624 (N_22624,N_20629,N_20686);
xor U22625 (N_22625,N_20877,N_21598);
or U22626 (N_22626,N_20934,N_21542);
xor U22627 (N_22627,N_20652,N_21146);
or U22628 (N_22628,N_20841,N_21220);
nand U22629 (N_22629,N_21550,N_20437);
or U22630 (N_22630,N_21247,N_20578);
xnor U22631 (N_22631,N_21319,N_20804);
xnor U22632 (N_22632,N_20835,N_21193);
or U22633 (N_22633,N_20909,N_20474);
or U22634 (N_22634,N_21219,N_20850);
nor U22635 (N_22635,N_20601,N_20718);
nand U22636 (N_22636,N_20664,N_20754);
nor U22637 (N_22637,N_21332,N_21493);
nor U22638 (N_22638,N_21003,N_21414);
nand U22639 (N_22639,N_21564,N_21443);
or U22640 (N_22640,N_21147,N_20546);
nand U22641 (N_22641,N_20564,N_21431);
nand U22642 (N_22642,N_20936,N_20438);
nand U22643 (N_22643,N_21040,N_20789);
and U22644 (N_22644,N_20868,N_21368);
nand U22645 (N_22645,N_20752,N_21134);
xnor U22646 (N_22646,N_21280,N_20593);
xnor U22647 (N_22647,N_21576,N_20827);
nor U22648 (N_22648,N_20687,N_20469);
nand U22649 (N_22649,N_21262,N_21583);
xnor U22650 (N_22650,N_21191,N_20819);
xor U22651 (N_22651,N_20938,N_21318);
xnor U22652 (N_22652,N_21465,N_20836);
and U22653 (N_22653,N_20403,N_21073);
nor U22654 (N_22654,N_20796,N_21254);
or U22655 (N_22655,N_21146,N_21415);
or U22656 (N_22656,N_21444,N_21583);
xor U22657 (N_22657,N_21218,N_21484);
or U22658 (N_22658,N_21586,N_21136);
nand U22659 (N_22659,N_20898,N_21083);
nand U22660 (N_22660,N_21281,N_20566);
or U22661 (N_22661,N_20965,N_21341);
and U22662 (N_22662,N_21545,N_21596);
nor U22663 (N_22663,N_20757,N_21374);
nor U22664 (N_22664,N_21460,N_21093);
or U22665 (N_22665,N_21470,N_21397);
nand U22666 (N_22666,N_21108,N_20500);
or U22667 (N_22667,N_20889,N_20696);
and U22668 (N_22668,N_20481,N_20432);
nand U22669 (N_22669,N_20501,N_20526);
xor U22670 (N_22670,N_21010,N_20481);
nand U22671 (N_22671,N_20542,N_21251);
nand U22672 (N_22672,N_20592,N_20980);
nor U22673 (N_22673,N_20498,N_21474);
xor U22674 (N_22674,N_20445,N_20416);
nor U22675 (N_22675,N_20494,N_20724);
nor U22676 (N_22676,N_20957,N_21000);
and U22677 (N_22677,N_20797,N_21436);
xor U22678 (N_22678,N_20881,N_20905);
xor U22679 (N_22679,N_21068,N_21340);
or U22680 (N_22680,N_21071,N_21334);
and U22681 (N_22681,N_21106,N_20976);
or U22682 (N_22682,N_20589,N_21144);
nor U22683 (N_22683,N_21284,N_21169);
and U22684 (N_22684,N_20916,N_21026);
or U22685 (N_22685,N_20858,N_21250);
nand U22686 (N_22686,N_20886,N_20860);
nor U22687 (N_22687,N_20941,N_21324);
or U22688 (N_22688,N_21296,N_21163);
nand U22689 (N_22689,N_21538,N_20742);
or U22690 (N_22690,N_20907,N_21514);
nor U22691 (N_22691,N_20651,N_21286);
or U22692 (N_22692,N_20621,N_21245);
xnor U22693 (N_22693,N_21069,N_21001);
or U22694 (N_22694,N_20860,N_20898);
or U22695 (N_22695,N_21085,N_21416);
or U22696 (N_22696,N_21226,N_21164);
and U22697 (N_22697,N_20808,N_20693);
nand U22698 (N_22698,N_21305,N_20673);
and U22699 (N_22699,N_20849,N_20897);
nor U22700 (N_22700,N_21399,N_21071);
and U22701 (N_22701,N_21118,N_21315);
or U22702 (N_22702,N_20580,N_20751);
or U22703 (N_22703,N_21468,N_20939);
xor U22704 (N_22704,N_21110,N_20892);
and U22705 (N_22705,N_21264,N_20431);
xnor U22706 (N_22706,N_21392,N_21056);
nand U22707 (N_22707,N_20798,N_20712);
xor U22708 (N_22708,N_20459,N_20521);
xor U22709 (N_22709,N_21254,N_21030);
xnor U22710 (N_22710,N_20678,N_20623);
and U22711 (N_22711,N_20859,N_21473);
nand U22712 (N_22712,N_20815,N_21319);
nor U22713 (N_22713,N_20528,N_21109);
xnor U22714 (N_22714,N_20766,N_20786);
or U22715 (N_22715,N_21430,N_21291);
nor U22716 (N_22716,N_21510,N_20889);
nor U22717 (N_22717,N_21539,N_20585);
or U22718 (N_22718,N_21439,N_21317);
nor U22719 (N_22719,N_21139,N_20971);
nor U22720 (N_22720,N_21225,N_20872);
nor U22721 (N_22721,N_20520,N_21304);
or U22722 (N_22722,N_21075,N_20789);
nor U22723 (N_22723,N_20585,N_21295);
nand U22724 (N_22724,N_21198,N_20865);
or U22725 (N_22725,N_20440,N_21269);
and U22726 (N_22726,N_21228,N_20452);
nor U22727 (N_22727,N_21393,N_20490);
or U22728 (N_22728,N_21357,N_20498);
nand U22729 (N_22729,N_20553,N_21017);
and U22730 (N_22730,N_20788,N_20634);
and U22731 (N_22731,N_20705,N_21571);
or U22732 (N_22732,N_20772,N_20795);
nand U22733 (N_22733,N_20472,N_21378);
xnor U22734 (N_22734,N_21100,N_20573);
xnor U22735 (N_22735,N_20730,N_21074);
nor U22736 (N_22736,N_20851,N_20553);
and U22737 (N_22737,N_21467,N_21406);
and U22738 (N_22738,N_20617,N_21215);
or U22739 (N_22739,N_21049,N_21195);
or U22740 (N_22740,N_20722,N_20602);
and U22741 (N_22741,N_20556,N_21392);
or U22742 (N_22742,N_21008,N_20651);
nand U22743 (N_22743,N_20671,N_21072);
xor U22744 (N_22744,N_21333,N_21597);
nand U22745 (N_22745,N_21458,N_21248);
and U22746 (N_22746,N_20523,N_20991);
and U22747 (N_22747,N_20839,N_21153);
xor U22748 (N_22748,N_20504,N_21347);
nand U22749 (N_22749,N_20704,N_21442);
or U22750 (N_22750,N_21159,N_20459);
or U22751 (N_22751,N_21231,N_21535);
nor U22752 (N_22752,N_21282,N_20516);
and U22753 (N_22753,N_21088,N_21235);
xor U22754 (N_22754,N_20704,N_21587);
or U22755 (N_22755,N_21234,N_20427);
xnor U22756 (N_22756,N_21355,N_21308);
or U22757 (N_22757,N_21068,N_21442);
and U22758 (N_22758,N_21569,N_21415);
nor U22759 (N_22759,N_20887,N_20485);
and U22760 (N_22760,N_21348,N_20533);
nand U22761 (N_22761,N_20405,N_21510);
nand U22762 (N_22762,N_20798,N_20496);
xor U22763 (N_22763,N_21013,N_21400);
or U22764 (N_22764,N_20525,N_20592);
nor U22765 (N_22765,N_21446,N_20570);
nand U22766 (N_22766,N_21504,N_20724);
nand U22767 (N_22767,N_20884,N_21237);
nand U22768 (N_22768,N_21345,N_21327);
and U22769 (N_22769,N_20599,N_21121);
and U22770 (N_22770,N_20997,N_21522);
or U22771 (N_22771,N_21111,N_21358);
xnor U22772 (N_22772,N_21197,N_20501);
xor U22773 (N_22773,N_20885,N_20685);
xnor U22774 (N_22774,N_21594,N_21585);
nor U22775 (N_22775,N_21458,N_20589);
nor U22776 (N_22776,N_21458,N_20644);
nand U22777 (N_22777,N_20685,N_21115);
nor U22778 (N_22778,N_21428,N_21308);
and U22779 (N_22779,N_20622,N_20635);
or U22780 (N_22780,N_21542,N_20583);
or U22781 (N_22781,N_21166,N_20577);
or U22782 (N_22782,N_20672,N_20981);
and U22783 (N_22783,N_20681,N_20883);
nand U22784 (N_22784,N_21350,N_20456);
and U22785 (N_22785,N_20948,N_20525);
or U22786 (N_22786,N_21307,N_20860);
nor U22787 (N_22787,N_20589,N_21494);
nor U22788 (N_22788,N_20777,N_20685);
xnor U22789 (N_22789,N_21309,N_21415);
and U22790 (N_22790,N_20692,N_20583);
xnor U22791 (N_22791,N_20809,N_20916);
nand U22792 (N_22792,N_20886,N_21115);
nor U22793 (N_22793,N_21318,N_21018);
nor U22794 (N_22794,N_20916,N_21350);
nor U22795 (N_22795,N_20723,N_21247);
nand U22796 (N_22796,N_21217,N_20555);
xnor U22797 (N_22797,N_20968,N_20501);
or U22798 (N_22798,N_20552,N_20528);
or U22799 (N_22799,N_21560,N_21301);
nand U22800 (N_22800,N_22140,N_22541);
nor U22801 (N_22801,N_21896,N_22710);
and U22802 (N_22802,N_22186,N_21907);
and U22803 (N_22803,N_22074,N_22169);
nand U22804 (N_22804,N_22361,N_21842);
nand U22805 (N_22805,N_21795,N_22332);
and U22806 (N_22806,N_22257,N_22765);
nor U22807 (N_22807,N_22194,N_22201);
or U22808 (N_22808,N_21886,N_22077);
nor U22809 (N_22809,N_21669,N_22364);
xor U22810 (N_22810,N_22663,N_21953);
xor U22811 (N_22811,N_22320,N_22350);
or U22812 (N_22812,N_22282,N_22358);
and U22813 (N_22813,N_21961,N_21736);
and U22814 (N_22814,N_21879,N_22637);
nand U22815 (N_22815,N_22090,N_22153);
nand U22816 (N_22816,N_22382,N_21860);
xor U22817 (N_22817,N_22393,N_22344);
nor U22818 (N_22818,N_21902,N_22500);
xnor U22819 (N_22819,N_21648,N_21625);
xor U22820 (N_22820,N_22219,N_22260);
xnor U22821 (N_22821,N_22609,N_22235);
or U22822 (N_22822,N_21831,N_22237);
or U22823 (N_22823,N_22240,N_21812);
or U22824 (N_22824,N_21634,N_21877);
and U22825 (N_22825,N_21710,N_22189);
nand U22826 (N_22826,N_22013,N_22433);
nand U22827 (N_22827,N_21770,N_21702);
xnor U22828 (N_22828,N_22322,N_22071);
nor U22829 (N_22829,N_21999,N_22404);
nor U22830 (N_22830,N_22399,N_22751);
and U22831 (N_22831,N_22587,N_21682);
nand U22832 (N_22832,N_22111,N_22618);
nor U22833 (N_22833,N_22175,N_22577);
nand U22834 (N_22834,N_21765,N_21743);
xor U22835 (N_22835,N_22760,N_22634);
xor U22836 (N_22836,N_21676,N_22231);
nor U22837 (N_22837,N_21618,N_22465);
nor U22838 (N_22838,N_22308,N_22655);
nand U22839 (N_22839,N_21607,N_22701);
nor U22840 (N_22840,N_21819,N_22210);
nand U22841 (N_22841,N_21809,N_22418);
and U22842 (N_22842,N_22195,N_21853);
and U22843 (N_22843,N_22056,N_21735);
nor U22844 (N_22844,N_22177,N_22252);
nand U22845 (N_22845,N_22551,N_22471);
or U22846 (N_22846,N_22679,N_22487);
nor U22847 (N_22847,N_21733,N_22389);
xnor U22848 (N_22848,N_22114,N_22706);
nand U22849 (N_22849,N_22674,N_22455);
nor U22850 (N_22850,N_22375,N_21714);
nand U22851 (N_22851,N_22479,N_22758);
xor U22852 (N_22852,N_22146,N_21880);
or U22853 (N_22853,N_22176,N_21664);
nor U22854 (N_22854,N_22652,N_21950);
nor U22855 (N_22855,N_21711,N_22660);
nor U22856 (N_22856,N_22445,N_22324);
nor U22857 (N_22857,N_22070,N_22245);
xor U22858 (N_22858,N_22648,N_21967);
xor U22859 (N_22859,N_22702,N_22419);
xor U22860 (N_22860,N_22141,N_21752);
or U22861 (N_22861,N_21635,N_22520);
nor U22862 (N_22862,N_22403,N_22489);
nor U22863 (N_22863,N_22279,N_22430);
nor U22864 (N_22864,N_21988,N_22517);
xor U22865 (N_22865,N_22718,N_22695);
or U22866 (N_22866,N_22476,N_21940);
or U22867 (N_22867,N_22630,N_21695);
or U22868 (N_22868,N_22097,N_22456);
nand U22869 (N_22869,N_22728,N_21899);
or U22870 (N_22870,N_22147,N_21912);
nor U22871 (N_22871,N_22591,N_21933);
nor U22872 (N_22872,N_21643,N_22209);
xor U22873 (N_22873,N_22105,N_21621);
nand U22874 (N_22874,N_22287,N_21806);
nor U22875 (N_22875,N_22474,N_21734);
nand U22876 (N_22876,N_22553,N_21851);
and U22877 (N_22877,N_21615,N_22162);
or U22878 (N_22878,N_21926,N_22200);
and U22879 (N_22879,N_21982,N_22052);
nand U22880 (N_22880,N_22484,N_22396);
nor U22881 (N_22881,N_21675,N_22473);
xnor U22882 (N_22882,N_22116,N_21873);
or U22883 (N_22883,N_22133,N_22095);
and U22884 (N_22884,N_21986,N_22420);
nor U22885 (N_22885,N_22661,N_21740);
xor U22886 (N_22886,N_22023,N_22155);
or U22887 (N_22887,N_22646,N_22331);
xnor U22888 (N_22888,N_22565,N_21741);
xor U22889 (N_22889,N_21887,N_22451);
and U22890 (N_22890,N_21638,N_21766);
xor U22891 (N_22891,N_21647,N_22684);
or U22892 (N_22892,N_21852,N_22325);
and U22893 (N_22893,N_21874,N_21707);
nand U22894 (N_22894,N_22417,N_21833);
and U22895 (N_22895,N_21661,N_22271);
or U22896 (N_22896,N_21995,N_22767);
xor U22897 (N_22897,N_22062,N_22170);
and U22898 (N_22898,N_22622,N_22028);
xor U22899 (N_22899,N_22117,N_21946);
xor U22900 (N_22900,N_22590,N_22296);
and U22901 (N_22901,N_22126,N_21657);
or U22902 (N_22902,N_22686,N_21843);
xnor U22903 (N_22903,N_22672,N_21721);
nand U22904 (N_22904,N_22449,N_22136);
or U22905 (N_22905,N_22383,N_21700);
or U22906 (N_22906,N_21610,N_22464);
and U22907 (N_22907,N_22499,N_22319);
and U22908 (N_22908,N_22715,N_21768);
and U22909 (N_22909,N_21816,N_22472);
or U22910 (N_22910,N_21921,N_22190);
nand U22911 (N_22911,N_22341,N_22397);
nor U22912 (N_22912,N_22756,N_21849);
and U22913 (N_22913,N_22665,N_21709);
or U22914 (N_22914,N_22466,N_22079);
nor U22915 (N_22915,N_21901,N_21925);
nor U22916 (N_22916,N_22589,N_21913);
nand U22917 (N_22917,N_22619,N_22475);
xnor U22918 (N_22918,N_22318,N_21811);
nand U22919 (N_22919,N_22048,N_22168);
or U22920 (N_22920,N_22298,N_21628);
nor U22921 (N_22921,N_22478,N_22386);
and U22922 (N_22922,N_21959,N_22444);
nand U22923 (N_22923,N_22343,N_21885);
or U22924 (N_22924,N_22726,N_22447);
or U22925 (N_22925,N_22259,N_21878);
nand U22926 (N_22926,N_22680,N_22625);
and U22927 (N_22927,N_21841,N_22340);
nand U22928 (N_22928,N_22112,N_22067);
and U22929 (N_22929,N_22215,N_22503);
and U22930 (N_22930,N_22579,N_21723);
xnor U22931 (N_22931,N_22422,N_22171);
or U22932 (N_22932,N_22676,N_22534);
and U22933 (N_22933,N_22443,N_21780);
nand U22934 (N_22934,N_21951,N_22360);
and U22935 (N_22935,N_22003,N_22569);
and U22936 (N_22936,N_21759,N_22778);
xnor U22937 (N_22937,N_22390,N_22388);
nor U22938 (N_22938,N_21751,N_21781);
nand U22939 (N_22939,N_22301,N_22108);
nand U22940 (N_22940,N_21854,N_22394);
nand U22941 (N_22941,N_22083,N_22008);
nand U22942 (N_22942,N_22368,N_22697);
or U22943 (N_22943,N_21892,N_21685);
nand U22944 (N_22944,N_22239,N_22567);
xor U22945 (N_22945,N_21865,N_21651);
or U22946 (N_22946,N_21728,N_22303);
or U22947 (N_22947,N_21800,N_22167);
nor U22948 (N_22948,N_21970,N_22749);
nand U22949 (N_22949,N_22521,N_21928);
nand U22950 (N_22950,N_22039,N_22311);
nand U22951 (N_22951,N_21744,N_22234);
or U22952 (N_22952,N_21739,N_22440);
and U22953 (N_22953,N_22647,N_22086);
or U22954 (N_22954,N_22671,N_21775);
xor U22955 (N_22955,N_21726,N_21883);
nor U22956 (N_22956,N_22799,N_21964);
or U22957 (N_22957,N_22635,N_22599);
xor U22958 (N_22958,N_22542,N_21746);
and U22959 (N_22959,N_22532,N_22187);
nand U22960 (N_22960,N_21701,N_22531);
and U22961 (N_22961,N_22281,N_22562);
or U22962 (N_22962,N_21998,N_22429);
and U22963 (N_22963,N_22641,N_22624);
nand U22964 (N_22964,N_22104,N_21722);
nand U22965 (N_22965,N_22152,N_22119);
nor U22966 (N_22966,N_21801,N_21745);
and U22967 (N_22967,N_22255,N_22380);
or U22968 (N_22968,N_21972,N_22598);
or U22969 (N_22969,N_21924,N_22253);
nand U22970 (N_22970,N_22612,N_22300);
or U22971 (N_22971,N_22208,N_22722);
or U22972 (N_22972,N_22131,N_21905);
xor U22973 (N_22973,N_22144,N_21619);
xnor U22974 (N_22974,N_21965,N_21994);
nor U22975 (N_22975,N_22408,N_22110);
or U22976 (N_22976,N_22407,N_22063);
nand U22977 (N_22977,N_22065,N_22607);
and U22978 (N_22978,N_22258,N_21996);
or U22979 (N_22979,N_21835,N_22580);
nand U22980 (N_22980,N_22123,N_22485);
xor U22981 (N_22981,N_22091,N_22362);
xor U22982 (N_22982,N_22416,N_22782);
and U22983 (N_22983,N_21969,N_22154);
xor U22984 (N_22984,N_22164,N_22348);
and U22985 (N_22985,N_21891,N_22613);
xnor U22986 (N_22986,N_21720,N_21724);
nand U22987 (N_22987,N_22696,N_22727);
nor U22988 (N_22988,N_22582,N_22502);
xor U22989 (N_22989,N_21787,N_22349);
and U22990 (N_22990,N_22125,N_21927);
nand U22991 (N_22991,N_21798,N_22611);
xor U22992 (N_22992,N_21945,N_22304);
xnor U22993 (N_22993,N_22768,N_22224);
xor U22994 (N_22994,N_22431,N_22685);
or U22995 (N_22995,N_22351,N_22571);
nor U22996 (N_22996,N_22649,N_22267);
or U22997 (N_22997,N_22214,N_22524);
nand U22998 (N_22998,N_22101,N_21672);
and U22999 (N_22999,N_22497,N_21605);
or U23000 (N_23000,N_22174,N_22547);
xnor U23001 (N_23001,N_21850,N_22035);
nor U23002 (N_23002,N_21903,N_21861);
xor U23003 (N_23003,N_22716,N_22519);
or U23004 (N_23004,N_21642,N_22027);
or U23005 (N_23005,N_22313,N_22439);
nor U23006 (N_23006,N_22406,N_21976);
nor U23007 (N_23007,N_22772,N_22031);
nand U23008 (N_23008,N_22527,N_21606);
nor U23009 (N_23009,N_22160,N_22161);
or U23010 (N_23010,N_21698,N_21881);
nand U23011 (N_23011,N_22068,N_21949);
nor U23012 (N_23012,N_22277,N_22398);
nor U23013 (N_23013,N_21688,N_22078);
or U23014 (N_23014,N_22636,N_21977);
xnor U23015 (N_23015,N_22448,N_22436);
or U23016 (N_23016,N_22384,N_21670);
and U23017 (N_23017,N_22617,N_22558);
or U23018 (N_23018,N_22405,N_21987);
xnor U23019 (N_23019,N_21769,N_21825);
nand U23020 (N_23020,N_22034,N_22217);
xnor U23021 (N_23021,N_22335,N_21753);
xor U23022 (N_23022,N_22196,N_22230);
xor U23023 (N_23023,N_21920,N_22620);
and U23024 (N_23024,N_22453,N_21663);
nor U23025 (N_23025,N_21985,N_21867);
and U23026 (N_23026,N_21684,N_22481);
and U23027 (N_23027,N_22106,N_22583);
nor U23028 (N_23028,N_22411,N_21777);
or U23029 (N_23029,N_22206,N_21730);
and U23030 (N_23030,N_22738,N_22568);
xnor U23031 (N_23031,N_22514,N_21627);
or U23032 (N_23032,N_22033,N_21639);
nor U23033 (N_23033,N_22426,N_21620);
and U23034 (N_23034,N_22747,N_22712);
and U23035 (N_23035,N_22199,N_22310);
nand U23036 (N_23036,N_22080,N_21633);
and U23037 (N_23037,N_22461,N_22670);
nor U23038 (N_23038,N_22786,N_22272);
nand U23039 (N_23039,N_22072,N_22743);
nand U23040 (N_23040,N_21980,N_21983);
xor U23041 (N_23041,N_22606,N_21832);
and U23042 (N_23042,N_22379,N_22038);
xor U23043 (N_23043,N_22566,N_21857);
nor U23044 (N_23044,N_22793,N_22314);
and U23045 (N_23045,N_21629,N_22576);
nor U23046 (N_23046,N_22563,N_22020);
nor U23047 (N_23047,N_21750,N_22731);
xnor U23048 (N_23048,N_22191,N_22669);
nand U23049 (N_23049,N_21778,N_22007);
or U23050 (N_23050,N_21908,N_22525);
xor U23051 (N_23051,N_22069,N_22207);
or U23052 (N_23052,N_22243,N_21919);
nor U23053 (N_23053,N_22593,N_21824);
and U23054 (N_23054,N_22012,N_21821);
nor U23055 (N_23055,N_22051,N_22688);
nand U23056 (N_23056,N_22777,N_21757);
or U23057 (N_23057,N_22244,N_22694);
xor U23058 (N_23058,N_21703,N_21660);
nand U23059 (N_23059,N_22043,N_22729);
nand U23060 (N_23060,N_22184,N_22468);
xnor U23061 (N_23061,N_22204,N_22387);
nand U23062 (N_23062,N_21725,N_22796);
and U23063 (N_23063,N_21958,N_22357);
or U23064 (N_23064,N_22150,N_22507);
nand U23065 (N_23065,N_22554,N_22315);
nand U23066 (N_23066,N_21888,N_21943);
or U23067 (N_23067,N_22730,N_22528);
or U23068 (N_23068,N_22278,N_22100);
xor U23069 (N_23069,N_22347,N_21716);
nor U23070 (N_23070,N_22373,N_22640);
or U23071 (N_23071,N_22410,N_22604);
or U23072 (N_23072,N_21962,N_22442);
nor U23073 (N_23073,N_22365,N_22748);
or U23074 (N_23074,N_22011,N_21762);
nand U23075 (N_23075,N_21763,N_22266);
nand U23076 (N_23076,N_22783,N_21929);
and U23077 (N_23077,N_22306,N_22690);
and U23078 (N_23078,N_22494,N_21957);
xor U23079 (N_23079,N_21779,N_22668);
xnor U23080 (N_23080,N_22570,N_22228);
xor U23081 (N_23081,N_22700,N_22536);
nor U23082 (N_23082,N_22057,N_22797);
xnor U23083 (N_23083,N_22202,N_21845);
nor U23084 (N_23084,N_22401,N_22483);
nand U23085 (N_23085,N_22698,N_21782);
or U23086 (N_23086,N_22560,N_22014);
and U23087 (N_23087,N_22491,N_22276);
nand U23088 (N_23088,N_21646,N_22211);
xnor U23089 (N_23089,N_21917,N_21948);
xor U23090 (N_23090,N_22346,N_22791);
xor U23091 (N_23091,N_22610,N_22124);
nor U23092 (N_23092,N_21742,N_22022);
nand U23093 (N_23093,N_21715,N_22248);
nand U23094 (N_23094,N_21930,N_22629);
xnor U23095 (N_23095,N_21963,N_22032);
and U23096 (N_23096,N_22467,N_22400);
nor U23097 (N_23097,N_22412,N_21823);
nor U23098 (N_23098,N_22182,N_21894);
nand U23099 (N_23099,N_22653,N_22490);
and U23100 (N_23100,N_22754,N_22264);
xor U23101 (N_23101,N_22458,N_22724);
and U23102 (N_23102,N_22366,N_21805);
nor U23103 (N_23103,N_22042,N_22792);
nand U23104 (N_23104,N_21952,N_21810);
nor U23105 (N_23105,N_22076,N_22145);
xor U23106 (N_23106,N_22261,N_22530);
or U23107 (N_23107,N_22575,N_22220);
nor U23108 (N_23108,N_22691,N_22081);
nor U23109 (N_23109,N_22552,N_22293);
nand U23110 (N_23110,N_22678,N_21942);
or U23111 (N_23111,N_22621,N_22659);
nor U23112 (N_23112,N_22251,N_21838);
xnor U23113 (N_23113,N_22452,N_21704);
nand U23114 (N_23114,N_21679,N_22236);
xor U23115 (N_23115,N_22482,N_21937);
and U23116 (N_23116,N_22163,N_21612);
and U23117 (N_23117,N_22172,N_22626);
or U23118 (N_23118,N_22585,N_22723);
and U23119 (N_23119,N_22047,N_22055);
nor U23120 (N_23120,N_22638,N_22559);
xnor U23121 (N_23121,N_22795,N_21828);
and U23122 (N_23122,N_22075,N_21767);
nor U23123 (N_23123,N_21626,N_22283);
xor U23124 (N_23124,N_22798,N_21960);
nand U23125 (N_23125,N_21689,N_22292);
or U23126 (N_23126,N_22781,N_22486);
xnor U23127 (N_23127,N_22708,N_21956);
or U23128 (N_23128,N_22093,N_22717);
nor U23129 (N_23129,N_22581,N_22687);
nor U23130 (N_23130,N_21636,N_22066);
xor U23131 (N_23131,N_21922,N_22769);
or U23132 (N_23132,N_22516,N_22274);
nor U23133 (N_23133,N_21804,N_22683);
nor U23134 (N_23134,N_21673,N_22615);
nor U23135 (N_23135,N_21681,N_21749);
or U23136 (N_23136,N_22654,N_22302);
xnor U23137 (N_23137,N_22539,N_22165);
and U23138 (N_23138,N_22250,N_22735);
nor U23139 (N_23139,N_22509,N_21797);
nand U23140 (N_23140,N_22227,N_22385);
and U23141 (N_23141,N_21856,N_22006);
or U23142 (N_23142,N_22149,N_22492);
nand U23143 (N_23143,N_22699,N_21993);
xnor U23144 (N_23144,N_21844,N_21784);
xor U23145 (N_23145,N_22510,N_22773);
nand U23146 (N_23146,N_21882,N_21614);
and U23147 (N_23147,N_22233,N_22438);
nor U23148 (N_23148,N_22317,N_21788);
xnor U23149 (N_23149,N_21790,N_21674);
nor U23150 (N_23150,N_22381,N_22218);
and U23151 (N_23151,N_22435,N_22454);
or U23152 (N_23152,N_22413,N_22064);
xor U23153 (N_23153,N_21897,N_22098);
nor U23154 (N_23154,N_22290,N_22720);
and U23155 (N_23155,N_22739,N_22437);
and U23156 (N_23156,N_22732,N_22523);
nand U23157 (N_23157,N_21941,N_22040);
xor U23158 (N_23158,N_21813,N_22424);
xor U23159 (N_23159,N_21786,N_22143);
nand U23160 (N_23160,N_22601,N_21872);
xor U23161 (N_23161,N_21984,N_22774);
and U23162 (N_23162,N_21687,N_21654);
xnor U23163 (N_23163,N_22645,N_22297);
xor U23164 (N_23164,N_22273,N_21756);
xor U23165 (N_23165,N_22737,N_21755);
or U23166 (N_23166,N_21641,N_22657);
nor U23167 (N_23167,N_21616,N_22094);
and U23168 (N_23168,N_22460,N_22734);
nor U23169 (N_23169,N_22586,N_21791);
xnor U23170 (N_23170,N_22181,N_22212);
or U23171 (N_23171,N_22755,N_22321);
nor U23172 (N_23172,N_21659,N_22725);
nand U23173 (N_23173,N_22741,N_22102);
nand U23174 (N_23174,N_21658,N_22535);
xnor U23175 (N_23175,N_21822,N_22205);
nand U23176 (N_23176,N_22506,N_22584);
xnor U23177 (N_23177,N_22794,N_22339);
or U23178 (N_23178,N_21708,N_21678);
xor U23179 (N_23179,N_22021,N_21789);
xnor U23180 (N_23180,N_22639,N_21997);
xnor U23181 (N_23181,N_22254,N_22139);
nor U23182 (N_23182,N_21608,N_22462);
nand U23183 (N_23183,N_21692,N_21911);
nand U23184 (N_23184,N_21603,N_21771);
nor U23185 (N_23185,N_21655,N_22705);
nor U23186 (N_23186,N_21802,N_22395);
nand U23187 (N_23187,N_21827,N_21895);
nand U23188 (N_23188,N_21820,N_21826);
nand U23189 (N_23189,N_22330,N_22644);
xnor U23190 (N_23190,N_22628,N_22546);
or U23191 (N_23191,N_22323,N_22173);
nand U23192 (N_23192,N_22223,N_21694);
xnor U23193 (N_23193,N_22704,N_21859);
or U23194 (N_23194,N_22578,N_22221);
and U23195 (N_23195,N_22280,N_22017);
nand U23196 (N_23196,N_22498,N_22096);
xor U23197 (N_23197,N_21935,N_21760);
nand U23198 (N_23198,N_22024,N_22631);
nand U23199 (N_23199,N_22766,N_22049);
nor U23200 (N_23200,N_21989,N_22600);
and U23201 (N_23201,N_22511,N_21600);
and U23202 (N_23202,N_22544,N_22241);
nor U23203 (N_23203,N_21623,N_22441);
and U23204 (N_23204,N_22421,N_21632);
and U23205 (N_23205,N_22409,N_22496);
or U23206 (N_23206,N_22305,N_21936);
nor U23207 (N_23207,N_21737,N_22480);
xnor U23208 (N_23208,N_22713,N_22556);
and U23209 (N_23209,N_21990,N_22216);
or U23210 (N_23210,N_22785,N_22015);
nand U23211 (N_23211,N_22573,N_22651);
xnor U23212 (N_23212,N_21918,N_22001);
or U23213 (N_23213,N_22118,N_22675);
xor U23214 (N_23214,N_21712,N_22789);
and U23215 (N_23215,N_21869,N_21630);
xor U23216 (N_23216,N_22058,N_22434);
or U23217 (N_23217,N_22135,N_22477);
xor U23218 (N_23218,N_22295,N_21855);
or U23219 (N_23219,N_22089,N_21815);
nor U23220 (N_23220,N_21738,N_22092);
nand U23221 (N_23221,N_22120,N_22616);
xnor U23222 (N_23222,N_22329,N_22495);
nand U23223 (N_23223,N_22512,N_21814);
nor U23224 (N_23224,N_22763,N_22128);
xor U23225 (N_23225,N_22692,N_22656);
nor U23226 (N_23226,N_21971,N_21662);
xnor U23227 (N_23227,N_22423,N_22355);
nor U23228 (N_23228,N_21717,N_21904);
nor U23229 (N_23229,N_21764,N_21611);
and U23230 (N_23230,N_22750,N_22746);
and U23231 (N_23231,N_22225,N_22784);
nand U23232 (N_23232,N_21868,N_22603);
or U23233 (N_23233,N_21776,N_22529);
nor U23234 (N_23234,N_22005,N_21732);
nor U23235 (N_23235,N_22356,N_21975);
nand U23236 (N_23236,N_22336,N_22213);
or U23237 (N_23237,N_22197,N_22268);
or U23238 (N_23238,N_21796,N_22088);
nand U23239 (N_23239,N_22677,N_21898);
xnor U23240 (N_23240,N_21667,N_22522);
nor U23241 (N_23241,N_22770,N_22658);
nand U23242 (N_23242,N_22309,N_22371);
nor U23243 (N_23243,N_21893,N_22353);
nor U23244 (N_23244,N_22060,N_22642);
nor U23245 (N_23245,N_22391,N_21602);
nand U23246 (N_23246,N_22745,N_22369);
nor U23247 (N_23247,N_21829,N_22780);
and U23248 (N_23248,N_21840,N_22333);
or U23249 (N_23249,N_22134,N_21713);
and U23250 (N_23250,N_21680,N_22352);
xor U23251 (N_23251,N_21974,N_22122);
nor U23252 (N_23252,N_21624,N_22061);
xnor U23253 (N_23253,N_21938,N_22109);
nand U23254 (N_23254,N_22776,N_22312);
nand U23255 (N_23255,N_22469,N_21864);
and U23256 (N_23256,N_22130,N_21871);
xnor U23257 (N_23257,N_21656,N_21645);
nor U23258 (N_23258,N_22446,N_22374);
nor U23259 (N_23259,N_21808,N_22327);
nand U23260 (N_23260,N_21622,N_22085);
or U23261 (N_23261,N_21705,N_22178);
xor U23262 (N_23262,N_21683,N_22291);
xnor U23263 (N_23263,N_22608,N_21613);
and U23264 (N_23264,N_22082,N_22711);
or U23265 (N_23265,N_22650,N_22740);
and U23266 (N_23266,N_21848,N_22328);
nand U23267 (N_23267,N_22229,N_22761);
and U23268 (N_23268,N_22526,N_22148);
nand U23269 (N_23269,N_21916,N_22378);
xnor U23270 (N_23270,N_22354,N_22256);
xnor U23271 (N_23271,N_21890,N_22275);
nor U23272 (N_23272,N_22294,N_22370);
nand U23273 (N_23273,N_22103,N_22594);
or U23274 (N_23274,N_22463,N_21774);
and U23275 (N_23275,N_22508,N_22790);
or U23276 (N_23276,N_21665,N_21729);
and U23277 (N_23277,N_22030,N_21830);
or U23278 (N_23278,N_22543,N_22693);
nor U23279 (N_23279,N_21773,N_22107);
or U23280 (N_23280,N_22019,N_21915);
nor U23281 (N_23281,N_21617,N_22000);
xor U23282 (N_23282,N_21649,N_22753);
nand U23283 (N_23283,N_21637,N_22036);
and U23284 (N_23284,N_22719,N_21803);
xor U23285 (N_23285,N_22518,N_21601);
nor U23286 (N_23286,N_22285,N_22703);
and U23287 (N_23287,N_22156,N_22779);
xnor U23288 (N_23288,N_21910,N_22159);
or U23289 (N_23289,N_22359,N_22286);
or U23290 (N_23290,N_22151,N_22744);
xnor U23291 (N_23291,N_22428,N_22533);
xor U23292 (N_23292,N_21794,N_21793);
and U23293 (N_23293,N_21807,N_22759);
xor U23294 (N_23294,N_22029,N_21923);
and U23295 (N_23295,N_21668,N_21718);
nand U23296 (N_23296,N_22129,N_22084);
nand U23297 (N_23297,N_22721,N_21650);
nand U23298 (N_23298,N_22041,N_22376);
nand U23299 (N_23299,N_22307,N_22537);
and U23300 (N_23300,N_22180,N_22050);
and U23301 (N_23301,N_21693,N_22788);
and U23302 (N_23302,N_22538,N_22643);
or U23303 (N_23303,N_22002,N_21863);
nor U23304 (N_23304,N_22505,N_22338);
and U23305 (N_23305,N_21889,N_22284);
xor U23306 (N_23306,N_22775,N_22004);
xnor U23307 (N_23307,N_21870,N_21761);
and U23308 (N_23308,N_22113,N_21992);
nor U23309 (N_23309,N_22602,N_21834);
or U23310 (N_23310,N_22588,N_22054);
nand U23311 (N_23311,N_22137,N_22632);
and U23312 (N_23312,N_22242,N_22470);
and U23313 (N_23313,N_22762,N_21991);
nand U23314 (N_23314,N_22249,N_22166);
nor U23315 (N_23315,N_22226,N_21866);
and U23316 (N_23316,N_21783,N_22555);
xor U23317 (N_23317,N_22059,N_22709);
nand U23318 (N_23318,N_21671,N_22247);
nand U23319 (N_23319,N_22771,N_22627);
and U23320 (N_23320,N_22415,N_21884);
nand U23321 (N_23321,N_22053,N_22132);
and U23322 (N_23322,N_22246,N_22540);
nor U23323 (N_23323,N_21652,N_21690);
xor U23324 (N_23324,N_22115,N_21686);
nor U23325 (N_23325,N_22432,N_22367);
or U23326 (N_23326,N_22179,N_22757);
xor U23327 (N_23327,N_21747,N_22714);
and U23328 (N_23328,N_22742,N_22493);
nand U23329 (N_23329,N_22157,N_21696);
nand U23330 (N_23330,N_22402,N_21839);
xnor U23331 (N_23331,N_21677,N_22682);
nor U23332 (N_23332,N_22087,N_22736);
xnor U23333 (N_23333,N_22198,N_22138);
or U23334 (N_23334,N_21981,N_22673);
or U23335 (N_23335,N_22269,N_22504);
or U23336 (N_23336,N_21799,N_22363);
and U23337 (N_23337,N_21931,N_21666);
or U23338 (N_23338,N_22633,N_22414);
nand U23339 (N_23339,N_21876,N_22345);
and U23340 (N_23340,N_22188,N_22597);
or U23341 (N_23341,N_22010,N_22427);
and U23342 (N_23342,N_22623,N_22045);
and U23343 (N_23343,N_22450,N_22681);
nor U23344 (N_23344,N_21858,N_22425);
xnor U23345 (N_23345,N_22459,N_22513);
or U23346 (N_23346,N_22018,N_22142);
or U23347 (N_23347,N_21875,N_22009);
or U23348 (N_23348,N_22337,N_22222);
xor U23349 (N_23349,N_21944,N_22592);
and U23350 (N_23350,N_21900,N_22372);
xor U23351 (N_23351,N_21979,N_22614);
and U23352 (N_23352,N_22664,N_22334);
or U23353 (N_23353,N_21973,N_21653);
nor U23354 (N_23354,N_22016,N_22595);
and U23355 (N_23355,N_22764,N_22733);
and U23356 (N_23356,N_22501,N_21719);
or U23357 (N_23357,N_21785,N_22026);
nand U23358 (N_23358,N_22099,N_22662);
xnor U23359 (N_23359,N_21604,N_22073);
and U23360 (N_23360,N_21862,N_22044);
nor U23361 (N_23361,N_22262,N_21754);
xor U23362 (N_23362,N_22299,N_22787);
nand U23363 (N_23363,N_21846,N_22377);
or U23364 (N_23364,N_21748,N_22342);
nand U23365 (N_23365,N_22185,N_22689);
nand U23366 (N_23366,N_21727,N_22127);
nor U23367 (N_23367,N_21837,N_22158);
or U23368 (N_23368,N_22270,N_22667);
nand U23369 (N_23369,N_21699,N_22488);
nor U23370 (N_23370,N_21914,N_21772);
nor U23371 (N_23371,N_22289,N_22238);
nor U23372 (N_23372,N_21644,N_21978);
and U23373 (N_23373,N_22392,N_21932);
nor U23374 (N_23374,N_22192,N_22046);
nand U23375 (N_23375,N_21847,N_22265);
xnor U23376 (N_23376,N_21966,N_22515);
and U23377 (N_23377,N_22263,N_21691);
nor U23378 (N_23378,N_22203,N_22561);
or U23379 (N_23379,N_21731,N_22121);
nor U23380 (N_23380,N_22037,N_21955);
and U23381 (N_23381,N_22666,N_22752);
or U23382 (N_23382,N_21939,N_21818);
nor U23383 (N_23383,N_22596,N_21631);
and U23384 (N_23384,N_22574,N_22232);
xor U23385 (N_23385,N_21706,N_22545);
and U23386 (N_23386,N_22025,N_21968);
nor U23387 (N_23387,N_22288,N_22557);
and U23388 (N_23388,N_21906,N_22707);
nand U23389 (N_23389,N_22316,N_22572);
nor U23390 (N_23390,N_21817,N_21909);
nand U23391 (N_23391,N_22549,N_21758);
nor U23392 (N_23392,N_21609,N_21792);
or U23393 (N_23393,N_22457,N_21697);
xnor U23394 (N_23394,N_22605,N_21934);
xor U23395 (N_23395,N_22564,N_22548);
or U23396 (N_23396,N_21947,N_21836);
or U23397 (N_23397,N_22193,N_21954);
xor U23398 (N_23398,N_22183,N_21640);
nor U23399 (N_23399,N_22550,N_22326);
and U23400 (N_23400,N_22708,N_21918);
or U23401 (N_23401,N_22278,N_21835);
nor U23402 (N_23402,N_21991,N_21642);
or U23403 (N_23403,N_22461,N_22158);
xor U23404 (N_23404,N_22799,N_22742);
nor U23405 (N_23405,N_21754,N_22727);
xor U23406 (N_23406,N_21931,N_21974);
nand U23407 (N_23407,N_21959,N_22085);
nand U23408 (N_23408,N_22586,N_22227);
nand U23409 (N_23409,N_21799,N_22771);
xnor U23410 (N_23410,N_21837,N_21945);
nand U23411 (N_23411,N_22509,N_21647);
nand U23412 (N_23412,N_22338,N_21715);
or U23413 (N_23413,N_22663,N_22460);
xor U23414 (N_23414,N_21789,N_22524);
nand U23415 (N_23415,N_22056,N_22198);
and U23416 (N_23416,N_21888,N_21926);
nor U23417 (N_23417,N_21875,N_22737);
and U23418 (N_23418,N_22578,N_22512);
or U23419 (N_23419,N_22298,N_22647);
and U23420 (N_23420,N_22729,N_22124);
nor U23421 (N_23421,N_21803,N_21608);
nand U23422 (N_23422,N_21642,N_22340);
and U23423 (N_23423,N_22167,N_22484);
xor U23424 (N_23424,N_22652,N_22464);
nand U23425 (N_23425,N_22079,N_22178);
nor U23426 (N_23426,N_22560,N_21618);
and U23427 (N_23427,N_22164,N_22628);
nor U23428 (N_23428,N_21643,N_21899);
xor U23429 (N_23429,N_22406,N_22546);
nand U23430 (N_23430,N_22309,N_22531);
and U23431 (N_23431,N_22749,N_22305);
nand U23432 (N_23432,N_22663,N_22473);
nand U23433 (N_23433,N_22197,N_22063);
and U23434 (N_23434,N_21872,N_21882);
and U23435 (N_23435,N_21963,N_22055);
or U23436 (N_23436,N_22460,N_22777);
xor U23437 (N_23437,N_22209,N_22275);
or U23438 (N_23438,N_21704,N_21932);
nor U23439 (N_23439,N_22069,N_22333);
or U23440 (N_23440,N_21781,N_21951);
xnor U23441 (N_23441,N_22293,N_21783);
or U23442 (N_23442,N_21783,N_22574);
and U23443 (N_23443,N_22199,N_21801);
nand U23444 (N_23444,N_22582,N_22330);
nor U23445 (N_23445,N_21615,N_21917);
nor U23446 (N_23446,N_22016,N_21725);
or U23447 (N_23447,N_22520,N_21860);
nand U23448 (N_23448,N_22017,N_21955);
xor U23449 (N_23449,N_22760,N_22430);
xnor U23450 (N_23450,N_21818,N_22073);
xnor U23451 (N_23451,N_22241,N_22785);
xor U23452 (N_23452,N_22086,N_22103);
nand U23453 (N_23453,N_22128,N_21984);
or U23454 (N_23454,N_21845,N_21680);
xor U23455 (N_23455,N_22062,N_22784);
or U23456 (N_23456,N_22157,N_21961);
nand U23457 (N_23457,N_22162,N_22308);
xnor U23458 (N_23458,N_21822,N_22327);
and U23459 (N_23459,N_22781,N_21861);
nor U23460 (N_23460,N_21754,N_21915);
xor U23461 (N_23461,N_21681,N_22609);
xor U23462 (N_23462,N_22558,N_22040);
xor U23463 (N_23463,N_22682,N_22557);
or U23464 (N_23464,N_21951,N_21820);
or U23465 (N_23465,N_21793,N_22493);
nor U23466 (N_23466,N_21909,N_22123);
xnor U23467 (N_23467,N_21960,N_22139);
nor U23468 (N_23468,N_21845,N_22719);
or U23469 (N_23469,N_21912,N_22279);
xnor U23470 (N_23470,N_22770,N_22478);
or U23471 (N_23471,N_22440,N_21863);
nor U23472 (N_23472,N_22012,N_22024);
and U23473 (N_23473,N_22549,N_22603);
or U23474 (N_23474,N_21613,N_22794);
xor U23475 (N_23475,N_21772,N_22773);
nand U23476 (N_23476,N_21695,N_22746);
or U23477 (N_23477,N_21788,N_21648);
or U23478 (N_23478,N_21992,N_22392);
nand U23479 (N_23479,N_21613,N_22380);
nand U23480 (N_23480,N_22292,N_21935);
nor U23481 (N_23481,N_22158,N_22495);
nand U23482 (N_23482,N_22354,N_22108);
nand U23483 (N_23483,N_21836,N_22581);
xor U23484 (N_23484,N_22788,N_22572);
nor U23485 (N_23485,N_22031,N_22367);
xor U23486 (N_23486,N_21956,N_22254);
and U23487 (N_23487,N_22718,N_22350);
and U23488 (N_23488,N_22691,N_22153);
nor U23489 (N_23489,N_22409,N_21749);
and U23490 (N_23490,N_21631,N_21851);
or U23491 (N_23491,N_22302,N_22601);
nor U23492 (N_23492,N_22628,N_22595);
and U23493 (N_23493,N_22150,N_22463);
or U23494 (N_23494,N_21808,N_21782);
nor U23495 (N_23495,N_21701,N_22189);
xnor U23496 (N_23496,N_22751,N_22643);
and U23497 (N_23497,N_22322,N_21874);
or U23498 (N_23498,N_22049,N_22567);
xor U23499 (N_23499,N_22472,N_21628);
nand U23500 (N_23500,N_22222,N_21980);
or U23501 (N_23501,N_22497,N_22268);
nor U23502 (N_23502,N_21750,N_21978);
and U23503 (N_23503,N_22686,N_21885);
or U23504 (N_23504,N_21696,N_21684);
xnor U23505 (N_23505,N_22042,N_22641);
nor U23506 (N_23506,N_21633,N_22293);
nand U23507 (N_23507,N_22407,N_22501);
or U23508 (N_23508,N_21885,N_22757);
xor U23509 (N_23509,N_21916,N_21889);
nand U23510 (N_23510,N_22196,N_21628);
or U23511 (N_23511,N_22095,N_22461);
and U23512 (N_23512,N_22544,N_21952);
nor U23513 (N_23513,N_22242,N_21795);
xor U23514 (N_23514,N_22179,N_21901);
and U23515 (N_23515,N_22699,N_22167);
or U23516 (N_23516,N_21751,N_21965);
and U23517 (N_23517,N_21730,N_22104);
or U23518 (N_23518,N_21850,N_22595);
or U23519 (N_23519,N_22503,N_21845);
nor U23520 (N_23520,N_22106,N_22565);
nor U23521 (N_23521,N_21779,N_22026);
nand U23522 (N_23522,N_22324,N_22009);
xnor U23523 (N_23523,N_21968,N_22144);
nand U23524 (N_23524,N_22781,N_21828);
or U23525 (N_23525,N_22212,N_22360);
xor U23526 (N_23526,N_22518,N_21667);
nor U23527 (N_23527,N_22154,N_21670);
xor U23528 (N_23528,N_22756,N_22111);
nor U23529 (N_23529,N_21977,N_22422);
or U23530 (N_23530,N_21815,N_21647);
nand U23531 (N_23531,N_21852,N_21810);
nor U23532 (N_23532,N_21967,N_22376);
or U23533 (N_23533,N_22723,N_22575);
nand U23534 (N_23534,N_22029,N_21690);
nand U23535 (N_23535,N_21973,N_22743);
nand U23536 (N_23536,N_22078,N_22736);
or U23537 (N_23537,N_22553,N_21683);
nor U23538 (N_23538,N_22775,N_21666);
nor U23539 (N_23539,N_21911,N_22262);
nor U23540 (N_23540,N_21603,N_22743);
or U23541 (N_23541,N_21718,N_22317);
and U23542 (N_23542,N_21881,N_22326);
and U23543 (N_23543,N_21697,N_21703);
nor U23544 (N_23544,N_22390,N_22334);
and U23545 (N_23545,N_21791,N_22492);
nand U23546 (N_23546,N_22664,N_22772);
nor U23547 (N_23547,N_22752,N_22632);
nand U23548 (N_23548,N_22206,N_22218);
xor U23549 (N_23549,N_22665,N_22558);
and U23550 (N_23550,N_21606,N_22275);
nor U23551 (N_23551,N_22566,N_22485);
nand U23552 (N_23552,N_22538,N_22212);
or U23553 (N_23553,N_22716,N_22062);
and U23554 (N_23554,N_21669,N_22500);
or U23555 (N_23555,N_22775,N_21865);
nor U23556 (N_23556,N_22503,N_22135);
and U23557 (N_23557,N_22188,N_22118);
or U23558 (N_23558,N_22407,N_21786);
nand U23559 (N_23559,N_22285,N_22328);
xnor U23560 (N_23560,N_21983,N_22759);
xor U23561 (N_23561,N_22497,N_22402);
and U23562 (N_23562,N_22156,N_22386);
and U23563 (N_23563,N_22764,N_22449);
nand U23564 (N_23564,N_21727,N_21904);
nor U23565 (N_23565,N_22780,N_22100);
xor U23566 (N_23566,N_22105,N_21623);
nand U23567 (N_23567,N_22564,N_21774);
nor U23568 (N_23568,N_22611,N_22792);
xnor U23569 (N_23569,N_22315,N_21873);
and U23570 (N_23570,N_22140,N_21652);
or U23571 (N_23571,N_22418,N_22759);
and U23572 (N_23572,N_22338,N_22543);
and U23573 (N_23573,N_21984,N_21665);
nor U23574 (N_23574,N_21742,N_22521);
xor U23575 (N_23575,N_21931,N_21971);
nand U23576 (N_23576,N_22143,N_21684);
xnor U23577 (N_23577,N_22560,N_22410);
or U23578 (N_23578,N_22479,N_22590);
xor U23579 (N_23579,N_21672,N_21966);
or U23580 (N_23580,N_22134,N_21871);
and U23581 (N_23581,N_22558,N_22404);
nand U23582 (N_23582,N_21938,N_21877);
or U23583 (N_23583,N_22118,N_21672);
and U23584 (N_23584,N_21865,N_22283);
nor U23585 (N_23585,N_22359,N_21701);
and U23586 (N_23586,N_22640,N_21732);
and U23587 (N_23587,N_22637,N_22601);
xnor U23588 (N_23588,N_21870,N_22039);
nand U23589 (N_23589,N_22495,N_22211);
xnor U23590 (N_23590,N_22199,N_22076);
nand U23591 (N_23591,N_22186,N_22152);
xnor U23592 (N_23592,N_21965,N_22088);
nand U23593 (N_23593,N_22551,N_22208);
xnor U23594 (N_23594,N_21601,N_22001);
nor U23595 (N_23595,N_21799,N_21621);
nand U23596 (N_23596,N_21736,N_22456);
or U23597 (N_23597,N_21941,N_22791);
nor U23598 (N_23598,N_22459,N_22690);
or U23599 (N_23599,N_21730,N_22173);
nor U23600 (N_23600,N_22334,N_22611);
xor U23601 (N_23601,N_22510,N_22312);
or U23602 (N_23602,N_22382,N_22205);
and U23603 (N_23603,N_21953,N_22795);
xnor U23604 (N_23604,N_22675,N_22678);
or U23605 (N_23605,N_22602,N_22743);
nand U23606 (N_23606,N_21866,N_22247);
xor U23607 (N_23607,N_21860,N_22241);
xnor U23608 (N_23608,N_21924,N_22203);
nand U23609 (N_23609,N_21644,N_21932);
or U23610 (N_23610,N_22021,N_22507);
nand U23611 (N_23611,N_22352,N_22055);
or U23612 (N_23612,N_21982,N_22424);
and U23613 (N_23613,N_22314,N_21894);
nor U23614 (N_23614,N_21631,N_22468);
and U23615 (N_23615,N_22737,N_22066);
nor U23616 (N_23616,N_21688,N_22432);
nand U23617 (N_23617,N_22653,N_22626);
nand U23618 (N_23618,N_22468,N_22101);
nand U23619 (N_23619,N_21794,N_22473);
or U23620 (N_23620,N_22134,N_22060);
nand U23621 (N_23621,N_22077,N_22146);
or U23622 (N_23622,N_22456,N_21649);
and U23623 (N_23623,N_22612,N_22684);
nand U23624 (N_23624,N_22710,N_21655);
or U23625 (N_23625,N_21705,N_22355);
and U23626 (N_23626,N_22601,N_22294);
nand U23627 (N_23627,N_21788,N_22100);
xnor U23628 (N_23628,N_22365,N_22233);
nor U23629 (N_23629,N_21634,N_22529);
nand U23630 (N_23630,N_22237,N_22425);
xnor U23631 (N_23631,N_22255,N_22582);
nor U23632 (N_23632,N_22567,N_21923);
or U23633 (N_23633,N_21922,N_22589);
xnor U23634 (N_23634,N_21813,N_21924);
xnor U23635 (N_23635,N_22144,N_22285);
or U23636 (N_23636,N_22476,N_21971);
or U23637 (N_23637,N_22473,N_21831);
nand U23638 (N_23638,N_22252,N_21948);
or U23639 (N_23639,N_21750,N_22472);
and U23640 (N_23640,N_21663,N_21697);
and U23641 (N_23641,N_22144,N_22578);
xor U23642 (N_23642,N_22545,N_21887);
and U23643 (N_23643,N_21829,N_22528);
and U23644 (N_23644,N_22097,N_22445);
or U23645 (N_23645,N_22785,N_22355);
or U23646 (N_23646,N_22324,N_21741);
or U23647 (N_23647,N_22695,N_22612);
nor U23648 (N_23648,N_21748,N_22316);
nand U23649 (N_23649,N_21745,N_22604);
xnor U23650 (N_23650,N_22364,N_22132);
nor U23651 (N_23651,N_21623,N_22603);
xor U23652 (N_23652,N_22534,N_22388);
or U23653 (N_23653,N_21756,N_22231);
nand U23654 (N_23654,N_22157,N_22044);
or U23655 (N_23655,N_21627,N_21865);
xnor U23656 (N_23656,N_21817,N_22377);
nand U23657 (N_23657,N_22679,N_21844);
nor U23658 (N_23658,N_22288,N_21978);
or U23659 (N_23659,N_21757,N_22724);
and U23660 (N_23660,N_21915,N_22472);
and U23661 (N_23661,N_22154,N_22465);
or U23662 (N_23662,N_22227,N_22567);
nor U23663 (N_23663,N_21827,N_22441);
nand U23664 (N_23664,N_21876,N_22703);
nand U23665 (N_23665,N_21601,N_22643);
or U23666 (N_23666,N_21852,N_22579);
or U23667 (N_23667,N_22599,N_22461);
nor U23668 (N_23668,N_22306,N_22423);
and U23669 (N_23669,N_21602,N_22193);
xor U23670 (N_23670,N_22195,N_21639);
xor U23671 (N_23671,N_21868,N_22200);
nor U23672 (N_23672,N_22030,N_22436);
nand U23673 (N_23673,N_22346,N_22198);
xnor U23674 (N_23674,N_22335,N_22257);
and U23675 (N_23675,N_21696,N_22463);
and U23676 (N_23676,N_22755,N_22406);
xor U23677 (N_23677,N_22055,N_21626);
and U23678 (N_23678,N_22416,N_21804);
and U23679 (N_23679,N_22610,N_22458);
nor U23680 (N_23680,N_21748,N_22725);
and U23681 (N_23681,N_22484,N_21772);
nand U23682 (N_23682,N_22137,N_22357);
nand U23683 (N_23683,N_22700,N_22240);
or U23684 (N_23684,N_22644,N_22713);
and U23685 (N_23685,N_22753,N_21608);
or U23686 (N_23686,N_21615,N_22732);
xnor U23687 (N_23687,N_22339,N_22730);
nor U23688 (N_23688,N_21971,N_22228);
or U23689 (N_23689,N_22201,N_22645);
and U23690 (N_23690,N_21968,N_21652);
nor U23691 (N_23691,N_21797,N_22009);
nand U23692 (N_23692,N_22437,N_22542);
or U23693 (N_23693,N_22549,N_21625);
nand U23694 (N_23694,N_21794,N_22100);
nor U23695 (N_23695,N_22490,N_21635);
xnor U23696 (N_23696,N_21980,N_21992);
nor U23697 (N_23697,N_21959,N_22697);
or U23698 (N_23698,N_22514,N_22377);
or U23699 (N_23699,N_22633,N_22748);
nor U23700 (N_23700,N_22464,N_22169);
nor U23701 (N_23701,N_21629,N_21857);
xnor U23702 (N_23702,N_22165,N_22746);
and U23703 (N_23703,N_21909,N_21940);
or U23704 (N_23704,N_21999,N_22774);
xnor U23705 (N_23705,N_21608,N_22189);
or U23706 (N_23706,N_22368,N_22096);
xor U23707 (N_23707,N_22056,N_22337);
or U23708 (N_23708,N_22206,N_22179);
or U23709 (N_23709,N_22473,N_22177);
or U23710 (N_23710,N_22359,N_22529);
nand U23711 (N_23711,N_22207,N_22301);
or U23712 (N_23712,N_21946,N_22622);
nand U23713 (N_23713,N_22432,N_22238);
xor U23714 (N_23714,N_21910,N_22685);
or U23715 (N_23715,N_22782,N_21655);
or U23716 (N_23716,N_21935,N_22401);
xnor U23717 (N_23717,N_22488,N_22635);
and U23718 (N_23718,N_22047,N_21853);
xnor U23719 (N_23719,N_22508,N_22064);
and U23720 (N_23720,N_22529,N_22545);
nand U23721 (N_23721,N_22223,N_22450);
xnor U23722 (N_23722,N_22551,N_22093);
nand U23723 (N_23723,N_22713,N_21677);
xor U23724 (N_23724,N_22687,N_21673);
xnor U23725 (N_23725,N_22710,N_22555);
nand U23726 (N_23726,N_22009,N_22659);
nand U23727 (N_23727,N_22580,N_22450);
or U23728 (N_23728,N_22155,N_22479);
or U23729 (N_23729,N_22748,N_22142);
nand U23730 (N_23730,N_22268,N_22753);
or U23731 (N_23731,N_22798,N_21951);
nand U23732 (N_23732,N_22656,N_22307);
nand U23733 (N_23733,N_21722,N_22475);
nor U23734 (N_23734,N_21719,N_21945);
or U23735 (N_23735,N_21982,N_22498);
or U23736 (N_23736,N_22708,N_22523);
nor U23737 (N_23737,N_22367,N_21935);
nand U23738 (N_23738,N_21793,N_22684);
nand U23739 (N_23739,N_21900,N_21660);
nand U23740 (N_23740,N_22041,N_21916);
nor U23741 (N_23741,N_22389,N_22077);
nand U23742 (N_23742,N_22156,N_21871);
or U23743 (N_23743,N_22365,N_21609);
and U23744 (N_23744,N_22334,N_22281);
nand U23745 (N_23745,N_21983,N_22019);
nand U23746 (N_23746,N_22745,N_22609);
and U23747 (N_23747,N_21763,N_22730);
or U23748 (N_23748,N_21644,N_22503);
nand U23749 (N_23749,N_22070,N_21943);
nand U23750 (N_23750,N_21813,N_22120);
and U23751 (N_23751,N_22608,N_22525);
nand U23752 (N_23752,N_22709,N_22150);
or U23753 (N_23753,N_22074,N_21615);
xnor U23754 (N_23754,N_21740,N_21854);
nor U23755 (N_23755,N_22542,N_22166);
or U23756 (N_23756,N_22140,N_22427);
or U23757 (N_23757,N_22396,N_22240);
or U23758 (N_23758,N_22324,N_21657);
nand U23759 (N_23759,N_22563,N_22587);
xnor U23760 (N_23760,N_22779,N_21765);
nor U23761 (N_23761,N_21782,N_22488);
or U23762 (N_23762,N_21754,N_22486);
xor U23763 (N_23763,N_22034,N_22317);
xor U23764 (N_23764,N_22743,N_22258);
nor U23765 (N_23765,N_22513,N_22054);
nand U23766 (N_23766,N_21666,N_22405);
nand U23767 (N_23767,N_21712,N_21669);
nand U23768 (N_23768,N_21795,N_22482);
xnor U23769 (N_23769,N_22388,N_22370);
nor U23770 (N_23770,N_21652,N_21913);
or U23771 (N_23771,N_21801,N_21645);
and U23772 (N_23772,N_22661,N_21746);
nor U23773 (N_23773,N_21869,N_22172);
nand U23774 (N_23774,N_22603,N_22180);
xnor U23775 (N_23775,N_21987,N_22507);
nor U23776 (N_23776,N_21656,N_21842);
or U23777 (N_23777,N_22025,N_22555);
and U23778 (N_23778,N_21998,N_22025);
or U23779 (N_23779,N_21621,N_22170);
or U23780 (N_23780,N_21615,N_22443);
nand U23781 (N_23781,N_22703,N_22004);
xor U23782 (N_23782,N_22097,N_21815);
nor U23783 (N_23783,N_22626,N_21614);
or U23784 (N_23784,N_22447,N_22677);
nor U23785 (N_23785,N_22205,N_21899);
and U23786 (N_23786,N_21887,N_22165);
and U23787 (N_23787,N_22011,N_21738);
or U23788 (N_23788,N_21648,N_21844);
xnor U23789 (N_23789,N_21827,N_22336);
xnor U23790 (N_23790,N_22082,N_21961);
nand U23791 (N_23791,N_22680,N_22609);
xnor U23792 (N_23792,N_22128,N_22247);
xor U23793 (N_23793,N_22435,N_22754);
nand U23794 (N_23794,N_21969,N_21773);
xor U23795 (N_23795,N_22653,N_22755);
or U23796 (N_23796,N_21744,N_22402);
nor U23797 (N_23797,N_22325,N_21826);
and U23798 (N_23798,N_22045,N_22021);
or U23799 (N_23799,N_22071,N_21877);
nor U23800 (N_23800,N_21987,N_21902);
nand U23801 (N_23801,N_22063,N_22145);
and U23802 (N_23802,N_22289,N_21989);
or U23803 (N_23803,N_21867,N_22330);
or U23804 (N_23804,N_22248,N_21800);
xor U23805 (N_23805,N_22585,N_22022);
nor U23806 (N_23806,N_22057,N_22734);
nor U23807 (N_23807,N_22771,N_22416);
nor U23808 (N_23808,N_22547,N_22212);
nor U23809 (N_23809,N_21961,N_22340);
nor U23810 (N_23810,N_22751,N_21981);
nand U23811 (N_23811,N_21621,N_21932);
nand U23812 (N_23812,N_22429,N_22603);
and U23813 (N_23813,N_22259,N_22416);
xnor U23814 (N_23814,N_21870,N_21705);
or U23815 (N_23815,N_22145,N_21735);
xnor U23816 (N_23816,N_22663,N_22353);
nor U23817 (N_23817,N_21812,N_21703);
xnor U23818 (N_23818,N_22259,N_21767);
nor U23819 (N_23819,N_21716,N_21801);
nand U23820 (N_23820,N_22523,N_22653);
and U23821 (N_23821,N_22681,N_22095);
nor U23822 (N_23822,N_22735,N_22205);
and U23823 (N_23823,N_21864,N_21893);
nand U23824 (N_23824,N_22621,N_22142);
xor U23825 (N_23825,N_22509,N_21666);
or U23826 (N_23826,N_21720,N_22794);
and U23827 (N_23827,N_22187,N_22242);
and U23828 (N_23828,N_22468,N_21707);
or U23829 (N_23829,N_21824,N_22110);
xnor U23830 (N_23830,N_22007,N_22429);
or U23831 (N_23831,N_21815,N_22168);
and U23832 (N_23832,N_22726,N_22279);
nor U23833 (N_23833,N_21677,N_22360);
nor U23834 (N_23834,N_22622,N_22159);
nor U23835 (N_23835,N_21799,N_22283);
and U23836 (N_23836,N_22660,N_21747);
nor U23837 (N_23837,N_22267,N_21838);
xnor U23838 (N_23838,N_22417,N_22549);
nand U23839 (N_23839,N_22697,N_22490);
nand U23840 (N_23840,N_22202,N_22195);
and U23841 (N_23841,N_22728,N_22716);
or U23842 (N_23842,N_22576,N_22186);
nor U23843 (N_23843,N_22582,N_22275);
xor U23844 (N_23844,N_22707,N_21863);
nor U23845 (N_23845,N_21869,N_21765);
nor U23846 (N_23846,N_22174,N_22644);
xor U23847 (N_23847,N_22746,N_22297);
and U23848 (N_23848,N_22019,N_22364);
or U23849 (N_23849,N_21734,N_22611);
xor U23850 (N_23850,N_22505,N_21816);
or U23851 (N_23851,N_21773,N_22165);
or U23852 (N_23852,N_21690,N_22554);
and U23853 (N_23853,N_21963,N_22715);
nor U23854 (N_23854,N_22421,N_22084);
or U23855 (N_23855,N_22782,N_22138);
nor U23856 (N_23856,N_21975,N_22708);
nand U23857 (N_23857,N_21648,N_22499);
nor U23858 (N_23858,N_21902,N_21956);
nand U23859 (N_23859,N_22633,N_21902);
nand U23860 (N_23860,N_22197,N_22668);
and U23861 (N_23861,N_22203,N_21670);
xor U23862 (N_23862,N_21838,N_21834);
nor U23863 (N_23863,N_22412,N_22190);
and U23864 (N_23864,N_22641,N_21875);
or U23865 (N_23865,N_22283,N_22138);
or U23866 (N_23866,N_22564,N_22466);
nand U23867 (N_23867,N_22673,N_22557);
xnor U23868 (N_23868,N_22280,N_22432);
nand U23869 (N_23869,N_22071,N_22791);
xnor U23870 (N_23870,N_21602,N_22511);
nor U23871 (N_23871,N_22263,N_22627);
nand U23872 (N_23872,N_22437,N_22635);
nor U23873 (N_23873,N_22341,N_22674);
and U23874 (N_23874,N_21884,N_22337);
nand U23875 (N_23875,N_22151,N_22416);
and U23876 (N_23876,N_21750,N_22570);
xor U23877 (N_23877,N_21653,N_21877);
nor U23878 (N_23878,N_22132,N_22697);
and U23879 (N_23879,N_21621,N_21769);
or U23880 (N_23880,N_21764,N_21722);
nand U23881 (N_23881,N_21913,N_22317);
and U23882 (N_23882,N_21943,N_21715);
nor U23883 (N_23883,N_22772,N_22025);
nand U23884 (N_23884,N_22410,N_22102);
xnor U23885 (N_23885,N_22583,N_22484);
or U23886 (N_23886,N_22069,N_22052);
xnor U23887 (N_23887,N_22006,N_22723);
and U23888 (N_23888,N_22655,N_22261);
xor U23889 (N_23889,N_22722,N_21774);
nor U23890 (N_23890,N_22595,N_22677);
or U23891 (N_23891,N_21743,N_22392);
nand U23892 (N_23892,N_22509,N_21929);
xnor U23893 (N_23893,N_22761,N_21865);
nor U23894 (N_23894,N_21809,N_21897);
nor U23895 (N_23895,N_22199,N_22078);
nor U23896 (N_23896,N_21897,N_22120);
or U23897 (N_23897,N_22092,N_22757);
or U23898 (N_23898,N_22795,N_22115);
xnor U23899 (N_23899,N_22629,N_21931);
nor U23900 (N_23900,N_22480,N_22040);
nand U23901 (N_23901,N_22660,N_22258);
and U23902 (N_23902,N_22729,N_22177);
xor U23903 (N_23903,N_22153,N_22342);
and U23904 (N_23904,N_22052,N_22607);
and U23905 (N_23905,N_21898,N_21825);
xor U23906 (N_23906,N_22568,N_22628);
and U23907 (N_23907,N_22352,N_21871);
and U23908 (N_23908,N_22191,N_22405);
nand U23909 (N_23909,N_22604,N_22684);
xor U23910 (N_23910,N_22562,N_22352);
nor U23911 (N_23911,N_22095,N_22781);
xnor U23912 (N_23912,N_21784,N_22619);
xnor U23913 (N_23913,N_22020,N_22713);
nor U23914 (N_23914,N_22081,N_22476);
or U23915 (N_23915,N_22382,N_22321);
or U23916 (N_23916,N_22287,N_21912);
nor U23917 (N_23917,N_22665,N_21991);
nor U23918 (N_23918,N_22552,N_22396);
and U23919 (N_23919,N_22534,N_21729);
nand U23920 (N_23920,N_21781,N_21657);
xor U23921 (N_23921,N_21785,N_21720);
or U23922 (N_23922,N_22502,N_21792);
or U23923 (N_23923,N_21601,N_22417);
xor U23924 (N_23924,N_21891,N_21917);
and U23925 (N_23925,N_21724,N_22525);
xor U23926 (N_23926,N_22697,N_22749);
nor U23927 (N_23927,N_21990,N_22176);
nand U23928 (N_23928,N_22089,N_21654);
nand U23929 (N_23929,N_21634,N_22018);
or U23930 (N_23930,N_22799,N_22365);
nor U23931 (N_23931,N_21683,N_22184);
nand U23932 (N_23932,N_22481,N_22318);
nand U23933 (N_23933,N_22686,N_22797);
nor U23934 (N_23934,N_21706,N_22455);
or U23935 (N_23935,N_21876,N_21802);
xor U23936 (N_23936,N_22337,N_22505);
xnor U23937 (N_23937,N_22135,N_22388);
xor U23938 (N_23938,N_22264,N_21848);
xnor U23939 (N_23939,N_22069,N_22154);
and U23940 (N_23940,N_22623,N_22524);
nor U23941 (N_23941,N_21631,N_21897);
nand U23942 (N_23942,N_22578,N_22297);
and U23943 (N_23943,N_21893,N_22389);
and U23944 (N_23944,N_22211,N_22046);
xor U23945 (N_23945,N_22482,N_21791);
nor U23946 (N_23946,N_21990,N_21834);
and U23947 (N_23947,N_21652,N_21965);
and U23948 (N_23948,N_21702,N_21871);
or U23949 (N_23949,N_21835,N_22129);
nor U23950 (N_23950,N_21957,N_22503);
or U23951 (N_23951,N_22018,N_21961);
and U23952 (N_23952,N_22004,N_22429);
or U23953 (N_23953,N_22595,N_22776);
or U23954 (N_23954,N_22262,N_22746);
nand U23955 (N_23955,N_22167,N_22136);
nor U23956 (N_23956,N_21713,N_22218);
and U23957 (N_23957,N_22052,N_22355);
and U23958 (N_23958,N_22698,N_22380);
nand U23959 (N_23959,N_21766,N_22535);
xor U23960 (N_23960,N_21939,N_22722);
nand U23961 (N_23961,N_22291,N_22461);
or U23962 (N_23962,N_22098,N_21936);
nor U23963 (N_23963,N_22047,N_22617);
and U23964 (N_23964,N_22273,N_22456);
nor U23965 (N_23965,N_22638,N_22599);
nor U23966 (N_23966,N_21693,N_21950);
xnor U23967 (N_23967,N_21638,N_21653);
and U23968 (N_23968,N_21897,N_22137);
nand U23969 (N_23969,N_21682,N_22634);
and U23970 (N_23970,N_21799,N_21964);
xnor U23971 (N_23971,N_22105,N_22640);
and U23972 (N_23972,N_22468,N_22364);
nor U23973 (N_23973,N_22056,N_22263);
xor U23974 (N_23974,N_21784,N_21800);
or U23975 (N_23975,N_21848,N_21966);
and U23976 (N_23976,N_22657,N_22121);
xor U23977 (N_23977,N_22302,N_22295);
or U23978 (N_23978,N_22578,N_22422);
nor U23979 (N_23979,N_22524,N_22391);
xor U23980 (N_23980,N_21993,N_22657);
or U23981 (N_23981,N_21834,N_21772);
xor U23982 (N_23982,N_22326,N_22409);
or U23983 (N_23983,N_22220,N_22379);
and U23984 (N_23984,N_22569,N_22160);
and U23985 (N_23985,N_22644,N_22005);
or U23986 (N_23986,N_22536,N_22330);
and U23987 (N_23987,N_22474,N_21652);
nor U23988 (N_23988,N_22402,N_21862);
nand U23989 (N_23989,N_21814,N_22793);
xnor U23990 (N_23990,N_21608,N_22219);
or U23991 (N_23991,N_22297,N_22494);
xnor U23992 (N_23992,N_21766,N_22670);
nor U23993 (N_23993,N_21698,N_21679);
xor U23994 (N_23994,N_22053,N_22610);
or U23995 (N_23995,N_22771,N_22751);
and U23996 (N_23996,N_22491,N_22311);
xnor U23997 (N_23997,N_21731,N_22238);
nand U23998 (N_23998,N_22607,N_22258);
xor U23999 (N_23999,N_21960,N_22250);
nand U24000 (N_24000,N_23772,N_23552);
xor U24001 (N_24001,N_23469,N_23053);
nand U24002 (N_24002,N_22904,N_23684);
nand U24003 (N_24003,N_23606,N_23457);
or U24004 (N_24004,N_22974,N_23612);
and U24005 (N_24005,N_22906,N_23449);
and U24006 (N_24006,N_23926,N_23556);
nand U24007 (N_24007,N_23463,N_23398);
nand U24008 (N_24008,N_22867,N_23784);
and U24009 (N_24009,N_22905,N_23117);
and U24010 (N_24010,N_23145,N_23204);
xor U24011 (N_24011,N_22954,N_23789);
nor U24012 (N_24012,N_22957,N_22824);
nand U24013 (N_24013,N_22962,N_23685);
or U24014 (N_24014,N_23374,N_23705);
nand U24015 (N_24015,N_23339,N_22861);
and U24016 (N_24016,N_23063,N_23151);
xor U24017 (N_24017,N_23293,N_23477);
or U24018 (N_24018,N_23871,N_23119);
nand U24019 (N_24019,N_22915,N_23758);
and U24020 (N_24020,N_23370,N_22990);
and U24021 (N_24021,N_22951,N_23137);
nand U24022 (N_24022,N_23541,N_23620);
xor U24023 (N_24023,N_23351,N_23386);
nor U24024 (N_24024,N_23898,N_23610);
or U24025 (N_24025,N_23762,N_23257);
and U24026 (N_24026,N_23847,N_23909);
or U24027 (N_24027,N_23795,N_22830);
and U24028 (N_24028,N_22891,N_23336);
or U24029 (N_24029,N_23460,N_23216);
xnor U24030 (N_24030,N_22925,N_23225);
or U24031 (N_24031,N_22923,N_23717);
and U24032 (N_24032,N_23098,N_23450);
and U24033 (N_24033,N_22980,N_23706);
nand U24034 (N_24034,N_23945,N_23852);
nor U24035 (N_24035,N_23008,N_23628);
or U24036 (N_24036,N_23454,N_23694);
and U24037 (N_24037,N_23292,N_23380);
or U24038 (N_24038,N_23962,N_23046);
nor U24039 (N_24039,N_23433,N_22916);
xnor U24040 (N_24040,N_23050,N_23482);
or U24041 (N_24041,N_23496,N_23208);
and U24042 (N_24042,N_23333,N_23172);
or U24043 (N_24043,N_23271,N_23657);
or U24044 (N_24044,N_23600,N_22963);
and U24045 (N_24045,N_23415,N_23550);
nor U24046 (N_24046,N_23207,N_23180);
xor U24047 (N_24047,N_23273,N_23437);
or U24048 (N_24048,N_23199,N_23782);
or U24049 (N_24049,N_23918,N_23313);
xor U24050 (N_24050,N_23362,N_23341);
or U24051 (N_24051,N_23501,N_23507);
or U24052 (N_24052,N_23078,N_23422);
xnor U24053 (N_24053,N_23448,N_23786);
nand U24054 (N_24054,N_22937,N_23956);
nand U24055 (N_24055,N_22931,N_23618);
xnor U24056 (N_24056,N_23889,N_22947);
nand U24057 (N_24057,N_23551,N_23820);
and U24058 (N_24058,N_23827,N_23754);
or U24059 (N_24059,N_23314,N_23730);
or U24060 (N_24060,N_23049,N_23752);
xor U24061 (N_24061,N_23958,N_22908);
or U24062 (N_24062,N_22973,N_22943);
xnor U24063 (N_24063,N_22953,N_23783);
or U24064 (N_24064,N_22983,N_23083);
and U24065 (N_24065,N_23737,N_23921);
or U24066 (N_24066,N_23838,N_22894);
or U24067 (N_24067,N_23619,N_23653);
xnor U24068 (N_24068,N_22875,N_23245);
xnor U24069 (N_24069,N_22878,N_23082);
nand U24070 (N_24070,N_23868,N_23069);
and U24071 (N_24071,N_23572,N_23532);
xor U24072 (N_24072,N_23294,N_23340);
nand U24073 (N_24073,N_23807,N_23246);
or U24074 (N_24074,N_23139,N_22853);
and U24075 (N_24075,N_23322,N_22800);
or U24076 (N_24076,N_23387,N_23933);
nor U24077 (N_24077,N_22805,N_23116);
or U24078 (N_24078,N_23502,N_23219);
nor U24079 (N_24079,N_22920,N_23989);
nor U24080 (N_24080,N_23179,N_23295);
nor U24081 (N_24081,N_23356,N_23240);
xor U24082 (N_24082,N_23022,N_23335);
xor U24083 (N_24083,N_22985,N_23215);
or U24084 (N_24084,N_23875,N_23006);
xnor U24085 (N_24085,N_22809,N_23344);
xor U24086 (N_24086,N_23138,N_23607);
nand U24087 (N_24087,N_23776,N_23263);
xor U24088 (N_24088,N_23638,N_23744);
nor U24089 (N_24089,N_22834,N_23756);
and U24090 (N_24090,N_23920,N_22949);
nor U24091 (N_24091,N_23315,N_23191);
and U24092 (N_24092,N_23557,N_23650);
or U24093 (N_24093,N_23061,N_23753);
xnor U24094 (N_24094,N_23305,N_23318);
or U24095 (N_24095,N_23939,N_22868);
and U24096 (N_24096,N_23074,N_23656);
nor U24097 (N_24097,N_22892,N_23671);
or U24098 (N_24098,N_23603,N_23359);
and U24099 (N_24099,N_23495,N_22967);
nand U24100 (N_24100,N_22929,N_23916);
and U24101 (N_24101,N_23522,N_23384);
or U24102 (N_24102,N_23743,N_22804);
nor U24103 (N_24103,N_22895,N_23520);
nor U24104 (N_24104,N_23382,N_22932);
nor U24105 (N_24105,N_23913,N_23678);
xor U24106 (N_24106,N_23128,N_23809);
or U24107 (N_24107,N_23017,N_23835);
or U24108 (N_24108,N_23160,N_23876);
xor U24109 (N_24109,N_23662,N_23690);
and U24110 (N_24110,N_23521,N_23000);
and U24111 (N_24111,N_23676,N_23045);
xor U24112 (N_24112,N_23964,N_23709);
and U24113 (N_24113,N_23815,N_23692);
nor U24114 (N_24114,N_23134,N_23252);
nand U24115 (N_24115,N_23330,N_23951);
or U24116 (N_24116,N_22958,N_23093);
nand U24117 (N_24117,N_23872,N_23757);
or U24118 (N_24118,N_23161,N_22907);
and U24119 (N_24119,N_23819,N_23724);
nand U24120 (N_24120,N_23105,N_22910);
and U24121 (N_24121,N_22996,N_23817);
or U24122 (N_24122,N_23652,N_23192);
xnor U24123 (N_24123,N_23266,N_23411);
or U24124 (N_24124,N_23791,N_23251);
and U24125 (N_24125,N_23511,N_23900);
nand U24126 (N_24126,N_23961,N_23354);
or U24127 (N_24127,N_23696,N_23106);
nor U24128 (N_24128,N_23531,N_23682);
nor U24129 (N_24129,N_23476,N_23641);
xor U24130 (N_24130,N_23970,N_22811);
xnor U24131 (N_24131,N_23987,N_23693);
nand U24132 (N_24132,N_23584,N_23133);
and U24133 (N_24133,N_23170,N_23033);
nand U24134 (N_24134,N_23400,N_23887);
or U24135 (N_24135,N_23186,N_22909);
or U24136 (N_24136,N_23242,N_22917);
xor U24137 (N_24137,N_23767,N_23862);
nor U24138 (N_24138,N_23475,N_23338);
and U24139 (N_24139,N_23915,N_23129);
or U24140 (N_24140,N_23930,N_23052);
xor U24141 (N_24141,N_23558,N_22955);
nor U24142 (N_24142,N_23484,N_23513);
xnor U24143 (N_24143,N_23158,N_23923);
xor U24144 (N_24144,N_22820,N_23850);
nor U24145 (N_24145,N_23416,N_22897);
nor U24146 (N_24146,N_22825,N_23393);
nand U24147 (N_24147,N_23394,N_22857);
nand U24148 (N_24148,N_23068,N_23543);
nor U24149 (N_24149,N_23472,N_23894);
nor U24150 (N_24150,N_23542,N_23094);
nand U24151 (N_24151,N_23614,N_23159);
or U24152 (N_24152,N_23683,N_23878);
nor U24153 (N_24153,N_22912,N_23927);
xor U24154 (N_24154,N_23218,N_23593);
nand U24155 (N_24155,N_23658,N_23831);
xnor U24156 (N_24156,N_23514,N_23932);
and U24157 (N_24157,N_22961,N_23494);
and U24158 (N_24158,N_23589,N_23903);
nor U24159 (N_24159,N_23715,N_22968);
nor U24160 (N_24160,N_23585,N_23250);
and U24161 (N_24161,N_23588,N_23402);
and U24162 (N_24162,N_22933,N_23804);
or U24163 (N_24163,N_22810,N_23524);
and U24164 (N_24164,N_23763,N_23282);
and U24165 (N_24165,N_23721,N_23761);
xnor U24166 (N_24166,N_23267,N_23210);
and U24167 (N_24167,N_23481,N_22815);
nor U24168 (N_24168,N_23467,N_22976);
and U24169 (N_24169,N_23197,N_23404);
nor U24170 (N_24170,N_23892,N_23781);
or U24171 (N_24171,N_23539,N_22888);
xor U24172 (N_24172,N_23109,N_23283);
nand U24173 (N_24173,N_23397,N_23734);
nand U24174 (N_24174,N_23981,N_23713);
and U24175 (N_24175,N_22884,N_23195);
nor U24176 (N_24176,N_23566,N_23028);
or U24177 (N_24177,N_23190,N_23978);
or U24178 (N_24178,N_22900,N_23857);
nand U24179 (N_24179,N_22992,N_23451);
and U24180 (N_24180,N_23143,N_23741);
xor U24181 (N_24181,N_23243,N_22986);
nor U24182 (N_24182,N_23675,N_23081);
nand U24183 (N_24183,N_23306,N_22975);
nand U24184 (N_24184,N_23358,N_23001);
nor U24185 (N_24185,N_22972,N_23071);
nand U24186 (N_24186,N_23428,N_23256);
or U24187 (N_24187,N_23591,N_23239);
nand U24188 (N_24188,N_22948,N_23908);
xnor U24189 (N_24189,N_23347,N_23931);
xnor U24190 (N_24190,N_22839,N_23258);
nand U24191 (N_24191,N_23381,N_23301);
xor U24192 (N_24192,N_23714,N_23812);
nand U24193 (N_24193,N_23486,N_23136);
or U24194 (N_24194,N_23794,N_23536);
nand U24195 (N_24195,N_23244,N_23132);
nor U24196 (N_24196,N_23984,N_23544);
nor U24197 (N_24197,N_23147,N_23226);
xor U24198 (N_24198,N_23598,N_23740);
or U24199 (N_24199,N_23048,N_23466);
and U24200 (N_24200,N_22879,N_23429);
nand U24201 (N_24201,N_23639,N_23910);
nand U24202 (N_24202,N_23332,N_23439);
nand U24203 (N_24203,N_23773,N_23198);
xnor U24204 (N_24204,N_23655,N_22881);
nand U24205 (N_24205,N_23072,N_23221);
xor U24206 (N_24206,N_23044,N_23785);
or U24207 (N_24207,N_23442,N_23957);
and U24208 (N_24208,N_23473,N_23453);
and U24209 (N_24209,N_23169,N_23560);
xor U24210 (N_24210,N_23506,N_22964);
and U24211 (N_24211,N_23919,N_23943);
nand U24212 (N_24212,N_22993,N_23980);
xnor U24213 (N_24213,N_23667,N_23084);
nor U24214 (N_24214,N_22886,N_23888);
nand U24215 (N_24215,N_23275,N_23329);
and U24216 (N_24216,N_23311,N_23372);
nor U24217 (N_24217,N_23581,N_23162);
xor U24218 (N_24218,N_23038,N_23366);
nor U24219 (N_24219,N_23260,N_23259);
nor U24220 (N_24220,N_23493,N_22944);
nand U24221 (N_24221,N_22952,N_23201);
xnor U24222 (N_24222,N_23241,N_22858);
or U24223 (N_24223,N_23327,N_23942);
and U24224 (N_24224,N_23976,N_23924);
nand U24225 (N_24225,N_23893,N_22965);
nand U24226 (N_24226,N_23371,N_23051);
or U24227 (N_24227,N_22859,N_23262);
nor U24228 (N_24228,N_23669,N_23582);
xnor U24229 (N_24229,N_23991,N_23220);
nand U24230 (N_24230,N_22987,N_23751);
nand U24231 (N_24231,N_23302,N_23624);
xor U24232 (N_24232,N_23548,N_23851);
xor U24233 (N_24233,N_23565,N_23175);
xnor U24234 (N_24234,N_23408,N_22819);
or U24235 (N_24235,N_23019,N_23176);
nand U24236 (N_24236,N_23613,N_23016);
xor U24237 (N_24237,N_22840,N_23883);
and U24238 (N_24238,N_23316,N_23719);
and U24239 (N_24239,N_23879,N_23825);
xnor U24240 (N_24240,N_23077,N_23352);
nand U24241 (N_24241,N_23444,N_23024);
or U24242 (N_24242,N_23023,N_23181);
xnor U24243 (N_24243,N_23007,N_22940);
or U24244 (N_24244,N_23525,N_23659);
xnor U24245 (N_24245,N_23731,N_23914);
and U24246 (N_24246,N_22849,N_23014);
and U24247 (N_24247,N_22818,N_23649);
nor U24248 (N_24248,N_22913,N_23523);
and U24249 (N_24249,N_23011,N_23745);
xnor U24250 (N_24250,N_23085,N_23108);
nor U24251 (N_24251,N_23056,N_23748);
or U24252 (N_24252,N_22919,N_23228);
xnor U24253 (N_24253,N_22882,N_23080);
nor U24254 (N_24254,N_23399,N_22994);
nand U24255 (N_24255,N_23563,N_23829);
nor U24256 (N_24256,N_23934,N_23065);
xnor U24257 (N_24257,N_22981,N_23342);
or U24258 (N_24258,N_23284,N_23645);
and U24259 (N_24259,N_23421,N_22866);
xor U24260 (N_24260,N_23882,N_23157);
nor U24261 (N_24261,N_23774,N_23264);
nand U24262 (N_24262,N_22883,N_23661);
xnor U24263 (N_24263,N_23518,N_23654);
and U24264 (N_24264,N_23261,N_23103);
and U24265 (N_24265,N_23235,N_23845);
xnor U24266 (N_24266,N_23086,N_23559);
and U24267 (N_24267,N_23944,N_23123);
nand U24268 (N_24268,N_23146,N_23974);
and U24269 (N_24269,N_23505,N_23018);
or U24270 (N_24270,N_22869,N_23529);
nor U24271 (N_24271,N_22828,N_23826);
and U24272 (N_24272,N_22971,N_23867);
and U24273 (N_24273,N_23247,N_23487);
and U24274 (N_24274,N_23609,N_23647);
nor U24275 (N_24275,N_23597,N_23034);
nand U24276 (N_24276,N_23971,N_23615);
or U24277 (N_24277,N_23378,N_23632);
nand U24278 (N_24278,N_23113,N_23200);
nand U24279 (N_24279,N_23902,N_23296);
or U24280 (N_24280,N_23955,N_23674);
nor U24281 (N_24281,N_23746,N_23095);
nor U24282 (N_24282,N_23097,N_23073);
xor U24283 (N_24283,N_23854,N_23577);
and U24284 (N_24284,N_23839,N_23012);
xor U24285 (N_24285,N_23604,N_23977);
and U24286 (N_24286,N_23840,N_23602);
nand U24287 (N_24287,N_23142,N_23222);
nand U24288 (N_24288,N_23237,N_23363);
nor U24289 (N_24289,N_23720,N_22803);
or U24290 (N_24290,N_23039,N_23096);
nand U24291 (N_24291,N_23324,N_23594);
and U24292 (N_24292,N_23935,N_23122);
nand U24293 (N_24293,N_22832,N_23206);
or U24294 (N_24294,N_23688,N_23886);
xnor U24295 (N_24295,N_23365,N_23427);
nor U24296 (N_24296,N_23156,N_23979);
and U24297 (N_24297,N_23861,N_23841);
nor U24298 (N_24298,N_23070,N_23837);
xnor U24299 (N_24299,N_23515,N_23834);
xnor U24300 (N_24300,N_23403,N_23568);
nand U24301 (N_24301,N_23855,N_23698);
nand U24302 (N_24302,N_23865,N_23623);
or U24303 (N_24303,N_23707,N_23822);
nor U24304 (N_24304,N_23575,N_23443);
xor U24305 (N_24305,N_23312,N_23631);
nor U24306 (N_24306,N_23742,N_22960);
xnor U24307 (N_24307,N_23278,N_23303);
nand U24308 (N_24308,N_23229,N_23968);
or U24309 (N_24309,N_23127,N_23736);
nand U24310 (N_24310,N_23379,N_23885);
nor U24311 (N_24311,N_22885,N_23853);
or U24312 (N_24312,N_23066,N_23323);
nor U24313 (N_24313,N_23777,N_23574);
xnor U24314 (N_24314,N_23465,N_23643);
xor U24315 (N_24315,N_23104,N_23897);
or U24316 (N_24316,N_22872,N_23986);
or U24317 (N_24317,N_22842,N_23739);
nand U24318 (N_24318,N_23291,N_23995);
nor U24319 (N_24319,N_23504,N_22847);
nand U24320 (N_24320,N_23355,N_23771);
xnor U24321 (N_24321,N_23832,N_23027);
xnor U24322 (N_24322,N_23478,N_23140);
xnor U24323 (N_24323,N_22848,N_23067);
nand U24324 (N_24324,N_23032,N_23925);
nor U24325 (N_24325,N_23184,N_23182);
nor U24326 (N_24326,N_23953,N_23174);
nand U24327 (N_24327,N_23155,N_23899);
xor U24328 (N_24328,N_23360,N_23966);
nor U24329 (N_24329,N_23567,N_23031);
nor U24330 (N_24330,N_23249,N_22833);
or U24331 (N_24331,N_22978,N_23842);
nor U24332 (N_24332,N_23177,N_23877);
nor U24333 (N_24333,N_23859,N_22856);
nand U24334 (N_24334,N_23409,N_23972);
nor U24335 (N_24335,N_23004,N_23759);
nor U24336 (N_24336,N_23747,N_23858);
or U24337 (N_24337,N_23223,N_23490);
nand U24338 (N_24338,N_23418,N_23948);
nor U24339 (N_24339,N_23874,N_23406);
nor U24340 (N_24340,N_23232,N_23230);
or U24341 (N_24341,N_23405,N_23592);
or U24342 (N_24342,N_23111,N_23990);
nor U24343 (N_24343,N_22852,N_23349);
nor U24344 (N_24344,N_23153,N_23664);
nor U24345 (N_24345,N_23555,N_23281);
or U24346 (N_24346,N_23700,N_23485);
nand U24347 (N_24347,N_23905,N_23873);
nor U24348 (N_24348,N_23407,N_22841);
nor U24349 (N_24349,N_22922,N_23689);
nor U24350 (N_24350,N_23447,N_22870);
and U24351 (N_24351,N_22873,N_23430);
and U24352 (N_24352,N_23843,N_23124);
nor U24353 (N_24353,N_23670,N_22999);
nand U24354 (N_24354,N_23488,N_23992);
or U24355 (N_24355,N_23704,N_23985);
nor U24356 (N_24356,N_23361,N_23265);
nand U24357 (N_24357,N_22807,N_23131);
or U24358 (N_24358,N_23666,N_23092);
nor U24359 (N_24359,N_23716,N_23346);
xnor U24360 (N_24360,N_23954,N_23441);
and U24361 (N_24361,N_23663,N_22934);
or U24362 (N_24362,N_23797,N_23168);
nor U24363 (N_24363,N_23383,N_23489);
nor U24364 (N_24364,N_23491,N_23634);
xor U24365 (N_24365,N_23937,N_23075);
nor U24366 (N_24366,N_23385,N_23648);
and U24367 (N_24367,N_23870,N_23540);
nand U24368 (N_24368,N_23564,N_22889);
nor U24369 (N_24369,N_23665,N_23280);
or U24370 (N_24370,N_23483,N_23579);
nand U24371 (N_24371,N_22821,N_23946);
xnor U24372 (N_24372,N_23076,N_23963);
and U24373 (N_24373,N_23286,N_23248);
and U24374 (N_24374,N_23107,N_23770);
nand U24375 (N_24375,N_23462,N_22814);
and U24376 (N_24376,N_23254,N_23456);
nor U24377 (N_24377,N_23035,N_23672);
nor U24378 (N_24378,N_23432,N_23679);
and U24379 (N_24379,N_23644,N_23596);
xnor U24380 (N_24380,N_23860,N_23193);
nand U24381 (N_24381,N_23571,N_23517);
or U24382 (N_24382,N_23534,N_23152);
or U24383 (N_24383,N_23712,N_23202);
or U24384 (N_24384,N_23725,N_23320);
or U24385 (N_24385,N_23446,N_23499);
or U24386 (N_24386,N_22854,N_23578);
nor U24387 (N_24387,N_23390,N_23723);
and U24388 (N_24388,N_23880,N_23020);
and U24389 (N_24389,N_23114,N_23060);
or U24390 (N_24390,N_23464,N_23765);
nor U24391 (N_24391,N_23760,N_23695);
and U24392 (N_24392,N_23535,N_23189);
nor U24393 (N_24393,N_22860,N_23805);
xnor U24394 (N_24394,N_23553,N_23255);
or U24395 (N_24395,N_22855,N_23642);
nand U24396 (N_24396,N_23426,N_23947);
nor U24397 (N_24397,N_22823,N_23792);
and U24398 (N_24398,N_23425,N_23969);
nor U24399 (N_24399,N_23509,N_23755);
xnor U24400 (N_24400,N_22813,N_23345);
xnor U24401 (N_24401,N_22837,N_23010);
xor U24402 (N_24402,N_23884,N_22843);
xnor U24403 (N_24403,N_23952,N_23279);
and U24404 (N_24404,N_23328,N_23288);
xnor U24405 (N_24405,N_23125,N_23587);
and U24406 (N_24406,N_23479,N_23808);
and U24407 (N_24407,N_23766,N_23605);
and U24408 (N_24408,N_23270,N_23196);
nand U24409 (N_24409,N_23090,N_23410);
nor U24410 (N_24410,N_23940,N_23586);
or U24411 (N_24411,N_23431,N_23621);
nand U24412 (N_24412,N_23468,N_23732);
nor U24413 (N_24413,N_23120,N_23144);
and U24414 (N_24414,N_23994,N_23848);
xor U24415 (N_24415,N_23445,N_22801);
nor U24416 (N_24416,N_23824,N_23608);
nand U24417 (N_24417,N_23167,N_23800);
nor U24418 (N_24418,N_23203,N_23205);
nor U24419 (N_24419,N_22942,N_23996);
xnor U24420 (N_24420,N_23764,N_23419);
and U24421 (N_24421,N_23901,N_23891);
or U24422 (N_24422,N_23993,N_23735);
and U24423 (N_24423,N_23680,N_22880);
and U24424 (N_24424,N_23836,N_23304);
nand U24425 (N_24425,N_23750,N_23611);
or U24426 (N_24426,N_23321,N_23059);
or U24427 (N_24427,N_22890,N_23164);
xor U24428 (N_24428,N_23627,N_22808);
and U24429 (N_24429,N_22816,N_23527);
xor U24430 (N_24430,N_23959,N_23058);
xnor U24431 (N_24431,N_23570,N_23165);
or U24432 (N_24432,N_22850,N_23769);
and U24433 (N_24433,N_23300,N_23194);
nand U24434 (N_24434,N_23391,N_22864);
nand U24435 (N_24435,N_23150,N_23965);
and U24436 (N_24436,N_23348,N_23710);
xnor U24437 (N_24437,N_23434,N_23091);
nor U24438 (N_24438,N_22903,N_22938);
xnor U24439 (N_24439,N_23949,N_23101);
nor U24440 (N_24440,N_23021,N_23691);
or U24441 (N_24441,N_22935,N_22984);
nand U24442 (N_24442,N_22926,N_23003);
nor U24443 (N_24443,N_23864,N_22902);
nand U24444 (N_24444,N_23461,N_23526);
nand U24445 (N_24445,N_23796,N_23554);
and U24446 (N_24446,N_23519,N_23799);
or U24447 (N_24447,N_23537,N_23154);
nand U24448 (N_24448,N_23420,N_23890);
nand U24449 (N_24449,N_23616,N_23811);
or U24450 (N_24450,N_23790,N_23508);
xor U24451 (N_24451,N_23814,N_23213);
xor U24452 (N_24452,N_23178,N_23929);
nor U24453 (N_24453,N_23112,N_23436);
and U24454 (N_24454,N_23546,N_23089);
and U24455 (N_24455,N_23576,N_23029);
nand U24456 (N_24456,N_23833,N_23801);
and U24457 (N_24457,N_23497,N_22802);
or U24458 (N_24458,N_23810,N_23997);
nand U24459 (N_24459,N_23896,N_23274);
xnor U24460 (N_24460,N_23630,N_23701);
or U24461 (N_24461,N_23907,N_22991);
nor U24462 (N_24462,N_23268,N_23928);
and U24463 (N_24463,N_23780,N_23573);
xnor U24464 (N_24464,N_23806,N_23087);
nor U24465 (N_24465,N_23788,N_23310);
xor U24466 (N_24466,N_23064,N_23396);
nand U24467 (N_24467,N_22863,N_23726);
nand U24468 (N_24468,N_23470,N_23768);
nor U24469 (N_24469,N_23037,N_23459);
nor U24470 (N_24470,N_22862,N_22941);
and U24471 (N_24471,N_23936,N_23043);
xor U24472 (N_24472,N_22956,N_22876);
nor U24473 (N_24473,N_23171,N_23917);
and U24474 (N_24474,N_22817,N_22844);
or U24475 (N_24475,N_23285,N_22901);
and U24476 (N_24476,N_23622,N_23212);
nand U24477 (N_24477,N_23500,N_23054);
nand U24478 (N_24478,N_23601,N_22822);
nand U24479 (N_24479,N_23738,N_23417);
or U24480 (N_24480,N_23042,N_23036);
and U24481 (N_24481,N_22970,N_22977);
nand U24482 (N_24482,N_22995,N_23778);
nand U24483 (N_24483,N_23369,N_23299);
or U24484 (N_24484,N_23115,N_23277);
xor U24485 (N_24485,N_23368,N_22928);
and U24486 (N_24486,N_23912,N_22829);
nor U24487 (N_24487,N_23287,N_23492);
and U24488 (N_24488,N_23307,N_23562);
xnor U24489 (N_24489,N_23816,N_23395);
nor U24490 (N_24490,N_23561,N_23471);
or U24491 (N_24491,N_23635,N_23435);
or U24492 (N_24492,N_23163,N_23727);
nor U24493 (N_24493,N_23269,N_23002);
xor U24494 (N_24494,N_23099,N_23135);
or U24495 (N_24495,N_23583,N_23775);
or U24496 (N_24496,N_22827,N_23238);
or U24497 (N_24497,N_23828,N_23530);
xnor U24498 (N_24498,N_22826,N_22946);
and U24499 (N_24499,N_23538,N_22936);
nor U24500 (N_24500,N_22989,N_23389);
xor U24501 (N_24501,N_23906,N_23687);
and U24502 (N_24502,N_23510,N_23697);
nor U24503 (N_24503,N_22997,N_23149);
and U24504 (N_24504,N_23062,N_23413);
or U24505 (N_24505,N_23376,N_23319);
nor U24506 (N_24506,N_23802,N_23057);
or U24507 (N_24507,N_23334,N_23326);
xnor U24508 (N_24508,N_23231,N_23331);
nand U24509 (N_24509,N_23636,N_22838);
xnor U24510 (N_24510,N_23309,N_22806);
nor U24511 (N_24511,N_23121,N_23224);
nand U24512 (N_24512,N_23474,N_23272);
nand U24513 (N_24513,N_23458,N_23599);
nand U24514 (N_24514,N_23998,N_23660);
xor U24515 (N_24515,N_23227,N_23187);
xnor U24516 (N_24516,N_22969,N_23729);
and U24517 (N_24517,N_23846,N_23733);
nor U24518 (N_24518,N_23547,N_23173);
nor U24519 (N_24519,N_23015,N_23633);
xnor U24520 (N_24520,N_23983,N_23549);
nor U24521 (N_24521,N_23708,N_23749);
xor U24522 (N_24522,N_23988,N_23999);
nor U24523 (N_24523,N_23343,N_23424);
and U24524 (N_24524,N_23337,N_23722);
nand U24525 (N_24525,N_23025,N_22911);
nand U24526 (N_24526,N_23452,N_23214);
or U24527 (N_24527,N_23026,N_23699);
nand U24528 (N_24528,N_22851,N_23911);
nand U24529 (N_24529,N_23677,N_22914);
nand U24530 (N_24530,N_23364,N_23813);
and U24531 (N_24531,N_23148,N_23569);
nand U24532 (N_24532,N_22899,N_22896);
or U24533 (N_24533,N_23787,N_23185);
nand U24534 (N_24534,N_23686,N_22927);
and U24535 (N_24535,N_23440,N_23233);
and U24536 (N_24536,N_23118,N_23625);
and U24537 (N_24537,N_23545,N_23844);
xor U24538 (N_24538,N_23702,N_23126);
xor U24539 (N_24539,N_22959,N_23088);
nand U24540 (N_24540,N_23881,N_23590);
and U24541 (N_24541,N_23005,N_22898);
nor U24542 (N_24542,N_23960,N_22887);
nor U24543 (N_24543,N_23030,N_23373);
nand U24544 (N_24544,N_23941,N_23668);
xor U24545 (N_24545,N_23102,N_23289);
nand U24546 (N_24546,N_23498,N_22835);
or U24547 (N_24547,N_22950,N_23166);
or U24548 (N_24548,N_23866,N_23357);
nor U24549 (N_24549,N_23350,N_23367);
or U24550 (N_24550,N_23617,N_23253);
xor U24551 (N_24551,N_22812,N_23793);
nor U24552 (N_24552,N_23401,N_23438);
nor U24553 (N_24553,N_23629,N_22966);
and U24554 (N_24554,N_22831,N_23234);
or U24555 (N_24555,N_23950,N_23798);
or U24556 (N_24556,N_23895,N_23353);
xor U24557 (N_24557,N_23703,N_23141);
nor U24558 (N_24558,N_23297,N_22846);
or U24559 (N_24559,N_23718,N_23681);
nand U24560 (N_24560,N_23728,N_23188);
and U24561 (N_24561,N_22998,N_23975);
nand U24562 (N_24562,N_23480,N_23183);
xor U24563 (N_24563,N_23803,N_22982);
and U24564 (N_24564,N_23130,N_23211);
xnor U24565 (N_24565,N_23388,N_23041);
nor U24566 (N_24566,N_22918,N_23856);
or U24567 (N_24567,N_22877,N_23711);
or U24568 (N_24568,N_23973,N_23640);
or U24569 (N_24569,N_22924,N_23528);
and U24570 (N_24570,N_23217,N_23308);
xnor U24571 (N_24571,N_22921,N_23013);
xor U24572 (N_24572,N_23423,N_23849);
or U24573 (N_24573,N_23512,N_23414);
xnor U24574 (N_24574,N_22893,N_23673);
and U24575 (N_24575,N_23595,N_23276);
xor U24576 (N_24576,N_23209,N_23533);
or U24577 (N_24577,N_23412,N_23580);
xnor U24578 (N_24578,N_23455,N_23009);
nor U24579 (N_24579,N_22865,N_22979);
or U24580 (N_24580,N_23375,N_23040);
xor U24581 (N_24581,N_23317,N_23055);
or U24582 (N_24582,N_23047,N_23904);
and U24583 (N_24583,N_23823,N_22871);
and U24584 (N_24584,N_23392,N_23626);
xnor U24585 (N_24585,N_23079,N_23503);
nand U24586 (N_24586,N_23982,N_23646);
and U24587 (N_24587,N_22845,N_23938);
nor U24588 (N_24588,N_22988,N_23236);
nor U24589 (N_24589,N_23325,N_23290);
and U24590 (N_24590,N_23922,N_23298);
nand U24591 (N_24591,N_23863,N_23818);
nor U24592 (N_24592,N_23830,N_23967);
and U24593 (N_24593,N_23100,N_23651);
nor U24594 (N_24594,N_23637,N_23821);
nor U24595 (N_24595,N_22930,N_22939);
nor U24596 (N_24596,N_23779,N_23869);
nor U24597 (N_24597,N_23516,N_23377);
and U24598 (N_24598,N_22836,N_22945);
nand U24599 (N_24599,N_23110,N_22874);
nor U24600 (N_24600,N_23461,N_23554);
nand U24601 (N_24601,N_22858,N_23877);
nand U24602 (N_24602,N_23418,N_22997);
and U24603 (N_24603,N_23354,N_23340);
and U24604 (N_24604,N_23353,N_23991);
xor U24605 (N_24605,N_23714,N_23808);
or U24606 (N_24606,N_23485,N_22841);
and U24607 (N_24607,N_23698,N_23228);
and U24608 (N_24608,N_22859,N_23408);
nor U24609 (N_24609,N_23074,N_23644);
xor U24610 (N_24610,N_23953,N_23757);
nand U24611 (N_24611,N_23874,N_23345);
or U24612 (N_24612,N_23172,N_22955);
and U24613 (N_24613,N_23895,N_22808);
and U24614 (N_24614,N_23302,N_23210);
and U24615 (N_24615,N_23381,N_23837);
nor U24616 (N_24616,N_22906,N_23533);
or U24617 (N_24617,N_23018,N_23826);
xnor U24618 (N_24618,N_23367,N_23505);
xor U24619 (N_24619,N_23966,N_23182);
xnor U24620 (N_24620,N_23609,N_23545);
or U24621 (N_24621,N_23097,N_23660);
or U24622 (N_24622,N_23518,N_23609);
xnor U24623 (N_24623,N_23960,N_23463);
or U24624 (N_24624,N_23795,N_22872);
xor U24625 (N_24625,N_23500,N_23654);
nor U24626 (N_24626,N_23473,N_23010);
xnor U24627 (N_24627,N_23406,N_23123);
and U24628 (N_24628,N_23884,N_23380);
nor U24629 (N_24629,N_23950,N_23630);
or U24630 (N_24630,N_23963,N_23365);
xor U24631 (N_24631,N_23597,N_23949);
nor U24632 (N_24632,N_23967,N_23996);
or U24633 (N_24633,N_23665,N_23941);
or U24634 (N_24634,N_23415,N_23524);
nor U24635 (N_24635,N_23240,N_23911);
xnor U24636 (N_24636,N_23518,N_23435);
nor U24637 (N_24637,N_23776,N_23872);
or U24638 (N_24638,N_22880,N_23555);
nor U24639 (N_24639,N_23802,N_23505);
or U24640 (N_24640,N_23710,N_23044);
xnor U24641 (N_24641,N_23923,N_22859);
xor U24642 (N_24642,N_23044,N_23088);
nor U24643 (N_24643,N_23591,N_23963);
and U24644 (N_24644,N_23774,N_23445);
nor U24645 (N_24645,N_23519,N_23574);
xor U24646 (N_24646,N_22864,N_23613);
nor U24647 (N_24647,N_23793,N_23628);
xnor U24648 (N_24648,N_23535,N_23660);
or U24649 (N_24649,N_23671,N_22807);
nor U24650 (N_24650,N_23703,N_23914);
nor U24651 (N_24651,N_23551,N_23932);
xnor U24652 (N_24652,N_23697,N_23787);
nand U24653 (N_24653,N_23195,N_23500);
nor U24654 (N_24654,N_23661,N_22937);
nand U24655 (N_24655,N_23283,N_23491);
or U24656 (N_24656,N_23316,N_23271);
xnor U24657 (N_24657,N_23603,N_23852);
nand U24658 (N_24658,N_23463,N_23011);
nor U24659 (N_24659,N_23094,N_23727);
or U24660 (N_24660,N_22916,N_23484);
nor U24661 (N_24661,N_22881,N_22883);
nor U24662 (N_24662,N_23925,N_23277);
or U24663 (N_24663,N_23408,N_23523);
or U24664 (N_24664,N_23244,N_23777);
xnor U24665 (N_24665,N_23594,N_23290);
xor U24666 (N_24666,N_22996,N_22954);
and U24667 (N_24667,N_23269,N_23495);
nor U24668 (N_24668,N_23594,N_23195);
xnor U24669 (N_24669,N_23644,N_23822);
nand U24670 (N_24670,N_23396,N_23050);
nand U24671 (N_24671,N_23412,N_23022);
nor U24672 (N_24672,N_23197,N_23706);
xor U24673 (N_24673,N_23285,N_23920);
and U24674 (N_24674,N_23965,N_23249);
nand U24675 (N_24675,N_23876,N_23500);
nor U24676 (N_24676,N_23540,N_23484);
nand U24677 (N_24677,N_23919,N_23772);
and U24678 (N_24678,N_23005,N_23393);
and U24679 (N_24679,N_23922,N_23054);
or U24680 (N_24680,N_23793,N_23213);
and U24681 (N_24681,N_23510,N_23004);
xnor U24682 (N_24682,N_23449,N_23442);
xor U24683 (N_24683,N_23821,N_23647);
nand U24684 (N_24684,N_23385,N_23548);
or U24685 (N_24685,N_23548,N_23193);
or U24686 (N_24686,N_23998,N_23825);
nand U24687 (N_24687,N_22878,N_23480);
nand U24688 (N_24688,N_23980,N_22994);
nand U24689 (N_24689,N_23490,N_23801);
and U24690 (N_24690,N_23829,N_23754);
xnor U24691 (N_24691,N_23501,N_23941);
nor U24692 (N_24692,N_23161,N_23954);
xnor U24693 (N_24693,N_23303,N_23691);
nor U24694 (N_24694,N_22988,N_23734);
nand U24695 (N_24695,N_23606,N_23731);
nor U24696 (N_24696,N_23347,N_22825);
nor U24697 (N_24697,N_22919,N_22832);
nor U24698 (N_24698,N_23737,N_23611);
or U24699 (N_24699,N_23786,N_23164);
nor U24700 (N_24700,N_23802,N_23475);
xnor U24701 (N_24701,N_23878,N_22901);
or U24702 (N_24702,N_22875,N_22893);
nand U24703 (N_24703,N_23453,N_23342);
and U24704 (N_24704,N_23042,N_23396);
nor U24705 (N_24705,N_22966,N_23061);
and U24706 (N_24706,N_23962,N_23660);
or U24707 (N_24707,N_22922,N_23253);
nor U24708 (N_24708,N_23454,N_23435);
nor U24709 (N_24709,N_23205,N_23547);
or U24710 (N_24710,N_23060,N_23467);
nand U24711 (N_24711,N_23621,N_23122);
xor U24712 (N_24712,N_23127,N_23941);
and U24713 (N_24713,N_23608,N_23814);
nand U24714 (N_24714,N_23668,N_23588);
and U24715 (N_24715,N_23057,N_23506);
nand U24716 (N_24716,N_23231,N_22829);
and U24717 (N_24717,N_23181,N_23010);
and U24718 (N_24718,N_23739,N_23974);
and U24719 (N_24719,N_23143,N_23040);
nor U24720 (N_24720,N_23504,N_23119);
nor U24721 (N_24721,N_23436,N_23060);
nand U24722 (N_24722,N_23602,N_23907);
and U24723 (N_24723,N_23635,N_23900);
xor U24724 (N_24724,N_23351,N_23214);
nor U24725 (N_24725,N_23051,N_23035);
xnor U24726 (N_24726,N_23296,N_23708);
nor U24727 (N_24727,N_23398,N_23027);
and U24728 (N_24728,N_22973,N_23526);
nor U24729 (N_24729,N_23626,N_23163);
or U24730 (N_24730,N_23071,N_23058);
or U24731 (N_24731,N_23920,N_23396);
nor U24732 (N_24732,N_23466,N_23962);
xor U24733 (N_24733,N_23263,N_23052);
nor U24734 (N_24734,N_23626,N_23596);
nor U24735 (N_24735,N_23225,N_23209);
xor U24736 (N_24736,N_23616,N_23693);
or U24737 (N_24737,N_23979,N_22920);
or U24738 (N_24738,N_22817,N_23574);
and U24739 (N_24739,N_23219,N_22897);
and U24740 (N_24740,N_23910,N_22807);
or U24741 (N_24741,N_23529,N_23803);
xnor U24742 (N_24742,N_23140,N_23063);
nand U24743 (N_24743,N_23010,N_23969);
xor U24744 (N_24744,N_23308,N_23523);
nand U24745 (N_24745,N_23497,N_23015);
and U24746 (N_24746,N_23675,N_23630);
nor U24747 (N_24747,N_22853,N_23603);
xnor U24748 (N_24748,N_23153,N_23401);
nand U24749 (N_24749,N_23566,N_23935);
or U24750 (N_24750,N_23193,N_23909);
and U24751 (N_24751,N_23004,N_23153);
or U24752 (N_24752,N_22837,N_23999);
nor U24753 (N_24753,N_23301,N_23941);
or U24754 (N_24754,N_23684,N_23222);
nand U24755 (N_24755,N_23636,N_23675);
nand U24756 (N_24756,N_23477,N_23521);
xnor U24757 (N_24757,N_23644,N_23560);
xor U24758 (N_24758,N_23634,N_23888);
or U24759 (N_24759,N_23312,N_23252);
nor U24760 (N_24760,N_23092,N_23135);
or U24761 (N_24761,N_23819,N_23042);
and U24762 (N_24762,N_23391,N_23578);
or U24763 (N_24763,N_23720,N_22932);
nor U24764 (N_24764,N_23045,N_23776);
and U24765 (N_24765,N_23343,N_23560);
nand U24766 (N_24766,N_23169,N_22955);
xor U24767 (N_24767,N_23007,N_22910);
xor U24768 (N_24768,N_23316,N_23054);
or U24769 (N_24769,N_23009,N_23847);
and U24770 (N_24770,N_23840,N_22983);
and U24771 (N_24771,N_23012,N_23788);
and U24772 (N_24772,N_23897,N_23471);
nand U24773 (N_24773,N_23612,N_23917);
xor U24774 (N_24774,N_23750,N_22823);
nand U24775 (N_24775,N_23994,N_23265);
nor U24776 (N_24776,N_23747,N_22881);
nand U24777 (N_24777,N_23838,N_23568);
or U24778 (N_24778,N_23277,N_23773);
or U24779 (N_24779,N_23034,N_22899);
nand U24780 (N_24780,N_23008,N_23423);
nor U24781 (N_24781,N_23082,N_22846);
xnor U24782 (N_24782,N_23966,N_23207);
xnor U24783 (N_24783,N_23853,N_23274);
or U24784 (N_24784,N_23047,N_23857);
nor U24785 (N_24785,N_23687,N_23276);
and U24786 (N_24786,N_23509,N_23559);
xnor U24787 (N_24787,N_23651,N_22851);
xnor U24788 (N_24788,N_23541,N_23776);
and U24789 (N_24789,N_23522,N_23149);
and U24790 (N_24790,N_23565,N_23101);
nand U24791 (N_24791,N_23237,N_22930);
nor U24792 (N_24792,N_23155,N_22971);
nor U24793 (N_24793,N_23738,N_23669);
xor U24794 (N_24794,N_23013,N_23363);
nand U24795 (N_24795,N_23575,N_23714);
nor U24796 (N_24796,N_23798,N_23704);
xnor U24797 (N_24797,N_23208,N_23133);
or U24798 (N_24798,N_23425,N_23150);
nor U24799 (N_24799,N_23793,N_23241);
xnor U24800 (N_24800,N_23146,N_23327);
or U24801 (N_24801,N_22953,N_23422);
nand U24802 (N_24802,N_23493,N_22954);
or U24803 (N_24803,N_23271,N_23850);
and U24804 (N_24804,N_23268,N_23872);
xor U24805 (N_24805,N_23082,N_23731);
nand U24806 (N_24806,N_23304,N_23531);
or U24807 (N_24807,N_22862,N_23175);
or U24808 (N_24808,N_22939,N_23025);
or U24809 (N_24809,N_23432,N_23608);
nor U24810 (N_24810,N_23784,N_23889);
nor U24811 (N_24811,N_23413,N_22899);
or U24812 (N_24812,N_23621,N_23048);
or U24813 (N_24813,N_23029,N_23198);
nor U24814 (N_24814,N_22875,N_23662);
nand U24815 (N_24815,N_22868,N_23538);
nor U24816 (N_24816,N_22983,N_23434);
nor U24817 (N_24817,N_22890,N_23715);
xnor U24818 (N_24818,N_23552,N_23227);
and U24819 (N_24819,N_23688,N_22975);
nor U24820 (N_24820,N_23653,N_23028);
xnor U24821 (N_24821,N_22990,N_22866);
or U24822 (N_24822,N_23920,N_23794);
or U24823 (N_24823,N_23506,N_23073);
nor U24824 (N_24824,N_23446,N_23241);
nand U24825 (N_24825,N_23543,N_23766);
nand U24826 (N_24826,N_22862,N_23949);
or U24827 (N_24827,N_23446,N_23452);
or U24828 (N_24828,N_23228,N_22934);
or U24829 (N_24829,N_23095,N_23561);
and U24830 (N_24830,N_23903,N_23719);
nor U24831 (N_24831,N_23270,N_23850);
or U24832 (N_24832,N_23615,N_23614);
xnor U24833 (N_24833,N_22853,N_23438);
or U24834 (N_24834,N_23340,N_23495);
xor U24835 (N_24835,N_22967,N_22989);
nand U24836 (N_24836,N_23296,N_23886);
or U24837 (N_24837,N_22852,N_23438);
nor U24838 (N_24838,N_23647,N_22865);
and U24839 (N_24839,N_23982,N_23816);
nor U24840 (N_24840,N_23592,N_23623);
or U24841 (N_24841,N_23495,N_23926);
nand U24842 (N_24842,N_23685,N_23097);
xnor U24843 (N_24843,N_23539,N_23853);
nand U24844 (N_24844,N_23506,N_23624);
nor U24845 (N_24845,N_23875,N_23985);
xnor U24846 (N_24846,N_22833,N_23292);
and U24847 (N_24847,N_23447,N_23994);
nor U24848 (N_24848,N_23363,N_23550);
or U24849 (N_24849,N_23108,N_22906);
xor U24850 (N_24850,N_22928,N_23447);
and U24851 (N_24851,N_23043,N_22932);
or U24852 (N_24852,N_23573,N_23713);
nor U24853 (N_24853,N_23689,N_23000);
nand U24854 (N_24854,N_22840,N_23128);
nand U24855 (N_24855,N_23872,N_23730);
or U24856 (N_24856,N_23548,N_23711);
xor U24857 (N_24857,N_23021,N_23081);
or U24858 (N_24858,N_22979,N_23658);
nor U24859 (N_24859,N_23811,N_23891);
xnor U24860 (N_24860,N_22953,N_22902);
nand U24861 (N_24861,N_23965,N_23351);
nand U24862 (N_24862,N_23801,N_23541);
or U24863 (N_24863,N_23179,N_22894);
nor U24864 (N_24864,N_23692,N_23901);
and U24865 (N_24865,N_23157,N_23974);
xnor U24866 (N_24866,N_23152,N_23623);
xnor U24867 (N_24867,N_22911,N_23632);
nor U24868 (N_24868,N_22992,N_22914);
or U24869 (N_24869,N_22886,N_22824);
nand U24870 (N_24870,N_23404,N_22882);
xor U24871 (N_24871,N_23512,N_23246);
nor U24872 (N_24872,N_22996,N_22857);
and U24873 (N_24873,N_23991,N_23762);
xor U24874 (N_24874,N_23258,N_23220);
or U24875 (N_24875,N_23931,N_22956);
xnor U24876 (N_24876,N_23434,N_22902);
nor U24877 (N_24877,N_22912,N_22870);
nor U24878 (N_24878,N_23574,N_23495);
and U24879 (N_24879,N_23956,N_23233);
xnor U24880 (N_24880,N_23183,N_23586);
and U24881 (N_24881,N_23943,N_23663);
nor U24882 (N_24882,N_23397,N_23881);
or U24883 (N_24883,N_23298,N_23642);
nand U24884 (N_24884,N_23793,N_23707);
or U24885 (N_24885,N_22849,N_23799);
xor U24886 (N_24886,N_23513,N_22891);
xor U24887 (N_24887,N_23529,N_23723);
nand U24888 (N_24888,N_23431,N_22959);
or U24889 (N_24889,N_22831,N_23614);
xor U24890 (N_24890,N_22941,N_22853);
and U24891 (N_24891,N_23453,N_22840);
xor U24892 (N_24892,N_23888,N_23287);
or U24893 (N_24893,N_23315,N_22810);
nor U24894 (N_24894,N_23461,N_22933);
nor U24895 (N_24895,N_23159,N_23439);
nand U24896 (N_24896,N_23686,N_23614);
and U24897 (N_24897,N_23148,N_23945);
or U24898 (N_24898,N_22929,N_23624);
and U24899 (N_24899,N_23621,N_23923);
xnor U24900 (N_24900,N_23346,N_23874);
xor U24901 (N_24901,N_22858,N_23447);
nor U24902 (N_24902,N_23817,N_23240);
or U24903 (N_24903,N_23614,N_23250);
and U24904 (N_24904,N_23609,N_22982);
or U24905 (N_24905,N_23563,N_23026);
xor U24906 (N_24906,N_23560,N_23730);
or U24907 (N_24907,N_23995,N_23865);
nor U24908 (N_24908,N_23870,N_23906);
nor U24909 (N_24909,N_23858,N_23895);
nand U24910 (N_24910,N_23813,N_23682);
nor U24911 (N_24911,N_23342,N_23701);
nand U24912 (N_24912,N_23553,N_22868);
nand U24913 (N_24913,N_23269,N_23534);
nor U24914 (N_24914,N_23584,N_23050);
and U24915 (N_24915,N_23880,N_22976);
nand U24916 (N_24916,N_23806,N_23866);
or U24917 (N_24917,N_23297,N_23294);
nand U24918 (N_24918,N_23850,N_23336);
xnor U24919 (N_24919,N_22938,N_23531);
nor U24920 (N_24920,N_23332,N_23700);
nor U24921 (N_24921,N_22870,N_22964);
or U24922 (N_24922,N_23673,N_22810);
xnor U24923 (N_24923,N_23019,N_22974);
and U24924 (N_24924,N_23616,N_23741);
xnor U24925 (N_24925,N_23478,N_23880);
nand U24926 (N_24926,N_23168,N_23463);
and U24927 (N_24927,N_23006,N_23205);
nand U24928 (N_24928,N_23893,N_23007);
xor U24929 (N_24929,N_23721,N_23895);
nor U24930 (N_24930,N_23702,N_23809);
nor U24931 (N_24931,N_23186,N_22949);
or U24932 (N_24932,N_23749,N_23532);
or U24933 (N_24933,N_23124,N_22930);
xor U24934 (N_24934,N_23593,N_23817);
or U24935 (N_24935,N_23268,N_22972);
xor U24936 (N_24936,N_22969,N_23139);
and U24937 (N_24937,N_23303,N_23338);
nor U24938 (N_24938,N_23942,N_23257);
nand U24939 (N_24939,N_23720,N_23781);
and U24940 (N_24940,N_23699,N_22993);
or U24941 (N_24941,N_23265,N_23018);
and U24942 (N_24942,N_23270,N_23910);
nand U24943 (N_24943,N_23299,N_22945);
nor U24944 (N_24944,N_23114,N_23326);
xor U24945 (N_24945,N_23872,N_23159);
nand U24946 (N_24946,N_23212,N_22813);
and U24947 (N_24947,N_23821,N_23167);
or U24948 (N_24948,N_22994,N_23179);
nor U24949 (N_24949,N_23748,N_22940);
nand U24950 (N_24950,N_23029,N_23927);
or U24951 (N_24951,N_23744,N_23144);
xnor U24952 (N_24952,N_23212,N_22842);
nand U24953 (N_24953,N_22926,N_23127);
nor U24954 (N_24954,N_23976,N_23034);
nor U24955 (N_24955,N_23749,N_22858);
nand U24956 (N_24956,N_23625,N_23778);
and U24957 (N_24957,N_22878,N_23027);
xnor U24958 (N_24958,N_23832,N_22910);
xor U24959 (N_24959,N_23885,N_23317);
and U24960 (N_24960,N_23112,N_23760);
and U24961 (N_24961,N_23369,N_23170);
or U24962 (N_24962,N_23732,N_23353);
and U24963 (N_24963,N_22917,N_23804);
or U24964 (N_24964,N_22984,N_23686);
nand U24965 (N_24965,N_23148,N_23732);
nand U24966 (N_24966,N_23393,N_23073);
nor U24967 (N_24967,N_22996,N_23652);
xor U24968 (N_24968,N_23414,N_23898);
nor U24969 (N_24969,N_23908,N_22897);
nor U24970 (N_24970,N_23841,N_23962);
nand U24971 (N_24971,N_22882,N_23092);
and U24972 (N_24972,N_23148,N_23371);
nand U24973 (N_24973,N_23972,N_23313);
or U24974 (N_24974,N_23605,N_23234);
nand U24975 (N_24975,N_23158,N_23072);
or U24976 (N_24976,N_23530,N_23117);
nand U24977 (N_24977,N_23070,N_23782);
nor U24978 (N_24978,N_23535,N_23356);
xnor U24979 (N_24979,N_23842,N_23720);
nor U24980 (N_24980,N_23564,N_23495);
or U24981 (N_24981,N_22950,N_23602);
nand U24982 (N_24982,N_23220,N_22912);
nand U24983 (N_24983,N_22906,N_23987);
or U24984 (N_24984,N_23250,N_23253);
nand U24985 (N_24985,N_22800,N_23721);
xnor U24986 (N_24986,N_23919,N_23954);
or U24987 (N_24987,N_23798,N_23963);
and U24988 (N_24988,N_23313,N_22844);
and U24989 (N_24989,N_23238,N_23878);
or U24990 (N_24990,N_23950,N_23041);
nor U24991 (N_24991,N_23619,N_23723);
xor U24992 (N_24992,N_23182,N_23591);
nor U24993 (N_24993,N_23743,N_23207);
or U24994 (N_24994,N_23743,N_23106);
nand U24995 (N_24995,N_22837,N_23910);
nand U24996 (N_24996,N_23537,N_23603);
and U24997 (N_24997,N_23468,N_22820);
and U24998 (N_24998,N_23242,N_23907);
and U24999 (N_24999,N_23480,N_23081);
or U25000 (N_25000,N_23168,N_23675);
xor U25001 (N_25001,N_23665,N_23303);
nor U25002 (N_25002,N_23030,N_22826);
nand U25003 (N_25003,N_23098,N_22946);
nor U25004 (N_25004,N_23820,N_23022);
and U25005 (N_25005,N_23234,N_23321);
nor U25006 (N_25006,N_22814,N_23692);
nor U25007 (N_25007,N_23577,N_23583);
nor U25008 (N_25008,N_23572,N_22994);
nor U25009 (N_25009,N_22800,N_23725);
and U25010 (N_25010,N_23720,N_23452);
nand U25011 (N_25011,N_23952,N_22963);
or U25012 (N_25012,N_23841,N_22826);
or U25013 (N_25013,N_22894,N_23521);
nand U25014 (N_25014,N_23698,N_23284);
nor U25015 (N_25015,N_23691,N_23675);
or U25016 (N_25016,N_23217,N_23530);
nor U25017 (N_25017,N_23629,N_22834);
xnor U25018 (N_25018,N_23165,N_22955);
nor U25019 (N_25019,N_23188,N_22904);
nor U25020 (N_25020,N_23764,N_23636);
and U25021 (N_25021,N_23650,N_23697);
nand U25022 (N_25022,N_23738,N_22971);
or U25023 (N_25023,N_23122,N_23002);
nand U25024 (N_25024,N_22857,N_23088);
nand U25025 (N_25025,N_23173,N_23023);
and U25026 (N_25026,N_23073,N_23370);
and U25027 (N_25027,N_23917,N_22950);
xor U25028 (N_25028,N_23958,N_23111);
nand U25029 (N_25029,N_23234,N_23995);
nor U25030 (N_25030,N_23052,N_23819);
and U25031 (N_25031,N_23341,N_23334);
nor U25032 (N_25032,N_23330,N_23766);
nand U25033 (N_25033,N_23499,N_23822);
nand U25034 (N_25034,N_23369,N_23657);
and U25035 (N_25035,N_23654,N_22867);
and U25036 (N_25036,N_23010,N_23255);
nor U25037 (N_25037,N_22883,N_23895);
nor U25038 (N_25038,N_23384,N_23654);
xor U25039 (N_25039,N_23561,N_23686);
xor U25040 (N_25040,N_23103,N_23193);
xnor U25041 (N_25041,N_23766,N_23045);
nand U25042 (N_25042,N_23421,N_23467);
nor U25043 (N_25043,N_23041,N_22982);
xor U25044 (N_25044,N_23589,N_23366);
nor U25045 (N_25045,N_23755,N_23302);
nand U25046 (N_25046,N_22951,N_23314);
and U25047 (N_25047,N_23740,N_23638);
or U25048 (N_25048,N_23682,N_23737);
nor U25049 (N_25049,N_23926,N_22846);
and U25050 (N_25050,N_23168,N_23230);
nor U25051 (N_25051,N_23287,N_22920);
and U25052 (N_25052,N_23424,N_23717);
nand U25053 (N_25053,N_23055,N_23839);
xor U25054 (N_25054,N_23714,N_23538);
xor U25055 (N_25055,N_23582,N_23340);
nand U25056 (N_25056,N_23272,N_23152);
xor U25057 (N_25057,N_23900,N_23086);
nor U25058 (N_25058,N_22906,N_23283);
nor U25059 (N_25059,N_23241,N_23196);
or U25060 (N_25060,N_23641,N_23648);
xnor U25061 (N_25061,N_23870,N_23764);
xor U25062 (N_25062,N_22864,N_23169);
nor U25063 (N_25063,N_23900,N_22957);
or U25064 (N_25064,N_23375,N_23008);
nand U25065 (N_25065,N_23031,N_23121);
xor U25066 (N_25066,N_23213,N_22929);
nand U25067 (N_25067,N_23307,N_23311);
or U25068 (N_25068,N_23194,N_23355);
and U25069 (N_25069,N_23012,N_23373);
nand U25070 (N_25070,N_23899,N_23844);
and U25071 (N_25071,N_23711,N_23105);
nand U25072 (N_25072,N_23042,N_23588);
nor U25073 (N_25073,N_23611,N_23081);
xnor U25074 (N_25074,N_22805,N_23036);
nand U25075 (N_25075,N_23177,N_23954);
nor U25076 (N_25076,N_23598,N_23903);
xor U25077 (N_25077,N_23943,N_23486);
or U25078 (N_25078,N_23586,N_23257);
or U25079 (N_25079,N_23558,N_23661);
and U25080 (N_25080,N_22858,N_23679);
nor U25081 (N_25081,N_23714,N_23961);
or U25082 (N_25082,N_22945,N_23786);
nand U25083 (N_25083,N_22870,N_23650);
xnor U25084 (N_25084,N_23823,N_23680);
nand U25085 (N_25085,N_23620,N_23568);
or U25086 (N_25086,N_23682,N_23799);
nor U25087 (N_25087,N_23001,N_23248);
xor U25088 (N_25088,N_23693,N_22918);
nor U25089 (N_25089,N_22916,N_23275);
nand U25090 (N_25090,N_23645,N_22981);
and U25091 (N_25091,N_23418,N_23203);
and U25092 (N_25092,N_22933,N_23343);
nand U25093 (N_25093,N_23576,N_23969);
nor U25094 (N_25094,N_23572,N_23032);
nand U25095 (N_25095,N_23066,N_22920);
or U25096 (N_25096,N_23339,N_23691);
nor U25097 (N_25097,N_22957,N_23418);
nand U25098 (N_25098,N_23200,N_23147);
xor U25099 (N_25099,N_23053,N_22823);
or U25100 (N_25100,N_23454,N_23198);
xor U25101 (N_25101,N_22813,N_23690);
nor U25102 (N_25102,N_23693,N_23326);
nor U25103 (N_25103,N_23062,N_23094);
nor U25104 (N_25104,N_23252,N_23032);
or U25105 (N_25105,N_23940,N_23032);
and U25106 (N_25106,N_23840,N_23978);
or U25107 (N_25107,N_23544,N_23575);
nor U25108 (N_25108,N_23094,N_22999);
xnor U25109 (N_25109,N_23302,N_23197);
xor U25110 (N_25110,N_23492,N_22894);
and U25111 (N_25111,N_23017,N_23291);
or U25112 (N_25112,N_22964,N_23055);
nor U25113 (N_25113,N_23350,N_23717);
and U25114 (N_25114,N_23880,N_23772);
and U25115 (N_25115,N_23033,N_23286);
nand U25116 (N_25116,N_23754,N_23372);
and U25117 (N_25117,N_23780,N_23077);
nand U25118 (N_25118,N_23365,N_23232);
xnor U25119 (N_25119,N_23846,N_23036);
xnor U25120 (N_25120,N_23209,N_23594);
and U25121 (N_25121,N_23923,N_23603);
and U25122 (N_25122,N_23731,N_23724);
nand U25123 (N_25123,N_23655,N_23260);
nand U25124 (N_25124,N_22881,N_22894);
xor U25125 (N_25125,N_22962,N_23376);
xnor U25126 (N_25126,N_23795,N_23927);
or U25127 (N_25127,N_23238,N_23439);
and U25128 (N_25128,N_23306,N_22817);
nand U25129 (N_25129,N_23352,N_23553);
or U25130 (N_25130,N_23300,N_23711);
nor U25131 (N_25131,N_22807,N_22966);
nand U25132 (N_25132,N_23297,N_23483);
nor U25133 (N_25133,N_23097,N_22910);
or U25134 (N_25134,N_23183,N_22803);
or U25135 (N_25135,N_23287,N_23479);
or U25136 (N_25136,N_22938,N_23318);
or U25137 (N_25137,N_23586,N_22805);
xor U25138 (N_25138,N_23341,N_22832);
nand U25139 (N_25139,N_23333,N_23785);
and U25140 (N_25140,N_23888,N_22910);
nand U25141 (N_25141,N_22961,N_22951);
xor U25142 (N_25142,N_23791,N_22950);
or U25143 (N_25143,N_23427,N_23283);
xnor U25144 (N_25144,N_23323,N_23068);
xnor U25145 (N_25145,N_23348,N_23506);
xor U25146 (N_25146,N_23960,N_23896);
and U25147 (N_25147,N_23388,N_23411);
or U25148 (N_25148,N_23903,N_23372);
nand U25149 (N_25149,N_23167,N_23750);
nand U25150 (N_25150,N_23570,N_23337);
xnor U25151 (N_25151,N_23887,N_23348);
or U25152 (N_25152,N_23837,N_23323);
nand U25153 (N_25153,N_23080,N_22977);
xnor U25154 (N_25154,N_22897,N_23278);
nand U25155 (N_25155,N_23355,N_23453);
or U25156 (N_25156,N_23059,N_23204);
nor U25157 (N_25157,N_23046,N_23253);
nor U25158 (N_25158,N_23704,N_23205);
nand U25159 (N_25159,N_23783,N_23642);
nor U25160 (N_25160,N_23037,N_22860);
xor U25161 (N_25161,N_23340,N_23559);
and U25162 (N_25162,N_22802,N_23120);
and U25163 (N_25163,N_23897,N_23831);
or U25164 (N_25164,N_23095,N_23742);
nand U25165 (N_25165,N_22940,N_23885);
nand U25166 (N_25166,N_22984,N_23695);
and U25167 (N_25167,N_22942,N_23930);
nand U25168 (N_25168,N_23236,N_23172);
xor U25169 (N_25169,N_23755,N_23481);
and U25170 (N_25170,N_22809,N_23140);
or U25171 (N_25171,N_23791,N_23331);
xnor U25172 (N_25172,N_22989,N_22948);
nand U25173 (N_25173,N_23204,N_23719);
nand U25174 (N_25174,N_23680,N_23911);
nand U25175 (N_25175,N_23997,N_23838);
nand U25176 (N_25176,N_23153,N_23656);
nand U25177 (N_25177,N_23113,N_22912);
and U25178 (N_25178,N_23326,N_22938);
nand U25179 (N_25179,N_23075,N_23415);
or U25180 (N_25180,N_22822,N_22821);
and U25181 (N_25181,N_23539,N_23857);
xor U25182 (N_25182,N_23374,N_23538);
nand U25183 (N_25183,N_23210,N_23142);
and U25184 (N_25184,N_23394,N_23913);
nand U25185 (N_25185,N_23954,N_23226);
and U25186 (N_25186,N_23039,N_23021);
nor U25187 (N_25187,N_23288,N_23444);
nor U25188 (N_25188,N_23549,N_23490);
and U25189 (N_25189,N_23102,N_23598);
xnor U25190 (N_25190,N_23290,N_22847);
or U25191 (N_25191,N_23499,N_23448);
nor U25192 (N_25192,N_23046,N_23015);
xor U25193 (N_25193,N_23778,N_23991);
nand U25194 (N_25194,N_23556,N_23134);
xnor U25195 (N_25195,N_23414,N_23339);
or U25196 (N_25196,N_23131,N_23983);
and U25197 (N_25197,N_23388,N_23098);
and U25198 (N_25198,N_23780,N_23428);
or U25199 (N_25199,N_23075,N_23964);
or U25200 (N_25200,N_24319,N_24935);
xor U25201 (N_25201,N_25042,N_24462);
nand U25202 (N_25202,N_24815,N_24519);
nand U25203 (N_25203,N_25054,N_24060);
or U25204 (N_25204,N_25145,N_24370);
or U25205 (N_25205,N_24418,N_25104);
or U25206 (N_25206,N_24716,N_25010);
or U25207 (N_25207,N_24910,N_24177);
nor U25208 (N_25208,N_24276,N_25172);
nand U25209 (N_25209,N_24544,N_25113);
nor U25210 (N_25210,N_24832,N_24942);
xor U25211 (N_25211,N_24753,N_24627);
xnor U25212 (N_25212,N_25147,N_24708);
xor U25213 (N_25213,N_25080,N_24775);
and U25214 (N_25214,N_24358,N_24904);
nand U25215 (N_25215,N_24897,N_24514);
nand U25216 (N_25216,N_25081,N_24950);
and U25217 (N_25217,N_24699,N_24140);
and U25218 (N_25218,N_25166,N_24311);
and U25219 (N_25219,N_24485,N_24448);
xor U25220 (N_25220,N_24978,N_24503);
xnor U25221 (N_25221,N_24908,N_24092);
nor U25222 (N_25222,N_24947,N_24575);
nand U25223 (N_25223,N_24703,N_24261);
nand U25224 (N_25224,N_24141,N_24839);
nor U25225 (N_25225,N_24225,N_24731);
xor U25226 (N_25226,N_24618,N_24610);
nand U25227 (N_25227,N_24638,N_24714);
nor U25228 (N_25228,N_24718,N_24201);
nor U25229 (N_25229,N_24037,N_24310);
nand U25230 (N_25230,N_24326,N_24659);
or U25231 (N_25231,N_24873,N_25032);
and U25232 (N_25232,N_24946,N_24142);
and U25233 (N_25233,N_24899,N_24607);
nand U25234 (N_25234,N_24224,N_24269);
or U25235 (N_25235,N_24337,N_24664);
xor U25236 (N_25236,N_24720,N_24119);
xor U25237 (N_25237,N_24958,N_24341);
or U25238 (N_25238,N_24994,N_24582);
nor U25239 (N_25239,N_24138,N_24343);
nand U25240 (N_25240,N_24813,N_24153);
xor U25241 (N_25241,N_24482,N_24905);
nand U25242 (N_25242,N_24327,N_24307);
and U25243 (N_25243,N_24635,N_24325);
xnor U25244 (N_25244,N_24324,N_24650);
nor U25245 (N_25245,N_24233,N_24205);
and U25246 (N_25246,N_25100,N_25000);
nand U25247 (N_25247,N_24644,N_25001);
nand U25248 (N_25248,N_24314,N_24105);
nand U25249 (N_25249,N_25159,N_24881);
xnor U25250 (N_25250,N_25163,N_24235);
nor U25251 (N_25251,N_24255,N_24968);
or U25252 (N_25252,N_24901,N_24374);
and U25253 (N_25253,N_24967,N_24126);
nand U25254 (N_25254,N_25011,N_24795);
nand U25255 (N_25255,N_24003,N_24336);
or U25256 (N_25256,N_24289,N_24766);
nor U25257 (N_25257,N_24214,N_24260);
nand U25258 (N_25258,N_24471,N_24675);
and U25259 (N_25259,N_24601,N_24554);
nand U25260 (N_25260,N_24211,N_24015);
nand U25261 (N_25261,N_25109,N_24587);
nor U25262 (N_25262,N_24781,N_25021);
nor U25263 (N_25263,N_24856,N_24393);
or U25264 (N_25264,N_24019,N_25112);
xor U25265 (N_25265,N_25075,N_24814);
nand U25266 (N_25266,N_24401,N_25108);
xnor U25267 (N_25267,N_24208,N_24786);
xnor U25268 (N_25268,N_25139,N_24990);
xor U25269 (N_25269,N_24243,N_24769);
and U25270 (N_25270,N_25095,N_24288);
or U25271 (N_25271,N_24646,N_24934);
or U25272 (N_25272,N_24479,N_24085);
nor U25273 (N_25273,N_24363,N_24517);
and U25274 (N_25274,N_24615,N_24980);
nor U25275 (N_25275,N_24641,N_24604);
or U25276 (N_25276,N_24427,N_25127);
xnor U25277 (N_25277,N_24398,N_24102);
and U25278 (N_25278,N_24173,N_24828);
or U25279 (N_25279,N_24898,N_24522);
xor U25280 (N_25280,N_24704,N_25162);
xor U25281 (N_25281,N_24249,N_24649);
or U25282 (N_25282,N_24526,N_24570);
or U25283 (N_25283,N_24230,N_24217);
nand U25284 (N_25284,N_25061,N_24972);
or U25285 (N_25285,N_24933,N_24316);
or U25286 (N_25286,N_24939,N_25168);
nand U25287 (N_25287,N_24512,N_24344);
xnor U25288 (N_25288,N_24606,N_25071);
xor U25289 (N_25289,N_24265,N_24889);
or U25290 (N_25290,N_24549,N_24069);
nor U25291 (N_25291,N_24868,N_25092);
xor U25292 (N_25292,N_24315,N_24189);
xor U25293 (N_25293,N_25170,N_25178);
or U25294 (N_25294,N_24473,N_24413);
nor U25295 (N_25295,N_24912,N_24500);
nor U25296 (N_25296,N_24568,N_24874);
or U25297 (N_25297,N_24981,N_24867);
nand U25298 (N_25298,N_24982,N_24932);
nand U25299 (N_25299,N_24080,N_24555);
and U25300 (N_25300,N_24672,N_24789);
nor U25301 (N_25301,N_24835,N_24228);
nor U25302 (N_25302,N_24164,N_25089);
xnor U25303 (N_25303,N_24847,N_24861);
nand U25304 (N_25304,N_24882,N_24780);
xor U25305 (N_25305,N_24262,N_24090);
xnor U25306 (N_25306,N_24452,N_24422);
nor U25307 (N_25307,N_25114,N_24109);
nor U25308 (N_25308,N_25124,N_24876);
or U25309 (N_25309,N_24654,N_24879);
or U25310 (N_25310,N_25155,N_24317);
xnor U25311 (N_25311,N_24812,N_24097);
nand U25312 (N_25312,N_24375,N_25137);
nor U25313 (N_25313,N_24588,N_24450);
nor U25314 (N_25314,N_24000,N_24497);
nor U25315 (N_25315,N_24134,N_24521);
or U25316 (N_25316,N_25188,N_24018);
xor U25317 (N_25317,N_24022,N_24902);
or U25318 (N_25318,N_24330,N_24447);
nand U25319 (N_25319,N_24490,N_24278);
nor U25320 (N_25320,N_24251,N_24464);
or U25321 (N_25321,N_25036,N_24169);
nand U25322 (N_25322,N_24166,N_24806);
nor U25323 (N_25323,N_24058,N_24425);
nor U25324 (N_25324,N_24884,N_25189);
and U25325 (N_25325,N_25173,N_24199);
or U25326 (N_25326,N_25142,N_24545);
or U25327 (N_25327,N_24747,N_25176);
nor U25328 (N_25328,N_24309,N_24928);
xnor U25329 (N_25329,N_24429,N_24320);
nand U25330 (N_25330,N_24062,N_24459);
or U25331 (N_25331,N_24687,N_25103);
and U25332 (N_25332,N_24361,N_24507);
and U25333 (N_25333,N_25086,N_24550);
or U25334 (N_25334,N_24200,N_24053);
nor U25335 (N_25335,N_24352,N_24987);
nor U25336 (N_25336,N_24347,N_24959);
nand U25337 (N_25337,N_24525,N_25161);
nor U25338 (N_25338,N_25070,N_24732);
nor U25339 (N_25339,N_24693,N_24602);
nor U25340 (N_25340,N_24547,N_24415);
and U25341 (N_25341,N_24880,N_24364);
or U25342 (N_25342,N_24996,N_24171);
or U25343 (N_25343,N_24963,N_25144);
nor U25344 (N_25344,N_25045,N_24074);
xnor U25345 (N_25345,N_25143,N_24700);
nand U25346 (N_25346,N_25184,N_24081);
nand U25347 (N_25347,N_25033,N_24697);
or U25348 (N_25348,N_24843,N_24213);
nor U25349 (N_25349,N_24438,N_24378);
or U25350 (N_25350,N_24841,N_24698);
or U25351 (N_25351,N_24472,N_24756);
or U25352 (N_25352,N_25041,N_24002);
nand U25353 (N_25353,N_24299,N_24871);
nor U25354 (N_25354,N_24945,N_24923);
nor U25355 (N_25355,N_24245,N_24094);
or U25356 (N_25356,N_24365,N_24660);
xor U25357 (N_25357,N_24160,N_24059);
nor U25358 (N_25358,N_24726,N_25039);
nand U25359 (N_25359,N_24976,N_24630);
nor U25360 (N_25360,N_24345,N_25116);
xnor U25361 (N_25361,N_24135,N_25122);
nor U25362 (N_25362,N_24253,N_24332);
nor U25363 (N_25363,N_24564,N_25044);
xnor U25364 (N_25364,N_24241,N_24095);
nand U25365 (N_25365,N_24748,N_24424);
or U25366 (N_25366,N_24397,N_24844);
nor U25367 (N_25367,N_24655,N_24055);
nor U25368 (N_25368,N_24285,N_24678);
and U25369 (N_25369,N_24215,N_24773);
xnor U25370 (N_25370,N_24966,N_24670);
nand U25371 (N_25371,N_24983,N_25026);
nor U25372 (N_25372,N_24875,N_24721);
and U25373 (N_25373,N_24457,N_24106);
and U25374 (N_25374,N_24724,N_25098);
nand U25375 (N_25375,N_24962,N_24076);
and U25376 (N_25376,N_24229,N_24740);
nand U25377 (N_25377,N_24758,N_24096);
nand U25378 (N_25378,N_24301,N_25187);
or U25379 (N_25379,N_25183,N_24395);
or U25380 (N_25380,N_24416,N_24368);
nand U25381 (N_25381,N_24657,N_24536);
and U25382 (N_25382,N_24648,N_24639);
xor U25383 (N_25383,N_24772,N_25028);
nor U25384 (N_25384,N_24308,N_24535);
xor U25385 (N_25385,N_24498,N_25119);
and U25386 (N_25386,N_24098,N_24154);
and U25387 (N_25387,N_24466,N_24662);
and U25388 (N_25388,N_24159,N_24725);
nor U25389 (N_25389,N_24072,N_24210);
xor U25390 (N_25390,N_24187,N_25007);
and U25391 (N_25391,N_24136,N_24194);
nor U25392 (N_25392,N_24865,N_24122);
and U25393 (N_25393,N_24888,N_24803);
and U25394 (N_25394,N_24799,N_24121);
and U25395 (N_25395,N_24297,N_24198);
nor U25396 (N_25396,N_24869,N_24842);
nand U25397 (N_25397,N_24656,N_25079);
and U25398 (N_25398,N_24409,N_24175);
nand U25399 (N_25399,N_24516,N_24776);
or U25400 (N_25400,N_25153,N_24917);
and U25401 (N_25401,N_24454,N_24054);
nor U25402 (N_25402,N_24673,N_24957);
and U25403 (N_25403,N_24465,N_24007);
nor U25404 (N_25404,N_24284,N_24252);
nor U25405 (N_25405,N_24480,N_24763);
xor U25406 (N_25406,N_24562,N_24470);
or U25407 (N_25407,N_24710,N_24954);
xnor U25408 (N_25408,N_25192,N_24783);
nor U25409 (N_25409,N_24050,N_24614);
nor U25410 (N_25410,N_24290,N_24811);
xnor U25411 (N_25411,N_24203,N_24247);
nand U25412 (N_25412,N_24162,N_25193);
and U25413 (N_25413,N_25151,N_25195);
xor U25414 (N_25414,N_25102,N_24546);
or U25415 (N_25415,N_24633,N_24569);
or U25416 (N_25416,N_24524,N_25020);
xor U25417 (N_25417,N_24127,N_24351);
nand U25418 (N_25418,N_25072,N_24563);
nand U25419 (N_25419,N_24688,N_24283);
and U25420 (N_25420,N_24254,N_24752);
nor U25421 (N_25421,N_25034,N_24366);
nand U25422 (N_25422,N_24383,N_24681);
and U25423 (N_25423,N_24271,N_24689);
and U25424 (N_25424,N_24218,N_24491);
or U25425 (N_25425,N_24272,N_24608);
xor U25426 (N_25426,N_24951,N_24565);
xor U25427 (N_25427,N_25074,N_24174);
or U25428 (N_25428,N_24446,N_24711);
nand U25429 (N_25429,N_24674,N_24866);
nor U25430 (N_25430,N_25179,N_24116);
nand U25431 (N_25431,N_24191,N_24543);
nor U25432 (N_25432,N_24823,N_24042);
or U25433 (N_25433,N_25059,N_24858);
nand U25434 (N_25434,N_24791,N_24423);
nor U25435 (N_25435,N_25101,N_24571);
nor U25436 (N_25436,N_24103,N_24690);
and U25437 (N_25437,N_25146,N_24304);
or U25438 (N_25438,N_24400,N_25171);
nand U25439 (N_25439,N_24281,N_24151);
and U25440 (N_25440,N_25134,N_24834);
nand U25441 (N_25441,N_25065,N_24067);
nand U25442 (N_25442,N_24997,N_24044);
xnor U25443 (N_25443,N_24282,N_24508);
nor U25444 (N_25444,N_24146,N_24988);
nand U25445 (N_25445,N_24077,N_24808);
nor U25446 (N_25446,N_24830,N_24286);
nand U25447 (N_25447,N_24770,N_24071);
nor U25448 (N_25448,N_24035,N_24335);
xor U25449 (N_25449,N_24955,N_24590);
or U25450 (N_25450,N_24864,N_24020);
xnor U25451 (N_25451,N_24616,N_25197);
xor U25452 (N_25452,N_24960,N_24321);
or U25453 (N_25453,N_24765,N_25175);
nand U25454 (N_25454,N_25160,N_24930);
or U25455 (N_25455,N_24645,N_24825);
and U25456 (N_25456,N_24736,N_24014);
nand U25457 (N_25457,N_24114,N_24576);
nor U25458 (N_25458,N_24837,N_24768);
and U25459 (N_25459,N_24914,N_25133);
xnor U25460 (N_25460,N_25148,N_24040);
or U25461 (N_25461,N_25076,N_25047);
or U25462 (N_25462,N_24691,N_25149);
xnor U25463 (N_25463,N_24513,N_24206);
nand U25464 (N_25464,N_25083,N_24685);
xor U25465 (N_25465,N_24755,N_24029);
and U25466 (N_25466,N_25164,N_25130);
nand U25467 (N_25467,N_24086,N_24860);
nor U25468 (N_25468,N_24651,N_25005);
and U25469 (N_25469,N_24801,N_24157);
nand U25470 (N_25470,N_25199,N_24158);
nor U25471 (N_25471,N_24439,N_25174);
xnor U25472 (N_25472,N_24111,N_24350);
and U25473 (N_25473,N_24057,N_24197);
nor U25474 (N_25474,N_24779,N_24984);
nand U25475 (N_25475,N_24394,N_24782);
nand U25476 (N_25476,N_24739,N_24956);
and U25477 (N_25477,N_24440,N_25012);
or U25478 (N_25478,N_24677,N_24373);
xnor U25479 (N_25479,N_24354,N_24181);
nor U25480 (N_25480,N_24167,N_24030);
xor U25481 (N_25481,N_24551,N_25056);
xor U25482 (N_25482,N_24207,N_24192);
nand U25483 (N_25483,N_24918,N_24117);
nor U25484 (N_25484,N_24622,N_24494);
and U25485 (N_25485,N_24743,N_24730);
and U25486 (N_25486,N_24150,N_24113);
or U25487 (N_25487,N_25030,N_25129);
nor U25488 (N_25488,N_24745,N_24038);
and U25489 (N_25489,N_24531,N_24371);
nand U25490 (N_25490,N_24515,N_25106);
nand U25491 (N_25491,N_24455,N_24056);
or U25492 (N_25492,N_24405,N_24561);
nand U25493 (N_25493,N_25120,N_24430);
nand U25494 (N_25494,N_25132,N_24147);
nand U25495 (N_25495,N_24817,N_24125);
nor U25496 (N_25496,N_24529,N_24617);
nor U25497 (N_25497,N_24891,N_25087);
nor U25498 (N_25498,N_24991,N_25027);
xor U25499 (N_25499,N_24468,N_24172);
nor U25500 (N_25500,N_24937,N_24195);
nand U25501 (N_25501,N_24144,N_25023);
and U25502 (N_25502,N_24872,N_24107);
or U25503 (N_25503,N_24883,N_24051);
or U25504 (N_25504,N_24595,N_25085);
xnor U25505 (N_25505,N_24790,N_24534);
nand U25506 (N_25506,N_24734,N_25190);
xnor U25507 (N_25507,N_24467,N_24183);
and U25508 (N_25508,N_24139,N_24810);
nand U25509 (N_25509,N_24999,N_24481);
xnor U25510 (N_25510,N_25121,N_25055);
nor U25511 (N_25511,N_24762,N_24759);
and U25512 (N_25512,N_24886,N_25017);
and U25513 (N_25513,N_24652,N_24684);
nor U25514 (N_25514,N_24093,N_24611);
nand U25515 (N_25515,N_24658,N_24636);
nand U25516 (N_25516,N_25068,N_24026);
nor U25517 (N_25517,N_24985,N_25107);
or U25518 (N_25518,N_24100,N_24737);
xnor U25519 (N_25519,N_24896,N_24148);
and U25520 (N_25520,N_24819,N_24403);
nand U25521 (N_25521,N_24266,N_24804);
and U25522 (N_25522,N_24893,N_24073);
and U25523 (N_25523,N_24444,N_24671);
nor U25524 (N_25524,N_25004,N_24577);
or U25525 (N_25525,N_24303,N_24623);
nor U25526 (N_25526,N_24391,N_24537);
and U25527 (N_25527,N_24637,N_24155);
or U25528 (N_25528,N_24046,N_25117);
nand U25529 (N_25529,N_24973,N_24031);
nand U25530 (N_25530,N_24702,N_24298);
xor U25531 (N_25531,N_24302,N_24433);
nor U25532 (N_25532,N_24442,N_24927);
nand U25533 (N_25533,N_24190,N_24965);
and U25534 (N_25534,N_24665,N_24082);
nand U25535 (N_25535,N_24993,N_24360);
nor U25536 (N_25536,N_24246,N_24944);
or U25537 (N_25537,N_24802,N_24108);
nor U25538 (N_25538,N_25097,N_24989);
or U25539 (N_25539,N_24746,N_24853);
nand U25540 (N_25540,N_24419,N_24717);
nor U25541 (N_25541,N_24520,N_24406);
xor U25542 (N_25542,N_24389,N_24428);
xnor U25543 (N_25543,N_24949,N_24824);
nor U25544 (N_25544,N_25186,N_25196);
xor U25545 (N_25545,N_24676,N_25110);
xor U25546 (N_25546,N_24349,N_24385);
and U25547 (N_25547,N_24004,N_24083);
nand U25548 (N_25548,N_25191,N_25078);
nand U25549 (N_25549,N_24542,N_24906);
nand U25550 (N_25550,N_25157,N_24242);
nand U25551 (N_25551,N_24331,N_24256);
nor U25552 (N_25552,N_25158,N_25111);
or U25553 (N_25553,N_24539,N_24008);
nor U25554 (N_25554,N_24862,N_25031);
nor U25555 (N_25555,N_24104,N_24527);
and U25556 (N_25556,N_25037,N_24212);
nand U25557 (N_25557,N_24476,N_24408);
xor U25558 (N_25558,N_24919,N_24407);
xnor U25559 (N_25559,N_24248,N_24712);
or U25560 (N_25560,N_24800,N_24895);
and U25561 (N_25561,N_24574,N_24632);
and U25562 (N_25562,N_24456,N_24892);
xnor U25563 (N_25563,N_24631,N_24793);
nor U25564 (N_25564,N_24557,N_24585);
and U25565 (N_25565,N_24478,N_24367);
xor U25566 (N_25566,N_25019,N_24796);
nand U25567 (N_25567,N_24975,N_24161);
or U25568 (N_25568,N_24063,N_25040);
nand U25569 (N_25569,N_24952,N_24572);
xnor U25570 (N_25570,N_24694,N_24971);
xor U25571 (N_25571,N_24221,N_25067);
or U25572 (N_25572,N_24735,N_25049);
nand U25573 (N_25573,N_25118,N_24511);
nand U25574 (N_25574,N_24451,N_24701);
and U25575 (N_25575,N_24530,N_24043);
xnor U25576 (N_25576,N_24469,N_24822);
nand U25577 (N_25577,N_24483,N_24578);
xor U25578 (N_25578,N_24915,N_24909);
xnor U25579 (N_25579,N_24168,N_24499);
or U25580 (N_25580,N_25029,N_24232);
and U25581 (N_25581,N_24066,N_24133);
nor U25582 (N_25582,N_24669,N_25135);
or U25583 (N_25583,N_24010,N_24931);
nor U25584 (N_25584,N_24719,N_24850);
or U25585 (N_25585,N_24900,N_25008);
or U25586 (N_25586,N_24238,N_25181);
and U25587 (N_25587,N_25136,N_25022);
xor U25588 (N_25588,N_24270,N_25141);
nor U25589 (N_25589,N_24540,N_24329);
xnor U25590 (N_25590,N_24774,N_24432);
and U25591 (N_25591,N_24598,N_24584);
and U25592 (N_25592,N_25156,N_24475);
and U25593 (N_25593,N_24722,N_24061);
nand U25594 (N_25594,N_25115,N_24589);
nor U25595 (N_25595,N_24493,N_24761);
or U25596 (N_25596,N_24680,N_25006);
or U25597 (N_25597,N_24390,N_24084);
nor U25598 (N_25598,N_24346,N_24663);
nor U25599 (N_25599,N_24929,N_24411);
and U25600 (N_25600,N_24392,N_24305);
or U25601 (N_25601,N_24274,N_24940);
or U25602 (N_25602,N_24859,N_25096);
xnor U25603 (N_25603,N_25088,N_24333);
and U25604 (N_25604,N_24234,N_24489);
and U25605 (N_25605,N_24553,N_24357);
and U25606 (N_25606,N_24223,N_24560);
xor U25607 (N_25607,N_24129,N_24548);
nand U25608 (N_25608,N_24749,N_24137);
and U25609 (N_25609,N_25002,N_24556);
nand U25610 (N_25610,N_24412,N_24048);
and U25611 (N_25611,N_24836,N_24006);
nand U25612 (N_25612,N_24421,N_24964);
nand U25613 (N_25613,N_24580,N_24599);
nand U25614 (N_25614,N_25123,N_24064);
nand U25615 (N_25615,N_24816,N_24130);
nand U25616 (N_25616,N_25152,N_24313);
nand U25617 (N_25617,N_24292,N_24359);
or U25618 (N_25618,N_24339,N_24532);
or U25619 (N_25619,N_24001,N_24713);
nor U25620 (N_25620,N_24894,N_24821);
xor U25621 (N_25621,N_24170,N_25091);
nor U25622 (N_25622,N_24065,N_24435);
xnor U25623 (N_25623,N_24380,N_24620);
and U25624 (N_25624,N_24193,N_24953);
nand U25625 (N_25625,N_24566,N_24696);
nand U25626 (N_25626,N_25077,N_24088);
or U25627 (N_25627,N_24204,N_24510);
xnor U25628 (N_25628,N_24099,N_24826);
or U25629 (N_25629,N_24705,N_24437);
or U25630 (N_25630,N_24922,N_24642);
xnor U25631 (N_25631,N_24805,N_24443);
nor U25632 (N_25632,N_24244,N_24079);
nand U25633 (N_25633,N_24013,N_25043);
or U25634 (N_25634,N_24504,N_24727);
xnor U25635 (N_25635,N_24609,N_24754);
and U25636 (N_25636,N_24907,N_25167);
nand U25637 (N_25637,N_25169,N_25062);
xnor U25638 (N_25638,N_25015,N_24101);
and U25639 (N_25639,N_24692,N_24024);
and U25640 (N_25640,N_24145,N_24182);
or U25641 (N_25641,N_24523,N_25194);
or U25642 (N_25642,N_24668,N_24399);
and U25643 (N_25643,N_24979,N_24686);
or U25644 (N_25644,N_24268,N_24091);
or U25645 (N_25645,N_24120,N_24666);
nand U25646 (N_25646,N_25060,N_24878);
nor U25647 (N_25647,N_24179,N_25046);
xnor U25648 (N_25648,N_24025,N_24621);
or U25649 (N_25649,N_24741,N_24227);
and U25650 (N_25650,N_24829,N_24300);
xnor U25651 (N_25651,N_24913,N_24362);
or U25652 (N_25652,N_24231,N_24683);
xnor U25653 (N_25653,N_24477,N_24961);
nand U25654 (N_25654,N_24920,N_25140);
nand U25655 (N_25655,N_25165,N_24047);
nor U25656 (N_25656,N_24306,N_24764);
nand U25657 (N_25657,N_25126,N_24977);
nor U25658 (N_25658,N_24558,N_24992);
xor U25659 (N_25659,N_24846,N_24760);
nor U25660 (N_25660,N_24924,N_24414);
nor U25661 (N_25661,N_24372,N_24463);
or U25662 (N_25662,N_24124,N_24597);
nor U25663 (N_25663,N_25138,N_24287);
or U25664 (N_25664,N_24280,N_24180);
nand U25665 (N_25665,N_24827,N_24296);
and U25666 (N_25666,N_24936,N_24591);
nor U25667 (N_25667,N_24970,N_24857);
and U25668 (N_25668,N_24123,N_24533);
nand U25669 (N_25669,N_24852,N_25024);
xnor U25670 (N_25670,N_24593,N_24009);
nand U25671 (N_25671,N_24236,N_24369);
xor U25672 (N_25672,N_25057,N_24239);
and U25673 (N_25673,N_25073,N_24176);
and U25674 (N_25674,N_24706,N_24032);
or U25675 (N_25675,N_24382,N_24613);
nor U25676 (N_25676,N_24643,N_24328);
xor U25677 (N_25677,N_24851,N_24379);
and U25678 (N_25678,N_24012,N_24388);
nor U25679 (N_25679,N_24528,N_24903);
or U25680 (N_25680,N_24277,N_24707);
nor U25681 (N_25681,N_24318,N_24626);
nor U25682 (N_25682,N_25198,N_24039);
nand U25683 (N_25683,N_24634,N_24870);
and U25684 (N_25684,N_24036,N_24628);
and U25685 (N_25685,N_24948,N_24295);
nor U25686 (N_25686,N_24818,N_24115);
and U25687 (N_25687,N_25003,N_25053);
or U25688 (N_25688,N_24041,N_25093);
nand U25689 (N_25689,N_24679,N_24460);
nand U25690 (N_25690,N_24552,N_24667);
xor U25691 (N_25691,N_24925,N_25084);
nor U25692 (N_25692,N_24807,N_25094);
and U25693 (N_25693,N_24156,N_24188);
or U25694 (N_25694,N_24312,N_24128);
nor U25695 (N_25695,N_25069,N_24186);
or U25696 (N_25696,N_24938,N_24738);
nand U25697 (N_25697,N_24612,N_24600);
or U25698 (N_25698,N_24943,N_24744);
or U25699 (N_25699,N_24356,N_24629);
nor U25700 (N_25700,N_24506,N_24695);
nor U25701 (N_25701,N_24222,N_24855);
or U25702 (N_25702,N_24797,N_24263);
xnor U25703 (N_25703,N_24974,N_24887);
xnor U25704 (N_25704,N_24209,N_24845);
nand U25705 (N_25705,N_24921,N_25014);
or U25706 (N_25706,N_24788,N_25013);
nor U25707 (N_25707,N_24023,N_24291);
and U25708 (N_25708,N_24021,N_24434);
or U25709 (N_25709,N_25009,N_24340);
nor U25710 (N_25710,N_24492,N_24750);
nor U25711 (N_25711,N_25185,N_24998);
xor U25712 (N_25712,N_24838,N_24833);
and U25713 (N_25713,N_24495,N_24005);
nand U25714 (N_25714,N_24995,N_24715);
nand U25715 (N_25715,N_24353,N_24404);
nor U25716 (N_25716,N_24916,N_24220);
nand U25717 (N_25717,N_24216,N_24293);
xor U25718 (N_25718,N_24820,N_24541);
nor U25719 (N_25719,N_24723,N_24596);
nor U25720 (N_25720,N_24033,N_25154);
nor U25721 (N_25721,N_24474,N_25150);
and U25722 (N_25722,N_24334,N_24131);
nand U25723 (N_25723,N_24027,N_25038);
and U25724 (N_25724,N_24034,N_25051);
or U25725 (N_25725,N_24586,N_24376);
or U25726 (N_25726,N_25035,N_24259);
nand U25727 (N_25727,N_24848,N_25082);
xnor U25728 (N_25728,N_25128,N_24863);
xnor U25729 (N_25729,N_24461,N_24787);
and U25730 (N_25730,N_24016,N_24402);
nor U25731 (N_25731,N_24488,N_24342);
and U25732 (N_25732,N_24417,N_24089);
nor U25733 (N_25733,N_24453,N_24396);
xnor U25734 (N_25734,N_24486,N_25048);
nor U25735 (N_25735,N_24625,N_24647);
nor U25736 (N_25736,N_24387,N_24579);
xnor U25737 (N_25737,N_24410,N_24849);
nand U25738 (N_25738,N_24785,N_24250);
xor U25739 (N_25739,N_24237,N_24594);
or U25740 (N_25740,N_24986,N_24163);
xor U25741 (N_25741,N_24226,N_24911);
nor U25742 (N_25742,N_25063,N_24728);
and U25743 (N_25743,N_24068,N_24559);
or U25744 (N_25744,N_24431,N_24449);
xor U25745 (N_25745,N_24219,N_24484);
nand U25746 (N_25746,N_24045,N_24784);
nand U25747 (N_25747,N_25182,N_24640);
nor U25748 (N_25748,N_24771,N_24505);
and U25749 (N_25749,N_24798,N_24877);
or U25750 (N_25750,N_25052,N_24840);
or U25751 (N_25751,N_24078,N_24294);
nand U25752 (N_25752,N_24573,N_24132);
and U25753 (N_25753,N_25131,N_25090);
and U25754 (N_25754,N_24496,N_24941);
and U25755 (N_25755,N_24733,N_24441);
or U25756 (N_25756,N_24087,N_24969);
nand U25757 (N_25757,N_24264,N_24377);
or U25758 (N_25758,N_25177,N_24890);
and U25759 (N_25759,N_24661,N_24778);
xor U25760 (N_25760,N_24386,N_25066);
and U25761 (N_25761,N_24751,N_24809);
nor U25762 (N_25762,N_24767,N_25180);
or U25763 (N_25763,N_25050,N_24885);
and U25764 (N_25764,N_24624,N_24275);
nor U25765 (N_25765,N_24426,N_24605);
and U25766 (N_25766,N_24487,N_24458);
nor U25767 (N_25767,N_24420,N_24436);
nor U25768 (N_25768,N_24682,N_24348);
or U25769 (N_25769,N_24538,N_24501);
xor U25770 (N_25770,N_24258,N_24323);
xor U25771 (N_25771,N_24240,N_24854);
and U25772 (N_25772,N_25125,N_24152);
xnor U25773 (N_25773,N_24070,N_24581);
nor U25774 (N_25774,N_25018,N_24185);
and U25775 (N_25775,N_24049,N_24583);
nand U25776 (N_25776,N_24653,N_24355);
and U25777 (N_25777,N_25025,N_24509);
xor U25778 (N_25778,N_24792,N_24742);
nand U25779 (N_25779,N_24926,N_24709);
nand U25780 (N_25780,N_24381,N_24196);
nand U25781 (N_25781,N_25058,N_24052);
nand U25782 (N_25782,N_24518,N_24184);
xnor U25783 (N_25783,N_24028,N_24143);
xor U25784 (N_25784,N_24110,N_24202);
nor U25785 (N_25785,N_24149,N_24729);
xnor U25786 (N_25786,N_24338,N_24445);
nor U25787 (N_25787,N_24011,N_24112);
xnor U25788 (N_25788,N_24794,N_25099);
nand U25789 (N_25789,N_24273,N_24603);
nor U25790 (N_25790,N_24384,N_24257);
nor U25791 (N_25791,N_24267,N_25105);
or U25792 (N_25792,N_24831,N_24279);
nand U25793 (N_25793,N_24619,N_24322);
nand U25794 (N_25794,N_24592,N_24075);
nand U25795 (N_25795,N_25064,N_24502);
and U25796 (N_25796,N_24178,N_24777);
and U25797 (N_25797,N_25016,N_24757);
and U25798 (N_25798,N_24165,N_24017);
nor U25799 (N_25799,N_24118,N_24567);
nand U25800 (N_25800,N_24928,N_24291);
or U25801 (N_25801,N_24905,N_24432);
nor U25802 (N_25802,N_24688,N_24605);
xor U25803 (N_25803,N_24784,N_24111);
nor U25804 (N_25804,N_24366,N_25189);
nand U25805 (N_25805,N_24592,N_24071);
nor U25806 (N_25806,N_24514,N_24495);
xor U25807 (N_25807,N_24970,N_24876);
or U25808 (N_25808,N_24890,N_24489);
xor U25809 (N_25809,N_24201,N_24578);
nor U25810 (N_25810,N_24408,N_24902);
nor U25811 (N_25811,N_24697,N_24391);
xnor U25812 (N_25812,N_24255,N_25068);
or U25813 (N_25813,N_24158,N_24586);
nand U25814 (N_25814,N_24526,N_24172);
nand U25815 (N_25815,N_24052,N_24527);
and U25816 (N_25816,N_24225,N_24782);
or U25817 (N_25817,N_24061,N_24591);
or U25818 (N_25818,N_24492,N_24412);
or U25819 (N_25819,N_24440,N_24192);
xor U25820 (N_25820,N_25108,N_24677);
nand U25821 (N_25821,N_24559,N_24011);
and U25822 (N_25822,N_25109,N_24557);
nor U25823 (N_25823,N_25048,N_25083);
nand U25824 (N_25824,N_24163,N_24743);
xor U25825 (N_25825,N_25059,N_24591);
and U25826 (N_25826,N_24637,N_24069);
nor U25827 (N_25827,N_24522,N_25035);
nand U25828 (N_25828,N_24079,N_24013);
or U25829 (N_25829,N_24077,N_24356);
xor U25830 (N_25830,N_24930,N_25101);
and U25831 (N_25831,N_24356,N_24522);
nand U25832 (N_25832,N_24395,N_24547);
nor U25833 (N_25833,N_25122,N_24702);
xnor U25834 (N_25834,N_24521,N_24320);
nor U25835 (N_25835,N_25131,N_24358);
and U25836 (N_25836,N_25144,N_24934);
nand U25837 (N_25837,N_24931,N_24909);
and U25838 (N_25838,N_24095,N_24773);
and U25839 (N_25839,N_24905,N_24666);
or U25840 (N_25840,N_24085,N_24690);
or U25841 (N_25841,N_24849,N_24942);
or U25842 (N_25842,N_24199,N_24622);
xnor U25843 (N_25843,N_25099,N_24815);
xor U25844 (N_25844,N_25141,N_24673);
or U25845 (N_25845,N_24143,N_24487);
or U25846 (N_25846,N_24875,N_24720);
and U25847 (N_25847,N_24209,N_24027);
or U25848 (N_25848,N_25030,N_24078);
or U25849 (N_25849,N_24095,N_24247);
nand U25850 (N_25850,N_24772,N_24887);
nand U25851 (N_25851,N_24363,N_25168);
and U25852 (N_25852,N_25193,N_24492);
or U25853 (N_25853,N_24836,N_24096);
nor U25854 (N_25854,N_25180,N_24309);
or U25855 (N_25855,N_24509,N_24521);
nand U25856 (N_25856,N_24145,N_24506);
or U25857 (N_25857,N_24934,N_24650);
nor U25858 (N_25858,N_24376,N_24050);
xnor U25859 (N_25859,N_24721,N_24281);
xor U25860 (N_25860,N_24734,N_24578);
or U25861 (N_25861,N_25112,N_24178);
nor U25862 (N_25862,N_25023,N_24050);
and U25863 (N_25863,N_24011,N_25193);
nand U25864 (N_25864,N_24319,N_24980);
or U25865 (N_25865,N_24493,N_24898);
or U25866 (N_25866,N_24114,N_24462);
nor U25867 (N_25867,N_24192,N_25066);
and U25868 (N_25868,N_24616,N_24839);
or U25869 (N_25869,N_24021,N_24499);
xor U25870 (N_25870,N_25129,N_25115);
nor U25871 (N_25871,N_25065,N_24378);
and U25872 (N_25872,N_24136,N_24345);
nor U25873 (N_25873,N_24642,N_24322);
nand U25874 (N_25874,N_24291,N_24139);
or U25875 (N_25875,N_24969,N_24612);
nor U25876 (N_25876,N_24949,N_24757);
nand U25877 (N_25877,N_24328,N_24423);
nor U25878 (N_25878,N_24872,N_24861);
nand U25879 (N_25879,N_24335,N_24846);
xnor U25880 (N_25880,N_25155,N_24503);
or U25881 (N_25881,N_24323,N_24400);
and U25882 (N_25882,N_24393,N_25183);
xnor U25883 (N_25883,N_24762,N_25162);
nand U25884 (N_25884,N_25040,N_24570);
or U25885 (N_25885,N_25178,N_25159);
or U25886 (N_25886,N_24027,N_24341);
nor U25887 (N_25887,N_24522,N_24181);
and U25888 (N_25888,N_24589,N_24999);
or U25889 (N_25889,N_24422,N_25067);
nor U25890 (N_25890,N_24351,N_24852);
or U25891 (N_25891,N_24620,N_25010);
xor U25892 (N_25892,N_25048,N_24570);
nand U25893 (N_25893,N_24265,N_24456);
and U25894 (N_25894,N_24138,N_25163);
nor U25895 (N_25895,N_24961,N_24698);
and U25896 (N_25896,N_24875,N_24249);
nor U25897 (N_25897,N_24312,N_24110);
nand U25898 (N_25898,N_24518,N_24953);
nand U25899 (N_25899,N_24752,N_24389);
or U25900 (N_25900,N_24021,N_24222);
nor U25901 (N_25901,N_25143,N_25145);
or U25902 (N_25902,N_24063,N_24995);
xor U25903 (N_25903,N_24888,N_25114);
nand U25904 (N_25904,N_24189,N_25096);
or U25905 (N_25905,N_25090,N_24425);
nand U25906 (N_25906,N_24955,N_24073);
nor U25907 (N_25907,N_24507,N_24885);
or U25908 (N_25908,N_24274,N_24770);
xor U25909 (N_25909,N_24487,N_24280);
or U25910 (N_25910,N_25055,N_24740);
and U25911 (N_25911,N_25137,N_24939);
or U25912 (N_25912,N_24717,N_24957);
or U25913 (N_25913,N_24263,N_25057);
xor U25914 (N_25914,N_24884,N_24699);
or U25915 (N_25915,N_25002,N_24359);
nand U25916 (N_25916,N_24311,N_24697);
nand U25917 (N_25917,N_24776,N_24613);
or U25918 (N_25918,N_24217,N_24097);
and U25919 (N_25919,N_24306,N_24257);
nand U25920 (N_25920,N_24736,N_24206);
and U25921 (N_25921,N_25067,N_24674);
and U25922 (N_25922,N_24890,N_24385);
or U25923 (N_25923,N_24873,N_24588);
and U25924 (N_25924,N_24696,N_24512);
nand U25925 (N_25925,N_24898,N_24439);
xor U25926 (N_25926,N_24832,N_24267);
xor U25927 (N_25927,N_24016,N_25131);
and U25928 (N_25928,N_24316,N_24959);
nand U25929 (N_25929,N_24782,N_24857);
xnor U25930 (N_25930,N_24580,N_24115);
nor U25931 (N_25931,N_25189,N_24052);
and U25932 (N_25932,N_24350,N_24001);
nand U25933 (N_25933,N_24929,N_24074);
nor U25934 (N_25934,N_24678,N_24650);
nand U25935 (N_25935,N_24058,N_24895);
and U25936 (N_25936,N_24224,N_24533);
and U25937 (N_25937,N_24395,N_24102);
nor U25938 (N_25938,N_24143,N_24518);
xor U25939 (N_25939,N_24017,N_24708);
xnor U25940 (N_25940,N_24592,N_24001);
xor U25941 (N_25941,N_24636,N_24441);
or U25942 (N_25942,N_25101,N_24083);
and U25943 (N_25943,N_24081,N_24594);
or U25944 (N_25944,N_25012,N_24398);
nand U25945 (N_25945,N_24595,N_25122);
xnor U25946 (N_25946,N_24643,N_25185);
and U25947 (N_25947,N_24969,N_24347);
xnor U25948 (N_25948,N_25185,N_24767);
nand U25949 (N_25949,N_24014,N_24792);
nor U25950 (N_25950,N_24661,N_24377);
and U25951 (N_25951,N_24578,N_24008);
nand U25952 (N_25952,N_25024,N_24446);
or U25953 (N_25953,N_24178,N_24419);
nand U25954 (N_25954,N_24776,N_25191);
and U25955 (N_25955,N_24151,N_24906);
and U25956 (N_25956,N_24563,N_24063);
xnor U25957 (N_25957,N_25009,N_24299);
or U25958 (N_25958,N_24814,N_24512);
nor U25959 (N_25959,N_24914,N_24587);
xor U25960 (N_25960,N_25025,N_25017);
and U25961 (N_25961,N_24259,N_24992);
nor U25962 (N_25962,N_25118,N_24667);
and U25963 (N_25963,N_24969,N_25148);
and U25964 (N_25964,N_24097,N_25126);
nand U25965 (N_25965,N_24593,N_24372);
xnor U25966 (N_25966,N_24478,N_24754);
nand U25967 (N_25967,N_24725,N_24074);
nand U25968 (N_25968,N_24229,N_25012);
xnor U25969 (N_25969,N_24829,N_25024);
and U25970 (N_25970,N_24753,N_24053);
or U25971 (N_25971,N_25195,N_24727);
nand U25972 (N_25972,N_24228,N_24253);
or U25973 (N_25973,N_24572,N_25178);
nor U25974 (N_25974,N_24214,N_25170);
nor U25975 (N_25975,N_24079,N_24266);
nor U25976 (N_25976,N_24452,N_24307);
and U25977 (N_25977,N_24700,N_24778);
xnor U25978 (N_25978,N_24105,N_24981);
xnor U25979 (N_25979,N_24816,N_24877);
xnor U25980 (N_25980,N_24468,N_25098);
nand U25981 (N_25981,N_24663,N_24231);
nor U25982 (N_25982,N_24039,N_25159);
nor U25983 (N_25983,N_24637,N_24869);
nor U25984 (N_25984,N_24678,N_24667);
and U25985 (N_25985,N_24910,N_24738);
or U25986 (N_25986,N_24845,N_24814);
nand U25987 (N_25987,N_24847,N_24115);
or U25988 (N_25988,N_24423,N_24501);
xor U25989 (N_25989,N_24262,N_24568);
nor U25990 (N_25990,N_24254,N_24326);
and U25991 (N_25991,N_25157,N_24165);
xor U25992 (N_25992,N_25038,N_24051);
nor U25993 (N_25993,N_24563,N_24723);
or U25994 (N_25994,N_24381,N_24368);
nor U25995 (N_25995,N_24327,N_24869);
nor U25996 (N_25996,N_24172,N_25020);
and U25997 (N_25997,N_24538,N_24143);
nor U25998 (N_25998,N_24383,N_25077);
and U25999 (N_25999,N_24585,N_24236);
nand U26000 (N_26000,N_24450,N_24668);
xor U26001 (N_26001,N_24683,N_24587);
nor U26002 (N_26002,N_24583,N_24447);
nand U26003 (N_26003,N_24513,N_24691);
nor U26004 (N_26004,N_25182,N_24290);
nor U26005 (N_26005,N_24649,N_24682);
or U26006 (N_26006,N_24353,N_24615);
or U26007 (N_26007,N_24034,N_24784);
and U26008 (N_26008,N_24996,N_25190);
nor U26009 (N_26009,N_25012,N_24561);
xor U26010 (N_26010,N_24180,N_24944);
and U26011 (N_26011,N_24318,N_24110);
nor U26012 (N_26012,N_24131,N_24124);
xor U26013 (N_26013,N_24100,N_24885);
or U26014 (N_26014,N_24976,N_24653);
nor U26015 (N_26015,N_24950,N_24973);
or U26016 (N_26016,N_24605,N_24621);
and U26017 (N_26017,N_24493,N_24381);
or U26018 (N_26018,N_24411,N_24136);
and U26019 (N_26019,N_24455,N_24871);
nor U26020 (N_26020,N_24368,N_24297);
xnor U26021 (N_26021,N_24724,N_24211);
or U26022 (N_26022,N_25128,N_24924);
xnor U26023 (N_26023,N_24997,N_24458);
and U26024 (N_26024,N_25191,N_24033);
nand U26025 (N_26025,N_24424,N_24619);
nand U26026 (N_26026,N_25149,N_25190);
or U26027 (N_26027,N_24834,N_24672);
and U26028 (N_26028,N_24076,N_24250);
or U26029 (N_26029,N_24968,N_24386);
nor U26030 (N_26030,N_24950,N_24117);
or U26031 (N_26031,N_24585,N_24587);
nand U26032 (N_26032,N_24580,N_24878);
or U26033 (N_26033,N_24049,N_25083);
xor U26034 (N_26034,N_24530,N_25015);
xnor U26035 (N_26035,N_24994,N_24372);
and U26036 (N_26036,N_24789,N_24477);
nor U26037 (N_26037,N_24365,N_24655);
or U26038 (N_26038,N_25112,N_24402);
xnor U26039 (N_26039,N_24192,N_24987);
and U26040 (N_26040,N_24335,N_25146);
nand U26041 (N_26041,N_24668,N_24051);
and U26042 (N_26042,N_24709,N_24573);
nor U26043 (N_26043,N_24098,N_24959);
or U26044 (N_26044,N_24568,N_24336);
or U26045 (N_26045,N_24485,N_25102);
nand U26046 (N_26046,N_25166,N_24461);
or U26047 (N_26047,N_24941,N_24009);
and U26048 (N_26048,N_24532,N_24211);
nand U26049 (N_26049,N_24980,N_24380);
and U26050 (N_26050,N_25036,N_25017);
and U26051 (N_26051,N_24636,N_25035);
nand U26052 (N_26052,N_24410,N_24736);
and U26053 (N_26053,N_24798,N_24794);
nor U26054 (N_26054,N_24571,N_25190);
nand U26055 (N_26055,N_25011,N_24716);
nand U26056 (N_26056,N_24957,N_24603);
and U26057 (N_26057,N_25069,N_24175);
and U26058 (N_26058,N_24664,N_24380);
xnor U26059 (N_26059,N_24633,N_24533);
nand U26060 (N_26060,N_25151,N_24194);
xor U26061 (N_26061,N_24693,N_24608);
or U26062 (N_26062,N_24776,N_24358);
and U26063 (N_26063,N_24505,N_24065);
nor U26064 (N_26064,N_25106,N_24150);
xnor U26065 (N_26065,N_25100,N_24485);
or U26066 (N_26066,N_24972,N_24107);
and U26067 (N_26067,N_24104,N_24000);
nand U26068 (N_26068,N_24547,N_25140);
nor U26069 (N_26069,N_24678,N_24996);
nand U26070 (N_26070,N_24645,N_25012);
and U26071 (N_26071,N_24366,N_24086);
or U26072 (N_26072,N_25077,N_24869);
xnor U26073 (N_26073,N_24819,N_24691);
and U26074 (N_26074,N_24571,N_24780);
and U26075 (N_26075,N_24611,N_24257);
nand U26076 (N_26076,N_25012,N_25006);
nor U26077 (N_26077,N_24310,N_24359);
xnor U26078 (N_26078,N_24111,N_24462);
and U26079 (N_26079,N_25004,N_24225);
or U26080 (N_26080,N_24455,N_24075);
nand U26081 (N_26081,N_24166,N_24769);
or U26082 (N_26082,N_24510,N_24418);
and U26083 (N_26083,N_24155,N_24383);
nand U26084 (N_26084,N_24650,N_24470);
nand U26085 (N_26085,N_25061,N_25161);
nand U26086 (N_26086,N_24846,N_24962);
or U26087 (N_26087,N_24509,N_24485);
nor U26088 (N_26088,N_24925,N_24698);
and U26089 (N_26089,N_24056,N_24121);
nand U26090 (N_26090,N_24787,N_24464);
nand U26091 (N_26091,N_24432,N_24941);
xnor U26092 (N_26092,N_24454,N_24882);
or U26093 (N_26093,N_24071,N_24571);
nand U26094 (N_26094,N_24325,N_25178);
nor U26095 (N_26095,N_25132,N_24845);
nor U26096 (N_26096,N_25183,N_24815);
and U26097 (N_26097,N_24414,N_24267);
xnor U26098 (N_26098,N_24645,N_24387);
and U26099 (N_26099,N_24042,N_24760);
and U26100 (N_26100,N_24824,N_24554);
nor U26101 (N_26101,N_24616,N_24426);
xor U26102 (N_26102,N_24816,N_24870);
nand U26103 (N_26103,N_24164,N_24065);
xor U26104 (N_26104,N_24138,N_24711);
nand U26105 (N_26105,N_24871,N_24236);
nor U26106 (N_26106,N_24558,N_24505);
nand U26107 (N_26107,N_24079,N_24576);
nand U26108 (N_26108,N_24318,N_24002);
nor U26109 (N_26109,N_24110,N_24556);
xor U26110 (N_26110,N_24436,N_24337);
and U26111 (N_26111,N_24766,N_24562);
nand U26112 (N_26112,N_25068,N_25017);
xnor U26113 (N_26113,N_24225,N_24978);
nor U26114 (N_26114,N_24517,N_24008);
xnor U26115 (N_26115,N_24482,N_24307);
and U26116 (N_26116,N_24759,N_25108);
nor U26117 (N_26117,N_24919,N_24703);
nor U26118 (N_26118,N_24881,N_24268);
and U26119 (N_26119,N_24714,N_24892);
and U26120 (N_26120,N_24658,N_24568);
and U26121 (N_26121,N_25055,N_24408);
xor U26122 (N_26122,N_24448,N_25126);
and U26123 (N_26123,N_24660,N_25153);
or U26124 (N_26124,N_24078,N_24359);
nor U26125 (N_26125,N_24627,N_25077);
or U26126 (N_26126,N_25066,N_24577);
nand U26127 (N_26127,N_24844,N_24459);
nand U26128 (N_26128,N_24301,N_24485);
nor U26129 (N_26129,N_24277,N_24788);
and U26130 (N_26130,N_24456,N_25034);
xnor U26131 (N_26131,N_24787,N_24693);
or U26132 (N_26132,N_24598,N_24097);
nand U26133 (N_26133,N_24068,N_24621);
and U26134 (N_26134,N_24145,N_24071);
nand U26135 (N_26135,N_24704,N_24919);
or U26136 (N_26136,N_25183,N_24237);
nand U26137 (N_26137,N_24930,N_25128);
nor U26138 (N_26138,N_24256,N_24617);
and U26139 (N_26139,N_24823,N_24664);
xnor U26140 (N_26140,N_24197,N_24995);
or U26141 (N_26141,N_24114,N_24067);
nand U26142 (N_26142,N_24474,N_24599);
or U26143 (N_26143,N_24952,N_24561);
nor U26144 (N_26144,N_24002,N_24782);
or U26145 (N_26145,N_24486,N_24073);
and U26146 (N_26146,N_24397,N_24394);
xor U26147 (N_26147,N_24002,N_25020);
nor U26148 (N_26148,N_25046,N_24705);
or U26149 (N_26149,N_24534,N_24059);
xor U26150 (N_26150,N_24695,N_25108);
nor U26151 (N_26151,N_24232,N_24041);
nand U26152 (N_26152,N_24156,N_24997);
and U26153 (N_26153,N_24464,N_24344);
nor U26154 (N_26154,N_25006,N_24108);
nor U26155 (N_26155,N_24688,N_24596);
or U26156 (N_26156,N_24337,N_24241);
xor U26157 (N_26157,N_24633,N_24976);
nand U26158 (N_26158,N_24533,N_24928);
and U26159 (N_26159,N_24770,N_25079);
nand U26160 (N_26160,N_24461,N_24922);
and U26161 (N_26161,N_25110,N_24521);
xor U26162 (N_26162,N_25083,N_24908);
or U26163 (N_26163,N_24468,N_24605);
and U26164 (N_26164,N_24235,N_24669);
or U26165 (N_26165,N_24220,N_24677);
nor U26166 (N_26166,N_24129,N_24403);
nand U26167 (N_26167,N_25102,N_25165);
or U26168 (N_26168,N_24943,N_24551);
nand U26169 (N_26169,N_24619,N_24764);
nand U26170 (N_26170,N_24576,N_24496);
or U26171 (N_26171,N_24990,N_24216);
nor U26172 (N_26172,N_25175,N_25083);
xnor U26173 (N_26173,N_25136,N_24721);
and U26174 (N_26174,N_24678,N_24694);
or U26175 (N_26175,N_24167,N_24152);
and U26176 (N_26176,N_24196,N_25167);
nor U26177 (N_26177,N_24280,N_24221);
or U26178 (N_26178,N_24794,N_24806);
xnor U26179 (N_26179,N_24044,N_25189);
nor U26180 (N_26180,N_24351,N_24976);
nand U26181 (N_26181,N_24337,N_24675);
nor U26182 (N_26182,N_24280,N_24633);
and U26183 (N_26183,N_25187,N_25057);
xor U26184 (N_26184,N_24244,N_24699);
and U26185 (N_26185,N_24112,N_24612);
and U26186 (N_26186,N_24897,N_24658);
and U26187 (N_26187,N_24932,N_24407);
or U26188 (N_26188,N_24579,N_24282);
xor U26189 (N_26189,N_24115,N_24973);
and U26190 (N_26190,N_24189,N_24367);
xor U26191 (N_26191,N_24437,N_24681);
nand U26192 (N_26192,N_24718,N_24978);
and U26193 (N_26193,N_24263,N_24568);
nor U26194 (N_26194,N_24064,N_24004);
nor U26195 (N_26195,N_24171,N_24636);
or U26196 (N_26196,N_25164,N_24353);
and U26197 (N_26197,N_24383,N_24126);
or U26198 (N_26198,N_24708,N_24565);
nand U26199 (N_26199,N_24178,N_24745);
and U26200 (N_26200,N_24961,N_25162);
or U26201 (N_26201,N_24095,N_24045);
nor U26202 (N_26202,N_24991,N_24046);
nand U26203 (N_26203,N_25006,N_24702);
and U26204 (N_26204,N_24309,N_24193);
nor U26205 (N_26205,N_24240,N_24205);
nor U26206 (N_26206,N_24333,N_24899);
and U26207 (N_26207,N_24630,N_24757);
nand U26208 (N_26208,N_24021,N_25051);
and U26209 (N_26209,N_24413,N_24595);
or U26210 (N_26210,N_24249,N_24368);
or U26211 (N_26211,N_24400,N_25050);
xor U26212 (N_26212,N_24023,N_25050);
xor U26213 (N_26213,N_24312,N_24656);
or U26214 (N_26214,N_24368,N_25070);
or U26215 (N_26215,N_24645,N_25072);
nor U26216 (N_26216,N_24824,N_24079);
nand U26217 (N_26217,N_24279,N_25101);
and U26218 (N_26218,N_24827,N_25127);
xnor U26219 (N_26219,N_24894,N_24028);
xnor U26220 (N_26220,N_24471,N_25007);
or U26221 (N_26221,N_24906,N_25190);
nor U26222 (N_26222,N_24636,N_24867);
or U26223 (N_26223,N_24818,N_25128);
nand U26224 (N_26224,N_24316,N_24667);
nand U26225 (N_26225,N_24488,N_24766);
or U26226 (N_26226,N_24365,N_24720);
nor U26227 (N_26227,N_24158,N_24439);
nor U26228 (N_26228,N_24350,N_24331);
or U26229 (N_26229,N_24809,N_25150);
nor U26230 (N_26230,N_24164,N_24892);
nand U26231 (N_26231,N_24757,N_24665);
xnor U26232 (N_26232,N_24416,N_24977);
xor U26233 (N_26233,N_24235,N_24827);
and U26234 (N_26234,N_24485,N_24093);
and U26235 (N_26235,N_24721,N_24086);
or U26236 (N_26236,N_24922,N_24560);
nor U26237 (N_26237,N_24139,N_25070);
or U26238 (N_26238,N_24707,N_24179);
or U26239 (N_26239,N_25150,N_24297);
nor U26240 (N_26240,N_24995,N_24589);
or U26241 (N_26241,N_24606,N_25198);
nor U26242 (N_26242,N_24665,N_24332);
xnor U26243 (N_26243,N_24355,N_24383);
and U26244 (N_26244,N_24105,N_24119);
and U26245 (N_26245,N_24179,N_24768);
or U26246 (N_26246,N_24674,N_24973);
or U26247 (N_26247,N_25018,N_24158);
and U26248 (N_26248,N_24233,N_24760);
nor U26249 (N_26249,N_24714,N_25115);
and U26250 (N_26250,N_25007,N_24015);
nor U26251 (N_26251,N_24542,N_24974);
xor U26252 (N_26252,N_24119,N_24983);
xnor U26253 (N_26253,N_24376,N_24226);
nand U26254 (N_26254,N_24186,N_24972);
and U26255 (N_26255,N_24257,N_24277);
and U26256 (N_26256,N_24142,N_25166);
nand U26257 (N_26257,N_25130,N_24287);
or U26258 (N_26258,N_24852,N_24088);
nor U26259 (N_26259,N_24873,N_24620);
or U26260 (N_26260,N_24223,N_24345);
and U26261 (N_26261,N_24613,N_24001);
or U26262 (N_26262,N_24796,N_24877);
and U26263 (N_26263,N_24064,N_24570);
nand U26264 (N_26264,N_24918,N_24131);
nand U26265 (N_26265,N_24363,N_24045);
or U26266 (N_26266,N_24294,N_24004);
nor U26267 (N_26267,N_24273,N_24998);
nand U26268 (N_26268,N_24347,N_24158);
nor U26269 (N_26269,N_24729,N_24335);
xnor U26270 (N_26270,N_24338,N_24321);
xor U26271 (N_26271,N_24034,N_24060);
xor U26272 (N_26272,N_24234,N_24837);
nand U26273 (N_26273,N_24888,N_24703);
xor U26274 (N_26274,N_24295,N_24593);
xor U26275 (N_26275,N_24798,N_24708);
xnor U26276 (N_26276,N_24357,N_24485);
nor U26277 (N_26277,N_24704,N_24794);
xnor U26278 (N_26278,N_24128,N_24937);
and U26279 (N_26279,N_24963,N_24232);
xor U26280 (N_26280,N_24325,N_24703);
and U26281 (N_26281,N_24678,N_25182);
or U26282 (N_26282,N_24121,N_24342);
and U26283 (N_26283,N_24618,N_24982);
and U26284 (N_26284,N_24400,N_24658);
and U26285 (N_26285,N_25058,N_24275);
or U26286 (N_26286,N_24628,N_24586);
or U26287 (N_26287,N_24754,N_24916);
or U26288 (N_26288,N_24219,N_24563);
or U26289 (N_26289,N_24381,N_24732);
nor U26290 (N_26290,N_24578,N_25092);
and U26291 (N_26291,N_24219,N_24543);
xor U26292 (N_26292,N_24249,N_24996);
and U26293 (N_26293,N_24989,N_24106);
and U26294 (N_26294,N_24687,N_25133);
and U26295 (N_26295,N_24780,N_24216);
nor U26296 (N_26296,N_24776,N_24779);
or U26297 (N_26297,N_24645,N_24595);
or U26298 (N_26298,N_24765,N_24348);
nand U26299 (N_26299,N_24562,N_24866);
and U26300 (N_26300,N_24916,N_24816);
nand U26301 (N_26301,N_24844,N_24204);
and U26302 (N_26302,N_25078,N_24177);
or U26303 (N_26303,N_24331,N_25009);
nand U26304 (N_26304,N_24216,N_24738);
nor U26305 (N_26305,N_24630,N_24320);
xor U26306 (N_26306,N_24929,N_24521);
and U26307 (N_26307,N_24872,N_24572);
nor U26308 (N_26308,N_24370,N_24133);
or U26309 (N_26309,N_24836,N_24092);
or U26310 (N_26310,N_24146,N_24210);
nand U26311 (N_26311,N_25155,N_24433);
nor U26312 (N_26312,N_25005,N_25035);
nand U26313 (N_26313,N_24800,N_24682);
nor U26314 (N_26314,N_25153,N_24689);
xor U26315 (N_26315,N_24150,N_24786);
nand U26316 (N_26316,N_24141,N_24607);
and U26317 (N_26317,N_25140,N_24108);
nand U26318 (N_26318,N_24955,N_24665);
nor U26319 (N_26319,N_25084,N_24931);
or U26320 (N_26320,N_24618,N_24665);
nor U26321 (N_26321,N_24578,N_24869);
nand U26322 (N_26322,N_24553,N_24191);
xnor U26323 (N_26323,N_24077,N_25006);
nand U26324 (N_26324,N_24749,N_24591);
nand U26325 (N_26325,N_24758,N_24429);
and U26326 (N_26326,N_24712,N_24675);
or U26327 (N_26327,N_24137,N_24194);
and U26328 (N_26328,N_24598,N_24683);
nor U26329 (N_26329,N_24387,N_24447);
nor U26330 (N_26330,N_24923,N_24850);
and U26331 (N_26331,N_24711,N_24964);
xor U26332 (N_26332,N_24447,N_24966);
nand U26333 (N_26333,N_25198,N_24217);
nor U26334 (N_26334,N_24100,N_24730);
or U26335 (N_26335,N_24209,N_24296);
or U26336 (N_26336,N_24526,N_24448);
or U26337 (N_26337,N_24034,N_24217);
xor U26338 (N_26338,N_24256,N_24313);
xor U26339 (N_26339,N_24500,N_24418);
nand U26340 (N_26340,N_24041,N_24597);
and U26341 (N_26341,N_24461,N_24145);
nor U26342 (N_26342,N_24096,N_24136);
nand U26343 (N_26343,N_24164,N_24837);
or U26344 (N_26344,N_24679,N_24863);
nor U26345 (N_26345,N_24163,N_24142);
xnor U26346 (N_26346,N_24130,N_24930);
nor U26347 (N_26347,N_24896,N_25106);
or U26348 (N_26348,N_24119,N_24894);
nand U26349 (N_26349,N_24083,N_24578);
nor U26350 (N_26350,N_25079,N_24600);
nand U26351 (N_26351,N_25042,N_24888);
nor U26352 (N_26352,N_24992,N_24582);
nand U26353 (N_26353,N_24603,N_25128);
and U26354 (N_26354,N_24367,N_24554);
nand U26355 (N_26355,N_24180,N_24430);
nand U26356 (N_26356,N_24840,N_24182);
and U26357 (N_26357,N_25095,N_24075);
or U26358 (N_26358,N_25026,N_24832);
nor U26359 (N_26359,N_24108,N_24174);
nor U26360 (N_26360,N_24852,N_24806);
xnor U26361 (N_26361,N_25082,N_24468);
nor U26362 (N_26362,N_24723,N_24318);
nor U26363 (N_26363,N_24742,N_24947);
or U26364 (N_26364,N_24650,N_24333);
nor U26365 (N_26365,N_25113,N_24441);
and U26366 (N_26366,N_24407,N_24050);
nor U26367 (N_26367,N_24937,N_24102);
and U26368 (N_26368,N_24221,N_24551);
nor U26369 (N_26369,N_24458,N_24899);
or U26370 (N_26370,N_24599,N_24800);
nor U26371 (N_26371,N_25066,N_25115);
or U26372 (N_26372,N_25184,N_25016);
and U26373 (N_26373,N_24312,N_25150);
nand U26374 (N_26374,N_24986,N_24700);
and U26375 (N_26375,N_24706,N_24372);
nor U26376 (N_26376,N_24319,N_24990);
nand U26377 (N_26377,N_24472,N_24262);
nor U26378 (N_26378,N_24275,N_24956);
nand U26379 (N_26379,N_24371,N_24045);
or U26380 (N_26380,N_24653,N_24233);
nand U26381 (N_26381,N_24213,N_24426);
or U26382 (N_26382,N_24471,N_24073);
nand U26383 (N_26383,N_25013,N_24527);
or U26384 (N_26384,N_24579,N_24071);
or U26385 (N_26385,N_24276,N_24426);
and U26386 (N_26386,N_24119,N_24369);
nand U26387 (N_26387,N_24912,N_24713);
nor U26388 (N_26388,N_24988,N_24219);
nor U26389 (N_26389,N_24091,N_24839);
or U26390 (N_26390,N_24409,N_25023);
xnor U26391 (N_26391,N_24673,N_24946);
or U26392 (N_26392,N_25182,N_24628);
nor U26393 (N_26393,N_24038,N_24008);
xor U26394 (N_26394,N_24538,N_24268);
and U26395 (N_26395,N_24801,N_25081);
nand U26396 (N_26396,N_24639,N_24406);
and U26397 (N_26397,N_24022,N_24550);
or U26398 (N_26398,N_24034,N_24626);
or U26399 (N_26399,N_24532,N_25142);
xor U26400 (N_26400,N_25730,N_25366);
xor U26401 (N_26401,N_25758,N_25279);
nand U26402 (N_26402,N_25639,N_25235);
or U26403 (N_26403,N_25455,N_25899);
and U26404 (N_26404,N_25516,N_25264);
nand U26405 (N_26405,N_25253,N_25781);
nand U26406 (N_26406,N_25221,N_25607);
xnor U26407 (N_26407,N_25316,N_25827);
xnor U26408 (N_26408,N_26112,N_25356);
xnor U26409 (N_26409,N_26250,N_26300);
nor U26410 (N_26410,N_26232,N_25724);
and U26411 (N_26411,N_26394,N_25991);
and U26412 (N_26412,N_26120,N_26380);
or U26413 (N_26413,N_25473,N_25289);
or U26414 (N_26414,N_25663,N_26248);
and U26415 (N_26415,N_25780,N_26230);
nor U26416 (N_26416,N_26385,N_25201);
nand U26417 (N_26417,N_25904,N_26395);
nand U26418 (N_26418,N_26007,N_26314);
xor U26419 (N_26419,N_26275,N_25964);
and U26420 (N_26420,N_26301,N_25840);
nor U26421 (N_26421,N_25797,N_26029);
and U26422 (N_26422,N_26281,N_25761);
or U26423 (N_26423,N_25450,N_25882);
or U26424 (N_26424,N_26286,N_26043);
nand U26425 (N_26425,N_25677,N_25521);
nand U26426 (N_26426,N_25465,N_26060);
or U26427 (N_26427,N_25265,N_25843);
or U26428 (N_26428,N_25210,N_25658);
and U26429 (N_26429,N_26332,N_25898);
or U26430 (N_26430,N_25272,N_26073);
xor U26431 (N_26431,N_26303,N_25218);
or U26432 (N_26432,N_26276,N_25349);
xor U26433 (N_26433,N_25337,N_25969);
or U26434 (N_26434,N_25492,N_26016);
and U26435 (N_26435,N_25872,N_25255);
nor U26436 (N_26436,N_25354,N_25252);
nand U26437 (N_26437,N_25951,N_25963);
xor U26438 (N_26438,N_25747,N_25393);
or U26439 (N_26439,N_25546,N_25748);
or U26440 (N_26440,N_25223,N_25438);
or U26441 (N_26441,N_26117,N_26199);
and U26442 (N_26442,N_26200,N_25905);
and U26443 (N_26443,N_26165,N_25869);
nor U26444 (N_26444,N_25359,N_25352);
xnor U26445 (N_26445,N_26113,N_26134);
xnor U26446 (N_26446,N_25555,N_25286);
nor U26447 (N_26447,N_25595,N_25412);
xor U26448 (N_26448,N_25532,N_26090);
nor U26449 (N_26449,N_25541,N_26126);
xnor U26450 (N_26450,N_25609,N_25915);
and U26451 (N_26451,N_25824,N_25529);
xor U26452 (N_26452,N_25849,N_25464);
nor U26453 (N_26453,N_25788,N_26004);
or U26454 (N_26454,N_26040,N_25580);
or U26455 (N_26455,N_25665,N_25929);
and U26456 (N_26456,N_25912,N_25416);
or U26457 (N_26457,N_26186,N_25628);
xnor U26458 (N_26458,N_26168,N_26012);
or U26459 (N_26459,N_26274,N_25340);
and U26460 (N_26460,N_25706,N_25925);
nor U26461 (N_26461,N_25254,N_25568);
or U26462 (N_26462,N_26325,N_26384);
nor U26463 (N_26463,N_26291,N_26202);
nand U26464 (N_26464,N_25791,N_25950);
and U26465 (N_26465,N_25792,N_26098);
or U26466 (N_26466,N_26011,N_26082);
or U26467 (N_26467,N_25533,N_25530);
nor U26468 (N_26468,N_26035,N_26141);
or U26469 (N_26469,N_25859,N_25268);
nor U26470 (N_26470,N_25461,N_25996);
nor U26471 (N_26471,N_25266,N_25673);
xor U26472 (N_26472,N_25491,N_25680);
and U26473 (N_26473,N_25392,N_25604);
nor U26474 (N_26474,N_26024,N_25570);
xnor U26475 (N_26475,N_25752,N_25594);
xor U26476 (N_26476,N_26344,N_25755);
nor U26477 (N_26477,N_26270,N_25696);
and U26478 (N_26478,N_25861,N_26118);
nor U26479 (N_26479,N_25717,N_26062);
nand U26480 (N_26480,N_25232,N_25686);
nand U26481 (N_26481,N_25917,N_26234);
or U26482 (N_26482,N_25224,N_25308);
and U26483 (N_26483,N_25795,N_25679);
nand U26484 (N_26484,N_26310,N_25575);
and U26485 (N_26485,N_25848,N_25259);
nand U26486 (N_26486,N_25886,N_25208);
xnor U26487 (N_26487,N_25338,N_26006);
nand U26488 (N_26488,N_25466,N_25207);
xor U26489 (N_26489,N_25376,N_26175);
nor U26490 (N_26490,N_25468,N_25962);
nor U26491 (N_26491,N_25343,N_26026);
and U26492 (N_26492,N_26107,N_25972);
or U26493 (N_26493,N_25275,N_25411);
or U26494 (N_26494,N_25344,N_26137);
nand U26495 (N_26495,N_25514,N_25754);
xnor U26496 (N_26496,N_25690,N_26143);
xnor U26497 (N_26497,N_25321,N_26241);
or U26498 (N_26498,N_25767,N_26072);
xnor U26499 (N_26499,N_25378,N_25811);
or U26500 (N_26500,N_25787,N_26002);
xnor U26501 (N_26501,N_25261,N_25612);
nand U26502 (N_26502,N_25834,N_25428);
or U26503 (N_26503,N_26280,N_25652);
or U26504 (N_26504,N_26321,N_25558);
and U26505 (N_26505,N_26162,N_26256);
and U26506 (N_26506,N_25688,N_26139);
nor U26507 (N_26507,N_25992,N_25336);
or U26508 (N_26508,N_25852,N_25676);
or U26509 (N_26509,N_26214,N_25870);
or U26510 (N_26510,N_25236,N_25425);
nand U26511 (N_26511,N_25407,N_25641);
or U26512 (N_26512,N_26338,N_25248);
or U26513 (N_26513,N_26309,N_26375);
and U26514 (N_26514,N_26263,N_26316);
nand U26515 (N_26515,N_25814,N_25273);
xor U26516 (N_26516,N_25726,N_25550);
xnor U26517 (N_26517,N_25484,N_25556);
or U26518 (N_26518,N_25744,N_25368);
and U26519 (N_26519,N_25957,N_25683);
nand U26520 (N_26520,N_25889,N_25858);
nor U26521 (N_26521,N_26224,N_26179);
nor U26522 (N_26522,N_25333,N_25678);
nor U26523 (N_26523,N_25485,N_25241);
nor U26524 (N_26524,N_26071,N_25311);
and U26525 (N_26525,N_26324,N_26292);
xor U26526 (N_26526,N_25495,N_26068);
and U26527 (N_26527,N_26238,N_26251);
or U26528 (N_26528,N_26272,N_25472);
xor U26529 (N_26529,N_25624,N_26271);
nand U26530 (N_26530,N_25574,N_25384);
nand U26531 (N_26531,N_25524,N_25672);
xor U26532 (N_26532,N_25206,N_26067);
nor U26533 (N_26533,N_25545,N_25305);
nor U26534 (N_26534,N_25290,N_25507);
and U26535 (N_26535,N_25990,N_26302);
or U26536 (N_26536,N_25256,N_25871);
or U26537 (N_26537,N_25939,N_26099);
and U26538 (N_26538,N_25816,N_26336);
or U26539 (N_26539,N_26086,N_26294);
or U26540 (N_26540,N_26180,N_25757);
nand U26541 (N_26541,N_26084,N_25271);
nand U26542 (N_26542,N_26153,N_25613);
and U26543 (N_26543,N_26341,N_26299);
xor U26544 (N_26544,N_26381,N_25267);
xnor U26545 (N_26545,N_25937,N_26279);
nor U26546 (N_26546,N_25999,N_26081);
or U26547 (N_26547,N_26064,N_26282);
xor U26548 (N_26548,N_25711,N_25723);
nand U26549 (N_26549,N_25873,N_25225);
nor U26550 (N_26550,N_25629,N_25238);
and U26551 (N_26551,N_25260,N_25847);
nor U26552 (N_26552,N_25681,N_25597);
or U26553 (N_26553,N_26017,N_26221);
and U26554 (N_26554,N_25883,N_25978);
or U26555 (N_26555,N_25875,N_25371);
nand U26556 (N_26556,N_25935,N_25650);
or U26557 (N_26557,N_25421,N_25874);
nand U26558 (N_26558,N_25328,N_25535);
nor U26559 (N_26559,N_25348,N_25908);
and U26560 (N_26560,N_25429,N_25245);
nor U26561 (N_26561,N_26036,N_25487);
or U26562 (N_26562,N_26323,N_25638);
xor U26563 (N_26563,N_25893,N_25299);
xor U26564 (N_26564,N_26111,N_25561);
nor U26565 (N_26565,N_26041,N_26167);
or U26566 (N_26566,N_25435,N_25394);
or U26567 (N_26567,N_25388,N_26399);
nor U26568 (N_26568,N_26397,N_25242);
xnor U26569 (N_26569,N_26236,N_25948);
xnor U26570 (N_26570,N_25621,N_26097);
nor U26571 (N_26571,N_25590,N_25572);
and U26572 (N_26572,N_26161,N_25775);
nor U26573 (N_26573,N_25903,N_25581);
xor U26574 (N_26574,N_25810,N_25285);
or U26575 (N_26575,N_26362,N_26034);
nor U26576 (N_26576,N_25405,N_26019);
and U26577 (N_26577,N_25800,N_25857);
xor U26578 (N_26578,N_25911,N_25721);
xnor U26579 (N_26579,N_25578,N_25988);
and U26580 (N_26580,N_25569,N_25505);
and U26581 (N_26581,N_25370,N_25941);
nand U26582 (N_26582,N_25377,N_26229);
nand U26583 (N_26583,N_26258,N_26374);
or U26584 (N_26584,N_26094,N_25630);
and U26585 (N_26585,N_25325,N_26077);
xor U26586 (N_26586,N_26049,N_25753);
xor U26587 (N_26587,N_26315,N_26003);
and U26588 (N_26588,N_26208,N_26212);
nand U26589 (N_26589,N_25646,N_25975);
or U26590 (N_26590,N_25654,N_25804);
nand U26591 (N_26591,N_25387,N_25430);
or U26592 (N_26592,N_25458,N_25353);
and U26593 (N_26593,N_25719,N_25381);
and U26594 (N_26594,N_25436,N_25651);
and U26595 (N_26595,N_25296,N_25949);
xnor U26596 (N_26596,N_25854,N_25291);
nand U26597 (N_26597,N_25868,N_26340);
and U26598 (N_26598,N_25486,N_25973);
xor U26599 (N_26599,N_26259,N_26185);
and U26600 (N_26600,N_25283,N_25965);
nor U26601 (N_26601,N_26023,N_25821);
xor U26602 (N_26602,N_26377,N_25801);
nor U26603 (N_26603,N_25398,N_26151);
nor U26604 (N_26604,N_25924,N_26135);
and U26605 (N_26605,N_25923,N_26158);
nor U26606 (N_26606,N_25234,N_25667);
and U26607 (N_26607,N_26376,N_26237);
nand U26608 (N_26608,N_25300,N_25361);
nor U26609 (N_26609,N_26193,N_25853);
xor U26610 (N_26610,N_26104,N_26218);
nand U26611 (N_26611,N_25863,N_26222);
xor U26612 (N_26612,N_25502,N_25576);
or U26613 (N_26613,N_25961,N_26354);
xnor U26614 (N_26614,N_25549,N_25608);
nor U26615 (N_26615,N_25482,N_26345);
or U26616 (N_26616,N_26176,N_25312);
xnor U26617 (N_26617,N_26333,N_25735);
or U26618 (N_26618,N_26014,N_25790);
xor U26619 (N_26619,N_25895,N_25481);
nor U26620 (N_26620,N_26058,N_25213);
and U26621 (N_26621,N_26327,N_26391);
nand U26622 (N_26622,N_25986,N_25557);
nand U26623 (N_26623,N_25825,N_25441);
xnor U26624 (N_26624,N_25842,N_26116);
nor U26625 (N_26625,N_25479,N_25776);
nor U26626 (N_26626,N_25669,N_25523);
and U26627 (N_26627,N_25415,N_26147);
or U26628 (N_26628,N_26129,N_26089);
and U26629 (N_26629,N_25226,N_26051);
and U26630 (N_26630,N_25866,N_25439);
xor U26631 (N_26631,N_25729,N_26095);
nand U26632 (N_26632,N_25771,N_25940);
nor U26633 (N_26633,N_25709,N_26273);
xor U26634 (N_26634,N_25692,N_25513);
nand U26635 (N_26635,N_26030,N_25701);
or U26636 (N_26636,N_25577,N_25860);
nand U26637 (N_26637,N_25540,N_25918);
nor U26638 (N_26638,N_25768,N_26061);
and U26639 (N_26639,N_25967,N_25725);
nor U26640 (N_26640,N_25262,N_25548);
nor U26641 (N_26641,N_25712,N_26226);
and U26642 (N_26642,N_26288,N_26210);
and U26643 (N_26643,N_25876,N_26239);
xnor U26644 (N_26644,N_25317,N_25520);
nand U26645 (N_26645,N_26293,N_25622);
nor U26646 (N_26646,N_25298,N_26265);
nor U26647 (N_26647,N_25553,N_25329);
nand U26648 (N_26648,N_26046,N_26289);
nand U26649 (N_26649,N_25503,N_25508);
xor U26650 (N_26650,N_26055,N_26266);
nand U26651 (N_26651,N_26219,N_25644);
nor U26652 (N_26652,N_25304,N_25471);
xnor U26653 (N_26653,N_25433,N_25326);
nand U26654 (N_26654,N_26181,N_25493);
nor U26655 (N_26655,N_26021,N_25350);
nor U26656 (N_26656,N_25976,N_26109);
or U26657 (N_26657,N_25534,N_26205);
or U26658 (N_26658,N_26198,N_25240);
xnor U26659 (N_26659,N_25380,N_26196);
nor U26660 (N_26660,N_25227,N_26177);
nand U26661 (N_26661,N_25539,N_26370);
nor U26662 (N_26662,N_26102,N_26353);
or U26663 (N_26663,N_26096,N_26393);
or U26664 (N_26664,N_25704,N_26308);
and U26665 (N_26665,N_26169,N_25422);
nor U26666 (N_26666,N_25634,N_25382);
nand U26667 (N_26667,N_25896,N_25664);
and U26668 (N_26668,N_26334,N_26190);
nor U26669 (N_26669,N_26038,N_26243);
and U26670 (N_26670,N_26110,N_25258);
nand U26671 (N_26671,N_25391,N_25922);
nor U26672 (N_26672,N_25647,N_25799);
nor U26673 (N_26673,N_25426,N_25611);
xnor U26674 (N_26674,N_25718,N_25734);
nand U26675 (N_26675,N_25246,N_26351);
or U26676 (N_26676,N_25635,N_26093);
nor U26677 (N_26677,N_25274,N_25499);
nor U26678 (N_26678,N_26298,N_25462);
and U26679 (N_26679,N_25987,N_25537);
nor U26680 (N_26680,N_25947,N_25884);
xor U26681 (N_26681,N_25442,N_25528);
xnor U26682 (N_26682,N_26010,N_26028);
or U26683 (N_26683,N_25307,N_25294);
nor U26684 (N_26684,N_26080,N_25313);
nor U26685 (N_26685,N_25803,N_26358);
and U26686 (N_26686,N_26356,N_25865);
xnor U26687 (N_26687,N_25983,N_25456);
or U26688 (N_26688,N_25440,N_25731);
nor U26689 (N_26689,N_26152,N_26382);
nor U26690 (N_26690,N_25897,N_25902);
nor U26691 (N_26691,N_26059,N_25832);
and U26692 (N_26692,N_26159,N_25280);
and U26693 (N_26693,N_26048,N_25765);
or U26694 (N_26694,N_25817,N_25292);
and U26695 (N_26695,N_25997,N_25542);
or U26696 (N_26696,N_25603,N_25447);
nor U26697 (N_26697,N_25355,N_26335);
or U26698 (N_26698,N_26204,N_25457);
or U26699 (N_26699,N_26357,N_25977);
nor U26700 (N_26700,N_25373,N_26203);
and U26701 (N_26701,N_25879,N_26262);
nand U26702 (N_26702,N_26398,N_25510);
or U26703 (N_26703,N_25203,N_25693);
nand U26704 (N_26704,N_25489,N_25599);
xor U26705 (N_26705,N_26087,N_25829);
xor U26706 (N_26706,N_25494,N_25470);
or U26707 (N_26707,N_25501,N_26170);
xnor U26708 (N_26708,N_25971,N_26331);
or U26709 (N_26709,N_26085,N_25217);
nor U26710 (N_26710,N_26296,N_25877);
and U26711 (N_26711,N_25400,N_25600);
or U26712 (N_26712,N_25362,N_25878);
nand U26713 (N_26713,N_25293,N_25661);
xnor U26714 (N_26714,N_26148,N_25623);
and U26715 (N_26715,N_25845,N_26386);
and U26716 (N_26716,N_26027,N_25714);
and U26717 (N_26717,N_25695,N_25566);
xnor U26718 (N_26718,N_25324,N_25741);
and U26719 (N_26719,N_25547,N_25943);
and U26720 (N_26720,N_25200,N_25270);
xnor U26721 (N_26721,N_25921,N_25383);
or U26722 (N_26722,N_25946,N_25443);
nor U26723 (N_26723,N_25367,N_25815);
and U26724 (N_26724,N_26305,N_25490);
xor U26725 (N_26725,N_25675,N_26131);
nand U26726 (N_26726,N_25389,N_26240);
and U26727 (N_26727,N_26031,N_25985);
or U26728 (N_26728,N_25579,N_25615);
nor U26729 (N_26729,N_25617,N_25360);
xnor U26730 (N_26730,N_25331,N_26150);
xor U26731 (N_26731,N_25739,N_25998);
and U26732 (N_26732,N_25297,N_25610);
nand U26733 (N_26733,N_26389,N_25424);
and U26734 (N_26734,N_25320,N_25759);
and U26735 (N_26735,N_25284,N_26235);
xor U26736 (N_26736,N_25205,N_25419);
nor U26737 (N_26737,N_25894,N_25584);
nand U26738 (N_26738,N_25784,N_25928);
nand U26739 (N_26739,N_25335,N_25809);
xor U26740 (N_26740,N_25525,N_25710);
and U26741 (N_26741,N_25907,N_25705);
nand U26742 (N_26742,N_25365,N_25666);
or U26743 (N_26743,N_26368,N_25993);
and U26744 (N_26744,N_26092,N_26105);
nor U26745 (N_26745,N_26330,N_26146);
and U26746 (N_26746,N_25526,N_25636);
and U26747 (N_26747,N_25850,N_25431);
or U26748 (N_26748,N_25720,N_26290);
xnor U26749 (N_26749,N_25209,N_26171);
nand U26750 (N_26750,N_26337,N_26268);
nand U26751 (N_26751,N_25633,N_25645);
nor U26752 (N_26752,N_25480,N_25745);
or U26753 (N_26753,N_25216,N_25778);
nor U26754 (N_26754,N_25760,N_26254);
xor U26755 (N_26755,N_25958,N_26350);
xnor U26756 (N_26756,N_25698,N_26194);
and U26757 (N_26757,N_26020,N_25229);
nand U26758 (N_26758,N_25970,N_25420);
or U26759 (N_26759,N_26339,N_26363);
nor U26760 (N_26760,N_26255,N_25732);
xnor U26761 (N_26761,N_25750,N_25979);
nand U26762 (N_26762,N_26145,N_25498);
nor U26763 (N_26763,N_25269,N_26253);
and U26764 (N_26764,N_25995,N_26053);
or U26765 (N_26765,N_25257,N_26378);
and U26766 (N_26766,N_25880,N_25914);
and U26767 (N_26767,N_26065,N_25397);
nor U26768 (N_26768,N_26388,N_25589);
xnor U26769 (N_26769,N_25697,N_26367);
xnor U26770 (N_26770,N_25427,N_26192);
and U26771 (N_26771,N_25315,N_25451);
xnor U26772 (N_26772,N_26039,N_25782);
nand U26773 (N_26773,N_26366,N_25944);
or U26774 (N_26774,N_25806,N_25476);
xnor U26775 (N_26775,N_25445,N_26127);
xor U26776 (N_26776,N_25864,N_25437);
or U26777 (N_26777,N_25770,N_25418);
nor U26778 (N_26778,N_26312,N_26283);
nand U26779 (N_26779,N_26361,N_25909);
and U26780 (N_26780,N_25214,N_25994);
nand U26781 (N_26781,N_25694,N_25601);
and U26782 (N_26782,N_25945,N_25452);
xnor U26783 (N_26783,N_25682,N_26343);
xor U26784 (N_26784,N_26249,N_25934);
xnor U26785 (N_26785,N_25777,N_25737);
nand U26786 (N_26786,N_25385,N_25459);
nand U26787 (N_26787,N_25567,N_25571);
nor U26788 (N_26788,N_26297,N_25277);
and U26789 (N_26789,N_25318,N_25736);
nor U26790 (N_26790,N_26184,N_26128);
nand U26791 (N_26791,N_25512,N_25469);
nand U26792 (N_26792,N_25700,N_25231);
xnor U26793 (N_26793,N_25543,N_26033);
and U26794 (N_26794,N_26018,N_26042);
nand U26795 (N_26795,N_26233,N_26140);
nand U26796 (N_26796,N_25478,N_26130);
and U26797 (N_26797,N_25616,N_26285);
nand U26798 (N_26798,N_26326,N_25808);
and U26799 (N_26799,N_26242,N_26227);
and U26800 (N_26800,N_25938,N_26217);
nand U26801 (N_26801,N_25786,N_26245);
and U26802 (N_26802,N_25358,N_25497);
and U26803 (N_26803,N_25984,N_26342);
or U26804 (N_26804,N_25506,N_25341);
xnor U26805 (N_26805,N_25793,N_26329);
nand U26806 (N_26806,N_26057,N_25685);
or U26807 (N_26807,N_25762,N_25743);
or U26808 (N_26808,N_26075,N_26246);
xor U26809 (N_26809,N_25715,N_26121);
xor U26810 (N_26810,N_26348,N_25432);
or U26811 (N_26811,N_25835,N_25504);
nand U26812 (N_26812,N_25774,N_25386);
and U26813 (N_26813,N_25867,N_25942);
and U26814 (N_26814,N_25802,N_25891);
and U26815 (N_26815,N_26304,N_26088);
and U26816 (N_26816,N_26247,N_26063);
or U26817 (N_26817,N_26083,N_25538);
or U26818 (N_26818,N_25454,N_26213);
xor U26819 (N_26819,N_25372,N_25822);
xor U26820 (N_26820,N_25332,N_25374);
and U26821 (N_26821,N_25851,N_25892);
nor U26822 (N_26822,N_25831,N_26122);
and U26823 (N_26823,N_26277,N_25306);
and U26824 (N_26824,N_25310,N_25295);
or U26825 (N_26825,N_26396,N_26373);
and U26826 (N_26826,N_25763,N_25573);
and U26827 (N_26827,N_25837,N_26307);
nand U26828 (N_26828,N_26347,N_26076);
nor U26829 (N_26829,N_25733,N_26101);
nand U26830 (N_26830,N_25563,N_25363);
nand U26831 (N_26831,N_26000,N_25239);
and U26832 (N_26832,N_26009,N_26360);
nand U26833 (N_26833,N_26133,N_26015);
and U26834 (N_26834,N_25444,N_25519);
or U26835 (N_26835,N_25544,N_25954);
nor U26836 (N_26836,N_25467,N_26001);
nand U26837 (N_26837,N_26178,N_26317);
or U26838 (N_26838,N_26022,N_25631);
xor U26839 (N_26839,N_26164,N_25900);
xnor U26840 (N_26840,N_26187,N_25278);
nand U26841 (N_26841,N_26392,N_26163);
xnor U26842 (N_26842,N_26149,N_26079);
or U26843 (N_26843,N_25281,N_26005);
xor U26844 (N_26844,N_26056,N_25766);
nor U26845 (N_26845,N_25772,N_25779);
and U26846 (N_26846,N_26166,N_25417);
nand U26847 (N_26847,N_25828,N_26295);
and U26848 (N_26848,N_25346,N_25689);
xor U26849 (N_26849,N_25856,N_25659);
nand U26850 (N_26850,N_25475,N_25906);
nand U26851 (N_26851,N_25602,N_26138);
nor U26852 (N_26852,N_25322,N_25204);
nor U26853 (N_26853,N_25794,N_26114);
nor U26854 (N_26854,N_25598,N_25233);
nor U26855 (N_26855,N_25699,N_26188);
or U26856 (N_26856,N_26284,N_25395);
nor U26857 (N_26857,N_25327,N_25660);
nor U26858 (N_26858,N_25727,N_25740);
nand U26859 (N_26859,N_25583,N_26264);
or U26860 (N_26860,N_25703,N_25565);
xnor U26861 (N_26861,N_26108,N_25674);
nor U26862 (N_26862,N_25930,N_26201);
xor U26863 (N_26863,N_25536,N_25742);
xnor U26864 (N_26864,N_25477,N_25423);
xor U26865 (N_26865,N_25404,N_25926);
xor U26866 (N_26866,N_26244,N_25403);
nor U26867 (N_26867,N_25756,N_25463);
xnor U26868 (N_26868,N_25769,N_25913);
nand U26869 (N_26869,N_25656,N_25846);
xnor U26870 (N_26870,N_25955,N_25627);
nor U26871 (N_26871,N_25862,N_25936);
nor U26872 (N_26872,N_26223,N_25968);
and U26873 (N_26873,N_25396,N_26372);
nand U26874 (N_26874,N_26013,N_26050);
and U26875 (N_26875,N_25632,N_25890);
nand U26876 (N_26876,N_25881,N_25989);
nor U26877 (N_26877,N_25562,N_25369);
and U26878 (N_26878,N_26359,N_25215);
and U26879 (N_26879,N_26206,N_25222);
xnor U26880 (N_26880,N_26069,N_26106);
xnor U26881 (N_26881,N_26225,N_25818);
nand U26882 (N_26882,N_25956,N_25728);
and U26883 (N_26883,N_25836,N_26349);
xnor U26884 (N_26884,N_25687,N_26125);
nand U26885 (N_26885,N_26364,N_26261);
nand U26886 (N_26886,N_26123,N_26231);
xnor U26887 (N_26887,N_25515,N_26154);
nor U26888 (N_26888,N_25596,N_25798);
or U26889 (N_26889,N_26355,N_25982);
nor U26890 (N_26890,N_25531,N_26365);
nor U26891 (N_26891,N_25713,N_25522);
xnor U26892 (N_26892,N_25981,N_25564);
xnor U26893 (N_26893,N_25960,N_25345);
xor U26894 (N_26894,N_26195,N_26115);
nand U26895 (N_26895,N_25402,N_25764);
nand U26896 (N_26896,N_25244,N_26025);
nor U26897 (N_26897,N_25309,N_25406);
nand U26898 (N_26898,N_25500,N_25707);
nor U26899 (N_26899,N_25483,N_25605);
nor U26900 (N_26900,N_25640,N_25657);
xor U26901 (N_26901,N_25276,N_25953);
nor U26902 (N_26902,N_25585,N_25287);
nand U26903 (N_26903,N_25474,N_26189);
xor U26904 (N_26904,N_25807,N_25342);
and U26905 (N_26905,N_25805,N_26100);
and U26906 (N_26906,N_26191,N_26346);
nand U26907 (N_26907,N_26320,N_25751);
or U26908 (N_26908,N_26103,N_25448);
and U26909 (N_26909,N_25554,N_26311);
and U26910 (N_26910,N_25974,N_25927);
nor U26911 (N_26911,N_25746,N_25749);
nor U26912 (N_26912,N_26371,N_25830);
nand U26913 (N_26913,N_26278,N_26070);
xnor U26914 (N_26914,N_25347,N_26215);
and U26915 (N_26915,N_26078,N_26044);
nor U26916 (N_26916,N_25409,N_25488);
nand U26917 (N_26917,N_26091,N_25844);
and U26918 (N_26918,N_25219,N_25684);
xnor U26919 (N_26919,N_26174,N_25560);
or U26920 (N_26920,N_25357,N_25351);
xor U26921 (N_26921,N_26054,N_25582);
xnor U26922 (N_26922,N_25716,N_26352);
nand U26923 (N_26923,N_25648,N_25250);
nand U26924 (N_26924,N_25901,N_25401);
or U26925 (N_26925,N_25933,N_25334);
and U26926 (N_26926,N_26379,N_25920);
nand U26927 (N_26927,N_25820,N_26252);
nor U26928 (N_26928,N_25919,N_26136);
or U26929 (N_26929,N_25434,N_26197);
xor U26930 (N_26930,N_26132,N_25303);
nor U26931 (N_26931,N_25453,N_25263);
nor U26932 (N_26932,N_25399,N_25551);
or U26933 (N_26933,N_25789,N_25237);
xnor U26934 (N_26934,N_25625,N_26269);
nand U26935 (N_26935,N_25211,N_25288);
xnor U26936 (N_26936,N_25247,N_26322);
or U26937 (N_26937,N_25243,N_25888);
nand U26938 (N_26938,N_25773,N_25228);
or U26939 (N_26939,N_25379,N_25511);
or U26940 (N_26940,N_26328,N_25410);
nor U26941 (N_26941,N_25855,N_25819);
nor U26942 (N_26942,N_25375,N_25212);
nand U26943 (N_26943,N_25323,N_26319);
and U26944 (N_26944,N_26045,N_25826);
and U26945 (N_26945,N_25980,N_25413);
nand U26946 (N_26946,N_25614,N_25642);
and U26947 (N_26947,N_25620,N_26267);
and U26948 (N_26948,N_25414,N_25885);
xor U26949 (N_26949,N_25449,N_25587);
and U26950 (N_26950,N_25702,N_25796);
and U26951 (N_26951,N_26228,N_26156);
and U26952 (N_26952,N_25588,N_26032);
or U26953 (N_26953,N_25552,N_26124);
or U26954 (N_26954,N_25606,N_26066);
or U26955 (N_26955,N_25653,N_25282);
nand U26956 (N_26956,N_25662,N_25301);
and U26957 (N_26957,N_26047,N_26220);
nand U26958 (N_26958,N_25839,N_25841);
xor U26959 (N_26959,N_25527,N_25586);
nor U26960 (N_26960,N_25649,N_25959);
or U26961 (N_26961,N_25931,N_25643);
nand U26962 (N_26962,N_25932,N_26260);
nand U26963 (N_26963,N_25619,N_26119);
xor U26964 (N_26964,N_26160,N_25966);
and U26965 (N_26965,N_25823,N_25812);
nand U26966 (N_26966,N_25670,N_25783);
xor U26967 (N_26967,N_26207,N_25668);
xnor U26968 (N_26968,N_25671,N_25626);
and U26969 (N_26969,N_25408,N_25364);
nor U26970 (N_26970,N_25446,N_26173);
nor U26971 (N_26971,N_25593,N_25509);
xnor U26972 (N_26972,N_25591,N_26369);
xor U26973 (N_26973,N_25838,N_25496);
or U26974 (N_26974,N_25251,N_25330);
nand U26975 (N_26975,N_26387,N_26008);
or U26976 (N_26976,N_26383,N_26216);
nor U26977 (N_26977,N_26155,N_25813);
nand U26978 (N_26978,N_26157,N_25230);
or U26979 (N_26979,N_26142,N_26209);
nand U26980 (N_26980,N_25559,N_26074);
xnor U26981 (N_26981,N_26037,N_26287);
and U26982 (N_26982,N_26172,N_26211);
or U26983 (N_26983,N_25249,N_25910);
nor U26984 (N_26984,N_25302,N_26183);
nor U26985 (N_26985,N_25390,N_25655);
nand U26986 (N_26986,N_25708,N_26052);
or U26987 (N_26987,N_26257,N_25637);
and U26988 (N_26988,N_25517,N_25319);
nor U26989 (N_26989,N_25618,N_25785);
nand U26990 (N_26990,N_26144,N_26182);
xnor U26991 (N_26991,N_25220,N_25887);
xor U26992 (N_26992,N_25833,N_25592);
nor U26993 (N_26993,N_25518,N_26318);
nand U26994 (N_26994,N_25916,N_26306);
nand U26995 (N_26995,N_25460,N_25202);
and U26996 (N_26996,N_25314,N_25691);
nand U26997 (N_26997,N_26313,N_25339);
xor U26998 (N_26998,N_25738,N_25722);
or U26999 (N_26999,N_26390,N_25952);
and U27000 (N_27000,N_25906,N_26204);
xor U27001 (N_27001,N_25996,N_25348);
or U27002 (N_27002,N_26084,N_25549);
or U27003 (N_27003,N_26260,N_25976);
xor U27004 (N_27004,N_25798,N_25683);
xnor U27005 (N_27005,N_26001,N_25491);
nor U27006 (N_27006,N_26042,N_25465);
xnor U27007 (N_27007,N_25527,N_25347);
or U27008 (N_27008,N_25584,N_26329);
or U27009 (N_27009,N_25772,N_26343);
nor U27010 (N_27010,N_26048,N_25457);
xor U27011 (N_27011,N_25465,N_25243);
or U27012 (N_27012,N_25962,N_25745);
nand U27013 (N_27013,N_26172,N_25893);
or U27014 (N_27014,N_25586,N_26357);
or U27015 (N_27015,N_25446,N_26199);
or U27016 (N_27016,N_25884,N_25762);
or U27017 (N_27017,N_25870,N_25932);
and U27018 (N_27018,N_25438,N_25735);
and U27019 (N_27019,N_25680,N_25401);
and U27020 (N_27020,N_25813,N_25271);
nor U27021 (N_27021,N_25372,N_26362);
or U27022 (N_27022,N_25965,N_25798);
xnor U27023 (N_27023,N_25626,N_26175);
nor U27024 (N_27024,N_25302,N_25313);
and U27025 (N_27025,N_25866,N_25465);
xnor U27026 (N_27026,N_25907,N_25855);
nand U27027 (N_27027,N_25677,N_26195);
nand U27028 (N_27028,N_25414,N_26342);
nand U27029 (N_27029,N_25247,N_26394);
and U27030 (N_27030,N_25354,N_25276);
nand U27031 (N_27031,N_26063,N_26124);
nand U27032 (N_27032,N_26083,N_25668);
or U27033 (N_27033,N_26236,N_25214);
xor U27034 (N_27034,N_25228,N_25605);
or U27035 (N_27035,N_26333,N_25209);
nand U27036 (N_27036,N_26163,N_25560);
nand U27037 (N_27037,N_25624,N_26035);
nand U27038 (N_27038,N_25292,N_26038);
and U27039 (N_27039,N_25228,N_25587);
xor U27040 (N_27040,N_26299,N_26202);
nor U27041 (N_27041,N_25822,N_26220);
nand U27042 (N_27042,N_25794,N_25748);
nor U27043 (N_27043,N_25824,N_25796);
and U27044 (N_27044,N_26378,N_26098);
nand U27045 (N_27045,N_26158,N_25482);
nand U27046 (N_27046,N_25674,N_25945);
nand U27047 (N_27047,N_25779,N_25225);
or U27048 (N_27048,N_25890,N_25367);
nand U27049 (N_27049,N_25740,N_25855);
nor U27050 (N_27050,N_26225,N_26200);
nor U27051 (N_27051,N_25280,N_26134);
or U27052 (N_27052,N_26140,N_25760);
xnor U27053 (N_27053,N_25830,N_25826);
nand U27054 (N_27054,N_26376,N_26162);
nor U27055 (N_27055,N_26130,N_26216);
nand U27056 (N_27056,N_26121,N_26362);
and U27057 (N_27057,N_25371,N_25926);
or U27058 (N_27058,N_26296,N_25638);
nand U27059 (N_27059,N_25368,N_25559);
and U27060 (N_27060,N_25892,N_25335);
and U27061 (N_27061,N_26372,N_25752);
or U27062 (N_27062,N_25817,N_25826);
nor U27063 (N_27063,N_25859,N_25984);
or U27064 (N_27064,N_25432,N_25799);
nor U27065 (N_27065,N_25738,N_26258);
nand U27066 (N_27066,N_26237,N_25891);
or U27067 (N_27067,N_26076,N_26162);
and U27068 (N_27068,N_25304,N_25981);
xnor U27069 (N_27069,N_25638,N_25431);
xnor U27070 (N_27070,N_25892,N_26103);
xnor U27071 (N_27071,N_25297,N_26036);
xnor U27072 (N_27072,N_25927,N_25936);
nand U27073 (N_27073,N_26271,N_25457);
and U27074 (N_27074,N_25290,N_26166);
and U27075 (N_27075,N_25223,N_26338);
and U27076 (N_27076,N_25332,N_26313);
nor U27077 (N_27077,N_25362,N_26276);
or U27078 (N_27078,N_25678,N_25434);
xnor U27079 (N_27079,N_25921,N_26087);
and U27080 (N_27080,N_26112,N_25817);
or U27081 (N_27081,N_25907,N_26275);
nor U27082 (N_27082,N_26308,N_26046);
xnor U27083 (N_27083,N_25399,N_26123);
and U27084 (N_27084,N_25807,N_25438);
and U27085 (N_27085,N_25581,N_26243);
xnor U27086 (N_27086,N_26345,N_25400);
and U27087 (N_27087,N_25686,N_25736);
nand U27088 (N_27088,N_25791,N_26337);
or U27089 (N_27089,N_25292,N_26103);
or U27090 (N_27090,N_25922,N_25781);
nor U27091 (N_27091,N_26284,N_26156);
nand U27092 (N_27092,N_26044,N_25676);
xnor U27093 (N_27093,N_26128,N_25892);
xnor U27094 (N_27094,N_25778,N_25325);
and U27095 (N_27095,N_26225,N_25559);
nor U27096 (N_27096,N_25586,N_25602);
and U27097 (N_27097,N_25330,N_26092);
and U27098 (N_27098,N_25921,N_25310);
nand U27099 (N_27099,N_25277,N_25382);
nor U27100 (N_27100,N_26245,N_25310);
nand U27101 (N_27101,N_26232,N_25311);
xor U27102 (N_27102,N_25781,N_25269);
and U27103 (N_27103,N_25391,N_25587);
nor U27104 (N_27104,N_25589,N_25632);
xor U27105 (N_27105,N_25697,N_25724);
xnor U27106 (N_27106,N_25680,N_25714);
and U27107 (N_27107,N_25431,N_26186);
nor U27108 (N_27108,N_26116,N_26151);
or U27109 (N_27109,N_25501,N_25771);
xor U27110 (N_27110,N_26058,N_25610);
or U27111 (N_27111,N_25781,N_25434);
or U27112 (N_27112,N_25548,N_25868);
nand U27113 (N_27113,N_25923,N_25999);
or U27114 (N_27114,N_25624,N_26202);
or U27115 (N_27115,N_25698,N_25433);
or U27116 (N_27116,N_25522,N_25232);
nand U27117 (N_27117,N_25762,N_26181);
nand U27118 (N_27118,N_25511,N_25507);
nand U27119 (N_27119,N_25840,N_25750);
or U27120 (N_27120,N_26269,N_25270);
and U27121 (N_27121,N_25954,N_26190);
nand U27122 (N_27122,N_25500,N_25398);
nor U27123 (N_27123,N_25381,N_26335);
nor U27124 (N_27124,N_25935,N_25639);
and U27125 (N_27125,N_25296,N_25303);
xnor U27126 (N_27126,N_25804,N_25622);
xor U27127 (N_27127,N_25573,N_25378);
nor U27128 (N_27128,N_25804,N_25889);
nor U27129 (N_27129,N_25825,N_25811);
nand U27130 (N_27130,N_25948,N_26057);
nand U27131 (N_27131,N_26390,N_25893);
nand U27132 (N_27132,N_25658,N_25365);
nand U27133 (N_27133,N_26140,N_25596);
xnor U27134 (N_27134,N_26179,N_26213);
or U27135 (N_27135,N_25236,N_26261);
or U27136 (N_27136,N_26299,N_25207);
xor U27137 (N_27137,N_25608,N_26054);
and U27138 (N_27138,N_25349,N_25315);
nand U27139 (N_27139,N_26236,N_25856);
xor U27140 (N_27140,N_25645,N_25486);
xnor U27141 (N_27141,N_25643,N_26225);
and U27142 (N_27142,N_25611,N_26365);
xor U27143 (N_27143,N_26022,N_26294);
or U27144 (N_27144,N_26002,N_26149);
nor U27145 (N_27145,N_25959,N_26045);
or U27146 (N_27146,N_25486,N_25785);
xor U27147 (N_27147,N_26224,N_25370);
xor U27148 (N_27148,N_25543,N_25467);
nor U27149 (N_27149,N_25882,N_26146);
and U27150 (N_27150,N_26142,N_25442);
xnor U27151 (N_27151,N_25439,N_25959);
and U27152 (N_27152,N_25638,N_25822);
nor U27153 (N_27153,N_25549,N_26278);
xor U27154 (N_27154,N_25624,N_26325);
nand U27155 (N_27155,N_25817,N_26012);
xor U27156 (N_27156,N_25623,N_25965);
xnor U27157 (N_27157,N_25710,N_26156);
xnor U27158 (N_27158,N_26265,N_26310);
nand U27159 (N_27159,N_25455,N_25696);
nor U27160 (N_27160,N_25919,N_26279);
nor U27161 (N_27161,N_25479,N_26156);
nand U27162 (N_27162,N_26248,N_25383);
nand U27163 (N_27163,N_26079,N_25302);
xnor U27164 (N_27164,N_26395,N_25682);
nor U27165 (N_27165,N_26287,N_25960);
and U27166 (N_27166,N_26087,N_25452);
and U27167 (N_27167,N_25955,N_25377);
or U27168 (N_27168,N_26151,N_26393);
xor U27169 (N_27169,N_26274,N_25241);
nor U27170 (N_27170,N_25905,N_25304);
or U27171 (N_27171,N_26170,N_25576);
xor U27172 (N_27172,N_26312,N_25744);
xnor U27173 (N_27173,N_25962,N_26246);
or U27174 (N_27174,N_25999,N_25791);
and U27175 (N_27175,N_25347,N_25681);
nor U27176 (N_27176,N_25246,N_25923);
and U27177 (N_27177,N_25649,N_26352);
or U27178 (N_27178,N_25456,N_25904);
xnor U27179 (N_27179,N_25864,N_25410);
or U27180 (N_27180,N_26253,N_26271);
nand U27181 (N_27181,N_25596,N_25374);
nand U27182 (N_27182,N_25772,N_26308);
xnor U27183 (N_27183,N_25449,N_25697);
nand U27184 (N_27184,N_26314,N_25995);
and U27185 (N_27185,N_25656,N_25808);
nor U27186 (N_27186,N_26036,N_25518);
nand U27187 (N_27187,N_25999,N_26105);
nor U27188 (N_27188,N_25743,N_26292);
xnor U27189 (N_27189,N_26215,N_25822);
xor U27190 (N_27190,N_25645,N_25887);
or U27191 (N_27191,N_25738,N_25859);
or U27192 (N_27192,N_25730,N_25642);
xor U27193 (N_27193,N_25548,N_25893);
nand U27194 (N_27194,N_26010,N_25479);
nor U27195 (N_27195,N_25509,N_25775);
or U27196 (N_27196,N_25884,N_25264);
xnor U27197 (N_27197,N_25991,N_25850);
or U27198 (N_27198,N_25963,N_25843);
nand U27199 (N_27199,N_25202,N_25772);
and U27200 (N_27200,N_26251,N_25549);
and U27201 (N_27201,N_25966,N_25311);
or U27202 (N_27202,N_25245,N_25894);
or U27203 (N_27203,N_26091,N_26197);
and U27204 (N_27204,N_25694,N_26114);
and U27205 (N_27205,N_25664,N_25831);
and U27206 (N_27206,N_25240,N_26154);
nor U27207 (N_27207,N_26119,N_25968);
xor U27208 (N_27208,N_25389,N_25813);
nor U27209 (N_27209,N_26153,N_25390);
or U27210 (N_27210,N_25206,N_25286);
xor U27211 (N_27211,N_25825,N_25440);
nor U27212 (N_27212,N_25585,N_26107);
xnor U27213 (N_27213,N_25335,N_25503);
nand U27214 (N_27214,N_25332,N_25272);
and U27215 (N_27215,N_26188,N_25927);
nor U27216 (N_27216,N_25586,N_26223);
xor U27217 (N_27217,N_25396,N_25849);
and U27218 (N_27218,N_26174,N_25491);
nor U27219 (N_27219,N_25220,N_25624);
and U27220 (N_27220,N_25470,N_26375);
xnor U27221 (N_27221,N_25684,N_26019);
xor U27222 (N_27222,N_25799,N_26370);
xor U27223 (N_27223,N_26230,N_25762);
nand U27224 (N_27224,N_25219,N_26383);
nand U27225 (N_27225,N_25790,N_25858);
nand U27226 (N_27226,N_25840,N_26007);
or U27227 (N_27227,N_26016,N_25205);
nand U27228 (N_27228,N_25657,N_25206);
nand U27229 (N_27229,N_25863,N_25686);
nand U27230 (N_27230,N_26383,N_25516);
xnor U27231 (N_27231,N_25459,N_26165);
and U27232 (N_27232,N_25686,N_25992);
nand U27233 (N_27233,N_26167,N_25624);
xnor U27234 (N_27234,N_25605,N_25402);
and U27235 (N_27235,N_25709,N_25473);
and U27236 (N_27236,N_26091,N_25926);
nand U27237 (N_27237,N_25587,N_25266);
nand U27238 (N_27238,N_25568,N_25794);
nor U27239 (N_27239,N_25993,N_25265);
nor U27240 (N_27240,N_26294,N_26003);
nand U27241 (N_27241,N_25708,N_25800);
xor U27242 (N_27242,N_25509,N_26293);
nand U27243 (N_27243,N_25694,N_25829);
xor U27244 (N_27244,N_25524,N_25403);
nand U27245 (N_27245,N_26246,N_25298);
and U27246 (N_27246,N_25275,N_26395);
nand U27247 (N_27247,N_25264,N_25990);
nand U27248 (N_27248,N_26102,N_25245);
and U27249 (N_27249,N_26071,N_25266);
xor U27250 (N_27250,N_26345,N_25331);
xor U27251 (N_27251,N_25820,N_26179);
xor U27252 (N_27252,N_26394,N_26225);
or U27253 (N_27253,N_25412,N_25223);
xor U27254 (N_27254,N_26357,N_25475);
xnor U27255 (N_27255,N_26209,N_25574);
or U27256 (N_27256,N_26058,N_25667);
or U27257 (N_27257,N_26165,N_25782);
nor U27258 (N_27258,N_25528,N_25513);
xnor U27259 (N_27259,N_26261,N_26155);
or U27260 (N_27260,N_25740,N_26165);
or U27261 (N_27261,N_26202,N_25858);
nor U27262 (N_27262,N_26306,N_26395);
xnor U27263 (N_27263,N_25652,N_25773);
nand U27264 (N_27264,N_25339,N_25437);
nor U27265 (N_27265,N_26046,N_25225);
or U27266 (N_27266,N_25869,N_25718);
and U27267 (N_27267,N_26170,N_26362);
nor U27268 (N_27268,N_26104,N_26336);
and U27269 (N_27269,N_25529,N_26257);
nand U27270 (N_27270,N_25822,N_25776);
or U27271 (N_27271,N_26011,N_25826);
and U27272 (N_27272,N_25326,N_26306);
and U27273 (N_27273,N_26104,N_26284);
and U27274 (N_27274,N_25475,N_26127);
xnor U27275 (N_27275,N_26121,N_25964);
and U27276 (N_27276,N_26076,N_25742);
or U27277 (N_27277,N_26020,N_26382);
nor U27278 (N_27278,N_25208,N_26170);
or U27279 (N_27279,N_26034,N_25289);
nand U27280 (N_27280,N_26399,N_26394);
nand U27281 (N_27281,N_25584,N_25886);
and U27282 (N_27282,N_26210,N_25833);
or U27283 (N_27283,N_25374,N_26378);
and U27284 (N_27284,N_25416,N_25737);
nor U27285 (N_27285,N_25657,N_25471);
nand U27286 (N_27286,N_26098,N_25583);
xor U27287 (N_27287,N_26233,N_25594);
nor U27288 (N_27288,N_25413,N_25559);
nand U27289 (N_27289,N_25679,N_26135);
or U27290 (N_27290,N_25448,N_25592);
nand U27291 (N_27291,N_25308,N_26262);
xnor U27292 (N_27292,N_25332,N_25733);
nor U27293 (N_27293,N_26226,N_26212);
or U27294 (N_27294,N_25550,N_25809);
and U27295 (N_27295,N_25654,N_25243);
xor U27296 (N_27296,N_25830,N_25793);
and U27297 (N_27297,N_26323,N_25603);
and U27298 (N_27298,N_25718,N_25656);
and U27299 (N_27299,N_25351,N_25257);
and U27300 (N_27300,N_25943,N_25864);
or U27301 (N_27301,N_25890,N_26145);
or U27302 (N_27302,N_25966,N_25877);
xor U27303 (N_27303,N_25717,N_25526);
and U27304 (N_27304,N_25857,N_26354);
nor U27305 (N_27305,N_25689,N_25420);
nand U27306 (N_27306,N_26053,N_25353);
and U27307 (N_27307,N_25562,N_25957);
and U27308 (N_27308,N_25654,N_25577);
nand U27309 (N_27309,N_26256,N_26226);
and U27310 (N_27310,N_25947,N_25618);
or U27311 (N_27311,N_25724,N_26182);
and U27312 (N_27312,N_26273,N_25815);
xor U27313 (N_27313,N_25243,N_26194);
nand U27314 (N_27314,N_25314,N_25713);
or U27315 (N_27315,N_25762,N_25608);
or U27316 (N_27316,N_25583,N_25474);
nor U27317 (N_27317,N_26348,N_25446);
and U27318 (N_27318,N_25842,N_25840);
nand U27319 (N_27319,N_25632,N_26125);
or U27320 (N_27320,N_26086,N_25436);
xor U27321 (N_27321,N_25687,N_25821);
and U27322 (N_27322,N_26363,N_25401);
and U27323 (N_27323,N_25494,N_25459);
nor U27324 (N_27324,N_25722,N_26272);
and U27325 (N_27325,N_25577,N_25836);
and U27326 (N_27326,N_25458,N_25527);
xnor U27327 (N_27327,N_25723,N_25466);
and U27328 (N_27328,N_26204,N_26216);
nor U27329 (N_27329,N_26392,N_25593);
xnor U27330 (N_27330,N_26201,N_26041);
or U27331 (N_27331,N_26240,N_26034);
xor U27332 (N_27332,N_26398,N_25677);
nor U27333 (N_27333,N_25298,N_25647);
xor U27334 (N_27334,N_25404,N_26200);
or U27335 (N_27335,N_25764,N_25587);
xor U27336 (N_27336,N_26352,N_25294);
and U27337 (N_27337,N_26117,N_25683);
nand U27338 (N_27338,N_25667,N_25805);
or U27339 (N_27339,N_25389,N_25872);
xor U27340 (N_27340,N_25939,N_26002);
nor U27341 (N_27341,N_26211,N_25709);
nor U27342 (N_27342,N_26140,N_25728);
or U27343 (N_27343,N_26015,N_26359);
and U27344 (N_27344,N_26199,N_25937);
nand U27345 (N_27345,N_25998,N_25981);
nand U27346 (N_27346,N_26089,N_26237);
xnor U27347 (N_27347,N_26301,N_25786);
nor U27348 (N_27348,N_25328,N_26281);
or U27349 (N_27349,N_26241,N_25475);
or U27350 (N_27350,N_26344,N_26051);
and U27351 (N_27351,N_25527,N_25374);
nor U27352 (N_27352,N_26030,N_25517);
xnor U27353 (N_27353,N_26137,N_25870);
nor U27354 (N_27354,N_25985,N_25769);
xnor U27355 (N_27355,N_26385,N_25425);
and U27356 (N_27356,N_26197,N_25484);
and U27357 (N_27357,N_25406,N_25800);
and U27358 (N_27358,N_25501,N_26100);
nor U27359 (N_27359,N_25570,N_26265);
and U27360 (N_27360,N_26201,N_25621);
and U27361 (N_27361,N_26375,N_26260);
xor U27362 (N_27362,N_26332,N_25255);
nand U27363 (N_27363,N_26178,N_25406);
nor U27364 (N_27364,N_25229,N_25544);
nor U27365 (N_27365,N_26029,N_25530);
and U27366 (N_27366,N_26260,N_26217);
nand U27367 (N_27367,N_25749,N_25503);
nand U27368 (N_27368,N_25904,N_26199);
xor U27369 (N_27369,N_26375,N_25328);
nor U27370 (N_27370,N_26267,N_25669);
xor U27371 (N_27371,N_26398,N_25717);
nand U27372 (N_27372,N_25347,N_26174);
and U27373 (N_27373,N_25704,N_25465);
and U27374 (N_27374,N_25565,N_26029);
nor U27375 (N_27375,N_25213,N_26167);
and U27376 (N_27376,N_25472,N_25663);
xnor U27377 (N_27377,N_25460,N_26135);
nand U27378 (N_27378,N_26323,N_25870);
nor U27379 (N_27379,N_25981,N_26049);
nor U27380 (N_27380,N_26211,N_25805);
xor U27381 (N_27381,N_25464,N_25726);
nor U27382 (N_27382,N_26091,N_25942);
and U27383 (N_27383,N_25626,N_25716);
xor U27384 (N_27384,N_26174,N_25705);
and U27385 (N_27385,N_25841,N_26372);
nor U27386 (N_27386,N_26307,N_26221);
nand U27387 (N_27387,N_25733,N_25552);
xnor U27388 (N_27388,N_25280,N_25344);
xor U27389 (N_27389,N_26200,N_25387);
xnor U27390 (N_27390,N_26312,N_26015);
nor U27391 (N_27391,N_26397,N_26007);
and U27392 (N_27392,N_26019,N_25895);
and U27393 (N_27393,N_25719,N_25435);
and U27394 (N_27394,N_25545,N_26051);
nand U27395 (N_27395,N_25336,N_25470);
nor U27396 (N_27396,N_25618,N_25747);
nor U27397 (N_27397,N_25688,N_25606);
and U27398 (N_27398,N_25668,N_26396);
nor U27399 (N_27399,N_25332,N_26032);
or U27400 (N_27400,N_26048,N_25724);
or U27401 (N_27401,N_25827,N_25260);
or U27402 (N_27402,N_25364,N_25813);
nand U27403 (N_27403,N_25257,N_25430);
nand U27404 (N_27404,N_25984,N_26078);
xor U27405 (N_27405,N_26319,N_26243);
or U27406 (N_27406,N_25899,N_25656);
xnor U27407 (N_27407,N_25245,N_25390);
and U27408 (N_27408,N_26110,N_25202);
nand U27409 (N_27409,N_25649,N_25455);
and U27410 (N_27410,N_25419,N_25429);
or U27411 (N_27411,N_25487,N_26138);
nor U27412 (N_27412,N_26343,N_26108);
nor U27413 (N_27413,N_26128,N_25427);
nand U27414 (N_27414,N_25624,N_25210);
and U27415 (N_27415,N_25586,N_25544);
and U27416 (N_27416,N_25553,N_26347);
nor U27417 (N_27417,N_26316,N_26266);
nand U27418 (N_27418,N_25710,N_25591);
xor U27419 (N_27419,N_26314,N_26048);
and U27420 (N_27420,N_26058,N_26173);
nand U27421 (N_27421,N_26142,N_25605);
nand U27422 (N_27422,N_25880,N_26075);
and U27423 (N_27423,N_25433,N_25251);
and U27424 (N_27424,N_26112,N_25971);
xnor U27425 (N_27425,N_25242,N_25787);
or U27426 (N_27426,N_25358,N_25483);
xor U27427 (N_27427,N_26093,N_25669);
or U27428 (N_27428,N_25259,N_26373);
or U27429 (N_27429,N_25897,N_25795);
nor U27430 (N_27430,N_26089,N_25328);
or U27431 (N_27431,N_25492,N_25893);
nor U27432 (N_27432,N_26373,N_25559);
or U27433 (N_27433,N_25605,N_26277);
and U27434 (N_27434,N_25897,N_26115);
nand U27435 (N_27435,N_25879,N_26034);
or U27436 (N_27436,N_25526,N_25637);
xnor U27437 (N_27437,N_25348,N_26046);
or U27438 (N_27438,N_25340,N_25822);
nor U27439 (N_27439,N_25793,N_25905);
nor U27440 (N_27440,N_25236,N_25606);
nor U27441 (N_27441,N_25629,N_25338);
xnor U27442 (N_27442,N_26238,N_25958);
and U27443 (N_27443,N_26113,N_25776);
nor U27444 (N_27444,N_25371,N_25808);
nor U27445 (N_27445,N_26047,N_26107);
xor U27446 (N_27446,N_25485,N_26380);
or U27447 (N_27447,N_25770,N_25980);
nor U27448 (N_27448,N_25348,N_25663);
xnor U27449 (N_27449,N_25746,N_26039);
nor U27450 (N_27450,N_25950,N_25257);
xnor U27451 (N_27451,N_25284,N_25947);
and U27452 (N_27452,N_25437,N_25316);
xnor U27453 (N_27453,N_25521,N_25940);
nand U27454 (N_27454,N_26287,N_25734);
or U27455 (N_27455,N_25283,N_25662);
or U27456 (N_27456,N_25541,N_26315);
nand U27457 (N_27457,N_25859,N_25805);
nand U27458 (N_27458,N_25884,N_25370);
and U27459 (N_27459,N_25364,N_25625);
nand U27460 (N_27460,N_26330,N_25409);
xnor U27461 (N_27461,N_25330,N_26209);
xnor U27462 (N_27462,N_25397,N_26205);
nand U27463 (N_27463,N_26263,N_25635);
xnor U27464 (N_27464,N_25609,N_25928);
nor U27465 (N_27465,N_26000,N_26275);
or U27466 (N_27466,N_25638,N_26157);
and U27467 (N_27467,N_25704,N_26292);
nand U27468 (N_27468,N_25888,N_25445);
nand U27469 (N_27469,N_26205,N_25598);
and U27470 (N_27470,N_25547,N_25252);
nor U27471 (N_27471,N_26384,N_26142);
nor U27472 (N_27472,N_26136,N_25689);
and U27473 (N_27473,N_25528,N_26101);
xor U27474 (N_27474,N_25940,N_25537);
xor U27475 (N_27475,N_25820,N_25664);
or U27476 (N_27476,N_26037,N_25386);
and U27477 (N_27477,N_26024,N_25347);
xnor U27478 (N_27478,N_25883,N_25214);
and U27479 (N_27479,N_25548,N_25592);
nor U27480 (N_27480,N_25339,N_25704);
or U27481 (N_27481,N_26080,N_26016);
nand U27482 (N_27482,N_25792,N_25937);
nand U27483 (N_27483,N_25632,N_25544);
nand U27484 (N_27484,N_26119,N_25354);
nand U27485 (N_27485,N_25894,N_26125);
xnor U27486 (N_27486,N_25958,N_25358);
nand U27487 (N_27487,N_26108,N_25882);
or U27488 (N_27488,N_26309,N_25434);
and U27489 (N_27489,N_25596,N_25903);
xor U27490 (N_27490,N_25240,N_26250);
or U27491 (N_27491,N_25933,N_25838);
nand U27492 (N_27492,N_26339,N_25960);
or U27493 (N_27493,N_26268,N_25830);
and U27494 (N_27494,N_25645,N_26237);
nand U27495 (N_27495,N_26338,N_26357);
nor U27496 (N_27496,N_26045,N_25903);
and U27497 (N_27497,N_25457,N_25727);
xnor U27498 (N_27498,N_26189,N_26155);
nor U27499 (N_27499,N_25687,N_25880);
nand U27500 (N_27500,N_26256,N_25661);
nand U27501 (N_27501,N_25815,N_25472);
or U27502 (N_27502,N_25426,N_26093);
nor U27503 (N_27503,N_25902,N_25613);
nand U27504 (N_27504,N_25574,N_26333);
or U27505 (N_27505,N_25801,N_25563);
and U27506 (N_27506,N_25951,N_25378);
nand U27507 (N_27507,N_25818,N_25953);
nand U27508 (N_27508,N_25302,N_25392);
nand U27509 (N_27509,N_25847,N_25725);
and U27510 (N_27510,N_25879,N_25756);
or U27511 (N_27511,N_25738,N_25380);
xor U27512 (N_27512,N_26268,N_25492);
xnor U27513 (N_27513,N_25461,N_26393);
nand U27514 (N_27514,N_25703,N_26317);
or U27515 (N_27515,N_26256,N_25565);
nor U27516 (N_27516,N_26225,N_26290);
xor U27517 (N_27517,N_25581,N_25950);
xor U27518 (N_27518,N_25933,N_25772);
and U27519 (N_27519,N_26037,N_25765);
and U27520 (N_27520,N_26175,N_25645);
nand U27521 (N_27521,N_25995,N_25395);
nand U27522 (N_27522,N_26363,N_26377);
nand U27523 (N_27523,N_25905,N_26324);
nor U27524 (N_27524,N_25454,N_25946);
and U27525 (N_27525,N_25500,N_26196);
xor U27526 (N_27526,N_25771,N_25717);
nor U27527 (N_27527,N_26169,N_25698);
nor U27528 (N_27528,N_26195,N_26077);
xor U27529 (N_27529,N_25503,N_25461);
nor U27530 (N_27530,N_25738,N_25267);
or U27531 (N_27531,N_25557,N_25618);
xnor U27532 (N_27532,N_25801,N_25666);
and U27533 (N_27533,N_25622,N_25759);
and U27534 (N_27534,N_26311,N_25864);
nor U27535 (N_27535,N_25966,N_25764);
or U27536 (N_27536,N_25596,N_25725);
nor U27537 (N_27537,N_25281,N_26149);
nand U27538 (N_27538,N_25511,N_25746);
nor U27539 (N_27539,N_25726,N_25923);
nor U27540 (N_27540,N_25260,N_26382);
or U27541 (N_27541,N_26088,N_25752);
or U27542 (N_27542,N_26384,N_25271);
xor U27543 (N_27543,N_25329,N_25474);
nand U27544 (N_27544,N_25740,N_26389);
or U27545 (N_27545,N_26135,N_26100);
xnor U27546 (N_27546,N_25397,N_25634);
and U27547 (N_27547,N_26303,N_26234);
nand U27548 (N_27548,N_25434,N_25342);
xnor U27549 (N_27549,N_25831,N_25917);
nand U27550 (N_27550,N_25729,N_25959);
and U27551 (N_27551,N_26288,N_25291);
and U27552 (N_27552,N_25281,N_25578);
nor U27553 (N_27553,N_25788,N_25366);
nor U27554 (N_27554,N_26065,N_25509);
nand U27555 (N_27555,N_25565,N_25271);
nand U27556 (N_27556,N_25788,N_26061);
or U27557 (N_27557,N_25799,N_26214);
nand U27558 (N_27558,N_25601,N_25530);
nand U27559 (N_27559,N_25435,N_25575);
nor U27560 (N_27560,N_26180,N_25925);
or U27561 (N_27561,N_25431,N_25587);
or U27562 (N_27562,N_25328,N_26001);
or U27563 (N_27563,N_25669,N_25815);
and U27564 (N_27564,N_26340,N_26234);
and U27565 (N_27565,N_25415,N_25746);
and U27566 (N_27566,N_26336,N_25956);
nand U27567 (N_27567,N_25298,N_25664);
nor U27568 (N_27568,N_25503,N_26336);
xor U27569 (N_27569,N_26107,N_25479);
nor U27570 (N_27570,N_26357,N_26065);
and U27571 (N_27571,N_26084,N_25763);
or U27572 (N_27572,N_25412,N_25314);
xor U27573 (N_27573,N_26373,N_26326);
nor U27574 (N_27574,N_26391,N_25593);
nand U27575 (N_27575,N_25201,N_25858);
and U27576 (N_27576,N_25221,N_26233);
nor U27577 (N_27577,N_26044,N_25937);
xor U27578 (N_27578,N_25994,N_25814);
nor U27579 (N_27579,N_25431,N_25416);
or U27580 (N_27580,N_25698,N_25793);
or U27581 (N_27581,N_25271,N_25598);
xor U27582 (N_27582,N_25405,N_25751);
and U27583 (N_27583,N_26220,N_25817);
nor U27584 (N_27584,N_25225,N_26223);
or U27585 (N_27585,N_26275,N_25331);
or U27586 (N_27586,N_25994,N_25499);
and U27587 (N_27587,N_26219,N_26227);
or U27588 (N_27588,N_25268,N_25464);
xnor U27589 (N_27589,N_25990,N_25928);
nand U27590 (N_27590,N_26372,N_25890);
nand U27591 (N_27591,N_25622,N_25277);
xnor U27592 (N_27592,N_26087,N_26108);
nand U27593 (N_27593,N_25727,N_25599);
nand U27594 (N_27594,N_26293,N_26166);
xor U27595 (N_27595,N_26335,N_25642);
and U27596 (N_27596,N_25988,N_26018);
xnor U27597 (N_27597,N_25696,N_25537);
or U27598 (N_27598,N_26205,N_25655);
xnor U27599 (N_27599,N_25391,N_26106);
nor U27600 (N_27600,N_27392,N_26513);
or U27601 (N_27601,N_27191,N_26765);
or U27602 (N_27602,N_27314,N_26533);
nand U27603 (N_27603,N_26708,N_26622);
or U27604 (N_27604,N_26406,N_26656);
nor U27605 (N_27605,N_26947,N_26985);
nand U27606 (N_27606,N_26600,N_26537);
or U27607 (N_27607,N_26788,N_26632);
or U27608 (N_27608,N_27576,N_26847);
nor U27609 (N_27609,N_27172,N_27410);
xnor U27610 (N_27610,N_27484,N_27434);
and U27611 (N_27611,N_27458,N_26450);
and U27612 (N_27612,N_27217,N_26785);
or U27613 (N_27613,N_27194,N_26875);
xor U27614 (N_27614,N_26799,N_27534);
and U27615 (N_27615,N_26786,N_26640);
and U27616 (N_27616,N_27402,N_27425);
or U27617 (N_27617,N_26635,N_26978);
or U27618 (N_27618,N_26793,N_27090);
nor U27619 (N_27619,N_26721,N_26924);
xor U27620 (N_27620,N_26581,N_26912);
nor U27621 (N_27621,N_27127,N_27150);
nor U27622 (N_27622,N_26869,N_26745);
nor U27623 (N_27623,N_27240,N_27334);
xor U27624 (N_27624,N_26530,N_26698);
and U27625 (N_27625,N_26454,N_26510);
xnor U27626 (N_27626,N_26848,N_27514);
xor U27627 (N_27627,N_26752,N_27417);
or U27628 (N_27628,N_26538,N_27498);
or U27629 (N_27629,N_27069,N_27506);
nor U27630 (N_27630,N_27561,N_27259);
and U27631 (N_27631,N_26994,N_26572);
nor U27632 (N_27632,N_26954,N_27221);
nand U27633 (N_27633,N_26951,N_27012);
or U27634 (N_27634,N_27236,N_26753);
nand U27635 (N_27635,N_27253,N_26995);
or U27636 (N_27636,N_27547,N_26644);
xnor U27637 (N_27637,N_27360,N_27499);
or U27638 (N_27638,N_27429,N_27503);
nand U27639 (N_27639,N_26589,N_26509);
nand U27640 (N_27640,N_26953,N_26929);
or U27641 (N_27641,N_27214,N_27423);
xnor U27642 (N_27642,N_26700,N_27120);
xnor U27643 (N_27643,N_27256,N_27472);
or U27644 (N_27644,N_27368,N_26996);
nand U27645 (N_27645,N_26420,N_27473);
nand U27646 (N_27646,N_26901,N_27289);
nand U27647 (N_27647,N_27528,N_27571);
and U27648 (N_27648,N_27496,N_26933);
xor U27649 (N_27649,N_26828,N_26737);
nand U27650 (N_27650,N_26521,N_26870);
and U27651 (N_27651,N_27193,N_26651);
xnor U27652 (N_27652,N_26895,N_26902);
nand U27653 (N_27653,N_26527,N_26528);
xor U27654 (N_27654,N_27273,N_26952);
nor U27655 (N_27655,N_27470,N_26990);
and U27656 (N_27656,N_26487,N_27167);
xor U27657 (N_27657,N_26976,N_26941);
xor U27658 (N_27658,N_27296,N_27445);
and U27659 (N_27659,N_26403,N_26404);
nor U27660 (N_27660,N_26891,N_27076);
and U27661 (N_27661,N_26775,N_27192);
and U27662 (N_27662,N_26770,N_26546);
nor U27663 (N_27663,N_26673,N_26787);
xor U27664 (N_27664,N_27269,N_26879);
or U27665 (N_27665,N_27451,N_27482);
or U27666 (N_27666,N_26865,N_27294);
nand U27667 (N_27667,N_26439,N_26919);
or U27668 (N_27668,N_27138,N_27001);
xnor U27669 (N_27669,N_26411,N_26922);
or U27670 (N_27670,N_26518,N_26429);
nand U27671 (N_27671,N_27276,N_27185);
xor U27672 (N_27672,N_26970,N_26629);
and U27673 (N_27673,N_27340,N_27375);
xnor U27674 (N_27674,N_27320,N_26498);
and U27675 (N_27675,N_26474,N_27306);
nand U27676 (N_27676,N_27311,N_27208);
nand U27677 (N_27677,N_26797,N_26664);
nor U27678 (N_27678,N_26423,N_26713);
and U27679 (N_27679,N_26961,N_27501);
or U27680 (N_27680,N_26586,N_27045);
or U27681 (N_27681,N_26531,N_26419);
and U27682 (N_27682,N_27546,N_26832);
nand U27683 (N_27683,N_27050,N_26571);
or U27684 (N_27684,N_27562,N_27421);
and U27685 (N_27685,N_26926,N_26611);
and U27686 (N_27686,N_26499,N_27517);
nor U27687 (N_27687,N_27397,N_26490);
or U27688 (N_27688,N_27080,N_27513);
and U27689 (N_27689,N_26637,N_26859);
nand U27690 (N_27690,N_27223,N_27394);
nand U27691 (N_27691,N_26433,N_27309);
and U27692 (N_27692,N_27188,N_27122);
xnor U27693 (N_27693,N_26905,N_27074);
and U27694 (N_27694,N_27084,N_27516);
or U27695 (N_27695,N_26957,N_26437);
and U27696 (N_27696,N_26465,N_27131);
nand U27697 (N_27697,N_27021,N_27545);
nor U27698 (N_27698,N_26723,N_27293);
and U27699 (N_27699,N_26790,N_27333);
and U27700 (N_27700,N_27290,N_26958);
nor U27701 (N_27701,N_27175,N_26407);
and U27702 (N_27702,N_27366,N_27526);
nor U27703 (N_27703,N_26885,N_26772);
nor U27704 (N_27704,N_27485,N_27005);
and U27705 (N_27705,N_27380,N_27181);
and U27706 (N_27706,N_26892,N_27089);
or U27707 (N_27707,N_27251,N_26712);
or U27708 (N_27708,N_27298,N_27108);
nor U27709 (N_27709,N_27180,N_27572);
or U27710 (N_27710,N_27075,N_27337);
nor U27711 (N_27711,N_27107,N_26678);
nand U27712 (N_27712,N_27478,N_26615);
or U27713 (N_27713,N_26925,N_26727);
or U27714 (N_27714,N_27072,N_27464);
or U27715 (N_27715,N_27250,N_27406);
xnor U27716 (N_27716,N_26565,N_26866);
nand U27717 (N_27717,N_27297,N_26583);
nand U27718 (N_27718,N_27169,N_26427);
xor U27719 (N_27719,N_26401,N_26967);
nor U27720 (N_27720,N_27207,N_26900);
and U27721 (N_27721,N_26872,N_27153);
nand U27722 (N_27722,N_26762,N_27411);
xnor U27723 (N_27723,N_26956,N_26830);
nand U27724 (N_27724,N_26883,N_26938);
and U27725 (N_27725,N_27047,N_26541);
xor U27726 (N_27726,N_27585,N_27344);
xnor U27727 (N_27727,N_26795,N_27044);
and U27728 (N_27728,N_26648,N_26858);
nor U27729 (N_27729,N_26681,N_26677);
nor U27730 (N_27730,N_26544,N_26945);
xnor U27731 (N_27731,N_27203,N_26857);
xnor U27732 (N_27732,N_26837,N_26558);
xor U27733 (N_27733,N_26587,N_27178);
and U27734 (N_27734,N_27227,N_27575);
and U27735 (N_27735,N_26405,N_26861);
nand U27736 (N_27736,N_27565,N_27201);
nand U27737 (N_27737,N_27324,N_27121);
nand U27738 (N_27738,N_27128,N_26973);
nor U27739 (N_27739,N_27145,N_27525);
and U27740 (N_27740,N_26594,N_26524);
nor U27741 (N_27741,N_26687,N_26626);
nor U27742 (N_27742,N_27522,N_26868);
nor U27743 (N_27743,N_27376,N_26460);
or U27744 (N_27744,N_26904,N_27568);
and U27745 (N_27745,N_26710,N_27307);
and U27746 (N_27746,N_27031,N_26576);
nor U27747 (N_27747,N_26827,N_26817);
or U27748 (N_27748,N_27384,N_27286);
nor U27749 (N_27749,N_26841,N_27596);
xor U27750 (N_27750,N_27291,N_27468);
nand U27751 (N_27751,N_27186,N_26694);
nand U27752 (N_27752,N_26466,N_26998);
nand U27753 (N_27753,N_27404,N_26823);
and U27754 (N_27754,N_27148,N_26562);
xnor U27755 (N_27755,N_27039,N_27454);
or U27756 (N_27756,N_27521,N_26934);
nand U27757 (N_27757,N_27532,N_26894);
xnor U27758 (N_27758,N_27002,N_27594);
xor U27759 (N_27759,N_26602,N_26556);
or U27760 (N_27760,N_26864,N_27530);
nand U27761 (N_27761,N_27364,N_26627);
nor U27762 (N_27762,N_27379,N_26500);
and U27763 (N_27763,N_27209,N_27117);
nor U27764 (N_27764,N_26819,N_26728);
nor U27765 (N_27765,N_27246,N_27233);
and U27766 (N_27766,N_27502,N_26605);
and U27767 (N_27767,N_27556,N_26824);
and U27768 (N_27768,N_27222,N_26932);
xor U27769 (N_27769,N_26993,N_26791);
nand U27770 (N_27770,N_26624,N_26833);
or U27771 (N_27771,N_27096,N_26741);
nand U27772 (N_27772,N_26969,N_26472);
or U27773 (N_27773,N_26944,N_26689);
nand U27774 (N_27774,N_26997,N_26580);
or U27775 (N_27775,N_27056,N_27064);
nor U27776 (N_27776,N_27539,N_27059);
and U27777 (N_27777,N_26732,N_26874);
nand U27778 (N_27778,N_26992,N_26748);
xor U27779 (N_27779,N_27126,N_26489);
and U27780 (N_27780,N_27137,N_26886);
xor U27781 (N_27781,N_26884,N_27537);
xor U27782 (N_27782,N_26647,N_26504);
nand U27783 (N_27783,N_26796,N_26746);
nand U27784 (N_27784,N_27563,N_26826);
xor U27785 (N_27785,N_26496,N_26692);
nor U27786 (N_27786,N_26764,N_26598);
or U27787 (N_27787,N_26804,N_27319);
and U27788 (N_27788,N_26890,N_27474);
nand U27789 (N_27789,N_26669,N_27164);
xor U27790 (N_27790,N_26942,N_27010);
nor U27791 (N_27791,N_27582,N_26989);
and U27792 (N_27792,N_26485,N_26812);
and U27793 (N_27793,N_26911,N_26747);
and U27794 (N_27794,N_26876,N_27331);
xnor U27795 (N_27795,N_27466,N_26421);
nor U27796 (N_27796,N_26610,N_27141);
and U27797 (N_27797,N_27447,N_26853);
nor U27798 (N_27798,N_26761,N_27373);
nand U27799 (N_27799,N_27544,N_26452);
xor U27800 (N_27800,N_27285,N_27538);
xor U27801 (N_27801,N_26554,N_27100);
nor U27802 (N_27802,N_27341,N_26715);
nor U27803 (N_27803,N_27023,N_26693);
and U27804 (N_27804,N_27431,N_27370);
nor U27805 (N_27805,N_27212,N_27157);
nand U27806 (N_27806,N_27367,N_26688);
nand U27807 (N_27807,N_27211,N_27261);
or U27808 (N_27808,N_26609,N_27439);
nand U27809 (N_27809,N_27555,N_26968);
and U27810 (N_27810,N_27430,N_26893);
nand U27811 (N_27811,N_27265,N_27094);
xnor U27812 (N_27812,N_27197,N_26735);
nand U27813 (N_27813,N_27409,N_26523);
xor U27814 (N_27814,N_26810,N_27151);
or U27815 (N_27815,N_26691,N_27550);
and U27816 (N_27816,N_27245,N_26914);
and U27817 (N_27817,N_27398,N_27529);
nor U27818 (N_27818,N_26671,N_26940);
xnor U27819 (N_27819,N_27554,N_27266);
nor U27820 (N_27820,N_27213,N_26604);
nand U27821 (N_27821,N_27424,N_26878);
nor U27822 (N_27822,N_26749,N_27486);
or U27823 (N_27823,N_26972,N_27548);
and U27824 (N_27824,N_27016,N_26494);
or U27825 (N_27825,N_26923,N_26779);
nor U27826 (N_27826,N_26540,N_27543);
and U27827 (N_27827,N_26674,N_26711);
or U27828 (N_27828,N_26468,N_27357);
nor U27829 (N_27829,N_27280,N_26570);
or U27830 (N_27830,N_27219,N_27237);
nand U27831 (N_27831,N_27351,N_26578);
nand U27832 (N_27832,N_27564,N_27598);
nand U27833 (N_27833,N_26943,N_26739);
or U27834 (N_27834,N_27098,N_27196);
or U27835 (N_27835,N_26559,N_26734);
and U27836 (N_27836,N_26939,N_26966);
xor U27837 (N_27837,N_26470,N_26809);
and U27838 (N_27838,N_27457,N_26888);
xnor U27839 (N_27839,N_26769,N_27267);
xor U27840 (N_27840,N_27224,N_26596);
nand U27841 (N_27841,N_27102,N_27020);
or U27842 (N_27842,N_26442,N_27007);
nand U27843 (N_27843,N_26740,N_27279);
nor U27844 (N_27844,N_26755,N_27216);
nor U27845 (N_27845,N_27284,N_27133);
xnor U27846 (N_27846,N_27132,N_26738);
or U27847 (N_27847,N_27113,N_27463);
nor U27848 (N_27848,N_26999,N_27046);
and U27849 (N_27849,N_26873,N_27597);
nand U27850 (N_27850,N_26616,N_26843);
nand U27851 (N_27851,N_26814,N_27385);
and U27852 (N_27852,N_26657,N_27130);
or U27853 (N_27853,N_27495,N_26601);
and U27854 (N_27854,N_26898,N_27308);
or U27855 (N_27855,N_26889,N_26816);
nand U27856 (N_27856,N_27432,N_27415);
nand U27857 (N_27857,N_26806,N_27436);
nand U27858 (N_27858,N_27347,N_27025);
nor U27859 (N_27859,N_27206,N_27389);
nand U27860 (N_27860,N_26758,N_27234);
or U27861 (N_27861,N_27275,N_26836);
nand U27862 (N_27862,N_26493,N_26424);
xor U27863 (N_27863,N_26621,N_27299);
or U27864 (N_27864,N_27058,N_26974);
and U27865 (N_27865,N_27026,N_26906);
and U27866 (N_27866,N_27184,N_26545);
xor U27867 (N_27867,N_26516,N_27330);
and U27868 (N_27868,N_26881,N_26630);
or U27869 (N_27869,N_27471,N_26931);
nor U27870 (N_27870,N_27238,N_27099);
and U27871 (N_27871,N_27479,N_27317);
or U27872 (N_27872,N_26410,N_27358);
nor U27873 (N_27873,N_26851,N_26402);
xnor U27874 (N_27874,N_27179,N_26773);
nor U27875 (N_27875,N_27242,N_26766);
and U27876 (N_27876,N_27119,N_27264);
nand U27877 (N_27877,N_27321,N_26896);
and U27878 (N_27878,N_27362,N_26899);
xnor U27879 (N_27879,N_27599,N_26459);
or U27880 (N_27880,N_26486,N_27450);
or U27881 (N_27881,N_27190,N_26502);
nor U27882 (N_27882,N_26654,N_26453);
or U27883 (N_27883,N_26451,N_27028);
nor U27884 (N_27884,N_26921,N_27262);
and U27885 (N_27885,N_26449,N_27052);
and U27886 (N_27886,N_26930,N_26432);
or U27887 (N_27887,N_27302,N_26834);
nor U27888 (N_27888,N_27204,N_26573);
xor U27889 (N_27889,N_27412,N_26461);
nor U27890 (N_27890,N_26794,N_27480);
and U27891 (N_27891,N_27263,N_27159);
xor U27892 (N_27892,N_27004,N_26927);
and U27893 (N_27893,N_26699,N_27490);
or U27894 (N_27894,N_27115,N_26628);
and U27895 (N_27895,N_27006,N_27042);
and U27896 (N_27896,N_27249,N_26917);
nand U27897 (N_27897,N_26910,N_27318);
nor U27898 (N_27898,N_26962,N_27198);
nand U27899 (N_27899,N_26431,N_26807);
nand U27900 (N_27900,N_27442,N_27063);
xnor U27901 (N_27901,N_26488,N_27523);
and U27902 (N_27902,N_26641,N_26763);
nand U27903 (N_27903,N_27413,N_26959);
nor U27904 (N_27904,N_26636,N_27504);
nor U27905 (N_27905,N_27325,N_27166);
nand U27906 (N_27906,N_27062,N_26903);
nand U27907 (N_27907,N_26719,N_27034);
or U27908 (N_27908,N_26789,N_26520);
and U27909 (N_27909,N_26638,N_26760);
and U27910 (N_27910,N_27027,N_27032);
and U27911 (N_27911,N_26682,N_26606);
nand U27912 (N_27912,N_27114,N_27123);
or U27913 (N_27913,N_27595,N_27374);
nand U27914 (N_27914,N_27313,N_27553);
or U27915 (N_27915,N_27218,N_26588);
xor U27916 (N_27916,N_27158,N_27066);
or U27917 (N_27917,N_26986,N_26491);
nor U27918 (N_27918,N_27041,N_27510);
or U27919 (N_27919,N_26730,N_26800);
or U27920 (N_27920,N_26733,N_26643);
or U27921 (N_27921,N_27228,N_27149);
or U27922 (N_27922,N_26582,N_26482);
and U27923 (N_27923,N_27252,N_27139);
or U27924 (N_27924,N_27549,N_26553);
nand U27925 (N_27925,N_26477,N_27241);
and U27926 (N_27926,N_26667,N_27356);
or U27927 (N_27927,N_27051,N_27215);
and U27928 (N_27928,N_26983,N_27282);
and U27929 (N_27929,N_27584,N_27176);
nor U27930 (N_27930,N_27414,N_26532);
and U27931 (N_27931,N_27444,N_27390);
xnor U27932 (N_27932,N_27254,N_26620);
or U27933 (N_27933,N_26820,N_26652);
xor U27934 (N_27934,N_27422,N_27029);
and U27935 (N_27935,N_27230,N_26754);
nor U27936 (N_27936,N_27581,N_26808);
nor U27937 (N_27937,N_26850,N_27182);
nand U27938 (N_27938,N_26503,N_26928);
or U27939 (N_27939,N_26463,N_27391);
nor U27940 (N_27940,N_26655,N_27533);
or U27941 (N_27941,N_27578,N_26849);
xnor U27942 (N_27942,N_26436,N_27465);
or U27943 (N_27943,N_26547,N_27512);
xnor U27944 (N_27944,N_26412,N_27061);
xnor U27945 (N_27945,N_27152,N_26457);
xnor U27946 (N_27946,N_27350,N_26846);
or U27947 (N_27947,N_27082,N_26455);
xnor U27948 (N_27948,N_27205,N_27287);
nand U27949 (N_27949,N_27443,N_26703);
nor U27950 (N_27950,N_27382,N_26430);
xnor U27951 (N_27951,N_26963,N_27336);
nand U27952 (N_27952,N_27093,N_27569);
or U27953 (N_27953,N_27500,N_26722);
nand U27954 (N_27954,N_26511,N_27369);
xnor U27955 (N_27955,N_27483,N_26913);
nor U27956 (N_27956,N_27277,N_26650);
or U27957 (N_27957,N_26844,N_27377);
nor U27958 (N_27958,N_26731,N_27271);
and U27959 (N_27959,N_26702,N_27455);
and U27960 (N_27960,N_27146,N_27541);
nor U27961 (N_27961,N_26592,N_26639);
or U27962 (N_27962,N_27278,N_26668);
or U27963 (N_27963,N_26774,N_26633);
nand U27964 (N_27964,N_27449,N_27140);
nand U27965 (N_27965,N_27144,N_26991);
and U27966 (N_27966,N_26566,N_27511);
nand U27967 (N_27967,N_26977,N_26550);
or U27968 (N_27968,N_27124,N_27452);
xor U27969 (N_27969,N_26458,N_26909);
nor U27970 (N_27970,N_27590,N_27393);
and U27971 (N_27971,N_27327,N_26464);
nand U27972 (N_27972,N_27118,N_27258);
xor U27973 (N_27973,N_26937,N_27303);
or U27974 (N_27974,N_27078,N_27038);
and U27975 (N_27975,N_26949,N_27349);
or U27976 (N_27976,N_27339,N_27505);
xnor U27977 (N_27977,N_27009,N_26574);
nor U27978 (N_27978,N_26623,N_27428);
or U27979 (N_27979,N_26670,N_27365);
xnor U27980 (N_27980,N_26736,N_26984);
and U27981 (N_27981,N_27515,N_27247);
xnor U27982 (N_27982,N_26805,N_26936);
and U27983 (N_27983,N_26663,N_27035);
or U27984 (N_27984,N_27519,N_26982);
xor U27985 (N_27985,N_26975,N_26417);
and U27986 (N_27986,N_26916,N_27295);
and U27987 (N_27987,N_27110,N_26852);
and U27988 (N_27988,N_26987,N_27426);
nor U27989 (N_27989,N_26517,N_26508);
nand U27990 (N_27990,N_26776,N_27387);
nand U27991 (N_27991,N_27405,N_27156);
and U27992 (N_27992,N_27372,N_27248);
xnor U27993 (N_27993,N_27155,N_26557);
and U27994 (N_27994,N_27577,N_27260);
nand U27995 (N_27995,N_27408,N_26686);
xor U27996 (N_27996,N_27135,N_26751);
or U27997 (N_27997,N_27288,N_26979);
or U27998 (N_27998,N_27040,N_27085);
nand U27999 (N_27999,N_26676,N_26863);
nor U28000 (N_28000,N_26434,N_26707);
xnor U28001 (N_28001,N_27573,N_27520);
and U28002 (N_28002,N_27559,N_27070);
or U28003 (N_28003,N_27147,N_27416);
or U28004 (N_28004,N_27048,N_27202);
nor U28005 (N_28005,N_26416,N_27022);
nor U28006 (N_28006,N_26897,N_26778);
nor U28007 (N_28007,N_26918,N_26591);
and U28008 (N_28008,N_26642,N_27557);
nand U28009 (N_28009,N_26679,N_26955);
or U28010 (N_28010,N_27491,N_26475);
nand U28011 (N_28011,N_26448,N_27312);
xnor U28012 (N_28012,N_27477,N_27332);
or U28013 (N_28013,N_26683,N_26709);
nor U28014 (N_28014,N_27551,N_26479);
xor U28015 (N_28015,N_26780,N_27446);
and U28016 (N_28016,N_27077,N_26696);
xnor U28017 (N_28017,N_26980,N_26418);
or U28018 (N_28018,N_26441,N_26965);
xnor U28019 (N_28019,N_27587,N_26704);
nand U28020 (N_28020,N_27014,N_26782);
nor U28021 (N_28021,N_26666,N_26428);
nand U28022 (N_28022,N_27328,N_27343);
xnor U28023 (N_28023,N_26880,N_27030);
nor U28024 (N_28024,N_26815,N_26759);
and U28025 (N_28025,N_27283,N_27225);
xnor U28026 (N_28026,N_27109,N_26792);
or U28027 (N_28027,N_27154,N_27560);
xnor U28028 (N_28028,N_26855,N_26964);
xor U28029 (N_28029,N_26535,N_26481);
nor U28030 (N_28030,N_27106,N_26658);
nand U28031 (N_28031,N_26435,N_26882);
xor U28032 (N_28032,N_27257,N_26484);
nor U28033 (N_28033,N_26645,N_27338);
nand U28034 (N_28034,N_26767,N_26569);
and U28035 (N_28035,N_27015,N_27593);
or U28036 (N_28036,N_26946,N_26539);
or U28037 (N_28037,N_26552,N_27494);
xnor U28038 (N_28038,N_26564,N_26744);
nor U28039 (N_28039,N_26413,N_26920);
or U28040 (N_28040,N_27535,N_27111);
or U28041 (N_28041,N_27440,N_27427);
or U28042 (N_28042,N_27087,N_26501);
xnor U28043 (N_28043,N_27104,N_27177);
xnor U28044 (N_28044,N_27274,N_26634);
nor U28045 (N_28045,N_26818,N_27588);
and U28046 (N_28046,N_27460,N_27243);
and U28047 (N_28047,N_26473,N_26476);
and U28048 (N_28048,N_27136,N_27335);
xor U28049 (N_28049,N_26618,N_26811);
or U28050 (N_28050,N_26801,N_26821);
or U28051 (N_28051,N_27013,N_26988);
xnor U28052 (N_28052,N_26716,N_26750);
xnor U28053 (N_28053,N_26597,N_27235);
or U28054 (N_28054,N_26577,N_27361);
or U28055 (N_28055,N_26768,N_26724);
xnor U28056 (N_28056,N_26529,N_27315);
or U28057 (N_28057,N_26515,N_27011);
nand U28058 (N_28058,N_26462,N_27527);
xnor U28059 (N_28059,N_26860,N_27101);
nand U28060 (N_28060,N_27542,N_26948);
and U28061 (N_28061,N_26555,N_26608);
and U28062 (N_28062,N_27210,N_26725);
and U28063 (N_28063,N_27453,N_26697);
and U28064 (N_28064,N_27068,N_27438);
xnor U28065 (N_28065,N_27170,N_26612);
nor U28066 (N_28066,N_27226,N_26695);
xor U28067 (N_28067,N_27008,N_27165);
nor U28068 (N_28068,N_27270,N_26614);
and U28069 (N_28069,N_26567,N_26497);
nor U28070 (N_28070,N_27049,N_27518);
xnor U28071 (N_28071,N_26512,N_27054);
and U28072 (N_28072,N_26777,N_27088);
nand U28073 (N_28073,N_26659,N_26593);
or U28074 (N_28074,N_27189,N_26492);
xnor U28075 (N_28075,N_27433,N_27345);
nand U28076 (N_28076,N_27395,N_27129);
nand U28077 (N_28077,N_26590,N_27509);
xnor U28078 (N_28078,N_26471,N_27272);
nor U28079 (N_28079,N_27134,N_27301);
nor U28080 (N_28080,N_27469,N_26579);
nand U28081 (N_28081,N_26714,N_27043);
nor U28082 (N_28082,N_27401,N_27079);
xnor U28083 (N_28083,N_26798,N_27017);
or U28084 (N_28084,N_27057,N_27419);
xor U28085 (N_28085,N_26575,N_27037);
or U28086 (N_28086,N_26757,N_26829);
and U28087 (N_28087,N_27323,N_27329);
nand U28088 (N_28088,N_27036,N_27195);
xnor U28089 (N_28089,N_27310,N_27018);
xnor U28090 (N_28090,N_26584,N_26469);
xnor U28091 (N_28091,N_27024,N_26595);
nand U28092 (N_28092,N_26854,N_27160);
and U28093 (N_28093,N_26783,N_26915);
and U28094 (N_28094,N_27232,N_26603);
xor U28095 (N_28095,N_26446,N_27591);
and U28096 (N_28096,N_27407,N_26646);
or U28097 (N_28097,N_27073,N_27352);
xor U28098 (N_28098,N_27383,N_26981);
nor U28099 (N_28099,N_26835,N_26525);
and U28100 (N_28100,N_27229,N_26526);
and U28101 (N_28101,N_26718,N_27200);
nand U28102 (N_28102,N_27570,N_26720);
and U28103 (N_28103,N_27019,N_26548);
or U28104 (N_28104,N_26551,N_26685);
nor U28105 (N_28105,N_27448,N_27354);
or U28106 (N_28106,N_26831,N_27566);
and U28107 (N_28107,N_26701,N_26649);
nand U28108 (N_28108,N_27183,N_26680);
xnor U28109 (N_28109,N_26617,N_26867);
nor U28110 (N_28110,N_26507,N_26661);
and U28111 (N_28111,N_27244,N_26771);
or U28112 (N_28112,N_27531,N_26480);
and U28113 (N_28113,N_26425,N_26887);
nand U28114 (N_28114,N_26822,N_27199);
nor U28115 (N_28115,N_27467,N_26506);
xor U28116 (N_28116,N_26729,N_26549);
nand U28117 (N_28117,N_27396,N_27508);
xnor U28118 (N_28118,N_27095,N_27187);
and U28119 (N_28119,N_27060,N_26426);
nor U28120 (N_28120,N_27355,N_26563);
and U28121 (N_28121,N_26907,N_27388);
and U28122 (N_28122,N_26690,N_27300);
nor U28123 (N_28123,N_26877,N_27507);
nor U28124 (N_28124,N_27418,N_27524);
and U28125 (N_28125,N_27371,N_27441);
nand U28126 (N_28126,N_27255,N_27220);
and U28127 (N_28127,N_27116,N_26613);
nor U28128 (N_28128,N_27558,N_27281);
nor U28129 (N_28129,N_26825,N_27459);
or U28130 (N_28130,N_26440,N_27053);
or U28131 (N_28131,N_27378,N_26781);
nor U28132 (N_28132,N_27348,N_27497);
and U28133 (N_28133,N_27143,N_27586);
nand U28134 (N_28134,N_27125,N_27536);
or U28135 (N_28135,N_27488,N_26478);
or U28136 (N_28136,N_26756,N_27000);
xnor U28137 (N_28137,N_26971,N_26675);
nor U28138 (N_28138,N_27487,N_26585);
nand U28139 (N_28139,N_26908,N_26813);
xor U28140 (N_28140,N_26717,N_26534);
and U28141 (N_28141,N_26619,N_27475);
or U28142 (N_28142,N_27574,N_27363);
nor U28143 (N_28143,N_26684,N_27071);
and U28144 (N_28144,N_27003,N_27092);
nand U28145 (N_28145,N_27579,N_27161);
xor U28146 (N_28146,N_26514,N_27305);
xnor U28147 (N_28147,N_26742,N_26653);
nand U28148 (N_28148,N_27359,N_26802);
or U28149 (N_28149,N_27173,N_27105);
nor U28150 (N_28150,N_26803,N_26561);
or U28151 (N_28151,N_27326,N_27055);
xor U28152 (N_28152,N_26522,N_26660);
nor U28153 (N_28153,N_27481,N_26560);
and U28154 (N_28154,N_26467,N_27083);
nor U28155 (N_28155,N_27476,N_27580);
xor U28156 (N_28156,N_26607,N_26409);
nand U28157 (N_28157,N_26495,N_27097);
xor U28158 (N_28158,N_27346,N_26568);
or U28159 (N_28159,N_27489,N_27552);
nor U28160 (N_28160,N_27589,N_27112);
nand U28161 (N_28161,N_26543,N_26444);
and U28162 (N_28162,N_26415,N_26599);
or U28163 (N_28163,N_27142,N_26456);
or U28164 (N_28164,N_27420,N_26536);
xnor U28165 (N_28165,N_27067,N_26414);
nor U28166 (N_28166,N_27353,N_26784);
xor U28167 (N_28167,N_26706,N_26935);
nand U28168 (N_28168,N_27342,N_27033);
nor U28169 (N_28169,N_26842,N_26672);
nor U28170 (N_28170,N_27493,N_26856);
or U28171 (N_28171,N_26422,N_26871);
or U28172 (N_28172,N_27583,N_27168);
and U28173 (N_28173,N_26665,N_27171);
xnor U28174 (N_28174,N_26443,N_27304);
xnor U28175 (N_28175,N_27316,N_27174);
and U28176 (N_28176,N_26519,N_27461);
xor U28177 (N_28177,N_27462,N_26542);
or U28178 (N_28178,N_27163,N_27381);
nor U28179 (N_28179,N_26505,N_26408);
nand U28180 (N_28180,N_26625,N_27086);
nor U28181 (N_28181,N_27403,N_27567);
xnor U28182 (N_28182,N_27456,N_27231);
nand U28183 (N_28183,N_26438,N_26840);
xor U28184 (N_28184,N_26838,N_26845);
or U28185 (N_28185,N_26445,N_27162);
nor U28186 (N_28186,N_27239,N_27103);
nor U28187 (N_28187,N_26447,N_26950);
xor U28188 (N_28188,N_27268,N_27592);
xnor U28189 (N_28189,N_27065,N_27540);
nor U28190 (N_28190,N_27091,N_27400);
and U28191 (N_28191,N_26705,N_26400);
nand U28192 (N_28192,N_27386,N_27399);
nand U28193 (N_28193,N_26662,N_26839);
nor U28194 (N_28194,N_26726,N_27492);
and U28195 (N_28195,N_26743,N_26631);
nand U28196 (N_28196,N_27322,N_26862);
nor U28197 (N_28197,N_27081,N_27292);
nor U28198 (N_28198,N_26960,N_27435);
xnor U28199 (N_28199,N_26483,N_27437);
xnor U28200 (N_28200,N_26611,N_26852);
nand U28201 (N_28201,N_26613,N_26655);
nor U28202 (N_28202,N_27364,N_26573);
nor U28203 (N_28203,N_27281,N_27473);
and U28204 (N_28204,N_26937,N_26954);
or U28205 (N_28205,N_27000,N_26407);
xnor U28206 (N_28206,N_26780,N_27381);
and U28207 (N_28207,N_26476,N_27270);
or U28208 (N_28208,N_26997,N_26733);
nor U28209 (N_28209,N_27563,N_26729);
xnor U28210 (N_28210,N_27110,N_26617);
and U28211 (N_28211,N_26779,N_27526);
or U28212 (N_28212,N_26505,N_26786);
nor U28213 (N_28213,N_26808,N_26924);
nor U28214 (N_28214,N_26578,N_27519);
nand U28215 (N_28215,N_27072,N_27158);
xnor U28216 (N_28216,N_26505,N_26506);
nand U28217 (N_28217,N_27598,N_27064);
or U28218 (N_28218,N_26607,N_27215);
nor U28219 (N_28219,N_27475,N_27083);
and U28220 (N_28220,N_26580,N_26980);
xor U28221 (N_28221,N_27198,N_27538);
xor U28222 (N_28222,N_27279,N_26540);
xnor U28223 (N_28223,N_26902,N_26768);
xnor U28224 (N_28224,N_27056,N_27364);
nor U28225 (N_28225,N_27245,N_26792);
or U28226 (N_28226,N_27310,N_27028);
and U28227 (N_28227,N_26950,N_26660);
nand U28228 (N_28228,N_27348,N_26477);
and U28229 (N_28229,N_26424,N_26762);
nor U28230 (N_28230,N_26671,N_26889);
nand U28231 (N_28231,N_27433,N_26908);
and U28232 (N_28232,N_27156,N_27567);
or U28233 (N_28233,N_27189,N_27173);
nor U28234 (N_28234,N_26465,N_27210);
or U28235 (N_28235,N_27569,N_26944);
nand U28236 (N_28236,N_26529,N_27130);
and U28237 (N_28237,N_27378,N_26929);
nor U28238 (N_28238,N_27161,N_26595);
and U28239 (N_28239,N_26542,N_27436);
nand U28240 (N_28240,N_26924,N_26918);
nor U28241 (N_28241,N_26511,N_26453);
nor U28242 (N_28242,N_27031,N_27007);
nand U28243 (N_28243,N_26925,N_27284);
or U28244 (N_28244,N_27463,N_27357);
xor U28245 (N_28245,N_26985,N_27183);
nand U28246 (N_28246,N_27283,N_27210);
xnor U28247 (N_28247,N_27296,N_27134);
and U28248 (N_28248,N_26489,N_27580);
xnor U28249 (N_28249,N_27174,N_26667);
and U28250 (N_28250,N_27055,N_27578);
xnor U28251 (N_28251,N_27502,N_26942);
and U28252 (N_28252,N_26873,N_26782);
or U28253 (N_28253,N_26832,N_26697);
or U28254 (N_28254,N_26472,N_26591);
nand U28255 (N_28255,N_26764,N_27087);
and U28256 (N_28256,N_26473,N_26998);
nor U28257 (N_28257,N_27188,N_26872);
and U28258 (N_28258,N_26636,N_26817);
nand U28259 (N_28259,N_26682,N_27377);
xnor U28260 (N_28260,N_26707,N_27288);
nor U28261 (N_28261,N_26557,N_26543);
nor U28262 (N_28262,N_27276,N_27494);
or U28263 (N_28263,N_26892,N_27579);
nand U28264 (N_28264,N_27552,N_26935);
xnor U28265 (N_28265,N_27031,N_27043);
and U28266 (N_28266,N_26764,N_26556);
nor U28267 (N_28267,N_27149,N_26900);
xnor U28268 (N_28268,N_26626,N_26513);
nor U28269 (N_28269,N_26937,N_27117);
xnor U28270 (N_28270,N_26764,N_26603);
and U28271 (N_28271,N_26614,N_26799);
and U28272 (N_28272,N_26956,N_26743);
or U28273 (N_28273,N_27010,N_27482);
or U28274 (N_28274,N_26814,N_26914);
and U28275 (N_28275,N_26668,N_27464);
or U28276 (N_28276,N_27296,N_26946);
or U28277 (N_28277,N_27019,N_27211);
xnor U28278 (N_28278,N_26526,N_26713);
xnor U28279 (N_28279,N_27095,N_26661);
nor U28280 (N_28280,N_26713,N_26668);
and U28281 (N_28281,N_26637,N_26650);
or U28282 (N_28282,N_27430,N_27220);
xnor U28283 (N_28283,N_26432,N_26846);
and U28284 (N_28284,N_26655,N_26846);
nand U28285 (N_28285,N_27292,N_26624);
xnor U28286 (N_28286,N_26781,N_26953);
or U28287 (N_28287,N_27306,N_26924);
nand U28288 (N_28288,N_27169,N_26814);
nand U28289 (N_28289,N_27386,N_27285);
and U28290 (N_28290,N_26889,N_26897);
nor U28291 (N_28291,N_26724,N_26989);
or U28292 (N_28292,N_27308,N_27222);
or U28293 (N_28293,N_27384,N_27573);
and U28294 (N_28294,N_27085,N_27223);
xnor U28295 (N_28295,N_26917,N_27329);
or U28296 (N_28296,N_27384,N_27245);
xor U28297 (N_28297,N_26814,N_27582);
nand U28298 (N_28298,N_27163,N_27485);
or U28299 (N_28299,N_26673,N_27345);
or U28300 (N_28300,N_26750,N_26902);
nor U28301 (N_28301,N_27107,N_27118);
or U28302 (N_28302,N_26482,N_27156);
and U28303 (N_28303,N_27017,N_27209);
nand U28304 (N_28304,N_27211,N_27430);
and U28305 (N_28305,N_27050,N_26600);
or U28306 (N_28306,N_26951,N_26979);
nor U28307 (N_28307,N_27291,N_27063);
or U28308 (N_28308,N_26980,N_27289);
nand U28309 (N_28309,N_26822,N_26840);
and U28310 (N_28310,N_26694,N_27117);
nor U28311 (N_28311,N_27260,N_26571);
xnor U28312 (N_28312,N_26688,N_26794);
nor U28313 (N_28313,N_27227,N_26906);
nand U28314 (N_28314,N_27147,N_27471);
nor U28315 (N_28315,N_26827,N_27533);
nor U28316 (N_28316,N_26869,N_27325);
and U28317 (N_28317,N_27267,N_27196);
nor U28318 (N_28318,N_27484,N_27273);
xnor U28319 (N_28319,N_27078,N_27046);
xor U28320 (N_28320,N_27443,N_27022);
nor U28321 (N_28321,N_26717,N_26482);
xnor U28322 (N_28322,N_27417,N_27014);
and U28323 (N_28323,N_27294,N_27571);
or U28324 (N_28324,N_27317,N_26824);
or U28325 (N_28325,N_27113,N_26836);
and U28326 (N_28326,N_26902,N_26799);
xnor U28327 (N_28327,N_26980,N_26513);
xor U28328 (N_28328,N_27504,N_27366);
xnor U28329 (N_28329,N_26953,N_27069);
or U28330 (N_28330,N_26744,N_27445);
nand U28331 (N_28331,N_27058,N_27373);
nand U28332 (N_28332,N_26715,N_27356);
or U28333 (N_28333,N_27161,N_27496);
or U28334 (N_28334,N_26637,N_27016);
or U28335 (N_28335,N_26785,N_26513);
or U28336 (N_28336,N_27128,N_27586);
nand U28337 (N_28337,N_27486,N_27007);
nor U28338 (N_28338,N_26728,N_27467);
nand U28339 (N_28339,N_27207,N_26836);
nand U28340 (N_28340,N_26892,N_27204);
xnor U28341 (N_28341,N_27357,N_26428);
xor U28342 (N_28342,N_27101,N_27456);
and U28343 (N_28343,N_26795,N_27331);
nand U28344 (N_28344,N_27546,N_27428);
xor U28345 (N_28345,N_27578,N_27407);
xnor U28346 (N_28346,N_26937,N_27043);
nor U28347 (N_28347,N_27551,N_26814);
or U28348 (N_28348,N_26520,N_27259);
nor U28349 (N_28349,N_27060,N_27263);
and U28350 (N_28350,N_27415,N_27326);
nand U28351 (N_28351,N_26540,N_26553);
nor U28352 (N_28352,N_26633,N_27484);
nor U28353 (N_28353,N_27216,N_26880);
nor U28354 (N_28354,N_27434,N_26426);
nand U28355 (N_28355,N_26584,N_26509);
or U28356 (N_28356,N_27418,N_26678);
and U28357 (N_28357,N_27342,N_26533);
nor U28358 (N_28358,N_26744,N_27090);
nor U28359 (N_28359,N_26612,N_26917);
or U28360 (N_28360,N_27135,N_26436);
xnor U28361 (N_28361,N_27524,N_26835);
or U28362 (N_28362,N_26848,N_26832);
and U28363 (N_28363,N_27132,N_27391);
nor U28364 (N_28364,N_27455,N_27444);
nor U28365 (N_28365,N_27020,N_26646);
and U28366 (N_28366,N_27290,N_27409);
xnor U28367 (N_28367,N_27001,N_26992);
nand U28368 (N_28368,N_26654,N_27148);
or U28369 (N_28369,N_27292,N_27384);
xor U28370 (N_28370,N_27414,N_26913);
or U28371 (N_28371,N_26876,N_26864);
or U28372 (N_28372,N_27303,N_27158);
or U28373 (N_28373,N_26662,N_26941);
xor U28374 (N_28374,N_27201,N_27252);
xnor U28375 (N_28375,N_27385,N_26976);
nor U28376 (N_28376,N_27081,N_27539);
xnor U28377 (N_28377,N_26635,N_27075);
xor U28378 (N_28378,N_27596,N_26660);
xnor U28379 (N_28379,N_26410,N_26754);
xnor U28380 (N_28380,N_27222,N_26905);
nor U28381 (N_28381,N_27472,N_27061);
or U28382 (N_28382,N_27438,N_27217);
nand U28383 (N_28383,N_26767,N_27476);
nand U28384 (N_28384,N_26430,N_26590);
nand U28385 (N_28385,N_26945,N_26958);
or U28386 (N_28386,N_27582,N_26799);
xnor U28387 (N_28387,N_27572,N_27130);
and U28388 (N_28388,N_26422,N_27123);
nand U28389 (N_28389,N_26884,N_26916);
nor U28390 (N_28390,N_26555,N_26454);
xnor U28391 (N_28391,N_27518,N_27196);
and U28392 (N_28392,N_27353,N_27113);
and U28393 (N_28393,N_27038,N_26553);
nand U28394 (N_28394,N_26479,N_26511);
xor U28395 (N_28395,N_27063,N_26991);
nand U28396 (N_28396,N_26936,N_26566);
and U28397 (N_28397,N_26474,N_27597);
nor U28398 (N_28398,N_26479,N_26534);
xnor U28399 (N_28399,N_26986,N_27292);
and U28400 (N_28400,N_27052,N_27050);
xnor U28401 (N_28401,N_27273,N_26943);
or U28402 (N_28402,N_27215,N_27499);
xor U28403 (N_28403,N_27285,N_26807);
or U28404 (N_28404,N_26980,N_26474);
or U28405 (N_28405,N_26727,N_26585);
nand U28406 (N_28406,N_27132,N_26670);
or U28407 (N_28407,N_27375,N_27453);
or U28408 (N_28408,N_26731,N_26561);
nand U28409 (N_28409,N_26686,N_26535);
nor U28410 (N_28410,N_26416,N_27380);
nand U28411 (N_28411,N_26844,N_26679);
or U28412 (N_28412,N_26745,N_26604);
or U28413 (N_28413,N_27404,N_26584);
nor U28414 (N_28414,N_26957,N_26895);
nor U28415 (N_28415,N_27077,N_26647);
or U28416 (N_28416,N_27175,N_27572);
nor U28417 (N_28417,N_27367,N_27454);
and U28418 (N_28418,N_26620,N_26788);
nand U28419 (N_28419,N_26826,N_27197);
nand U28420 (N_28420,N_26858,N_26479);
nand U28421 (N_28421,N_27091,N_27280);
nand U28422 (N_28422,N_26752,N_27407);
or U28423 (N_28423,N_27384,N_26506);
and U28424 (N_28424,N_27317,N_27061);
nor U28425 (N_28425,N_27149,N_26925);
nand U28426 (N_28426,N_27268,N_26411);
or U28427 (N_28427,N_26921,N_27495);
xor U28428 (N_28428,N_26956,N_27112);
xnor U28429 (N_28429,N_26876,N_26853);
or U28430 (N_28430,N_27301,N_26760);
or U28431 (N_28431,N_26425,N_26577);
nor U28432 (N_28432,N_27124,N_27531);
xor U28433 (N_28433,N_27511,N_27490);
xnor U28434 (N_28434,N_27160,N_26573);
nor U28435 (N_28435,N_26650,N_27425);
nand U28436 (N_28436,N_27112,N_27229);
xor U28437 (N_28437,N_27004,N_26833);
and U28438 (N_28438,N_27234,N_26982);
xor U28439 (N_28439,N_26665,N_27079);
nand U28440 (N_28440,N_26787,N_26747);
nand U28441 (N_28441,N_26784,N_26782);
or U28442 (N_28442,N_26751,N_26685);
xnor U28443 (N_28443,N_26545,N_26986);
or U28444 (N_28444,N_27465,N_27010);
or U28445 (N_28445,N_26720,N_27180);
nand U28446 (N_28446,N_26841,N_27018);
xor U28447 (N_28447,N_26471,N_26897);
xor U28448 (N_28448,N_26950,N_27060);
nand U28449 (N_28449,N_26800,N_26647);
or U28450 (N_28450,N_27306,N_27575);
and U28451 (N_28451,N_26672,N_27406);
and U28452 (N_28452,N_26805,N_27033);
nand U28453 (N_28453,N_27056,N_26457);
or U28454 (N_28454,N_26629,N_26974);
xor U28455 (N_28455,N_26862,N_26762);
nand U28456 (N_28456,N_26484,N_26936);
or U28457 (N_28457,N_26809,N_27220);
and U28458 (N_28458,N_26749,N_26528);
xor U28459 (N_28459,N_27145,N_26520);
nand U28460 (N_28460,N_26830,N_27232);
xnor U28461 (N_28461,N_26561,N_26780);
nand U28462 (N_28462,N_26593,N_27211);
and U28463 (N_28463,N_27061,N_26912);
nand U28464 (N_28464,N_27033,N_26430);
nor U28465 (N_28465,N_26989,N_26702);
nor U28466 (N_28466,N_27075,N_26907);
and U28467 (N_28467,N_26765,N_26734);
and U28468 (N_28468,N_27056,N_27265);
nand U28469 (N_28469,N_27492,N_26961);
or U28470 (N_28470,N_27163,N_26698);
nor U28471 (N_28471,N_26644,N_26968);
or U28472 (N_28472,N_26490,N_26877);
nor U28473 (N_28473,N_26541,N_26814);
xnor U28474 (N_28474,N_27498,N_27219);
nand U28475 (N_28475,N_27219,N_26641);
or U28476 (N_28476,N_27552,N_27148);
xnor U28477 (N_28477,N_27488,N_27493);
nor U28478 (N_28478,N_27587,N_26750);
nand U28479 (N_28479,N_26949,N_27092);
or U28480 (N_28480,N_27310,N_26560);
and U28481 (N_28481,N_27182,N_27449);
nor U28482 (N_28482,N_26947,N_26619);
and U28483 (N_28483,N_27498,N_26736);
xnor U28484 (N_28484,N_26832,N_27423);
or U28485 (N_28485,N_26762,N_26724);
nor U28486 (N_28486,N_27331,N_26487);
nand U28487 (N_28487,N_26708,N_26445);
and U28488 (N_28488,N_27102,N_26565);
xor U28489 (N_28489,N_26589,N_26577);
nor U28490 (N_28490,N_27218,N_27487);
xnor U28491 (N_28491,N_27385,N_26889);
and U28492 (N_28492,N_27246,N_27189);
and U28493 (N_28493,N_27556,N_27596);
nand U28494 (N_28494,N_27281,N_27046);
nand U28495 (N_28495,N_27100,N_27026);
or U28496 (N_28496,N_26556,N_26726);
and U28497 (N_28497,N_26949,N_27585);
nand U28498 (N_28498,N_26714,N_27191);
nor U28499 (N_28499,N_27187,N_26997);
xor U28500 (N_28500,N_26805,N_26943);
and U28501 (N_28501,N_27539,N_26511);
nor U28502 (N_28502,N_27092,N_27459);
or U28503 (N_28503,N_26909,N_27556);
or U28504 (N_28504,N_26925,N_26767);
xor U28505 (N_28505,N_27421,N_26973);
nor U28506 (N_28506,N_27453,N_26671);
or U28507 (N_28507,N_27594,N_26521);
and U28508 (N_28508,N_26596,N_26480);
or U28509 (N_28509,N_27437,N_26622);
xnor U28510 (N_28510,N_26924,N_26587);
and U28511 (N_28511,N_26612,N_27123);
and U28512 (N_28512,N_27353,N_26643);
and U28513 (N_28513,N_27456,N_26757);
or U28514 (N_28514,N_27462,N_26884);
nand U28515 (N_28515,N_27566,N_26705);
or U28516 (N_28516,N_26810,N_27477);
or U28517 (N_28517,N_26910,N_27101);
and U28518 (N_28518,N_26968,N_27412);
nor U28519 (N_28519,N_27463,N_26793);
or U28520 (N_28520,N_27428,N_27107);
nor U28521 (N_28521,N_27487,N_26774);
xnor U28522 (N_28522,N_27480,N_26639);
and U28523 (N_28523,N_26733,N_26889);
nor U28524 (N_28524,N_26701,N_26864);
and U28525 (N_28525,N_26808,N_26804);
xor U28526 (N_28526,N_26615,N_27085);
nand U28527 (N_28527,N_27002,N_26731);
or U28528 (N_28528,N_27167,N_27415);
nand U28529 (N_28529,N_27435,N_26912);
or U28530 (N_28530,N_26961,N_26677);
nand U28531 (N_28531,N_26667,N_27547);
and U28532 (N_28532,N_26959,N_26772);
or U28533 (N_28533,N_26972,N_27448);
or U28534 (N_28534,N_27485,N_27387);
or U28535 (N_28535,N_26622,N_26737);
nand U28536 (N_28536,N_27063,N_27393);
nor U28537 (N_28537,N_26490,N_26438);
xnor U28538 (N_28538,N_27418,N_26984);
nand U28539 (N_28539,N_27144,N_26446);
nor U28540 (N_28540,N_26426,N_26757);
or U28541 (N_28541,N_26906,N_27580);
nor U28542 (N_28542,N_26799,N_27066);
nand U28543 (N_28543,N_26956,N_26887);
or U28544 (N_28544,N_27007,N_27161);
xor U28545 (N_28545,N_27286,N_27547);
and U28546 (N_28546,N_27160,N_27266);
and U28547 (N_28547,N_27376,N_27252);
nand U28548 (N_28548,N_26608,N_26431);
nand U28549 (N_28549,N_26651,N_27213);
nand U28550 (N_28550,N_27407,N_26892);
nand U28551 (N_28551,N_27434,N_27140);
nand U28552 (N_28552,N_27031,N_27510);
nand U28553 (N_28553,N_27369,N_26535);
or U28554 (N_28554,N_26627,N_27119);
nand U28555 (N_28555,N_26681,N_27553);
nor U28556 (N_28556,N_27199,N_26907);
xnor U28557 (N_28557,N_26558,N_27234);
xnor U28558 (N_28558,N_27178,N_27510);
xor U28559 (N_28559,N_27041,N_26854);
nor U28560 (N_28560,N_26801,N_26941);
xnor U28561 (N_28561,N_26655,N_26651);
xnor U28562 (N_28562,N_26733,N_26608);
nand U28563 (N_28563,N_26789,N_27189);
xor U28564 (N_28564,N_26803,N_26666);
and U28565 (N_28565,N_27158,N_27491);
xor U28566 (N_28566,N_26781,N_26809);
and U28567 (N_28567,N_27377,N_26636);
nand U28568 (N_28568,N_27276,N_27527);
and U28569 (N_28569,N_26709,N_27521);
or U28570 (N_28570,N_26652,N_27578);
and U28571 (N_28571,N_26881,N_26409);
nor U28572 (N_28572,N_26570,N_27535);
xnor U28573 (N_28573,N_26969,N_27335);
nor U28574 (N_28574,N_27059,N_27555);
xor U28575 (N_28575,N_27359,N_27107);
nand U28576 (N_28576,N_27214,N_26813);
or U28577 (N_28577,N_27468,N_27023);
xor U28578 (N_28578,N_27020,N_27142);
or U28579 (N_28579,N_26866,N_27402);
and U28580 (N_28580,N_26649,N_27236);
or U28581 (N_28581,N_27249,N_26437);
and U28582 (N_28582,N_27311,N_27188);
xor U28583 (N_28583,N_27451,N_27324);
or U28584 (N_28584,N_27550,N_26861);
xnor U28585 (N_28585,N_27323,N_26472);
nor U28586 (N_28586,N_27129,N_26835);
xor U28587 (N_28587,N_27560,N_26439);
or U28588 (N_28588,N_27074,N_26565);
nor U28589 (N_28589,N_27506,N_27157);
and U28590 (N_28590,N_26801,N_27423);
or U28591 (N_28591,N_27432,N_27394);
or U28592 (N_28592,N_27590,N_26506);
xor U28593 (N_28593,N_27361,N_27294);
or U28594 (N_28594,N_26945,N_26853);
xnor U28595 (N_28595,N_27095,N_27394);
nor U28596 (N_28596,N_27075,N_26513);
nand U28597 (N_28597,N_26926,N_27533);
nand U28598 (N_28598,N_26766,N_27408);
or U28599 (N_28599,N_26429,N_27349);
nor U28600 (N_28600,N_27532,N_26701);
nand U28601 (N_28601,N_27442,N_26583);
xor U28602 (N_28602,N_27452,N_27515);
and U28603 (N_28603,N_27036,N_26422);
xor U28604 (N_28604,N_26508,N_26638);
and U28605 (N_28605,N_27398,N_26473);
and U28606 (N_28606,N_26692,N_27468);
nand U28607 (N_28607,N_27194,N_27480);
and U28608 (N_28608,N_26604,N_26773);
xnor U28609 (N_28609,N_27045,N_26875);
nand U28610 (N_28610,N_26731,N_26530);
nand U28611 (N_28611,N_27566,N_26558);
nand U28612 (N_28612,N_27179,N_27019);
nor U28613 (N_28613,N_27282,N_27357);
nor U28614 (N_28614,N_27391,N_26549);
and U28615 (N_28615,N_26464,N_27198);
xor U28616 (N_28616,N_27002,N_26698);
or U28617 (N_28617,N_27326,N_26501);
or U28618 (N_28618,N_27318,N_27583);
or U28619 (N_28619,N_26415,N_27152);
nand U28620 (N_28620,N_27400,N_26733);
nand U28621 (N_28621,N_27278,N_27217);
nor U28622 (N_28622,N_27575,N_26948);
nor U28623 (N_28623,N_27486,N_27138);
nor U28624 (N_28624,N_26680,N_26594);
nor U28625 (N_28625,N_27302,N_26817);
xor U28626 (N_28626,N_27046,N_26487);
nor U28627 (N_28627,N_27322,N_27255);
xor U28628 (N_28628,N_27005,N_27360);
or U28629 (N_28629,N_27316,N_26710);
nand U28630 (N_28630,N_26449,N_27036);
and U28631 (N_28631,N_26641,N_27356);
or U28632 (N_28632,N_26858,N_27001);
nand U28633 (N_28633,N_27232,N_27060);
nand U28634 (N_28634,N_26899,N_27039);
nand U28635 (N_28635,N_27592,N_26443);
xnor U28636 (N_28636,N_26917,N_26875);
xor U28637 (N_28637,N_27299,N_27374);
nor U28638 (N_28638,N_27243,N_26977);
and U28639 (N_28639,N_27144,N_26457);
nand U28640 (N_28640,N_27189,N_27024);
nand U28641 (N_28641,N_27212,N_26777);
and U28642 (N_28642,N_27318,N_27307);
xor U28643 (N_28643,N_26707,N_26940);
and U28644 (N_28644,N_27355,N_27085);
nor U28645 (N_28645,N_27004,N_26589);
and U28646 (N_28646,N_26707,N_26837);
xor U28647 (N_28647,N_27541,N_27339);
nor U28648 (N_28648,N_27361,N_26489);
xnor U28649 (N_28649,N_26706,N_27489);
xnor U28650 (N_28650,N_27306,N_27492);
nand U28651 (N_28651,N_27269,N_27125);
nor U28652 (N_28652,N_26840,N_26582);
or U28653 (N_28653,N_27365,N_26513);
xor U28654 (N_28654,N_26784,N_26409);
xor U28655 (N_28655,N_27030,N_27401);
nand U28656 (N_28656,N_26663,N_27534);
nor U28657 (N_28657,N_26662,N_27452);
nand U28658 (N_28658,N_26926,N_27551);
nand U28659 (N_28659,N_26549,N_27547);
or U28660 (N_28660,N_27523,N_26738);
nor U28661 (N_28661,N_27060,N_26663);
or U28662 (N_28662,N_27272,N_26486);
or U28663 (N_28663,N_26769,N_27080);
and U28664 (N_28664,N_26470,N_27288);
nor U28665 (N_28665,N_26519,N_26627);
nand U28666 (N_28666,N_26747,N_26448);
xnor U28667 (N_28667,N_26670,N_26533);
xor U28668 (N_28668,N_26964,N_27092);
or U28669 (N_28669,N_26725,N_26806);
xnor U28670 (N_28670,N_27093,N_26785);
or U28671 (N_28671,N_27064,N_27236);
xor U28672 (N_28672,N_27446,N_27032);
xnor U28673 (N_28673,N_27354,N_27280);
xor U28674 (N_28674,N_26493,N_26868);
and U28675 (N_28675,N_27244,N_26848);
xnor U28676 (N_28676,N_27269,N_27112);
xor U28677 (N_28677,N_26829,N_27129);
xnor U28678 (N_28678,N_26905,N_27308);
xnor U28679 (N_28679,N_26723,N_26511);
or U28680 (N_28680,N_27598,N_26945);
or U28681 (N_28681,N_26411,N_27239);
or U28682 (N_28682,N_26681,N_27403);
or U28683 (N_28683,N_26894,N_26581);
nand U28684 (N_28684,N_27452,N_26897);
xor U28685 (N_28685,N_26622,N_27107);
xnor U28686 (N_28686,N_26413,N_27183);
nor U28687 (N_28687,N_26903,N_26740);
nor U28688 (N_28688,N_26998,N_26820);
or U28689 (N_28689,N_26712,N_26748);
nand U28690 (N_28690,N_27389,N_27357);
xor U28691 (N_28691,N_26932,N_27489);
or U28692 (N_28692,N_26833,N_27150);
and U28693 (N_28693,N_26561,N_27402);
or U28694 (N_28694,N_27482,N_26415);
nand U28695 (N_28695,N_26728,N_26674);
xor U28696 (N_28696,N_27280,N_26471);
xnor U28697 (N_28697,N_26423,N_27513);
xor U28698 (N_28698,N_27437,N_26786);
nand U28699 (N_28699,N_27475,N_27205);
or U28700 (N_28700,N_27008,N_27589);
nand U28701 (N_28701,N_26573,N_26669);
nand U28702 (N_28702,N_26806,N_27420);
nor U28703 (N_28703,N_27392,N_26572);
nor U28704 (N_28704,N_27498,N_26461);
or U28705 (N_28705,N_26670,N_27512);
or U28706 (N_28706,N_26701,N_27044);
nor U28707 (N_28707,N_26852,N_27548);
nand U28708 (N_28708,N_27560,N_27582);
nor U28709 (N_28709,N_26839,N_26850);
nand U28710 (N_28710,N_27002,N_27219);
and U28711 (N_28711,N_27296,N_27409);
or U28712 (N_28712,N_27153,N_27328);
nand U28713 (N_28713,N_27212,N_26669);
nor U28714 (N_28714,N_26400,N_27317);
nand U28715 (N_28715,N_26478,N_27162);
nor U28716 (N_28716,N_27047,N_27398);
nand U28717 (N_28717,N_27537,N_27094);
or U28718 (N_28718,N_27078,N_26798);
or U28719 (N_28719,N_27504,N_26923);
nor U28720 (N_28720,N_27281,N_27170);
nor U28721 (N_28721,N_27483,N_27479);
nand U28722 (N_28722,N_26409,N_27297);
nand U28723 (N_28723,N_27109,N_26875);
nor U28724 (N_28724,N_26654,N_26586);
nor U28725 (N_28725,N_26405,N_26491);
or U28726 (N_28726,N_26422,N_26893);
xor U28727 (N_28727,N_26642,N_26765);
or U28728 (N_28728,N_27577,N_27412);
and U28729 (N_28729,N_26621,N_26506);
xor U28730 (N_28730,N_26855,N_26799);
or U28731 (N_28731,N_27445,N_27064);
nor U28732 (N_28732,N_27404,N_26567);
and U28733 (N_28733,N_27261,N_26856);
xnor U28734 (N_28734,N_26435,N_26784);
nand U28735 (N_28735,N_26729,N_27292);
xor U28736 (N_28736,N_27518,N_26586);
nand U28737 (N_28737,N_27556,N_26989);
xor U28738 (N_28738,N_27216,N_27414);
xor U28739 (N_28739,N_26641,N_27155);
nand U28740 (N_28740,N_27452,N_27366);
xnor U28741 (N_28741,N_26672,N_26861);
xnor U28742 (N_28742,N_27577,N_26972);
nor U28743 (N_28743,N_27121,N_26920);
nand U28744 (N_28744,N_26435,N_26497);
xor U28745 (N_28745,N_27564,N_27204);
nand U28746 (N_28746,N_27480,N_26847);
or U28747 (N_28747,N_27516,N_26808);
nand U28748 (N_28748,N_26492,N_27343);
and U28749 (N_28749,N_27161,N_26567);
nor U28750 (N_28750,N_26913,N_27511);
nand U28751 (N_28751,N_26965,N_27075);
xnor U28752 (N_28752,N_26525,N_27380);
or U28753 (N_28753,N_27315,N_27266);
or U28754 (N_28754,N_27114,N_27425);
xnor U28755 (N_28755,N_27274,N_27255);
xor U28756 (N_28756,N_26928,N_26580);
or U28757 (N_28757,N_27419,N_26400);
nand U28758 (N_28758,N_26555,N_26537);
nand U28759 (N_28759,N_27307,N_27469);
and U28760 (N_28760,N_27580,N_27207);
nand U28761 (N_28761,N_27089,N_26769);
and U28762 (N_28762,N_26791,N_27458);
nor U28763 (N_28763,N_27598,N_27599);
nand U28764 (N_28764,N_26607,N_26615);
nor U28765 (N_28765,N_27557,N_27384);
nand U28766 (N_28766,N_26975,N_26713);
and U28767 (N_28767,N_27472,N_27097);
nand U28768 (N_28768,N_26466,N_27224);
nor U28769 (N_28769,N_27563,N_27582);
xor U28770 (N_28770,N_26436,N_26529);
nor U28771 (N_28771,N_26575,N_27554);
xnor U28772 (N_28772,N_27575,N_27330);
xor U28773 (N_28773,N_27218,N_27488);
or U28774 (N_28774,N_26408,N_27523);
xor U28775 (N_28775,N_27057,N_26891);
nor U28776 (N_28776,N_26973,N_26464);
and U28777 (N_28777,N_27447,N_26728);
nor U28778 (N_28778,N_27016,N_26756);
nor U28779 (N_28779,N_27581,N_26463);
and U28780 (N_28780,N_26774,N_26873);
or U28781 (N_28781,N_27230,N_27069);
and U28782 (N_28782,N_26540,N_27562);
and U28783 (N_28783,N_26823,N_27074);
and U28784 (N_28784,N_27372,N_26973);
xnor U28785 (N_28785,N_26935,N_27289);
nor U28786 (N_28786,N_27410,N_26603);
or U28787 (N_28787,N_27268,N_26501);
nor U28788 (N_28788,N_26698,N_26550);
nand U28789 (N_28789,N_26640,N_27274);
and U28790 (N_28790,N_26624,N_27255);
and U28791 (N_28791,N_26742,N_26991);
nand U28792 (N_28792,N_26970,N_27564);
xor U28793 (N_28793,N_27034,N_27472);
and U28794 (N_28794,N_27169,N_27128);
nor U28795 (N_28795,N_27261,N_27517);
nor U28796 (N_28796,N_26691,N_26994);
and U28797 (N_28797,N_26811,N_26701);
nor U28798 (N_28798,N_26816,N_27287);
xnor U28799 (N_28799,N_27165,N_26978);
nand U28800 (N_28800,N_27888,N_27701);
xnor U28801 (N_28801,N_27666,N_27804);
nor U28802 (N_28802,N_28057,N_28086);
or U28803 (N_28803,N_28421,N_28129);
xnor U28804 (N_28804,N_28009,N_28371);
nand U28805 (N_28805,N_28203,N_27866);
and U28806 (N_28806,N_28730,N_28352);
nand U28807 (N_28807,N_27688,N_28109);
xor U28808 (N_28808,N_27803,N_27747);
xnor U28809 (N_28809,N_28073,N_28466);
xnor U28810 (N_28810,N_27644,N_28735);
xnor U28811 (N_28811,N_27626,N_28170);
nor U28812 (N_28812,N_28494,N_28445);
nand U28813 (N_28813,N_28161,N_28070);
nand U28814 (N_28814,N_28159,N_27630);
or U28815 (N_28815,N_28052,N_28343);
and U28816 (N_28816,N_28484,N_27749);
nor U28817 (N_28817,N_28426,N_28797);
nand U28818 (N_28818,N_27730,N_28675);
and U28819 (N_28819,N_28523,N_27836);
nor U28820 (N_28820,N_28672,N_28464);
nor U28821 (N_28821,N_28493,N_27713);
nor U28822 (N_28822,N_27825,N_28166);
nand U28823 (N_28823,N_27754,N_28011);
and U28824 (N_28824,N_27760,N_28568);
or U28825 (N_28825,N_27895,N_28134);
or U28826 (N_28826,N_28754,N_28604);
or U28827 (N_28827,N_28409,N_28624);
nor U28828 (N_28828,N_27673,N_27812);
nand U28829 (N_28829,N_27896,N_28255);
xor U28830 (N_28830,N_27704,N_27627);
nand U28831 (N_28831,N_28220,N_27671);
xor U28832 (N_28832,N_28405,N_28686);
xor U28833 (N_28833,N_27853,N_27699);
nor U28834 (N_28834,N_28776,N_28289);
nor U28835 (N_28835,N_27654,N_28571);
xnor U28836 (N_28836,N_27988,N_28152);
xnor U28837 (N_28837,N_28689,N_27722);
nand U28838 (N_28838,N_27905,N_28185);
and U28839 (N_28839,N_28591,N_27632);
nand U28840 (N_28840,N_28279,N_28027);
nand U28841 (N_28841,N_27822,N_27649);
or U28842 (N_28842,N_28507,N_27882);
xor U28843 (N_28843,N_28490,N_28463);
and U28844 (N_28844,N_28432,N_28475);
xor U28845 (N_28845,N_28457,N_27807);
and U28846 (N_28846,N_28277,N_28098);
or U28847 (N_28847,N_28721,N_28003);
xor U28848 (N_28848,N_27603,N_28626);
xnor U28849 (N_28849,N_27952,N_28211);
and U28850 (N_28850,N_27916,N_28154);
or U28851 (N_28851,N_28381,N_28276);
or U28852 (N_28852,N_28422,N_28094);
xor U28853 (N_28853,N_27799,N_28008);
or U28854 (N_28854,N_28573,N_27879);
xnor U28855 (N_28855,N_28254,N_28734);
nand U28856 (N_28856,N_27867,N_27748);
and U28857 (N_28857,N_28376,N_27857);
xnor U28858 (N_28858,N_27631,N_28497);
or U28859 (N_28859,N_28048,N_27765);
or U28860 (N_28860,N_28291,N_27979);
or U28861 (N_28861,N_28508,N_28299);
nand U28862 (N_28862,N_28112,N_27848);
and U28863 (N_28863,N_28582,N_27623);
xor U28864 (N_28864,N_28664,N_28329);
nor U28865 (N_28865,N_28026,N_28054);
and U28866 (N_28866,N_28130,N_28419);
nor U28867 (N_28867,N_28654,N_27665);
xnor U28868 (N_28868,N_27772,N_28715);
xnor U28869 (N_28869,N_27908,N_27615);
nand U28870 (N_28870,N_28013,N_27851);
or U28871 (N_28871,N_28058,N_27625);
nand U28872 (N_28872,N_28212,N_28088);
and U28873 (N_28873,N_28526,N_28439);
xnor U28874 (N_28874,N_28586,N_28521);
or U28875 (N_28875,N_28554,N_28183);
and U28876 (N_28876,N_28580,N_28035);
and U28877 (N_28877,N_28320,N_28744);
nand U28878 (N_28878,N_28075,N_28190);
xor U28879 (N_28879,N_28613,N_28179);
nor U28880 (N_28880,N_27697,N_27775);
nand U28881 (N_28881,N_27948,N_28794);
xnor U28882 (N_28882,N_28780,N_27845);
and U28883 (N_28883,N_27787,N_28551);
and U28884 (N_28884,N_28017,N_27993);
nand U28885 (N_28885,N_28180,N_27852);
or U28886 (N_28886,N_28694,N_28657);
nor U28887 (N_28887,N_27633,N_27849);
nand U28888 (N_28888,N_28216,N_27801);
xor U28889 (N_28889,N_27725,N_27756);
and U28890 (N_28890,N_28340,N_28728);
nand U28891 (N_28891,N_28652,N_28135);
or U28892 (N_28892,N_27683,N_28296);
nor U28893 (N_28893,N_28393,N_28782);
nand U28894 (N_28894,N_28483,N_28798);
nor U28895 (N_28895,N_27741,N_27838);
or U28896 (N_28896,N_28512,N_27911);
and U28897 (N_28897,N_28372,N_28007);
nand U28898 (N_28898,N_28060,N_27808);
nor U28899 (N_28899,N_27998,N_28459);
nor U28900 (N_28900,N_27921,N_28128);
nand U28901 (N_28901,N_28690,N_28682);
xnor U28902 (N_28902,N_28369,N_28022);
nand U28903 (N_28903,N_27717,N_27913);
xnor U28904 (N_28904,N_27823,N_27659);
nor U28905 (N_28905,N_28337,N_27777);
and U28906 (N_28906,N_28326,N_28449);
xor U28907 (N_28907,N_28074,N_27681);
and U28908 (N_28908,N_27837,N_27862);
nor U28909 (N_28909,N_28676,N_28127);
xor U28910 (N_28910,N_28383,N_27707);
xnor U28911 (N_28911,N_27985,N_28097);
nand U28912 (N_28912,N_28325,N_28479);
xor U28913 (N_28913,N_27859,N_28033);
or U28914 (N_28914,N_28763,N_28228);
nor U28915 (N_28915,N_27685,N_28710);
xor U28916 (N_28916,N_28537,N_28498);
xor U28917 (N_28917,N_27664,N_28010);
nor U28918 (N_28918,N_27931,N_27710);
nand U28919 (N_28919,N_28015,N_28647);
or U28920 (N_28920,N_28261,N_28217);
xnor U28921 (N_28921,N_28759,N_28608);
nor U28922 (N_28922,N_28633,N_28745);
nand U28923 (N_28923,N_28727,N_27968);
or U28924 (N_28924,N_27915,N_28062);
nand U28925 (N_28925,N_28614,N_27613);
and U28926 (N_28926,N_27820,N_27767);
and U28927 (N_28927,N_28142,N_27910);
xnor U28928 (N_28928,N_28565,N_28758);
or U28929 (N_28929,N_27796,N_27675);
or U28930 (N_28930,N_28321,N_28746);
nand U28931 (N_28931,N_28666,N_28595);
or U28932 (N_28932,N_28558,N_28160);
xnor U28933 (N_28933,N_28594,N_28413);
or U28934 (N_28934,N_28144,N_28367);
or U28935 (N_28935,N_27978,N_27800);
or U28936 (N_28936,N_27668,N_28462);
xnor U28937 (N_28937,N_27780,N_28082);
xor U28938 (N_28938,N_28430,N_28306);
nor U28939 (N_28939,N_27651,N_28729);
or U28940 (N_28940,N_28342,N_28638);
and U28941 (N_28941,N_27956,N_27745);
and U28942 (N_28942,N_28197,N_27719);
xnor U28943 (N_28943,N_28333,N_28678);
or U28944 (N_28944,N_27621,N_28083);
xnor U28945 (N_28945,N_27989,N_27709);
xnor U28946 (N_28946,N_28205,N_27642);
and U28947 (N_28947,N_28717,N_28605);
xor U28948 (N_28948,N_28742,N_27677);
or U28949 (N_28949,N_27770,N_28401);
nor U28950 (N_28950,N_28307,N_28467);
xnor U28951 (N_28951,N_28025,N_27661);
and U28952 (N_28952,N_28168,N_27903);
or U28953 (N_28953,N_28716,N_28520);
or U28954 (N_28954,N_28460,N_28324);
nor U28955 (N_28955,N_27983,N_28303);
nor U28956 (N_28956,N_28576,N_27794);
and U28957 (N_28957,N_28762,N_28514);
nor U28958 (N_28958,N_27815,N_28601);
nor U28959 (N_28959,N_28194,N_27982);
nand U28960 (N_28960,N_27928,N_27637);
nor U28961 (N_28961,N_28380,N_28028);
xor U28962 (N_28962,N_28093,N_28757);
nor U28963 (N_28963,N_28042,N_28519);
and U28964 (N_28964,N_28091,N_28038);
and U28965 (N_28965,N_28724,N_28646);
xnor U28966 (N_28966,N_28562,N_28767);
and U28967 (N_28967,N_28714,N_27698);
or U28968 (N_28968,N_28505,N_28612);
nor U28969 (N_28969,N_27616,N_27977);
nand U28970 (N_28970,N_28072,N_27892);
and U28971 (N_28971,N_28691,N_28698);
xor U28972 (N_28972,N_28719,N_28793);
or U28973 (N_28973,N_28773,N_28100);
nor U28974 (N_28974,N_28408,N_27889);
and U28975 (N_28975,N_28037,N_27758);
nor U28976 (N_28976,N_27899,N_28799);
or U28977 (N_28977,N_28471,N_28748);
nand U28978 (N_28978,N_28178,N_28473);
xnor U28979 (N_28979,N_28294,N_28014);
nor U28980 (N_28980,N_28566,N_28428);
xnor U28981 (N_28981,N_28658,N_27640);
nor U28982 (N_28982,N_27609,N_28029);
nor U28983 (N_28983,N_28359,N_28377);
and U28984 (N_28984,N_27716,N_28363);
and U28985 (N_28985,N_28740,N_27755);
and U28986 (N_28986,N_27648,N_28344);
or U28987 (N_28987,N_28561,N_27764);
xor U28988 (N_28988,N_28287,N_27774);
nand U28989 (N_28989,N_28396,N_27861);
xnor U28990 (N_28990,N_28442,N_28378);
or U28991 (N_28991,N_27940,N_27680);
or U28992 (N_28992,N_28310,N_28309);
and U28993 (N_28993,N_28567,N_27843);
or U28994 (N_28994,N_28739,N_28531);
or U28995 (N_28995,N_28140,N_28628);
or U28996 (N_28996,N_28547,N_28090);
nor U28997 (N_28997,N_27810,N_28575);
xnor U28998 (N_28998,N_28084,N_27802);
xor U28999 (N_28999,N_28769,N_27779);
or U29000 (N_29000,N_28214,N_28618);
nand U29001 (N_29001,N_28360,N_28248);
nor U29002 (N_29002,N_28670,N_28796);
or U29003 (N_29003,N_28468,N_28511);
xor U29004 (N_29004,N_27976,N_27693);
and U29005 (N_29005,N_27833,N_28684);
xnor U29006 (N_29006,N_28671,N_28357);
or U29007 (N_29007,N_28592,N_28712);
or U29008 (N_29008,N_27742,N_28024);
nor U29009 (N_29009,N_28673,N_28236);
xnor U29010 (N_29010,N_28019,N_28263);
nor U29011 (N_29011,N_28641,N_28315);
or U29012 (N_29012,N_28107,N_28031);
and U29013 (N_29013,N_28313,N_28574);
xor U29014 (N_29014,N_28208,N_28437);
xnor U29015 (N_29015,N_28785,N_28195);
or U29016 (N_29016,N_27686,N_28662);
and U29017 (N_29017,N_28262,N_28223);
nor U29018 (N_29018,N_28176,N_27721);
or U29019 (N_29019,N_28385,N_28499);
nand U29020 (N_29020,N_28219,N_28124);
and U29021 (N_29021,N_28650,N_28151);
or U29022 (N_29022,N_28132,N_28645);
xor U29023 (N_29023,N_28242,N_27737);
or U29024 (N_29024,N_28659,N_27938);
nand U29025 (N_29025,N_27925,N_28527);
nor U29026 (N_29026,N_27739,N_28032);
nand U29027 (N_29027,N_28111,N_27986);
and U29028 (N_29028,N_28105,N_28136);
or U29029 (N_29029,N_28260,N_27768);
nor U29030 (N_29030,N_28761,N_28751);
and U29031 (N_29031,N_27718,N_28541);
and U29032 (N_29032,N_28373,N_28725);
nor U29033 (N_29033,N_28472,N_27955);
and U29034 (N_29034,N_27622,N_28162);
or U29035 (N_29035,N_28210,N_28713);
or U29036 (N_29036,N_28397,N_28200);
nor U29037 (N_29037,N_28187,N_28529);
nand U29038 (N_29038,N_28685,N_28012);
or U29039 (N_29039,N_27792,N_28192);
xor U29040 (N_29040,N_28516,N_27893);
or U29041 (N_29041,N_28607,N_28317);
or U29042 (N_29042,N_28587,N_28298);
or U29043 (N_29043,N_28102,N_28427);
and U29044 (N_29044,N_27856,N_28726);
nand U29045 (N_29045,N_27670,N_28593);
nor U29046 (N_29046,N_28723,N_28133);
nor U29047 (N_29047,N_28224,N_28598);
nor U29048 (N_29048,N_28655,N_28441);
or U29049 (N_29049,N_27782,N_28648);
nor U29050 (N_29050,N_27620,N_27994);
or U29051 (N_29051,N_27639,N_27964);
xnor U29052 (N_29052,N_27924,N_27824);
or U29053 (N_29053,N_27904,N_28186);
xnor U29054 (N_29054,N_28538,N_28201);
and U29055 (N_29055,N_27865,N_28403);
nor U29056 (N_29056,N_28335,N_28006);
xor U29057 (N_29057,N_28524,N_28181);
and U29058 (N_29058,N_27814,N_28143);
and U29059 (N_29059,N_27846,N_27734);
nand U29060 (N_29060,N_28450,N_27869);
or U29061 (N_29061,N_28669,N_27963);
nor U29062 (N_29062,N_28485,N_28579);
nor U29063 (N_29063,N_28199,N_28354);
or U29064 (N_29064,N_28622,N_28774);
nor U29065 (N_29065,N_27771,N_28384);
nor U29066 (N_29066,N_28584,N_27682);
or U29067 (N_29067,N_28051,N_28544);
nand U29068 (N_29068,N_28632,N_28665);
nor U29069 (N_29069,N_28044,N_28046);
nor U29070 (N_29070,N_27635,N_28771);
or U29071 (N_29071,N_28522,N_27847);
nand U29072 (N_29072,N_28274,N_28681);
xor U29073 (N_29073,N_28602,N_28517);
nand U29074 (N_29074,N_27929,N_28731);
xor U29075 (N_29075,N_28451,N_27607);
and U29076 (N_29076,N_27645,N_28288);
nor U29077 (N_29077,N_28280,N_28709);
or U29078 (N_29078,N_28634,N_28259);
and U29079 (N_29079,N_28066,N_28000);
and U29080 (N_29080,N_27798,N_28703);
and U29081 (N_29081,N_27970,N_28290);
nand U29082 (N_29082,N_28600,N_28569);
or U29083 (N_29083,N_28271,N_28415);
xnor U29084 (N_29084,N_28314,N_28753);
or U29085 (N_29085,N_28533,N_28068);
and U29086 (N_29086,N_28244,N_27608);
xor U29087 (N_29087,N_28174,N_28452);
nand U29088 (N_29088,N_28610,N_28470);
nor U29089 (N_29089,N_28241,N_28080);
or U29090 (N_29090,N_28777,N_27981);
xnor U29091 (N_29091,N_28282,N_28707);
and U29092 (N_29092,N_27954,N_27712);
nor U29093 (N_29093,N_28747,N_28268);
nor U29094 (N_29094,N_27898,N_28117);
and U29095 (N_29095,N_27711,N_27695);
nor U29096 (N_29096,N_27936,N_28620);
and U29097 (N_29097,N_28394,N_28131);
and U29098 (N_29098,N_28433,N_28589);
and U29099 (N_29099,N_28518,N_27902);
nand U29100 (N_29100,N_28175,N_28379);
nand U29101 (N_29101,N_28424,N_28229);
or U29102 (N_29102,N_28559,N_28150);
nand U29103 (N_29103,N_28071,N_27678);
or U29104 (N_29104,N_28251,N_27870);
and U29105 (N_29105,N_28596,N_28041);
nand U29106 (N_29106,N_27927,N_28043);
or U29107 (N_29107,N_28103,N_28693);
nand U29108 (N_29108,N_27646,N_28458);
xor U29109 (N_29109,N_27900,N_27650);
nor U29110 (N_29110,N_28504,N_28704);
nand U29111 (N_29111,N_28273,N_28546);
nand U29112 (N_29112,N_27858,N_27990);
and U29113 (N_29113,N_27696,N_28651);
nor U29114 (N_29114,N_28264,N_28119);
or U29115 (N_29115,N_27844,N_28674);
or U29116 (N_29116,N_28115,N_27669);
xor U29117 (N_29117,N_28267,N_28435);
nor U29118 (N_29118,N_28619,N_28050);
or U29119 (N_29119,N_28350,N_27992);
nand U29120 (N_29120,N_27941,N_28525);
nor U29121 (N_29121,N_27880,N_27726);
xnor U29122 (N_29122,N_27660,N_28145);
xnor U29123 (N_29123,N_27687,N_28049);
nand U29124 (N_29124,N_28079,N_28249);
xnor U29125 (N_29125,N_28487,N_28482);
xor U29126 (N_29126,N_28137,N_28304);
and U29127 (N_29127,N_28030,N_28169);
xnor U29128 (N_29128,N_27818,N_27995);
nand U29129 (N_29129,N_28156,N_28440);
nand U29130 (N_29130,N_27934,N_28722);
nand U29131 (N_29131,N_27881,N_27652);
nand U29132 (N_29132,N_28346,N_28322);
nor U29133 (N_29133,N_27932,N_28697);
and U29134 (N_29134,N_27636,N_27984);
and U29135 (N_29135,N_28741,N_28540);
and U29136 (N_29136,N_28153,N_28486);
xor U29137 (N_29137,N_27723,N_28149);
nand U29138 (N_29138,N_28636,N_28085);
and U29139 (N_29139,N_28055,N_28680);
xor U29140 (N_29140,N_28238,N_27887);
nor U29141 (N_29141,N_28171,N_27624);
or U29142 (N_29142,N_28338,N_27731);
and U29143 (N_29143,N_27789,N_28496);
nand U29144 (N_29144,N_28345,N_27876);
xor U29145 (N_29145,N_28417,N_28077);
xor U29146 (N_29146,N_28474,N_27914);
xor U29147 (N_29147,N_28283,N_28364);
nand U29148 (N_29148,N_27735,N_28502);
xnor U29149 (N_29149,N_27702,N_28772);
or U29150 (N_29150,N_28549,N_28184);
nand U29151 (N_29151,N_28163,N_28755);
or U29152 (N_29152,N_28786,N_27841);
nand U29153 (N_29153,N_27816,N_28300);
nor U29154 (N_29154,N_28640,N_28114);
nand U29155 (N_29155,N_28695,N_28791);
and U29156 (N_29156,N_27871,N_28534);
or U29157 (N_29157,N_28063,N_28067);
nor U29158 (N_29158,N_28756,N_28705);
xor U29159 (N_29159,N_27872,N_27805);
nor U29160 (N_29160,N_28588,N_28234);
or U29161 (N_29161,N_27602,N_28056);
nand U29162 (N_29162,N_27811,N_28362);
or U29163 (N_29163,N_27834,N_28766);
or U29164 (N_29164,N_28765,N_28256);
xnor U29165 (N_29165,N_27829,N_28316);
nor U29166 (N_29166,N_28778,N_28366);
and U29167 (N_29167,N_27855,N_28631);
nor U29168 (N_29168,N_28456,N_28410);
xor U29169 (N_29169,N_27894,N_27667);
or U29170 (N_29170,N_28095,N_28461);
xnor U29171 (N_29171,N_28232,N_28311);
and U29172 (N_29172,N_28454,N_28065);
or U29173 (N_29173,N_27918,N_27647);
xor U29174 (N_29174,N_27766,N_28198);
and U29175 (N_29175,N_28609,N_28661);
and U29176 (N_29176,N_28683,N_28545);
or U29177 (N_29177,N_28089,N_28370);
xnor U29178 (N_29178,N_28209,N_27923);
and U29179 (N_29179,N_28790,N_28349);
or U29180 (N_29180,N_28500,N_28110);
nand U29181 (N_29181,N_28692,N_28227);
and U29182 (N_29182,N_27877,N_28365);
or U29183 (N_29183,N_28503,N_27891);
or U29184 (N_29184,N_28222,N_28202);
or U29185 (N_29185,N_27835,N_27655);
nor U29186 (N_29186,N_28611,N_27935);
nand U29187 (N_29187,N_28557,N_28061);
xor U29188 (N_29188,N_27944,N_28361);
nand U29189 (N_29189,N_27676,N_28539);
nand U29190 (N_29190,N_28585,N_28688);
nor U29191 (N_29191,N_28578,N_27689);
and U29192 (N_29192,N_28447,N_28718);
nand U29193 (N_29193,N_27732,N_28278);
xor U29194 (N_29194,N_27953,N_27875);
xor U29195 (N_29195,N_27634,N_28020);
and U29196 (N_29196,N_28436,N_28699);
nor U29197 (N_29197,N_28218,N_27863);
nand U29198 (N_29198,N_27919,N_28243);
nor U29199 (N_29199,N_28528,N_28226);
and U29200 (N_29200,N_28284,N_28590);
xor U29201 (N_29201,N_27897,N_28334);
nor U29202 (N_29202,N_28481,N_27657);
and U29203 (N_29203,N_28318,N_28301);
xor U29204 (N_29204,N_28501,N_27819);
xor U29205 (N_29205,N_28572,N_28305);
and U29206 (N_29206,N_27662,N_27753);
nor U29207 (N_29207,N_27720,N_27797);
and U29208 (N_29208,N_28630,N_28649);
nor U29209 (N_29209,N_28126,N_28548);
xor U29210 (N_29210,N_27750,N_28101);
nor U29211 (N_29211,N_27945,N_28275);
nand U29212 (N_29212,N_28489,N_28270);
nand U29213 (N_29213,N_28016,N_27864);
nor U29214 (N_29214,N_28668,N_28550);
nor U29215 (N_29215,N_28792,N_28687);
or U29216 (N_29216,N_27757,N_28087);
nand U29217 (N_29217,N_27920,N_28347);
xnor U29218 (N_29218,N_27949,N_28491);
or U29219 (N_29219,N_28239,N_28002);
and U29220 (N_29220,N_27878,N_28444);
or U29221 (N_29221,N_28297,N_27672);
xnor U29222 (N_29222,N_28420,N_28642);
nand U29223 (N_29223,N_28116,N_28789);
nand U29224 (N_29224,N_28700,N_28005);
or U29225 (N_29225,N_28480,N_28250);
nand U29226 (N_29226,N_28542,N_27705);
or U29227 (N_29227,N_28230,N_28059);
nand U29228 (N_29228,N_28099,N_28108);
xnor U29229 (N_29229,N_28768,N_27656);
nor U29230 (N_29230,N_27950,N_28553);
nor U29231 (N_29231,N_28375,N_28615);
and U29232 (N_29232,N_28412,N_28237);
or U29233 (N_29233,N_27684,N_28775);
nand U29234 (N_29234,N_28076,N_27874);
nor U29235 (N_29235,N_28193,N_28532);
and U29236 (N_29236,N_28530,N_27761);
xnor U29237 (N_29237,N_28233,N_27809);
and U29238 (N_29238,N_28509,N_28231);
nor U29239 (N_29239,N_27738,N_28737);
or U29240 (N_29240,N_28123,N_27769);
xnor U29241 (N_29241,N_27980,N_28269);
and U29242 (N_29242,N_27641,N_27907);
nor U29243 (N_29243,N_27612,N_27744);
and U29244 (N_29244,N_27600,N_27972);
nand U29245 (N_29245,N_27778,N_27885);
or U29246 (N_29246,N_27961,N_28312);
nor U29247 (N_29247,N_27715,N_28147);
and U29248 (N_29248,N_28382,N_28783);
and U29249 (N_29249,N_28328,N_27691);
nor U29250 (N_29250,N_28355,N_27965);
or U29251 (N_29251,N_28660,N_28599);
and U29252 (N_29252,N_28696,N_28779);
nor U29253 (N_29253,N_28506,N_28749);
nand U29254 (N_29254,N_28390,N_27793);
and U29255 (N_29255,N_27604,N_28711);
or U29256 (N_29256,N_28387,N_27724);
nor U29257 (N_29257,N_28146,N_28395);
nor U29258 (N_29258,N_28515,N_28570);
nand U29259 (N_29259,N_28281,N_28351);
nor U29260 (N_29260,N_28398,N_28787);
xor U29261 (N_29261,N_28701,N_27912);
nor U29262 (N_29262,N_27839,N_27997);
xnor U29263 (N_29263,N_28760,N_28606);
and U29264 (N_29264,N_28583,N_28252);
or U29265 (N_29265,N_27746,N_27813);
xor U29266 (N_29266,N_27773,N_28556);
or U29267 (N_29267,N_28167,N_28603);
xor U29268 (N_29268,N_27806,N_27901);
and U29269 (N_29269,N_28577,N_27628);
and U29270 (N_29270,N_27930,N_27991);
and U29271 (N_29271,N_27643,N_28004);
and U29272 (N_29272,N_28510,N_27614);
nand U29273 (N_29273,N_27832,N_27751);
xnor U29274 (N_29274,N_28627,N_28411);
or U29275 (N_29275,N_28391,N_27939);
or U29276 (N_29276,N_27909,N_28327);
xnor U29277 (N_29277,N_28443,N_27943);
nor U29278 (N_29278,N_27840,N_28406);
or U29279 (N_29279,N_28448,N_28720);
nor U29280 (N_29280,N_27617,N_28122);
nor U29281 (N_29281,N_27960,N_27854);
nand U29282 (N_29282,N_28253,N_27618);
and U29283 (N_29283,N_27690,N_28356);
or U29284 (N_29284,N_28469,N_28285);
or U29285 (N_29285,N_27860,N_27850);
and U29286 (N_29286,N_27728,N_28348);
nand U29287 (N_29287,N_28045,N_28096);
nor U29288 (N_29288,N_28106,N_28563);
xnor U29289 (N_29289,N_28138,N_28743);
and U29290 (N_29290,N_28555,N_28784);
or U29291 (N_29291,N_28207,N_27922);
and U29292 (N_29292,N_27974,N_27601);
xor U29293 (N_29293,N_27763,N_28018);
xnor U29294 (N_29294,N_28247,N_27759);
or U29295 (N_29295,N_28139,N_27679);
or U29296 (N_29296,N_27830,N_27951);
xnor U29297 (N_29297,N_27842,N_28302);
and U29298 (N_29298,N_27937,N_27933);
nor U29299 (N_29299,N_27886,N_27791);
xor U29300 (N_29300,N_28308,N_28182);
and U29301 (N_29301,N_28643,N_27714);
nand U29302 (N_29302,N_28323,N_28039);
or U29303 (N_29303,N_28332,N_28629);
or U29304 (N_29304,N_28639,N_28221);
and U29305 (N_29305,N_28092,N_28266);
nor U29306 (N_29306,N_27692,N_27653);
or U29307 (N_29307,N_28165,N_28191);
and U29308 (N_29308,N_27828,N_27827);
xnor U29309 (N_29309,N_27966,N_28155);
xor U29310 (N_29310,N_28141,N_28418);
nand U29311 (N_29311,N_27817,N_28478);
nor U29312 (N_29312,N_28189,N_28021);
nor U29313 (N_29313,N_28120,N_27826);
nand U29314 (N_29314,N_28495,N_28621);
xor U29315 (N_29315,N_28431,N_28225);
nor U29316 (N_29316,N_28286,N_28679);
nand U29317 (N_29317,N_28173,N_28113);
xor U29318 (N_29318,N_27999,N_28069);
or U29319 (N_29319,N_28341,N_27781);
nand U29320 (N_29320,N_28036,N_28616);
nor U29321 (N_29321,N_27629,N_28121);
nor U29322 (N_29322,N_28023,N_28295);
or U29323 (N_29323,N_27873,N_27606);
xor U29324 (N_29324,N_28386,N_27785);
or U29325 (N_29325,N_28564,N_28764);
nand U29326 (N_29326,N_28177,N_28118);
or U29327 (N_29327,N_27740,N_28752);
nand U29328 (N_29328,N_28402,N_28438);
xor U29329 (N_29329,N_28240,N_27946);
nand U29330 (N_29330,N_28374,N_27906);
nand U29331 (N_29331,N_28477,N_28272);
or U29332 (N_29332,N_28001,N_28733);
nor U29333 (N_29333,N_27821,N_27795);
nor U29334 (N_29334,N_28081,N_28235);
nand U29335 (N_29335,N_28206,N_28635);
xor U29336 (N_29336,N_27638,N_28158);
nor U29337 (N_29337,N_28513,N_27962);
nand U29338 (N_29338,N_28788,N_27708);
nor U29339 (N_29339,N_28246,N_27790);
or U29340 (N_29340,N_28732,N_28623);
nand U29341 (N_29341,N_27700,N_27729);
and U29342 (N_29342,N_28414,N_27776);
nand U29343 (N_29343,N_28407,N_27663);
nor U29344 (N_29344,N_27727,N_28617);
xor U29345 (N_29345,N_28404,N_28392);
nor U29346 (N_29346,N_28319,N_28637);
xor U29347 (N_29347,N_27959,N_27975);
nor U29348 (N_29348,N_28172,N_28388);
nand U29349 (N_29349,N_28560,N_28148);
and U29350 (N_29350,N_28750,N_28795);
and U29351 (N_29351,N_27605,N_28677);
nand U29352 (N_29352,N_28781,N_28258);
and U29353 (N_29353,N_28353,N_27958);
xor U29354 (N_29354,N_27967,N_28265);
nor U29355 (N_29355,N_27694,N_28157);
and U29356 (N_29356,N_28164,N_28389);
nor U29357 (N_29357,N_28453,N_28213);
xnor U29358 (N_29358,N_28104,N_28429);
and U29359 (N_29359,N_28245,N_27736);
and U29360 (N_29360,N_27619,N_28416);
nor U29361 (N_29361,N_27947,N_27917);
and U29362 (N_29362,N_28488,N_27752);
and U29363 (N_29363,N_27969,N_28663);
xnor U29364 (N_29364,N_27762,N_28625);
nor U29365 (N_29365,N_27957,N_28331);
or U29366 (N_29366,N_27788,N_28257);
nand U29367 (N_29367,N_27884,N_28425);
nand U29368 (N_29368,N_28204,N_28597);
or U29369 (N_29369,N_28455,N_27783);
or U29370 (N_29370,N_27610,N_28644);
or U29371 (N_29371,N_28339,N_28656);
or U29372 (N_29372,N_27987,N_28125);
or U29373 (N_29373,N_27706,N_28581);
nand U29374 (N_29374,N_27611,N_28465);
and U29375 (N_29375,N_27942,N_28667);
nand U29376 (N_29376,N_28330,N_27674);
nor U29377 (N_29377,N_27868,N_27883);
nand U29378 (N_29378,N_28293,N_28736);
xor U29379 (N_29379,N_27733,N_28196);
nand U29380 (N_29380,N_27658,N_28400);
nand U29381 (N_29381,N_28492,N_28653);
nand U29382 (N_29382,N_28706,N_27971);
or U29383 (N_29383,N_28078,N_27703);
and U29384 (N_29384,N_27784,N_28399);
and U29385 (N_29385,N_28423,N_28738);
xnor U29386 (N_29386,N_28476,N_28708);
and U29387 (N_29387,N_28040,N_27743);
and U29388 (N_29388,N_28034,N_27786);
xor U29389 (N_29389,N_28215,N_28536);
nand U29390 (N_29390,N_28047,N_27890);
xor U29391 (N_29391,N_28535,N_28368);
and U29392 (N_29392,N_28358,N_28543);
xor U29393 (N_29393,N_28292,N_27973);
nor U29394 (N_29394,N_28770,N_28188);
or U29395 (N_29395,N_28336,N_27831);
or U29396 (N_29396,N_28053,N_27926);
and U29397 (N_29397,N_28064,N_28434);
nand U29398 (N_29398,N_28702,N_28446);
and U29399 (N_29399,N_27996,N_28552);
nor U29400 (N_29400,N_27772,N_28487);
or U29401 (N_29401,N_28145,N_28480);
xnor U29402 (N_29402,N_28501,N_28293);
xor U29403 (N_29403,N_27975,N_28691);
nand U29404 (N_29404,N_28526,N_28423);
nor U29405 (N_29405,N_27876,N_28014);
or U29406 (N_29406,N_28431,N_27665);
or U29407 (N_29407,N_27600,N_27938);
nor U29408 (N_29408,N_28316,N_28693);
nand U29409 (N_29409,N_28034,N_28363);
xor U29410 (N_29410,N_27643,N_27998);
or U29411 (N_29411,N_27639,N_28422);
xnor U29412 (N_29412,N_28385,N_28213);
and U29413 (N_29413,N_28304,N_27907);
nand U29414 (N_29414,N_28456,N_28097);
and U29415 (N_29415,N_28347,N_27953);
nor U29416 (N_29416,N_28478,N_28756);
xor U29417 (N_29417,N_28010,N_28667);
or U29418 (N_29418,N_27615,N_28521);
xnor U29419 (N_29419,N_28779,N_27958);
xor U29420 (N_29420,N_28324,N_27934);
and U29421 (N_29421,N_27987,N_27947);
nand U29422 (N_29422,N_28329,N_28253);
nand U29423 (N_29423,N_28079,N_28758);
and U29424 (N_29424,N_28313,N_27689);
or U29425 (N_29425,N_27822,N_27923);
nand U29426 (N_29426,N_27619,N_28694);
nor U29427 (N_29427,N_28198,N_28605);
nand U29428 (N_29428,N_28560,N_27789);
nor U29429 (N_29429,N_28279,N_27809);
xnor U29430 (N_29430,N_28654,N_27879);
nand U29431 (N_29431,N_28073,N_28009);
and U29432 (N_29432,N_27978,N_28788);
or U29433 (N_29433,N_27745,N_27801);
nand U29434 (N_29434,N_27994,N_28175);
or U29435 (N_29435,N_28248,N_28039);
nor U29436 (N_29436,N_27804,N_27967);
or U29437 (N_29437,N_28605,N_28209);
and U29438 (N_29438,N_27884,N_28236);
xnor U29439 (N_29439,N_28789,N_28738);
and U29440 (N_29440,N_27762,N_28279);
or U29441 (N_29441,N_28038,N_27767);
xnor U29442 (N_29442,N_28036,N_27764);
nand U29443 (N_29443,N_28143,N_28704);
nand U29444 (N_29444,N_28092,N_27744);
nand U29445 (N_29445,N_27769,N_28107);
and U29446 (N_29446,N_28342,N_28598);
and U29447 (N_29447,N_28561,N_27941);
nor U29448 (N_29448,N_28507,N_28760);
and U29449 (N_29449,N_27959,N_28186);
and U29450 (N_29450,N_28787,N_28115);
xor U29451 (N_29451,N_28504,N_27981);
nand U29452 (N_29452,N_28609,N_27888);
and U29453 (N_29453,N_28516,N_28689);
and U29454 (N_29454,N_28774,N_28129);
and U29455 (N_29455,N_28082,N_27968);
and U29456 (N_29456,N_28761,N_28506);
xnor U29457 (N_29457,N_28484,N_27752);
nor U29458 (N_29458,N_28294,N_28631);
and U29459 (N_29459,N_28228,N_27912);
nand U29460 (N_29460,N_27943,N_28065);
and U29461 (N_29461,N_28208,N_27992);
nor U29462 (N_29462,N_27702,N_28105);
xnor U29463 (N_29463,N_28604,N_27671);
nand U29464 (N_29464,N_27898,N_28571);
nor U29465 (N_29465,N_28370,N_28389);
nor U29466 (N_29466,N_28299,N_28345);
nand U29467 (N_29467,N_27653,N_28735);
nor U29468 (N_29468,N_28793,N_27886);
or U29469 (N_29469,N_28274,N_28499);
or U29470 (N_29470,N_27874,N_28350);
or U29471 (N_29471,N_27983,N_28609);
nand U29472 (N_29472,N_28466,N_27697);
nand U29473 (N_29473,N_28417,N_27978);
or U29474 (N_29474,N_28187,N_27821);
xor U29475 (N_29475,N_28239,N_28033);
xnor U29476 (N_29476,N_28525,N_28406);
and U29477 (N_29477,N_28488,N_27941);
nor U29478 (N_29478,N_27983,N_27760);
xnor U29479 (N_29479,N_27852,N_28284);
and U29480 (N_29480,N_27672,N_28436);
nand U29481 (N_29481,N_27818,N_27654);
or U29482 (N_29482,N_27871,N_28594);
nor U29483 (N_29483,N_28120,N_28203);
nor U29484 (N_29484,N_28443,N_27703);
and U29485 (N_29485,N_28146,N_27601);
xor U29486 (N_29486,N_28000,N_28257);
xor U29487 (N_29487,N_28061,N_28676);
nor U29488 (N_29488,N_27747,N_28160);
nand U29489 (N_29489,N_28717,N_28160);
nor U29490 (N_29490,N_27897,N_28724);
nor U29491 (N_29491,N_28303,N_28415);
or U29492 (N_29492,N_28776,N_28190);
nor U29493 (N_29493,N_27781,N_28750);
nor U29494 (N_29494,N_28445,N_27691);
and U29495 (N_29495,N_28548,N_28328);
xnor U29496 (N_29496,N_28019,N_27819);
or U29497 (N_29497,N_28638,N_27922);
nand U29498 (N_29498,N_28069,N_27656);
or U29499 (N_29499,N_28514,N_27702);
nor U29500 (N_29500,N_27814,N_28768);
nor U29501 (N_29501,N_28350,N_28428);
xor U29502 (N_29502,N_28384,N_28489);
or U29503 (N_29503,N_27651,N_28376);
or U29504 (N_29504,N_27848,N_27605);
or U29505 (N_29505,N_28402,N_27742);
and U29506 (N_29506,N_28473,N_27886);
nor U29507 (N_29507,N_28730,N_28478);
or U29508 (N_29508,N_27762,N_27983);
nand U29509 (N_29509,N_28135,N_28022);
xnor U29510 (N_29510,N_27629,N_28018);
xor U29511 (N_29511,N_28515,N_28343);
and U29512 (N_29512,N_27625,N_28617);
nand U29513 (N_29513,N_27651,N_28377);
or U29514 (N_29514,N_27887,N_27789);
xor U29515 (N_29515,N_27935,N_28169);
and U29516 (N_29516,N_28347,N_28417);
nor U29517 (N_29517,N_28089,N_27959);
nor U29518 (N_29518,N_28175,N_28531);
and U29519 (N_29519,N_27872,N_28322);
nand U29520 (N_29520,N_28626,N_28385);
and U29521 (N_29521,N_28573,N_28373);
nand U29522 (N_29522,N_27747,N_28761);
xor U29523 (N_29523,N_28391,N_27670);
nor U29524 (N_29524,N_28058,N_28272);
or U29525 (N_29525,N_27954,N_27706);
nor U29526 (N_29526,N_27663,N_28193);
and U29527 (N_29527,N_27909,N_27972);
nor U29528 (N_29528,N_27751,N_27760);
xor U29529 (N_29529,N_27721,N_28643);
nor U29530 (N_29530,N_27865,N_27898);
nor U29531 (N_29531,N_28437,N_28300);
or U29532 (N_29532,N_28110,N_27770);
nand U29533 (N_29533,N_28323,N_28003);
nor U29534 (N_29534,N_28267,N_28015);
nor U29535 (N_29535,N_28066,N_27760);
and U29536 (N_29536,N_28395,N_28645);
or U29537 (N_29537,N_28450,N_27863);
xnor U29538 (N_29538,N_27881,N_27765);
xor U29539 (N_29539,N_28292,N_28416);
nand U29540 (N_29540,N_27910,N_27627);
or U29541 (N_29541,N_27930,N_27979);
xor U29542 (N_29542,N_27659,N_28427);
xnor U29543 (N_29543,N_28138,N_27676);
nand U29544 (N_29544,N_28599,N_28010);
nor U29545 (N_29545,N_27967,N_27842);
or U29546 (N_29546,N_27885,N_28521);
nand U29547 (N_29547,N_27897,N_28356);
xor U29548 (N_29548,N_27791,N_28415);
or U29549 (N_29549,N_28143,N_28165);
nand U29550 (N_29550,N_28137,N_27664);
nand U29551 (N_29551,N_28299,N_27886);
xnor U29552 (N_29552,N_28421,N_28480);
nor U29553 (N_29553,N_28552,N_28705);
xnor U29554 (N_29554,N_28190,N_28605);
or U29555 (N_29555,N_28589,N_27858);
and U29556 (N_29556,N_28069,N_28583);
or U29557 (N_29557,N_28420,N_28153);
nor U29558 (N_29558,N_28779,N_28520);
nand U29559 (N_29559,N_28253,N_27960);
nor U29560 (N_29560,N_28783,N_28771);
nor U29561 (N_29561,N_28418,N_28381);
xor U29562 (N_29562,N_28280,N_28675);
and U29563 (N_29563,N_28725,N_27807);
or U29564 (N_29564,N_27801,N_28531);
and U29565 (N_29565,N_28399,N_28138);
or U29566 (N_29566,N_27969,N_27646);
and U29567 (N_29567,N_28667,N_27630);
xnor U29568 (N_29568,N_28266,N_28214);
and U29569 (N_29569,N_27714,N_28066);
and U29570 (N_29570,N_27849,N_28177);
nor U29571 (N_29571,N_27905,N_27722);
or U29572 (N_29572,N_27813,N_27613);
nand U29573 (N_29573,N_28491,N_27743);
or U29574 (N_29574,N_28680,N_28760);
or U29575 (N_29575,N_28766,N_28757);
and U29576 (N_29576,N_27654,N_28343);
nand U29577 (N_29577,N_27649,N_28627);
nand U29578 (N_29578,N_28660,N_28722);
xor U29579 (N_29579,N_28077,N_28323);
or U29580 (N_29580,N_28701,N_28280);
or U29581 (N_29581,N_28319,N_28516);
and U29582 (N_29582,N_28780,N_27939);
xnor U29583 (N_29583,N_28194,N_27669);
nor U29584 (N_29584,N_28089,N_28585);
or U29585 (N_29585,N_28549,N_28775);
xor U29586 (N_29586,N_28282,N_28186);
nor U29587 (N_29587,N_28782,N_27650);
nand U29588 (N_29588,N_27609,N_28572);
nand U29589 (N_29589,N_28135,N_28387);
and U29590 (N_29590,N_27925,N_28431);
and U29591 (N_29591,N_28711,N_27820);
nand U29592 (N_29592,N_28595,N_27758);
and U29593 (N_29593,N_28743,N_27773);
and U29594 (N_29594,N_27718,N_28160);
and U29595 (N_29595,N_27942,N_27844);
xor U29596 (N_29596,N_28028,N_28341);
nor U29597 (N_29597,N_28251,N_28137);
and U29598 (N_29598,N_28757,N_27931);
and U29599 (N_29599,N_27819,N_28262);
nand U29600 (N_29600,N_28474,N_28746);
xnor U29601 (N_29601,N_28511,N_28024);
nor U29602 (N_29602,N_27651,N_28692);
nor U29603 (N_29603,N_27610,N_28475);
or U29604 (N_29604,N_28529,N_27726);
nor U29605 (N_29605,N_27889,N_28573);
nand U29606 (N_29606,N_27982,N_28603);
xnor U29607 (N_29607,N_28508,N_27715);
nor U29608 (N_29608,N_27768,N_27711);
nor U29609 (N_29609,N_28595,N_28590);
xnor U29610 (N_29610,N_28630,N_28558);
or U29611 (N_29611,N_28400,N_27947);
nor U29612 (N_29612,N_28502,N_28525);
nor U29613 (N_29613,N_28788,N_27757);
nor U29614 (N_29614,N_27705,N_28215);
nand U29615 (N_29615,N_27951,N_28650);
nand U29616 (N_29616,N_28357,N_28710);
xor U29617 (N_29617,N_28405,N_28787);
nor U29618 (N_29618,N_28768,N_27698);
nand U29619 (N_29619,N_28729,N_28423);
nor U29620 (N_29620,N_28192,N_28021);
nor U29621 (N_29621,N_28257,N_28579);
or U29622 (N_29622,N_27716,N_27738);
or U29623 (N_29623,N_27617,N_28650);
or U29624 (N_29624,N_28210,N_27686);
nand U29625 (N_29625,N_27883,N_28013);
xnor U29626 (N_29626,N_28775,N_28081);
nand U29627 (N_29627,N_28259,N_28443);
or U29628 (N_29628,N_28118,N_28209);
nor U29629 (N_29629,N_28582,N_27842);
nor U29630 (N_29630,N_28778,N_28349);
or U29631 (N_29631,N_28088,N_28462);
nor U29632 (N_29632,N_28235,N_27773);
and U29633 (N_29633,N_28764,N_28778);
xnor U29634 (N_29634,N_28423,N_28360);
xnor U29635 (N_29635,N_28740,N_28452);
xnor U29636 (N_29636,N_28102,N_28656);
nand U29637 (N_29637,N_28335,N_28549);
nor U29638 (N_29638,N_28215,N_28239);
nand U29639 (N_29639,N_28003,N_27756);
nand U29640 (N_29640,N_28497,N_27989);
or U29641 (N_29641,N_27784,N_28642);
and U29642 (N_29642,N_28007,N_28184);
or U29643 (N_29643,N_28179,N_28353);
xnor U29644 (N_29644,N_28628,N_27840);
nand U29645 (N_29645,N_27822,N_28631);
xnor U29646 (N_29646,N_27949,N_27830);
or U29647 (N_29647,N_28544,N_27854);
or U29648 (N_29648,N_28207,N_27945);
nor U29649 (N_29649,N_28512,N_28258);
nand U29650 (N_29650,N_27812,N_28339);
or U29651 (N_29651,N_28156,N_28395);
nand U29652 (N_29652,N_27690,N_28737);
xor U29653 (N_29653,N_27646,N_27835);
xnor U29654 (N_29654,N_28155,N_27642);
xor U29655 (N_29655,N_28286,N_28031);
or U29656 (N_29656,N_27797,N_28229);
nor U29657 (N_29657,N_27985,N_27627);
or U29658 (N_29658,N_28013,N_27710);
nand U29659 (N_29659,N_27725,N_27870);
and U29660 (N_29660,N_28234,N_28485);
or U29661 (N_29661,N_28232,N_28257);
xnor U29662 (N_29662,N_28689,N_27978);
and U29663 (N_29663,N_28624,N_28155);
and U29664 (N_29664,N_28566,N_28496);
nor U29665 (N_29665,N_28394,N_27814);
nand U29666 (N_29666,N_28198,N_28482);
xor U29667 (N_29667,N_28537,N_27823);
xnor U29668 (N_29668,N_27614,N_28063);
xor U29669 (N_29669,N_28693,N_27934);
and U29670 (N_29670,N_28040,N_28060);
nor U29671 (N_29671,N_28304,N_28766);
xor U29672 (N_29672,N_28301,N_28409);
and U29673 (N_29673,N_28590,N_28454);
and U29674 (N_29674,N_28123,N_27988);
xnor U29675 (N_29675,N_27997,N_27952);
nor U29676 (N_29676,N_27778,N_28361);
and U29677 (N_29677,N_28694,N_28380);
and U29678 (N_29678,N_28559,N_28222);
nand U29679 (N_29679,N_28128,N_27825);
and U29680 (N_29680,N_27890,N_27869);
and U29681 (N_29681,N_27809,N_27759);
and U29682 (N_29682,N_28085,N_28067);
xnor U29683 (N_29683,N_28506,N_28119);
nor U29684 (N_29684,N_27780,N_28129);
nand U29685 (N_29685,N_28414,N_28531);
xnor U29686 (N_29686,N_28028,N_28288);
and U29687 (N_29687,N_28461,N_28195);
nor U29688 (N_29688,N_28267,N_27990);
and U29689 (N_29689,N_27600,N_28575);
nor U29690 (N_29690,N_28154,N_28699);
and U29691 (N_29691,N_28214,N_28105);
or U29692 (N_29692,N_28042,N_27741);
nand U29693 (N_29693,N_28017,N_28087);
xnor U29694 (N_29694,N_28709,N_28680);
nor U29695 (N_29695,N_28300,N_28608);
nand U29696 (N_29696,N_28746,N_27883);
and U29697 (N_29697,N_27705,N_28778);
nor U29698 (N_29698,N_27933,N_27883);
xor U29699 (N_29699,N_28281,N_28225);
nor U29700 (N_29700,N_28093,N_28726);
nor U29701 (N_29701,N_27695,N_27796);
nor U29702 (N_29702,N_28364,N_28213);
and U29703 (N_29703,N_27622,N_28198);
nand U29704 (N_29704,N_28103,N_28247);
xnor U29705 (N_29705,N_27802,N_27775);
or U29706 (N_29706,N_28094,N_28486);
and U29707 (N_29707,N_28344,N_28786);
or U29708 (N_29708,N_28594,N_27957);
nand U29709 (N_29709,N_28626,N_28517);
or U29710 (N_29710,N_28177,N_27901);
nor U29711 (N_29711,N_28284,N_28373);
nor U29712 (N_29712,N_28671,N_28510);
nand U29713 (N_29713,N_28014,N_28234);
xnor U29714 (N_29714,N_28655,N_27799);
nand U29715 (N_29715,N_27923,N_28333);
or U29716 (N_29716,N_28218,N_28588);
or U29717 (N_29717,N_28764,N_27772);
xnor U29718 (N_29718,N_28453,N_27752);
xnor U29719 (N_29719,N_28142,N_27630);
and U29720 (N_29720,N_27709,N_28320);
xor U29721 (N_29721,N_28450,N_27794);
or U29722 (N_29722,N_27987,N_28695);
or U29723 (N_29723,N_27814,N_27843);
nor U29724 (N_29724,N_28799,N_27658);
nand U29725 (N_29725,N_27683,N_28124);
or U29726 (N_29726,N_28718,N_28698);
and U29727 (N_29727,N_28600,N_27703);
nor U29728 (N_29728,N_28030,N_28774);
or U29729 (N_29729,N_28341,N_28165);
nand U29730 (N_29730,N_28782,N_27728);
xor U29731 (N_29731,N_28479,N_28766);
nor U29732 (N_29732,N_27673,N_27622);
and U29733 (N_29733,N_28237,N_27827);
or U29734 (N_29734,N_27952,N_28022);
nand U29735 (N_29735,N_28697,N_27801);
or U29736 (N_29736,N_27800,N_28233);
nand U29737 (N_29737,N_28282,N_28031);
xnor U29738 (N_29738,N_28177,N_27769);
xnor U29739 (N_29739,N_28651,N_28758);
and U29740 (N_29740,N_28481,N_28236);
nor U29741 (N_29741,N_28717,N_28490);
nand U29742 (N_29742,N_28263,N_27689);
and U29743 (N_29743,N_28698,N_28676);
nor U29744 (N_29744,N_27721,N_28166);
or U29745 (N_29745,N_27614,N_27785);
and U29746 (N_29746,N_27660,N_27999);
nand U29747 (N_29747,N_27941,N_28222);
nor U29748 (N_29748,N_27853,N_27883);
nand U29749 (N_29749,N_27975,N_27928);
and U29750 (N_29750,N_28242,N_28041);
nor U29751 (N_29751,N_28369,N_27646);
nor U29752 (N_29752,N_27889,N_27910);
and U29753 (N_29753,N_27866,N_28672);
or U29754 (N_29754,N_28735,N_28321);
nor U29755 (N_29755,N_28246,N_27793);
and U29756 (N_29756,N_28311,N_27939);
xnor U29757 (N_29757,N_28346,N_28542);
or U29758 (N_29758,N_28401,N_28480);
nor U29759 (N_29759,N_27878,N_28239);
and U29760 (N_29760,N_28061,N_27941);
or U29761 (N_29761,N_27695,N_28795);
nand U29762 (N_29762,N_28128,N_27600);
xnor U29763 (N_29763,N_28131,N_28762);
and U29764 (N_29764,N_27771,N_28309);
and U29765 (N_29765,N_28443,N_27741);
nor U29766 (N_29766,N_28717,N_27793);
nand U29767 (N_29767,N_28563,N_27652);
nor U29768 (N_29768,N_28502,N_28201);
xnor U29769 (N_29769,N_28458,N_27999);
and U29770 (N_29770,N_28715,N_28316);
or U29771 (N_29771,N_27874,N_28735);
xnor U29772 (N_29772,N_27775,N_28624);
nand U29773 (N_29773,N_27644,N_28634);
and U29774 (N_29774,N_28721,N_28609);
and U29775 (N_29775,N_27917,N_28628);
nand U29776 (N_29776,N_28680,N_27696);
or U29777 (N_29777,N_27857,N_28778);
nand U29778 (N_29778,N_28104,N_28048);
xor U29779 (N_29779,N_27653,N_28385);
nor U29780 (N_29780,N_27983,N_28126);
nor U29781 (N_29781,N_27610,N_28088);
nand U29782 (N_29782,N_28772,N_28061);
xor U29783 (N_29783,N_27905,N_28469);
nand U29784 (N_29784,N_28471,N_28454);
and U29785 (N_29785,N_28126,N_28532);
or U29786 (N_29786,N_28549,N_28742);
nand U29787 (N_29787,N_27849,N_28701);
nor U29788 (N_29788,N_28775,N_28214);
and U29789 (N_29789,N_28430,N_28265);
nor U29790 (N_29790,N_28241,N_27966);
or U29791 (N_29791,N_27678,N_28722);
nand U29792 (N_29792,N_27627,N_28101);
or U29793 (N_29793,N_27728,N_28595);
and U29794 (N_29794,N_28014,N_27647);
and U29795 (N_29795,N_28066,N_27932);
xnor U29796 (N_29796,N_28444,N_28716);
xor U29797 (N_29797,N_28698,N_27810);
and U29798 (N_29798,N_27904,N_27630);
xnor U29799 (N_29799,N_28035,N_27960);
xor U29800 (N_29800,N_28438,N_28512);
or U29801 (N_29801,N_27976,N_28347);
or U29802 (N_29802,N_28798,N_28365);
or U29803 (N_29803,N_27912,N_28709);
nand U29804 (N_29804,N_27973,N_28589);
xor U29805 (N_29805,N_28362,N_28790);
xnor U29806 (N_29806,N_27732,N_28139);
xor U29807 (N_29807,N_27770,N_28220);
or U29808 (N_29808,N_27940,N_28644);
xnor U29809 (N_29809,N_28032,N_28509);
nor U29810 (N_29810,N_28086,N_27881);
nand U29811 (N_29811,N_28192,N_28580);
nand U29812 (N_29812,N_28156,N_27835);
xnor U29813 (N_29813,N_28088,N_28296);
xnor U29814 (N_29814,N_27994,N_28152);
nor U29815 (N_29815,N_28697,N_28682);
nand U29816 (N_29816,N_27879,N_28432);
or U29817 (N_29817,N_27992,N_27902);
or U29818 (N_29818,N_27949,N_27974);
nand U29819 (N_29819,N_27621,N_28402);
or U29820 (N_29820,N_28259,N_28193);
xnor U29821 (N_29821,N_28516,N_27669);
xnor U29822 (N_29822,N_28222,N_27733);
xnor U29823 (N_29823,N_28724,N_27846);
or U29824 (N_29824,N_28770,N_27901);
nor U29825 (N_29825,N_28153,N_28463);
nand U29826 (N_29826,N_27994,N_27787);
nand U29827 (N_29827,N_28218,N_27881);
nand U29828 (N_29828,N_28332,N_27679);
and U29829 (N_29829,N_28180,N_28447);
and U29830 (N_29830,N_28584,N_28018);
nand U29831 (N_29831,N_27601,N_28689);
nand U29832 (N_29832,N_28411,N_28525);
or U29833 (N_29833,N_28341,N_27847);
nand U29834 (N_29834,N_28747,N_27742);
or U29835 (N_29835,N_27767,N_28614);
or U29836 (N_29836,N_28097,N_28736);
and U29837 (N_29837,N_28522,N_27934);
or U29838 (N_29838,N_28513,N_28553);
xnor U29839 (N_29839,N_28598,N_27864);
or U29840 (N_29840,N_27797,N_28490);
or U29841 (N_29841,N_28276,N_28609);
xnor U29842 (N_29842,N_28507,N_27906);
and U29843 (N_29843,N_27937,N_28300);
and U29844 (N_29844,N_28781,N_28274);
nand U29845 (N_29845,N_28757,N_28261);
nand U29846 (N_29846,N_27699,N_28226);
xor U29847 (N_29847,N_28001,N_27900);
and U29848 (N_29848,N_28133,N_28684);
or U29849 (N_29849,N_27620,N_28060);
and U29850 (N_29850,N_28179,N_27803);
nor U29851 (N_29851,N_27747,N_28497);
or U29852 (N_29852,N_27902,N_28110);
nand U29853 (N_29853,N_28590,N_28113);
or U29854 (N_29854,N_28175,N_28618);
xnor U29855 (N_29855,N_28243,N_28799);
or U29856 (N_29856,N_27684,N_28527);
and U29857 (N_29857,N_27686,N_28546);
nand U29858 (N_29858,N_27721,N_28522);
xnor U29859 (N_29859,N_28438,N_27985);
nor U29860 (N_29860,N_28616,N_27744);
nand U29861 (N_29861,N_28372,N_28010);
nor U29862 (N_29862,N_28466,N_28453);
xnor U29863 (N_29863,N_28233,N_28014);
nor U29864 (N_29864,N_27677,N_27830);
nand U29865 (N_29865,N_28058,N_28087);
and U29866 (N_29866,N_27764,N_27951);
and U29867 (N_29867,N_28122,N_27755);
xor U29868 (N_29868,N_28746,N_28444);
nor U29869 (N_29869,N_27740,N_28378);
nor U29870 (N_29870,N_28550,N_28625);
or U29871 (N_29871,N_28774,N_28165);
xor U29872 (N_29872,N_27626,N_28031);
and U29873 (N_29873,N_28002,N_28253);
xor U29874 (N_29874,N_28712,N_27833);
and U29875 (N_29875,N_28092,N_28475);
xnor U29876 (N_29876,N_27790,N_28650);
xor U29877 (N_29877,N_28058,N_28780);
or U29878 (N_29878,N_28011,N_27603);
nor U29879 (N_29879,N_27906,N_27641);
or U29880 (N_29880,N_27804,N_28664);
xor U29881 (N_29881,N_27655,N_28313);
nand U29882 (N_29882,N_28476,N_27880);
nor U29883 (N_29883,N_27835,N_27959);
or U29884 (N_29884,N_28184,N_28381);
and U29885 (N_29885,N_27720,N_27660);
xor U29886 (N_29886,N_28191,N_28764);
nand U29887 (N_29887,N_28711,N_27840);
xor U29888 (N_29888,N_27679,N_28690);
nand U29889 (N_29889,N_28365,N_28563);
nand U29890 (N_29890,N_28530,N_27879);
nor U29891 (N_29891,N_28309,N_28396);
and U29892 (N_29892,N_27861,N_27982);
or U29893 (N_29893,N_28421,N_28712);
or U29894 (N_29894,N_27781,N_27972);
or U29895 (N_29895,N_28655,N_28432);
and U29896 (N_29896,N_28008,N_27825);
nand U29897 (N_29897,N_27625,N_27867);
nor U29898 (N_29898,N_28203,N_27782);
and U29899 (N_29899,N_28157,N_27848);
nand U29900 (N_29900,N_28559,N_28716);
and U29901 (N_29901,N_27894,N_28299);
xor U29902 (N_29902,N_27953,N_28113);
nor U29903 (N_29903,N_28327,N_27919);
or U29904 (N_29904,N_28423,N_28461);
nor U29905 (N_29905,N_28754,N_28495);
or U29906 (N_29906,N_27755,N_28601);
and U29907 (N_29907,N_27755,N_28737);
xor U29908 (N_29908,N_28623,N_28593);
nor U29909 (N_29909,N_28130,N_28461);
xor U29910 (N_29910,N_27613,N_28203);
and U29911 (N_29911,N_28320,N_28666);
and U29912 (N_29912,N_28265,N_28423);
or U29913 (N_29913,N_27996,N_27746);
nor U29914 (N_29914,N_27988,N_27605);
nand U29915 (N_29915,N_28621,N_28462);
nor U29916 (N_29916,N_28051,N_28308);
or U29917 (N_29917,N_27986,N_28243);
nand U29918 (N_29918,N_28780,N_27646);
and U29919 (N_29919,N_28030,N_28647);
xnor U29920 (N_29920,N_28380,N_28756);
or U29921 (N_29921,N_28633,N_27953);
nand U29922 (N_29922,N_28791,N_28002);
nor U29923 (N_29923,N_28362,N_28307);
xnor U29924 (N_29924,N_28193,N_28692);
or U29925 (N_29925,N_27702,N_27717);
or U29926 (N_29926,N_28066,N_27981);
xor U29927 (N_29927,N_28714,N_28789);
nor U29928 (N_29928,N_28274,N_28487);
or U29929 (N_29929,N_28592,N_27711);
nor U29930 (N_29930,N_28713,N_28268);
nor U29931 (N_29931,N_28506,N_28518);
nand U29932 (N_29932,N_27811,N_28287);
nand U29933 (N_29933,N_28588,N_27836);
or U29934 (N_29934,N_28767,N_27801);
and U29935 (N_29935,N_28246,N_27656);
xor U29936 (N_29936,N_28269,N_28538);
and U29937 (N_29937,N_28629,N_28530);
nand U29938 (N_29938,N_27676,N_27635);
or U29939 (N_29939,N_28333,N_28726);
nand U29940 (N_29940,N_27756,N_28206);
or U29941 (N_29941,N_28051,N_28636);
xnor U29942 (N_29942,N_28583,N_28175);
nand U29943 (N_29943,N_28204,N_27777);
and U29944 (N_29944,N_28194,N_28214);
nand U29945 (N_29945,N_27960,N_28146);
nor U29946 (N_29946,N_28087,N_28567);
or U29947 (N_29947,N_28546,N_28573);
nand U29948 (N_29948,N_28226,N_27651);
or U29949 (N_29949,N_27877,N_28073);
xnor U29950 (N_29950,N_27906,N_27934);
and U29951 (N_29951,N_27834,N_28726);
nand U29952 (N_29952,N_28577,N_28547);
or U29953 (N_29953,N_27733,N_27816);
nor U29954 (N_29954,N_28027,N_28449);
nand U29955 (N_29955,N_28470,N_28643);
or U29956 (N_29956,N_28636,N_28785);
xnor U29957 (N_29957,N_27709,N_27657);
or U29958 (N_29958,N_27747,N_28083);
or U29959 (N_29959,N_28753,N_28051);
nand U29960 (N_29960,N_27895,N_28708);
and U29961 (N_29961,N_28115,N_27689);
nand U29962 (N_29962,N_28026,N_28750);
and U29963 (N_29963,N_27729,N_27630);
or U29964 (N_29964,N_28697,N_28620);
xnor U29965 (N_29965,N_28060,N_27655);
nor U29966 (N_29966,N_28381,N_28685);
or U29967 (N_29967,N_28504,N_28545);
xor U29968 (N_29968,N_28001,N_28216);
xor U29969 (N_29969,N_27965,N_28733);
or U29970 (N_29970,N_28099,N_28310);
or U29971 (N_29971,N_28666,N_28600);
nand U29972 (N_29972,N_27848,N_28420);
or U29973 (N_29973,N_28255,N_28087);
or U29974 (N_29974,N_28553,N_27920);
and U29975 (N_29975,N_28036,N_28255);
nor U29976 (N_29976,N_28733,N_28375);
nand U29977 (N_29977,N_27831,N_27786);
nor U29978 (N_29978,N_28191,N_27632);
or U29979 (N_29979,N_28073,N_27649);
and U29980 (N_29980,N_28469,N_28157);
or U29981 (N_29981,N_28518,N_28100);
nand U29982 (N_29982,N_28128,N_27859);
nand U29983 (N_29983,N_28690,N_27835);
or U29984 (N_29984,N_28213,N_28045);
or U29985 (N_29985,N_28775,N_28278);
nand U29986 (N_29986,N_28194,N_28021);
nor U29987 (N_29987,N_28611,N_28250);
xnor U29988 (N_29988,N_28743,N_28263);
nor U29989 (N_29989,N_27636,N_27696);
xor U29990 (N_29990,N_28462,N_28687);
xor U29991 (N_29991,N_28534,N_28640);
xnor U29992 (N_29992,N_28450,N_27922);
or U29993 (N_29993,N_27978,N_28467);
nand U29994 (N_29994,N_28740,N_28250);
nor U29995 (N_29995,N_28451,N_27694);
nand U29996 (N_29996,N_27773,N_28158);
and U29997 (N_29997,N_28032,N_28353);
nor U29998 (N_29998,N_28407,N_27684);
nor U29999 (N_29999,N_28791,N_27727);
nand UO_0 (O_0,N_29581,N_29161);
nand UO_1 (O_1,N_28930,N_28896);
or UO_2 (O_2,N_29085,N_29696);
xnor UO_3 (O_3,N_29726,N_29140);
and UO_4 (O_4,N_29611,N_29612);
and UO_5 (O_5,N_29450,N_29947);
or UO_6 (O_6,N_29335,N_29151);
xnor UO_7 (O_7,N_29305,N_29339);
or UO_8 (O_8,N_28815,N_29863);
or UO_9 (O_9,N_29349,N_29606);
and UO_10 (O_10,N_29075,N_29482);
xor UO_11 (O_11,N_29650,N_29683);
and UO_12 (O_12,N_29087,N_29879);
and UO_13 (O_13,N_29752,N_29928);
and UO_14 (O_14,N_29435,N_29246);
nor UO_15 (O_15,N_28843,N_28857);
or UO_16 (O_16,N_29204,N_29854);
nand UO_17 (O_17,N_29320,N_28903);
or UO_18 (O_18,N_29155,N_29713);
nor UO_19 (O_19,N_29596,N_28914);
or UO_20 (O_20,N_28844,N_29266);
xnor UO_21 (O_21,N_29425,N_29795);
or UO_22 (O_22,N_29493,N_29990);
and UO_23 (O_23,N_29211,N_29836);
xnor UO_24 (O_24,N_29406,N_29171);
xnor UO_25 (O_25,N_29597,N_29167);
xnor UO_26 (O_26,N_29804,N_29277);
and UO_27 (O_27,N_29569,N_29258);
or UO_28 (O_28,N_29021,N_29945);
or UO_29 (O_29,N_29833,N_29391);
nand UO_30 (O_30,N_29269,N_29234);
nand UO_31 (O_31,N_28982,N_29851);
nor UO_32 (O_32,N_29102,N_28852);
and UO_33 (O_33,N_28824,N_29004);
and UO_34 (O_34,N_29438,N_29710);
nand UO_35 (O_35,N_29537,N_28855);
or UO_36 (O_36,N_29203,N_29826);
nor UO_37 (O_37,N_28970,N_29018);
nor UO_38 (O_38,N_28871,N_29379);
and UO_39 (O_39,N_29392,N_29940);
nand UO_40 (O_40,N_29638,N_29201);
xor UO_41 (O_41,N_29512,N_29012);
nand UO_42 (O_42,N_29785,N_29137);
or UO_43 (O_43,N_29646,N_29426);
or UO_44 (O_44,N_28868,N_28836);
xnor UO_45 (O_45,N_29427,N_29359);
or UO_46 (O_46,N_28864,N_29968);
or UO_47 (O_47,N_28999,N_28909);
nor UO_48 (O_48,N_29381,N_29421);
xnor UO_49 (O_49,N_29232,N_29236);
xnor UO_50 (O_50,N_29371,N_29434);
or UO_51 (O_51,N_29002,N_29995);
or UO_52 (O_52,N_28845,N_29964);
or UO_53 (O_53,N_29202,N_28819);
xnor UO_54 (O_54,N_29261,N_29496);
or UO_55 (O_55,N_29275,N_29858);
xnor UO_56 (O_56,N_29593,N_29505);
and UO_57 (O_57,N_29109,N_29896);
nor UO_58 (O_58,N_29924,N_29466);
nand UO_59 (O_59,N_29721,N_29189);
nor UO_60 (O_60,N_29300,N_29812);
nand UO_61 (O_61,N_29913,N_29692);
or UO_62 (O_62,N_29464,N_29460);
nand UO_63 (O_63,N_29264,N_29310);
and UO_64 (O_64,N_29338,N_29456);
and UO_65 (O_65,N_29552,N_29472);
xor UO_66 (O_66,N_28906,N_29626);
nor UO_67 (O_67,N_29322,N_29765);
or UO_68 (O_68,N_29191,N_29452);
and UO_69 (O_69,N_29374,N_29568);
nand UO_70 (O_70,N_29480,N_29759);
nand UO_71 (O_71,N_29748,N_29001);
and UO_72 (O_72,N_29554,N_29503);
nand UO_73 (O_73,N_29311,N_29429);
or UO_74 (O_74,N_29585,N_29390);
or UO_75 (O_75,N_28986,N_29690);
nor UO_76 (O_76,N_29788,N_29485);
xor UO_77 (O_77,N_29987,N_29797);
nand UO_78 (O_78,N_29048,N_29306);
or UO_79 (O_79,N_29570,N_29933);
xnor UO_80 (O_80,N_29294,N_28923);
and UO_81 (O_81,N_29011,N_28990);
or UO_82 (O_82,N_29756,N_29398);
nor UO_83 (O_83,N_29800,N_29601);
or UO_84 (O_84,N_29971,N_29342);
xnor UO_85 (O_85,N_29350,N_28885);
nor UO_86 (O_86,N_29817,N_29355);
nor UO_87 (O_87,N_29318,N_29367);
and UO_88 (O_88,N_28863,N_29509);
and UO_89 (O_89,N_29327,N_29571);
and UO_90 (O_90,N_29679,N_29681);
xor UO_91 (O_91,N_29985,N_28941);
nor UO_92 (O_92,N_29873,N_29285);
and UO_93 (O_93,N_28804,N_29813);
xnor UO_94 (O_94,N_29841,N_29044);
nand UO_95 (O_95,N_29187,N_29096);
xnor UO_96 (O_96,N_28908,N_28891);
xnor UO_97 (O_97,N_29963,N_29908);
nand UO_98 (O_98,N_29459,N_29885);
xnor UO_99 (O_99,N_29210,N_29418);
xnor UO_100 (O_100,N_29218,N_29592);
or UO_101 (O_101,N_28913,N_28883);
xor UO_102 (O_102,N_29378,N_29824);
nand UO_103 (O_103,N_29404,N_29637);
and UO_104 (O_104,N_29420,N_28818);
nand UO_105 (O_105,N_29206,N_29220);
xor UO_106 (O_106,N_29060,N_29746);
or UO_107 (O_107,N_28968,N_28873);
nor UO_108 (O_108,N_29702,N_29687);
and UO_109 (O_109,N_29556,N_29523);
nor UO_110 (O_110,N_29899,N_29869);
nand UO_111 (O_111,N_29081,N_29468);
xnor UO_112 (O_112,N_29634,N_29287);
xnor UO_113 (O_113,N_29159,N_29777);
nor UO_114 (O_114,N_29703,N_29775);
and UO_115 (O_115,N_29852,N_29572);
nand UO_116 (O_116,N_29307,N_29538);
xnor UO_117 (O_117,N_29991,N_29979);
xor UO_118 (O_118,N_29383,N_28847);
xnor UO_119 (O_119,N_29040,N_29877);
and UO_120 (O_120,N_29492,N_29844);
or UO_121 (O_121,N_29693,N_29790);
xnor UO_122 (O_122,N_29881,N_29528);
xnor UO_123 (O_123,N_29078,N_29400);
xor UO_124 (O_124,N_29967,N_29989);
nand UO_125 (O_125,N_29047,N_28835);
and UO_126 (O_126,N_28821,N_29674);
nor UO_127 (O_127,N_29639,N_29716);
nor UO_128 (O_128,N_29665,N_29225);
or UO_129 (O_129,N_29960,N_29317);
nand UO_130 (O_130,N_29781,N_29767);
nand UO_131 (O_131,N_29661,N_29892);
nand UO_132 (O_132,N_29445,N_29722);
nand UO_133 (O_133,N_29671,N_29165);
or UO_134 (O_134,N_29823,N_29544);
and UO_135 (O_135,N_29123,N_29988);
xor UO_136 (O_136,N_29501,N_29870);
and UO_137 (O_137,N_29032,N_29831);
nor UO_138 (O_138,N_29124,N_28833);
xnor UO_139 (O_139,N_28993,N_29992);
nor UO_140 (O_140,N_28983,N_29226);
or UO_141 (O_141,N_29208,N_29948);
nor UO_142 (O_142,N_29405,N_29997);
or UO_143 (O_143,N_29982,N_28838);
or UO_144 (O_144,N_29148,N_29799);
xnor UO_145 (O_145,N_29943,N_29701);
or UO_146 (O_146,N_29654,N_29677);
nor UO_147 (O_147,N_29931,N_29658);
nand UO_148 (O_148,N_29531,N_29782);
xor UO_149 (O_149,N_29022,N_29440);
and UO_150 (O_150,N_29006,N_29973);
or UO_151 (O_151,N_29778,N_29905);
and UO_152 (O_152,N_29498,N_28834);
nor UO_153 (O_153,N_29950,N_29893);
and UO_154 (O_154,N_29431,N_29672);
and UO_155 (O_155,N_29278,N_29645);
nor UO_156 (O_156,N_29895,N_29534);
or UO_157 (O_157,N_29640,N_29944);
and UO_158 (O_158,N_29173,N_29712);
xnor UO_159 (O_159,N_29680,N_29753);
nand UO_160 (O_160,N_29017,N_28933);
or UO_161 (O_161,N_29076,N_29197);
nor UO_162 (O_162,N_28928,N_29630);
xnor UO_163 (O_163,N_29631,N_29872);
xnor UO_164 (O_164,N_29112,N_29332);
nand UO_165 (O_165,N_29084,N_29825);
and UO_166 (O_166,N_29227,N_29600);
or UO_167 (O_167,N_29773,N_28837);
nand UO_168 (O_168,N_29740,N_29099);
nand UO_169 (O_169,N_29564,N_29362);
xnor UO_170 (O_170,N_29725,N_29104);
xnor UO_171 (O_171,N_28907,N_29432);
nor UO_172 (O_172,N_28975,N_29422);
nor UO_173 (O_173,N_28952,N_29558);
or UO_174 (O_174,N_29082,N_29441);
xnor UO_175 (O_175,N_29632,N_29053);
xor UO_176 (O_176,N_29070,N_29541);
xnor UO_177 (O_177,N_29412,N_29126);
nor UO_178 (O_178,N_29837,N_29163);
nand UO_179 (O_179,N_28915,N_29884);
and UO_180 (O_180,N_28965,N_29326);
nand UO_181 (O_181,N_28802,N_28840);
xor UO_182 (O_182,N_29442,N_29954);
nand UO_183 (O_183,N_29919,N_29845);
xnor UO_184 (O_184,N_28902,N_29563);
nand UO_185 (O_185,N_29957,N_29223);
xnor UO_186 (O_186,N_29849,N_29801);
and UO_187 (O_187,N_29682,N_29283);
nand UO_188 (O_188,N_29560,N_29014);
xnor UO_189 (O_189,N_29325,N_29621);
nor UO_190 (O_190,N_29100,N_29411);
xnor UO_191 (O_191,N_29750,N_28875);
xor UO_192 (O_192,N_29388,N_29424);
or UO_193 (O_193,N_29366,N_28985);
xor UO_194 (O_194,N_29546,N_29248);
nor UO_195 (O_195,N_29584,N_28960);
or UO_196 (O_196,N_29588,N_29708);
or UO_197 (O_197,N_29407,N_28946);
or UO_198 (O_198,N_29368,N_29545);
xor UO_199 (O_199,N_28851,N_29127);
nor UO_200 (O_200,N_29952,N_28878);
xor UO_201 (O_201,N_29779,N_28816);
and UO_202 (O_202,N_29871,N_29265);
nor UO_203 (O_203,N_29276,N_28803);
nand UO_204 (O_204,N_29565,N_29056);
and UO_205 (O_205,N_29059,N_29808);
and UO_206 (O_206,N_29522,N_29499);
nor UO_207 (O_207,N_29914,N_29865);
and UO_208 (O_208,N_29793,N_29664);
nor UO_209 (O_209,N_29348,N_29548);
nand UO_210 (O_210,N_29513,N_29760);
or UO_211 (O_211,N_29254,N_29547);
or UO_212 (O_212,N_28848,N_29156);
or UO_213 (O_213,N_29365,N_29907);
or UO_214 (O_214,N_29994,N_29149);
nand UO_215 (O_215,N_29162,N_29771);
nor UO_216 (O_216,N_29524,N_28940);
xnor UO_217 (O_217,N_28935,N_29917);
xor UO_218 (O_218,N_28886,N_28846);
or UO_219 (O_219,N_29037,N_28832);
nand UO_220 (O_220,N_29243,N_29152);
xnor UO_221 (O_221,N_29819,N_29724);
nor UO_222 (O_222,N_29959,N_28995);
xnor UO_223 (O_223,N_29286,N_28973);
nand UO_224 (O_224,N_29280,N_29477);
nand UO_225 (O_225,N_29101,N_29655);
nor UO_226 (O_226,N_29700,N_29178);
nand UO_227 (O_227,N_29176,N_28822);
nand UO_228 (O_228,N_29316,N_29361);
or UO_229 (O_229,N_29755,N_28957);
xnor UO_230 (O_230,N_29590,N_29142);
nor UO_231 (O_231,N_29188,N_28879);
and UO_232 (O_232,N_29970,N_29587);
or UO_233 (O_233,N_29510,N_28810);
nor UO_234 (O_234,N_29138,N_28828);
or UO_235 (O_235,N_29706,N_29533);
and UO_236 (O_236,N_29515,N_29835);
or UO_237 (O_237,N_29312,N_29993);
or UO_238 (O_238,N_29372,N_29401);
nand UO_239 (O_239,N_28954,N_29652);
and UO_240 (O_240,N_29414,N_29471);
and UO_241 (O_241,N_29038,N_29489);
and UO_242 (O_242,N_29303,N_28805);
xnor UO_243 (O_243,N_28937,N_29238);
nor UO_244 (O_244,N_29216,N_29816);
nor UO_245 (O_245,N_29883,N_29986);
nand UO_246 (O_246,N_29641,N_29242);
and UO_247 (O_247,N_29798,N_29504);
or UO_248 (O_248,N_29610,N_29263);
and UO_249 (O_249,N_29615,N_29336);
and UO_250 (O_250,N_29484,N_29279);
nand UO_251 (O_251,N_29474,N_29031);
nor UO_252 (O_252,N_29268,N_29551);
xor UO_253 (O_253,N_29219,N_29250);
or UO_254 (O_254,N_29233,N_29939);
nand UO_255 (O_255,N_29091,N_29627);
xnor UO_256 (O_256,N_29670,N_28974);
xor UO_257 (O_257,N_29290,N_29071);
xor UO_258 (O_258,N_29315,N_29736);
or UO_259 (O_259,N_29007,N_29749);
xor UO_260 (O_260,N_29521,N_29302);
nor UO_261 (O_261,N_29864,N_29228);
and UO_262 (O_262,N_29281,N_29738);
or UO_263 (O_263,N_28842,N_29911);
nand UO_264 (O_264,N_28971,N_29354);
or UO_265 (O_265,N_29517,N_29763);
xor UO_266 (O_266,N_29063,N_28856);
nor UO_267 (O_267,N_29352,N_29026);
and UO_268 (O_268,N_29720,N_28992);
and UO_269 (O_269,N_29174,N_29304);
or UO_270 (O_270,N_29408,N_29927);
xnor UO_271 (O_271,N_28801,N_28934);
xnor UO_272 (O_272,N_29830,N_29244);
or UO_273 (O_273,N_29969,N_28984);
or UO_274 (O_274,N_28820,N_29984);
nor UO_275 (O_275,N_29399,N_29900);
and UO_276 (O_276,N_29920,N_29678);
and UO_277 (O_277,N_29618,N_29791);
nand UO_278 (O_278,N_29818,N_28884);
nand UO_279 (O_279,N_29622,N_29577);
xnor UO_280 (O_280,N_29451,N_29860);
and UO_281 (O_281,N_29262,N_29105);
nand UO_282 (O_282,N_29376,N_29673);
or UO_283 (O_283,N_29333,N_29301);
nor UO_284 (O_284,N_29848,N_29550);
and UO_285 (O_285,N_28912,N_28859);
nor UO_286 (O_286,N_28817,N_29935);
xor UO_287 (O_287,N_29814,N_28964);
and UO_288 (O_288,N_29043,N_29614);
and UO_289 (O_289,N_29586,N_29095);
nand UO_290 (O_290,N_29363,N_29386);
nor UO_291 (O_291,N_29956,N_29444);
nor UO_292 (O_292,N_29953,N_28904);
or UO_293 (O_293,N_29734,N_29805);
nor UO_294 (O_294,N_29481,N_29055);
and UO_295 (O_295,N_29200,N_29049);
or UO_296 (O_296,N_28929,N_29072);
or UO_297 (O_297,N_29874,N_29542);
or UO_298 (O_298,N_28932,N_29134);
nor UO_299 (O_299,N_29526,N_29393);
and UO_300 (O_300,N_29921,N_29008);
xor UO_301 (O_301,N_29118,N_29131);
nand UO_302 (O_302,N_29579,N_29462);
nand UO_303 (O_303,N_29446,N_29128);
or UO_304 (O_304,N_29635,N_29834);
and UO_305 (O_305,N_28897,N_29867);
or UO_306 (O_306,N_29483,N_29212);
nor UO_307 (O_307,N_29599,N_28877);
nor UO_308 (O_308,N_29604,N_28861);
nand UO_309 (O_309,N_29347,N_29506);
or UO_310 (O_310,N_29097,N_29025);
or UO_311 (O_311,N_29465,N_29794);
and UO_312 (O_312,N_29714,N_29253);
nand UO_313 (O_313,N_29052,N_29083);
nor UO_314 (O_314,N_29475,N_29229);
xor UO_315 (O_315,N_29274,N_29981);
nor UO_316 (O_316,N_29602,N_29685);
nand UO_317 (O_317,N_28959,N_29416);
xor UO_318 (O_318,N_29185,N_29882);
nor UO_319 (O_319,N_29027,N_29000);
or UO_320 (O_320,N_28892,N_29974);
or UO_321 (O_321,N_29976,N_29669);
and UO_322 (O_322,N_29643,N_29230);
nand UO_323 (O_323,N_29235,N_29941);
nand UO_324 (O_324,N_29811,N_28809);
and UO_325 (O_325,N_28917,N_29925);
or UO_326 (O_326,N_29010,N_29132);
nand UO_327 (O_327,N_29983,N_29309);
and UO_328 (O_328,N_29843,N_29497);
nor UO_329 (O_329,N_28963,N_29942);
nor UO_330 (O_330,N_29961,N_29769);
and UO_331 (O_331,N_28866,N_29257);
xnor UO_332 (O_332,N_29743,N_29494);
xnor UO_333 (O_333,N_29747,N_29146);
xor UO_334 (O_334,N_29154,N_29419);
nand UO_335 (O_335,N_28811,N_29897);
nor UO_336 (O_336,N_29291,N_29946);
or UO_337 (O_337,N_29135,N_29413);
and UO_338 (O_338,N_29215,N_29036);
and UO_339 (O_339,N_29491,N_29092);
or UO_340 (O_340,N_29241,N_29358);
or UO_341 (O_341,N_29886,N_28949);
nand UO_342 (O_342,N_29770,N_29158);
xnor UO_343 (O_343,N_28874,N_29486);
and UO_344 (O_344,N_29133,N_29539);
nand UO_345 (O_345,N_29820,N_29853);
and UO_346 (O_346,N_29757,N_29878);
or UO_347 (O_347,N_28827,N_29346);
and UO_348 (O_348,N_29727,N_29186);
or UO_349 (O_349,N_29862,N_29120);
or UO_350 (O_350,N_28890,N_29423);
xnor UO_351 (O_351,N_29530,N_29296);
xnor UO_352 (O_352,N_29744,N_29996);
xor UO_353 (O_353,N_29783,N_29057);
nor UO_354 (O_354,N_29536,N_29741);
nand UO_355 (O_355,N_29328,N_29576);
or UO_356 (O_356,N_29447,N_28950);
xnor UO_357 (O_357,N_29821,N_28989);
nor UO_358 (O_358,N_29205,N_29803);
or UO_359 (O_359,N_28920,N_29439);
and UO_360 (O_360,N_29394,N_29842);
and UO_361 (O_361,N_28981,N_29802);
and UO_362 (O_362,N_29175,N_29323);
nand UO_363 (O_363,N_29520,N_28841);
or UO_364 (O_364,N_29088,N_29718);
xor UO_365 (O_365,N_29567,N_28887);
or UO_366 (O_366,N_29169,N_29508);
and UO_367 (O_367,N_29113,N_28831);
or UO_368 (O_368,N_29792,N_29345);
nor UO_369 (O_369,N_29256,N_29479);
and UO_370 (O_370,N_29389,N_28916);
xnor UO_371 (O_371,N_29566,N_29894);
and UO_372 (O_372,N_29573,N_28865);
or UO_373 (O_373,N_29433,N_29181);
and UO_374 (O_374,N_29377,N_29535);
or UO_375 (O_375,N_29240,N_29916);
xor UO_376 (O_376,N_29766,N_29005);
xnor UO_377 (O_377,N_28893,N_29912);
xor UO_378 (O_378,N_29436,N_29659);
xnor UO_379 (O_379,N_29583,N_29272);
nand UO_380 (O_380,N_29768,N_29351);
nor UO_381 (O_381,N_29013,N_29633);
nand UO_382 (O_382,N_29107,N_29511);
and UO_383 (O_383,N_29694,N_29397);
xor UO_384 (O_384,N_29732,N_28931);
xor UO_385 (O_385,N_29540,N_29415);
nand UO_386 (O_386,N_29589,N_28988);
or UO_387 (O_387,N_29932,N_29838);
nand UO_388 (O_388,N_29255,N_29364);
or UO_389 (O_389,N_29666,N_28961);
or UO_390 (O_390,N_28858,N_29695);
xnor UO_391 (O_391,N_29730,N_28854);
and UO_392 (O_392,N_29245,N_28979);
or UO_393 (O_393,N_29663,N_29966);
and UO_394 (O_394,N_29660,N_29050);
nand UO_395 (O_395,N_29103,N_29448);
or UO_396 (O_396,N_28980,N_29898);
xor UO_397 (O_397,N_29143,N_29090);
and UO_398 (O_398,N_29086,N_28944);
or UO_399 (O_399,N_29199,N_29527);
nand UO_400 (O_400,N_29029,N_29409);
and UO_401 (O_401,N_29516,N_29815);
and UO_402 (O_402,N_29514,N_29136);
and UO_403 (O_403,N_29651,N_29866);
nand UO_404 (O_404,N_29139,N_29094);
xnor UO_405 (O_405,N_29252,N_29478);
nor UO_406 (O_406,N_29089,N_29875);
nor UO_407 (O_407,N_29529,N_29938);
nor UO_408 (O_408,N_29787,N_29473);
or UO_409 (O_409,N_29313,N_29653);
nor UO_410 (O_410,N_29889,N_29273);
nor UO_411 (O_411,N_29129,N_29839);
xnor UO_412 (O_412,N_29457,N_29469);
xnor UO_413 (O_413,N_29373,N_29282);
and UO_414 (O_414,N_29613,N_28966);
or UO_415 (O_415,N_29074,N_28939);
nor UO_416 (O_416,N_29595,N_29754);
or UO_417 (O_417,N_29723,N_28922);
nand UO_418 (O_418,N_28994,N_28888);
xor UO_419 (O_419,N_29789,N_28898);
and UO_420 (O_420,N_29574,N_29458);
or UO_421 (O_421,N_29192,N_28853);
or UO_422 (O_422,N_28882,N_28967);
or UO_423 (O_423,N_29041,N_28808);
and UO_424 (O_424,N_29319,N_29647);
nand UO_425 (O_425,N_29918,N_29553);
nor UO_426 (O_426,N_29951,N_29170);
nand UO_427 (O_427,N_29344,N_29668);
and UO_428 (O_428,N_29122,N_29962);
and UO_429 (O_429,N_29114,N_28825);
or UO_430 (O_430,N_29453,N_29237);
nor UO_431 (O_431,N_29251,N_29902);
and UO_432 (O_432,N_29308,N_29121);
xor UO_433 (O_433,N_28905,N_29906);
xor UO_434 (O_434,N_28977,N_28978);
or UO_435 (O_435,N_29607,N_29594);
nor UO_436 (O_436,N_28867,N_29045);
xnor UO_437 (O_437,N_28869,N_29698);
xnor UO_438 (O_438,N_29901,N_29809);
and UO_439 (O_439,N_29857,N_29157);
or UO_440 (O_440,N_29249,N_28925);
xnor UO_441 (O_441,N_29784,N_29314);
nand UO_442 (O_442,N_29758,N_28870);
xnor UO_443 (O_443,N_29507,N_28987);
or UO_444 (O_444,N_28895,N_29035);
or UO_445 (O_445,N_29561,N_29910);
or UO_446 (O_446,N_29636,N_29575);
and UO_447 (O_447,N_29487,N_29222);
xnor UO_448 (O_448,N_29689,N_28936);
xnor UO_449 (O_449,N_29196,N_29737);
nor UO_450 (O_450,N_28997,N_29195);
nand UO_451 (O_451,N_29780,N_29179);
or UO_452 (O_452,N_29578,N_29697);
or UO_453 (O_453,N_29184,N_29729);
xor UO_454 (O_454,N_29370,N_28813);
nand UO_455 (O_455,N_29106,N_29020);
xor UO_456 (O_456,N_29267,N_29868);
nor UO_457 (O_457,N_28889,N_29147);
xnor UO_458 (O_458,N_29648,N_29180);
xnor UO_459 (O_459,N_29271,N_29922);
and UO_460 (O_460,N_29353,N_29019);
or UO_461 (O_461,N_29608,N_29064);
nor UO_462 (O_462,N_29023,N_29357);
nor UO_463 (O_463,N_29340,N_29217);
and UO_464 (O_464,N_29145,N_29402);
nor UO_465 (O_465,N_29073,N_28862);
nand UO_466 (O_466,N_29616,N_28849);
or UO_467 (O_467,N_28947,N_29810);
nor UO_468 (O_468,N_29289,N_29936);
nand UO_469 (O_469,N_28899,N_28823);
nand UO_470 (O_470,N_29428,N_28910);
xor UO_471 (O_471,N_29125,N_28880);
xor UO_472 (O_472,N_29930,N_29965);
nand UO_473 (O_473,N_28927,N_29003);
nor UO_474 (O_474,N_29270,N_28996);
nor UO_475 (O_475,N_29260,N_29904);
nand UO_476 (O_476,N_29822,N_29840);
nand UO_477 (O_477,N_29688,N_29656);
xnor UO_478 (O_478,N_29463,N_29476);
xor UO_479 (O_479,N_29209,N_29024);
nor UO_480 (O_480,N_29876,N_29117);
xor UO_481 (O_481,N_28807,N_29828);
or UO_482 (O_482,N_29686,N_28972);
xor UO_483 (O_483,N_28826,N_29772);
xor UO_484 (O_484,N_29343,N_28881);
xor UO_485 (O_485,N_28956,N_29193);
or UO_486 (O_486,N_29331,N_29559);
xnor UO_487 (O_487,N_29880,N_29705);
nand UO_488 (O_488,N_29728,N_29735);
nor UO_489 (O_489,N_29009,N_29609);
nor UO_490 (O_490,N_29888,N_29676);
nand UO_491 (O_491,N_29467,N_29380);
and UO_492 (O_492,N_29980,N_28901);
or UO_493 (O_493,N_29806,N_28900);
xnor UO_494 (O_494,N_29324,N_29949);
nor UO_495 (O_495,N_29166,N_29829);
xnor UO_496 (O_496,N_29046,N_29620);
nand UO_497 (O_497,N_29582,N_29691);
nand UO_498 (O_498,N_29847,N_29360);
and UO_499 (O_499,N_29958,N_29731);
nand UO_500 (O_500,N_29454,N_29684);
or UO_501 (O_501,N_29042,N_29827);
nand UO_502 (O_502,N_29329,N_29410);
and UO_503 (O_503,N_29915,N_29667);
xor UO_504 (O_504,N_29532,N_29067);
nand UO_505 (O_505,N_29183,N_29239);
or UO_506 (O_506,N_29115,N_29715);
and UO_507 (O_507,N_29111,N_29642);
and UO_508 (O_508,N_29733,N_29855);
or UO_509 (O_509,N_29657,N_29649);
nand UO_510 (O_510,N_29334,N_29926);
xor UO_511 (O_511,N_29321,N_29080);
nor UO_512 (O_512,N_29034,N_29625);
and UO_513 (O_513,N_28924,N_29077);
and UO_514 (O_514,N_29603,N_29069);
and UO_515 (O_515,N_29488,N_29079);
and UO_516 (O_516,N_29623,N_29030);
xor UO_517 (O_517,N_29403,N_29382);
xnor UO_518 (O_518,N_28806,N_29617);
or UO_519 (O_519,N_29224,N_29937);
nand UO_520 (O_520,N_29624,N_29375);
xnor UO_521 (O_521,N_29745,N_29160);
and UO_522 (O_522,N_29776,N_29062);
and UO_523 (O_523,N_29742,N_28860);
and UO_524 (O_524,N_29093,N_29709);
xnor UO_525 (O_525,N_29028,N_29699);
or UO_526 (O_526,N_29033,N_29891);
and UO_527 (O_527,N_29707,N_28926);
xnor UO_528 (O_528,N_29039,N_28918);
nand UO_529 (O_529,N_29972,N_29861);
nor UO_530 (O_530,N_29299,N_29061);
nor UO_531 (O_531,N_29518,N_29519);
xnor UO_532 (O_532,N_29016,N_29221);
nor UO_533 (O_533,N_28976,N_29437);
and UO_534 (O_534,N_29150,N_29214);
nand UO_535 (O_535,N_29890,N_29977);
nor UO_536 (O_536,N_29443,N_29108);
xor UO_537 (O_537,N_29856,N_29396);
nand UO_538 (O_538,N_29194,N_28953);
nand UO_539 (O_539,N_29177,N_28969);
and UO_540 (O_540,N_29934,N_29182);
nor UO_541 (O_541,N_29430,N_29461);
nand UO_542 (O_542,N_29337,N_29288);
and UO_543 (O_543,N_29711,N_29119);
or UO_544 (O_544,N_29591,N_28800);
xnor UO_545 (O_545,N_29213,N_29385);
xnor UO_546 (O_546,N_29470,N_29999);
and UO_547 (O_547,N_29065,N_29978);
nand UO_548 (O_548,N_29384,N_29644);
nand UO_549 (O_549,N_28839,N_29417);
xor UO_550 (O_550,N_29846,N_28945);
and UO_551 (O_551,N_29975,N_29284);
nand UO_552 (O_552,N_28872,N_29098);
xor UO_553 (O_553,N_29502,N_29500);
xor UO_554 (O_554,N_29449,N_29598);
xor UO_555 (O_555,N_29130,N_29297);
or UO_556 (O_556,N_29555,N_29058);
xnor UO_557 (O_557,N_29675,N_28943);
nor UO_558 (O_558,N_28894,N_28876);
nand UO_559 (O_559,N_29455,N_29247);
or UO_560 (O_560,N_29141,N_29292);
and UO_561 (O_561,N_29066,N_28812);
xnor UO_562 (O_562,N_29998,N_29796);
xnor UO_563 (O_563,N_29929,N_29543);
or UO_564 (O_564,N_29761,N_28919);
nor UO_565 (O_565,N_29739,N_29330);
xnor UO_566 (O_566,N_29190,N_29629);
nor UO_567 (O_567,N_28958,N_29580);
nor UO_568 (O_568,N_29909,N_29164);
and UO_569 (O_569,N_29172,N_29887);
or UO_570 (O_570,N_29495,N_29786);
and UO_571 (O_571,N_28991,N_29295);
or UO_572 (O_572,N_29605,N_29859);
or UO_573 (O_573,N_28921,N_29619);
and UO_574 (O_574,N_29850,N_29525);
xor UO_575 (O_575,N_29168,N_29549);
nor UO_576 (O_576,N_29395,N_29923);
nand UO_577 (O_577,N_29051,N_29110);
xnor UO_578 (O_578,N_28850,N_29832);
nor UO_579 (O_579,N_29153,N_29490);
nor UO_580 (O_580,N_28942,N_29704);
and UO_581 (O_581,N_29807,N_28948);
xor UO_582 (O_582,N_28951,N_29116);
xor UO_583 (O_583,N_29369,N_29903);
and UO_584 (O_584,N_29341,N_29717);
or UO_585 (O_585,N_29719,N_29955);
and UO_586 (O_586,N_29774,N_29015);
or UO_587 (O_587,N_29144,N_28998);
nor UO_588 (O_588,N_29387,N_28830);
xor UO_589 (O_589,N_28911,N_29356);
nand UO_590 (O_590,N_29764,N_29557);
and UO_591 (O_591,N_28938,N_29751);
xnor UO_592 (O_592,N_29207,N_29562);
xor UO_593 (O_593,N_29198,N_29762);
and UO_594 (O_594,N_28814,N_29298);
or UO_595 (O_595,N_28955,N_29068);
xnor UO_596 (O_596,N_29628,N_29259);
or UO_597 (O_597,N_29662,N_28829);
xnor UO_598 (O_598,N_28962,N_29293);
and UO_599 (O_599,N_29054,N_29231);
nand UO_600 (O_600,N_29214,N_29529);
xor UO_601 (O_601,N_29083,N_29011);
or UO_602 (O_602,N_28983,N_29892);
and UO_603 (O_603,N_29635,N_29865);
nand UO_604 (O_604,N_29639,N_29794);
or UO_605 (O_605,N_29322,N_29695);
and UO_606 (O_606,N_29039,N_29193);
or UO_607 (O_607,N_28963,N_29730);
or UO_608 (O_608,N_29389,N_29524);
xnor UO_609 (O_609,N_29131,N_29500);
and UO_610 (O_610,N_29386,N_29850);
xor UO_611 (O_611,N_29445,N_28946);
and UO_612 (O_612,N_29021,N_29077);
or UO_613 (O_613,N_29229,N_28861);
and UO_614 (O_614,N_29092,N_29688);
and UO_615 (O_615,N_29914,N_29436);
xor UO_616 (O_616,N_29533,N_29936);
nor UO_617 (O_617,N_28984,N_29062);
nand UO_618 (O_618,N_29038,N_29061);
and UO_619 (O_619,N_29016,N_29922);
and UO_620 (O_620,N_29924,N_29427);
or UO_621 (O_621,N_29207,N_29360);
or UO_622 (O_622,N_29788,N_29731);
or UO_623 (O_623,N_28963,N_28842);
and UO_624 (O_624,N_28812,N_29988);
xnor UO_625 (O_625,N_29428,N_29167);
nor UO_626 (O_626,N_29099,N_29462);
nor UO_627 (O_627,N_28865,N_29357);
nand UO_628 (O_628,N_29597,N_29659);
or UO_629 (O_629,N_29028,N_29767);
nor UO_630 (O_630,N_29129,N_29488);
and UO_631 (O_631,N_29213,N_29367);
nor UO_632 (O_632,N_29541,N_29956);
nand UO_633 (O_633,N_29369,N_29847);
nor UO_634 (O_634,N_29473,N_28856);
and UO_635 (O_635,N_29565,N_29387);
nand UO_636 (O_636,N_29114,N_29450);
nor UO_637 (O_637,N_28967,N_29316);
or UO_638 (O_638,N_29009,N_28867);
and UO_639 (O_639,N_28954,N_28955);
or UO_640 (O_640,N_29468,N_29838);
nor UO_641 (O_641,N_29940,N_29195);
nor UO_642 (O_642,N_29395,N_28869);
and UO_643 (O_643,N_29935,N_28892);
nor UO_644 (O_644,N_29359,N_28829);
nand UO_645 (O_645,N_29257,N_29848);
and UO_646 (O_646,N_28947,N_29637);
nand UO_647 (O_647,N_29096,N_29021);
xnor UO_648 (O_648,N_28875,N_29313);
nor UO_649 (O_649,N_28837,N_29657);
nand UO_650 (O_650,N_29873,N_29715);
or UO_651 (O_651,N_29596,N_29278);
nand UO_652 (O_652,N_29888,N_29228);
nor UO_653 (O_653,N_29869,N_29315);
and UO_654 (O_654,N_28927,N_29500);
or UO_655 (O_655,N_28973,N_29768);
nor UO_656 (O_656,N_28849,N_29864);
and UO_657 (O_657,N_28847,N_29414);
and UO_658 (O_658,N_29148,N_29176);
nand UO_659 (O_659,N_29556,N_29670);
nand UO_660 (O_660,N_29928,N_29432);
nor UO_661 (O_661,N_28993,N_29126);
nand UO_662 (O_662,N_29830,N_29692);
nand UO_663 (O_663,N_29836,N_29287);
or UO_664 (O_664,N_29081,N_29118);
and UO_665 (O_665,N_29884,N_29936);
xnor UO_666 (O_666,N_28963,N_29772);
or UO_667 (O_667,N_29792,N_29922);
and UO_668 (O_668,N_29079,N_29930);
xnor UO_669 (O_669,N_29745,N_29045);
or UO_670 (O_670,N_29611,N_28863);
nand UO_671 (O_671,N_29484,N_29297);
or UO_672 (O_672,N_28883,N_29297);
or UO_673 (O_673,N_29904,N_29615);
nand UO_674 (O_674,N_29028,N_29156);
nand UO_675 (O_675,N_29915,N_29606);
or UO_676 (O_676,N_29375,N_29991);
and UO_677 (O_677,N_28862,N_29127);
nand UO_678 (O_678,N_29330,N_29735);
xnor UO_679 (O_679,N_28939,N_28987);
xor UO_680 (O_680,N_29812,N_29343);
nor UO_681 (O_681,N_29668,N_29776);
nor UO_682 (O_682,N_29475,N_29632);
and UO_683 (O_683,N_28897,N_29177);
and UO_684 (O_684,N_29318,N_28828);
or UO_685 (O_685,N_29660,N_29259);
xnor UO_686 (O_686,N_29591,N_28816);
xnor UO_687 (O_687,N_29524,N_28861);
nor UO_688 (O_688,N_29437,N_29887);
nand UO_689 (O_689,N_29252,N_28856);
xnor UO_690 (O_690,N_29258,N_29889);
nor UO_691 (O_691,N_29308,N_29605);
nor UO_692 (O_692,N_29200,N_29701);
nor UO_693 (O_693,N_29268,N_29119);
nand UO_694 (O_694,N_29776,N_29695);
or UO_695 (O_695,N_29571,N_29885);
nand UO_696 (O_696,N_29063,N_29082);
or UO_697 (O_697,N_29537,N_29542);
nand UO_698 (O_698,N_29805,N_29354);
and UO_699 (O_699,N_29853,N_28931);
xnor UO_700 (O_700,N_28954,N_29031);
nand UO_701 (O_701,N_29715,N_28894);
xnor UO_702 (O_702,N_28864,N_29420);
xnor UO_703 (O_703,N_29696,N_28982);
or UO_704 (O_704,N_29498,N_29559);
or UO_705 (O_705,N_29626,N_29624);
nand UO_706 (O_706,N_29611,N_28992);
nor UO_707 (O_707,N_29229,N_29784);
nor UO_708 (O_708,N_29808,N_29482);
xor UO_709 (O_709,N_28892,N_29844);
or UO_710 (O_710,N_29118,N_29681);
nor UO_711 (O_711,N_29614,N_29359);
nor UO_712 (O_712,N_28855,N_29302);
nand UO_713 (O_713,N_28925,N_29372);
or UO_714 (O_714,N_29768,N_29712);
xnor UO_715 (O_715,N_29065,N_28926);
nand UO_716 (O_716,N_29431,N_29250);
xor UO_717 (O_717,N_28941,N_29570);
xor UO_718 (O_718,N_28975,N_29936);
and UO_719 (O_719,N_29881,N_29491);
nand UO_720 (O_720,N_29022,N_29041);
nor UO_721 (O_721,N_29465,N_29298);
or UO_722 (O_722,N_29468,N_28909);
xor UO_723 (O_723,N_28806,N_29816);
nand UO_724 (O_724,N_29309,N_29459);
and UO_725 (O_725,N_29997,N_28862);
xnor UO_726 (O_726,N_29638,N_29432);
xor UO_727 (O_727,N_28909,N_29051);
and UO_728 (O_728,N_29068,N_29863);
nand UO_729 (O_729,N_28820,N_28972);
nand UO_730 (O_730,N_29760,N_28881);
xor UO_731 (O_731,N_29189,N_28912);
or UO_732 (O_732,N_28955,N_29658);
and UO_733 (O_733,N_29036,N_29980);
xor UO_734 (O_734,N_29308,N_29467);
nand UO_735 (O_735,N_28847,N_28971);
nand UO_736 (O_736,N_29443,N_29911);
and UO_737 (O_737,N_29695,N_29813);
nor UO_738 (O_738,N_29565,N_29330);
nand UO_739 (O_739,N_29529,N_29221);
nand UO_740 (O_740,N_29701,N_29570);
or UO_741 (O_741,N_29487,N_29168);
nor UO_742 (O_742,N_29371,N_29502);
nand UO_743 (O_743,N_29194,N_29970);
nor UO_744 (O_744,N_29324,N_29349);
xor UO_745 (O_745,N_29661,N_29579);
nor UO_746 (O_746,N_29414,N_29049);
or UO_747 (O_747,N_29472,N_29688);
nor UO_748 (O_748,N_29685,N_29813);
nand UO_749 (O_749,N_29829,N_29876);
nand UO_750 (O_750,N_29492,N_29039);
and UO_751 (O_751,N_29064,N_29975);
nor UO_752 (O_752,N_29056,N_29851);
and UO_753 (O_753,N_28936,N_28814);
nor UO_754 (O_754,N_29805,N_29435);
nor UO_755 (O_755,N_29583,N_29008);
xor UO_756 (O_756,N_29808,N_29130);
nand UO_757 (O_757,N_29689,N_29575);
nor UO_758 (O_758,N_29468,N_29880);
nor UO_759 (O_759,N_28969,N_29483);
nand UO_760 (O_760,N_29309,N_29935);
nand UO_761 (O_761,N_29226,N_29004);
and UO_762 (O_762,N_29451,N_29340);
or UO_763 (O_763,N_29819,N_29850);
and UO_764 (O_764,N_29344,N_28830);
and UO_765 (O_765,N_29513,N_29213);
nand UO_766 (O_766,N_29535,N_28971);
or UO_767 (O_767,N_29478,N_29339);
and UO_768 (O_768,N_29213,N_29713);
nand UO_769 (O_769,N_29864,N_28985);
and UO_770 (O_770,N_29249,N_29173);
xor UO_771 (O_771,N_29401,N_29550);
or UO_772 (O_772,N_29686,N_28990);
nand UO_773 (O_773,N_29971,N_28813);
xor UO_774 (O_774,N_29325,N_28886);
nor UO_775 (O_775,N_28867,N_29903);
nor UO_776 (O_776,N_29041,N_29480);
nand UO_777 (O_777,N_29565,N_29815);
and UO_778 (O_778,N_28821,N_29727);
and UO_779 (O_779,N_29194,N_28904);
nor UO_780 (O_780,N_29996,N_29653);
or UO_781 (O_781,N_29876,N_29560);
nand UO_782 (O_782,N_29161,N_29432);
and UO_783 (O_783,N_29907,N_28882);
xor UO_784 (O_784,N_29827,N_29770);
xor UO_785 (O_785,N_29959,N_29525);
xor UO_786 (O_786,N_29815,N_29704);
xor UO_787 (O_787,N_29059,N_29698);
xor UO_788 (O_788,N_29753,N_29066);
nand UO_789 (O_789,N_29419,N_29675);
and UO_790 (O_790,N_29635,N_29159);
nand UO_791 (O_791,N_29818,N_29371);
xnor UO_792 (O_792,N_29659,N_29473);
nand UO_793 (O_793,N_29927,N_29554);
and UO_794 (O_794,N_29269,N_29687);
xnor UO_795 (O_795,N_29601,N_29305);
or UO_796 (O_796,N_29478,N_29116);
xor UO_797 (O_797,N_29663,N_29324);
and UO_798 (O_798,N_29877,N_29116);
xnor UO_799 (O_799,N_28873,N_29261);
or UO_800 (O_800,N_29646,N_29463);
xnor UO_801 (O_801,N_29744,N_29189);
xnor UO_802 (O_802,N_29258,N_28967);
and UO_803 (O_803,N_28982,N_29348);
or UO_804 (O_804,N_29521,N_29149);
and UO_805 (O_805,N_28932,N_29582);
xor UO_806 (O_806,N_28911,N_29614);
or UO_807 (O_807,N_29163,N_29582);
nor UO_808 (O_808,N_29726,N_29947);
nand UO_809 (O_809,N_29306,N_29009);
nor UO_810 (O_810,N_29056,N_29450);
xnor UO_811 (O_811,N_29560,N_29625);
or UO_812 (O_812,N_29666,N_29895);
and UO_813 (O_813,N_29954,N_28801);
and UO_814 (O_814,N_29454,N_29049);
or UO_815 (O_815,N_29269,N_29473);
or UO_816 (O_816,N_29881,N_28973);
or UO_817 (O_817,N_29361,N_29040);
nand UO_818 (O_818,N_29325,N_29253);
or UO_819 (O_819,N_29454,N_29057);
or UO_820 (O_820,N_29569,N_29799);
nor UO_821 (O_821,N_29276,N_29207);
nor UO_822 (O_822,N_29571,N_29287);
nor UO_823 (O_823,N_29201,N_29191);
and UO_824 (O_824,N_29369,N_29108);
nand UO_825 (O_825,N_29245,N_29730);
or UO_826 (O_826,N_29661,N_29500);
or UO_827 (O_827,N_29552,N_29261);
or UO_828 (O_828,N_29996,N_29268);
and UO_829 (O_829,N_29789,N_29874);
nand UO_830 (O_830,N_29394,N_29731);
nor UO_831 (O_831,N_29892,N_29896);
xnor UO_832 (O_832,N_29790,N_29662);
and UO_833 (O_833,N_29144,N_28937);
xor UO_834 (O_834,N_29458,N_29769);
and UO_835 (O_835,N_29285,N_29630);
or UO_836 (O_836,N_29943,N_29386);
nand UO_837 (O_837,N_29887,N_29986);
xor UO_838 (O_838,N_29653,N_29476);
and UO_839 (O_839,N_29410,N_29767);
nand UO_840 (O_840,N_29561,N_29453);
and UO_841 (O_841,N_29706,N_29901);
xnor UO_842 (O_842,N_29720,N_29796);
nor UO_843 (O_843,N_29010,N_29511);
nand UO_844 (O_844,N_29946,N_29584);
and UO_845 (O_845,N_29879,N_29767);
nor UO_846 (O_846,N_29428,N_29254);
or UO_847 (O_847,N_29657,N_29832);
nand UO_848 (O_848,N_28895,N_29854);
and UO_849 (O_849,N_29945,N_29517);
or UO_850 (O_850,N_29578,N_29800);
and UO_851 (O_851,N_28991,N_29860);
nor UO_852 (O_852,N_29256,N_29933);
and UO_853 (O_853,N_29277,N_29238);
nand UO_854 (O_854,N_29656,N_28815);
and UO_855 (O_855,N_29635,N_28902);
and UO_856 (O_856,N_29831,N_29669);
nand UO_857 (O_857,N_29181,N_29435);
nand UO_858 (O_858,N_29073,N_29173);
xnor UO_859 (O_859,N_29346,N_29018);
or UO_860 (O_860,N_29701,N_29215);
and UO_861 (O_861,N_29749,N_29394);
or UO_862 (O_862,N_28849,N_29072);
and UO_863 (O_863,N_29746,N_29279);
and UO_864 (O_864,N_29894,N_29359);
or UO_865 (O_865,N_29205,N_29093);
nor UO_866 (O_866,N_29195,N_29861);
and UO_867 (O_867,N_29217,N_29273);
xnor UO_868 (O_868,N_28817,N_29343);
nor UO_869 (O_869,N_29856,N_29732);
nor UO_870 (O_870,N_29773,N_29162);
or UO_871 (O_871,N_28843,N_29345);
and UO_872 (O_872,N_28869,N_29862);
and UO_873 (O_873,N_29833,N_29876);
nand UO_874 (O_874,N_29084,N_28917);
xor UO_875 (O_875,N_29688,N_29839);
and UO_876 (O_876,N_29693,N_29284);
nand UO_877 (O_877,N_29269,N_29527);
nor UO_878 (O_878,N_29210,N_28936);
and UO_879 (O_879,N_29153,N_29964);
nor UO_880 (O_880,N_29915,N_29046);
nor UO_881 (O_881,N_29260,N_29863);
or UO_882 (O_882,N_29799,N_29034);
nor UO_883 (O_883,N_29969,N_28863);
xnor UO_884 (O_884,N_29965,N_29083);
or UO_885 (O_885,N_29377,N_29647);
nand UO_886 (O_886,N_29497,N_29895);
or UO_887 (O_887,N_29311,N_29307);
or UO_888 (O_888,N_28894,N_29264);
nand UO_889 (O_889,N_29470,N_29435);
xor UO_890 (O_890,N_29564,N_29854);
or UO_891 (O_891,N_29961,N_29411);
and UO_892 (O_892,N_29994,N_29477);
or UO_893 (O_893,N_28910,N_28912);
or UO_894 (O_894,N_29513,N_29769);
or UO_895 (O_895,N_29903,N_29373);
nand UO_896 (O_896,N_29545,N_29982);
and UO_897 (O_897,N_29131,N_29818);
nor UO_898 (O_898,N_29440,N_29505);
nand UO_899 (O_899,N_28803,N_29959);
and UO_900 (O_900,N_29073,N_28985);
nor UO_901 (O_901,N_29147,N_29102);
xor UO_902 (O_902,N_29604,N_29924);
and UO_903 (O_903,N_28838,N_28886);
nand UO_904 (O_904,N_29332,N_29006);
nor UO_905 (O_905,N_29111,N_29208);
nor UO_906 (O_906,N_29062,N_29972);
xnor UO_907 (O_907,N_29676,N_29408);
nand UO_908 (O_908,N_29647,N_29679);
or UO_909 (O_909,N_29591,N_29517);
nand UO_910 (O_910,N_29615,N_29549);
nor UO_911 (O_911,N_29296,N_28899);
nand UO_912 (O_912,N_29139,N_29312);
and UO_913 (O_913,N_29737,N_28944);
xor UO_914 (O_914,N_29887,N_29643);
xor UO_915 (O_915,N_29186,N_28857);
xor UO_916 (O_916,N_29157,N_28949);
nor UO_917 (O_917,N_28993,N_29181);
nor UO_918 (O_918,N_29660,N_29946);
and UO_919 (O_919,N_29041,N_29759);
nand UO_920 (O_920,N_28836,N_29192);
and UO_921 (O_921,N_28981,N_28919);
xnor UO_922 (O_922,N_29303,N_29567);
nand UO_923 (O_923,N_28802,N_29317);
nor UO_924 (O_924,N_29285,N_29717);
xnor UO_925 (O_925,N_29136,N_29158);
nand UO_926 (O_926,N_29792,N_29775);
xor UO_927 (O_927,N_29769,N_29822);
nand UO_928 (O_928,N_29142,N_29751);
and UO_929 (O_929,N_29752,N_29657);
nor UO_930 (O_930,N_29884,N_29521);
xnor UO_931 (O_931,N_29236,N_28895);
nor UO_932 (O_932,N_29247,N_28919);
and UO_933 (O_933,N_29334,N_29626);
nor UO_934 (O_934,N_29893,N_29041);
and UO_935 (O_935,N_29225,N_28984);
nand UO_936 (O_936,N_29103,N_29888);
and UO_937 (O_937,N_29672,N_29460);
or UO_938 (O_938,N_29229,N_29600);
and UO_939 (O_939,N_29536,N_28864);
nand UO_940 (O_940,N_29039,N_29983);
or UO_941 (O_941,N_29107,N_29267);
xnor UO_942 (O_942,N_29608,N_29203);
or UO_943 (O_943,N_29205,N_29495);
xor UO_944 (O_944,N_29583,N_29991);
xor UO_945 (O_945,N_29003,N_28833);
nor UO_946 (O_946,N_29369,N_29002);
and UO_947 (O_947,N_29618,N_29934);
xor UO_948 (O_948,N_28948,N_29524);
and UO_949 (O_949,N_29448,N_29701);
nor UO_950 (O_950,N_29259,N_29640);
nor UO_951 (O_951,N_29121,N_28856);
and UO_952 (O_952,N_29321,N_29767);
xor UO_953 (O_953,N_29950,N_29275);
or UO_954 (O_954,N_29709,N_29859);
xor UO_955 (O_955,N_29096,N_29560);
nor UO_956 (O_956,N_29380,N_29890);
nand UO_957 (O_957,N_29501,N_29964);
nor UO_958 (O_958,N_29677,N_28853);
nand UO_959 (O_959,N_29513,N_29940);
and UO_960 (O_960,N_29283,N_29602);
nor UO_961 (O_961,N_28987,N_29745);
nand UO_962 (O_962,N_28973,N_29745);
xor UO_963 (O_963,N_29174,N_29281);
xnor UO_964 (O_964,N_29135,N_29102);
nor UO_965 (O_965,N_29221,N_29394);
or UO_966 (O_966,N_29660,N_28986);
nand UO_967 (O_967,N_29624,N_29338);
or UO_968 (O_968,N_29517,N_29908);
nand UO_969 (O_969,N_29845,N_29018);
or UO_970 (O_970,N_29128,N_29165);
nand UO_971 (O_971,N_29494,N_28958);
or UO_972 (O_972,N_29510,N_29122);
or UO_973 (O_973,N_29742,N_29137);
or UO_974 (O_974,N_29463,N_28969);
and UO_975 (O_975,N_29485,N_29882);
nand UO_976 (O_976,N_29801,N_28861);
or UO_977 (O_977,N_29299,N_29533);
xnor UO_978 (O_978,N_29019,N_29256);
nand UO_979 (O_979,N_29957,N_28863);
and UO_980 (O_980,N_28917,N_29572);
and UO_981 (O_981,N_29816,N_29116);
xnor UO_982 (O_982,N_29005,N_29070);
or UO_983 (O_983,N_29652,N_29591);
or UO_984 (O_984,N_29787,N_29052);
nand UO_985 (O_985,N_28946,N_29234);
and UO_986 (O_986,N_29390,N_29563);
or UO_987 (O_987,N_29135,N_29597);
and UO_988 (O_988,N_29622,N_29271);
nand UO_989 (O_989,N_29487,N_29476);
or UO_990 (O_990,N_29343,N_28823);
xor UO_991 (O_991,N_29727,N_29730);
or UO_992 (O_992,N_29702,N_29034);
nor UO_993 (O_993,N_29574,N_29160);
xor UO_994 (O_994,N_29629,N_29046);
and UO_995 (O_995,N_29526,N_29904);
and UO_996 (O_996,N_29991,N_29434);
or UO_997 (O_997,N_29847,N_29618);
nor UO_998 (O_998,N_29094,N_29252);
or UO_999 (O_999,N_29844,N_29227);
nor UO_1000 (O_1000,N_28814,N_28972);
and UO_1001 (O_1001,N_29607,N_29268);
nand UO_1002 (O_1002,N_28904,N_29440);
nand UO_1003 (O_1003,N_29285,N_29627);
nor UO_1004 (O_1004,N_29817,N_29083);
nand UO_1005 (O_1005,N_28944,N_29124);
xnor UO_1006 (O_1006,N_29926,N_29433);
and UO_1007 (O_1007,N_29019,N_29530);
nand UO_1008 (O_1008,N_29356,N_29460);
or UO_1009 (O_1009,N_28933,N_29193);
and UO_1010 (O_1010,N_29872,N_29470);
nor UO_1011 (O_1011,N_29416,N_29739);
or UO_1012 (O_1012,N_29159,N_29709);
xor UO_1013 (O_1013,N_29375,N_29645);
xor UO_1014 (O_1014,N_28962,N_29357);
xnor UO_1015 (O_1015,N_29443,N_29323);
and UO_1016 (O_1016,N_28978,N_29992);
nand UO_1017 (O_1017,N_28836,N_29353);
and UO_1018 (O_1018,N_29081,N_28902);
xor UO_1019 (O_1019,N_29113,N_28947);
and UO_1020 (O_1020,N_29759,N_29173);
or UO_1021 (O_1021,N_29828,N_28875);
and UO_1022 (O_1022,N_29611,N_28882);
nand UO_1023 (O_1023,N_29888,N_28871);
and UO_1024 (O_1024,N_29557,N_29158);
nand UO_1025 (O_1025,N_29422,N_29578);
nand UO_1026 (O_1026,N_29254,N_29194);
xnor UO_1027 (O_1027,N_29239,N_29157);
and UO_1028 (O_1028,N_29805,N_29548);
nand UO_1029 (O_1029,N_29309,N_29706);
or UO_1030 (O_1030,N_29250,N_29132);
xor UO_1031 (O_1031,N_29651,N_29753);
nor UO_1032 (O_1032,N_29223,N_29721);
nand UO_1033 (O_1033,N_29610,N_29996);
nand UO_1034 (O_1034,N_29981,N_29705);
nand UO_1035 (O_1035,N_29472,N_29421);
xnor UO_1036 (O_1036,N_29517,N_29379);
and UO_1037 (O_1037,N_28961,N_29282);
xor UO_1038 (O_1038,N_29121,N_29960);
nor UO_1039 (O_1039,N_29969,N_29798);
nand UO_1040 (O_1040,N_28912,N_29379);
and UO_1041 (O_1041,N_29938,N_29865);
nand UO_1042 (O_1042,N_29523,N_29134);
xnor UO_1043 (O_1043,N_29486,N_29947);
and UO_1044 (O_1044,N_29321,N_29869);
nor UO_1045 (O_1045,N_28875,N_29610);
and UO_1046 (O_1046,N_29883,N_29430);
nand UO_1047 (O_1047,N_28880,N_29694);
or UO_1048 (O_1048,N_28989,N_28945);
or UO_1049 (O_1049,N_29138,N_29201);
xor UO_1050 (O_1050,N_29130,N_28826);
nor UO_1051 (O_1051,N_29087,N_29841);
xor UO_1052 (O_1052,N_29543,N_29603);
nand UO_1053 (O_1053,N_29799,N_29326);
and UO_1054 (O_1054,N_29110,N_29377);
nor UO_1055 (O_1055,N_29537,N_29491);
nor UO_1056 (O_1056,N_29905,N_29744);
nor UO_1057 (O_1057,N_29890,N_28933);
nor UO_1058 (O_1058,N_29735,N_29251);
xor UO_1059 (O_1059,N_29930,N_29099);
xnor UO_1060 (O_1060,N_29739,N_28856);
xor UO_1061 (O_1061,N_29795,N_29259);
nand UO_1062 (O_1062,N_28878,N_29592);
nor UO_1063 (O_1063,N_29132,N_29632);
nand UO_1064 (O_1064,N_29006,N_29235);
nor UO_1065 (O_1065,N_29683,N_29716);
xor UO_1066 (O_1066,N_29005,N_29401);
nand UO_1067 (O_1067,N_28960,N_29332);
nor UO_1068 (O_1068,N_29370,N_29262);
or UO_1069 (O_1069,N_29713,N_29667);
and UO_1070 (O_1070,N_29221,N_29477);
and UO_1071 (O_1071,N_29394,N_29720);
and UO_1072 (O_1072,N_28818,N_29761);
xnor UO_1073 (O_1073,N_29496,N_29343);
xor UO_1074 (O_1074,N_29322,N_29892);
xor UO_1075 (O_1075,N_29936,N_28870);
xor UO_1076 (O_1076,N_29142,N_29869);
nor UO_1077 (O_1077,N_29609,N_29906);
and UO_1078 (O_1078,N_28940,N_29577);
or UO_1079 (O_1079,N_29958,N_29730);
and UO_1080 (O_1080,N_29057,N_29876);
nor UO_1081 (O_1081,N_29065,N_29583);
nor UO_1082 (O_1082,N_29101,N_29703);
or UO_1083 (O_1083,N_29837,N_29207);
and UO_1084 (O_1084,N_29157,N_29672);
xnor UO_1085 (O_1085,N_28923,N_29029);
nand UO_1086 (O_1086,N_29170,N_28952);
xor UO_1087 (O_1087,N_29939,N_28837);
or UO_1088 (O_1088,N_29842,N_29541);
nand UO_1089 (O_1089,N_29754,N_29850);
nand UO_1090 (O_1090,N_29252,N_29317);
nand UO_1091 (O_1091,N_29369,N_28824);
nand UO_1092 (O_1092,N_29848,N_28943);
xor UO_1093 (O_1093,N_29259,N_29684);
or UO_1094 (O_1094,N_28958,N_29862);
and UO_1095 (O_1095,N_29837,N_29999);
or UO_1096 (O_1096,N_28869,N_29633);
or UO_1097 (O_1097,N_29234,N_28981);
or UO_1098 (O_1098,N_29239,N_29801);
or UO_1099 (O_1099,N_29654,N_29907);
nand UO_1100 (O_1100,N_29702,N_29928);
or UO_1101 (O_1101,N_29859,N_29579);
xnor UO_1102 (O_1102,N_29453,N_28807);
nor UO_1103 (O_1103,N_29498,N_29422);
nor UO_1104 (O_1104,N_29383,N_29774);
nor UO_1105 (O_1105,N_29305,N_28897);
and UO_1106 (O_1106,N_29584,N_29070);
or UO_1107 (O_1107,N_29993,N_29953);
nand UO_1108 (O_1108,N_29597,N_29955);
nand UO_1109 (O_1109,N_29628,N_29358);
or UO_1110 (O_1110,N_28839,N_29404);
and UO_1111 (O_1111,N_29313,N_29152);
nand UO_1112 (O_1112,N_29373,N_28929);
nor UO_1113 (O_1113,N_29722,N_29728);
and UO_1114 (O_1114,N_29951,N_28954);
xnor UO_1115 (O_1115,N_28906,N_29943);
or UO_1116 (O_1116,N_29070,N_29635);
nand UO_1117 (O_1117,N_29816,N_29435);
or UO_1118 (O_1118,N_28980,N_28936);
xnor UO_1119 (O_1119,N_29417,N_29704);
or UO_1120 (O_1120,N_29560,N_29307);
and UO_1121 (O_1121,N_29607,N_29062);
nand UO_1122 (O_1122,N_29483,N_28881);
xor UO_1123 (O_1123,N_28936,N_28994);
and UO_1124 (O_1124,N_29312,N_29321);
nand UO_1125 (O_1125,N_28983,N_28988);
nor UO_1126 (O_1126,N_29084,N_29977);
or UO_1127 (O_1127,N_29167,N_29387);
and UO_1128 (O_1128,N_29198,N_28973);
nand UO_1129 (O_1129,N_29494,N_29480);
and UO_1130 (O_1130,N_29687,N_29518);
nor UO_1131 (O_1131,N_28904,N_29340);
or UO_1132 (O_1132,N_29889,N_29277);
and UO_1133 (O_1133,N_29284,N_29041);
nand UO_1134 (O_1134,N_29827,N_29503);
nor UO_1135 (O_1135,N_28920,N_29293);
nor UO_1136 (O_1136,N_29281,N_29847);
nor UO_1137 (O_1137,N_29469,N_29644);
nand UO_1138 (O_1138,N_29136,N_29833);
nand UO_1139 (O_1139,N_29997,N_29924);
xnor UO_1140 (O_1140,N_28878,N_29880);
and UO_1141 (O_1141,N_28887,N_28819);
and UO_1142 (O_1142,N_29913,N_28872);
and UO_1143 (O_1143,N_28879,N_29203);
and UO_1144 (O_1144,N_29035,N_29653);
or UO_1145 (O_1145,N_29050,N_28808);
nand UO_1146 (O_1146,N_29845,N_29211);
nand UO_1147 (O_1147,N_29479,N_29203);
nor UO_1148 (O_1148,N_29498,N_29814);
xnor UO_1149 (O_1149,N_29756,N_29840);
nor UO_1150 (O_1150,N_29670,N_29865);
nor UO_1151 (O_1151,N_29804,N_29377);
or UO_1152 (O_1152,N_28858,N_29651);
nor UO_1153 (O_1153,N_29673,N_29964);
nor UO_1154 (O_1154,N_29138,N_29743);
xor UO_1155 (O_1155,N_29145,N_29797);
and UO_1156 (O_1156,N_29925,N_29159);
and UO_1157 (O_1157,N_29380,N_29691);
xnor UO_1158 (O_1158,N_29262,N_29114);
nor UO_1159 (O_1159,N_28860,N_29572);
nor UO_1160 (O_1160,N_28816,N_29367);
xor UO_1161 (O_1161,N_29935,N_29617);
and UO_1162 (O_1162,N_29489,N_29158);
or UO_1163 (O_1163,N_28950,N_29043);
xor UO_1164 (O_1164,N_28874,N_29168);
nor UO_1165 (O_1165,N_29708,N_29827);
xor UO_1166 (O_1166,N_29057,N_29709);
xnor UO_1167 (O_1167,N_29263,N_28876);
xor UO_1168 (O_1168,N_29648,N_29449);
nand UO_1169 (O_1169,N_29571,N_29618);
xor UO_1170 (O_1170,N_29653,N_29898);
and UO_1171 (O_1171,N_29926,N_29967);
xor UO_1172 (O_1172,N_29696,N_28873);
or UO_1173 (O_1173,N_28800,N_29353);
or UO_1174 (O_1174,N_29860,N_29174);
xnor UO_1175 (O_1175,N_29588,N_29746);
nand UO_1176 (O_1176,N_29830,N_29192);
xnor UO_1177 (O_1177,N_29487,N_28934);
or UO_1178 (O_1178,N_29388,N_28914);
and UO_1179 (O_1179,N_29126,N_29771);
nor UO_1180 (O_1180,N_29244,N_29236);
and UO_1181 (O_1181,N_29551,N_29544);
and UO_1182 (O_1182,N_29836,N_29095);
and UO_1183 (O_1183,N_29022,N_29404);
xor UO_1184 (O_1184,N_28913,N_29190);
nand UO_1185 (O_1185,N_29080,N_29351);
xor UO_1186 (O_1186,N_29863,N_28848);
xor UO_1187 (O_1187,N_29331,N_29094);
nor UO_1188 (O_1188,N_29332,N_29052);
and UO_1189 (O_1189,N_29905,N_29439);
and UO_1190 (O_1190,N_29341,N_29625);
nor UO_1191 (O_1191,N_29969,N_29523);
and UO_1192 (O_1192,N_29335,N_28879);
nand UO_1193 (O_1193,N_29556,N_29126);
and UO_1194 (O_1194,N_28967,N_29827);
nor UO_1195 (O_1195,N_29337,N_29009);
and UO_1196 (O_1196,N_29668,N_29209);
nor UO_1197 (O_1197,N_28802,N_29759);
nor UO_1198 (O_1198,N_28915,N_29516);
nor UO_1199 (O_1199,N_28968,N_29775);
nand UO_1200 (O_1200,N_29139,N_29323);
nand UO_1201 (O_1201,N_29669,N_29192);
nand UO_1202 (O_1202,N_29954,N_29467);
xnor UO_1203 (O_1203,N_29473,N_29381);
and UO_1204 (O_1204,N_29899,N_29943);
nor UO_1205 (O_1205,N_29458,N_29137);
nand UO_1206 (O_1206,N_29394,N_29920);
and UO_1207 (O_1207,N_29126,N_29529);
xnor UO_1208 (O_1208,N_29067,N_29132);
and UO_1209 (O_1209,N_28927,N_29160);
or UO_1210 (O_1210,N_29195,N_29438);
and UO_1211 (O_1211,N_29239,N_29882);
nand UO_1212 (O_1212,N_29508,N_29686);
nor UO_1213 (O_1213,N_29621,N_29361);
and UO_1214 (O_1214,N_29589,N_29375);
nor UO_1215 (O_1215,N_29306,N_29754);
xor UO_1216 (O_1216,N_29910,N_29862);
xor UO_1217 (O_1217,N_28824,N_29532);
xor UO_1218 (O_1218,N_29660,N_28966);
nor UO_1219 (O_1219,N_28963,N_29598);
and UO_1220 (O_1220,N_29196,N_29604);
and UO_1221 (O_1221,N_29039,N_28935);
nand UO_1222 (O_1222,N_29372,N_29422);
xor UO_1223 (O_1223,N_29958,N_29118);
or UO_1224 (O_1224,N_29134,N_29145);
nor UO_1225 (O_1225,N_29746,N_29309);
nand UO_1226 (O_1226,N_29380,N_28968);
nand UO_1227 (O_1227,N_29176,N_29923);
nand UO_1228 (O_1228,N_29981,N_29578);
nand UO_1229 (O_1229,N_29503,N_29632);
nor UO_1230 (O_1230,N_29219,N_28817);
or UO_1231 (O_1231,N_28897,N_29084);
nor UO_1232 (O_1232,N_29743,N_29328);
xor UO_1233 (O_1233,N_29817,N_29905);
and UO_1234 (O_1234,N_29247,N_29389);
nor UO_1235 (O_1235,N_29321,N_29320);
xnor UO_1236 (O_1236,N_29095,N_29169);
xnor UO_1237 (O_1237,N_29541,N_29372);
nand UO_1238 (O_1238,N_29804,N_29452);
or UO_1239 (O_1239,N_29518,N_29869);
xnor UO_1240 (O_1240,N_29930,N_29294);
or UO_1241 (O_1241,N_28956,N_28821);
nand UO_1242 (O_1242,N_29009,N_28837);
or UO_1243 (O_1243,N_29201,N_29686);
nand UO_1244 (O_1244,N_29204,N_29542);
xor UO_1245 (O_1245,N_29403,N_29693);
and UO_1246 (O_1246,N_29318,N_28918);
nor UO_1247 (O_1247,N_29949,N_28825);
nand UO_1248 (O_1248,N_29693,N_29525);
nand UO_1249 (O_1249,N_29500,N_29373);
nand UO_1250 (O_1250,N_29091,N_29482);
xor UO_1251 (O_1251,N_29991,N_28863);
and UO_1252 (O_1252,N_29435,N_29827);
or UO_1253 (O_1253,N_29009,N_29149);
and UO_1254 (O_1254,N_29342,N_29007);
nor UO_1255 (O_1255,N_29464,N_29103);
xnor UO_1256 (O_1256,N_29891,N_29594);
xor UO_1257 (O_1257,N_29571,N_28921);
nor UO_1258 (O_1258,N_28981,N_28878);
nand UO_1259 (O_1259,N_29118,N_29176);
nor UO_1260 (O_1260,N_29993,N_29334);
xor UO_1261 (O_1261,N_29061,N_28981);
and UO_1262 (O_1262,N_29181,N_28836);
xnor UO_1263 (O_1263,N_29497,N_28856);
xnor UO_1264 (O_1264,N_29454,N_29000);
nand UO_1265 (O_1265,N_29917,N_29049);
nor UO_1266 (O_1266,N_28853,N_29465);
or UO_1267 (O_1267,N_29665,N_28951);
or UO_1268 (O_1268,N_28939,N_29467);
nand UO_1269 (O_1269,N_29108,N_29106);
and UO_1270 (O_1270,N_29568,N_29928);
or UO_1271 (O_1271,N_28944,N_29739);
nand UO_1272 (O_1272,N_29337,N_28942);
xnor UO_1273 (O_1273,N_29318,N_28945);
and UO_1274 (O_1274,N_29410,N_29501);
or UO_1275 (O_1275,N_29238,N_29522);
xor UO_1276 (O_1276,N_29798,N_28892);
nor UO_1277 (O_1277,N_29650,N_29547);
nand UO_1278 (O_1278,N_29776,N_29761);
and UO_1279 (O_1279,N_29850,N_28848);
and UO_1280 (O_1280,N_29939,N_29143);
or UO_1281 (O_1281,N_29261,N_28802);
and UO_1282 (O_1282,N_29794,N_29614);
and UO_1283 (O_1283,N_28866,N_29488);
or UO_1284 (O_1284,N_29394,N_29936);
or UO_1285 (O_1285,N_29325,N_29148);
xnor UO_1286 (O_1286,N_29110,N_28987);
or UO_1287 (O_1287,N_29666,N_29893);
nor UO_1288 (O_1288,N_29671,N_29059);
nand UO_1289 (O_1289,N_29402,N_29860);
xor UO_1290 (O_1290,N_29853,N_29443);
and UO_1291 (O_1291,N_29768,N_29675);
nor UO_1292 (O_1292,N_29578,N_29690);
nand UO_1293 (O_1293,N_29670,N_28993);
and UO_1294 (O_1294,N_28823,N_29223);
or UO_1295 (O_1295,N_29829,N_28892);
and UO_1296 (O_1296,N_28935,N_29047);
xnor UO_1297 (O_1297,N_29861,N_29227);
or UO_1298 (O_1298,N_29722,N_28857);
nand UO_1299 (O_1299,N_28880,N_29315);
and UO_1300 (O_1300,N_29602,N_29321);
nand UO_1301 (O_1301,N_29991,N_29609);
or UO_1302 (O_1302,N_29269,N_28829);
nand UO_1303 (O_1303,N_29543,N_29080);
nor UO_1304 (O_1304,N_29696,N_29922);
nor UO_1305 (O_1305,N_29199,N_29875);
and UO_1306 (O_1306,N_29029,N_29542);
xor UO_1307 (O_1307,N_29440,N_28894);
nand UO_1308 (O_1308,N_29396,N_28846);
xor UO_1309 (O_1309,N_28895,N_29075);
xor UO_1310 (O_1310,N_29735,N_29953);
and UO_1311 (O_1311,N_29311,N_29841);
xor UO_1312 (O_1312,N_29874,N_29558);
or UO_1313 (O_1313,N_29189,N_29619);
xnor UO_1314 (O_1314,N_29671,N_28959);
xor UO_1315 (O_1315,N_29495,N_29284);
nor UO_1316 (O_1316,N_29761,N_29705);
and UO_1317 (O_1317,N_29986,N_29640);
nand UO_1318 (O_1318,N_29246,N_29898);
xor UO_1319 (O_1319,N_29906,N_29669);
or UO_1320 (O_1320,N_28902,N_29790);
xor UO_1321 (O_1321,N_29521,N_29601);
xnor UO_1322 (O_1322,N_28959,N_29347);
nand UO_1323 (O_1323,N_29738,N_29828);
or UO_1324 (O_1324,N_29938,N_29877);
and UO_1325 (O_1325,N_29841,N_29991);
nor UO_1326 (O_1326,N_29585,N_29002);
or UO_1327 (O_1327,N_29735,N_29936);
nand UO_1328 (O_1328,N_29921,N_28974);
nor UO_1329 (O_1329,N_28945,N_29561);
xor UO_1330 (O_1330,N_29027,N_29060);
and UO_1331 (O_1331,N_29701,N_29378);
nand UO_1332 (O_1332,N_29290,N_29380);
xor UO_1333 (O_1333,N_29137,N_29312);
nor UO_1334 (O_1334,N_29989,N_29154);
or UO_1335 (O_1335,N_29634,N_29607);
or UO_1336 (O_1336,N_29162,N_29903);
nor UO_1337 (O_1337,N_29488,N_28988);
and UO_1338 (O_1338,N_29310,N_29976);
and UO_1339 (O_1339,N_29725,N_29238);
xor UO_1340 (O_1340,N_29586,N_29847);
or UO_1341 (O_1341,N_29146,N_28880);
or UO_1342 (O_1342,N_29708,N_29872);
xnor UO_1343 (O_1343,N_29329,N_28889);
and UO_1344 (O_1344,N_29569,N_29826);
and UO_1345 (O_1345,N_29287,N_29919);
nor UO_1346 (O_1346,N_29306,N_28984);
nand UO_1347 (O_1347,N_29168,N_29281);
xor UO_1348 (O_1348,N_29844,N_29957);
nor UO_1349 (O_1349,N_29828,N_29316);
nand UO_1350 (O_1350,N_29956,N_29520);
and UO_1351 (O_1351,N_28901,N_29498);
and UO_1352 (O_1352,N_29849,N_29828);
nand UO_1353 (O_1353,N_29894,N_29792);
and UO_1354 (O_1354,N_29224,N_29556);
nand UO_1355 (O_1355,N_29574,N_29860);
and UO_1356 (O_1356,N_29516,N_28927);
xor UO_1357 (O_1357,N_29823,N_29908);
and UO_1358 (O_1358,N_28960,N_28907);
or UO_1359 (O_1359,N_29786,N_29374);
or UO_1360 (O_1360,N_29418,N_29095);
or UO_1361 (O_1361,N_29221,N_29663);
nor UO_1362 (O_1362,N_29277,N_29102);
nand UO_1363 (O_1363,N_29526,N_29494);
or UO_1364 (O_1364,N_29709,N_29023);
xor UO_1365 (O_1365,N_29598,N_29716);
nand UO_1366 (O_1366,N_28836,N_29888);
and UO_1367 (O_1367,N_29019,N_29381);
xor UO_1368 (O_1368,N_29986,N_29728);
nor UO_1369 (O_1369,N_29584,N_29335);
nor UO_1370 (O_1370,N_29586,N_29912);
nand UO_1371 (O_1371,N_29655,N_28915);
or UO_1372 (O_1372,N_29809,N_29866);
xnor UO_1373 (O_1373,N_29201,N_29236);
nor UO_1374 (O_1374,N_29469,N_29906);
and UO_1375 (O_1375,N_29597,N_29080);
and UO_1376 (O_1376,N_29150,N_29269);
and UO_1377 (O_1377,N_29319,N_29538);
nor UO_1378 (O_1378,N_29752,N_29943);
xor UO_1379 (O_1379,N_28874,N_29718);
xnor UO_1380 (O_1380,N_29680,N_29176);
nand UO_1381 (O_1381,N_28943,N_29757);
nand UO_1382 (O_1382,N_29325,N_29750);
xnor UO_1383 (O_1383,N_29177,N_29578);
nand UO_1384 (O_1384,N_28966,N_29695);
nand UO_1385 (O_1385,N_28957,N_29416);
nand UO_1386 (O_1386,N_29079,N_29548);
xnor UO_1387 (O_1387,N_29818,N_29083);
nor UO_1388 (O_1388,N_29225,N_29873);
xor UO_1389 (O_1389,N_28986,N_29387);
nor UO_1390 (O_1390,N_29040,N_29996);
and UO_1391 (O_1391,N_29280,N_29335);
nand UO_1392 (O_1392,N_28908,N_29975);
or UO_1393 (O_1393,N_29973,N_29439);
nand UO_1394 (O_1394,N_29155,N_29401);
nor UO_1395 (O_1395,N_29848,N_29245);
and UO_1396 (O_1396,N_29888,N_29511);
and UO_1397 (O_1397,N_29737,N_29983);
nor UO_1398 (O_1398,N_29099,N_29382);
nor UO_1399 (O_1399,N_29404,N_29942);
nand UO_1400 (O_1400,N_29022,N_29572);
or UO_1401 (O_1401,N_28950,N_29401);
xor UO_1402 (O_1402,N_29215,N_29192);
or UO_1403 (O_1403,N_29592,N_29934);
and UO_1404 (O_1404,N_29378,N_29787);
nor UO_1405 (O_1405,N_29925,N_28953);
nand UO_1406 (O_1406,N_29606,N_29734);
nand UO_1407 (O_1407,N_28967,N_28832);
or UO_1408 (O_1408,N_29903,N_29234);
nor UO_1409 (O_1409,N_29613,N_29774);
or UO_1410 (O_1410,N_28989,N_29313);
xnor UO_1411 (O_1411,N_29509,N_29856);
nor UO_1412 (O_1412,N_29528,N_29898);
and UO_1413 (O_1413,N_29208,N_29346);
and UO_1414 (O_1414,N_28896,N_29058);
and UO_1415 (O_1415,N_29344,N_29644);
nor UO_1416 (O_1416,N_29364,N_28919);
nand UO_1417 (O_1417,N_29989,N_29098);
or UO_1418 (O_1418,N_29004,N_29824);
or UO_1419 (O_1419,N_29972,N_29365);
or UO_1420 (O_1420,N_29595,N_29414);
nor UO_1421 (O_1421,N_29768,N_28897);
or UO_1422 (O_1422,N_28977,N_29597);
xor UO_1423 (O_1423,N_29587,N_28833);
nor UO_1424 (O_1424,N_28916,N_29591);
or UO_1425 (O_1425,N_29828,N_29408);
and UO_1426 (O_1426,N_29762,N_29080);
or UO_1427 (O_1427,N_29882,N_29958);
and UO_1428 (O_1428,N_28857,N_29879);
or UO_1429 (O_1429,N_29347,N_29324);
nor UO_1430 (O_1430,N_28989,N_29024);
nor UO_1431 (O_1431,N_29540,N_29843);
nand UO_1432 (O_1432,N_29967,N_28857);
xor UO_1433 (O_1433,N_29720,N_28839);
xnor UO_1434 (O_1434,N_29840,N_29351);
and UO_1435 (O_1435,N_29217,N_29297);
xor UO_1436 (O_1436,N_29857,N_29320);
or UO_1437 (O_1437,N_29165,N_29736);
nor UO_1438 (O_1438,N_29827,N_29932);
nor UO_1439 (O_1439,N_29443,N_29235);
nor UO_1440 (O_1440,N_29653,N_29368);
or UO_1441 (O_1441,N_29699,N_29727);
nor UO_1442 (O_1442,N_28851,N_29768);
nand UO_1443 (O_1443,N_29133,N_28866);
xor UO_1444 (O_1444,N_29578,N_29588);
or UO_1445 (O_1445,N_29380,N_29458);
and UO_1446 (O_1446,N_29779,N_29887);
nand UO_1447 (O_1447,N_29737,N_29314);
nor UO_1448 (O_1448,N_29400,N_29557);
nor UO_1449 (O_1449,N_29041,N_28809);
nand UO_1450 (O_1450,N_28806,N_28938);
nor UO_1451 (O_1451,N_29103,N_29669);
and UO_1452 (O_1452,N_29805,N_29262);
or UO_1453 (O_1453,N_29180,N_29130);
or UO_1454 (O_1454,N_29971,N_29679);
or UO_1455 (O_1455,N_29595,N_29206);
nand UO_1456 (O_1456,N_29980,N_29278);
and UO_1457 (O_1457,N_29031,N_29938);
nand UO_1458 (O_1458,N_29645,N_29893);
or UO_1459 (O_1459,N_29789,N_29245);
nor UO_1460 (O_1460,N_29598,N_29772);
nor UO_1461 (O_1461,N_29123,N_29227);
and UO_1462 (O_1462,N_29114,N_28938);
nor UO_1463 (O_1463,N_29778,N_29775);
xor UO_1464 (O_1464,N_29588,N_29912);
or UO_1465 (O_1465,N_29139,N_29272);
and UO_1466 (O_1466,N_29319,N_29699);
nand UO_1467 (O_1467,N_29375,N_29361);
nand UO_1468 (O_1468,N_29557,N_29496);
or UO_1469 (O_1469,N_29741,N_28803);
and UO_1470 (O_1470,N_29735,N_29894);
nor UO_1471 (O_1471,N_29008,N_29202);
xnor UO_1472 (O_1472,N_29964,N_29005);
nor UO_1473 (O_1473,N_29757,N_29118);
nor UO_1474 (O_1474,N_29389,N_28875);
nor UO_1475 (O_1475,N_29724,N_29210);
nor UO_1476 (O_1476,N_29492,N_29213);
and UO_1477 (O_1477,N_29881,N_28944);
and UO_1478 (O_1478,N_29733,N_29376);
and UO_1479 (O_1479,N_29398,N_29205);
xnor UO_1480 (O_1480,N_29387,N_28955);
and UO_1481 (O_1481,N_29461,N_29792);
nand UO_1482 (O_1482,N_29742,N_29802);
xnor UO_1483 (O_1483,N_29645,N_29795);
or UO_1484 (O_1484,N_29873,N_29668);
and UO_1485 (O_1485,N_28892,N_28904);
nor UO_1486 (O_1486,N_29942,N_29485);
and UO_1487 (O_1487,N_29555,N_29393);
or UO_1488 (O_1488,N_29419,N_28808);
nand UO_1489 (O_1489,N_29061,N_29363);
or UO_1490 (O_1490,N_29072,N_29393);
and UO_1491 (O_1491,N_29146,N_29579);
xor UO_1492 (O_1492,N_29765,N_29602);
or UO_1493 (O_1493,N_29964,N_29484);
nor UO_1494 (O_1494,N_29101,N_28837);
nand UO_1495 (O_1495,N_28820,N_28826);
xor UO_1496 (O_1496,N_29347,N_28925);
nand UO_1497 (O_1497,N_29149,N_29238);
nor UO_1498 (O_1498,N_29833,N_29661);
and UO_1499 (O_1499,N_29221,N_29274);
xor UO_1500 (O_1500,N_28945,N_29169);
nand UO_1501 (O_1501,N_29888,N_29559);
nand UO_1502 (O_1502,N_28897,N_28872);
or UO_1503 (O_1503,N_29761,N_29132);
xnor UO_1504 (O_1504,N_29652,N_29558);
xor UO_1505 (O_1505,N_29108,N_29179);
nor UO_1506 (O_1506,N_29942,N_29354);
or UO_1507 (O_1507,N_28917,N_29770);
nor UO_1508 (O_1508,N_29438,N_29892);
or UO_1509 (O_1509,N_29774,N_29264);
nand UO_1510 (O_1510,N_29086,N_29160);
xnor UO_1511 (O_1511,N_29689,N_28927);
nand UO_1512 (O_1512,N_29853,N_29375);
and UO_1513 (O_1513,N_29489,N_29696);
xnor UO_1514 (O_1514,N_29682,N_29405);
and UO_1515 (O_1515,N_29800,N_28877);
and UO_1516 (O_1516,N_29693,N_29916);
xor UO_1517 (O_1517,N_29825,N_29596);
and UO_1518 (O_1518,N_28948,N_29043);
nand UO_1519 (O_1519,N_29434,N_29483);
and UO_1520 (O_1520,N_28878,N_29040);
and UO_1521 (O_1521,N_29965,N_29025);
nand UO_1522 (O_1522,N_29280,N_29926);
or UO_1523 (O_1523,N_28930,N_29958);
nand UO_1524 (O_1524,N_29376,N_29300);
nand UO_1525 (O_1525,N_29808,N_29468);
nand UO_1526 (O_1526,N_28973,N_29223);
nand UO_1527 (O_1527,N_29906,N_29358);
xor UO_1528 (O_1528,N_29149,N_29467);
nor UO_1529 (O_1529,N_29050,N_29523);
or UO_1530 (O_1530,N_29696,N_29397);
nand UO_1531 (O_1531,N_29348,N_29082);
or UO_1532 (O_1532,N_29368,N_29888);
nand UO_1533 (O_1533,N_28829,N_29375);
nor UO_1534 (O_1534,N_29490,N_29950);
and UO_1535 (O_1535,N_29413,N_29938);
or UO_1536 (O_1536,N_29731,N_29352);
and UO_1537 (O_1537,N_29306,N_29031);
and UO_1538 (O_1538,N_29499,N_29203);
xor UO_1539 (O_1539,N_29262,N_28806);
or UO_1540 (O_1540,N_29961,N_28929);
or UO_1541 (O_1541,N_29189,N_29426);
xnor UO_1542 (O_1542,N_29368,N_29592);
nor UO_1543 (O_1543,N_29158,N_29867);
nor UO_1544 (O_1544,N_28832,N_28958);
xor UO_1545 (O_1545,N_28954,N_29176);
or UO_1546 (O_1546,N_29010,N_29724);
xor UO_1547 (O_1547,N_29744,N_28836);
xor UO_1548 (O_1548,N_28826,N_29825);
nor UO_1549 (O_1549,N_29267,N_29840);
nand UO_1550 (O_1550,N_29249,N_29873);
nor UO_1551 (O_1551,N_29215,N_29943);
xor UO_1552 (O_1552,N_28998,N_29334);
nand UO_1553 (O_1553,N_29010,N_29422);
or UO_1554 (O_1554,N_28977,N_29654);
and UO_1555 (O_1555,N_29056,N_29571);
nor UO_1556 (O_1556,N_28887,N_29346);
or UO_1557 (O_1557,N_28860,N_29985);
nor UO_1558 (O_1558,N_29776,N_29956);
nand UO_1559 (O_1559,N_29180,N_28857);
nor UO_1560 (O_1560,N_29536,N_29163);
nor UO_1561 (O_1561,N_29295,N_29855);
nand UO_1562 (O_1562,N_29656,N_29581);
and UO_1563 (O_1563,N_29830,N_29429);
or UO_1564 (O_1564,N_28995,N_29844);
or UO_1565 (O_1565,N_29253,N_29102);
and UO_1566 (O_1566,N_29045,N_29597);
nand UO_1567 (O_1567,N_28836,N_28841);
and UO_1568 (O_1568,N_29270,N_29695);
or UO_1569 (O_1569,N_29708,N_29114);
nand UO_1570 (O_1570,N_29959,N_29511);
or UO_1571 (O_1571,N_29057,N_29013);
nand UO_1572 (O_1572,N_29712,N_29583);
nor UO_1573 (O_1573,N_29022,N_29357);
and UO_1574 (O_1574,N_28911,N_29623);
nand UO_1575 (O_1575,N_29113,N_29370);
nand UO_1576 (O_1576,N_29227,N_28899);
nand UO_1577 (O_1577,N_29307,N_29596);
nor UO_1578 (O_1578,N_29926,N_29163);
xor UO_1579 (O_1579,N_28998,N_29096);
nor UO_1580 (O_1580,N_29442,N_29417);
or UO_1581 (O_1581,N_29373,N_28898);
nor UO_1582 (O_1582,N_29732,N_29100);
or UO_1583 (O_1583,N_29266,N_29358);
nor UO_1584 (O_1584,N_29545,N_29609);
nand UO_1585 (O_1585,N_28912,N_29563);
nor UO_1586 (O_1586,N_28866,N_28963);
nand UO_1587 (O_1587,N_29844,N_29202);
and UO_1588 (O_1588,N_29384,N_29409);
nand UO_1589 (O_1589,N_29572,N_29021);
or UO_1590 (O_1590,N_29328,N_28805);
or UO_1591 (O_1591,N_29907,N_29024);
nand UO_1592 (O_1592,N_29179,N_28925);
xor UO_1593 (O_1593,N_29634,N_28905);
nor UO_1594 (O_1594,N_28991,N_29299);
nor UO_1595 (O_1595,N_29034,N_29125);
or UO_1596 (O_1596,N_29096,N_29909);
nor UO_1597 (O_1597,N_28980,N_29989);
xor UO_1598 (O_1598,N_29605,N_29870);
nand UO_1599 (O_1599,N_29391,N_29114);
or UO_1600 (O_1600,N_28873,N_28897);
xnor UO_1601 (O_1601,N_29489,N_29334);
or UO_1602 (O_1602,N_29073,N_28868);
xor UO_1603 (O_1603,N_29507,N_29017);
nor UO_1604 (O_1604,N_29770,N_28986);
or UO_1605 (O_1605,N_29193,N_29963);
and UO_1606 (O_1606,N_28806,N_29561);
nor UO_1607 (O_1607,N_28942,N_29791);
nand UO_1608 (O_1608,N_28952,N_29683);
nand UO_1609 (O_1609,N_29967,N_29012);
nor UO_1610 (O_1610,N_29200,N_29261);
nand UO_1611 (O_1611,N_28903,N_28875);
nor UO_1612 (O_1612,N_28960,N_29258);
nor UO_1613 (O_1613,N_29568,N_29512);
or UO_1614 (O_1614,N_29209,N_29552);
xnor UO_1615 (O_1615,N_29251,N_29150);
and UO_1616 (O_1616,N_29339,N_29898);
xnor UO_1617 (O_1617,N_29852,N_29123);
and UO_1618 (O_1618,N_29307,N_29677);
nor UO_1619 (O_1619,N_29096,N_29879);
or UO_1620 (O_1620,N_29324,N_29426);
xor UO_1621 (O_1621,N_29558,N_29112);
and UO_1622 (O_1622,N_29926,N_29780);
or UO_1623 (O_1623,N_29060,N_29716);
xnor UO_1624 (O_1624,N_29595,N_28870);
and UO_1625 (O_1625,N_29455,N_29497);
and UO_1626 (O_1626,N_29061,N_29068);
and UO_1627 (O_1627,N_29245,N_28813);
nor UO_1628 (O_1628,N_29419,N_29022);
nand UO_1629 (O_1629,N_28975,N_29850);
nand UO_1630 (O_1630,N_29058,N_29147);
xnor UO_1631 (O_1631,N_29871,N_29050);
or UO_1632 (O_1632,N_29515,N_29592);
and UO_1633 (O_1633,N_29095,N_29451);
xnor UO_1634 (O_1634,N_29479,N_29159);
or UO_1635 (O_1635,N_29580,N_29235);
xnor UO_1636 (O_1636,N_29692,N_29358);
xnor UO_1637 (O_1637,N_29302,N_29725);
and UO_1638 (O_1638,N_29036,N_28882);
nand UO_1639 (O_1639,N_29097,N_28863);
and UO_1640 (O_1640,N_29024,N_29643);
nor UO_1641 (O_1641,N_29973,N_29770);
and UO_1642 (O_1642,N_29703,N_29863);
xor UO_1643 (O_1643,N_29274,N_29601);
nor UO_1644 (O_1644,N_29225,N_29597);
or UO_1645 (O_1645,N_29345,N_29648);
or UO_1646 (O_1646,N_29431,N_29988);
nor UO_1647 (O_1647,N_29948,N_28965);
nand UO_1648 (O_1648,N_28832,N_29383);
nand UO_1649 (O_1649,N_28820,N_29524);
xor UO_1650 (O_1650,N_29200,N_29912);
nand UO_1651 (O_1651,N_28990,N_29664);
and UO_1652 (O_1652,N_29286,N_29310);
or UO_1653 (O_1653,N_29743,N_29869);
nand UO_1654 (O_1654,N_29219,N_28800);
xor UO_1655 (O_1655,N_29456,N_29305);
xor UO_1656 (O_1656,N_28879,N_29476);
or UO_1657 (O_1657,N_29089,N_29889);
nand UO_1658 (O_1658,N_29242,N_28852);
nor UO_1659 (O_1659,N_29391,N_29503);
or UO_1660 (O_1660,N_29313,N_29198);
nand UO_1661 (O_1661,N_29273,N_28945);
or UO_1662 (O_1662,N_29082,N_29366);
nand UO_1663 (O_1663,N_29029,N_29121);
and UO_1664 (O_1664,N_29065,N_28839);
or UO_1665 (O_1665,N_28892,N_28861);
or UO_1666 (O_1666,N_29124,N_28948);
nand UO_1667 (O_1667,N_29985,N_29607);
and UO_1668 (O_1668,N_29615,N_28832);
nand UO_1669 (O_1669,N_29954,N_29309);
xnor UO_1670 (O_1670,N_29553,N_29732);
or UO_1671 (O_1671,N_29049,N_29131);
and UO_1672 (O_1672,N_29187,N_29169);
nor UO_1673 (O_1673,N_29857,N_29191);
nand UO_1674 (O_1674,N_29924,N_29725);
and UO_1675 (O_1675,N_29925,N_29010);
nor UO_1676 (O_1676,N_29445,N_29960);
nand UO_1677 (O_1677,N_29930,N_29897);
xor UO_1678 (O_1678,N_29562,N_29586);
nor UO_1679 (O_1679,N_29946,N_29652);
and UO_1680 (O_1680,N_29652,N_29697);
or UO_1681 (O_1681,N_29847,N_29446);
nor UO_1682 (O_1682,N_29816,N_29448);
nor UO_1683 (O_1683,N_29463,N_28938);
and UO_1684 (O_1684,N_29467,N_29876);
xnor UO_1685 (O_1685,N_29502,N_29005);
or UO_1686 (O_1686,N_28900,N_28930);
nor UO_1687 (O_1687,N_29793,N_28803);
and UO_1688 (O_1688,N_28882,N_29859);
nand UO_1689 (O_1689,N_29117,N_29985);
xnor UO_1690 (O_1690,N_29418,N_29813);
xor UO_1691 (O_1691,N_28927,N_29877);
nand UO_1692 (O_1692,N_29677,N_29854);
and UO_1693 (O_1693,N_29826,N_29595);
and UO_1694 (O_1694,N_29643,N_29228);
xnor UO_1695 (O_1695,N_29706,N_29794);
or UO_1696 (O_1696,N_29707,N_29927);
nand UO_1697 (O_1697,N_29673,N_29457);
nand UO_1698 (O_1698,N_29142,N_29382);
nor UO_1699 (O_1699,N_29618,N_29285);
or UO_1700 (O_1700,N_29888,N_29619);
nand UO_1701 (O_1701,N_29069,N_29886);
nand UO_1702 (O_1702,N_29388,N_29963);
xnor UO_1703 (O_1703,N_29287,N_29309);
nand UO_1704 (O_1704,N_29885,N_29460);
nand UO_1705 (O_1705,N_29236,N_28814);
nand UO_1706 (O_1706,N_28853,N_28924);
or UO_1707 (O_1707,N_29293,N_29624);
and UO_1708 (O_1708,N_29064,N_28951);
or UO_1709 (O_1709,N_28970,N_29928);
and UO_1710 (O_1710,N_29418,N_29137);
nor UO_1711 (O_1711,N_28946,N_29803);
xor UO_1712 (O_1712,N_29501,N_29348);
nand UO_1713 (O_1713,N_29759,N_29490);
xor UO_1714 (O_1714,N_29246,N_28827);
or UO_1715 (O_1715,N_29939,N_29921);
nand UO_1716 (O_1716,N_29201,N_29482);
and UO_1717 (O_1717,N_29115,N_29939);
and UO_1718 (O_1718,N_29516,N_29219);
nor UO_1719 (O_1719,N_29296,N_29763);
nand UO_1720 (O_1720,N_28944,N_29131);
and UO_1721 (O_1721,N_29698,N_29747);
and UO_1722 (O_1722,N_29016,N_28900);
or UO_1723 (O_1723,N_29420,N_29686);
or UO_1724 (O_1724,N_29524,N_29646);
and UO_1725 (O_1725,N_28810,N_29877);
and UO_1726 (O_1726,N_29701,N_29476);
nand UO_1727 (O_1727,N_29750,N_29435);
xor UO_1728 (O_1728,N_29425,N_29790);
nor UO_1729 (O_1729,N_28840,N_29394);
nor UO_1730 (O_1730,N_29205,N_29103);
nand UO_1731 (O_1731,N_28951,N_29356);
nand UO_1732 (O_1732,N_29432,N_29833);
nand UO_1733 (O_1733,N_29925,N_29884);
and UO_1734 (O_1734,N_28959,N_29525);
xnor UO_1735 (O_1735,N_29534,N_28896);
and UO_1736 (O_1736,N_28957,N_29721);
xor UO_1737 (O_1737,N_29016,N_29353);
and UO_1738 (O_1738,N_29461,N_29879);
and UO_1739 (O_1739,N_29337,N_28933);
and UO_1740 (O_1740,N_29565,N_29578);
nand UO_1741 (O_1741,N_29252,N_28940);
nand UO_1742 (O_1742,N_28889,N_29195);
and UO_1743 (O_1743,N_29115,N_29255);
or UO_1744 (O_1744,N_29563,N_29674);
nand UO_1745 (O_1745,N_29429,N_29740);
nor UO_1746 (O_1746,N_28858,N_28998);
or UO_1747 (O_1747,N_28938,N_29076);
and UO_1748 (O_1748,N_29416,N_29436);
nand UO_1749 (O_1749,N_29260,N_29085);
nor UO_1750 (O_1750,N_29392,N_29087);
nand UO_1751 (O_1751,N_29374,N_29616);
xor UO_1752 (O_1752,N_28938,N_29207);
xor UO_1753 (O_1753,N_29519,N_29187);
xor UO_1754 (O_1754,N_29653,N_29947);
or UO_1755 (O_1755,N_29215,N_29963);
nand UO_1756 (O_1756,N_29906,N_29287);
or UO_1757 (O_1757,N_29004,N_29423);
nand UO_1758 (O_1758,N_29815,N_29059);
or UO_1759 (O_1759,N_29984,N_28893);
xor UO_1760 (O_1760,N_29482,N_29229);
or UO_1761 (O_1761,N_29420,N_29028);
and UO_1762 (O_1762,N_29460,N_29484);
nand UO_1763 (O_1763,N_28834,N_29157);
nand UO_1764 (O_1764,N_29460,N_29184);
nor UO_1765 (O_1765,N_29556,N_29443);
or UO_1766 (O_1766,N_29141,N_29271);
nor UO_1767 (O_1767,N_29300,N_29641);
nand UO_1768 (O_1768,N_29432,N_29108);
nand UO_1769 (O_1769,N_29763,N_29328);
nor UO_1770 (O_1770,N_29203,N_29564);
or UO_1771 (O_1771,N_29956,N_29491);
or UO_1772 (O_1772,N_29753,N_29454);
and UO_1773 (O_1773,N_28888,N_29418);
nor UO_1774 (O_1774,N_28956,N_29397);
nor UO_1775 (O_1775,N_29876,N_29394);
or UO_1776 (O_1776,N_29012,N_29822);
and UO_1777 (O_1777,N_29298,N_29822);
or UO_1778 (O_1778,N_28988,N_29474);
or UO_1779 (O_1779,N_29353,N_29637);
xnor UO_1780 (O_1780,N_29284,N_29232);
nor UO_1781 (O_1781,N_29962,N_29511);
nor UO_1782 (O_1782,N_29094,N_29484);
nor UO_1783 (O_1783,N_29281,N_29351);
or UO_1784 (O_1784,N_28856,N_29970);
or UO_1785 (O_1785,N_29376,N_29437);
xor UO_1786 (O_1786,N_29332,N_28983);
or UO_1787 (O_1787,N_29121,N_29466);
and UO_1788 (O_1788,N_29441,N_29566);
nor UO_1789 (O_1789,N_29215,N_29855);
and UO_1790 (O_1790,N_28928,N_29590);
or UO_1791 (O_1791,N_29795,N_29780);
and UO_1792 (O_1792,N_29130,N_29527);
and UO_1793 (O_1793,N_29219,N_29758);
nand UO_1794 (O_1794,N_29733,N_29021);
and UO_1795 (O_1795,N_28941,N_29789);
nand UO_1796 (O_1796,N_29507,N_29173);
nor UO_1797 (O_1797,N_28919,N_29339);
nand UO_1798 (O_1798,N_29078,N_29180);
nor UO_1799 (O_1799,N_29470,N_29476);
or UO_1800 (O_1800,N_29083,N_29830);
xor UO_1801 (O_1801,N_29338,N_29892);
nor UO_1802 (O_1802,N_29663,N_28908);
nor UO_1803 (O_1803,N_29589,N_29796);
nand UO_1804 (O_1804,N_29553,N_29126);
or UO_1805 (O_1805,N_28817,N_29402);
and UO_1806 (O_1806,N_29329,N_29508);
or UO_1807 (O_1807,N_29984,N_29493);
nand UO_1808 (O_1808,N_29905,N_29992);
nand UO_1809 (O_1809,N_29684,N_29035);
nor UO_1810 (O_1810,N_29194,N_29182);
or UO_1811 (O_1811,N_29182,N_29474);
or UO_1812 (O_1812,N_29037,N_29824);
or UO_1813 (O_1813,N_29177,N_28861);
nand UO_1814 (O_1814,N_29881,N_29903);
nor UO_1815 (O_1815,N_29914,N_28823);
nand UO_1816 (O_1816,N_29821,N_28988);
or UO_1817 (O_1817,N_29376,N_29819);
or UO_1818 (O_1818,N_29704,N_28820);
nand UO_1819 (O_1819,N_29936,N_29142);
nand UO_1820 (O_1820,N_29331,N_28852);
nor UO_1821 (O_1821,N_28927,N_29521);
or UO_1822 (O_1822,N_28946,N_28861);
xor UO_1823 (O_1823,N_29984,N_29869);
and UO_1824 (O_1824,N_29972,N_28924);
and UO_1825 (O_1825,N_29461,N_29102);
or UO_1826 (O_1826,N_29496,N_29205);
nand UO_1827 (O_1827,N_29417,N_29533);
nand UO_1828 (O_1828,N_29740,N_29200);
and UO_1829 (O_1829,N_29534,N_29999);
and UO_1830 (O_1830,N_29403,N_29780);
or UO_1831 (O_1831,N_29213,N_29420);
xnor UO_1832 (O_1832,N_29557,N_29659);
or UO_1833 (O_1833,N_29622,N_29858);
xor UO_1834 (O_1834,N_29482,N_29190);
nor UO_1835 (O_1835,N_29618,N_29388);
nand UO_1836 (O_1836,N_29027,N_29970);
nand UO_1837 (O_1837,N_29599,N_29049);
and UO_1838 (O_1838,N_29279,N_29458);
nor UO_1839 (O_1839,N_29287,N_29889);
nand UO_1840 (O_1840,N_29262,N_29570);
nor UO_1841 (O_1841,N_29479,N_28943);
nor UO_1842 (O_1842,N_29386,N_28837);
nor UO_1843 (O_1843,N_29910,N_29707);
or UO_1844 (O_1844,N_29462,N_28910);
xor UO_1845 (O_1845,N_29962,N_29243);
or UO_1846 (O_1846,N_29080,N_29814);
nor UO_1847 (O_1847,N_29963,N_28867);
nor UO_1848 (O_1848,N_29069,N_29511);
or UO_1849 (O_1849,N_29100,N_29992);
and UO_1850 (O_1850,N_29066,N_29097);
xnor UO_1851 (O_1851,N_28936,N_28926);
and UO_1852 (O_1852,N_29110,N_29700);
or UO_1853 (O_1853,N_29931,N_29220);
nor UO_1854 (O_1854,N_28902,N_28952);
nand UO_1855 (O_1855,N_29809,N_28870);
xnor UO_1856 (O_1856,N_29926,N_29400);
nand UO_1857 (O_1857,N_29238,N_29019);
nor UO_1858 (O_1858,N_29758,N_29186);
or UO_1859 (O_1859,N_29772,N_29931);
xnor UO_1860 (O_1860,N_29624,N_29435);
nor UO_1861 (O_1861,N_29922,N_28908);
and UO_1862 (O_1862,N_29329,N_29793);
xor UO_1863 (O_1863,N_29568,N_29183);
nor UO_1864 (O_1864,N_29060,N_29179);
or UO_1865 (O_1865,N_29880,N_29841);
nand UO_1866 (O_1866,N_29236,N_29798);
and UO_1867 (O_1867,N_28825,N_29676);
or UO_1868 (O_1868,N_29720,N_28825);
xor UO_1869 (O_1869,N_29017,N_29894);
and UO_1870 (O_1870,N_29566,N_29903);
nor UO_1871 (O_1871,N_28963,N_29211);
nand UO_1872 (O_1872,N_29215,N_29264);
nand UO_1873 (O_1873,N_28960,N_29406);
nor UO_1874 (O_1874,N_29676,N_29735);
nor UO_1875 (O_1875,N_29459,N_29436);
and UO_1876 (O_1876,N_29821,N_29785);
and UO_1877 (O_1877,N_29919,N_28878);
xor UO_1878 (O_1878,N_28960,N_29975);
nor UO_1879 (O_1879,N_29509,N_29705);
or UO_1880 (O_1880,N_29963,N_29452);
or UO_1881 (O_1881,N_29877,N_29874);
or UO_1882 (O_1882,N_28884,N_29072);
and UO_1883 (O_1883,N_29639,N_29770);
or UO_1884 (O_1884,N_29135,N_29407);
and UO_1885 (O_1885,N_29019,N_28855);
or UO_1886 (O_1886,N_28851,N_28887);
nor UO_1887 (O_1887,N_29729,N_28814);
nor UO_1888 (O_1888,N_29745,N_29200);
xor UO_1889 (O_1889,N_29278,N_29482);
or UO_1890 (O_1890,N_29192,N_29677);
or UO_1891 (O_1891,N_28857,N_29774);
and UO_1892 (O_1892,N_29666,N_29504);
and UO_1893 (O_1893,N_29671,N_29360);
and UO_1894 (O_1894,N_29640,N_29720);
and UO_1895 (O_1895,N_28884,N_29009);
xor UO_1896 (O_1896,N_28997,N_28993);
nand UO_1897 (O_1897,N_29089,N_29090);
nand UO_1898 (O_1898,N_29133,N_29000);
xnor UO_1899 (O_1899,N_29406,N_29541);
or UO_1900 (O_1900,N_29902,N_29374);
nor UO_1901 (O_1901,N_29735,N_29125);
and UO_1902 (O_1902,N_29793,N_29552);
or UO_1903 (O_1903,N_29082,N_29744);
nand UO_1904 (O_1904,N_29541,N_29566);
and UO_1905 (O_1905,N_29079,N_29701);
xnor UO_1906 (O_1906,N_29537,N_29249);
or UO_1907 (O_1907,N_29564,N_28990);
xor UO_1908 (O_1908,N_29096,N_29979);
nand UO_1909 (O_1909,N_29943,N_29396);
nor UO_1910 (O_1910,N_29202,N_29127);
and UO_1911 (O_1911,N_28968,N_29725);
nand UO_1912 (O_1912,N_29375,N_29724);
and UO_1913 (O_1913,N_29177,N_29266);
nor UO_1914 (O_1914,N_29024,N_29494);
nand UO_1915 (O_1915,N_29236,N_28975);
nand UO_1916 (O_1916,N_29307,N_29725);
and UO_1917 (O_1917,N_29218,N_29780);
nor UO_1918 (O_1918,N_29501,N_29533);
nand UO_1919 (O_1919,N_29988,N_29818);
xor UO_1920 (O_1920,N_29234,N_29609);
nor UO_1921 (O_1921,N_29413,N_29464);
or UO_1922 (O_1922,N_29963,N_29817);
nand UO_1923 (O_1923,N_29623,N_29097);
xnor UO_1924 (O_1924,N_29094,N_29505);
nor UO_1925 (O_1925,N_29178,N_29138);
nand UO_1926 (O_1926,N_29303,N_29030);
or UO_1927 (O_1927,N_29888,N_29066);
nor UO_1928 (O_1928,N_29345,N_29482);
xnor UO_1929 (O_1929,N_29702,N_29639);
nand UO_1930 (O_1930,N_29275,N_29268);
nand UO_1931 (O_1931,N_29804,N_29220);
or UO_1932 (O_1932,N_28961,N_29024);
or UO_1933 (O_1933,N_29707,N_29270);
or UO_1934 (O_1934,N_29234,N_29781);
nor UO_1935 (O_1935,N_29265,N_29100);
or UO_1936 (O_1936,N_29542,N_29615);
and UO_1937 (O_1937,N_29962,N_28883);
or UO_1938 (O_1938,N_29944,N_29594);
nor UO_1939 (O_1939,N_29633,N_29252);
xor UO_1940 (O_1940,N_29230,N_29219);
nand UO_1941 (O_1941,N_29676,N_29736);
nor UO_1942 (O_1942,N_29480,N_29902);
nor UO_1943 (O_1943,N_29820,N_29187);
nor UO_1944 (O_1944,N_29883,N_29874);
or UO_1945 (O_1945,N_28849,N_29130);
nor UO_1946 (O_1946,N_29966,N_29427);
nor UO_1947 (O_1947,N_29815,N_29643);
nor UO_1948 (O_1948,N_29333,N_29292);
nand UO_1949 (O_1949,N_29473,N_28883);
xnor UO_1950 (O_1950,N_28868,N_29013);
or UO_1951 (O_1951,N_29726,N_29161);
and UO_1952 (O_1952,N_29322,N_29361);
nor UO_1953 (O_1953,N_29361,N_29703);
or UO_1954 (O_1954,N_29722,N_29824);
nand UO_1955 (O_1955,N_29833,N_29503);
nand UO_1956 (O_1956,N_29569,N_29446);
nand UO_1957 (O_1957,N_29626,N_28867);
nor UO_1958 (O_1958,N_29988,N_29220);
or UO_1959 (O_1959,N_29806,N_29462);
or UO_1960 (O_1960,N_29386,N_29279);
xor UO_1961 (O_1961,N_29290,N_29438);
or UO_1962 (O_1962,N_29202,N_29485);
nand UO_1963 (O_1963,N_28967,N_29238);
or UO_1964 (O_1964,N_29405,N_29448);
nand UO_1965 (O_1965,N_29878,N_29404);
and UO_1966 (O_1966,N_29454,N_29574);
nor UO_1967 (O_1967,N_28994,N_29734);
nand UO_1968 (O_1968,N_28999,N_28908);
nor UO_1969 (O_1969,N_29840,N_29213);
and UO_1970 (O_1970,N_29712,N_29693);
or UO_1971 (O_1971,N_29411,N_28832);
nor UO_1972 (O_1972,N_29649,N_29476);
or UO_1973 (O_1973,N_29385,N_29663);
nand UO_1974 (O_1974,N_28941,N_28870);
and UO_1975 (O_1975,N_29571,N_29575);
and UO_1976 (O_1976,N_29112,N_28817);
xor UO_1977 (O_1977,N_29087,N_29580);
nand UO_1978 (O_1978,N_29033,N_29619);
and UO_1979 (O_1979,N_29770,N_29160);
and UO_1980 (O_1980,N_29026,N_28923);
or UO_1981 (O_1981,N_29105,N_29563);
nor UO_1982 (O_1982,N_28850,N_28973);
xnor UO_1983 (O_1983,N_29200,N_28916);
and UO_1984 (O_1984,N_29090,N_29103);
and UO_1985 (O_1985,N_29288,N_29228);
and UO_1986 (O_1986,N_29044,N_29074);
nand UO_1987 (O_1987,N_29892,N_29828);
or UO_1988 (O_1988,N_28923,N_28992);
and UO_1989 (O_1989,N_29199,N_29722);
and UO_1990 (O_1990,N_29155,N_29154);
nor UO_1991 (O_1991,N_29711,N_29227);
nor UO_1992 (O_1992,N_28818,N_29819);
nor UO_1993 (O_1993,N_28924,N_28890);
nand UO_1994 (O_1994,N_29292,N_29099);
nor UO_1995 (O_1995,N_28990,N_29078);
nand UO_1996 (O_1996,N_29934,N_29166);
xor UO_1997 (O_1997,N_29136,N_29788);
nor UO_1998 (O_1998,N_29550,N_29850);
xnor UO_1999 (O_1999,N_29546,N_29288);
nand UO_2000 (O_2000,N_28923,N_28891);
and UO_2001 (O_2001,N_29369,N_29284);
nor UO_2002 (O_2002,N_29607,N_29935);
nor UO_2003 (O_2003,N_29451,N_29744);
or UO_2004 (O_2004,N_29195,N_28974);
nor UO_2005 (O_2005,N_29173,N_29954);
or UO_2006 (O_2006,N_29521,N_29575);
nor UO_2007 (O_2007,N_29268,N_28999);
nand UO_2008 (O_2008,N_29909,N_29546);
and UO_2009 (O_2009,N_29650,N_29172);
nor UO_2010 (O_2010,N_28902,N_29586);
xnor UO_2011 (O_2011,N_29589,N_29935);
or UO_2012 (O_2012,N_29038,N_29329);
nand UO_2013 (O_2013,N_29778,N_29218);
nand UO_2014 (O_2014,N_29716,N_29600);
nor UO_2015 (O_2015,N_29122,N_29135);
and UO_2016 (O_2016,N_28975,N_29124);
and UO_2017 (O_2017,N_28929,N_28862);
or UO_2018 (O_2018,N_29620,N_29228);
and UO_2019 (O_2019,N_28937,N_29417);
or UO_2020 (O_2020,N_29307,N_28903);
or UO_2021 (O_2021,N_28808,N_29977);
nor UO_2022 (O_2022,N_29535,N_29998);
or UO_2023 (O_2023,N_29909,N_29298);
or UO_2024 (O_2024,N_29416,N_29840);
nand UO_2025 (O_2025,N_29493,N_29474);
or UO_2026 (O_2026,N_29803,N_29777);
nor UO_2027 (O_2027,N_29457,N_29002);
xnor UO_2028 (O_2028,N_29038,N_28938);
or UO_2029 (O_2029,N_29861,N_29352);
and UO_2030 (O_2030,N_29138,N_29248);
and UO_2031 (O_2031,N_29975,N_29738);
or UO_2032 (O_2032,N_29600,N_29427);
xnor UO_2033 (O_2033,N_29864,N_29965);
or UO_2034 (O_2034,N_29414,N_29979);
xnor UO_2035 (O_2035,N_28958,N_28985);
or UO_2036 (O_2036,N_29739,N_29169);
and UO_2037 (O_2037,N_29186,N_29148);
nand UO_2038 (O_2038,N_29595,N_29538);
nor UO_2039 (O_2039,N_29911,N_29704);
xor UO_2040 (O_2040,N_29835,N_29048);
nand UO_2041 (O_2041,N_29799,N_29006);
and UO_2042 (O_2042,N_29381,N_29537);
and UO_2043 (O_2043,N_29453,N_29652);
or UO_2044 (O_2044,N_29702,N_29787);
xnor UO_2045 (O_2045,N_29243,N_28847);
nor UO_2046 (O_2046,N_29391,N_28994);
nor UO_2047 (O_2047,N_29518,N_29699);
nand UO_2048 (O_2048,N_29722,N_29761);
nor UO_2049 (O_2049,N_29317,N_29413);
and UO_2050 (O_2050,N_29612,N_29132);
and UO_2051 (O_2051,N_28943,N_29288);
and UO_2052 (O_2052,N_29797,N_29394);
and UO_2053 (O_2053,N_29087,N_29142);
or UO_2054 (O_2054,N_29433,N_29008);
xnor UO_2055 (O_2055,N_29782,N_28826);
xor UO_2056 (O_2056,N_29787,N_29078);
and UO_2057 (O_2057,N_29275,N_29879);
xor UO_2058 (O_2058,N_29558,N_29004);
xor UO_2059 (O_2059,N_29985,N_29917);
or UO_2060 (O_2060,N_29733,N_28978);
and UO_2061 (O_2061,N_29004,N_29537);
nand UO_2062 (O_2062,N_29968,N_29883);
or UO_2063 (O_2063,N_29999,N_28992);
nand UO_2064 (O_2064,N_29952,N_28808);
and UO_2065 (O_2065,N_29230,N_29813);
and UO_2066 (O_2066,N_29405,N_28817);
or UO_2067 (O_2067,N_29211,N_29908);
xor UO_2068 (O_2068,N_29882,N_29826);
nand UO_2069 (O_2069,N_28844,N_29036);
nand UO_2070 (O_2070,N_29415,N_29517);
and UO_2071 (O_2071,N_29178,N_29421);
nor UO_2072 (O_2072,N_29691,N_28910);
or UO_2073 (O_2073,N_28935,N_29106);
xor UO_2074 (O_2074,N_29797,N_28923);
or UO_2075 (O_2075,N_29981,N_29447);
xnor UO_2076 (O_2076,N_28820,N_29360);
xor UO_2077 (O_2077,N_29737,N_29400);
nor UO_2078 (O_2078,N_29003,N_29073);
or UO_2079 (O_2079,N_29752,N_29857);
xor UO_2080 (O_2080,N_29919,N_29773);
or UO_2081 (O_2081,N_29122,N_29356);
nor UO_2082 (O_2082,N_29074,N_29173);
nand UO_2083 (O_2083,N_28974,N_28975);
and UO_2084 (O_2084,N_29003,N_29474);
nor UO_2085 (O_2085,N_29000,N_29628);
or UO_2086 (O_2086,N_29051,N_29584);
or UO_2087 (O_2087,N_29080,N_28808);
and UO_2088 (O_2088,N_29184,N_28973);
and UO_2089 (O_2089,N_29685,N_29937);
nor UO_2090 (O_2090,N_29087,N_29064);
xnor UO_2091 (O_2091,N_29062,N_29116);
xnor UO_2092 (O_2092,N_28950,N_29481);
nand UO_2093 (O_2093,N_29926,N_29308);
or UO_2094 (O_2094,N_28906,N_28926);
and UO_2095 (O_2095,N_29903,N_29865);
nand UO_2096 (O_2096,N_28905,N_29724);
and UO_2097 (O_2097,N_29495,N_29213);
nand UO_2098 (O_2098,N_29945,N_29469);
and UO_2099 (O_2099,N_29378,N_29306);
or UO_2100 (O_2100,N_29628,N_29304);
or UO_2101 (O_2101,N_29968,N_29203);
xor UO_2102 (O_2102,N_29113,N_29116);
xor UO_2103 (O_2103,N_28988,N_29239);
nor UO_2104 (O_2104,N_29470,N_29142);
nand UO_2105 (O_2105,N_28853,N_29373);
nand UO_2106 (O_2106,N_29306,N_29241);
or UO_2107 (O_2107,N_29770,N_28890);
and UO_2108 (O_2108,N_29723,N_29474);
nor UO_2109 (O_2109,N_29087,N_29518);
and UO_2110 (O_2110,N_29863,N_28895);
xor UO_2111 (O_2111,N_29388,N_28945);
nor UO_2112 (O_2112,N_29644,N_29835);
nor UO_2113 (O_2113,N_29032,N_28952);
and UO_2114 (O_2114,N_29507,N_29876);
nand UO_2115 (O_2115,N_29019,N_29817);
or UO_2116 (O_2116,N_29278,N_28963);
nand UO_2117 (O_2117,N_29593,N_29780);
or UO_2118 (O_2118,N_29390,N_29429);
nor UO_2119 (O_2119,N_29750,N_29976);
xor UO_2120 (O_2120,N_29387,N_28816);
nand UO_2121 (O_2121,N_28934,N_29135);
xor UO_2122 (O_2122,N_29361,N_29419);
nand UO_2123 (O_2123,N_29583,N_29811);
or UO_2124 (O_2124,N_29943,N_29235);
or UO_2125 (O_2125,N_28923,N_29754);
nand UO_2126 (O_2126,N_29080,N_29043);
or UO_2127 (O_2127,N_29854,N_28866);
or UO_2128 (O_2128,N_28991,N_29755);
nand UO_2129 (O_2129,N_29741,N_29190);
nor UO_2130 (O_2130,N_28834,N_29604);
and UO_2131 (O_2131,N_29420,N_29421);
xor UO_2132 (O_2132,N_29589,N_29465);
nand UO_2133 (O_2133,N_29913,N_29642);
nor UO_2134 (O_2134,N_29723,N_29294);
xor UO_2135 (O_2135,N_29765,N_29801);
xnor UO_2136 (O_2136,N_29731,N_29412);
and UO_2137 (O_2137,N_29693,N_29009);
or UO_2138 (O_2138,N_29669,N_29851);
nand UO_2139 (O_2139,N_29332,N_29735);
and UO_2140 (O_2140,N_28932,N_29774);
xor UO_2141 (O_2141,N_29031,N_29275);
and UO_2142 (O_2142,N_29387,N_29505);
or UO_2143 (O_2143,N_29658,N_28874);
xor UO_2144 (O_2144,N_29490,N_29713);
nand UO_2145 (O_2145,N_28858,N_29737);
and UO_2146 (O_2146,N_29690,N_29366);
nor UO_2147 (O_2147,N_29312,N_29545);
and UO_2148 (O_2148,N_28910,N_29090);
xnor UO_2149 (O_2149,N_29673,N_28866);
xor UO_2150 (O_2150,N_29699,N_29032);
or UO_2151 (O_2151,N_29846,N_29970);
nor UO_2152 (O_2152,N_29420,N_29754);
nand UO_2153 (O_2153,N_28864,N_29611);
xor UO_2154 (O_2154,N_29235,N_29051);
nor UO_2155 (O_2155,N_28867,N_29789);
nand UO_2156 (O_2156,N_29180,N_29557);
nand UO_2157 (O_2157,N_29103,N_28897);
xor UO_2158 (O_2158,N_29362,N_29086);
nor UO_2159 (O_2159,N_29092,N_28867);
nand UO_2160 (O_2160,N_29780,N_29577);
or UO_2161 (O_2161,N_29128,N_29272);
xnor UO_2162 (O_2162,N_28898,N_29459);
or UO_2163 (O_2163,N_29605,N_29900);
and UO_2164 (O_2164,N_28843,N_29641);
nor UO_2165 (O_2165,N_29490,N_29636);
and UO_2166 (O_2166,N_29259,N_29527);
or UO_2167 (O_2167,N_29229,N_28962);
or UO_2168 (O_2168,N_29721,N_29808);
nand UO_2169 (O_2169,N_29594,N_29566);
or UO_2170 (O_2170,N_29217,N_29456);
nand UO_2171 (O_2171,N_29571,N_29009);
nand UO_2172 (O_2172,N_28893,N_29658);
and UO_2173 (O_2173,N_29353,N_28848);
nor UO_2174 (O_2174,N_29805,N_29151);
nand UO_2175 (O_2175,N_29579,N_29779);
nor UO_2176 (O_2176,N_29053,N_29324);
nand UO_2177 (O_2177,N_29495,N_29233);
or UO_2178 (O_2178,N_29178,N_29062);
and UO_2179 (O_2179,N_29686,N_29540);
and UO_2180 (O_2180,N_29181,N_29364);
nand UO_2181 (O_2181,N_29510,N_29651);
or UO_2182 (O_2182,N_29905,N_29966);
and UO_2183 (O_2183,N_29425,N_29738);
xor UO_2184 (O_2184,N_29684,N_28952);
nor UO_2185 (O_2185,N_29766,N_29067);
or UO_2186 (O_2186,N_29553,N_29243);
or UO_2187 (O_2187,N_28978,N_29189);
nand UO_2188 (O_2188,N_29106,N_29163);
nand UO_2189 (O_2189,N_29846,N_28840);
or UO_2190 (O_2190,N_29242,N_29951);
nor UO_2191 (O_2191,N_29758,N_29476);
nand UO_2192 (O_2192,N_28901,N_29168);
xor UO_2193 (O_2193,N_29250,N_29203);
or UO_2194 (O_2194,N_29829,N_28956);
or UO_2195 (O_2195,N_29474,N_28946);
xnor UO_2196 (O_2196,N_29552,N_28858);
nor UO_2197 (O_2197,N_29542,N_29484);
nor UO_2198 (O_2198,N_28910,N_29447);
nand UO_2199 (O_2199,N_29688,N_29156);
nor UO_2200 (O_2200,N_29330,N_29649);
or UO_2201 (O_2201,N_29941,N_28951);
xor UO_2202 (O_2202,N_29149,N_29946);
xnor UO_2203 (O_2203,N_29036,N_28809);
or UO_2204 (O_2204,N_28993,N_29915);
xnor UO_2205 (O_2205,N_29045,N_29133);
nand UO_2206 (O_2206,N_29401,N_29049);
xor UO_2207 (O_2207,N_29139,N_29186);
xor UO_2208 (O_2208,N_29593,N_29807);
xor UO_2209 (O_2209,N_28826,N_29199);
xor UO_2210 (O_2210,N_29940,N_29514);
nand UO_2211 (O_2211,N_29675,N_29208);
xor UO_2212 (O_2212,N_29835,N_29410);
xor UO_2213 (O_2213,N_29573,N_29538);
nor UO_2214 (O_2214,N_29837,N_28899);
nand UO_2215 (O_2215,N_29155,N_29064);
and UO_2216 (O_2216,N_29782,N_29872);
nor UO_2217 (O_2217,N_29973,N_29110);
or UO_2218 (O_2218,N_29576,N_29162);
xnor UO_2219 (O_2219,N_29240,N_29337);
nor UO_2220 (O_2220,N_29249,N_29823);
nor UO_2221 (O_2221,N_29706,N_28934);
and UO_2222 (O_2222,N_29948,N_29590);
and UO_2223 (O_2223,N_29824,N_28863);
xor UO_2224 (O_2224,N_29198,N_28951);
or UO_2225 (O_2225,N_29810,N_29046);
or UO_2226 (O_2226,N_28830,N_29489);
or UO_2227 (O_2227,N_29703,N_29088);
or UO_2228 (O_2228,N_29123,N_29515);
or UO_2229 (O_2229,N_29790,N_29624);
nand UO_2230 (O_2230,N_28918,N_29823);
or UO_2231 (O_2231,N_28880,N_29459);
and UO_2232 (O_2232,N_29874,N_29159);
or UO_2233 (O_2233,N_28948,N_29141);
nor UO_2234 (O_2234,N_29427,N_29416);
nor UO_2235 (O_2235,N_29166,N_29158);
and UO_2236 (O_2236,N_29400,N_29203);
xnor UO_2237 (O_2237,N_29435,N_29712);
and UO_2238 (O_2238,N_29387,N_29196);
nor UO_2239 (O_2239,N_28834,N_28874);
or UO_2240 (O_2240,N_29516,N_29046);
xor UO_2241 (O_2241,N_29967,N_28996);
nor UO_2242 (O_2242,N_29407,N_29687);
or UO_2243 (O_2243,N_28962,N_29259);
or UO_2244 (O_2244,N_29151,N_29585);
xor UO_2245 (O_2245,N_29654,N_29291);
nor UO_2246 (O_2246,N_29317,N_29914);
nand UO_2247 (O_2247,N_29292,N_29145);
nor UO_2248 (O_2248,N_29248,N_29193);
nor UO_2249 (O_2249,N_29091,N_29203);
xor UO_2250 (O_2250,N_29324,N_29599);
nand UO_2251 (O_2251,N_29850,N_28856);
nor UO_2252 (O_2252,N_29561,N_29118);
xnor UO_2253 (O_2253,N_29302,N_29593);
nor UO_2254 (O_2254,N_29935,N_29888);
nand UO_2255 (O_2255,N_29706,N_29804);
nor UO_2256 (O_2256,N_28849,N_29199);
xor UO_2257 (O_2257,N_28814,N_29384);
xor UO_2258 (O_2258,N_29125,N_29308);
xnor UO_2259 (O_2259,N_29022,N_29296);
nand UO_2260 (O_2260,N_29592,N_29223);
nor UO_2261 (O_2261,N_28845,N_29560);
and UO_2262 (O_2262,N_29136,N_29027);
nor UO_2263 (O_2263,N_29456,N_28994);
nand UO_2264 (O_2264,N_29676,N_29266);
nand UO_2265 (O_2265,N_29670,N_29831);
nand UO_2266 (O_2266,N_29598,N_29839);
nand UO_2267 (O_2267,N_29596,N_29006);
nor UO_2268 (O_2268,N_29646,N_29319);
nand UO_2269 (O_2269,N_28802,N_29281);
xor UO_2270 (O_2270,N_29474,N_29148);
and UO_2271 (O_2271,N_29133,N_28888);
xor UO_2272 (O_2272,N_29192,N_28948);
nor UO_2273 (O_2273,N_29062,N_29391);
nand UO_2274 (O_2274,N_28813,N_29224);
xnor UO_2275 (O_2275,N_29084,N_29426);
and UO_2276 (O_2276,N_29148,N_29855);
nor UO_2277 (O_2277,N_29872,N_29826);
or UO_2278 (O_2278,N_29436,N_29902);
nor UO_2279 (O_2279,N_29663,N_28913);
nand UO_2280 (O_2280,N_29050,N_29571);
and UO_2281 (O_2281,N_29638,N_29998);
nand UO_2282 (O_2282,N_29966,N_29411);
and UO_2283 (O_2283,N_29228,N_29720);
nand UO_2284 (O_2284,N_29443,N_29138);
nand UO_2285 (O_2285,N_29949,N_29491);
nand UO_2286 (O_2286,N_29123,N_29861);
xnor UO_2287 (O_2287,N_29734,N_29251);
and UO_2288 (O_2288,N_29761,N_29106);
and UO_2289 (O_2289,N_29945,N_29572);
xnor UO_2290 (O_2290,N_29469,N_29116);
xnor UO_2291 (O_2291,N_29805,N_28812);
nand UO_2292 (O_2292,N_29933,N_28900);
nand UO_2293 (O_2293,N_29629,N_29494);
nor UO_2294 (O_2294,N_28867,N_29549);
nand UO_2295 (O_2295,N_29097,N_29698);
nor UO_2296 (O_2296,N_29037,N_28843);
xnor UO_2297 (O_2297,N_29126,N_29991);
nand UO_2298 (O_2298,N_28951,N_29409);
xor UO_2299 (O_2299,N_29617,N_28935);
xnor UO_2300 (O_2300,N_28865,N_29168);
nor UO_2301 (O_2301,N_29655,N_29501);
and UO_2302 (O_2302,N_29133,N_29608);
or UO_2303 (O_2303,N_28979,N_28928);
nand UO_2304 (O_2304,N_29836,N_29672);
nand UO_2305 (O_2305,N_28928,N_28956);
or UO_2306 (O_2306,N_29118,N_29501);
xnor UO_2307 (O_2307,N_29527,N_29988);
nor UO_2308 (O_2308,N_28807,N_29330);
and UO_2309 (O_2309,N_29848,N_29191);
nand UO_2310 (O_2310,N_29398,N_28921);
or UO_2311 (O_2311,N_29768,N_29760);
and UO_2312 (O_2312,N_28802,N_29485);
nand UO_2313 (O_2313,N_29016,N_29211);
and UO_2314 (O_2314,N_29989,N_29958);
nor UO_2315 (O_2315,N_28952,N_29536);
or UO_2316 (O_2316,N_29769,N_29445);
or UO_2317 (O_2317,N_29420,N_29757);
xor UO_2318 (O_2318,N_29168,N_29861);
and UO_2319 (O_2319,N_29121,N_28877);
or UO_2320 (O_2320,N_29198,N_29368);
nand UO_2321 (O_2321,N_29818,N_29746);
nand UO_2322 (O_2322,N_29167,N_29563);
or UO_2323 (O_2323,N_29005,N_29924);
or UO_2324 (O_2324,N_29527,N_29651);
and UO_2325 (O_2325,N_29369,N_29125);
xnor UO_2326 (O_2326,N_29721,N_29387);
nor UO_2327 (O_2327,N_29504,N_29222);
and UO_2328 (O_2328,N_29798,N_29105);
and UO_2329 (O_2329,N_29891,N_29647);
or UO_2330 (O_2330,N_29605,N_29567);
nor UO_2331 (O_2331,N_29378,N_29190);
nand UO_2332 (O_2332,N_29429,N_28953);
nor UO_2333 (O_2333,N_29492,N_29478);
and UO_2334 (O_2334,N_28974,N_29552);
xnor UO_2335 (O_2335,N_28810,N_29779);
nor UO_2336 (O_2336,N_29539,N_29526);
and UO_2337 (O_2337,N_28953,N_29978);
nor UO_2338 (O_2338,N_29890,N_28930);
or UO_2339 (O_2339,N_29931,N_29703);
nand UO_2340 (O_2340,N_29506,N_29929);
nor UO_2341 (O_2341,N_29158,N_29100);
nor UO_2342 (O_2342,N_29280,N_29830);
and UO_2343 (O_2343,N_29303,N_29947);
nor UO_2344 (O_2344,N_29276,N_29834);
xor UO_2345 (O_2345,N_28843,N_29719);
nand UO_2346 (O_2346,N_29813,N_29460);
nand UO_2347 (O_2347,N_29403,N_29264);
and UO_2348 (O_2348,N_29080,N_29190);
xnor UO_2349 (O_2349,N_29718,N_29040);
nor UO_2350 (O_2350,N_28933,N_29581);
and UO_2351 (O_2351,N_29189,N_29245);
nand UO_2352 (O_2352,N_29316,N_28921);
nand UO_2353 (O_2353,N_29591,N_29102);
and UO_2354 (O_2354,N_29781,N_29813);
nor UO_2355 (O_2355,N_29785,N_29779);
nor UO_2356 (O_2356,N_29889,N_29945);
xnor UO_2357 (O_2357,N_29384,N_28811);
xor UO_2358 (O_2358,N_29062,N_29170);
and UO_2359 (O_2359,N_29382,N_29644);
or UO_2360 (O_2360,N_28811,N_29117);
nor UO_2361 (O_2361,N_29030,N_29566);
and UO_2362 (O_2362,N_29651,N_29033);
xor UO_2363 (O_2363,N_29734,N_29716);
and UO_2364 (O_2364,N_28820,N_29077);
nand UO_2365 (O_2365,N_29615,N_29496);
or UO_2366 (O_2366,N_29821,N_28817);
and UO_2367 (O_2367,N_29860,N_29172);
or UO_2368 (O_2368,N_29709,N_29793);
or UO_2369 (O_2369,N_29610,N_29727);
and UO_2370 (O_2370,N_29304,N_28996);
xnor UO_2371 (O_2371,N_28849,N_29349);
and UO_2372 (O_2372,N_29393,N_29465);
xnor UO_2373 (O_2373,N_29774,N_29280);
or UO_2374 (O_2374,N_29070,N_28871);
nor UO_2375 (O_2375,N_29575,N_29164);
xnor UO_2376 (O_2376,N_29934,N_29259);
nand UO_2377 (O_2377,N_28930,N_29981);
and UO_2378 (O_2378,N_29014,N_29571);
nand UO_2379 (O_2379,N_29622,N_29313);
nor UO_2380 (O_2380,N_29381,N_29599);
nor UO_2381 (O_2381,N_29241,N_28828);
nor UO_2382 (O_2382,N_28807,N_29178);
and UO_2383 (O_2383,N_29684,N_29338);
or UO_2384 (O_2384,N_29930,N_29008);
xor UO_2385 (O_2385,N_29251,N_29091);
and UO_2386 (O_2386,N_29552,N_28933);
xnor UO_2387 (O_2387,N_29369,N_29190);
and UO_2388 (O_2388,N_29301,N_29948);
xor UO_2389 (O_2389,N_29722,N_29640);
nor UO_2390 (O_2390,N_29877,N_29619);
nor UO_2391 (O_2391,N_29175,N_28809);
xor UO_2392 (O_2392,N_28934,N_29986);
nor UO_2393 (O_2393,N_29359,N_29374);
nor UO_2394 (O_2394,N_29506,N_28841);
or UO_2395 (O_2395,N_29863,N_29939);
nand UO_2396 (O_2396,N_28919,N_29148);
or UO_2397 (O_2397,N_29443,N_29066);
nor UO_2398 (O_2398,N_29068,N_28878);
and UO_2399 (O_2399,N_29109,N_29680);
nand UO_2400 (O_2400,N_29473,N_29289);
nand UO_2401 (O_2401,N_28922,N_28999);
or UO_2402 (O_2402,N_29957,N_29485);
or UO_2403 (O_2403,N_29210,N_28969);
or UO_2404 (O_2404,N_29743,N_29787);
nand UO_2405 (O_2405,N_29518,N_29853);
and UO_2406 (O_2406,N_29983,N_29614);
or UO_2407 (O_2407,N_28872,N_29215);
or UO_2408 (O_2408,N_29947,N_29769);
nor UO_2409 (O_2409,N_29644,N_29680);
nor UO_2410 (O_2410,N_29203,N_29077);
nand UO_2411 (O_2411,N_29885,N_29287);
xor UO_2412 (O_2412,N_29184,N_29189);
nand UO_2413 (O_2413,N_29716,N_29050);
xnor UO_2414 (O_2414,N_29495,N_29658);
nor UO_2415 (O_2415,N_29778,N_29798);
xnor UO_2416 (O_2416,N_29792,N_29490);
xnor UO_2417 (O_2417,N_29860,N_29456);
and UO_2418 (O_2418,N_29462,N_29407);
or UO_2419 (O_2419,N_29142,N_29855);
nor UO_2420 (O_2420,N_29275,N_29633);
xnor UO_2421 (O_2421,N_28985,N_29478);
nor UO_2422 (O_2422,N_29534,N_29057);
xor UO_2423 (O_2423,N_29790,N_29652);
nand UO_2424 (O_2424,N_29778,N_28966);
and UO_2425 (O_2425,N_28957,N_29935);
or UO_2426 (O_2426,N_29534,N_29638);
and UO_2427 (O_2427,N_29170,N_29175);
nor UO_2428 (O_2428,N_29723,N_28982);
nor UO_2429 (O_2429,N_29098,N_29565);
nor UO_2430 (O_2430,N_29867,N_29046);
nor UO_2431 (O_2431,N_29520,N_28997);
xor UO_2432 (O_2432,N_29504,N_29465);
xnor UO_2433 (O_2433,N_29595,N_29241);
or UO_2434 (O_2434,N_29984,N_29571);
and UO_2435 (O_2435,N_29225,N_29114);
or UO_2436 (O_2436,N_29083,N_29523);
or UO_2437 (O_2437,N_29950,N_28980);
and UO_2438 (O_2438,N_29645,N_29474);
or UO_2439 (O_2439,N_29743,N_29674);
and UO_2440 (O_2440,N_29788,N_29862);
nor UO_2441 (O_2441,N_29918,N_28912);
xnor UO_2442 (O_2442,N_29693,N_29412);
xnor UO_2443 (O_2443,N_29694,N_29347);
or UO_2444 (O_2444,N_29183,N_29482);
and UO_2445 (O_2445,N_29698,N_29437);
nand UO_2446 (O_2446,N_29871,N_29953);
or UO_2447 (O_2447,N_29065,N_29588);
nor UO_2448 (O_2448,N_28802,N_29357);
nor UO_2449 (O_2449,N_29025,N_29888);
and UO_2450 (O_2450,N_29609,N_29391);
or UO_2451 (O_2451,N_29867,N_29595);
xnor UO_2452 (O_2452,N_29479,N_29268);
nor UO_2453 (O_2453,N_29174,N_29689);
or UO_2454 (O_2454,N_29181,N_29872);
and UO_2455 (O_2455,N_29716,N_29129);
nand UO_2456 (O_2456,N_29146,N_29641);
nand UO_2457 (O_2457,N_28990,N_29565);
xor UO_2458 (O_2458,N_28879,N_29223);
or UO_2459 (O_2459,N_29409,N_29217);
xnor UO_2460 (O_2460,N_28870,N_29485);
nand UO_2461 (O_2461,N_28976,N_29160);
xor UO_2462 (O_2462,N_28826,N_28952);
xnor UO_2463 (O_2463,N_29336,N_29178);
nor UO_2464 (O_2464,N_28846,N_29448);
and UO_2465 (O_2465,N_29155,N_28996);
and UO_2466 (O_2466,N_29829,N_29513);
nand UO_2467 (O_2467,N_29304,N_29908);
xor UO_2468 (O_2468,N_28859,N_29069);
xor UO_2469 (O_2469,N_28985,N_28820);
or UO_2470 (O_2470,N_28909,N_28958);
nand UO_2471 (O_2471,N_29437,N_29802);
xor UO_2472 (O_2472,N_29317,N_29910);
nand UO_2473 (O_2473,N_29912,N_29685);
xnor UO_2474 (O_2474,N_28866,N_29604);
or UO_2475 (O_2475,N_29814,N_29967);
or UO_2476 (O_2476,N_29065,N_29573);
xnor UO_2477 (O_2477,N_29670,N_29192);
nand UO_2478 (O_2478,N_29438,N_29698);
nor UO_2479 (O_2479,N_29052,N_28890);
xnor UO_2480 (O_2480,N_29714,N_29936);
xor UO_2481 (O_2481,N_29940,N_29688);
or UO_2482 (O_2482,N_29650,N_29489);
nand UO_2483 (O_2483,N_29631,N_29756);
xnor UO_2484 (O_2484,N_29913,N_29750);
xor UO_2485 (O_2485,N_28933,N_29939);
nor UO_2486 (O_2486,N_29471,N_29367);
or UO_2487 (O_2487,N_29265,N_29151);
or UO_2488 (O_2488,N_29351,N_29516);
and UO_2489 (O_2489,N_29061,N_29706);
or UO_2490 (O_2490,N_28809,N_29255);
or UO_2491 (O_2491,N_29533,N_29707);
or UO_2492 (O_2492,N_29087,N_29971);
or UO_2493 (O_2493,N_29177,N_29365);
nand UO_2494 (O_2494,N_28879,N_29356);
or UO_2495 (O_2495,N_29250,N_29070);
and UO_2496 (O_2496,N_29516,N_29412);
nor UO_2497 (O_2497,N_29107,N_29010);
xnor UO_2498 (O_2498,N_29320,N_29162);
xor UO_2499 (O_2499,N_29950,N_28876);
nor UO_2500 (O_2500,N_29347,N_29406);
xnor UO_2501 (O_2501,N_29983,N_29650);
nor UO_2502 (O_2502,N_29383,N_29507);
and UO_2503 (O_2503,N_28901,N_29014);
xnor UO_2504 (O_2504,N_29251,N_29757);
nor UO_2505 (O_2505,N_28933,N_29063);
xor UO_2506 (O_2506,N_29802,N_29461);
nor UO_2507 (O_2507,N_29289,N_29795);
or UO_2508 (O_2508,N_29646,N_29661);
nand UO_2509 (O_2509,N_29366,N_29677);
xnor UO_2510 (O_2510,N_29235,N_28810);
and UO_2511 (O_2511,N_29115,N_29408);
nor UO_2512 (O_2512,N_29587,N_29981);
and UO_2513 (O_2513,N_29827,N_29529);
and UO_2514 (O_2514,N_29715,N_28999);
nor UO_2515 (O_2515,N_29765,N_28872);
and UO_2516 (O_2516,N_29042,N_29278);
and UO_2517 (O_2517,N_29235,N_29956);
xnor UO_2518 (O_2518,N_29289,N_29524);
nor UO_2519 (O_2519,N_28968,N_29890);
xnor UO_2520 (O_2520,N_29193,N_29754);
and UO_2521 (O_2521,N_29398,N_29507);
nand UO_2522 (O_2522,N_29876,N_29564);
nor UO_2523 (O_2523,N_29811,N_29204);
nor UO_2524 (O_2524,N_29989,N_29188);
xor UO_2525 (O_2525,N_29152,N_29241);
or UO_2526 (O_2526,N_29827,N_29066);
xnor UO_2527 (O_2527,N_29525,N_29206);
nand UO_2528 (O_2528,N_28965,N_28888);
nor UO_2529 (O_2529,N_29374,N_29700);
xor UO_2530 (O_2530,N_28915,N_29976);
or UO_2531 (O_2531,N_29006,N_29976);
and UO_2532 (O_2532,N_29902,N_29978);
nand UO_2533 (O_2533,N_28819,N_29997);
xnor UO_2534 (O_2534,N_29938,N_29980);
nor UO_2535 (O_2535,N_29180,N_29269);
xnor UO_2536 (O_2536,N_29257,N_29437);
and UO_2537 (O_2537,N_29124,N_29621);
or UO_2538 (O_2538,N_29034,N_29709);
nand UO_2539 (O_2539,N_29754,N_29380);
nand UO_2540 (O_2540,N_28800,N_29936);
nand UO_2541 (O_2541,N_29487,N_29937);
nor UO_2542 (O_2542,N_29422,N_29417);
nor UO_2543 (O_2543,N_29451,N_29436);
xor UO_2544 (O_2544,N_29278,N_29943);
nor UO_2545 (O_2545,N_29173,N_29323);
and UO_2546 (O_2546,N_29868,N_29976);
and UO_2547 (O_2547,N_29972,N_29506);
nand UO_2548 (O_2548,N_29100,N_29753);
and UO_2549 (O_2549,N_29870,N_29389);
or UO_2550 (O_2550,N_29601,N_29894);
nor UO_2551 (O_2551,N_29882,N_28920);
and UO_2552 (O_2552,N_29964,N_29184);
xnor UO_2553 (O_2553,N_29842,N_29388);
xnor UO_2554 (O_2554,N_29465,N_29983);
nor UO_2555 (O_2555,N_29554,N_29531);
xor UO_2556 (O_2556,N_29931,N_29296);
and UO_2557 (O_2557,N_29784,N_28836);
nor UO_2558 (O_2558,N_29768,N_29337);
xor UO_2559 (O_2559,N_29057,N_29618);
nand UO_2560 (O_2560,N_29525,N_29866);
nor UO_2561 (O_2561,N_29204,N_28882);
or UO_2562 (O_2562,N_29014,N_29233);
and UO_2563 (O_2563,N_29462,N_29787);
nor UO_2564 (O_2564,N_29896,N_29806);
xnor UO_2565 (O_2565,N_29001,N_28892);
xnor UO_2566 (O_2566,N_29881,N_29032);
nand UO_2567 (O_2567,N_29770,N_29291);
nor UO_2568 (O_2568,N_29281,N_29920);
nor UO_2569 (O_2569,N_29418,N_29398);
nand UO_2570 (O_2570,N_29703,N_29308);
and UO_2571 (O_2571,N_29171,N_28973);
or UO_2572 (O_2572,N_29679,N_28931);
nor UO_2573 (O_2573,N_29868,N_29667);
or UO_2574 (O_2574,N_28922,N_28951);
or UO_2575 (O_2575,N_29739,N_29161);
nor UO_2576 (O_2576,N_29638,N_28851);
nor UO_2577 (O_2577,N_28911,N_29326);
nor UO_2578 (O_2578,N_28938,N_29488);
nand UO_2579 (O_2579,N_29945,N_29677);
and UO_2580 (O_2580,N_28884,N_29765);
or UO_2581 (O_2581,N_29886,N_29235);
nor UO_2582 (O_2582,N_28943,N_29101);
nor UO_2583 (O_2583,N_29584,N_29123);
nand UO_2584 (O_2584,N_29723,N_29148);
nand UO_2585 (O_2585,N_29104,N_29628);
nor UO_2586 (O_2586,N_29335,N_29739);
or UO_2587 (O_2587,N_29545,N_29427);
or UO_2588 (O_2588,N_28900,N_29699);
nand UO_2589 (O_2589,N_29814,N_29479);
and UO_2590 (O_2590,N_29703,N_29375);
nor UO_2591 (O_2591,N_29810,N_28820);
or UO_2592 (O_2592,N_29576,N_29171);
xor UO_2593 (O_2593,N_29079,N_29806);
and UO_2594 (O_2594,N_29986,N_29548);
or UO_2595 (O_2595,N_29013,N_29354);
and UO_2596 (O_2596,N_29265,N_29084);
and UO_2597 (O_2597,N_29536,N_29826);
or UO_2598 (O_2598,N_29435,N_29917);
xor UO_2599 (O_2599,N_29019,N_29230);
xnor UO_2600 (O_2600,N_28951,N_29147);
xor UO_2601 (O_2601,N_28999,N_29266);
xor UO_2602 (O_2602,N_29491,N_29772);
or UO_2603 (O_2603,N_29265,N_29165);
nand UO_2604 (O_2604,N_29457,N_28872);
or UO_2605 (O_2605,N_29748,N_29275);
xnor UO_2606 (O_2606,N_29558,N_29738);
nor UO_2607 (O_2607,N_28811,N_29108);
nor UO_2608 (O_2608,N_29687,N_29063);
or UO_2609 (O_2609,N_29731,N_28947);
nor UO_2610 (O_2610,N_29287,N_29984);
nor UO_2611 (O_2611,N_29147,N_29929);
xnor UO_2612 (O_2612,N_29903,N_29590);
xor UO_2613 (O_2613,N_29427,N_29169);
xnor UO_2614 (O_2614,N_28868,N_29275);
nand UO_2615 (O_2615,N_28897,N_29734);
and UO_2616 (O_2616,N_29712,N_29156);
and UO_2617 (O_2617,N_29211,N_29058);
nand UO_2618 (O_2618,N_29792,N_29234);
nor UO_2619 (O_2619,N_29247,N_29439);
nand UO_2620 (O_2620,N_29055,N_29606);
xor UO_2621 (O_2621,N_29196,N_29688);
and UO_2622 (O_2622,N_29305,N_28982);
and UO_2623 (O_2623,N_29580,N_29418);
nor UO_2624 (O_2624,N_29187,N_29304);
nor UO_2625 (O_2625,N_28931,N_29417);
or UO_2626 (O_2626,N_29926,N_29731);
or UO_2627 (O_2627,N_29379,N_29631);
nand UO_2628 (O_2628,N_29347,N_29552);
nor UO_2629 (O_2629,N_29683,N_29230);
nand UO_2630 (O_2630,N_29678,N_28946);
or UO_2631 (O_2631,N_29355,N_29228);
and UO_2632 (O_2632,N_29526,N_29622);
or UO_2633 (O_2633,N_29009,N_29343);
xnor UO_2634 (O_2634,N_29348,N_29303);
xor UO_2635 (O_2635,N_29068,N_29924);
nor UO_2636 (O_2636,N_29756,N_29001);
or UO_2637 (O_2637,N_29004,N_29805);
and UO_2638 (O_2638,N_28930,N_29416);
and UO_2639 (O_2639,N_28810,N_29173);
nor UO_2640 (O_2640,N_29180,N_29590);
nor UO_2641 (O_2641,N_29879,N_29105);
nand UO_2642 (O_2642,N_28871,N_29262);
xnor UO_2643 (O_2643,N_29561,N_29442);
nand UO_2644 (O_2644,N_29539,N_29729);
and UO_2645 (O_2645,N_29375,N_29963);
nand UO_2646 (O_2646,N_29933,N_29666);
or UO_2647 (O_2647,N_29751,N_29710);
nor UO_2648 (O_2648,N_29029,N_29380);
xnor UO_2649 (O_2649,N_29466,N_29813);
nand UO_2650 (O_2650,N_29579,N_29689);
xnor UO_2651 (O_2651,N_29631,N_29866);
nor UO_2652 (O_2652,N_29416,N_29970);
and UO_2653 (O_2653,N_28836,N_29025);
xnor UO_2654 (O_2654,N_29776,N_28875);
or UO_2655 (O_2655,N_28910,N_29008);
or UO_2656 (O_2656,N_29522,N_29004);
nor UO_2657 (O_2657,N_29091,N_29258);
xnor UO_2658 (O_2658,N_29700,N_28862);
xnor UO_2659 (O_2659,N_29334,N_29325);
or UO_2660 (O_2660,N_29957,N_29725);
nand UO_2661 (O_2661,N_29451,N_29701);
nand UO_2662 (O_2662,N_29813,N_29915);
xnor UO_2663 (O_2663,N_29252,N_29936);
nor UO_2664 (O_2664,N_29536,N_29679);
nor UO_2665 (O_2665,N_29118,N_29867);
xor UO_2666 (O_2666,N_29564,N_29806);
nor UO_2667 (O_2667,N_29760,N_28950);
and UO_2668 (O_2668,N_29393,N_29329);
nor UO_2669 (O_2669,N_29429,N_29119);
or UO_2670 (O_2670,N_29606,N_29644);
xnor UO_2671 (O_2671,N_28862,N_29973);
nand UO_2672 (O_2672,N_29430,N_28835);
xor UO_2673 (O_2673,N_29643,N_29436);
nor UO_2674 (O_2674,N_29516,N_28948);
xnor UO_2675 (O_2675,N_29001,N_29956);
nand UO_2676 (O_2676,N_29084,N_29111);
or UO_2677 (O_2677,N_29602,N_29114);
nand UO_2678 (O_2678,N_28929,N_29861);
nor UO_2679 (O_2679,N_28951,N_29962);
nor UO_2680 (O_2680,N_29313,N_29299);
and UO_2681 (O_2681,N_28805,N_29865);
nand UO_2682 (O_2682,N_29708,N_28908);
nand UO_2683 (O_2683,N_29884,N_29984);
xor UO_2684 (O_2684,N_29271,N_29277);
and UO_2685 (O_2685,N_29310,N_29768);
and UO_2686 (O_2686,N_29142,N_29784);
and UO_2687 (O_2687,N_29448,N_29446);
nand UO_2688 (O_2688,N_29035,N_29377);
and UO_2689 (O_2689,N_29089,N_29656);
and UO_2690 (O_2690,N_28818,N_29113);
nor UO_2691 (O_2691,N_29108,N_29425);
and UO_2692 (O_2692,N_29626,N_29549);
nand UO_2693 (O_2693,N_29631,N_29050);
and UO_2694 (O_2694,N_28951,N_29218);
nor UO_2695 (O_2695,N_29950,N_29992);
xnor UO_2696 (O_2696,N_28858,N_29430);
and UO_2697 (O_2697,N_29863,N_29376);
or UO_2698 (O_2698,N_29679,N_29427);
and UO_2699 (O_2699,N_29350,N_29234);
or UO_2700 (O_2700,N_29173,N_29099);
or UO_2701 (O_2701,N_29986,N_29571);
and UO_2702 (O_2702,N_29255,N_29518);
nor UO_2703 (O_2703,N_29529,N_29500);
nand UO_2704 (O_2704,N_29242,N_29958);
nand UO_2705 (O_2705,N_29719,N_29758);
xor UO_2706 (O_2706,N_29112,N_29562);
xnor UO_2707 (O_2707,N_29259,N_29463);
xnor UO_2708 (O_2708,N_29365,N_29220);
xor UO_2709 (O_2709,N_28977,N_29088);
xnor UO_2710 (O_2710,N_29170,N_29098);
and UO_2711 (O_2711,N_29630,N_28966);
or UO_2712 (O_2712,N_29357,N_29247);
xor UO_2713 (O_2713,N_29544,N_29804);
and UO_2714 (O_2714,N_29768,N_29771);
nand UO_2715 (O_2715,N_28966,N_29482);
and UO_2716 (O_2716,N_29728,N_28917);
or UO_2717 (O_2717,N_29487,N_29600);
or UO_2718 (O_2718,N_29925,N_29861);
nor UO_2719 (O_2719,N_29912,N_29214);
xor UO_2720 (O_2720,N_29625,N_29468);
or UO_2721 (O_2721,N_29960,N_29481);
and UO_2722 (O_2722,N_29213,N_28916);
or UO_2723 (O_2723,N_29688,N_29693);
or UO_2724 (O_2724,N_29578,N_28939);
or UO_2725 (O_2725,N_29901,N_29632);
or UO_2726 (O_2726,N_28959,N_28871);
nand UO_2727 (O_2727,N_29119,N_29106);
or UO_2728 (O_2728,N_28802,N_29778);
or UO_2729 (O_2729,N_29304,N_29488);
nor UO_2730 (O_2730,N_28944,N_29031);
nor UO_2731 (O_2731,N_29574,N_28933);
nor UO_2732 (O_2732,N_29618,N_29761);
and UO_2733 (O_2733,N_29812,N_29068);
and UO_2734 (O_2734,N_29907,N_29683);
or UO_2735 (O_2735,N_28859,N_29832);
or UO_2736 (O_2736,N_29506,N_29330);
nor UO_2737 (O_2737,N_28937,N_29399);
xnor UO_2738 (O_2738,N_29051,N_29375);
nor UO_2739 (O_2739,N_29294,N_28969);
and UO_2740 (O_2740,N_29634,N_29559);
or UO_2741 (O_2741,N_28946,N_29186);
xnor UO_2742 (O_2742,N_29134,N_29783);
xor UO_2743 (O_2743,N_29536,N_29650);
xor UO_2744 (O_2744,N_28985,N_29643);
nand UO_2745 (O_2745,N_29049,N_29976);
xnor UO_2746 (O_2746,N_29190,N_29357);
nor UO_2747 (O_2747,N_29214,N_29780);
nor UO_2748 (O_2748,N_29102,N_29204);
nor UO_2749 (O_2749,N_29001,N_29174);
xor UO_2750 (O_2750,N_29351,N_29505);
nand UO_2751 (O_2751,N_29304,N_29277);
nor UO_2752 (O_2752,N_28950,N_28981);
nand UO_2753 (O_2753,N_28868,N_29267);
xor UO_2754 (O_2754,N_29927,N_29774);
nand UO_2755 (O_2755,N_29314,N_28919);
nand UO_2756 (O_2756,N_28915,N_29800);
nor UO_2757 (O_2757,N_29532,N_29523);
or UO_2758 (O_2758,N_29440,N_29598);
nor UO_2759 (O_2759,N_28938,N_28977);
and UO_2760 (O_2760,N_29075,N_28846);
nor UO_2761 (O_2761,N_29936,N_29618);
nand UO_2762 (O_2762,N_29592,N_29239);
and UO_2763 (O_2763,N_29379,N_29581);
or UO_2764 (O_2764,N_29446,N_29874);
nand UO_2765 (O_2765,N_29511,N_29035);
nor UO_2766 (O_2766,N_29744,N_29683);
or UO_2767 (O_2767,N_29389,N_29836);
or UO_2768 (O_2768,N_29645,N_29651);
xnor UO_2769 (O_2769,N_29707,N_28831);
nand UO_2770 (O_2770,N_29224,N_29413);
or UO_2771 (O_2771,N_29911,N_29381);
nor UO_2772 (O_2772,N_29810,N_29504);
nor UO_2773 (O_2773,N_29408,N_29925);
or UO_2774 (O_2774,N_29531,N_29692);
and UO_2775 (O_2775,N_29895,N_29938);
nand UO_2776 (O_2776,N_29685,N_29415);
nor UO_2777 (O_2777,N_29445,N_29554);
nor UO_2778 (O_2778,N_29517,N_29309);
nand UO_2779 (O_2779,N_28980,N_29819);
or UO_2780 (O_2780,N_29799,N_29486);
nand UO_2781 (O_2781,N_29916,N_29268);
xnor UO_2782 (O_2782,N_29969,N_29510);
and UO_2783 (O_2783,N_29271,N_29548);
and UO_2784 (O_2784,N_28848,N_29846);
xnor UO_2785 (O_2785,N_29180,N_29620);
or UO_2786 (O_2786,N_29207,N_29258);
or UO_2787 (O_2787,N_29808,N_29926);
or UO_2788 (O_2788,N_28844,N_28942);
nand UO_2789 (O_2789,N_29693,N_29466);
and UO_2790 (O_2790,N_29782,N_29760);
or UO_2791 (O_2791,N_28960,N_29268);
and UO_2792 (O_2792,N_29729,N_29488);
xor UO_2793 (O_2793,N_29560,N_29344);
nand UO_2794 (O_2794,N_29372,N_29695);
and UO_2795 (O_2795,N_29650,N_28833);
and UO_2796 (O_2796,N_29892,N_29738);
xnor UO_2797 (O_2797,N_29189,N_29547);
nor UO_2798 (O_2798,N_29819,N_29152);
nand UO_2799 (O_2799,N_29088,N_29119);
nor UO_2800 (O_2800,N_29693,N_29942);
nand UO_2801 (O_2801,N_29748,N_28910);
xor UO_2802 (O_2802,N_29166,N_29437);
nand UO_2803 (O_2803,N_29900,N_29271);
nor UO_2804 (O_2804,N_29799,N_29952);
xor UO_2805 (O_2805,N_28939,N_29824);
nor UO_2806 (O_2806,N_29847,N_29563);
nor UO_2807 (O_2807,N_29677,N_29989);
or UO_2808 (O_2808,N_28911,N_28864);
xnor UO_2809 (O_2809,N_29837,N_28957);
and UO_2810 (O_2810,N_29760,N_29975);
or UO_2811 (O_2811,N_29576,N_29079);
nor UO_2812 (O_2812,N_29315,N_29936);
or UO_2813 (O_2813,N_28997,N_29145);
and UO_2814 (O_2814,N_29806,N_29627);
nand UO_2815 (O_2815,N_29795,N_28914);
nand UO_2816 (O_2816,N_29356,N_28805);
xor UO_2817 (O_2817,N_28928,N_29221);
or UO_2818 (O_2818,N_29769,N_29447);
xnor UO_2819 (O_2819,N_29138,N_29160);
or UO_2820 (O_2820,N_29798,N_29049);
or UO_2821 (O_2821,N_29142,N_29052);
xnor UO_2822 (O_2822,N_29678,N_29376);
xnor UO_2823 (O_2823,N_29981,N_29106);
nor UO_2824 (O_2824,N_29246,N_29420);
or UO_2825 (O_2825,N_29065,N_29369);
or UO_2826 (O_2826,N_29726,N_29668);
nand UO_2827 (O_2827,N_29294,N_29593);
or UO_2828 (O_2828,N_29445,N_29831);
nand UO_2829 (O_2829,N_29441,N_29912);
or UO_2830 (O_2830,N_29544,N_29981);
or UO_2831 (O_2831,N_29854,N_29428);
and UO_2832 (O_2832,N_29915,N_28951);
nand UO_2833 (O_2833,N_29968,N_29867);
or UO_2834 (O_2834,N_29289,N_29139);
or UO_2835 (O_2835,N_28989,N_29371);
xnor UO_2836 (O_2836,N_29470,N_29947);
nor UO_2837 (O_2837,N_29970,N_29860);
nor UO_2838 (O_2838,N_29427,N_28876);
nand UO_2839 (O_2839,N_29869,N_29961);
nand UO_2840 (O_2840,N_29833,N_29631);
and UO_2841 (O_2841,N_29121,N_29905);
or UO_2842 (O_2842,N_28820,N_29916);
or UO_2843 (O_2843,N_29618,N_29435);
xor UO_2844 (O_2844,N_29863,N_29227);
xnor UO_2845 (O_2845,N_29430,N_29747);
nor UO_2846 (O_2846,N_29689,N_29587);
nand UO_2847 (O_2847,N_29384,N_28895);
xor UO_2848 (O_2848,N_29849,N_29631);
and UO_2849 (O_2849,N_28904,N_28887);
xnor UO_2850 (O_2850,N_29180,N_28908);
and UO_2851 (O_2851,N_29024,N_29846);
or UO_2852 (O_2852,N_28810,N_29819);
xnor UO_2853 (O_2853,N_28822,N_28989);
nor UO_2854 (O_2854,N_29272,N_29858);
or UO_2855 (O_2855,N_29092,N_29849);
xnor UO_2856 (O_2856,N_29786,N_29179);
nor UO_2857 (O_2857,N_29625,N_29365);
nand UO_2858 (O_2858,N_29649,N_29810);
nand UO_2859 (O_2859,N_29850,N_29301);
nor UO_2860 (O_2860,N_29453,N_29310);
nor UO_2861 (O_2861,N_29523,N_29748);
nor UO_2862 (O_2862,N_29209,N_29040);
nand UO_2863 (O_2863,N_29687,N_29712);
xnor UO_2864 (O_2864,N_28921,N_29439);
nor UO_2865 (O_2865,N_29611,N_28818);
or UO_2866 (O_2866,N_29529,N_29229);
nand UO_2867 (O_2867,N_29125,N_29494);
or UO_2868 (O_2868,N_29240,N_28825);
nand UO_2869 (O_2869,N_29060,N_29644);
nor UO_2870 (O_2870,N_29365,N_29403);
xnor UO_2871 (O_2871,N_29011,N_29236);
and UO_2872 (O_2872,N_29369,N_29788);
or UO_2873 (O_2873,N_29207,N_29808);
xnor UO_2874 (O_2874,N_28849,N_28915);
nor UO_2875 (O_2875,N_29314,N_29215);
xor UO_2876 (O_2876,N_29475,N_29151);
and UO_2877 (O_2877,N_29372,N_28838);
nand UO_2878 (O_2878,N_29726,N_29138);
xnor UO_2879 (O_2879,N_29830,N_28941);
xor UO_2880 (O_2880,N_29060,N_29996);
and UO_2881 (O_2881,N_29896,N_29170);
nand UO_2882 (O_2882,N_29452,N_28833);
or UO_2883 (O_2883,N_29712,N_29205);
and UO_2884 (O_2884,N_29245,N_29095);
and UO_2885 (O_2885,N_29401,N_29447);
nand UO_2886 (O_2886,N_29584,N_29712);
and UO_2887 (O_2887,N_29596,N_28999);
xnor UO_2888 (O_2888,N_29239,N_28873);
xor UO_2889 (O_2889,N_29103,N_29946);
and UO_2890 (O_2890,N_29640,N_29401);
xor UO_2891 (O_2891,N_29307,N_28927);
or UO_2892 (O_2892,N_29359,N_29672);
and UO_2893 (O_2893,N_29514,N_29753);
or UO_2894 (O_2894,N_29954,N_29960);
nor UO_2895 (O_2895,N_29335,N_29922);
and UO_2896 (O_2896,N_29235,N_29806);
xnor UO_2897 (O_2897,N_29756,N_28944);
or UO_2898 (O_2898,N_29051,N_29162);
xnor UO_2899 (O_2899,N_29856,N_29707);
xnor UO_2900 (O_2900,N_28928,N_29094);
nand UO_2901 (O_2901,N_29995,N_29049);
nor UO_2902 (O_2902,N_29682,N_29158);
or UO_2903 (O_2903,N_29572,N_29728);
and UO_2904 (O_2904,N_29177,N_29282);
nand UO_2905 (O_2905,N_29373,N_29770);
or UO_2906 (O_2906,N_29153,N_29687);
xnor UO_2907 (O_2907,N_29057,N_29736);
and UO_2908 (O_2908,N_29408,N_29770);
or UO_2909 (O_2909,N_29415,N_29368);
nor UO_2910 (O_2910,N_28951,N_29180);
nor UO_2911 (O_2911,N_29212,N_29262);
nor UO_2912 (O_2912,N_29150,N_29506);
or UO_2913 (O_2913,N_29477,N_29789);
and UO_2914 (O_2914,N_29871,N_28972);
nand UO_2915 (O_2915,N_29315,N_29806);
xor UO_2916 (O_2916,N_28997,N_29027);
or UO_2917 (O_2917,N_29515,N_29729);
or UO_2918 (O_2918,N_29539,N_29821);
or UO_2919 (O_2919,N_28878,N_28835);
nand UO_2920 (O_2920,N_29838,N_28898);
or UO_2921 (O_2921,N_29996,N_28958);
xor UO_2922 (O_2922,N_28883,N_29114);
nor UO_2923 (O_2923,N_29952,N_29062);
or UO_2924 (O_2924,N_29019,N_29309);
or UO_2925 (O_2925,N_28914,N_29676);
and UO_2926 (O_2926,N_29222,N_29077);
nor UO_2927 (O_2927,N_29608,N_29929);
or UO_2928 (O_2928,N_29435,N_28918);
nand UO_2929 (O_2929,N_29510,N_29638);
or UO_2930 (O_2930,N_29530,N_29267);
and UO_2931 (O_2931,N_29803,N_29972);
nor UO_2932 (O_2932,N_29937,N_29858);
nor UO_2933 (O_2933,N_29141,N_29823);
nand UO_2934 (O_2934,N_28947,N_29207);
nand UO_2935 (O_2935,N_29734,N_29967);
nor UO_2936 (O_2936,N_29599,N_29140);
or UO_2937 (O_2937,N_29281,N_29745);
or UO_2938 (O_2938,N_29195,N_29850);
nor UO_2939 (O_2939,N_29005,N_29829);
and UO_2940 (O_2940,N_29521,N_29111);
nand UO_2941 (O_2941,N_29354,N_29355);
nor UO_2942 (O_2942,N_29350,N_29553);
and UO_2943 (O_2943,N_29539,N_29340);
nand UO_2944 (O_2944,N_28883,N_29700);
xnor UO_2945 (O_2945,N_28851,N_29043);
nor UO_2946 (O_2946,N_29650,N_29597);
nor UO_2947 (O_2947,N_29207,N_29576);
and UO_2948 (O_2948,N_29365,N_29163);
nand UO_2949 (O_2949,N_29695,N_29281);
xor UO_2950 (O_2950,N_29207,N_29079);
or UO_2951 (O_2951,N_29053,N_29432);
or UO_2952 (O_2952,N_29759,N_29850);
and UO_2953 (O_2953,N_29296,N_29959);
xor UO_2954 (O_2954,N_29126,N_29653);
and UO_2955 (O_2955,N_29094,N_29274);
xor UO_2956 (O_2956,N_29038,N_29115);
and UO_2957 (O_2957,N_29699,N_29414);
xor UO_2958 (O_2958,N_28982,N_29079);
or UO_2959 (O_2959,N_29530,N_29352);
xor UO_2960 (O_2960,N_28849,N_29839);
nand UO_2961 (O_2961,N_29876,N_29489);
or UO_2962 (O_2962,N_29821,N_29977);
and UO_2963 (O_2963,N_29573,N_29353);
nor UO_2964 (O_2964,N_29828,N_29997);
xor UO_2965 (O_2965,N_29897,N_28892);
nor UO_2966 (O_2966,N_29872,N_29535);
nand UO_2967 (O_2967,N_29305,N_29870);
or UO_2968 (O_2968,N_29441,N_29933);
nor UO_2969 (O_2969,N_29466,N_29826);
and UO_2970 (O_2970,N_29241,N_29704);
xor UO_2971 (O_2971,N_28887,N_29453);
nand UO_2972 (O_2972,N_29681,N_29200);
or UO_2973 (O_2973,N_29148,N_29108);
or UO_2974 (O_2974,N_29799,N_28851);
nand UO_2975 (O_2975,N_29581,N_29908);
nand UO_2976 (O_2976,N_28941,N_29993);
xnor UO_2977 (O_2977,N_29755,N_29186);
nor UO_2978 (O_2978,N_29610,N_29942);
nand UO_2979 (O_2979,N_29568,N_29605);
or UO_2980 (O_2980,N_28837,N_28856);
nand UO_2981 (O_2981,N_29042,N_29254);
nor UO_2982 (O_2982,N_29131,N_29192);
nor UO_2983 (O_2983,N_29334,N_28981);
nor UO_2984 (O_2984,N_29534,N_29171);
and UO_2985 (O_2985,N_29958,N_29820);
or UO_2986 (O_2986,N_29443,N_28867);
nor UO_2987 (O_2987,N_29892,N_29773);
xor UO_2988 (O_2988,N_29599,N_29058);
xnor UO_2989 (O_2989,N_29872,N_28868);
nor UO_2990 (O_2990,N_29774,N_29380);
nand UO_2991 (O_2991,N_29682,N_29449);
and UO_2992 (O_2992,N_29755,N_29087);
and UO_2993 (O_2993,N_29726,N_29380);
nor UO_2994 (O_2994,N_29475,N_29907);
nor UO_2995 (O_2995,N_29301,N_29387);
or UO_2996 (O_2996,N_28957,N_29662);
nor UO_2997 (O_2997,N_29734,N_29488);
nand UO_2998 (O_2998,N_29209,N_29891);
xnor UO_2999 (O_2999,N_29931,N_29605);
or UO_3000 (O_3000,N_29585,N_29594);
and UO_3001 (O_3001,N_29443,N_29900);
nand UO_3002 (O_3002,N_29114,N_29307);
nor UO_3003 (O_3003,N_29331,N_29366);
or UO_3004 (O_3004,N_29959,N_29420);
nor UO_3005 (O_3005,N_29804,N_29923);
nand UO_3006 (O_3006,N_28886,N_29478);
nor UO_3007 (O_3007,N_29421,N_28942);
or UO_3008 (O_3008,N_29690,N_29969);
and UO_3009 (O_3009,N_29165,N_29222);
nor UO_3010 (O_3010,N_29191,N_29955);
or UO_3011 (O_3011,N_28904,N_29882);
or UO_3012 (O_3012,N_29937,N_29266);
xor UO_3013 (O_3013,N_29952,N_29664);
nand UO_3014 (O_3014,N_29469,N_29693);
xnor UO_3015 (O_3015,N_28924,N_28858);
or UO_3016 (O_3016,N_29931,N_29589);
nor UO_3017 (O_3017,N_29819,N_29616);
xnor UO_3018 (O_3018,N_29520,N_28850);
nor UO_3019 (O_3019,N_29555,N_29533);
nor UO_3020 (O_3020,N_29370,N_29455);
xnor UO_3021 (O_3021,N_29148,N_29621);
and UO_3022 (O_3022,N_29023,N_29496);
and UO_3023 (O_3023,N_29875,N_28961);
nand UO_3024 (O_3024,N_29008,N_29387);
or UO_3025 (O_3025,N_29442,N_29163);
or UO_3026 (O_3026,N_28822,N_29079);
nor UO_3027 (O_3027,N_28929,N_29659);
and UO_3028 (O_3028,N_29360,N_29782);
xnor UO_3029 (O_3029,N_29019,N_29505);
and UO_3030 (O_3030,N_29718,N_29738);
nand UO_3031 (O_3031,N_28919,N_29516);
xnor UO_3032 (O_3032,N_29611,N_29545);
or UO_3033 (O_3033,N_29537,N_29241);
xor UO_3034 (O_3034,N_29954,N_29539);
xnor UO_3035 (O_3035,N_29371,N_29749);
xnor UO_3036 (O_3036,N_28826,N_29638);
or UO_3037 (O_3037,N_29680,N_29879);
nand UO_3038 (O_3038,N_29963,N_29640);
and UO_3039 (O_3039,N_29597,N_29039);
or UO_3040 (O_3040,N_29190,N_29381);
and UO_3041 (O_3041,N_29931,N_29426);
xnor UO_3042 (O_3042,N_29830,N_29393);
and UO_3043 (O_3043,N_29830,N_29420);
xor UO_3044 (O_3044,N_29624,N_29960);
xor UO_3045 (O_3045,N_29018,N_29151);
xnor UO_3046 (O_3046,N_28888,N_29672);
or UO_3047 (O_3047,N_29019,N_29991);
or UO_3048 (O_3048,N_29600,N_29059);
nand UO_3049 (O_3049,N_29724,N_29080);
nor UO_3050 (O_3050,N_29093,N_29055);
or UO_3051 (O_3051,N_28934,N_29159);
nand UO_3052 (O_3052,N_29090,N_29066);
nor UO_3053 (O_3053,N_28801,N_28884);
nor UO_3054 (O_3054,N_28957,N_29097);
xor UO_3055 (O_3055,N_29148,N_29600);
and UO_3056 (O_3056,N_28902,N_28986);
or UO_3057 (O_3057,N_29081,N_29553);
nor UO_3058 (O_3058,N_29482,N_29465);
or UO_3059 (O_3059,N_29164,N_29177);
and UO_3060 (O_3060,N_28947,N_29311);
nor UO_3061 (O_3061,N_29229,N_29033);
or UO_3062 (O_3062,N_29015,N_29025);
and UO_3063 (O_3063,N_29815,N_29015);
nor UO_3064 (O_3064,N_29593,N_29421);
nand UO_3065 (O_3065,N_29535,N_28844);
nand UO_3066 (O_3066,N_29435,N_29237);
nor UO_3067 (O_3067,N_29101,N_28869);
nor UO_3068 (O_3068,N_29110,N_29948);
nor UO_3069 (O_3069,N_29821,N_29741);
xnor UO_3070 (O_3070,N_29907,N_28921);
or UO_3071 (O_3071,N_29877,N_29125);
or UO_3072 (O_3072,N_29511,N_29453);
nor UO_3073 (O_3073,N_29437,N_29707);
or UO_3074 (O_3074,N_29960,N_29955);
or UO_3075 (O_3075,N_29724,N_29692);
nor UO_3076 (O_3076,N_29787,N_28926);
nor UO_3077 (O_3077,N_29274,N_29875);
xor UO_3078 (O_3078,N_29800,N_29983);
xor UO_3079 (O_3079,N_29509,N_29212);
and UO_3080 (O_3080,N_29783,N_29085);
xor UO_3081 (O_3081,N_29419,N_28983);
xnor UO_3082 (O_3082,N_28944,N_29268);
and UO_3083 (O_3083,N_29035,N_29841);
xnor UO_3084 (O_3084,N_29828,N_29136);
nand UO_3085 (O_3085,N_29909,N_28833);
and UO_3086 (O_3086,N_29165,N_29420);
xnor UO_3087 (O_3087,N_29318,N_29155);
or UO_3088 (O_3088,N_29923,N_29299);
and UO_3089 (O_3089,N_29911,N_29937);
and UO_3090 (O_3090,N_29841,N_29803);
xor UO_3091 (O_3091,N_29795,N_29503);
xor UO_3092 (O_3092,N_29379,N_28814);
xnor UO_3093 (O_3093,N_28911,N_29327);
nor UO_3094 (O_3094,N_29179,N_29305);
and UO_3095 (O_3095,N_29684,N_28902);
or UO_3096 (O_3096,N_28846,N_29461);
nor UO_3097 (O_3097,N_28822,N_29156);
or UO_3098 (O_3098,N_29505,N_29732);
and UO_3099 (O_3099,N_29027,N_29214);
and UO_3100 (O_3100,N_28993,N_29237);
and UO_3101 (O_3101,N_29672,N_29403);
or UO_3102 (O_3102,N_29487,N_28818);
nand UO_3103 (O_3103,N_29453,N_29803);
xnor UO_3104 (O_3104,N_28940,N_29024);
and UO_3105 (O_3105,N_29568,N_29407);
xor UO_3106 (O_3106,N_29458,N_28817);
or UO_3107 (O_3107,N_29520,N_29478);
nor UO_3108 (O_3108,N_29228,N_29286);
nor UO_3109 (O_3109,N_28821,N_29804);
xor UO_3110 (O_3110,N_28807,N_29955);
or UO_3111 (O_3111,N_29355,N_29327);
nor UO_3112 (O_3112,N_29551,N_29225);
nor UO_3113 (O_3113,N_29249,N_29253);
and UO_3114 (O_3114,N_28953,N_29655);
nand UO_3115 (O_3115,N_28803,N_29636);
or UO_3116 (O_3116,N_29369,N_29774);
and UO_3117 (O_3117,N_29991,N_29681);
nand UO_3118 (O_3118,N_29879,N_29532);
nor UO_3119 (O_3119,N_29584,N_28868);
or UO_3120 (O_3120,N_28805,N_29579);
nor UO_3121 (O_3121,N_29949,N_29438);
nand UO_3122 (O_3122,N_29051,N_29464);
xnor UO_3123 (O_3123,N_29492,N_29155);
nand UO_3124 (O_3124,N_29579,N_29270);
nor UO_3125 (O_3125,N_29929,N_29365);
and UO_3126 (O_3126,N_28912,N_29961);
and UO_3127 (O_3127,N_29040,N_29769);
and UO_3128 (O_3128,N_29404,N_29411);
xor UO_3129 (O_3129,N_29523,N_29487);
or UO_3130 (O_3130,N_28960,N_29521);
and UO_3131 (O_3131,N_29801,N_29960);
nor UO_3132 (O_3132,N_29940,N_29294);
nand UO_3133 (O_3133,N_28908,N_29593);
or UO_3134 (O_3134,N_29642,N_29561);
nand UO_3135 (O_3135,N_29603,N_29379);
or UO_3136 (O_3136,N_28909,N_29600);
or UO_3137 (O_3137,N_29824,N_29860);
and UO_3138 (O_3138,N_29724,N_28946);
nor UO_3139 (O_3139,N_29280,N_29974);
xor UO_3140 (O_3140,N_28897,N_29839);
or UO_3141 (O_3141,N_29158,N_29355);
or UO_3142 (O_3142,N_29668,N_28940);
nor UO_3143 (O_3143,N_29381,N_29948);
nand UO_3144 (O_3144,N_29812,N_29508);
and UO_3145 (O_3145,N_29434,N_29473);
or UO_3146 (O_3146,N_29202,N_28973);
nor UO_3147 (O_3147,N_29950,N_29496);
nand UO_3148 (O_3148,N_29783,N_29478);
or UO_3149 (O_3149,N_29300,N_29358);
and UO_3150 (O_3150,N_29296,N_29025);
or UO_3151 (O_3151,N_29179,N_29283);
xor UO_3152 (O_3152,N_28981,N_29460);
nand UO_3153 (O_3153,N_29549,N_29879);
and UO_3154 (O_3154,N_29773,N_28903);
or UO_3155 (O_3155,N_29543,N_29275);
or UO_3156 (O_3156,N_29461,N_29233);
xnor UO_3157 (O_3157,N_29889,N_29300);
or UO_3158 (O_3158,N_29108,N_29041);
nor UO_3159 (O_3159,N_28940,N_29266);
and UO_3160 (O_3160,N_28809,N_29148);
xnor UO_3161 (O_3161,N_28802,N_29024);
xnor UO_3162 (O_3162,N_29481,N_29211);
and UO_3163 (O_3163,N_28917,N_29870);
xnor UO_3164 (O_3164,N_28865,N_29528);
nand UO_3165 (O_3165,N_29626,N_29393);
nor UO_3166 (O_3166,N_29030,N_29585);
or UO_3167 (O_3167,N_29872,N_29684);
and UO_3168 (O_3168,N_29969,N_28927);
nand UO_3169 (O_3169,N_28856,N_29791);
nor UO_3170 (O_3170,N_29675,N_29360);
and UO_3171 (O_3171,N_29775,N_29925);
nand UO_3172 (O_3172,N_29676,N_29639);
and UO_3173 (O_3173,N_29380,N_29664);
and UO_3174 (O_3174,N_29663,N_29046);
nand UO_3175 (O_3175,N_29189,N_29831);
xnor UO_3176 (O_3176,N_28881,N_29285);
and UO_3177 (O_3177,N_29121,N_29489);
nand UO_3178 (O_3178,N_29669,N_29041);
and UO_3179 (O_3179,N_29834,N_29582);
nand UO_3180 (O_3180,N_29271,N_29557);
nand UO_3181 (O_3181,N_29623,N_29286);
or UO_3182 (O_3182,N_29068,N_29073);
xor UO_3183 (O_3183,N_29857,N_29092);
xor UO_3184 (O_3184,N_29620,N_29101);
xor UO_3185 (O_3185,N_29033,N_29044);
or UO_3186 (O_3186,N_29519,N_29249);
and UO_3187 (O_3187,N_28846,N_29307);
or UO_3188 (O_3188,N_29635,N_28897);
nand UO_3189 (O_3189,N_29558,N_29932);
xnor UO_3190 (O_3190,N_29201,N_29698);
and UO_3191 (O_3191,N_29689,N_29902);
and UO_3192 (O_3192,N_29373,N_29064);
xnor UO_3193 (O_3193,N_29229,N_28943);
nand UO_3194 (O_3194,N_29936,N_29472);
nand UO_3195 (O_3195,N_29464,N_29390);
and UO_3196 (O_3196,N_29142,N_29810);
nand UO_3197 (O_3197,N_29742,N_29763);
or UO_3198 (O_3198,N_29239,N_29768);
nor UO_3199 (O_3199,N_29137,N_29627);
or UO_3200 (O_3200,N_28936,N_28925);
nand UO_3201 (O_3201,N_28828,N_29117);
nand UO_3202 (O_3202,N_29807,N_29824);
nand UO_3203 (O_3203,N_29265,N_29680);
and UO_3204 (O_3204,N_29072,N_29428);
and UO_3205 (O_3205,N_29745,N_29114);
nand UO_3206 (O_3206,N_29556,N_29990);
and UO_3207 (O_3207,N_29427,N_29948);
nand UO_3208 (O_3208,N_28906,N_29875);
and UO_3209 (O_3209,N_29220,N_29888);
nand UO_3210 (O_3210,N_29941,N_29206);
nor UO_3211 (O_3211,N_29417,N_29733);
or UO_3212 (O_3212,N_29126,N_28818);
xor UO_3213 (O_3213,N_28883,N_29186);
xor UO_3214 (O_3214,N_28815,N_29104);
xor UO_3215 (O_3215,N_29772,N_29392);
or UO_3216 (O_3216,N_29617,N_29224);
and UO_3217 (O_3217,N_29235,N_29099);
nor UO_3218 (O_3218,N_29274,N_29038);
and UO_3219 (O_3219,N_29945,N_29101);
and UO_3220 (O_3220,N_29657,N_29953);
and UO_3221 (O_3221,N_28832,N_29332);
nand UO_3222 (O_3222,N_29967,N_29500);
or UO_3223 (O_3223,N_29875,N_29497);
nor UO_3224 (O_3224,N_29066,N_29824);
xor UO_3225 (O_3225,N_28872,N_29353);
and UO_3226 (O_3226,N_29715,N_29881);
nand UO_3227 (O_3227,N_28986,N_29787);
and UO_3228 (O_3228,N_29958,N_29785);
or UO_3229 (O_3229,N_29684,N_28850);
and UO_3230 (O_3230,N_29893,N_29435);
xnor UO_3231 (O_3231,N_29248,N_29200);
nor UO_3232 (O_3232,N_29540,N_29363);
or UO_3233 (O_3233,N_29578,N_29530);
nand UO_3234 (O_3234,N_29695,N_29370);
and UO_3235 (O_3235,N_29559,N_29328);
or UO_3236 (O_3236,N_29047,N_29752);
or UO_3237 (O_3237,N_29395,N_29290);
xor UO_3238 (O_3238,N_29691,N_28890);
and UO_3239 (O_3239,N_29108,N_29731);
xnor UO_3240 (O_3240,N_29855,N_29654);
or UO_3241 (O_3241,N_29116,N_28945);
xor UO_3242 (O_3242,N_28993,N_28837);
or UO_3243 (O_3243,N_28806,N_29266);
nor UO_3244 (O_3244,N_29404,N_29891);
and UO_3245 (O_3245,N_29264,N_29950);
xnor UO_3246 (O_3246,N_28938,N_29586);
nand UO_3247 (O_3247,N_29556,N_29785);
xnor UO_3248 (O_3248,N_29447,N_29229);
or UO_3249 (O_3249,N_29485,N_29099);
or UO_3250 (O_3250,N_29695,N_29383);
and UO_3251 (O_3251,N_29141,N_29262);
or UO_3252 (O_3252,N_29556,N_29807);
and UO_3253 (O_3253,N_29069,N_29818);
or UO_3254 (O_3254,N_29920,N_29762);
nor UO_3255 (O_3255,N_29620,N_29636);
xnor UO_3256 (O_3256,N_29151,N_29241);
xnor UO_3257 (O_3257,N_29150,N_29597);
or UO_3258 (O_3258,N_28982,N_29799);
nor UO_3259 (O_3259,N_29612,N_29114);
nand UO_3260 (O_3260,N_29953,N_29890);
nand UO_3261 (O_3261,N_29109,N_29547);
or UO_3262 (O_3262,N_29274,N_29593);
nor UO_3263 (O_3263,N_29516,N_29197);
and UO_3264 (O_3264,N_28810,N_29073);
xor UO_3265 (O_3265,N_29665,N_29012);
nor UO_3266 (O_3266,N_29344,N_29882);
or UO_3267 (O_3267,N_29660,N_29798);
and UO_3268 (O_3268,N_29465,N_29834);
nand UO_3269 (O_3269,N_29659,N_29964);
xor UO_3270 (O_3270,N_29188,N_29880);
and UO_3271 (O_3271,N_29058,N_29762);
xor UO_3272 (O_3272,N_29989,N_29436);
nor UO_3273 (O_3273,N_28901,N_29163);
xnor UO_3274 (O_3274,N_29817,N_29187);
and UO_3275 (O_3275,N_29881,N_29362);
or UO_3276 (O_3276,N_28912,N_29654);
or UO_3277 (O_3277,N_28994,N_29319);
nand UO_3278 (O_3278,N_29321,N_29847);
nor UO_3279 (O_3279,N_29787,N_29154);
nor UO_3280 (O_3280,N_28966,N_29433);
xor UO_3281 (O_3281,N_29825,N_29307);
xnor UO_3282 (O_3282,N_29056,N_29344);
nor UO_3283 (O_3283,N_29332,N_29594);
nand UO_3284 (O_3284,N_29553,N_29485);
and UO_3285 (O_3285,N_29462,N_29246);
nor UO_3286 (O_3286,N_29891,N_28980);
nand UO_3287 (O_3287,N_29464,N_29934);
and UO_3288 (O_3288,N_29871,N_29113);
nand UO_3289 (O_3289,N_29544,N_28951);
nand UO_3290 (O_3290,N_29486,N_28971);
nand UO_3291 (O_3291,N_29803,N_29059);
and UO_3292 (O_3292,N_29217,N_29339);
or UO_3293 (O_3293,N_29161,N_29967);
and UO_3294 (O_3294,N_29429,N_29727);
and UO_3295 (O_3295,N_28971,N_29713);
xnor UO_3296 (O_3296,N_28931,N_28993);
nor UO_3297 (O_3297,N_29150,N_29331);
or UO_3298 (O_3298,N_29820,N_29000);
nand UO_3299 (O_3299,N_29107,N_29392);
nand UO_3300 (O_3300,N_29130,N_29838);
and UO_3301 (O_3301,N_29158,N_29589);
xor UO_3302 (O_3302,N_29972,N_29267);
nand UO_3303 (O_3303,N_29909,N_28951);
nor UO_3304 (O_3304,N_29283,N_29804);
nand UO_3305 (O_3305,N_29159,N_29379);
or UO_3306 (O_3306,N_29307,N_29426);
and UO_3307 (O_3307,N_29408,N_29433);
nand UO_3308 (O_3308,N_28867,N_28897);
and UO_3309 (O_3309,N_29263,N_29676);
xnor UO_3310 (O_3310,N_29167,N_29244);
or UO_3311 (O_3311,N_29543,N_29266);
and UO_3312 (O_3312,N_29759,N_28879);
nand UO_3313 (O_3313,N_29511,N_29672);
or UO_3314 (O_3314,N_29868,N_28921);
nor UO_3315 (O_3315,N_29999,N_29199);
nor UO_3316 (O_3316,N_29715,N_29988);
nor UO_3317 (O_3317,N_29133,N_29961);
nand UO_3318 (O_3318,N_29780,N_29068);
and UO_3319 (O_3319,N_29615,N_29675);
nor UO_3320 (O_3320,N_28991,N_28985);
xor UO_3321 (O_3321,N_29708,N_29693);
xor UO_3322 (O_3322,N_28932,N_29986);
nor UO_3323 (O_3323,N_29500,N_29049);
nor UO_3324 (O_3324,N_29206,N_29618);
nor UO_3325 (O_3325,N_29219,N_29936);
and UO_3326 (O_3326,N_29250,N_28839);
xor UO_3327 (O_3327,N_29426,N_29218);
and UO_3328 (O_3328,N_29910,N_29270);
nor UO_3329 (O_3329,N_29570,N_29169);
nor UO_3330 (O_3330,N_28922,N_28966);
nand UO_3331 (O_3331,N_29989,N_29353);
and UO_3332 (O_3332,N_29914,N_29229);
xnor UO_3333 (O_3333,N_28843,N_29492);
nor UO_3334 (O_3334,N_29891,N_29625);
nand UO_3335 (O_3335,N_29359,N_29726);
xor UO_3336 (O_3336,N_28833,N_29950);
or UO_3337 (O_3337,N_29272,N_29921);
or UO_3338 (O_3338,N_29511,N_29295);
and UO_3339 (O_3339,N_29955,N_29425);
xor UO_3340 (O_3340,N_29464,N_29675);
and UO_3341 (O_3341,N_29454,N_29823);
nor UO_3342 (O_3342,N_29413,N_28976);
xnor UO_3343 (O_3343,N_29157,N_29282);
and UO_3344 (O_3344,N_29470,N_29199);
or UO_3345 (O_3345,N_28891,N_28933);
and UO_3346 (O_3346,N_28815,N_28950);
nand UO_3347 (O_3347,N_29247,N_29380);
nand UO_3348 (O_3348,N_28850,N_29946);
and UO_3349 (O_3349,N_28894,N_28974);
or UO_3350 (O_3350,N_29605,N_28846);
nor UO_3351 (O_3351,N_29494,N_29266);
or UO_3352 (O_3352,N_29219,N_28961);
or UO_3353 (O_3353,N_29820,N_29227);
nor UO_3354 (O_3354,N_29381,N_29385);
and UO_3355 (O_3355,N_29777,N_29735);
and UO_3356 (O_3356,N_29117,N_29105);
or UO_3357 (O_3357,N_29814,N_29879);
xnor UO_3358 (O_3358,N_29822,N_29481);
xor UO_3359 (O_3359,N_29410,N_29484);
or UO_3360 (O_3360,N_29029,N_29915);
nor UO_3361 (O_3361,N_29221,N_29999);
xnor UO_3362 (O_3362,N_28912,N_29582);
xnor UO_3363 (O_3363,N_29150,N_29309);
and UO_3364 (O_3364,N_29880,N_29050);
or UO_3365 (O_3365,N_29211,N_29307);
or UO_3366 (O_3366,N_29809,N_29637);
nand UO_3367 (O_3367,N_28837,N_29904);
xor UO_3368 (O_3368,N_29836,N_29452);
and UO_3369 (O_3369,N_28935,N_29902);
or UO_3370 (O_3370,N_29731,N_28815);
xnor UO_3371 (O_3371,N_29169,N_29409);
xnor UO_3372 (O_3372,N_29342,N_29165);
nand UO_3373 (O_3373,N_28813,N_29051);
nor UO_3374 (O_3374,N_28816,N_29921);
or UO_3375 (O_3375,N_29353,N_28917);
and UO_3376 (O_3376,N_29327,N_28981);
nand UO_3377 (O_3377,N_29577,N_28978);
and UO_3378 (O_3378,N_29903,N_29825);
nor UO_3379 (O_3379,N_28935,N_29495);
or UO_3380 (O_3380,N_28973,N_29121);
nand UO_3381 (O_3381,N_29207,N_29194);
nor UO_3382 (O_3382,N_29270,N_29226);
or UO_3383 (O_3383,N_29104,N_29125);
and UO_3384 (O_3384,N_29914,N_29336);
nand UO_3385 (O_3385,N_28903,N_29980);
nor UO_3386 (O_3386,N_29132,N_29741);
xor UO_3387 (O_3387,N_29830,N_28992);
nand UO_3388 (O_3388,N_29405,N_29014);
or UO_3389 (O_3389,N_29969,N_29572);
nand UO_3390 (O_3390,N_29027,N_29413);
and UO_3391 (O_3391,N_29874,N_28849);
xnor UO_3392 (O_3392,N_29356,N_29903);
and UO_3393 (O_3393,N_29837,N_29440);
nor UO_3394 (O_3394,N_28945,N_29688);
nand UO_3395 (O_3395,N_29951,N_29630);
xor UO_3396 (O_3396,N_28858,N_28928);
and UO_3397 (O_3397,N_29591,N_29162);
xor UO_3398 (O_3398,N_29620,N_29261);
nor UO_3399 (O_3399,N_29512,N_29364);
nor UO_3400 (O_3400,N_29443,N_29445);
or UO_3401 (O_3401,N_29580,N_29274);
nand UO_3402 (O_3402,N_29671,N_28863);
xor UO_3403 (O_3403,N_29964,N_29328);
nand UO_3404 (O_3404,N_29337,N_29479);
nor UO_3405 (O_3405,N_29809,N_28980);
or UO_3406 (O_3406,N_29527,N_29618);
xor UO_3407 (O_3407,N_29109,N_29149);
nor UO_3408 (O_3408,N_29821,N_29396);
xor UO_3409 (O_3409,N_29277,N_29005);
nand UO_3410 (O_3410,N_29532,N_29791);
or UO_3411 (O_3411,N_28919,N_29498);
nand UO_3412 (O_3412,N_29296,N_28958);
nor UO_3413 (O_3413,N_28840,N_29433);
xor UO_3414 (O_3414,N_29527,N_28924);
nand UO_3415 (O_3415,N_28977,N_29166);
and UO_3416 (O_3416,N_28936,N_28947);
and UO_3417 (O_3417,N_29606,N_29681);
nor UO_3418 (O_3418,N_29864,N_29589);
nor UO_3419 (O_3419,N_28936,N_29815);
or UO_3420 (O_3420,N_29832,N_29001);
nor UO_3421 (O_3421,N_29080,N_29322);
nand UO_3422 (O_3422,N_29692,N_29491);
nor UO_3423 (O_3423,N_29069,N_29941);
or UO_3424 (O_3424,N_29216,N_29208);
and UO_3425 (O_3425,N_28819,N_29257);
nor UO_3426 (O_3426,N_28887,N_29083);
nor UO_3427 (O_3427,N_29985,N_29668);
and UO_3428 (O_3428,N_29011,N_29312);
and UO_3429 (O_3429,N_29695,N_29304);
nor UO_3430 (O_3430,N_28969,N_29557);
or UO_3431 (O_3431,N_29523,N_29433);
nor UO_3432 (O_3432,N_29663,N_29048);
xor UO_3433 (O_3433,N_29607,N_29124);
nand UO_3434 (O_3434,N_28983,N_29075);
or UO_3435 (O_3435,N_29652,N_28841);
nand UO_3436 (O_3436,N_29471,N_29058);
or UO_3437 (O_3437,N_29391,N_29445);
and UO_3438 (O_3438,N_29766,N_29543);
nand UO_3439 (O_3439,N_29297,N_29924);
nand UO_3440 (O_3440,N_29069,N_28958);
nand UO_3441 (O_3441,N_28819,N_29910);
xnor UO_3442 (O_3442,N_28980,N_28905);
and UO_3443 (O_3443,N_29900,N_29812);
nor UO_3444 (O_3444,N_29884,N_29312);
nand UO_3445 (O_3445,N_28834,N_29072);
nor UO_3446 (O_3446,N_29552,N_28894);
or UO_3447 (O_3447,N_29818,N_29017);
and UO_3448 (O_3448,N_29803,N_29023);
nand UO_3449 (O_3449,N_29817,N_29641);
nor UO_3450 (O_3450,N_29875,N_29246);
or UO_3451 (O_3451,N_29230,N_29760);
and UO_3452 (O_3452,N_29115,N_28873);
or UO_3453 (O_3453,N_29129,N_28979);
nand UO_3454 (O_3454,N_29962,N_29015);
and UO_3455 (O_3455,N_28904,N_28919);
nand UO_3456 (O_3456,N_29570,N_29574);
or UO_3457 (O_3457,N_29224,N_29612);
or UO_3458 (O_3458,N_29569,N_29015);
nor UO_3459 (O_3459,N_29576,N_29923);
nor UO_3460 (O_3460,N_28930,N_29639);
and UO_3461 (O_3461,N_29604,N_29244);
and UO_3462 (O_3462,N_29425,N_29328);
and UO_3463 (O_3463,N_29154,N_29006);
or UO_3464 (O_3464,N_29120,N_29955);
or UO_3465 (O_3465,N_29213,N_29162);
nor UO_3466 (O_3466,N_29611,N_29401);
and UO_3467 (O_3467,N_29914,N_29314);
nand UO_3468 (O_3468,N_29719,N_29168);
or UO_3469 (O_3469,N_29950,N_29229);
nand UO_3470 (O_3470,N_29925,N_29916);
nand UO_3471 (O_3471,N_29766,N_28814);
and UO_3472 (O_3472,N_29014,N_29790);
or UO_3473 (O_3473,N_29987,N_29774);
nand UO_3474 (O_3474,N_29029,N_29687);
and UO_3475 (O_3475,N_28940,N_29345);
nand UO_3476 (O_3476,N_29692,N_28983);
and UO_3477 (O_3477,N_29360,N_29299);
nand UO_3478 (O_3478,N_29009,N_28879);
nor UO_3479 (O_3479,N_29293,N_29242);
xnor UO_3480 (O_3480,N_29239,N_29226);
nor UO_3481 (O_3481,N_29286,N_29172);
nor UO_3482 (O_3482,N_28838,N_28803);
or UO_3483 (O_3483,N_29894,N_28923);
and UO_3484 (O_3484,N_28853,N_29488);
and UO_3485 (O_3485,N_29030,N_29709);
or UO_3486 (O_3486,N_29770,N_29139);
nand UO_3487 (O_3487,N_29420,N_29045);
nand UO_3488 (O_3488,N_29148,N_29737);
xnor UO_3489 (O_3489,N_29227,N_29507);
or UO_3490 (O_3490,N_28842,N_29141);
xor UO_3491 (O_3491,N_29083,N_29136);
nor UO_3492 (O_3492,N_28869,N_28964);
nand UO_3493 (O_3493,N_29352,N_29031);
and UO_3494 (O_3494,N_29903,N_29327);
nor UO_3495 (O_3495,N_29281,N_29236);
and UO_3496 (O_3496,N_29874,N_29300);
nor UO_3497 (O_3497,N_29213,N_29031);
or UO_3498 (O_3498,N_29191,N_29040);
xor UO_3499 (O_3499,N_29809,N_29501);
endmodule