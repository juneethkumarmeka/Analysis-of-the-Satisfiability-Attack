module basic_500_3000_500_30_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_305,In_101);
or U1 (N_1,In_37,In_253);
and U2 (N_2,In_93,In_42);
or U3 (N_3,In_179,In_445);
nor U4 (N_4,In_23,In_149);
and U5 (N_5,In_489,In_429);
or U6 (N_6,In_237,In_312);
nor U7 (N_7,In_106,In_108);
nand U8 (N_8,In_21,In_89);
nand U9 (N_9,In_60,In_224);
and U10 (N_10,In_100,In_152);
nor U11 (N_11,In_255,In_47);
nor U12 (N_12,In_170,In_372);
nor U13 (N_13,In_308,In_168);
nor U14 (N_14,In_70,In_52);
nand U15 (N_15,In_370,In_322);
and U16 (N_16,In_307,In_7);
nor U17 (N_17,In_26,In_344);
or U18 (N_18,In_455,In_323);
nor U19 (N_19,In_466,In_135);
or U20 (N_20,In_490,In_86);
nand U21 (N_21,In_206,In_300);
nor U22 (N_22,In_494,In_109);
nand U23 (N_23,In_239,In_274);
or U24 (N_24,In_431,In_363);
xnor U25 (N_25,In_159,In_178);
or U26 (N_26,In_329,In_243);
and U27 (N_27,In_250,In_166);
or U28 (N_28,In_407,In_142);
nand U29 (N_29,In_81,In_53);
and U30 (N_30,In_215,In_20);
or U31 (N_31,In_43,In_175);
nand U32 (N_32,In_285,In_383);
and U33 (N_33,In_311,In_336);
nand U34 (N_34,In_485,In_90);
nor U35 (N_35,In_483,In_136);
or U36 (N_36,In_121,In_496);
nor U37 (N_37,In_48,In_337);
nor U38 (N_38,In_476,In_280);
and U39 (N_39,In_141,In_203);
and U40 (N_40,In_402,In_145);
or U41 (N_41,In_127,In_498);
and U42 (N_42,In_155,In_111);
and U43 (N_43,In_260,In_439);
nor U44 (N_44,In_408,In_479);
or U45 (N_45,In_176,In_5);
and U46 (N_46,In_392,In_193);
nor U47 (N_47,In_313,In_265);
nand U48 (N_48,In_218,In_341);
or U49 (N_49,In_73,In_33);
or U50 (N_50,In_474,In_443);
nand U51 (N_51,In_269,In_83);
or U52 (N_52,In_63,In_471);
and U53 (N_53,In_6,In_414);
or U54 (N_54,In_143,In_67);
or U55 (N_55,In_219,In_389);
nand U56 (N_56,In_378,In_434);
or U57 (N_57,In_197,In_477);
or U58 (N_58,In_2,In_314);
nor U59 (N_59,In_140,In_16);
nand U60 (N_60,In_281,In_126);
and U61 (N_61,In_147,In_78);
nand U62 (N_62,In_457,In_440);
or U63 (N_63,In_267,In_339);
and U64 (N_64,In_3,In_433);
nand U65 (N_65,In_475,In_430);
and U66 (N_66,In_229,In_347);
and U67 (N_67,In_411,In_317);
nand U68 (N_68,In_484,In_97);
or U69 (N_69,In_57,In_58);
nor U70 (N_70,In_211,In_491);
and U71 (N_71,In_130,In_299);
nand U72 (N_72,In_169,In_161);
nand U73 (N_73,In_92,In_330);
nand U74 (N_74,In_398,In_444);
nor U75 (N_75,In_117,In_374);
and U76 (N_76,In_74,In_188);
nor U77 (N_77,In_275,In_461);
and U78 (N_78,In_227,In_184);
nand U79 (N_79,In_55,In_25);
nor U80 (N_80,In_397,In_45);
nand U81 (N_81,In_316,In_172);
and U82 (N_82,In_278,In_12);
nand U83 (N_83,In_379,In_348);
and U84 (N_84,In_64,In_54);
or U85 (N_85,In_424,In_410);
nand U86 (N_86,In_72,In_115);
or U87 (N_87,In_191,In_375);
nor U88 (N_88,In_364,In_38);
and U89 (N_89,In_234,In_156);
nand U90 (N_90,In_85,In_387);
nor U91 (N_91,In_283,In_61);
nand U92 (N_92,In_456,In_263);
nor U93 (N_93,In_277,In_107);
nand U94 (N_94,In_76,In_436);
nor U95 (N_95,In_137,In_264);
and U96 (N_96,In_31,In_282);
nor U97 (N_97,In_332,In_244);
or U98 (N_98,In_196,In_200);
or U99 (N_99,In_353,In_349);
nor U100 (N_100,N_10,In_241);
and U101 (N_101,In_469,In_226);
nand U102 (N_102,In_376,In_238);
and U103 (N_103,In_257,In_315);
and U104 (N_104,In_301,In_134);
and U105 (N_105,In_105,In_185);
nand U106 (N_106,In_19,In_272);
or U107 (N_107,In_318,In_470);
and U108 (N_108,N_55,In_354);
nor U109 (N_109,In_463,In_15);
nand U110 (N_110,In_266,In_113);
nand U111 (N_111,In_325,In_319);
nor U112 (N_112,In_286,N_90);
and U113 (N_113,In_460,In_151);
or U114 (N_114,In_28,N_17);
nand U115 (N_115,In_119,In_157);
nand U116 (N_116,In_17,In_98);
or U117 (N_117,In_298,In_459);
and U118 (N_118,In_190,In_393);
nor U119 (N_119,In_452,N_65);
nand U120 (N_120,In_276,In_465);
or U121 (N_121,In_232,In_34);
and U122 (N_122,In_421,In_396);
or U123 (N_123,In_360,In_345);
or U124 (N_124,In_331,In_386);
or U125 (N_125,N_0,N_41);
and U126 (N_126,In_291,In_369);
xor U127 (N_127,N_7,In_79);
and U128 (N_128,In_390,In_8);
xor U129 (N_129,In_453,In_437);
nor U130 (N_130,N_19,In_419);
nand U131 (N_131,In_295,N_73);
nand U132 (N_132,In_423,In_468);
and U133 (N_133,In_118,N_95);
nand U134 (N_134,In_371,In_24);
xor U135 (N_135,In_36,In_217);
or U136 (N_136,In_56,In_230);
and U137 (N_137,In_65,In_368);
xnor U138 (N_138,N_33,N_68);
nand U139 (N_139,In_287,In_395);
and U140 (N_140,In_94,In_198);
or U141 (N_141,N_75,In_258);
nor U142 (N_142,In_488,In_9);
nand U143 (N_143,In_384,In_352);
nand U144 (N_144,In_138,In_248);
nand U145 (N_145,In_195,In_133);
nand U146 (N_146,In_228,In_448);
or U147 (N_147,In_449,N_83);
nor U148 (N_148,N_58,In_381);
nor U149 (N_149,In_139,N_20);
nor U150 (N_150,N_67,N_1);
or U151 (N_151,N_93,In_435);
nand U152 (N_152,N_14,In_427);
nand U153 (N_153,In_343,In_125);
and U154 (N_154,In_77,In_252);
and U155 (N_155,In_205,In_382);
or U156 (N_156,In_333,In_367);
or U157 (N_157,In_290,In_486);
and U158 (N_158,In_304,In_324);
nor U159 (N_159,In_404,In_405);
and U160 (N_160,N_94,In_44);
nand U161 (N_161,In_123,In_357);
and U162 (N_162,N_26,In_207);
or U163 (N_163,N_74,In_204);
nor U164 (N_164,In_245,In_428);
or U165 (N_165,In_365,In_432);
and U166 (N_166,N_47,N_78);
or U167 (N_167,In_189,N_13);
or U168 (N_168,In_46,In_165);
nand U169 (N_169,In_181,In_29);
nand U170 (N_170,N_80,In_99);
and U171 (N_171,In_492,In_262);
nor U172 (N_172,In_413,N_32);
and U173 (N_173,N_54,In_62);
and U174 (N_174,In_210,In_450);
and U175 (N_175,N_43,In_209);
or U176 (N_176,In_467,In_254);
and U177 (N_177,In_454,N_31);
or U178 (N_178,In_236,In_201);
nor U179 (N_179,In_293,N_69);
nand U180 (N_180,In_11,In_359);
nor U181 (N_181,In_103,In_14);
and U182 (N_182,In_270,N_4);
and U183 (N_183,In_481,N_76);
or U184 (N_184,In_220,In_388);
nor U185 (N_185,N_15,In_361);
nand U186 (N_186,N_23,In_199);
and U187 (N_187,In_32,In_223);
and U188 (N_188,In_75,In_403);
nand U189 (N_189,In_59,In_122);
nor U190 (N_190,In_242,In_473);
or U191 (N_191,N_61,N_63);
nor U192 (N_192,In_40,In_4);
nor U193 (N_193,In_124,In_292);
and U194 (N_194,N_40,In_91);
or U195 (N_195,In_240,In_114);
and U196 (N_196,In_183,In_116);
or U197 (N_197,N_79,In_321);
nor U198 (N_198,N_21,In_446);
nand U199 (N_199,In_87,In_102);
nor U200 (N_200,N_108,N_141);
or U201 (N_201,In_163,In_297);
nand U202 (N_202,N_86,N_99);
nor U203 (N_203,In_380,N_45);
nor U204 (N_204,N_137,N_113);
nor U205 (N_205,N_82,In_148);
or U206 (N_206,N_148,N_120);
or U207 (N_207,In_84,In_186);
nor U208 (N_208,N_138,In_212);
or U209 (N_209,In_146,N_174);
and U210 (N_210,In_328,N_64);
nand U211 (N_211,N_139,N_147);
nand U212 (N_212,In_373,N_133);
and U213 (N_213,N_38,N_168);
or U214 (N_214,In_49,In_409);
and U215 (N_215,In_51,In_50);
and U216 (N_216,N_188,In_271);
or U217 (N_217,N_117,In_458);
nand U218 (N_218,N_144,N_185);
nor U219 (N_219,In_326,In_164);
nor U220 (N_220,N_195,N_12);
or U221 (N_221,In_462,In_216);
or U222 (N_222,In_132,In_194);
and U223 (N_223,N_34,In_487);
nand U224 (N_224,N_158,In_400);
nor U225 (N_225,In_222,N_152);
or U226 (N_226,In_131,In_96);
and U227 (N_227,In_171,In_82);
nand U228 (N_228,In_377,N_132);
nor U229 (N_229,In_30,N_126);
or U230 (N_230,In_422,In_327);
or U231 (N_231,In_1,N_59);
or U232 (N_232,In_451,In_150);
nand U233 (N_233,N_198,N_53);
nand U234 (N_234,In_472,N_39);
or U235 (N_235,In_391,N_107);
or U236 (N_236,N_171,N_170);
nor U237 (N_237,N_44,In_0);
or U238 (N_238,N_2,In_310);
nand U239 (N_239,N_105,N_193);
or U240 (N_240,In_249,N_153);
nand U241 (N_241,In_426,N_123);
nand U242 (N_242,In_95,In_66);
and U243 (N_243,In_22,In_13);
and U244 (N_244,N_51,N_84);
and U245 (N_245,N_182,N_192);
or U246 (N_246,N_154,In_279);
nand U247 (N_247,N_197,In_213);
nor U248 (N_248,N_101,N_30);
and U249 (N_249,N_110,In_385);
nor U250 (N_250,In_41,N_96);
nor U251 (N_251,In_182,In_366);
nand U252 (N_252,N_6,N_163);
or U253 (N_253,N_114,N_111);
nand U254 (N_254,In_88,N_196);
nor U255 (N_255,In_18,In_480);
or U256 (N_256,In_202,In_173);
or U257 (N_257,In_192,N_89);
nand U258 (N_258,N_130,In_350);
nand U259 (N_259,N_166,In_356);
nor U260 (N_260,N_91,In_251);
or U261 (N_261,N_155,N_106);
nor U262 (N_262,In_464,In_362);
and U263 (N_263,In_417,N_134);
and U264 (N_264,N_183,N_177);
nand U265 (N_265,In_235,In_415);
nor U266 (N_266,In_303,N_131);
nand U267 (N_267,N_149,N_62);
nor U268 (N_268,N_27,N_194);
or U269 (N_269,N_159,N_36);
and U270 (N_270,In_162,In_10);
nand U271 (N_271,In_225,In_129);
nand U272 (N_272,In_334,N_24);
nor U273 (N_273,In_289,N_49);
or U274 (N_274,N_189,N_127);
and U275 (N_275,N_140,In_221);
nor U276 (N_276,N_52,N_16);
or U277 (N_277,In_112,N_191);
or U278 (N_278,In_478,N_146);
and U279 (N_279,In_358,N_28);
nor U280 (N_280,N_187,In_208);
nor U281 (N_281,N_181,N_167);
or U282 (N_282,N_135,In_154);
nor U283 (N_283,N_77,N_97);
nor U284 (N_284,In_153,In_288);
and U285 (N_285,In_68,N_102);
nand U286 (N_286,In_144,N_164);
and U287 (N_287,In_268,N_72);
nor U288 (N_288,In_261,In_306);
or U289 (N_289,In_120,In_187);
nand U290 (N_290,In_273,N_180);
and U291 (N_291,N_18,In_335);
or U292 (N_292,In_401,N_87);
or U293 (N_293,N_85,In_497);
or U294 (N_294,In_499,N_116);
or U295 (N_295,N_92,In_214);
and U296 (N_296,N_118,In_128);
and U297 (N_297,In_351,N_173);
or U298 (N_298,N_156,N_124);
nand U299 (N_299,In_259,N_29);
and U300 (N_300,N_219,N_224);
and U301 (N_301,N_288,N_202);
and U302 (N_302,N_281,N_208);
xnor U303 (N_303,N_279,N_243);
or U304 (N_304,In_110,In_416);
nor U305 (N_305,N_257,N_60);
and U306 (N_306,N_25,N_271);
and U307 (N_307,N_241,N_203);
nand U308 (N_308,N_88,In_256);
and U309 (N_309,N_254,N_5);
or U310 (N_310,N_273,N_244);
nand U311 (N_311,N_276,N_172);
or U312 (N_312,N_213,In_294);
nand U313 (N_313,N_220,In_302);
or U314 (N_314,N_184,N_176);
and U315 (N_315,In_27,N_50);
nor U316 (N_316,N_245,N_264);
or U317 (N_317,N_251,N_119);
nor U318 (N_318,N_157,N_81);
nand U319 (N_319,N_11,In_447);
and U320 (N_320,In_418,N_233);
nor U321 (N_321,N_42,N_272);
or U322 (N_322,In_284,N_269);
nor U323 (N_323,N_66,N_121);
and U324 (N_324,N_125,N_258);
and U325 (N_325,N_296,N_216);
nor U326 (N_326,N_206,N_293);
and U327 (N_327,N_290,N_299);
or U328 (N_328,N_250,In_340);
and U329 (N_329,N_275,N_265);
or U330 (N_330,N_205,N_283);
or U331 (N_331,N_270,N_98);
nor U332 (N_332,N_295,N_160);
nand U333 (N_333,In_231,N_35);
and U334 (N_334,N_225,N_129);
or U335 (N_335,N_222,N_260);
nand U336 (N_336,N_246,N_249);
nor U337 (N_337,N_223,In_441);
and U338 (N_338,N_37,N_103);
and U339 (N_339,N_8,N_9);
nor U340 (N_340,N_242,N_256);
nor U341 (N_341,N_112,N_143);
or U342 (N_342,In_355,N_56);
or U343 (N_343,N_214,N_136);
nor U344 (N_344,N_278,In_158);
nor U345 (N_345,N_268,N_70);
nand U346 (N_346,N_298,N_235);
nand U347 (N_347,N_240,In_35);
and U348 (N_348,N_266,N_255);
nand U349 (N_349,N_294,N_234);
and U350 (N_350,N_46,N_178);
or U351 (N_351,In_442,In_438);
nor U352 (N_352,N_252,N_277);
nor U353 (N_353,N_142,N_217);
nand U354 (N_354,In_39,N_229);
nand U355 (N_355,In_180,N_238);
and U356 (N_356,N_232,N_228);
and U357 (N_357,N_227,N_151);
nor U358 (N_358,In_104,N_212);
nand U359 (N_359,N_253,N_261);
nand U360 (N_360,In_495,N_226);
nor U361 (N_361,In_296,N_169);
or U362 (N_362,In_246,N_292);
or U363 (N_363,N_71,N_282);
nand U364 (N_364,N_179,N_218);
nand U365 (N_365,In_399,N_100);
nand U366 (N_366,N_211,N_201);
or U367 (N_367,In_160,N_150);
or U368 (N_368,N_48,In_394);
nor U369 (N_369,N_109,In_69);
or U370 (N_370,N_280,N_161);
or U371 (N_371,In_482,N_287);
nand U372 (N_372,N_165,In_177);
or U373 (N_373,In_309,N_162);
xor U374 (N_374,N_204,N_239);
or U375 (N_375,In_233,In_338);
or U376 (N_376,N_284,N_207);
and U377 (N_377,In_420,N_262);
nor U378 (N_378,N_230,In_425);
nand U379 (N_379,N_297,N_128);
or U380 (N_380,In_174,N_291);
and U381 (N_381,In_247,N_22);
nand U382 (N_382,N_200,N_248);
nand U383 (N_383,N_286,N_221);
or U384 (N_384,N_145,N_263);
nor U385 (N_385,In_320,In_346);
nand U386 (N_386,In_406,N_285);
and U387 (N_387,N_3,N_289);
nand U388 (N_388,In_71,N_267);
or U389 (N_389,N_247,In_167);
nor U390 (N_390,N_57,N_231);
and U391 (N_391,N_186,N_215);
nand U392 (N_392,N_199,In_412);
and U393 (N_393,N_209,In_80);
and U394 (N_394,N_236,In_493);
and U395 (N_395,N_122,N_274);
nor U396 (N_396,N_104,N_175);
nor U397 (N_397,In_342,N_210);
nor U398 (N_398,N_190,N_115);
nand U399 (N_399,N_259,N_237);
and U400 (N_400,N_396,N_347);
nand U401 (N_401,N_377,N_310);
nor U402 (N_402,N_337,N_336);
nor U403 (N_403,N_361,N_354);
nand U404 (N_404,N_344,N_366);
or U405 (N_405,N_340,N_376);
nand U406 (N_406,N_387,N_302);
or U407 (N_407,N_348,N_352);
nand U408 (N_408,N_343,N_317);
nand U409 (N_409,N_324,N_304);
and U410 (N_410,N_351,N_385);
nand U411 (N_411,N_319,N_322);
or U412 (N_412,N_355,N_350);
nand U413 (N_413,N_327,N_346);
or U414 (N_414,N_335,N_390);
or U415 (N_415,N_307,N_331);
nand U416 (N_416,N_378,N_392);
nor U417 (N_417,N_316,N_358);
and U418 (N_418,N_362,N_349);
nand U419 (N_419,N_332,N_395);
or U420 (N_420,N_370,N_393);
xnor U421 (N_421,N_338,N_359);
and U422 (N_422,N_380,N_368);
or U423 (N_423,N_364,N_308);
or U424 (N_424,N_315,N_379);
nand U425 (N_425,N_334,N_356);
nor U426 (N_426,N_373,N_345);
and U427 (N_427,N_329,N_367);
or U428 (N_428,N_305,N_328);
and U429 (N_429,N_325,N_333);
nor U430 (N_430,N_357,N_300);
or U431 (N_431,N_381,N_386);
nand U432 (N_432,N_375,N_369);
and U433 (N_433,N_342,N_321);
nor U434 (N_434,N_323,N_399);
xnor U435 (N_435,N_397,N_301);
and U436 (N_436,N_318,N_326);
and U437 (N_437,N_313,N_314);
nor U438 (N_438,N_374,N_306);
nand U439 (N_439,N_341,N_303);
and U440 (N_440,N_388,N_389);
nor U441 (N_441,N_384,N_372);
and U442 (N_442,N_391,N_383);
and U443 (N_443,N_365,N_398);
nor U444 (N_444,N_320,N_360);
xor U445 (N_445,N_363,N_309);
and U446 (N_446,N_394,N_312);
and U447 (N_447,N_353,N_311);
nor U448 (N_448,N_371,N_382);
nor U449 (N_449,N_330,N_339);
or U450 (N_450,N_374,N_394);
or U451 (N_451,N_350,N_395);
or U452 (N_452,N_385,N_334);
and U453 (N_453,N_376,N_368);
or U454 (N_454,N_386,N_371);
nor U455 (N_455,N_331,N_373);
and U456 (N_456,N_354,N_344);
or U457 (N_457,N_356,N_347);
or U458 (N_458,N_323,N_321);
or U459 (N_459,N_358,N_332);
and U460 (N_460,N_335,N_318);
or U461 (N_461,N_362,N_354);
and U462 (N_462,N_373,N_347);
or U463 (N_463,N_351,N_360);
and U464 (N_464,N_392,N_386);
nand U465 (N_465,N_304,N_340);
nor U466 (N_466,N_342,N_362);
or U467 (N_467,N_347,N_362);
or U468 (N_468,N_378,N_385);
nor U469 (N_469,N_392,N_325);
and U470 (N_470,N_327,N_369);
and U471 (N_471,N_389,N_374);
nand U472 (N_472,N_311,N_382);
nor U473 (N_473,N_376,N_377);
nor U474 (N_474,N_341,N_354);
or U475 (N_475,N_312,N_377);
nand U476 (N_476,N_373,N_362);
nor U477 (N_477,N_336,N_329);
nand U478 (N_478,N_360,N_368);
nor U479 (N_479,N_320,N_310);
nor U480 (N_480,N_396,N_339);
nor U481 (N_481,N_362,N_328);
nand U482 (N_482,N_321,N_358);
nand U483 (N_483,N_384,N_367);
nor U484 (N_484,N_305,N_369);
and U485 (N_485,N_387,N_373);
or U486 (N_486,N_335,N_349);
nor U487 (N_487,N_370,N_341);
and U488 (N_488,N_342,N_370);
and U489 (N_489,N_303,N_396);
nor U490 (N_490,N_315,N_316);
nor U491 (N_491,N_341,N_348);
or U492 (N_492,N_347,N_328);
nand U493 (N_493,N_392,N_345);
nor U494 (N_494,N_374,N_357);
nor U495 (N_495,N_370,N_344);
and U496 (N_496,N_342,N_316);
nor U497 (N_497,N_327,N_362);
or U498 (N_498,N_347,N_366);
nand U499 (N_499,N_345,N_321);
and U500 (N_500,N_427,N_419);
nand U501 (N_501,N_448,N_493);
nand U502 (N_502,N_449,N_423);
and U503 (N_503,N_435,N_457);
nand U504 (N_504,N_488,N_439);
nand U505 (N_505,N_472,N_462);
and U506 (N_506,N_407,N_422);
nand U507 (N_507,N_445,N_441);
nor U508 (N_508,N_492,N_494);
and U509 (N_509,N_402,N_425);
nand U510 (N_510,N_418,N_468);
nand U511 (N_511,N_491,N_459);
nor U512 (N_512,N_434,N_466);
and U513 (N_513,N_489,N_496);
and U514 (N_514,N_403,N_481);
or U515 (N_515,N_490,N_442);
or U516 (N_516,N_447,N_497);
or U517 (N_517,N_461,N_443);
or U518 (N_518,N_474,N_478);
nand U519 (N_519,N_438,N_485);
or U520 (N_520,N_495,N_436);
or U521 (N_521,N_486,N_456);
xor U522 (N_522,N_483,N_460);
nand U523 (N_523,N_475,N_455);
nor U524 (N_524,N_452,N_430);
and U525 (N_525,N_404,N_465);
or U526 (N_526,N_499,N_476);
or U527 (N_527,N_415,N_498);
or U528 (N_528,N_487,N_482);
and U529 (N_529,N_437,N_429);
or U530 (N_530,N_433,N_405);
nor U531 (N_531,N_484,N_479);
and U532 (N_532,N_408,N_432);
nand U533 (N_533,N_470,N_469);
nor U534 (N_534,N_428,N_473);
and U535 (N_535,N_454,N_471);
and U536 (N_536,N_414,N_421);
and U537 (N_537,N_440,N_417);
or U538 (N_538,N_412,N_446);
and U539 (N_539,N_453,N_411);
nand U540 (N_540,N_450,N_431);
nor U541 (N_541,N_416,N_409);
and U542 (N_542,N_413,N_477);
nor U543 (N_543,N_463,N_451);
nor U544 (N_544,N_401,N_444);
nand U545 (N_545,N_464,N_458);
nor U546 (N_546,N_420,N_480);
nand U547 (N_547,N_424,N_400);
or U548 (N_548,N_406,N_410);
and U549 (N_549,N_426,N_467);
or U550 (N_550,N_492,N_452);
nand U551 (N_551,N_414,N_468);
nand U552 (N_552,N_443,N_495);
nand U553 (N_553,N_475,N_466);
nor U554 (N_554,N_404,N_453);
or U555 (N_555,N_483,N_416);
xnor U556 (N_556,N_481,N_422);
nor U557 (N_557,N_445,N_466);
nand U558 (N_558,N_414,N_498);
nor U559 (N_559,N_443,N_414);
and U560 (N_560,N_417,N_434);
nor U561 (N_561,N_463,N_404);
or U562 (N_562,N_439,N_490);
and U563 (N_563,N_455,N_480);
nor U564 (N_564,N_474,N_457);
and U565 (N_565,N_441,N_483);
and U566 (N_566,N_489,N_483);
or U567 (N_567,N_475,N_439);
nor U568 (N_568,N_421,N_493);
and U569 (N_569,N_444,N_438);
or U570 (N_570,N_443,N_497);
nand U571 (N_571,N_430,N_486);
or U572 (N_572,N_452,N_497);
nor U573 (N_573,N_464,N_429);
or U574 (N_574,N_404,N_412);
or U575 (N_575,N_463,N_447);
and U576 (N_576,N_485,N_495);
nor U577 (N_577,N_445,N_453);
and U578 (N_578,N_428,N_436);
nor U579 (N_579,N_465,N_495);
nor U580 (N_580,N_437,N_456);
and U581 (N_581,N_426,N_429);
nand U582 (N_582,N_472,N_451);
nor U583 (N_583,N_490,N_466);
or U584 (N_584,N_414,N_491);
nor U585 (N_585,N_405,N_460);
nor U586 (N_586,N_490,N_410);
or U587 (N_587,N_463,N_411);
nor U588 (N_588,N_416,N_455);
and U589 (N_589,N_456,N_416);
nand U590 (N_590,N_428,N_414);
or U591 (N_591,N_473,N_416);
and U592 (N_592,N_451,N_433);
and U593 (N_593,N_464,N_497);
nand U594 (N_594,N_440,N_478);
nor U595 (N_595,N_450,N_410);
nand U596 (N_596,N_456,N_414);
nor U597 (N_597,N_417,N_499);
and U598 (N_598,N_471,N_414);
nor U599 (N_599,N_464,N_481);
or U600 (N_600,N_580,N_595);
nor U601 (N_601,N_558,N_510);
nor U602 (N_602,N_592,N_502);
or U603 (N_603,N_559,N_587);
or U604 (N_604,N_509,N_521);
nor U605 (N_605,N_537,N_599);
or U606 (N_606,N_542,N_544);
nor U607 (N_607,N_564,N_515);
or U608 (N_608,N_547,N_543);
and U609 (N_609,N_565,N_570);
or U610 (N_610,N_517,N_532);
or U611 (N_611,N_551,N_503);
and U612 (N_612,N_540,N_549);
nand U613 (N_613,N_562,N_577);
or U614 (N_614,N_561,N_576);
or U615 (N_615,N_512,N_504);
nand U616 (N_616,N_584,N_505);
nor U617 (N_617,N_591,N_583);
or U618 (N_618,N_585,N_508);
nand U619 (N_619,N_578,N_552);
and U620 (N_620,N_563,N_568);
nand U621 (N_621,N_569,N_524);
or U622 (N_622,N_574,N_523);
or U623 (N_623,N_556,N_534);
nor U624 (N_624,N_522,N_528);
and U625 (N_625,N_560,N_546);
nor U626 (N_626,N_582,N_571);
and U627 (N_627,N_518,N_527);
nor U628 (N_628,N_554,N_575);
nor U629 (N_629,N_557,N_525);
or U630 (N_630,N_597,N_593);
nor U631 (N_631,N_586,N_553);
or U632 (N_632,N_516,N_520);
nor U633 (N_633,N_513,N_514);
and U634 (N_634,N_539,N_526);
nor U635 (N_635,N_548,N_579);
or U636 (N_636,N_567,N_566);
nor U637 (N_637,N_535,N_550);
nor U638 (N_638,N_530,N_531);
nand U639 (N_639,N_500,N_533);
and U640 (N_640,N_590,N_511);
and U641 (N_641,N_506,N_545);
nand U642 (N_642,N_589,N_598);
or U643 (N_643,N_529,N_588);
nand U644 (N_644,N_541,N_596);
nor U645 (N_645,N_572,N_555);
nor U646 (N_646,N_501,N_573);
nor U647 (N_647,N_536,N_538);
and U648 (N_648,N_507,N_581);
nand U649 (N_649,N_519,N_594);
nor U650 (N_650,N_511,N_558);
nand U651 (N_651,N_583,N_544);
nor U652 (N_652,N_561,N_570);
and U653 (N_653,N_534,N_531);
nand U654 (N_654,N_502,N_575);
nor U655 (N_655,N_568,N_544);
or U656 (N_656,N_502,N_590);
nor U657 (N_657,N_562,N_555);
or U658 (N_658,N_592,N_522);
and U659 (N_659,N_530,N_511);
or U660 (N_660,N_520,N_519);
nor U661 (N_661,N_589,N_501);
nand U662 (N_662,N_521,N_574);
nand U663 (N_663,N_515,N_531);
or U664 (N_664,N_584,N_568);
nand U665 (N_665,N_585,N_588);
nor U666 (N_666,N_576,N_588);
nor U667 (N_667,N_506,N_591);
and U668 (N_668,N_587,N_595);
nor U669 (N_669,N_572,N_584);
nor U670 (N_670,N_583,N_566);
nor U671 (N_671,N_597,N_595);
and U672 (N_672,N_589,N_554);
or U673 (N_673,N_516,N_558);
and U674 (N_674,N_544,N_564);
and U675 (N_675,N_504,N_534);
nand U676 (N_676,N_509,N_548);
and U677 (N_677,N_588,N_501);
nor U678 (N_678,N_505,N_553);
or U679 (N_679,N_544,N_548);
and U680 (N_680,N_522,N_570);
and U681 (N_681,N_523,N_573);
nand U682 (N_682,N_505,N_570);
nand U683 (N_683,N_547,N_546);
or U684 (N_684,N_580,N_517);
and U685 (N_685,N_595,N_534);
or U686 (N_686,N_521,N_507);
nand U687 (N_687,N_575,N_560);
nor U688 (N_688,N_531,N_552);
nand U689 (N_689,N_551,N_560);
or U690 (N_690,N_597,N_534);
nand U691 (N_691,N_547,N_588);
or U692 (N_692,N_573,N_503);
nand U693 (N_693,N_540,N_537);
nor U694 (N_694,N_521,N_500);
nor U695 (N_695,N_544,N_508);
nor U696 (N_696,N_561,N_578);
and U697 (N_697,N_502,N_500);
or U698 (N_698,N_578,N_572);
or U699 (N_699,N_558,N_528);
and U700 (N_700,N_653,N_677);
nand U701 (N_701,N_603,N_684);
or U702 (N_702,N_664,N_636);
and U703 (N_703,N_692,N_620);
or U704 (N_704,N_663,N_674);
or U705 (N_705,N_654,N_633);
nand U706 (N_706,N_640,N_693);
and U707 (N_707,N_661,N_618);
nor U708 (N_708,N_662,N_670);
nand U709 (N_709,N_685,N_642);
and U710 (N_710,N_678,N_676);
or U711 (N_711,N_615,N_671);
nor U712 (N_712,N_611,N_600);
and U713 (N_713,N_699,N_672);
nor U714 (N_714,N_665,N_690);
and U715 (N_715,N_697,N_696);
or U716 (N_716,N_614,N_639);
nor U717 (N_717,N_624,N_617);
nor U718 (N_718,N_667,N_643);
nand U719 (N_719,N_608,N_622);
and U720 (N_720,N_646,N_632);
nand U721 (N_721,N_629,N_621);
nand U722 (N_722,N_645,N_648);
and U723 (N_723,N_698,N_656);
nor U724 (N_724,N_638,N_651);
nand U725 (N_725,N_605,N_637);
and U726 (N_726,N_679,N_655);
and U727 (N_727,N_631,N_659);
nand U728 (N_728,N_604,N_688);
nor U729 (N_729,N_669,N_602);
nor U730 (N_730,N_634,N_652);
nor U731 (N_731,N_613,N_657);
nor U732 (N_732,N_623,N_686);
and U733 (N_733,N_673,N_691);
nor U734 (N_734,N_658,N_650);
or U735 (N_735,N_612,N_689);
or U736 (N_736,N_627,N_635);
xnor U737 (N_737,N_630,N_681);
and U738 (N_738,N_606,N_625);
nor U739 (N_739,N_666,N_687);
nor U740 (N_740,N_668,N_601);
and U741 (N_741,N_610,N_626);
nor U742 (N_742,N_680,N_609);
xnor U743 (N_743,N_644,N_683);
and U744 (N_744,N_694,N_675);
nor U745 (N_745,N_647,N_616);
and U746 (N_746,N_619,N_695);
or U747 (N_747,N_607,N_628);
xor U748 (N_748,N_649,N_660);
or U749 (N_749,N_682,N_641);
or U750 (N_750,N_624,N_618);
or U751 (N_751,N_696,N_626);
nor U752 (N_752,N_619,N_648);
nand U753 (N_753,N_641,N_677);
nor U754 (N_754,N_675,N_698);
nor U755 (N_755,N_627,N_684);
nor U756 (N_756,N_680,N_673);
nand U757 (N_757,N_641,N_650);
or U758 (N_758,N_677,N_683);
nand U759 (N_759,N_610,N_611);
or U760 (N_760,N_614,N_681);
nand U761 (N_761,N_697,N_645);
nor U762 (N_762,N_671,N_673);
nand U763 (N_763,N_643,N_633);
or U764 (N_764,N_613,N_691);
and U765 (N_765,N_605,N_668);
xnor U766 (N_766,N_667,N_628);
nor U767 (N_767,N_666,N_629);
nor U768 (N_768,N_660,N_661);
and U769 (N_769,N_618,N_659);
or U770 (N_770,N_653,N_668);
or U771 (N_771,N_650,N_640);
and U772 (N_772,N_629,N_683);
and U773 (N_773,N_621,N_667);
and U774 (N_774,N_668,N_645);
or U775 (N_775,N_607,N_635);
nand U776 (N_776,N_696,N_681);
nand U777 (N_777,N_611,N_678);
nand U778 (N_778,N_661,N_687);
and U779 (N_779,N_670,N_603);
nand U780 (N_780,N_672,N_615);
nor U781 (N_781,N_674,N_603);
or U782 (N_782,N_600,N_697);
nand U783 (N_783,N_632,N_642);
nand U784 (N_784,N_660,N_698);
or U785 (N_785,N_611,N_658);
nand U786 (N_786,N_656,N_607);
or U787 (N_787,N_600,N_668);
nor U788 (N_788,N_603,N_677);
nor U789 (N_789,N_697,N_614);
nor U790 (N_790,N_689,N_631);
and U791 (N_791,N_675,N_606);
and U792 (N_792,N_604,N_631);
or U793 (N_793,N_617,N_673);
and U794 (N_794,N_642,N_650);
nor U795 (N_795,N_621,N_609);
nand U796 (N_796,N_693,N_670);
nand U797 (N_797,N_669,N_647);
nand U798 (N_798,N_644,N_697);
or U799 (N_799,N_607,N_612);
and U800 (N_800,N_715,N_736);
and U801 (N_801,N_779,N_768);
and U802 (N_802,N_777,N_788);
or U803 (N_803,N_733,N_794);
nand U804 (N_804,N_781,N_712);
nand U805 (N_805,N_741,N_738);
or U806 (N_806,N_707,N_764);
nand U807 (N_807,N_748,N_758);
nand U808 (N_808,N_792,N_772);
or U809 (N_809,N_744,N_753);
nand U810 (N_810,N_720,N_730);
nand U811 (N_811,N_785,N_767);
nand U812 (N_812,N_728,N_747);
nand U813 (N_813,N_766,N_765);
and U814 (N_814,N_756,N_722);
nor U815 (N_815,N_708,N_702);
or U816 (N_816,N_760,N_789);
or U817 (N_817,N_750,N_773);
nand U818 (N_818,N_787,N_752);
or U819 (N_819,N_740,N_795);
nor U820 (N_820,N_725,N_742);
and U821 (N_821,N_700,N_705);
or U822 (N_822,N_759,N_763);
and U823 (N_823,N_743,N_718);
nor U824 (N_824,N_726,N_737);
nand U825 (N_825,N_727,N_784);
or U826 (N_826,N_710,N_717);
and U827 (N_827,N_754,N_791);
nor U828 (N_828,N_783,N_778);
nor U829 (N_829,N_751,N_734);
and U830 (N_830,N_724,N_786);
and U831 (N_831,N_799,N_793);
nand U832 (N_832,N_735,N_775);
or U833 (N_833,N_755,N_723);
and U834 (N_834,N_704,N_732);
nor U835 (N_835,N_749,N_796);
nor U836 (N_836,N_701,N_721);
or U837 (N_837,N_713,N_782);
and U838 (N_838,N_745,N_757);
nor U839 (N_839,N_716,N_798);
and U840 (N_840,N_703,N_762);
nor U841 (N_841,N_719,N_729);
or U842 (N_842,N_769,N_714);
nor U843 (N_843,N_761,N_731);
nand U844 (N_844,N_739,N_746);
or U845 (N_845,N_774,N_770);
and U846 (N_846,N_780,N_797);
and U847 (N_847,N_709,N_790);
and U848 (N_848,N_771,N_706);
or U849 (N_849,N_776,N_711);
nand U850 (N_850,N_764,N_769);
and U851 (N_851,N_768,N_747);
nor U852 (N_852,N_740,N_711);
nor U853 (N_853,N_719,N_763);
nand U854 (N_854,N_711,N_785);
and U855 (N_855,N_763,N_736);
and U856 (N_856,N_713,N_780);
or U857 (N_857,N_778,N_725);
nand U858 (N_858,N_764,N_765);
nor U859 (N_859,N_774,N_702);
nor U860 (N_860,N_779,N_766);
or U861 (N_861,N_760,N_706);
or U862 (N_862,N_796,N_730);
or U863 (N_863,N_771,N_778);
nand U864 (N_864,N_792,N_731);
and U865 (N_865,N_757,N_782);
nor U866 (N_866,N_793,N_763);
nor U867 (N_867,N_725,N_792);
and U868 (N_868,N_789,N_751);
nor U869 (N_869,N_722,N_776);
and U870 (N_870,N_767,N_730);
nand U871 (N_871,N_725,N_746);
or U872 (N_872,N_773,N_776);
and U873 (N_873,N_705,N_769);
nand U874 (N_874,N_716,N_734);
and U875 (N_875,N_760,N_724);
nand U876 (N_876,N_766,N_759);
or U877 (N_877,N_778,N_764);
nor U878 (N_878,N_785,N_775);
and U879 (N_879,N_732,N_764);
and U880 (N_880,N_728,N_720);
nand U881 (N_881,N_707,N_748);
nand U882 (N_882,N_713,N_769);
nor U883 (N_883,N_732,N_788);
nand U884 (N_884,N_709,N_742);
or U885 (N_885,N_758,N_732);
nor U886 (N_886,N_764,N_754);
and U887 (N_887,N_776,N_783);
nor U888 (N_888,N_796,N_703);
nand U889 (N_889,N_796,N_759);
nand U890 (N_890,N_756,N_708);
or U891 (N_891,N_782,N_731);
and U892 (N_892,N_727,N_758);
nor U893 (N_893,N_721,N_772);
nor U894 (N_894,N_799,N_764);
nand U895 (N_895,N_793,N_746);
and U896 (N_896,N_785,N_758);
nand U897 (N_897,N_782,N_716);
nor U898 (N_898,N_736,N_794);
and U899 (N_899,N_737,N_731);
nand U900 (N_900,N_845,N_891);
or U901 (N_901,N_831,N_857);
or U902 (N_902,N_869,N_840);
nor U903 (N_903,N_828,N_830);
nor U904 (N_904,N_820,N_803);
and U905 (N_905,N_881,N_801);
and U906 (N_906,N_847,N_827);
or U907 (N_907,N_851,N_829);
nand U908 (N_908,N_874,N_855);
or U909 (N_909,N_841,N_808);
nand U910 (N_910,N_858,N_853);
nand U911 (N_911,N_863,N_868);
nor U912 (N_912,N_870,N_832);
or U913 (N_913,N_848,N_878);
nand U914 (N_914,N_873,N_814);
nand U915 (N_915,N_895,N_806);
and U916 (N_916,N_815,N_883);
xor U917 (N_917,N_896,N_835);
nor U918 (N_918,N_865,N_852);
and U919 (N_919,N_893,N_866);
and U920 (N_920,N_844,N_813);
and U921 (N_921,N_834,N_817);
and U922 (N_922,N_836,N_889);
or U923 (N_923,N_882,N_875);
nand U924 (N_924,N_876,N_862);
or U925 (N_925,N_879,N_850);
nor U926 (N_926,N_825,N_871);
nor U927 (N_927,N_884,N_838);
nor U928 (N_928,N_892,N_897);
nor U929 (N_929,N_854,N_821);
xor U930 (N_930,N_818,N_804);
or U931 (N_931,N_867,N_805);
or U932 (N_932,N_888,N_812);
and U933 (N_933,N_833,N_898);
or U934 (N_934,N_824,N_809);
nand U935 (N_935,N_885,N_886);
and U936 (N_936,N_899,N_819);
or U937 (N_937,N_846,N_877);
or U938 (N_938,N_864,N_856);
and U939 (N_939,N_823,N_810);
or U940 (N_940,N_861,N_860);
nor U941 (N_941,N_839,N_842);
nand U942 (N_942,N_872,N_826);
or U943 (N_943,N_887,N_807);
and U944 (N_944,N_822,N_843);
and U945 (N_945,N_816,N_890);
and U946 (N_946,N_811,N_859);
or U947 (N_947,N_802,N_880);
and U948 (N_948,N_837,N_894);
and U949 (N_949,N_849,N_800);
or U950 (N_950,N_886,N_860);
nor U951 (N_951,N_893,N_854);
or U952 (N_952,N_817,N_853);
nor U953 (N_953,N_817,N_842);
nor U954 (N_954,N_804,N_809);
nor U955 (N_955,N_872,N_854);
or U956 (N_956,N_866,N_844);
nand U957 (N_957,N_826,N_805);
nand U958 (N_958,N_802,N_803);
nor U959 (N_959,N_809,N_848);
and U960 (N_960,N_838,N_873);
nor U961 (N_961,N_873,N_819);
nor U962 (N_962,N_843,N_816);
or U963 (N_963,N_841,N_801);
and U964 (N_964,N_813,N_890);
nor U965 (N_965,N_864,N_851);
nor U966 (N_966,N_833,N_804);
nor U967 (N_967,N_898,N_856);
nor U968 (N_968,N_823,N_819);
or U969 (N_969,N_812,N_822);
or U970 (N_970,N_818,N_840);
or U971 (N_971,N_805,N_885);
nand U972 (N_972,N_849,N_844);
nand U973 (N_973,N_893,N_811);
or U974 (N_974,N_858,N_814);
and U975 (N_975,N_839,N_820);
nand U976 (N_976,N_863,N_870);
or U977 (N_977,N_879,N_847);
nor U978 (N_978,N_896,N_836);
or U979 (N_979,N_807,N_820);
nand U980 (N_980,N_845,N_821);
nand U981 (N_981,N_867,N_842);
or U982 (N_982,N_810,N_883);
and U983 (N_983,N_844,N_893);
nor U984 (N_984,N_828,N_843);
and U985 (N_985,N_898,N_808);
and U986 (N_986,N_816,N_840);
nor U987 (N_987,N_896,N_807);
nand U988 (N_988,N_837,N_831);
nor U989 (N_989,N_816,N_826);
and U990 (N_990,N_816,N_801);
nor U991 (N_991,N_828,N_851);
nor U992 (N_992,N_817,N_840);
nand U993 (N_993,N_833,N_881);
and U994 (N_994,N_854,N_806);
or U995 (N_995,N_850,N_866);
or U996 (N_996,N_807,N_859);
nand U997 (N_997,N_847,N_817);
or U998 (N_998,N_856,N_822);
or U999 (N_999,N_847,N_886);
xor U1000 (N_1000,N_964,N_909);
or U1001 (N_1001,N_915,N_902);
and U1002 (N_1002,N_978,N_918);
or U1003 (N_1003,N_998,N_951);
nor U1004 (N_1004,N_979,N_950);
nor U1005 (N_1005,N_935,N_931);
nand U1006 (N_1006,N_906,N_999);
and U1007 (N_1007,N_983,N_914);
nand U1008 (N_1008,N_997,N_928);
or U1009 (N_1009,N_993,N_985);
nor U1010 (N_1010,N_987,N_962);
nor U1011 (N_1011,N_900,N_940);
nor U1012 (N_1012,N_992,N_920);
nor U1013 (N_1013,N_986,N_965);
nor U1014 (N_1014,N_980,N_930);
and U1015 (N_1015,N_903,N_957);
or U1016 (N_1016,N_973,N_968);
or U1017 (N_1017,N_958,N_932);
and U1018 (N_1018,N_926,N_934);
or U1019 (N_1019,N_936,N_905);
nor U1020 (N_1020,N_982,N_911);
and U1021 (N_1021,N_946,N_921);
nand U1022 (N_1022,N_990,N_961);
or U1023 (N_1023,N_967,N_942);
xnor U1024 (N_1024,N_907,N_996);
nor U1025 (N_1025,N_922,N_971);
and U1026 (N_1026,N_904,N_948);
nor U1027 (N_1027,N_912,N_959);
or U1028 (N_1028,N_994,N_917);
nor U1029 (N_1029,N_974,N_953);
or U1030 (N_1030,N_916,N_970);
and U1031 (N_1031,N_960,N_989);
and U1032 (N_1032,N_913,N_919);
or U1033 (N_1033,N_945,N_910);
nor U1034 (N_1034,N_924,N_966);
nand U1035 (N_1035,N_943,N_956);
and U1036 (N_1036,N_954,N_977);
nor U1037 (N_1037,N_963,N_952);
or U1038 (N_1038,N_991,N_944);
or U1039 (N_1039,N_933,N_938);
nand U1040 (N_1040,N_927,N_955);
or U1041 (N_1041,N_908,N_981);
and U1042 (N_1042,N_925,N_988);
and U1043 (N_1043,N_947,N_923);
and U1044 (N_1044,N_975,N_949);
and U1045 (N_1045,N_976,N_972);
and U1046 (N_1046,N_969,N_929);
nor U1047 (N_1047,N_937,N_901);
or U1048 (N_1048,N_995,N_939);
and U1049 (N_1049,N_941,N_984);
nand U1050 (N_1050,N_923,N_922);
nand U1051 (N_1051,N_979,N_927);
nor U1052 (N_1052,N_998,N_950);
nand U1053 (N_1053,N_900,N_927);
or U1054 (N_1054,N_973,N_932);
or U1055 (N_1055,N_994,N_993);
nor U1056 (N_1056,N_917,N_914);
nand U1057 (N_1057,N_945,N_938);
and U1058 (N_1058,N_986,N_920);
and U1059 (N_1059,N_922,N_909);
and U1060 (N_1060,N_982,N_977);
nand U1061 (N_1061,N_988,N_930);
and U1062 (N_1062,N_993,N_918);
nor U1063 (N_1063,N_921,N_923);
nand U1064 (N_1064,N_904,N_951);
or U1065 (N_1065,N_902,N_996);
nand U1066 (N_1066,N_988,N_907);
and U1067 (N_1067,N_940,N_983);
nor U1068 (N_1068,N_952,N_945);
or U1069 (N_1069,N_909,N_904);
and U1070 (N_1070,N_932,N_938);
or U1071 (N_1071,N_962,N_981);
and U1072 (N_1072,N_942,N_986);
nand U1073 (N_1073,N_928,N_915);
nand U1074 (N_1074,N_990,N_952);
nor U1075 (N_1075,N_987,N_966);
nor U1076 (N_1076,N_946,N_913);
nand U1077 (N_1077,N_965,N_997);
and U1078 (N_1078,N_900,N_985);
nor U1079 (N_1079,N_936,N_948);
and U1080 (N_1080,N_901,N_945);
or U1081 (N_1081,N_964,N_968);
nand U1082 (N_1082,N_997,N_953);
or U1083 (N_1083,N_916,N_926);
and U1084 (N_1084,N_921,N_940);
and U1085 (N_1085,N_944,N_957);
nor U1086 (N_1086,N_971,N_937);
and U1087 (N_1087,N_934,N_985);
nand U1088 (N_1088,N_923,N_941);
or U1089 (N_1089,N_994,N_930);
nand U1090 (N_1090,N_929,N_983);
nand U1091 (N_1091,N_935,N_986);
or U1092 (N_1092,N_934,N_962);
nor U1093 (N_1093,N_951,N_900);
or U1094 (N_1094,N_993,N_902);
and U1095 (N_1095,N_930,N_948);
nor U1096 (N_1096,N_944,N_932);
nand U1097 (N_1097,N_988,N_908);
xor U1098 (N_1098,N_935,N_944);
nor U1099 (N_1099,N_975,N_973);
and U1100 (N_1100,N_1010,N_1075);
or U1101 (N_1101,N_1048,N_1009);
or U1102 (N_1102,N_1020,N_1095);
nand U1103 (N_1103,N_1094,N_1038);
and U1104 (N_1104,N_1053,N_1005);
nor U1105 (N_1105,N_1080,N_1070);
and U1106 (N_1106,N_1004,N_1090);
nand U1107 (N_1107,N_1049,N_1050);
nor U1108 (N_1108,N_1069,N_1067);
or U1109 (N_1109,N_1086,N_1076);
and U1110 (N_1110,N_1029,N_1024);
and U1111 (N_1111,N_1059,N_1011);
and U1112 (N_1112,N_1008,N_1033);
and U1113 (N_1113,N_1098,N_1035);
nor U1114 (N_1114,N_1021,N_1003);
nor U1115 (N_1115,N_1012,N_1045);
nor U1116 (N_1116,N_1044,N_1064);
or U1117 (N_1117,N_1071,N_1041);
and U1118 (N_1118,N_1072,N_1055);
and U1119 (N_1119,N_1017,N_1087);
and U1120 (N_1120,N_1062,N_1074);
nor U1121 (N_1121,N_1066,N_1007);
nor U1122 (N_1122,N_1068,N_1025);
and U1123 (N_1123,N_1063,N_1036);
nor U1124 (N_1124,N_1030,N_1027);
or U1125 (N_1125,N_1015,N_1037);
nor U1126 (N_1126,N_1023,N_1077);
and U1127 (N_1127,N_1052,N_1073);
nand U1128 (N_1128,N_1001,N_1078);
nand U1129 (N_1129,N_1043,N_1083);
and U1130 (N_1130,N_1054,N_1016);
and U1131 (N_1131,N_1002,N_1022);
nand U1132 (N_1132,N_1065,N_1032);
nand U1133 (N_1133,N_1096,N_1092);
and U1134 (N_1134,N_1000,N_1099);
nor U1135 (N_1135,N_1028,N_1014);
and U1136 (N_1136,N_1061,N_1047);
and U1137 (N_1137,N_1089,N_1026);
or U1138 (N_1138,N_1040,N_1039);
nor U1139 (N_1139,N_1019,N_1013);
nand U1140 (N_1140,N_1057,N_1006);
nor U1141 (N_1141,N_1097,N_1084);
nor U1142 (N_1142,N_1056,N_1093);
nand U1143 (N_1143,N_1081,N_1018);
nand U1144 (N_1144,N_1091,N_1088);
and U1145 (N_1145,N_1060,N_1082);
nand U1146 (N_1146,N_1058,N_1042);
nand U1147 (N_1147,N_1046,N_1085);
or U1148 (N_1148,N_1079,N_1034);
nand U1149 (N_1149,N_1031,N_1051);
nor U1150 (N_1150,N_1022,N_1055);
nand U1151 (N_1151,N_1060,N_1062);
or U1152 (N_1152,N_1067,N_1068);
or U1153 (N_1153,N_1083,N_1086);
and U1154 (N_1154,N_1090,N_1021);
or U1155 (N_1155,N_1062,N_1042);
nor U1156 (N_1156,N_1078,N_1079);
or U1157 (N_1157,N_1063,N_1085);
or U1158 (N_1158,N_1065,N_1078);
or U1159 (N_1159,N_1030,N_1023);
nor U1160 (N_1160,N_1013,N_1006);
or U1161 (N_1161,N_1050,N_1027);
nor U1162 (N_1162,N_1010,N_1019);
nor U1163 (N_1163,N_1071,N_1069);
or U1164 (N_1164,N_1057,N_1048);
or U1165 (N_1165,N_1093,N_1015);
xor U1166 (N_1166,N_1030,N_1048);
nor U1167 (N_1167,N_1047,N_1050);
nand U1168 (N_1168,N_1015,N_1076);
nor U1169 (N_1169,N_1095,N_1022);
nor U1170 (N_1170,N_1064,N_1097);
or U1171 (N_1171,N_1015,N_1062);
nor U1172 (N_1172,N_1037,N_1096);
nor U1173 (N_1173,N_1055,N_1087);
nand U1174 (N_1174,N_1070,N_1051);
nand U1175 (N_1175,N_1096,N_1011);
nand U1176 (N_1176,N_1064,N_1036);
nand U1177 (N_1177,N_1010,N_1021);
or U1178 (N_1178,N_1027,N_1017);
nor U1179 (N_1179,N_1065,N_1070);
nand U1180 (N_1180,N_1006,N_1062);
or U1181 (N_1181,N_1092,N_1080);
nor U1182 (N_1182,N_1076,N_1023);
and U1183 (N_1183,N_1000,N_1061);
or U1184 (N_1184,N_1021,N_1042);
or U1185 (N_1185,N_1054,N_1044);
nand U1186 (N_1186,N_1019,N_1051);
and U1187 (N_1187,N_1027,N_1010);
or U1188 (N_1188,N_1025,N_1042);
or U1189 (N_1189,N_1000,N_1016);
or U1190 (N_1190,N_1053,N_1088);
nand U1191 (N_1191,N_1042,N_1077);
xnor U1192 (N_1192,N_1054,N_1086);
and U1193 (N_1193,N_1083,N_1090);
nor U1194 (N_1194,N_1008,N_1083);
and U1195 (N_1195,N_1044,N_1089);
nand U1196 (N_1196,N_1082,N_1005);
or U1197 (N_1197,N_1083,N_1098);
and U1198 (N_1198,N_1083,N_1044);
and U1199 (N_1199,N_1085,N_1072);
or U1200 (N_1200,N_1149,N_1152);
or U1201 (N_1201,N_1178,N_1196);
and U1202 (N_1202,N_1127,N_1153);
nand U1203 (N_1203,N_1100,N_1108);
nand U1204 (N_1204,N_1135,N_1130);
and U1205 (N_1205,N_1176,N_1165);
nand U1206 (N_1206,N_1180,N_1117);
and U1207 (N_1207,N_1177,N_1116);
or U1208 (N_1208,N_1144,N_1118);
or U1209 (N_1209,N_1156,N_1133);
or U1210 (N_1210,N_1145,N_1143);
nand U1211 (N_1211,N_1147,N_1183);
nand U1212 (N_1212,N_1106,N_1174);
and U1213 (N_1213,N_1142,N_1187);
nor U1214 (N_1214,N_1131,N_1128);
and U1215 (N_1215,N_1105,N_1138);
and U1216 (N_1216,N_1120,N_1161);
nor U1217 (N_1217,N_1157,N_1181);
and U1218 (N_1218,N_1151,N_1129);
or U1219 (N_1219,N_1192,N_1172);
and U1220 (N_1220,N_1170,N_1164);
nand U1221 (N_1221,N_1115,N_1101);
and U1222 (N_1222,N_1122,N_1150);
nand U1223 (N_1223,N_1111,N_1182);
nor U1224 (N_1224,N_1195,N_1109);
or U1225 (N_1225,N_1102,N_1137);
or U1226 (N_1226,N_1191,N_1146);
nand U1227 (N_1227,N_1136,N_1175);
or U1228 (N_1228,N_1159,N_1162);
and U1229 (N_1229,N_1154,N_1167);
and U1230 (N_1230,N_1173,N_1123);
or U1231 (N_1231,N_1125,N_1107);
nand U1232 (N_1232,N_1158,N_1134);
or U1233 (N_1233,N_1140,N_1168);
and U1234 (N_1234,N_1199,N_1188);
and U1235 (N_1235,N_1194,N_1124);
and U1236 (N_1236,N_1179,N_1132);
nand U1237 (N_1237,N_1193,N_1103);
and U1238 (N_1238,N_1171,N_1197);
and U1239 (N_1239,N_1186,N_1190);
and U1240 (N_1240,N_1184,N_1189);
nor U1241 (N_1241,N_1119,N_1169);
and U1242 (N_1242,N_1141,N_1160);
or U1243 (N_1243,N_1114,N_1121);
and U1244 (N_1244,N_1113,N_1110);
nor U1245 (N_1245,N_1163,N_1148);
or U1246 (N_1246,N_1166,N_1104);
or U1247 (N_1247,N_1155,N_1126);
and U1248 (N_1248,N_1198,N_1139);
nor U1249 (N_1249,N_1112,N_1185);
nor U1250 (N_1250,N_1110,N_1191);
nand U1251 (N_1251,N_1198,N_1121);
or U1252 (N_1252,N_1159,N_1108);
and U1253 (N_1253,N_1131,N_1159);
or U1254 (N_1254,N_1162,N_1145);
nor U1255 (N_1255,N_1130,N_1150);
nand U1256 (N_1256,N_1113,N_1158);
nor U1257 (N_1257,N_1117,N_1133);
or U1258 (N_1258,N_1199,N_1154);
and U1259 (N_1259,N_1190,N_1160);
and U1260 (N_1260,N_1145,N_1182);
or U1261 (N_1261,N_1101,N_1139);
nand U1262 (N_1262,N_1137,N_1153);
nand U1263 (N_1263,N_1144,N_1150);
nor U1264 (N_1264,N_1152,N_1140);
nor U1265 (N_1265,N_1186,N_1183);
or U1266 (N_1266,N_1176,N_1192);
nor U1267 (N_1267,N_1192,N_1120);
or U1268 (N_1268,N_1154,N_1188);
and U1269 (N_1269,N_1162,N_1117);
nand U1270 (N_1270,N_1190,N_1168);
nor U1271 (N_1271,N_1135,N_1132);
nand U1272 (N_1272,N_1160,N_1121);
and U1273 (N_1273,N_1175,N_1119);
nor U1274 (N_1274,N_1139,N_1164);
nand U1275 (N_1275,N_1110,N_1178);
nand U1276 (N_1276,N_1169,N_1137);
nor U1277 (N_1277,N_1102,N_1131);
and U1278 (N_1278,N_1159,N_1169);
or U1279 (N_1279,N_1169,N_1160);
and U1280 (N_1280,N_1125,N_1116);
and U1281 (N_1281,N_1130,N_1195);
nand U1282 (N_1282,N_1140,N_1119);
and U1283 (N_1283,N_1113,N_1102);
nand U1284 (N_1284,N_1101,N_1147);
and U1285 (N_1285,N_1110,N_1108);
or U1286 (N_1286,N_1152,N_1151);
nor U1287 (N_1287,N_1188,N_1168);
nand U1288 (N_1288,N_1100,N_1103);
and U1289 (N_1289,N_1179,N_1151);
nor U1290 (N_1290,N_1108,N_1129);
nand U1291 (N_1291,N_1132,N_1168);
nor U1292 (N_1292,N_1199,N_1110);
nand U1293 (N_1293,N_1155,N_1191);
and U1294 (N_1294,N_1118,N_1136);
or U1295 (N_1295,N_1168,N_1147);
nor U1296 (N_1296,N_1155,N_1121);
and U1297 (N_1297,N_1183,N_1141);
nand U1298 (N_1298,N_1145,N_1127);
nand U1299 (N_1299,N_1140,N_1109);
nor U1300 (N_1300,N_1287,N_1231);
or U1301 (N_1301,N_1220,N_1272);
nor U1302 (N_1302,N_1201,N_1233);
and U1303 (N_1303,N_1210,N_1278);
nor U1304 (N_1304,N_1240,N_1243);
nand U1305 (N_1305,N_1236,N_1259);
nor U1306 (N_1306,N_1257,N_1224);
nand U1307 (N_1307,N_1211,N_1234);
nor U1308 (N_1308,N_1203,N_1217);
nor U1309 (N_1309,N_1265,N_1242);
and U1310 (N_1310,N_1291,N_1248);
or U1311 (N_1311,N_1268,N_1261);
nor U1312 (N_1312,N_1275,N_1232);
nor U1313 (N_1313,N_1239,N_1225);
nand U1314 (N_1314,N_1295,N_1271);
nor U1315 (N_1315,N_1237,N_1250);
or U1316 (N_1316,N_1222,N_1263);
and U1317 (N_1317,N_1200,N_1230);
nand U1318 (N_1318,N_1293,N_1204);
nand U1319 (N_1319,N_1245,N_1251);
or U1320 (N_1320,N_1267,N_1297);
or U1321 (N_1321,N_1282,N_1253);
and U1322 (N_1322,N_1256,N_1208);
and U1323 (N_1323,N_1213,N_1286);
or U1324 (N_1324,N_1254,N_1221);
or U1325 (N_1325,N_1266,N_1283);
nand U1326 (N_1326,N_1262,N_1216);
nand U1327 (N_1327,N_1247,N_1276);
and U1328 (N_1328,N_1264,N_1258);
or U1329 (N_1329,N_1207,N_1290);
nand U1330 (N_1330,N_1229,N_1289);
nand U1331 (N_1331,N_1284,N_1241);
or U1332 (N_1332,N_1285,N_1212);
or U1333 (N_1333,N_1255,N_1223);
nand U1334 (N_1334,N_1206,N_1246);
nand U1335 (N_1335,N_1281,N_1273);
nor U1336 (N_1336,N_1226,N_1277);
nand U1337 (N_1337,N_1235,N_1298);
nor U1338 (N_1338,N_1227,N_1209);
or U1339 (N_1339,N_1214,N_1260);
or U1340 (N_1340,N_1202,N_1279);
nand U1341 (N_1341,N_1218,N_1238);
nand U1342 (N_1342,N_1274,N_1294);
nor U1343 (N_1343,N_1228,N_1280);
nor U1344 (N_1344,N_1296,N_1292);
or U1345 (N_1345,N_1269,N_1288);
and U1346 (N_1346,N_1244,N_1299);
and U1347 (N_1347,N_1249,N_1219);
or U1348 (N_1348,N_1252,N_1205);
and U1349 (N_1349,N_1215,N_1270);
xnor U1350 (N_1350,N_1211,N_1268);
and U1351 (N_1351,N_1250,N_1277);
nand U1352 (N_1352,N_1202,N_1274);
nand U1353 (N_1353,N_1293,N_1212);
and U1354 (N_1354,N_1261,N_1229);
nor U1355 (N_1355,N_1288,N_1290);
and U1356 (N_1356,N_1266,N_1228);
nor U1357 (N_1357,N_1287,N_1232);
or U1358 (N_1358,N_1296,N_1260);
nor U1359 (N_1359,N_1215,N_1203);
and U1360 (N_1360,N_1289,N_1257);
and U1361 (N_1361,N_1283,N_1277);
and U1362 (N_1362,N_1286,N_1291);
nor U1363 (N_1363,N_1215,N_1247);
and U1364 (N_1364,N_1290,N_1248);
nor U1365 (N_1365,N_1265,N_1215);
nor U1366 (N_1366,N_1205,N_1273);
nand U1367 (N_1367,N_1292,N_1254);
nand U1368 (N_1368,N_1208,N_1273);
nor U1369 (N_1369,N_1215,N_1209);
nand U1370 (N_1370,N_1205,N_1218);
nand U1371 (N_1371,N_1271,N_1214);
or U1372 (N_1372,N_1223,N_1228);
nand U1373 (N_1373,N_1206,N_1277);
nor U1374 (N_1374,N_1225,N_1260);
and U1375 (N_1375,N_1216,N_1214);
or U1376 (N_1376,N_1269,N_1254);
or U1377 (N_1377,N_1212,N_1202);
nor U1378 (N_1378,N_1282,N_1209);
and U1379 (N_1379,N_1206,N_1270);
or U1380 (N_1380,N_1208,N_1240);
or U1381 (N_1381,N_1267,N_1299);
nor U1382 (N_1382,N_1264,N_1238);
or U1383 (N_1383,N_1231,N_1224);
xor U1384 (N_1384,N_1202,N_1272);
or U1385 (N_1385,N_1278,N_1261);
nor U1386 (N_1386,N_1237,N_1282);
or U1387 (N_1387,N_1211,N_1260);
and U1388 (N_1388,N_1267,N_1207);
or U1389 (N_1389,N_1223,N_1231);
or U1390 (N_1390,N_1249,N_1294);
or U1391 (N_1391,N_1212,N_1280);
and U1392 (N_1392,N_1248,N_1286);
and U1393 (N_1393,N_1279,N_1243);
nand U1394 (N_1394,N_1220,N_1247);
and U1395 (N_1395,N_1216,N_1292);
or U1396 (N_1396,N_1286,N_1274);
xnor U1397 (N_1397,N_1268,N_1226);
or U1398 (N_1398,N_1204,N_1225);
or U1399 (N_1399,N_1205,N_1261);
and U1400 (N_1400,N_1350,N_1394);
and U1401 (N_1401,N_1319,N_1383);
or U1402 (N_1402,N_1302,N_1326);
nand U1403 (N_1403,N_1354,N_1351);
nand U1404 (N_1404,N_1316,N_1338);
nor U1405 (N_1405,N_1344,N_1301);
nor U1406 (N_1406,N_1340,N_1311);
and U1407 (N_1407,N_1324,N_1332);
nand U1408 (N_1408,N_1317,N_1337);
nor U1409 (N_1409,N_1387,N_1361);
or U1410 (N_1410,N_1385,N_1365);
nor U1411 (N_1411,N_1359,N_1379);
and U1412 (N_1412,N_1305,N_1362);
and U1413 (N_1413,N_1306,N_1370);
nor U1414 (N_1414,N_1380,N_1352);
or U1415 (N_1415,N_1393,N_1347);
and U1416 (N_1416,N_1366,N_1349);
or U1417 (N_1417,N_1396,N_1390);
and U1418 (N_1418,N_1329,N_1377);
and U1419 (N_1419,N_1395,N_1348);
nor U1420 (N_1420,N_1307,N_1323);
nor U1421 (N_1421,N_1392,N_1309);
nand U1422 (N_1422,N_1388,N_1321);
nor U1423 (N_1423,N_1310,N_1355);
and U1424 (N_1424,N_1378,N_1357);
nand U1425 (N_1425,N_1334,N_1360);
nand U1426 (N_1426,N_1315,N_1368);
and U1427 (N_1427,N_1330,N_1322);
nor U1428 (N_1428,N_1364,N_1343);
nand U1429 (N_1429,N_1384,N_1325);
nor U1430 (N_1430,N_1318,N_1300);
nand U1431 (N_1431,N_1346,N_1372);
nand U1432 (N_1432,N_1399,N_1373);
or U1433 (N_1433,N_1371,N_1304);
or U1434 (N_1434,N_1333,N_1376);
or U1435 (N_1435,N_1327,N_1397);
or U1436 (N_1436,N_1342,N_1389);
nand U1437 (N_1437,N_1386,N_1341);
and U1438 (N_1438,N_1313,N_1382);
nand U1439 (N_1439,N_1369,N_1339);
nor U1440 (N_1440,N_1374,N_1312);
or U1441 (N_1441,N_1336,N_1363);
or U1442 (N_1442,N_1398,N_1367);
nand U1443 (N_1443,N_1314,N_1356);
and U1444 (N_1444,N_1320,N_1335);
or U1445 (N_1445,N_1358,N_1375);
nor U1446 (N_1446,N_1303,N_1331);
and U1447 (N_1447,N_1308,N_1353);
or U1448 (N_1448,N_1381,N_1345);
nor U1449 (N_1449,N_1391,N_1328);
nor U1450 (N_1450,N_1370,N_1360);
nand U1451 (N_1451,N_1303,N_1375);
nand U1452 (N_1452,N_1326,N_1304);
nor U1453 (N_1453,N_1378,N_1354);
and U1454 (N_1454,N_1374,N_1305);
nor U1455 (N_1455,N_1345,N_1317);
nand U1456 (N_1456,N_1395,N_1345);
nand U1457 (N_1457,N_1372,N_1347);
nor U1458 (N_1458,N_1365,N_1338);
and U1459 (N_1459,N_1368,N_1380);
and U1460 (N_1460,N_1350,N_1348);
nand U1461 (N_1461,N_1390,N_1371);
nand U1462 (N_1462,N_1374,N_1301);
nor U1463 (N_1463,N_1300,N_1385);
and U1464 (N_1464,N_1387,N_1301);
or U1465 (N_1465,N_1341,N_1323);
nor U1466 (N_1466,N_1316,N_1370);
and U1467 (N_1467,N_1345,N_1340);
and U1468 (N_1468,N_1381,N_1378);
or U1469 (N_1469,N_1325,N_1320);
or U1470 (N_1470,N_1328,N_1331);
nor U1471 (N_1471,N_1322,N_1325);
and U1472 (N_1472,N_1395,N_1325);
or U1473 (N_1473,N_1309,N_1365);
or U1474 (N_1474,N_1341,N_1371);
nand U1475 (N_1475,N_1390,N_1381);
and U1476 (N_1476,N_1384,N_1315);
nor U1477 (N_1477,N_1397,N_1313);
or U1478 (N_1478,N_1346,N_1351);
and U1479 (N_1479,N_1363,N_1361);
or U1480 (N_1480,N_1311,N_1309);
and U1481 (N_1481,N_1300,N_1398);
or U1482 (N_1482,N_1328,N_1342);
or U1483 (N_1483,N_1366,N_1322);
xor U1484 (N_1484,N_1346,N_1355);
nand U1485 (N_1485,N_1348,N_1356);
xor U1486 (N_1486,N_1347,N_1341);
nand U1487 (N_1487,N_1310,N_1356);
and U1488 (N_1488,N_1333,N_1368);
nor U1489 (N_1489,N_1384,N_1360);
nor U1490 (N_1490,N_1318,N_1399);
nand U1491 (N_1491,N_1324,N_1322);
and U1492 (N_1492,N_1325,N_1324);
nand U1493 (N_1493,N_1399,N_1345);
nand U1494 (N_1494,N_1366,N_1351);
nor U1495 (N_1495,N_1326,N_1365);
and U1496 (N_1496,N_1385,N_1354);
nor U1497 (N_1497,N_1376,N_1357);
nand U1498 (N_1498,N_1378,N_1335);
or U1499 (N_1499,N_1377,N_1374);
nor U1500 (N_1500,N_1406,N_1428);
or U1501 (N_1501,N_1498,N_1415);
and U1502 (N_1502,N_1496,N_1460);
nand U1503 (N_1503,N_1417,N_1416);
nand U1504 (N_1504,N_1434,N_1447);
nand U1505 (N_1505,N_1418,N_1450);
nand U1506 (N_1506,N_1432,N_1403);
and U1507 (N_1507,N_1412,N_1409);
nand U1508 (N_1508,N_1446,N_1471);
nand U1509 (N_1509,N_1454,N_1497);
nand U1510 (N_1510,N_1451,N_1469);
and U1511 (N_1511,N_1488,N_1429);
or U1512 (N_1512,N_1400,N_1492);
nand U1513 (N_1513,N_1458,N_1401);
and U1514 (N_1514,N_1455,N_1475);
or U1515 (N_1515,N_1440,N_1480);
nor U1516 (N_1516,N_1402,N_1425);
nor U1517 (N_1517,N_1491,N_1437);
nor U1518 (N_1518,N_1464,N_1421);
and U1519 (N_1519,N_1459,N_1482);
nand U1520 (N_1520,N_1404,N_1493);
and U1521 (N_1521,N_1473,N_1448);
and U1522 (N_1522,N_1445,N_1462);
and U1523 (N_1523,N_1481,N_1490);
and U1524 (N_1524,N_1463,N_1405);
nor U1525 (N_1525,N_1478,N_1472);
and U1526 (N_1526,N_1479,N_1433);
nor U1527 (N_1527,N_1430,N_1495);
nor U1528 (N_1528,N_1407,N_1453);
nand U1529 (N_1529,N_1443,N_1420);
nor U1530 (N_1530,N_1424,N_1499);
nand U1531 (N_1531,N_1423,N_1441);
nand U1532 (N_1532,N_1465,N_1452);
and U1533 (N_1533,N_1484,N_1467);
nand U1534 (N_1534,N_1466,N_1422);
and U1535 (N_1535,N_1477,N_1435);
xnor U1536 (N_1536,N_1494,N_1486);
nand U1537 (N_1537,N_1427,N_1487);
and U1538 (N_1538,N_1438,N_1449);
or U1539 (N_1539,N_1483,N_1468);
nand U1540 (N_1540,N_1439,N_1442);
nand U1541 (N_1541,N_1457,N_1436);
nor U1542 (N_1542,N_1474,N_1485);
nand U1543 (N_1543,N_1489,N_1408);
nand U1544 (N_1544,N_1413,N_1419);
and U1545 (N_1545,N_1410,N_1476);
or U1546 (N_1546,N_1461,N_1431);
nor U1547 (N_1547,N_1444,N_1426);
or U1548 (N_1548,N_1456,N_1470);
nand U1549 (N_1549,N_1414,N_1411);
and U1550 (N_1550,N_1421,N_1444);
or U1551 (N_1551,N_1416,N_1412);
xor U1552 (N_1552,N_1422,N_1493);
and U1553 (N_1553,N_1444,N_1432);
or U1554 (N_1554,N_1439,N_1440);
nand U1555 (N_1555,N_1430,N_1413);
nand U1556 (N_1556,N_1484,N_1453);
nand U1557 (N_1557,N_1462,N_1461);
and U1558 (N_1558,N_1441,N_1497);
and U1559 (N_1559,N_1498,N_1489);
and U1560 (N_1560,N_1474,N_1401);
nor U1561 (N_1561,N_1435,N_1445);
or U1562 (N_1562,N_1469,N_1448);
or U1563 (N_1563,N_1471,N_1429);
and U1564 (N_1564,N_1412,N_1441);
nor U1565 (N_1565,N_1474,N_1444);
nand U1566 (N_1566,N_1497,N_1434);
or U1567 (N_1567,N_1442,N_1468);
nand U1568 (N_1568,N_1469,N_1446);
nand U1569 (N_1569,N_1418,N_1447);
or U1570 (N_1570,N_1417,N_1401);
nand U1571 (N_1571,N_1426,N_1423);
and U1572 (N_1572,N_1474,N_1472);
nor U1573 (N_1573,N_1422,N_1438);
nand U1574 (N_1574,N_1489,N_1475);
and U1575 (N_1575,N_1419,N_1431);
and U1576 (N_1576,N_1436,N_1469);
or U1577 (N_1577,N_1458,N_1465);
and U1578 (N_1578,N_1438,N_1440);
or U1579 (N_1579,N_1437,N_1484);
nor U1580 (N_1580,N_1495,N_1466);
and U1581 (N_1581,N_1435,N_1413);
nor U1582 (N_1582,N_1493,N_1414);
nor U1583 (N_1583,N_1460,N_1461);
nand U1584 (N_1584,N_1453,N_1444);
xor U1585 (N_1585,N_1430,N_1421);
or U1586 (N_1586,N_1455,N_1402);
and U1587 (N_1587,N_1410,N_1430);
and U1588 (N_1588,N_1473,N_1490);
and U1589 (N_1589,N_1412,N_1496);
or U1590 (N_1590,N_1476,N_1458);
and U1591 (N_1591,N_1477,N_1408);
and U1592 (N_1592,N_1438,N_1460);
or U1593 (N_1593,N_1408,N_1472);
nand U1594 (N_1594,N_1460,N_1406);
nand U1595 (N_1595,N_1416,N_1466);
or U1596 (N_1596,N_1420,N_1461);
or U1597 (N_1597,N_1431,N_1464);
or U1598 (N_1598,N_1436,N_1484);
or U1599 (N_1599,N_1429,N_1482);
nand U1600 (N_1600,N_1531,N_1536);
and U1601 (N_1601,N_1507,N_1551);
and U1602 (N_1602,N_1532,N_1586);
or U1603 (N_1603,N_1535,N_1557);
xor U1604 (N_1604,N_1581,N_1588);
nand U1605 (N_1605,N_1528,N_1598);
nand U1606 (N_1606,N_1504,N_1589);
and U1607 (N_1607,N_1518,N_1526);
nand U1608 (N_1608,N_1582,N_1515);
and U1609 (N_1609,N_1546,N_1502);
and U1610 (N_1610,N_1570,N_1578);
nand U1611 (N_1611,N_1592,N_1508);
and U1612 (N_1612,N_1511,N_1549);
nor U1613 (N_1613,N_1556,N_1540);
and U1614 (N_1614,N_1571,N_1545);
nand U1615 (N_1615,N_1519,N_1501);
or U1616 (N_1616,N_1523,N_1568);
nor U1617 (N_1617,N_1553,N_1506);
nor U1618 (N_1618,N_1550,N_1560);
nor U1619 (N_1619,N_1559,N_1561);
and U1620 (N_1620,N_1513,N_1530);
and U1621 (N_1621,N_1580,N_1522);
and U1622 (N_1622,N_1579,N_1572);
nand U1623 (N_1623,N_1547,N_1577);
and U1624 (N_1624,N_1533,N_1525);
nor U1625 (N_1625,N_1599,N_1552);
or U1626 (N_1626,N_1583,N_1539);
and U1627 (N_1627,N_1529,N_1587);
and U1628 (N_1628,N_1542,N_1590);
or U1629 (N_1629,N_1521,N_1537);
nor U1630 (N_1630,N_1509,N_1524);
or U1631 (N_1631,N_1574,N_1543);
or U1632 (N_1632,N_1595,N_1569);
nand U1633 (N_1633,N_1510,N_1558);
and U1634 (N_1634,N_1576,N_1591);
and U1635 (N_1635,N_1562,N_1534);
or U1636 (N_1636,N_1548,N_1512);
and U1637 (N_1637,N_1503,N_1573);
nand U1638 (N_1638,N_1596,N_1585);
or U1639 (N_1639,N_1555,N_1593);
nand U1640 (N_1640,N_1597,N_1564);
and U1641 (N_1641,N_1516,N_1541);
or U1642 (N_1642,N_1575,N_1566);
and U1643 (N_1643,N_1567,N_1514);
nor U1644 (N_1644,N_1500,N_1584);
or U1645 (N_1645,N_1527,N_1563);
and U1646 (N_1646,N_1505,N_1554);
and U1647 (N_1647,N_1594,N_1544);
nor U1648 (N_1648,N_1517,N_1538);
nand U1649 (N_1649,N_1520,N_1565);
nand U1650 (N_1650,N_1532,N_1570);
and U1651 (N_1651,N_1586,N_1547);
and U1652 (N_1652,N_1507,N_1578);
nand U1653 (N_1653,N_1579,N_1515);
or U1654 (N_1654,N_1599,N_1593);
and U1655 (N_1655,N_1563,N_1510);
nor U1656 (N_1656,N_1521,N_1550);
and U1657 (N_1657,N_1523,N_1509);
nand U1658 (N_1658,N_1588,N_1528);
and U1659 (N_1659,N_1518,N_1592);
or U1660 (N_1660,N_1514,N_1598);
and U1661 (N_1661,N_1590,N_1568);
nor U1662 (N_1662,N_1587,N_1572);
and U1663 (N_1663,N_1570,N_1584);
nand U1664 (N_1664,N_1528,N_1567);
and U1665 (N_1665,N_1543,N_1566);
nand U1666 (N_1666,N_1500,N_1549);
and U1667 (N_1667,N_1573,N_1545);
and U1668 (N_1668,N_1559,N_1535);
nor U1669 (N_1669,N_1569,N_1593);
or U1670 (N_1670,N_1570,N_1556);
and U1671 (N_1671,N_1595,N_1567);
nand U1672 (N_1672,N_1571,N_1557);
or U1673 (N_1673,N_1567,N_1516);
nor U1674 (N_1674,N_1544,N_1531);
or U1675 (N_1675,N_1581,N_1529);
or U1676 (N_1676,N_1556,N_1583);
or U1677 (N_1677,N_1584,N_1572);
nor U1678 (N_1678,N_1586,N_1536);
or U1679 (N_1679,N_1574,N_1525);
nand U1680 (N_1680,N_1565,N_1552);
nor U1681 (N_1681,N_1520,N_1570);
nor U1682 (N_1682,N_1528,N_1586);
nand U1683 (N_1683,N_1565,N_1558);
nand U1684 (N_1684,N_1564,N_1555);
and U1685 (N_1685,N_1545,N_1553);
and U1686 (N_1686,N_1550,N_1508);
and U1687 (N_1687,N_1505,N_1567);
nand U1688 (N_1688,N_1578,N_1514);
nor U1689 (N_1689,N_1584,N_1547);
and U1690 (N_1690,N_1593,N_1537);
nor U1691 (N_1691,N_1542,N_1552);
nor U1692 (N_1692,N_1583,N_1518);
nor U1693 (N_1693,N_1598,N_1583);
nor U1694 (N_1694,N_1540,N_1502);
or U1695 (N_1695,N_1598,N_1577);
nor U1696 (N_1696,N_1580,N_1501);
or U1697 (N_1697,N_1536,N_1522);
and U1698 (N_1698,N_1519,N_1540);
nand U1699 (N_1699,N_1505,N_1562);
nand U1700 (N_1700,N_1689,N_1697);
nor U1701 (N_1701,N_1650,N_1694);
nand U1702 (N_1702,N_1661,N_1626);
nor U1703 (N_1703,N_1691,N_1649);
nor U1704 (N_1704,N_1682,N_1617);
nor U1705 (N_1705,N_1656,N_1605);
or U1706 (N_1706,N_1651,N_1623);
and U1707 (N_1707,N_1660,N_1642);
and U1708 (N_1708,N_1606,N_1653);
nor U1709 (N_1709,N_1628,N_1696);
xnor U1710 (N_1710,N_1679,N_1662);
or U1711 (N_1711,N_1670,N_1600);
and U1712 (N_1712,N_1686,N_1631);
nor U1713 (N_1713,N_1674,N_1609);
nor U1714 (N_1714,N_1699,N_1618);
nand U1715 (N_1715,N_1685,N_1610);
and U1716 (N_1716,N_1634,N_1629);
nand U1717 (N_1717,N_1627,N_1655);
nand U1718 (N_1718,N_1692,N_1636);
or U1719 (N_1719,N_1601,N_1615);
nor U1720 (N_1720,N_1666,N_1690);
or U1721 (N_1721,N_1652,N_1604);
nand U1722 (N_1722,N_1640,N_1668);
or U1723 (N_1723,N_1639,N_1641);
or U1724 (N_1724,N_1648,N_1683);
or U1725 (N_1725,N_1680,N_1616);
or U1726 (N_1726,N_1632,N_1693);
or U1727 (N_1727,N_1654,N_1676);
and U1728 (N_1728,N_1667,N_1664);
nor U1729 (N_1729,N_1647,N_1658);
nand U1730 (N_1730,N_1659,N_1621);
nand U1731 (N_1731,N_1671,N_1607);
and U1732 (N_1732,N_1638,N_1620);
nor U1733 (N_1733,N_1643,N_1669);
or U1734 (N_1734,N_1695,N_1675);
or U1735 (N_1735,N_1644,N_1614);
nand U1736 (N_1736,N_1602,N_1681);
nand U1737 (N_1737,N_1635,N_1612);
nor U1738 (N_1738,N_1698,N_1603);
nand U1739 (N_1739,N_1611,N_1646);
and U1740 (N_1740,N_1608,N_1630);
or U1741 (N_1741,N_1625,N_1619);
and U1742 (N_1742,N_1677,N_1622);
nor U1743 (N_1743,N_1672,N_1678);
or U1744 (N_1744,N_1687,N_1624);
nor U1745 (N_1745,N_1673,N_1645);
or U1746 (N_1746,N_1633,N_1665);
and U1747 (N_1747,N_1637,N_1613);
and U1748 (N_1748,N_1663,N_1684);
nand U1749 (N_1749,N_1688,N_1657);
and U1750 (N_1750,N_1684,N_1675);
nor U1751 (N_1751,N_1673,N_1657);
nand U1752 (N_1752,N_1694,N_1655);
and U1753 (N_1753,N_1645,N_1613);
or U1754 (N_1754,N_1611,N_1632);
nor U1755 (N_1755,N_1626,N_1638);
or U1756 (N_1756,N_1677,N_1667);
nor U1757 (N_1757,N_1697,N_1686);
or U1758 (N_1758,N_1605,N_1690);
or U1759 (N_1759,N_1603,N_1651);
or U1760 (N_1760,N_1613,N_1607);
xor U1761 (N_1761,N_1615,N_1695);
or U1762 (N_1762,N_1614,N_1610);
nor U1763 (N_1763,N_1619,N_1680);
nor U1764 (N_1764,N_1605,N_1697);
and U1765 (N_1765,N_1697,N_1644);
and U1766 (N_1766,N_1624,N_1691);
and U1767 (N_1767,N_1693,N_1628);
nor U1768 (N_1768,N_1609,N_1686);
and U1769 (N_1769,N_1650,N_1672);
nor U1770 (N_1770,N_1699,N_1695);
and U1771 (N_1771,N_1686,N_1622);
nor U1772 (N_1772,N_1661,N_1618);
nand U1773 (N_1773,N_1663,N_1620);
nand U1774 (N_1774,N_1649,N_1627);
nor U1775 (N_1775,N_1662,N_1649);
or U1776 (N_1776,N_1617,N_1693);
and U1777 (N_1777,N_1680,N_1675);
or U1778 (N_1778,N_1676,N_1606);
nand U1779 (N_1779,N_1649,N_1685);
nor U1780 (N_1780,N_1654,N_1664);
nor U1781 (N_1781,N_1648,N_1604);
nor U1782 (N_1782,N_1600,N_1673);
nand U1783 (N_1783,N_1659,N_1699);
nor U1784 (N_1784,N_1606,N_1654);
or U1785 (N_1785,N_1660,N_1662);
and U1786 (N_1786,N_1635,N_1662);
nand U1787 (N_1787,N_1668,N_1610);
nor U1788 (N_1788,N_1696,N_1691);
nand U1789 (N_1789,N_1621,N_1675);
and U1790 (N_1790,N_1670,N_1682);
or U1791 (N_1791,N_1671,N_1697);
nor U1792 (N_1792,N_1607,N_1644);
nand U1793 (N_1793,N_1668,N_1608);
nand U1794 (N_1794,N_1673,N_1601);
nand U1795 (N_1795,N_1690,N_1669);
or U1796 (N_1796,N_1692,N_1679);
nor U1797 (N_1797,N_1658,N_1666);
and U1798 (N_1798,N_1604,N_1684);
nor U1799 (N_1799,N_1655,N_1638);
nor U1800 (N_1800,N_1762,N_1722);
nor U1801 (N_1801,N_1753,N_1710);
nand U1802 (N_1802,N_1795,N_1781);
nand U1803 (N_1803,N_1770,N_1771);
and U1804 (N_1804,N_1767,N_1765);
and U1805 (N_1805,N_1769,N_1721);
and U1806 (N_1806,N_1768,N_1782);
and U1807 (N_1807,N_1793,N_1760);
and U1808 (N_1808,N_1706,N_1751);
nand U1809 (N_1809,N_1764,N_1754);
nand U1810 (N_1810,N_1750,N_1776);
nand U1811 (N_1811,N_1728,N_1787);
and U1812 (N_1812,N_1733,N_1743);
nand U1813 (N_1813,N_1708,N_1734);
nor U1814 (N_1814,N_1752,N_1718);
nand U1815 (N_1815,N_1703,N_1746);
or U1816 (N_1816,N_1784,N_1786);
and U1817 (N_1817,N_1789,N_1796);
nor U1818 (N_1818,N_1727,N_1731);
nand U1819 (N_1819,N_1741,N_1779);
and U1820 (N_1820,N_1740,N_1723);
and U1821 (N_1821,N_1792,N_1724);
nand U1822 (N_1822,N_1716,N_1713);
nand U1823 (N_1823,N_1707,N_1702);
and U1824 (N_1824,N_1778,N_1739);
nor U1825 (N_1825,N_1732,N_1711);
nor U1826 (N_1826,N_1730,N_1748);
nand U1827 (N_1827,N_1761,N_1749);
nor U1828 (N_1828,N_1799,N_1783);
or U1829 (N_1829,N_1775,N_1766);
and U1830 (N_1830,N_1705,N_1700);
or U1831 (N_1831,N_1758,N_1704);
or U1832 (N_1832,N_1709,N_1719);
and U1833 (N_1833,N_1735,N_1797);
nor U1834 (N_1834,N_1747,N_1772);
and U1835 (N_1835,N_1745,N_1798);
or U1836 (N_1836,N_1737,N_1744);
nand U1837 (N_1837,N_1780,N_1788);
or U1838 (N_1838,N_1791,N_1763);
nand U1839 (N_1839,N_1726,N_1773);
nor U1840 (N_1840,N_1714,N_1715);
and U1841 (N_1841,N_1712,N_1759);
and U1842 (N_1842,N_1794,N_1785);
and U1843 (N_1843,N_1738,N_1756);
and U1844 (N_1844,N_1777,N_1720);
or U1845 (N_1845,N_1725,N_1736);
and U1846 (N_1846,N_1790,N_1774);
nor U1847 (N_1847,N_1717,N_1755);
and U1848 (N_1848,N_1729,N_1701);
xnor U1849 (N_1849,N_1757,N_1742);
nand U1850 (N_1850,N_1729,N_1736);
nor U1851 (N_1851,N_1711,N_1722);
and U1852 (N_1852,N_1741,N_1785);
nand U1853 (N_1853,N_1738,N_1764);
nand U1854 (N_1854,N_1750,N_1783);
nand U1855 (N_1855,N_1710,N_1711);
nand U1856 (N_1856,N_1711,N_1733);
or U1857 (N_1857,N_1727,N_1769);
or U1858 (N_1858,N_1768,N_1798);
nor U1859 (N_1859,N_1796,N_1758);
nor U1860 (N_1860,N_1711,N_1764);
nand U1861 (N_1861,N_1763,N_1727);
and U1862 (N_1862,N_1754,N_1761);
nor U1863 (N_1863,N_1736,N_1717);
and U1864 (N_1864,N_1737,N_1726);
nor U1865 (N_1865,N_1728,N_1704);
or U1866 (N_1866,N_1704,N_1742);
or U1867 (N_1867,N_1781,N_1717);
or U1868 (N_1868,N_1766,N_1713);
xor U1869 (N_1869,N_1739,N_1763);
or U1870 (N_1870,N_1719,N_1720);
and U1871 (N_1871,N_1716,N_1718);
nand U1872 (N_1872,N_1792,N_1710);
nor U1873 (N_1873,N_1761,N_1785);
or U1874 (N_1874,N_1717,N_1763);
nand U1875 (N_1875,N_1797,N_1745);
nand U1876 (N_1876,N_1774,N_1766);
nand U1877 (N_1877,N_1709,N_1770);
or U1878 (N_1878,N_1770,N_1768);
and U1879 (N_1879,N_1799,N_1718);
and U1880 (N_1880,N_1768,N_1755);
and U1881 (N_1881,N_1748,N_1779);
nand U1882 (N_1882,N_1722,N_1725);
nand U1883 (N_1883,N_1769,N_1722);
nor U1884 (N_1884,N_1748,N_1782);
and U1885 (N_1885,N_1795,N_1729);
nor U1886 (N_1886,N_1755,N_1789);
nand U1887 (N_1887,N_1713,N_1733);
and U1888 (N_1888,N_1778,N_1788);
nand U1889 (N_1889,N_1722,N_1764);
or U1890 (N_1890,N_1797,N_1714);
nand U1891 (N_1891,N_1783,N_1716);
or U1892 (N_1892,N_1736,N_1706);
nor U1893 (N_1893,N_1767,N_1701);
nor U1894 (N_1894,N_1716,N_1749);
nor U1895 (N_1895,N_1769,N_1701);
nor U1896 (N_1896,N_1781,N_1789);
nand U1897 (N_1897,N_1793,N_1710);
and U1898 (N_1898,N_1748,N_1750);
nand U1899 (N_1899,N_1755,N_1745);
or U1900 (N_1900,N_1827,N_1850);
or U1901 (N_1901,N_1885,N_1819);
and U1902 (N_1902,N_1846,N_1876);
or U1903 (N_1903,N_1899,N_1849);
or U1904 (N_1904,N_1825,N_1894);
and U1905 (N_1905,N_1816,N_1860);
nand U1906 (N_1906,N_1802,N_1869);
and U1907 (N_1907,N_1809,N_1810);
or U1908 (N_1908,N_1853,N_1844);
and U1909 (N_1909,N_1858,N_1896);
nor U1910 (N_1910,N_1892,N_1866);
nand U1911 (N_1911,N_1882,N_1807);
nand U1912 (N_1912,N_1804,N_1837);
nor U1913 (N_1913,N_1891,N_1898);
and U1914 (N_1914,N_1886,N_1842);
or U1915 (N_1915,N_1887,N_1874);
nand U1916 (N_1916,N_1834,N_1867);
nor U1917 (N_1917,N_1832,N_1862);
or U1918 (N_1918,N_1868,N_1841);
nand U1919 (N_1919,N_1880,N_1871);
nand U1920 (N_1920,N_1838,N_1889);
and U1921 (N_1921,N_1839,N_1812);
nand U1922 (N_1922,N_1878,N_1830);
or U1923 (N_1923,N_1888,N_1813);
or U1924 (N_1924,N_1847,N_1895);
and U1925 (N_1925,N_1826,N_1861);
and U1926 (N_1926,N_1836,N_1856);
nor U1927 (N_1927,N_1835,N_1873);
nor U1928 (N_1928,N_1877,N_1852);
and U1929 (N_1929,N_1855,N_1884);
nand U1930 (N_1930,N_1821,N_1863);
nor U1931 (N_1931,N_1875,N_1801);
or U1932 (N_1932,N_1859,N_1897);
or U1933 (N_1933,N_1800,N_1851);
or U1934 (N_1934,N_1865,N_1811);
nor U1935 (N_1935,N_1833,N_1824);
nand U1936 (N_1936,N_1808,N_1870);
and U1937 (N_1937,N_1848,N_1840);
and U1938 (N_1938,N_1818,N_1814);
nand U1939 (N_1939,N_1879,N_1817);
nor U1940 (N_1940,N_1890,N_1854);
nand U1941 (N_1941,N_1805,N_1843);
nor U1942 (N_1942,N_1803,N_1815);
nor U1943 (N_1943,N_1829,N_1823);
or U1944 (N_1944,N_1883,N_1872);
nand U1945 (N_1945,N_1820,N_1828);
or U1946 (N_1946,N_1831,N_1857);
or U1947 (N_1947,N_1893,N_1822);
nor U1948 (N_1948,N_1845,N_1806);
and U1949 (N_1949,N_1864,N_1881);
and U1950 (N_1950,N_1895,N_1878);
and U1951 (N_1951,N_1850,N_1867);
or U1952 (N_1952,N_1899,N_1802);
nor U1953 (N_1953,N_1884,N_1865);
nor U1954 (N_1954,N_1888,N_1894);
nand U1955 (N_1955,N_1808,N_1854);
nor U1956 (N_1956,N_1880,N_1808);
nor U1957 (N_1957,N_1850,N_1885);
nor U1958 (N_1958,N_1820,N_1886);
nor U1959 (N_1959,N_1872,N_1821);
nand U1960 (N_1960,N_1872,N_1897);
or U1961 (N_1961,N_1890,N_1885);
or U1962 (N_1962,N_1854,N_1848);
or U1963 (N_1963,N_1880,N_1848);
and U1964 (N_1964,N_1874,N_1891);
nor U1965 (N_1965,N_1837,N_1898);
and U1966 (N_1966,N_1831,N_1850);
nand U1967 (N_1967,N_1892,N_1898);
nand U1968 (N_1968,N_1803,N_1843);
and U1969 (N_1969,N_1882,N_1892);
nand U1970 (N_1970,N_1889,N_1845);
and U1971 (N_1971,N_1801,N_1871);
and U1972 (N_1972,N_1887,N_1855);
or U1973 (N_1973,N_1896,N_1816);
nor U1974 (N_1974,N_1820,N_1894);
and U1975 (N_1975,N_1895,N_1893);
nand U1976 (N_1976,N_1845,N_1833);
nand U1977 (N_1977,N_1832,N_1813);
nand U1978 (N_1978,N_1829,N_1876);
or U1979 (N_1979,N_1826,N_1863);
nand U1980 (N_1980,N_1887,N_1898);
or U1981 (N_1981,N_1891,N_1856);
nand U1982 (N_1982,N_1816,N_1807);
nand U1983 (N_1983,N_1821,N_1874);
nor U1984 (N_1984,N_1858,N_1824);
nand U1985 (N_1985,N_1883,N_1858);
or U1986 (N_1986,N_1882,N_1822);
and U1987 (N_1987,N_1847,N_1864);
nand U1988 (N_1988,N_1815,N_1847);
nand U1989 (N_1989,N_1838,N_1800);
or U1990 (N_1990,N_1894,N_1879);
nand U1991 (N_1991,N_1809,N_1846);
and U1992 (N_1992,N_1836,N_1896);
or U1993 (N_1993,N_1842,N_1884);
nand U1994 (N_1994,N_1870,N_1814);
nor U1995 (N_1995,N_1808,N_1865);
or U1996 (N_1996,N_1823,N_1830);
nand U1997 (N_1997,N_1817,N_1834);
nor U1998 (N_1998,N_1848,N_1860);
and U1999 (N_1999,N_1890,N_1894);
nand U2000 (N_2000,N_1936,N_1903);
nand U2001 (N_2001,N_1912,N_1904);
nor U2002 (N_2002,N_1984,N_1971);
nand U2003 (N_2003,N_1929,N_1902);
and U2004 (N_2004,N_1958,N_1909);
or U2005 (N_2005,N_1908,N_1963);
nand U2006 (N_2006,N_1911,N_1906);
and U2007 (N_2007,N_1942,N_1919);
nand U2008 (N_2008,N_1914,N_1989);
nand U2009 (N_2009,N_1927,N_1955);
or U2010 (N_2010,N_1994,N_1953);
nand U2011 (N_2011,N_1920,N_1925);
or U2012 (N_2012,N_1900,N_1923);
and U2013 (N_2013,N_1934,N_1937);
or U2014 (N_2014,N_1944,N_1951);
nand U2015 (N_2015,N_1907,N_1940);
nor U2016 (N_2016,N_1975,N_1967);
or U2017 (N_2017,N_1957,N_1997);
nand U2018 (N_2018,N_1924,N_1974);
or U2019 (N_2019,N_1946,N_1910);
and U2020 (N_2020,N_1948,N_1986);
and U2021 (N_2021,N_1970,N_1996);
or U2022 (N_2022,N_1964,N_1983);
nor U2023 (N_2023,N_1995,N_1941);
and U2024 (N_2024,N_1965,N_1998);
and U2025 (N_2025,N_1999,N_1933);
and U2026 (N_2026,N_1921,N_1991);
and U2027 (N_2027,N_1915,N_1972);
nor U2028 (N_2028,N_1992,N_1961);
nand U2029 (N_2029,N_1930,N_1943);
xor U2030 (N_2030,N_1962,N_1959);
or U2031 (N_2031,N_1966,N_1922);
and U2032 (N_2032,N_1990,N_1932);
nor U2033 (N_2033,N_1993,N_1945);
nor U2034 (N_2034,N_1905,N_1952);
or U2035 (N_2035,N_1985,N_1980);
or U2036 (N_2036,N_1913,N_1960);
nor U2037 (N_2037,N_1926,N_1968);
and U2038 (N_2038,N_1916,N_1935);
or U2039 (N_2039,N_1981,N_1954);
or U2040 (N_2040,N_1928,N_1987);
or U2041 (N_2041,N_1939,N_1949);
or U2042 (N_2042,N_1938,N_1950);
and U2043 (N_2043,N_1982,N_1976);
or U2044 (N_2044,N_1918,N_1917);
or U2045 (N_2045,N_1973,N_1969);
nor U2046 (N_2046,N_1988,N_1901);
nand U2047 (N_2047,N_1947,N_1978);
or U2048 (N_2048,N_1977,N_1979);
or U2049 (N_2049,N_1931,N_1956);
nor U2050 (N_2050,N_1924,N_1952);
or U2051 (N_2051,N_1913,N_1978);
or U2052 (N_2052,N_1976,N_1972);
or U2053 (N_2053,N_1946,N_1998);
and U2054 (N_2054,N_1965,N_1980);
nand U2055 (N_2055,N_1987,N_1947);
nor U2056 (N_2056,N_1938,N_1969);
nand U2057 (N_2057,N_1953,N_1999);
nor U2058 (N_2058,N_1975,N_1991);
nor U2059 (N_2059,N_1998,N_1958);
nand U2060 (N_2060,N_1969,N_1958);
or U2061 (N_2061,N_1988,N_1958);
nor U2062 (N_2062,N_1986,N_1916);
nand U2063 (N_2063,N_1968,N_1976);
nor U2064 (N_2064,N_1963,N_1912);
and U2065 (N_2065,N_1994,N_1947);
nor U2066 (N_2066,N_1950,N_1990);
or U2067 (N_2067,N_1991,N_1971);
or U2068 (N_2068,N_1928,N_1986);
or U2069 (N_2069,N_1995,N_1939);
and U2070 (N_2070,N_1979,N_1936);
nand U2071 (N_2071,N_1957,N_1933);
or U2072 (N_2072,N_1943,N_1971);
and U2073 (N_2073,N_1904,N_1945);
and U2074 (N_2074,N_1988,N_1927);
nor U2075 (N_2075,N_1920,N_1934);
nand U2076 (N_2076,N_1929,N_1984);
nor U2077 (N_2077,N_1966,N_1959);
or U2078 (N_2078,N_1969,N_1919);
or U2079 (N_2079,N_1910,N_1957);
or U2080 (N_2080,N_1914,N_1957);
nand U2081 (N_2081,N_1902,N_1934);
nand U2082 (N_2082,N_1996,N_1977);
and U2083 (N_2083,N_1934,N_1988);
nand U2084 (N_2084,N_1964,N_1943);
nor U2085 (N_2085,N_1965,N_1976);
or U2086 (N_2086,N_1905,N_1942);
or U2087 (N_2087,N_1939,N_1948);
or U2088 (N_2088,N_1947,N_1983);
and U2089 (N_2089,N_1900,N_1904);
and U2090 (N_2090,N_1996,N_1948);
nand U2091 (N_2091,N_1916,N_1978);
nor U2092 (N_2092,N_1957,N_1994);
nand U2093 (N_2093,N_1983,N_1926);
and U2094 (N_2094,N_1952,N_1969);
nand U2095 (N_2095,N_1901,N_1983);
or U2096 (N_2096,N_1959,N_1905);
nand U2097 (N_2097,N_1948,N_1930);
and U2098 (N_2098,N_1948,N_1951);
nor U2099 (N_2099,N_1989,N_1977);
or U2100 (N_2100,N_2007,N_2029);
or U2101 (N_2101,N_2004,N_2018);
or U2102 (N_2102,N_2008,N_2022);
nand U2103 (N_2103,N_2047,N_2044);
nand U2104 (N_2104,N_2003,N_2011);
or U2105 (N_2105,N_2091,N_2060);
nand U2106 (N_2106,N_2016,N_2028);
nor U2107 (N_2107,N_2039,N_2059);
nand U2108 (N_2108,N_2079,N_2077);
nand U2109 (N_2109,N_2019,N_2048);
xnor U2110 (N_2110,N_2055,N_2010);
and U2111 (N_2111,N_2057,N_2051);
nand U2112 (N_2112,N_2025,N_2001);
nor U2113 (N_2113,N_2075,N_2081);
or U2114 (N_2114,N_2084,N_2023);
nor U2115 (N_2115,N_2046,N_2072);
and U2116 (N_2116,N_2020,N_2017);
nand U2117 (N_2117,N_2089,N_2099);
nand U2118 (N_2118,N_2096,N_2033);
nand U2119 (N_2119,N_2086,N_2093);
and U2120 (N_2120,N_2066,N_2095);
nand U2121 (N_2121,N_2024,N_2054);
nand U2122 (N_2122,N_2002,N_2034);
or U2123 (N_2123,N_2053,N_2082);
or U2124 (N_2124,N_2026,N_2042);
and U2125 (N_2125,N_2049,N_2040);
nor U2126 (N_2126,N_2068,N_2092);
or U2127 (N_2127,N_2071,N_2076);
or U2128 (N_2128,N_2006,N_2000);
nand U2129 (N_2129,N_2061,N_2045);
or U2130 (N_2130,N_2074,N_2041);
and U2131 (N_2131,N_2043,N_2038);
nor U2132 (N_2132,N_2021,N_2064);
or U2133 (N_2133,N_2087,N_2085);
nand U2134 (N_2134,N_2094,N_2027);
nor U2135 (N_2135,N_2030,N_2088);
nand U2136 (N_2136,N_2073,N_2069);
and U2137 (N_2137,N_2098,N_2013);
and U2138 (N_2138,N_2058,N_2065);
and U2139 (N_2139,N_2009,N_2083);
nand U2140 (N_2140,N_2050,N_2031);
nor U2141 (N_2141,N_2052,N_2090);
or U2142 (N_2142,N_2036,N_2097);
nor U2143 (N_2143,N_2035,N_2005);
and U2144 (N_2144,N_2012,N_2067);
or U2145 (N_2145,N_2032,N_2015);
or U2146 (N_2146,N_2070,N_2080);
and U2147 (N_2147,N_2078,N_2014);
or U2148 (N_2148,N_2037,N_2063);
and U2149 (N_2149,N_2056,N_2062);
nor U2150 (N_2150,N_2064,N_2095);
and U2151 (N_2151,N_2077,N_2038);
nand U2152 (N_2152,N_2053,N_2028);
nand U2153 (N_2153,N_2024,N_2073);
and U2154 (N_2154,N_2008,N_2088);
nor U2155 (N_2155,N_2061,N_2006);
or U2156 (N_2156,N_2025,N_2061);
or U2157 (N_2157,N_2079,N_2056);
nand U2158 (N_2158,N_2028,N_2063);
nand U2159 (N_2159,N_2033,N_2010);
nand U2160 (N_2160,N_2060,N_2097);
and U2161 (N_2161,N_2094,N_2060);
and U2162 (N_2162,N_2000,N_2020);
or U2163 (N_2163,N_2008,N_2089);
nand U2164 (N_2164,N_2080,N_2082);
or U2165 (N_2165,N_2094,N_2005);
or U2166 (N_2166,N_2014,N_2039);
and U2167 (N_2167,N_2054,N_2073);
nor U2168 (N_2168,N_2048,N_2067);
or U2169 (N_2169,N_2018,N_2095);
nor U2170 (N_2170,N_2027,N_2018);
or U2171 (N_2171,N_2079,N_2075);
nor U2172 (N_2172,N_2057,N_2056);
nand U2173 (N_2173,N_2030,N_2011);
and U2174 (N_2174,N_2055,N_2085);
nand U2175 (N_2175,N_2065,N_2013);
or U2176 (N_2176,N_2076,N_2056);
and U2177 (N_2177,N_2032,N_2040);
or U2178 (N_2178,N_2078,N_2095);
nand U2179 (N_2179,N_2053,N_2081);
or U2180 (N_2180,N_2065,N_2076);
nor U2181 (N_2181,N_2080,N_2002);
and U2182 (N_2182,N_2081,N_2007);
and U2183 (N_2183,N_2079,N_2071);
nand U2184 (N_2184,N_2004,N_2072);
nand U2185 (N_2185,N_2090,N_2016);
or U2186 (N_2186,N_2014,N_2022);
nand U2187 (N_2187,N_2089,N_2002);
nor U2188 (N_2188,N_2019,N_2078);
nand U2189 (N_2189,N_2093,N_2095);
nor U2190 (N_2190,N_2089,N_2044);
nor U2191 (N_2191,N_2003,N_2046);
or U2192 (N_2192,N_2052,N_2020);
nand U2193 (N_2193,N_2021,N_2096);
or U2194 (N_2194,N_2095,N_2036);
and U2195 (N_2195,N_2023,N_2005);
and U2196 (N_2196,N_2001,N_2055);
and U2197 (N_2197,N_2007,N_2068);
nor U2198 (N_2198,N_2036,N_2018);
and U2199 (N_2199,N_2003,N_2071);
or U2200 (N_2200,N_2150,N_2127);
or U2201 (N_2201,N_2184,N_2129);
and U2202 (N_2202,N_2120,N_2151);
and U2203 (N_2203,N_2159,N_2142);
and U2204 (N_2204,N_2190,N_2180);
nand U2205 (N_2205,N_2105,N_2118);
nor U2206 (N_2206,N_2155,N_2146);
nor U2207 (N_2207,N_2199,N_2136);
and U2208 (N_2208,N_2109,N_2141);
xnor U2209 (N_2209,N_2167,N_2169);
nand U2210 (N_2210,N_2154,N_2137);
nand U2211 (N_2211,N_2134,N_2152);
or U2212 (N_2212,N_2124,N_2174);
or U2213 (N_2213,N_2157,N_2189);
nor U2214 (N_2214,N_2108,N_2188);
and U2215 (N_2215,N_2172,N_2158);
and U2216 (N_2216,N_2104,N_2107);
nor U2217 (N_2217,N_2133,N_2193);
nor U2218 (N_2218,N_2126,N_2183);
and U2219 (N_2219,N_2162,N_2138);
and U2220 (N_2220,N_2166,N_2194);
or U2221 (N_2221,N_2170,N_2186);
and U2222 (N_2222,N_2187,N_2149);
and U2223 (N_2223,N_2101,N_2177);
or U2224 (N_2224,N_2139,N_2128);
nor U2225 (N_2225,N_2198,N_2163);
nand U2226 (N_2226,N_2123,N_2195);
and U2227 (N_2227,N_2114,N_2112);
or U2228 (N_2228,N_2122,N_2176);
nor U2229 (N_2229,N_2147,N_2115);
and U2230 (N_2230,N_2135,N_2132);
nand U2231 (N_2231,N_2164,N_2110);
nor U2232 (N_2232,N_2140,N_2121);
nand U2233 (N_2233,N_2191,N_2111);
and U2234 (N_2234,N_2130,N_2160);
nand U2235 (N_2235,N_2145,N_2148);
and U2236 (N_2236,N_2117,N_2168);
or U2237 (N_2237,N_2178,N_2102);
or U2238 (N_2238,N_2143,N_2106);
nand U2239 (N_2239,N_2119,N_2179);
nand U2240 (N_2240,N_2175,N_2171);
nand U2241 (N_2241,N_2192,N_2196);
or U2242 (N_2242,N_2100,N_2165);
nor U2243 (N_2243,N_2173,N_2156);
and U2244 (N_2244,N_2144,N_2161);
and U2245 (N_2245,N_2182,N_2125);
nand U2246 (N_2246,N_2116,N_2103);
nand U2247 (N_2247,N_2197,N_2185);
nor U2248 (N_2248,N_2153,N_2181);
nand U2249 (N_2249,N_2131,N_2113);
and U2250 (N_2250,N_2186,N_2115);
nor U2251 (N_2251,N_2167,N_2174);
nand U2252 (N_2252,N_2103,N_2129);
and U2253 (N_2253,N_2163,N_2156);
and U2254 (N_2254,N_2162,N_2189);
or U2255 (N_2255,N_2117,N_2194);
or U2256 (N_2256,N_2181,N_2109);
or U2257 (N_2257,N_2140,N_2139);
xnor U2258 (N_2258,N_2137,N_2138);
nor U2259 (N_2259,N_2133,N_2146);
and U2260 (N_2260,N_2159,N_2189);
nand U2261 (N_2261,N_2134,N_2147);
nand U2262 (N_2262,N_2163,N_2112);
or U2263 (N_2263,N_2172,N_2162);
nor U2264 (N_2264,N_2140,N_2120);
nand U2265 (N_2265,N_2135,N_2161);
nor U2266 (N_2266,N_2149,N_2161);
and U2267 (N_2267,N_2156,N_2188);
nand U2268 (N_2268,N_2119,N_2107);
and U2269 (N_2269,N_2105,N_2169);
or U2270 (N_2270,N_2148,N_2100);
and U2271 (N_2271,N_2128,N_2154);
and U2272 (N_2272,N_2183,N_2124);
nand U2273 (N_2273,N_2182,N_2105);
or U2274 (N_2274,N_2151,N_2144);
nor U2275 (N_2275,N_2181,N_2103);
and U2276 (N_2276,N_2191,N_2190);
and U2277 (N_2277,N_2199,N_2174);
nand U2278 (N_2278,N_2190,N_2138);
nor U2279 (N_2279,N_2198,N_2102);
nand U2280 (N_2280,N_2142,N_2161);
nor U2281 (N_2281,N_2198,N_2108);
and U2282 (N_2282,N_2159,N_2158);
and U2283 (N_2283,N_2156,N_2152);
or U2284 (N_2284,N_2133,N_2139);
xor U2285 (N_2285,N_2140,N_2103);
nor U2286 (N_2286,N_2118,N_2178);
and U2287 (N_2287,N_2174,N_2114);
and U2288 (N_2288,N_2126,N_2138);
and U2289 (N_2289,N_2199,N_2147);
nor U2290 (N_2290,N_2157,N_2186);
or U2291 (N_2291,N_2185,N_2195);
or U2292 (N_2292,N_2151,N_2197);
nor U2293 (N_2293,N_2165,N_2133);
or U2294 (N_2294,N_2196,N_2169);
nor U2295 (N_2295,N_2101,N_2148);
and U2296 (N_2296,N_2118,N_2103);
nor U2297 (N_2297,N_2147,N_2191);
and U2298 (N_2298,N_2129,N_2101);
nor U2299 (N_2299,N_2186,N_2183);
nor U2300 (N_2300,N_2289,N_2261);
nor U2301 (N_2301,N_2272,N_2248);
nor U2302 (N_2302,N_2260,N_2288);
nand U2303 (N_2303,N_2268,N_2292);
nand U2304 (N_2304,N_2224,N_2209);
or U2305 (N_2305,N_2259,N_2225);
xor U2306 (N_2306,N_2204,N_2231);
and U2307 (N_2307,N_2283,N_2249);
nand U2308 (N_2308,N_2233,N_2297);
nand U2309 (N_2309,N_2230,N_2208);
and U2310 (N_2310,N_2223,N_2293);
nand U2311 (N_2311,N_2280,N_2212);
or U2312 (N_2312,N_2213,N_2250);
and U2313 (N_2313,N_2253,N_2243);
and U2314 (N_2314,N_2277,N_2242);
nor U2315 (N_2315,N_2252,N_2235);
or U2316 (N_2316,N_2274,N_2281);
and U2317 (N_2317,N_2264,N_2211);
nand U2318 (N_2318,N_2271,N_2298);
nor U2319 (N_2319,N_2227,N_2270);
or U2320 (N_2320,N_2247,N_2279);
nand U2321 (N_2321,N_2291,N_2275);
and U2322 (N_2322,N_2236,N_2202);
or U2323 (N_2323,N_2256,N_2285);
or U2324 (N_2324,N_2255,N_2206);
nand U2325 (N_2325,N_2251,N_2232);
and U2326 (N_2326,N_2215,N_2237);
nand U2327 (N_2327,N_2205,N_2296);
nor U2328 (N_2328,N_2258,N_2295);
nand U2329 (N_2329,N_2262,N_2226);
nand U2330 (N_2330,N_2220,N_2214);
or U2331 (N_2331,N_2276,N_2287);
and U2332 (N_2332,N_2239,N_2269);
nand U2333 (N_2333,N_2246,N_2265);
nand U2334 (N_2334,N_2221,N_2228);
or U2335 (N_2335,N_2241,N_2278);
or U2336 (N_2336,N_2284,N_2294);
nand U2337 (N_2337,N_2222,N_2200);
and U2338 (N_2338,N_2290,N_2229);
nand U2339 (N_2339,N_2286,N_2207);
or U2340 (N_2340,N_2234,N_2257);
nor U2341 (N_2341,N_2254,N_2299);
nor U2342 (N_2342,N_2218,N_2267);
or U2343 (N_2343,N_2201,N_2266);
and U2344 (N_2344,N_2240,N_2245);
nor U2345 (N_2345,N_2217,N_2219);
nor U2346 (N_2346,N_2210,N_2216);
nor U2347 (N_2347,N_2238,N_2263);
or U2348 (N_2348,N_2282,N_2244);
nor U2349 (N_2349,N_2273,N_2203);
nor U2350 (N_2350,N_2258,N_2294);
nor U2351 (N_2351,N_2269,N_2245);
or U2352 (N_2352,N_2274,N_2239);
or U2353 (N_2353,N_2265,N_2254);
and U2354 (N_2354,N_2237,N_2261);
and U2355 (N_2355,N_2205,N_2243);
or U2356 (N_2356,N_2233,N_2287);
or U2357 (N_2357,N_2295,N_2203);
nor U2358 (N_2358,N_2201,N_2277);
and U2359 (N_2359,N_2222,N_2226);
xor U2360 (N_2360,N_2237,N_2258);
and U2361 (N_2361,N_2201,N_2209);
and U2362 (N_2362,N_2226,N_2211);
nand U2363 (N_2363,N_2295,N_2219);
nor U2364 (N_2364,N_2206,N_2211);
nor U2365 (N_2365,N_2298,N_2276);
and U2366 (N_2366,N_2213,N_2264);
and U2367 (N_2367,N_2274,N_2242);
or U2368 (N_2368,N_2280,N_2274);
nand U2369 (N_2369,N_2216,N_2226);
and U2370 (N_2370,N_2234,N_2204);
and U2371 (N_2371,N_2208,N_2289);
nand U2372 (N_2372,N_2254,N_2200);
nand U2373 (N_2373,N_2233,N_2252);
nor U2374 (N_2374,N_2214,N_2242);
and U2375 (N_2375,N_2223,N_2212);
xor U2376 (N_2376,N_2252,N_2238);
and U2377 (N_2377,N_2220,N_2280);
and U2378 (N_2378,N_2250,N_2208);
or U2379 (N_2379,N_2205,N_2249);
nand U2380 (N_2380,N_2224,N_2241);
nor U2381 (N_2381,N_2231,N_2226);
nand U2382 (N_2382,N_2278,N_2254);
nor U2383 (N_2383,N_2205,N_2242);
or U2384 (N_2384,N_2298,N_2245);
or U2385 (N_2385,N_2225,N_2212);
or U2386 (N_2386,N_2219,N_2260);
or U2387 (N_2387,N_2260,N_2252);
nor U2388 (N_2388,N_2283,N_2267);
nor U2389 (N_2389,N_2299,N_2236);
and U2390 (N_2390,N_2282,N_2277);
nor U2391 (N_2391,N_2294,N_2268);
nor U2392 (N_2392,N_2230,N_2268);
or U2393 (N_2393,N_2271,N_2268);
nor U2394 (N_2394,N_2210,N_2247);
nor U2395 (N_2395,N_2214,N_2276);
nor U2396 (N_2396,N_2235,N_2201);
nor U2397 (N_2397,N_2268,N_2213);
or U2398 (N_2398,N_2239,N_2266);
nor U2399 (N_2399,N_2231,N_2291);
nand U2400 (N_2400,N_2331,N_2333);
nor U2401 (N_2401,N_2345,N_2318);
nand U2402 (N_2402,N_2387,N_2395);
or U2403 (N_2403,N_2366,N_2334);
nor U2404 (N_2404,N_2390,N_2356);
nor U2405 (N_2405,N_2327,N_2321);
nor U2406 (N_2406,N_2379,N_2351);
and U2407 (N_2407,N_2363,N_2368);
and U2408 (N_2408,N_2360,N_2330);
or U2409 (N_2409,N_2341,N_2310);
or U2410 (N_2410,N_2306,N_2309);
nand U2411 (N_2411,N_2324,N_2373);
nor U2412 (N_2412,N_2393,N_2343);
and U2413 (N_2413,N_2301,N_2399);
or U2414 (N_2414,N_2388,N_2339);
and U2415 (N_2415,N_2349,N_2305);
nor U2416 (N_2416,N_2348,N_2340);
and U2417 (N_2417,N_2374,N_2385);
or U2418 (N_2418,N_2326,N_2347);
nor U2419 (N_2419,N_2365,N_2323);
nor U2420 (N_2420,N_2382,N_2378);
nand U2421 (N_2421,N_2342,N_2370);
or U2422 (N_2422,N_2376,N_2308);
nor U2423 (N_2423,N_2352,N_2302);
nor U2424 (N_2424,N_2383,N_2337);
nand U2425 (N_2425,N_2335,N_2317);
nand U2426 (N_2426,N_2367,N_2307);
nor U2427 (N_2427,N_2358,N_2344);
nand U2428 (N_2428,N_2396,N_2329);
nand U2429 (N_2429,N_2369,N_2338);
nor U2430 (N_2430,N_2353,N_2386);
nand U2431 (N_2431,N_2394,N_2355);
and U2432 (N_2432,N_2313,N_2314);
and U2433 (N_2433,N_2357,N_2371);
and U2434 (N_2434,N_2304,N_2380);
nand U2435 (N_2435,N_2397,N_2325);
nor U2436 (N_2436,N_2361,N_2336);
and U2437 (N_2437,N_2372,N_2384);
nor U2438 (N_2438,N_2303,N_2375);
and U2439 (N_2439,N_2350,N_2398);
nor U2440 (N_2440,N_2315,N_2377);
or U2441 (N_2441,N_2312,N_2359);
and U2442 (N_2442,N_2316,N_2362);
and U2443 (N_2443,N_2311,N_2354);
nor U2444 (N_2444,N_2364,N_2389);
nand U2445 (N_2445,N_2319,N_2328);
and U2446 (N_2446,N_2381,N_2322);
nor U2447 (N_2447,N_2391,N_2332);
nand U2448 (N_2448,N_2300,N_2392);
nand U2449 (N_2449,N_2320,N_2346);
and U2450 (N_2450,N_2310,N_2364);
nor U2451 (N_2451,N_2372,N_2390);
nor U2452 (N_2452,N_2318,N_2304);
nor U2453 (N_2453,N_2300,N_2384);
nor U2454 (N_2454,N_2330,N_2356);
nor U2455 (N_2455,N_2395,N_2386);
xor U2456 (N_2456,N_2381,N_2353);
nand U2457 (N_2457,N_2319,N_2353);
or U2458 (N_2458,N_2352,N_2356);
nand U2459 (N_2459,N_2365,N_2364);
nor U2460 (N_2460,N_2387,N_2339);
nor U2461 (N_2461,N_2377,N_2347);
and U2462 (N_2462,N_2341,N_2354);
nand U2463 (N_2463,N_2397,N_2386);
or U2464 (N_2464,N_2338,N_2337);
nor U2465 (N_2465,N_2392,N_2321);
nand U2466 (N_2466,N_2325,N_2348);
nand U2467 (N_2467,N_2301,N_2316);
nand U2468 (N_2468,N_2354,N_2330);
or U2469 (N_2469,N_2301,N_2318);
nor U2470 (N_2470,N_2386,N_2375);
and U2471 (N_2471,N_2359,N_2398);
or U2472 (N_2472,N_2362,N_2365);
nor U2473 (N_2473,N_2328,N_2398);
and U2474 (N_2474,N_2333,N_2334);
or U2475 (N_2475,N_2315,N_2347);
nor U2476 (N_2476,N_2301,N_2375);
or U2477 (N_2477,N_2385,N_2311);
or U2478 (N_2478,N_2346,N_2336);
nand U2479 (N_2479,N_2386,N_2333);
or U2480 (N_2480,N_2326,N_2325);
nand U2481 (N_2481,N_2310,N_2378);
and U2482 (N_2482,N_2332,N_2371);
nor U2483 (N_2483,N_2339,N_2360);
and U2484 (N_2484,N_2354,N_2378);
nor U2485 (N_2485,N_2350,N_2328);
or U2486 (N_2486,N_2319,N_2306);
nor U2487 (N_2487,N_2349,N_2343);
or U2488 (N_2488,N_2355,N_2331);
and U2489 (N_2489,N_2331,N_2300);
and U2490 (N_2490,N_2326,N_2382);
nor U2491 (N_2491,N_2341,N_2398);
nand U2492 (N_2492,N_2392,N_2361);
or U2493 (N_2493,N_2309,N_2316);
or U2494 (N_2494,N_2349,N_2348);
nor U2495 (N_2495,N_2395,N_2318);
nand U2496 (N_2496,N_2324,N_2338);
and U2497 (N_2497,N_2381,N_2331);
nand U2498 (N_2498,N_2314,N_2315);
nand U2499 (N_2499,N_2331,N_2323);
or U2500 (N_2500,N_2459,N_2403);
or U2501 (N_2501,N_2493,N_2407);
nor U2502 (N_2502,N_2415,N_2451);
or U2503 (N_2503,N_2448,N_2409);
xor U2504 (N_2504,N_2436,N_2410);
nor U2505 (N_2505,N_2430,N_2425);
nand U2506 (N_2506,N_2457,N_2440);
nor U2507 (N_2507,N_2414,N_2439);
or U2508 (N_2508,N_2486,N_2472);
or U2509 (N_2509,N_2480,N_2428);
nand U2510 (N_2510,N_2438,N_2456);
or U2511 (N_2511,N_2490,N_2495);
and U2512 (N_2512,N_2467,N_2421);
nor U2513 (N_2513,N_2411,N_2482);
nand U2514 (N_2514,N_2468,N_2460);
or U2515 (N_2515,N_2427,N_2449);
nand U2516 (N_2516,N_2412,N_2406);
or U2517 (N_2517,N_2432,N_2494);
nor U2518 (N_2518,N_2470,N_2462);
or U2519 (N_2519,N_2446,N_2469);
nor U2520 (N_2520,N_2465,N_2497);
xor U2521 (N_2521,N_2496,N_2473);
nand U2522 (N_2522,N_2499,N_2492);
nor U2523 (N_2523,N_2426,N_2488);
nand U2524 (N_2524,N_2420,N_2464);
or U2525 (N_2525,N_2447,N_2404);
nand U2526 (N_2526,N_2458,N_2483);
or U2527 (N_2527,N_2408,N_2434);
and U2528 (N_2528,N_2498,N_2419);
and U2529 (N_2529,N_2423,N_2453);
nor U2530 (N_2530,N_2476,N_2444);
and U2531 (N_2531,N_2477,N_2416);
nor U2532 (N_2532,N_2429,N_2413);
and U2533 (N_2533,N_2484,N_2400);
and U2534 (N_2534,N_2475,N_2445);
or U2535 (N_2535,N_2491,N_2431);
and U2536 (N_2536,N_2437,N_2478);
and U2537 (N_2537,N_2401,N_2479);
nor U2538 (N_2538,N_2466,N_2433);
nor U2539 (N_2539,N_2463,N_2417);
and U2540 (N_2540,N_2442,N_2441);
nor U2541 (N_2541,N_2461,N_2452);
and U2542 (N_2542,N_2474,N_2489);
and U2543 (N_2543,N_2450,N_2402);
nand U2544 (N_2544,N_2422,N_2418);
and U2545 (N_2545,N_2443,N_2471);
nand U2546 (N_2546,N_2405,N_2485);
and U2547 (N_2547,N_2481,N_2424);
and U2548 (N_2548,N_2454,N_2487);
or U2549 (N_2549,N_2455,N_2435);
and U2550 (N_2550,N_2474,N_2478);
or U2551 (N_2551,N_2494,N_2418);
and U2552 (N_2552,N_2470,N_2410);
or U2553 (N_2553,N_2471,N_2425);
nand U2554 (N_2554,N_2457,N_2481);
and U2555 (N_2555,N_2436,N_2453);
nand U2556 (N_2556,N_2497,N_2410);
or U2557 (N_2557,N_2453,N_2487);
nand U2558 (N_2558,N_2432,N_2423);
or U2559 (N_2559,N_2431,N_2446);
nor U2560 (N_2560,N_2406,N_2455);
nor U2561 (N_2561,N_2452,N_2437);
and U2562 (N_2562,N_2429,N_2495);
and U2563 (N_2563,N_2483,N_2449);
xnor U2564 (N_2564,N_2493,N_2450);
and U2565 (N_2565,N_2459,N_2497);
nor U2566 (N_2566,N_2415,N_2414);
nor U2567 (N_2567,N_2481,N_2468);
or U2568 (N_2568,N_2465,N_2436);
nand U2569 (N_2569,N_2475,N_2419);
and U2570 (N_2570,N_2469,N_2497);
or U2571 (N_2571,N_2453,N_2430);
xnor U2572 (N_2572,N_2474,N_2436);
nor U2573 (N_2573,N_2411,N_2495);
nor U2574 (N_2574,N_2438,N_2421);
and U2575 (N_2575,N_2496,N_2478);
or U2576 (N_2576,N_2428,N_2473);
or U2577 (N_2577,N_2461,N_2421);
or U2578 (N_2578,N_2458,N_2476);
nor U2579 (N_2579,N_2428,N_2403);
nand U2580 (N_2580,N_2415,N_2412);
nand U2581 (N_2581,N_2422,N_2434);
nand U2582 (N_2582,N_2443,N_2499);
or U2583 (N_2583,N_2462,N_2404);
and U2584 (N_2584,N_2441,N_2447);
or U2585 (N_2585,N_2467,N_2420);
nor U2586 (N_2586,N_2481,N_2408);
nor U2587 (N_2587,N_2431,N_2424);
nor U2588 (N_2588,N_2482,N_2496);
and U2589 (N_2589,N_2496,N_2464);
or U2590 (N_2590,N_2410,N_2474);
and U2591 (N_2591,N_2447,N_2475);
nand U2592 (N_2592,N_2413,N_2442);
and U2593 (N_2593,N_2468,N_2408);
nand U2594 (N_2594,N_2441,N_2472);
nand U2595 (N_2595,N_2414,N_2487);
or U2596 (N_2596,N_2409,N_2479);
or U2597 (N_2597,N_2463,N_2455);
or U2598 (N_2598,N_2473,N_2424);
nor U2599 (N_2599,N_2482,N_2452);
or U2600 (N_2600,N_2566,N_2597);
or U2601 (N_2601,N_2522,N_2599);
or U2602 (N_2602,N_2542,N_2520);
nor U2603 (N_2603,N_2554,N_2569);
or U2604 (N_2604,N_2585,N_2563);
nor U2605 (N_2605,N_2532,N_2593);
and U2606 (N_2606,N_2518,N_2571);
or U2607 (N_2607,N_2552,N_2596);
and U2608 (N_2608,N_2513,N_2515);
nor U2609 (N_2609,N_2573,N_2533);
or U2610 (N_2610,N_2519,N_2592);
nand U2611 (N_2611,N_2529,N_2583);
or U2612 (N_2612,N_2536,N_2557);
nor U2613 (N_2613,N_2523,N_2595);
or U2614 (N_2614,N_2505,N_2509);
and U2615 (N_2615,N_2579,N_2591);
nand U2616 (N_2616,N_2582,N_2551);
nor U2617 (N_2617,N_2512,N_2568);
or U2618 (N_2618,N_2545,N_2553);
nor U2619 (N_2619,N_2560,N_2503);
nand U2620 (N_2620,N_2528,N_2580);
nand U2621 (N_2621,N_2508,N_2581);
nand U2622 (N_2622,N_2500,N_2538);
nor U2623 (N_2623,N_2549,N_2548);
or U2624 (N_2624,N_2501,N_2544);
nand U2625 (N_2625,N_2562,N_2524);
or U2626 (N_2626,N_2511,N_2556);
nor U2627 (N_2627,N_2506,N_2530);
nor U2628 (N_2628,N_2577,N_2540);
and U2629 (N_2629,N_2594,N_2584);
or U2630 (N_2630,N_2575,N_2504);
or U2631 (N_2631,N_2590,N_2555);
nand U2632 (N_2632,N_2565,N_2517);
and U2633 (N_2633,N_2578,N_2537);
or U2634 (N_2634,N_2539,N_2586);
nor U2635 (N_2635,N_2527,N_2576);
nand U2636 (N_2636,N_2507,N_2550);
or U2637 (N_2637,N_2502,N_2525);
or U2638 (N_2638,N_2561,N_2574);
or U2639 (N_2639,N_2516,N_2567);
or U2640 (N_2640,N_2543,N_2514);
and U2641 (N_2641,N_2521,N_2531);
or U2642 (N_2642,N_2564,N_2547);
nor U2643 (N_2643,N_2572,N_2589);
nand U2644 (N_2644,N_2546,N_2588);
nand U2645 (N_2645,N_2526,N_2598);
or U2646 (N_2646,N_2510,N_2587);
nand U2647 (N_2647,N_2534,N_2570);
and U2648 (N_2648,N_2559,N_2535);
and U2649 (N_2649,N_2541,N_2558);
nor U2650 (N_2650,N_2594,N_2548);
and U2651 (N_2651,N_2582,N_2576);
and U2652 (N_2652,N_2548,N_2571);
and U2653 (N_2653,N_2509,N_2577);
and U2654 (N_2654,N_2513,N_2503);
nor U2655 (N_2655,N_2573,N_2542);
nor U2656 (N_2656,N_2511,N_2504);
or U2657 (N_2657,N_2514,N_2558);
nor U2658 (N_2658,N_2583,N_2518);
and U2659 (N_2659,N_2571,N_2559);
nand U2660 (N_2660,N_2533,N_2524);
nand U2661 (N_2661,N_2545,N_2590);
nor U2662 (N_2662,N_2542,N_2555);
or U2663 (N_2663,N_2573,N_2582);
or U2664 (N_2664,N_2544,N_2541);
nor U2665 (N_2665,N_2555,N_2505);
and U2666 (N_2666,N_2597,N_2503);
and U2667 (N_2667,N_2501,N_2525);
or U2668 (N_2668,N_2566,N_2501);
or U2669 (N_2669,N_2548,N_2599);
nor U2670 (N_2670,N_2592,N_2504);
or U2671 (N_2671,N_2597,N_2574);
or U2672 (N_2672,N_2592,N_2530);
and U2673 (N_2673,N_2504,N_2548);
or U2674 (N_2674,N_2522,N_2564);
and U2675 (N_2675,N_2509,N_2561);
or U2676 (N_2676,N_2552,N_2516);
and U2677 (N_2677,N_2563,N_2541);
and U2678 (N_2678,N_2569,N_2505);
nand U2679 (N_2679,N_2583,N_2539);
nand U2680 (N_2680,N_2589,N_2561);
and U2681 (N_2681,N_2500,N_2519);
and U2682 (N_2682,N_2580,N_2583);
nand U2683 (N_2683,N_2573,N_2577);
or U2684 (N_2684,N_2509,N_2549);
nand U2685 (N_2685,N_2558,N_2523);
or U2686 (N_2686,N_2535,N_2553);
nand U2687 (N_2687,N_2502,N_2522);
nand U2688 (N_2688,N_2518,N_2504);
and U2689 (N_2689,N_2519,N_2504);
nand U2690 (N_2690,N_2564,N_2512);
xor U2691 (N_2691,N_2565,N_2555);
nor U2692 (N_2692,N_2542,N_2524);
nand U2693 (N_2693,N_2568,N_2552);
and U2694 (N_2694,N_2589,N_2586);
nor U2695 (N_2695,N_2572,N_2579);
nor U2696 (N_2696,N_2568,N_2536);
or U2697 (N_2697,N_2598,N_2589);
nor U2698 (N_2698,N_2550,N_2563);
or U2699 (N_2699,N_2590,N_2591);
nand U2700 (N_2700,N_2602,N_2697);
nor U2701 (N_2701,N_2691,N_2696);
xnor U2702 (N_2702,N_2605,N_2655);
and U2703 (N_2703,N_2681,N_2634);
nand U2704 (N_2704,N_2695,N_2631);
nor U2705 (N_2705,N_2671,N_2693);
or U2706 (N_2706,N_2651,N_2659);
and U2707 (N_2707,N_2660,N_2606);
and U2708 (N_2708,N_2646,N_2641);
nor U2709 (N_2709,N_2652,N_2694);
and U2710 (N_2710,N_2688,N_2658);
or U2711 (N_2711,N_2630,N_2601);
or U2712 (N_2712,N_2640,N_2668);
or U2713 (N_2713,N_2686,N_2650);
or U2714 (N_2714,N_2620,N_2621);
or U2715 (N_2715,N_2679,N_2636);
or U2716 (N_2716,N_2667,N_2662);
nor U2717 (N_2717,N_2626,N_2632);
nand U2718 (N_2718,N_2666,N_2647);
nor U2719 (N_2719,N_2616,N_2683);
nor U2720 (N_2720,N_2649,N_2669);
nand U2721 (N_2721,N_2633,N_2644);
nand U2722 (N_2722,N_2675,N_2614);
and U2723 (N_2723,N_2692,N_2623);
nand U2724 (N_2724,N_2627,N_2612);
or U2725 (N_2725,N_2648,N_2653);
nor U2726 (N_2726,N_2642,N_2611);
nor U2727 (N_2727,N_2609,N_2604);
nor U2728 (N_2728,N_2628,N_2645);
and U2729 (N_2729,N_2638,N_2619);
nor U2730 (N_2730,N_2680,N_2689);
or U2731 (N_2731,N_2643,N_2656);
and U2732 (N_2732,N_2685,N_2613);
and U2733 (N_2733,N_2657,N_2622);
and U2734 (N_2734,N_2699,N_2678);
or U2735 (N_2735,N_2639,N_2654);
nand U2736 (N_2736,N_2607,N_2676);
and U2737 (N_2737,N_2603,N_2687);
or U2738 (N_2738,N_2661,N_2677);
xnor U2739 (N_2739,N_2617,N_2672);
and U2740 (N_2740,N_2608,N_2673);
nor U2741 (N_2741,N_2664,N_2698);
nor U2742 (N_2742,N_2610,N_2637);
nor U2743 (N_2743,N_2684,N_2624);
nor U2744 (N_2744,N_2615,N_2663);
or U2745 (N_2745,N_2682,N_2670);
nor U2746 (N_2746,N_2665,N_2618);
and U2747 (N_2747,N_2600,N_2629);
or U2748 (N_2748,N_2674,N_2625);
or U2749 (N_2749,N_2635,N_2690);
or U2750 (N_2750,N_2626,N_2675);
and U2751 (N_2751,N_2643,N_2611);
or U2752 (N_2752,N_2615,N_2690);
nor U2753 (N_2753,N_2647,N_2650);
or U2754 (N_2754,N_2641,N_2600);
nand U2755 (N_2755,N_2630,N_2603);
or U2756 (N_2756,N_2686,N_2693);
and U2757 (N_2757,N_2616,N_2618);
nand U2758 (N_2758,N_2630,N_2615);
nor U2759 (N_2759,N_2645,N_2607);
or U2760 (N_2760,N_2647,N_2612);
and U2761 (N_2761,N_2617,N_2600);
and U2762 (N_2762,N_2642,N_2622);
or U2763 (N_2763,N_2680,N_2696);
nor U2764 (N_2764,N_2650,N_2607);
nor U2765 (N_2765,N_2650,N_2603);
or U2766 (N_2766,N_2650,N_2657);
xnor U2767 (N_2767,N_2644,N_2626);
nor U2768 (N_2768,N_2640,N_2662);
nand U2769 (N_2769,N_2693,N_2680);
and U2770 (N_2770,N_2642,N_2636);
nand U2771 (N_2771,N_2623,N_2641);
or U2772 (N_2772,N_2692,N_2648);
nor U2773 (N_2773,N_2632,N_2649);
and U2774 (N_2774,N_2601,N_2658);
and U2775 (N_2775,N_2657,N_2687);
and U2776 (N_2776,N_2613,N_2663);
nor U2777 (N_2777,N_2611,N_2687);
and U2778 (N_2778,N_2613,N_2629);
nand U2779 (N_2779,N_2631,N_2602);
nor U2780 (N_2780,N_2662,N_2639);
and U2781 (N_2781,N_2617,N_2671);
xor U2782 (N_2782,N_2643,N_2650);
nor U2783 (N_2783,N_2607,N_2661);
or U2784 (N_2784,N_2668,N_2690);
nand U2785 (N_2785,N_2621,N_2611);
or U2786 (N_2786,N_2601,N_2681);
xor U2787 (N_2787,N_2630,N_2680);
and U2788 (N_2788,N_2623,N_2642);
nand U2789 (N_2789,N_2624,N_2660);
nand U2790 (N_2790,N_2665,N_2637);
and U2791 (N_2791,N_2614,N_2660);
and U2792 (N_2792,N_2661,N_2603);
nor U2793 (N_2793,N_2610,N_2667);
and U2794 (N_2794,N_2673,N_2631);
nand U2795 (N_2795,N_2676,N_2621);
nand U2796 (N_2796,N_2678,N_2624);
or U2797 (N_2797,N_2649,N_2670);
nor U2798 (N_2798,N_2636,N_2674);
and U2799 (N_2799,N_2615,N_2637);
and U2800 (N_2800,N_2734,N_2761);
nor U2801 (N_2801,N_2731,N_2771);
nor U2802 (N_2802,N_2756,N_2723);
or U2803 (N_2803,N_2781,N_2719);
and U2804 (N_2804,N_2728,N_2721);
nand U2805 (N_2805,N_2766,N_2789);
or U2806 (N_2806,N_2787,N_2726);
nor U2807 (N_2807,N_2782,N_2733);
nand U2808 (N_2808,N_2709,N_2745);
or U2809 (N_2809,N_2737,N_2704);
or U2810 (N_2810,N_2780,N_2739);
nand U2811 (N_2811,N_2788,N_2767);
nor U2812 (N_2812,N_2770,N_2748);
and U2813 (N_2813,N_2703,N_2779);
nand U2814 (N_2814,N_2729,N_2755);
nand U2815 (N_2815,N_2706,N_2762);
nor U2816 (N_2816,N_2778,N_2713);
nand U2817 (N_2817,N_2774,N_2792);
or U2818 (N_2818,N_2753,N_2705);
nor U2819 (N_2819,N_2783,N_2724);
and U2820 (N_2820,N_2736,N_2769);
nand U2821 (N_2821,N_2754,N_2740);
and U2822 (N_2822,N_2785,N_2711);
or U2823 (N_2823,N_2773,N_2790);
or U2824 (N_2824,N_2797,N_2795);
and U2825 (N_2825,N_2714,N_2720);
nand U2826 (N_2826,N_2730,N_2735);
nor U2827 (N_2827,N_2749,N_2799);
or U2828 (N_2828,N_2702,N_2747);
or U2829 (N_2829,N_2707,N_2765);
and U2830 (N_2830,N_2741,N_2752);
nor U2831 (N_2831,N_2722,N_2744);
and U2832 (N_2832,N_2772,N_2751);
and U2833 (N_2833,N_2718,N_2700);
nor U2834 (N_2834,N_2775,N_2738);
and U2835 (N_2835,N_2764,N_2768);
nor U2836 (N_2836,N_2716,N_2758);
and U2837 (N_2837,N_2791,N_2727);
and U2838 (N_2838,N_2708,N_2757);
nand U2839 (N_2839,N_2784,N_2712);
or U2840 (N_2840,N_2763,N_2777);
and U2841 (N_2841,N_2710,N_2786);
xor U2842 (N_2842,N_2793,N_2715);
or U2843 (N_2843,N_2794,N_2742);
nand U2844 (N_2844,N_2760,N_2732);
or U2845 (N_2845,N_2759,N_2796);
or U2846 (N_2846,N_2746,N_2750);
nor U2847 (N_2847,N_2701,N_2776);
nand U2848 (N_2848,N_2725,N_2743);
or U2849 (N_2849,N_2717,N_2798);
or U2850 (N_2850,N_2784,N_2794);
nand U2851 (N_2851,N_2785,N_2770);
nor U2852 (N_2852,N_2734,N_2779);
or U2853 (N_2853,N_2777,N_2701);
nand U2854 (N_2854,N_2742,N_2702);
and U2855 (N_2855,N_2777,N_2754);
nor U2856 (N_2856,N_2771,N_2737);
nand U2857 (N_2857,N_2746,N_2763);
nor U2858 (N_2858,N_2796,N_2729);
nor U2859 (N_2859,N_2779,N_2776);
or U2860 (N_2860,N_2757,N_2756);
nor U2861 (N_2861,N_2720,N_2737);
or U2862 (N_2862,N_2733,N_2767);
and U2863 (N_2863,N_2702,N_2736);
nor U2864 (N_2864,N_2734,N_2706);
or U2865 (N_2865,N_2739,N_2704);
and U2866 (N_2866,N_2738,N_2709);
nor U2867 (N_2867,N_2756,N_2751);
and U2868 (N_2868,N_2742,N_2736);
nor U2869 (N_2869,N_2798,N_2768);
nor U2870 (N_2870,N_2750,N_2792);
nand U2871 (N_2871,N_2724,N_2713);
and U2872 (N_2872,N_2788,N_2734);
and U2873 (N_2873,N_2754,N_2729);
nand U2874 (N_2874,N_2757,N_2767);
nand U2875 (N_2875,N_2772,N_2779);
or U2876 (N_2876,N_2749,N_2760);
and U2877 (N_2877,N_2722,N_2700);
nand U2878 (N_2878,N_2777,N_2711);
and U2879 (N_2879,N_2764,N_2792);
or U2880 (N_2880,N_2777,N_2756);
and U2881 (N_2881,N_2790,N_2737);
nand U2882 (N_2882,N_2781,N_2744);
nor U2883 (N_2883,N_2735,N_2718);
xnor U2884 (N_2884,N_2703,N_2786);
nor U2885 (N_2885,N_2772,N_2704);
nand U2886 (N_2886,N_2769,N_2771);
or U2887 (N_2887,N_2795,N_2794);
nor U2888 (N_2888,N_2756,N_2730);
nand U2889 (N_2889,N_2724,N_2791);
nand U2890 (N_2890,N_2731,N_2763);
nand U2891 (N_2891,N_2782,N_2791);
or U2892 (N_2892,N_2772,N_2797);
and U2893 (N_2893,N_2753,N_2761);
and U2894 (N_2894,N_2743,N_2788);
and U2895 (N_2895,N_2730,N_2768);
nor U2896 (N_2896,N_2720,N_2732);
and U2897 (N_2897,N_2787,N_2776);
nor U2898 (N_2898,N_2711,N_2737);
nand U2899 (N_2899,N_2767,N_2711);
nor U2900 (N_2900,N_2887,N_2863);
and U2901 (N_2901,N_2835,N_2831);
or U2902 (N_2902,N_2823,N_2867);
nand U2903 (N_2903,N_2848,N_2827);
or U2904 (N_2904,N_2860,N_2881);
or U2905 (N_2905,N_2876,N_2882);
nor U2906 (N_2906,N_2837,N_2818);
or U2907 (N_2907,N_2836,N_2806);
nand U2908 (N_2908,N_2841,N_2869);
and U2909 (N_2909,N_2898,N_2897);
nor U2910 (N_2910,N_2815,N_2850);
or U2911 (N_2911,N_2875,N_2822);
or U2912 (N_2912,N_2880,N_2840);
nand U2913 (N_2913,N_2808,N_2885);
and U2914 (N_2914,N_2899,N_2828);
nand U2915 (N_2915,N_2866,N_2892);
and U2916 (N_2916,N_2856,N_2858);
or U2917 (N_2917,N_2816,N_2834);
and U2918 (N_2918,N_2811,N_2853);
and U2919 (N_2919,N_2883,N_2855);
nor U2920 (N_2920,N_2810,N_2888);
nand U2921 (N_2921,N_2896,N_2809);
and U2922 (N_2922,N_2819,N_2894);
or U2923 (N_2923,N_2862,N_2844);
and U2924 (N_2924,N_2807,N_2801);
and U2925 (N_2925,N_2873,N_2849);
or U2926 (N_2926,N_2879,N_2890);
and U2927 (N_2927,N_2800,N_2839);
nand U2928 (N_2928,N_2846,N_2859);
or U2929 (N_2929,N_2893,N_2830);
nor U2930 (N_2930,N_2845,N_2878);
or U2931 (N_2931,N_2854,N_2826);
nor U2932 (N_2932,N_2842,N_2821);
and U2933 (N_2933,N_2864,N_2857);
nor U2934 (N_2934,N_2865,N_2891);
xor U2935 (N_2935,N_2804,N_2851);
or U2936 (N_2936,N_2877,N_2872);
nor U2937 (N_2937,N_2829,N_2884);
and U2938 (N_2938,N_2847,N_2812);
nor U2939 (N_2939,N_2833,N_2889);
or U2940 (N_2940,N_2805,N_2843);
nor U2941 (N_2941,N_2832,N_2825);
and U2942 (N_2942,N_2871,N_2868);
or U2943 (N_2943,N_2802,N_2817);
nor U2944 (N_2944,N_2838,N_2813);
nor U2945 (N_2945,N_2874,N_2895);
and U2946 (N_2946,N_2861,N_2814);
or U2947 (N_2947,N_2886,N_2820);
nor U2948 (N_2948,N_2870,N_2852);
or U2949 (N_2949,N_2824,N_2803);
nor U2950 (N_2950,N_2877,N_2807);
nor U2951 (N_2951,N_2804,N_2847);
nor U2952 (N_2952,N_2813,N_2873);
nand U2953 (N_2953,N_2891,N_2884);
or U2954 (N_2954,N_2858,N_2820);
nand U2955 (N_2955,N_2831,N_2805);
nand U2956 (N_2956,N_2822,N_2850);
or U2957 (N_2957,N_2853,N_2896);
or U2958 (N_2958,N_2830,N_2899);
nand U2959 (N_2959,N_2838,N_2867);
nand U2960 (N_2960,N_2817,N_2842);
or U2961 (N_2961,N_2818,N_2836);
or U2962 (N_2962,N_2876,N_2817);
or U2963 (N_2963,N_2897,N_2802);
or U2964 (N_2964,N_2858,N_2847);
nor U2965 (N_2965,N_2896,N_2815);
nand U2966 (N_2966,N_2807,N_2820);
or U2967 (N_2967,N_2862,N_2835);
or U2968 (N_2968,N_2817,N_2865);
and U2969 (N_2969,N_2880,N_2828);
nand U2970 (N_2970,N_2835,N_2810);
nor U2971 (N_2971,N_2898,N_2834);
or U2972 (N_2972,N_2810,N_2823);
nor U2973 (N_2973,N_2877,N_2849);
and U2974 (N_2974,N_2886,N_2882);
nor U2975 (N_2975,N_2812,N_2809);
nand U2976 (N_2976,N_2824,N_2848);
nor U2977 (N_2977,N_2837,N_2814);
or U2978 (N_2978,N_2838,N_2814);
or U2979 (N_2979,N_2859,N_2878);
nor U2980 (N_2980,N_2893,N_2805);
nor U2981 (N_2981,N_2824,N_2836);
and U2982 (N_2982,N_2854,N_2882);
nand U2983 (N_2983,N_2852,N_2811);
nand U2984 (N_2984,N_2833,N_2807);
nor U2985 (N_2985,N_2887,N_2886);
nor U2986 (N_2986,N_2836,N_2832);
nor U2987 (N_2987,N_2803,N_2863);
and U2988 (N_2988,N_2873,N_2810);
nor U2989 (N_2989,N_2804,N_2866);
and U2990 (N_2990,N_2855,N_2871);
nor U2991 (N_2991,N_2827,N_2884);
nor U2992 (N_2992,N_2891,N_2829);
nand U2993 (N_2993,N_2881,N_2889);
nor U2994 (N_2994,N_2884,N_2815);
and U2995 (N_2995,N_2824,N_2869);
and U2996 (N_2996,N_2858,N_2827);
nor U2997 (N_2997,N_2801,N_2814);
or U2998 (N_2998,N_2870,N_2821);
nor U2999 (N_2999,N_2817,N_2861);
nand UO_0 (O_0,N_2987,N_2966);
or UO_1 (O_1,N_2943,N_2910);
nand UO_2 (O_2,N_2914,N_2908);
and UO_3 (O_3,N_2948,N_2977);
and UO_4 (O_4,N_2936,N_2973);
and UO_5 (O_5,N_2985,N_2965);
and UO_6 (O_6,N_2902,N_2916);
nand UO_7 (O_7,N_2996,N_2976);
and UO_8 (O_8,N_2970,N_2992);
nand UO_9 (O_9,N_2999,N_2912);
nor UO_10 (O_10,N_2901,N_2930);
or UO_11 (O_11,N_2969,N_2991);
or UO_12 (O_12,N_2931,N_2920);
or UO_13 (O_13,N_2903,N_2941);
and UO_14 (O_14,N_2974,N_2958);
and UO_15 (O_15,N_2967,N_2993);
and UO_16 (O_16,N_2937,N_2904);
nor UO_17 (O_17,N_2907,N_2997);
and UO_18 (O_18,N_2925,N_2942);
nand UO_19 (O_19,N_2935,N_2972);
or UO_20 (O_20,N_2909,N_2954);
or UO_21 (O_21,N_2968,N_2900);
or UO_22 (O_22,N_2905,N_2949);
or UO_23 (O_23,N_2950,N_2984);
or UO_24 (O_24,N_2911,N_2951);
and UO_25 (O_25,N_2945,N_2932);
and UO_26 (O_26,N_2921,N_2981);
nand UO_27 (O_27,N_2922,N_2913);
nor UO_28 (O_28,N_2906,N_2989);
nand UO_29 (O_29,N_2947,N_2952);
nand UO_30 (O_30,N_2928,N_2923);
nand UO_31 (O_31,N_2983,N_2924);
or UO_32 (O_32,N_2938,N_2963);
or UO_33 (O_33,N_2982,N_2934);
nand UO_34 (O_34,N_2995,N_2915);
nor UO_35 (O_35,N_2918,N_2933);
or UO_36 (O_36,N_2975,N_2990);
or UO_37 (O_37,N_2956,N_2980);
nor UO_38 (O_38,N_2940,N_2917);
and UO_39 (O_39,N_2962,N_2986);
or UO_40 (O_40,N_2979,N_2961);
and UO_41 (O_41,N_2944,N_2929);
nor UO_42 (O_42,N_2971,N_2957);
or UO_43 (O_43,N_2959,N_2927);
or UO_44 (O_44,N_2994,N_2926);
nor UO_45 (O_45,N_2939,N_2955);
nor UO_46 (O_46,N_2946,N_2953);
and UO_47 (O_47,N_2919,N_2988);
or UO_48 (O_48,N_2998,N_2964);
nand UO_49 (O_49,N_2960,N_2978);
nor UO_50 (O_50,N_2936,N_2998);
nor UO_51 (O_51,N_2988,N_2926);
and UO_52 (O_52,N_2988,N_2916);
and UO_53 (O_53,N_2987,N_2939);
or UO_54 (O_54,N_2923,N_2908);
and UO_55 (O_55,N_2974,N_2944);
or UO_56 (O_56,N_2979,N_2915);
nand UO_57 (O_57,N_2915,N_2902);
and UO_58 (O_58,N_2936,N_2930);
and UO_59 (O_59,N_2937,N_2912);
nor UO_60 (O_60,N_2941,N_2925);
or UO_61 (O_61,N_2933,N_2963);
and UO_62 (O_62,N_2945,N_2948);
nor UO_63 (O_63,N_2953,N_2999);
nor UO_64 (O_64,N_2921,N_2909);
or UO_65 (O_65,N_2936,N_2993);
nor UO_66 (O_66,N_2986,N_2901);
nor UO_67 (O_67,N_2925,N_2963);
nor UO_68 (O_68,N_2999,N_2960);
and UO_69 (O_69,N_2931,N_2957);
and UO_70 (O_70,N_2943,N_2996);
or UO_71 (O_71,N_2936,N_2934);
nor UO_72 (O_72,N_2991,N_2953);
nand UO_73 (O_73,N_2965,N_2910);
or UO_74 (O_74,N_2956,N_2994);
nand UO_75 (O_75,N_2906,N_2956);
and UO_76 (O_76,N_2987,N_2986);
or UO_77 (O_77,N_2974,N_2916);
or UO_78 (O_78,N_2937,N_2936);
nand UO_79 (O_79,N_2944,N_2994);
and UO_80 (O_80,N_2920,N_2935);
and UO_81 (O_81,N_2918,N_2907);
nand UO_82 (O_82,N_2912,N_2984);
and UO_83 (O_83,N_2920,N_2977);
nor UO_84 (O_84,N_2977,N_2973);
and UO_85 (O_85,N_2975,N_2927);
and UO_86 (O_86,N_2989,N_2985);
nor UO_87 (O_87,N_2957,N_2913);
nand UO_88 (O_88,N_2948,N_2970);
or UO_89 (O_89,N_2962,N_2943);
and UO_90 (O_90,N_2901,N_2961);
or UO_91 (O_91,N_2955,N_2940);
nand UO_92 (O_92,N_2984,N_2961);
nor UO_93 (O_93,N_2932,N_2925);
and UO_94 (O_94,N_2954,N_2920);
nand UO_95 (O_95,N_2994,N_2976);
xor UO_96 (O_96,N_2970,N_2962);
nor UO_97 (O_97,N_2966,N_2914);
and UO_98 (O_98,N_2982,N_2930);
nor UO_99 (O_99,N_2975,N_2923);
and UO_100 (O_100,N_2999,N_2983);
and UO_101 (O_101,N_2937,N_2972);
nor UO_102 (O_102,N_2907,N_2963);
nand UO_103 (O_103,N_2972,N_2940);
or UO_104 (O_104,N_2914,N_2976);
nor UO_105 (O_105,N_2935,N_2971);
or UO_106 (O_106,N_2901,N_2976);
or UO_107 (O_107,N_2954,N_2928);
or UO_108 (O_108,N_2957,N_2919);
or UO_109 (O_109,N_2930,N_2925);
or UO_110 (O_110,N_2921,N_2993);
and UO_111 (O_111,N_2907,N_2965);
nand UO_112 (O_112,N_2987,N_2990);
nor UO_113 (O_113,N_2980,N_2976);
or UO_114 (O_114,N_2909,N_2981);
and UO_115 (O_115,N_2997,N_2931);
and UO_116 (O_116,N_2955,N_2977);
nor UO_117 (O_117,N_2994,N_2904);
nand UO_118 (O_118,N_2900,N_2990);
nor UO_119 (O_119,N_2906,N_2936);
nand UO_120 (O_120,N_2932,N_2910);
and UO_121 (O_121,N_2900,N_2969);
nor UO_122 (O_122,N_2947,N_2905);
nor UO_123 (O_123,N_2940,N_2902);
xnor UO_124 (O_124,N_2972,N_2992);
and UO_125 (O_125,N_2911,N_2947);
or UO_126 (O_126,N_2907,N_2913);
and UO_127 (O_127,N_2917,N_2982);
nand UO_128 (O_128,N_2950,N_2979);
nor UO_129 (O_129,N_2962,N_2917);
and UO_130 (O_130,N_2968,N_2993);
nor UO_131 (O_131,N_2995,N_2949);
and UO_132 (O_132,N_2957,N_2950);
and UO_133 (O_133,N_2911,N_2974);
or UO_134 (O_134,N_2950,N_2906);
nor UO_135 (O_135,N_2961,N_2935);
nor UO_136 (O_136,N_2909,N_2910);
and UO_137 (O_137,N_2924,N_2941);
and UO_138 (O_138,N_2975,N_2980);
and UO_139 (O_139,N_2950,N_2983);
nor UO_140 (O_140,N_2918,N_2936);
and UO_141 (O_141,N_2913,N_2959);
and UO_142 (O_142,N_2904,N_2988);
nor UO_143 (O_143,N_2959,N_2976);
nand UO_144 (O_144,N_2923,N_2993);
and UO_145 (O_145,N_2904,N_2978);
and UO_146 (O_146,N_2980,N_2910);
or UO_147 (O_147,N_2942,N_2977);
nor UO_148 (O_148,N_2973,N_2975);
or UO_149 (O_149,N_2901,N_2984);
or UO_150 (O_150,N_2946,N_2959);
nor UO_151 (O_151,N_2903,N_2958);
and UO_152 (O_152,N_2937,N_2975);
or UO_153 (O_153,N_2927,N_2968);
nor UO_154 (O_154,N_2942,N_2963);
nor UO_155 (O_155,N_2955,N_2936);
nor UO_156 (O_156,N_2948,N_2902);
nand UO_157 (O_157,N_2959,N_2948);
nor UO_158 (O_158,N_2990,N_2991);
nor UO_159 (O_159,N_2970,N_2915);
and UO_160 (O_160,N_2957,N_2917);
or UO_161 (O_161,N_2976,N_2998);
nor UO_162 (O_162,N_2941,N_2977);
nor UO_163 (O_163,N_2935,N_2965);
or UO_164 (O_164,N_2966,N_2942);
or UO_165 (O_165,N_2926,N_2925);
nor UO_166 (O_166,N_2932,N_2921);
and UO_167 (O_167,N_2959,N_2939);
nor UO_168 (O_168,N_2969,N_2990);
and UO_169 (O_169,N_2975,N_2931);
xor UO_170 (O_170,N_2984,N_2929);
nor UO_171 (O_171,N_2992,N_2931);
and UO_172 (O_172,N_2914,N_2917);
nor UO_173 (O_173,N_2944,N_2928);
nand UO_174 (O_174,N_2940,N_2997);
nand UO_175 (O_175,N_2917,N_2906);
nor UO_176 (O_176,N_2943,N_2965);
nor UO_177 (O_177,N_2938,N_2958);
nand UO_178 (O_178,N_2976,N_2921);
nor UO_179 (O_179,N_2910,N_2963);
or UO_180 (O_180,N_2957,N_2910);
nor UO_181 (O_181,N_2926,N_2972);
nand UO_182 (O_182,N_2940,N_2937);
nand UO_183 (O_183,N_2991,N_2976);
nor UO_184 (O_184,N_2978,N_2947);
nor UO_185 (O_185,N_2935,N_2948);
nor UO_186 (O_186,N_2913,N_2969);
nor UO_187 (O_187,N_2945,N_2939);
and UO_188 (O_188,N_2934,N_2962);
and UO_189 (O_189,N_2972,N_2964);
or UO_190 (O_190,N_2909,N_2984);
nand UO_191 (O_191,N_2945,N_2959);
nand UO_192 (O_192,N_2982,N_2964);
nand UO_193 (O_193,N_2924,N_2913);
nand UO_194 (O_194,N_2943,N_2952);
nand UO_195 (O_195,N_2904,N_2991);
xor UO_196 (O_196,N_2953,N_2970);
nor UO_197 (O_197,N_2955,N_2994);
or UO_198 (O_198,N_2986,N_2927);
and UO_199 (O_199,N_2998,N_2983);
and UO_200 (O_200,N_2912,N_2922);
or UO_201 (O_201,N_2920,N_2925);
and UO_202 (O_202,N_2992,N_2925);
or UO_203 (O_203,N_2956,N_2950);
nor UO_204 (O_204,N_2964,N_2930);
nand UO_205 (O_205,N_2910,N_2919);
nand UO_206 (O_206,N_2900,N_2928);
and UO_207 (O_207,N_2985,N_2981);
nand UO_208 (O_208,N_2927,N_2900);
nor UO_209 (O_209,N_2919,N_2900);
nor UO_210 (O_210,N_2911,N_2962);
nand UO_211 (O_211,N_2921,N_2968);
and UO_212 (O_212,N_2949,N_2978);
or UO_213 (O_213,N_2941,N_2946);
or UO_214 (O_214,N_2982,N_2938);
nor UO_215 (O_215,N_2956,N_2908);
or UO_216 (O_216,N_2902,N_2920);
nand UO_217 (O_217,N_2945,N_2957);
or UO_218 (O_218,N_2990,N_2992);
and UO_219 (O_219,N_2908,N_2974);
nor UO_220 (O_220,N_2961,N_2992);
nand UO_221 (O_221,N_2918,N_2986);
or UO_222 (O_222,N_2901,N_2948);
nor UO_223 (O_223,N_2963,N_2931);
or UO_224 (O_224,N_2943,N_2931);
xnor UO_225 (O_225,N_2968,N_2902);
and UO_226 (O_226,N_2963,N_2980);
and UO_227 (O_227,N_2968,N_2946);
or UO_228 (O_228,N_2968,N_2961);
nor UO_229 (O_229,N_2935,N_2950);
nor UO_230 (O_230,N_2932,N_2998);
or UO_231 (O_231,N_2905,N_2922);
or UO_232 (O_232,N_2942,N_2935);
xnor UO_233 (O_233,N_2972,N_2932);
or UO_234 (O_234,N_2954,N_2902);
nand UO_235 (O_235,N_2991,N_2977);
and UO_236 (O_236,N_2948,N_2983);
nor UO_237 (O_237,N_2915,N_2948);
and UO_238 (O_238,N_2981,N_2970);
and UO_239 (O_239,N_2916,N_2934);
or UO_240 (O_240,N_2904,N_2993);
nand UO_241 (O_241,N_2903,N_2994);
nand UO_242 (O_242,N_2912,N_2962);
nand UO_243 (O_243,N_2968,N_2944);
nand UO_244 (O_244,N_2944,N_2971);
nor UO_245 (O_245,N_2953,N_2962);
nand UO_246 (O_246,N_2966,N_2968);
nor UO_247 (O_247,N_2901,N_2903);
and UO_248 (O_248,N_2948,N_2988);
and UO_249 (O_249,N_2955,N_2929);
and UO_250 (O_250,N_2966,N_2999);
or UO_251 (O_251,N_2924,N_2994);
nand UO_252 (O_252,N_2937,N_2977);
nor UO_253 (O_253,N_2937,N_2956);
nand UO_254 (O_254,N_2976,N_2966);
nor UO_255 (O_255,N_2948,N_2929);
or UO_256 (O_256,N_2999,N_2982);
and UO_257 (O_257,N_2911,N_2941);
or UO_258 (O_258,N_2907,N_2902);
and UO_259 (O_259,N_2942,N_2980);
and UO_260 (O_260,N_2944,N_2904);
and UO_261 (O_261,N_2989,N_2954);
nand UO_262 (O_262,N_2953,N_2943);
or UO_263 (O_263,N_2955,N_2968);
or UO_264 (O_264,N_2957,N_2935);
nand UO_265 (O_265,N_2976,N_2964);
xor UO_266 (O_266,N_2938,N_2951);
nor UO_267 (O_267,N_2984,N_2974);
nand UO_268 (O_268,N_2926,N_2930);
or UO_269 (O_269,N_2978,N_2994);
and UO_270 (O_270,N_2935,N_2983);
and UO_271 (O_271,N_2934,N_2964);
and UO_272 (O_272,N_2913,N_2960);
nand UO_273 (O_273,N_2975,N_2946);
and UO_274 (O_274,N_2926,N_2981);
or UO_275 (O_275,N_2988,N_2900);
and UO_276 (O_276,N_2959,N_2909);
or UO_277 (O_277,N_2922,N_2963);
nor UO_278 (O_278,N_2906,N_2939);
or UO_279 (O_279,N_2998,N_2999);
or UO_280 (O_280,N_2913,N_2923);
nor UO_281 (O_281,N_2929,N_2911);
and UO_282 (O_282,N_2992,N_2936);
and UO_283 (O_283,N_2951,N_2925);
nand UO_284 (O_284,N_2920,N_2962);
and UO_285 (O_285,N_2917,N_2924);
or UO_286 (O_286,N_2919,N_2972);
and UO_287 (O_287,N_2904,N_2908);
or UO_288 (O_288,N_2955,N_2917);
nor UO_289 (O_289,N_2987,N_2934);
nand UO_290 (O_290,N_2941,N_2960);
nor UO_291 (O_291,N_2987,N_2973);
and UO_292 (O_292,N_2913,N_2914);
nand UO_293 (O_293,N_2981,N_2906);
nand UO_294 (O_294,N_2925,N_2918);
and UO_295 (O_295,N_2993,N_2961);
nand UO_296 (O_296,N_2984,N_2992);
and UO_297 (O_297,N_2950,N_2909);
nor UO_298 (O_298,N_2916,N_2970);
and UO_299 (O_299,N_2933,N_2917);
or UO_300 (O_300,N_2933,N_2914);
nor UO_301 (O_301,N_2997,N_2943);
and UO_302 (O_302,N_2947,N_2907);
or UO_303 (O_303,N_2989,N_2915);
nor UO_304 (O_304,N_2900,N_2972);
nor UO_305 (O_305,N_2975,N_2944);
or UO_306 (O_306,N_2998,N_2942);
or UO_307 (O_307,N_2991,N_2948);
nand UO_308 (O_308,N_2935,N_2990);
or UO_309 (O_309,N_2995,N_2901);
nor UO_310 (O_310,N_2938,N_2949);
nor UO_311 (O_311,N_2946,N_2982);
nor UO_312 (O_312,N_2954,N_2900);
nor UO_313 (O_313,N_2951,N_2949);
nor UO_314 (O_314,N_2973,N_2916);
nor UO_315 (O_315,N_2916,N_2924);
nand UO_316 (O_316,N_2989,N_2931);
xor UO_317 (O_317,N_2955,N_2904);
or UO_318 (O_318,N_2987,N_2918);
nand UO_319 (O_319,N_2976,N_2981);
nand UO_320 (O_320,N_2910,N_2960);
and UO_321 (O_321,N_2955,N_2945);
nand UO_322 (O_322,N_2965,N_2992);
nor UO_323 (O_323,N_2991,N_2960);
nand UO_324 (O_324,N_2932,N_2971);
and UO_325 (O_325,N_2943,N_2960);
or UO_326 (O_326,N_2990,N_2952);
or UO_327 (O_327,N_2992,N_2944);
or UO_328 (O_328,N_2928,N_2955);
and UO_329 (O_329,N_2960,N_2907);
nand UO_330 (O_330,N_2904,N_2934);
xnor UO_331 (O_331,N_2985,N_2906);
and UO_332 (O_332,N_2988,N_2930);
or UO_333 (O_333,N_2922,N_2936);
and UO_334 (O_334,N_2987,N_2948);
nand UO_335 (O_335,N_2998,N_2927);
and UO_336 (O_336,N_2917,N_2913);
nand UO_337 (O_337,N_2902,N_2910);
nand UO_338 (O_338,N_2957,N_2987);
nor UO_339 (O_339,N_2939,N_2924);
nand UO_340 (O_340,N_2957,N_2929);
nor UO_341 (O_341,N_2923,N_2932);
nor UO_342 (O_342,N_2902,N_2998);
or UO_343 (O_343,N_2916,N_2942);
nand UO_344 (O_344,N_2920,N_2981);
nor UO_345 (O_345,N_2956,N_2953);
and UO_346 (O_346,N_2960,N_2958);
or UO_347 (O_347,N_2918,N_2908);
nor UO_348 (O_348,N_2944,N_2931);
nor UO_349 (O_349,N_2975,N_2915);
or UO_350 (O_350,N_2951,N_2992);
nor UO_351 (O_351,N_2944,N_2912);
or UO_352 (O_352,N_2966,N_2932);
and UO_353 (O_353,N_2903,N_2934);
or UO_354 (O_354,N_2992,N_2926);
nand UO_355 (O_355,N_2915,N_2933);
and UO_356 (O_356,N_2929,N_2924);
nor UO_357 (O_357,N_2931,N_2936);
and UO_358 (O_358,N_2939,N_2967);
or UO_359 (O_359,N_2900,N_2936);
and UO_360 (O_360,N_2968,N_2935);
and UO_361 (O_361,N_2937,N_2982);
or UO_362 (O_362,N_2982,N_2925);
nand UO_363 (O_363,N_2916,N_2946);
and UO_364 (O_364,N_2947,N_2927);
or UO_365 (O_365,N_2988,N_2905);
and UO_366 (O_366,N_2926,N_2939);
and UO_367 (O_367,N_2943,N_2991);
and UO_368 (O_368,N_2924,N_2998);
or UO_369 (O_369,N_2982,N_2902);
and UO_370 (O_370,N_2916,N_2959);
and UO_371 (O_371,N_2949,N_2976);
nor UO_372 (O_372,N_2960,N_2939);
or UO_373 (O_373,N_2983,N_2927);
or UO_374 (O_374,N_2913,N_2990);
nand UO_375 (O_375,N_2967,N_2990);
or UO_376 (O_376,N_2968,N_2930);
or UO_377 (O_377,N_2935,N_2967);
or UO_378 (O_378,N_2985,N_2913);
xnor UO_379 (O_379,N_2981,N_2975);
or UO_380 (O_380,N_2969,N_2930);
and UO_381 (O_381,N_2943,N_2994);
nor UO_382 (O_382,N_2960,N_2912);
nand UO_383 (O_383,N_2932,N_2976);
and UO_384 (O_384,N_2926,N_2901);
nand UO_385 (O_385,N_2979,N_2959);
or UO_386 (O_386,N_2904,N_2985);
nor UO_387 (O_387,N_2987,N_2955);
nor UO_388 (O_388,N_2900,N_2942);
nand UO_389 (O_389,N_2943,N_2916);
nand UO_390 (O_390,N_2909,N_2957);
nor UO_391 (O_391,N_2923,N_2967);
nor UO_392 (O_392,N_2987,N_2999);
nor UO_393 (O_393,N_2945,N_2962);
nand UO_394 (O_394,N_2968,N_2939);
and UO_395 (O_395,N_2906,N_2922);
nor UO_396 (O_396,N_2999,N_2996);
and UO_397 (O_397,N_2939,N_2986);
and UO_398 (O_398,N_2974,N_2979);
xnor UO_399 (O_399,N_2955,N_2907);
nor UO_400 (O_400,N_2947,N_2944);
and UO_401 (O_401,N_2959,N_2949);
and UO_402 (O_402,N_2954,N_2974);
and UO_403 (O_403,N_2966,N_2929);
and UO_404 (O_404,N_2946,N_2924);
and UO_405 (O_405,N_2989,N_2922);
nand UO_406 (O_406,N_2974,N_2949);
nor UO_407 (O_407,N_2947,N_2923);
and UO_408 (O_408,N_2938,N_2999);
nor UO_409 (O_409,N_2981,N_2900);
and UO_410 (O_410,N_2991,N_2959);
and UO_411 (O_411,N_2945,N_2976);
xor UO_412 (O_412,N_2988,N_2956);
or UO_413 (O_413,N_2956,N_2983);
or UO_414 (O_414,N_2903,N_2912);
and UO_415 (O_415,N_2946,N_2933);
nand UO_416 (O_416,N_2953,N_2944);
nand UO_417 (O_417,N_2925,N_2965);
nor UO_418 (O_418,N_2935,N_2921);
and UO_419 (O_419,N_2940,N_2971);
or UO_420 (O_420,N_2914,N_2920);
or UO_421 (O_421,N_2938,N_2927);
nor UO_422 (O_422,N_2905,N_2917);
or UO_423 (O_423,N_2942,N_2910);
nor UO_424 (O_424,N_2900,N_2908);
and UO_425 (O_425,N_2978,N_2912);
nand UO_426 (O_426,N_2937,N_2947);
nand UO_427 (O_427,N_2966,N_2972);
or UO_428 (O_428,N_2962,N_2928);
nor UO_429 (O_429,N_2922,N_2986);
or UO_430 (O_430,N_2997,N_2993);
and UO_431 (O_431,N_2977,N_2996);
or UO_432 (O_432,N_2944,N_2906);
nand UO_433 (O_433,N_2949,N_2975);
and UO_434 (O_434,N_2982,N_2991);
and UO_435 (O_435,N_2921,N_2913);
or UO_436 (O_436,N_2975,N_2951);
and UO_437 (O_437,N_2960,N_2918);
and UO_438 (O_438,N_2939,N_2999);
or UO_439 (O_439,N_2929,N_2963);
or UO_440 (O_440,N_2964,N_2941);
and UO_441 (O_441,N_2924,N_2904);
and UO_442 (O_442,N_2916,N_2940);
nor UO_443 (O_443,N_2994,N_2951);
nor UO_444 (O_444,N_2946,N_2990);
nand UO_445 (O_445,N_2934,N_2911);
or UO_446 (O_446,N_2996,N_2964);
nand UO_447 (O_447,N_2933,N_2912);
nor UO_448 (O_448,N_2952,N_2909);
and UO_449 (O_449,N_2930,N_2966);
nor UO_450 (O_450,N_2972,N_2908);
or UO_451 (O_451,N_2946,N_2958);
nor UO_452 (O_452,N_2992,N_2953);
or UO_453 (O_453,N_2941,N_2962);
or UO_454 (O_454,N_2955,N_2983);
nand UO_455 (O_455,N_2935,N_2995);
and UO_456 (O_456,N_2998,N_2904);
or UO_457 (O_457,N_2926,N_2978);
nor UO_458 (O_458,N_2974,N_2918);
nand UO_459 (O_459,N_2906,N_2977);
or UO_460 (O_460,N_2994,N_2934);
nor UO_461 (O_461,N_2987,N_2994);
or UO_462 (O_462,N_2920,N_2973);
or UO_463 (O_463,N_2943,N_2993);
or UO_464 (O_464,N_2912,N_2917);
nor UO_465 (O_465,N_2973,N_2934);
or UO_466 (O_466,N_2904,N_2987);
xor UO_467 (O_467,N_2950,N_2943);
nand UO_468 (O_468,N_2939,N_2923);
or UO_469 (O_469,N_2940,N_2911);
nand UO_470 (O_470,N_2915,N_2957);
nor UO_471 (O_471,N_2966,N_2997);
or UO_472 (O_472,N_2976,N_2926);
and UO_473 (O_473,N_2963,N_2941);
or UO_474 (O_474,N_2930,N_2975);
nor UO_475 (O_475,N_2943,N_2905);
and UO_476 (O_476,N_2914,N_2961);
nor UO_477 (O_477,N_2968,N_2947);
nand UO_478 (O_478,N_2907,N_2904);
nor UO_479 (O_479,N_2998,N_2920);
or UO_480 (O_480,N_2971,N_2978);
and UO_481 (O_481,N_2922,N_2923);
nand UO_482 (O_482,N_2911,N_2978);
nand UO_483 (O_483,N_2981,N_2998);
nand UO_484 (O_484,N_2993,N_2929);
nand UO_485 (O_485,N_2991,N_2905);
nand UO_486 (O_486,N_2904,N_2932);
nand UO_487 (O_487,N_2995,N_2980);
nor UO_488 (O_488,N_2920,N_2911);
nor UO_489 (O_489,N_2924,N_2961);
or UO_490 (O_490,N_2946,N_2986);
nor UO_491 (O_491,N_2995,N_2997);
nand UO_492 (O_492,N_2971,N_2921);
nand UO_493 (O_493,N_2975,N_2943);
or UO_494 (O_494,N_2953,N_2915);
or UO_495 (O_495,N_2915,N_2913);
and UO_496 (O_496,N_2928,N_2991);
or UO_497 (O_497,N_2973,N_2942);
or UO_498 (O_498,N_2951,N_2963);
or UO_499 (O_499,N_2913,N_2929);
endmodule