module basic_2500_25000_3000_4_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18772,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18990,N_18991,N_18992,N_18993,N_18994,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19174,N_19176,N_19177,N_19178,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19378,N_19379,N_19380,N_19381,N_19382,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19668,N_19670,N_19671,N_19672,N_19673,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19880,N_19881,N_19882,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20038,N_20039,N_20040,N_20041,N_20042,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20249,N_20250,N_20251,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20457,N_20458,N_20459,N_20460,N_20461,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20506,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20537,N_20538,N_20540,N_20541,N_20542,N_20543,N_20544,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20582,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20713,N_20714,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20747,N_20748,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21383,N_21384,N_21385,N_21386,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21705,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21854,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22001,N_22002,N_22003,N_22004,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22156,N_22157,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22225,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22403,N_22404,N_22405,N_22406,N_22407,N_22409,N_22410,N_22411,N_22412,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22759,N_22760,N_22761,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22998,N_22999,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23184,N_23185,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23378,N_23379,N_23381,N_23382,N_23383,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23537,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23578,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23636,N_23637,N_23638,N_23639,N_23640,N_23642,N_23643,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23800,N_23801,N_23802,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23895,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24159,N_24160,N_24161,N_24162,N_24163,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24328,N_24329,N_24330,N_24331,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24374,N_24375,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24480,N_24481,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24541,N_24542,N_24543,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_835,In_1704);
nand U1 (N_1,In_1731,In_2079);
nand U2 (N_2,In_1734,In_285);
and U3 (N_3,In_2363,In_2110);
xnor U4 (N_4,In_1653,In_1745);
xor U5 (N_5,In_1730,In_920);
nand U6 (N_6,In_785,In_1167);
nor U7 (N_7,In_563,In_1763);
or U8 (N_8,In_1508,In_1794);
xor U9 (N_9,In_2217,In_1785);
nand U10 (N_10,In_2207,In_196);
or U11 (N_11,In_1275,In_152);
or U12 (N_12,In_1257,In_1598);
and U13 (N_13,In_2286,In_259);
nand U14 (N_14,In_654,In_1907);
nor U15 (N_15,In_1185,In_1437);
xor U16 (N_16,In_990,In_1507);
xor U17 (N_17,In_2461,In_1778);
xor U18 (N_18,In_1912,In_2174);
or U19 (N_19,In_1897,In_967);
nand U20 (N_20,In_2230,In_72);
and U21 (N_21,In_1203,In_1925);
and U22 (N_22,In_2308,In_959);
nand U23 (N_23,In_495,In_1408);
and U24 (N_24,In_1069,In_870);
nand U25 (N_25,In_614,In_104);
xnor U26 (N_26,In_1736,In_1890);
and U27 (N_27,In_481,In_483);
xor U28 (N_28,In_1122,In_406);
xnor U29 (N_29,In_637,In_1909);
nor U30 (N_30,In_162,In_305);
and U31 (N_31,In_701,In_743);
xnor U32 (N_32,In_1978,In_295);
and U33 (N_33,In_1087,In_274);
or U34 (N_34,In_574,In_2419);
or U35 (N_35,In_1593,In_880);
xnor U36 (N_36,In_1748,In_1093);
nor U37 (N_37,In_331,In_1461);
xor U38 (N_38,In_961,In_245);
or U39 (N_39,In_1086,In_1877);
xor U40 (N_40,In_2245,In_1921);
nand U41 (N_41,In_2172,In_474);
or U42 (N_42,In_348,In_461);
nor U43 (N_43,In_268,In_144);
nand U44 (N_44,In_2190,In_43);
and U45 (N_45,In_1563,In_1654);
nor U46 (N_46,In_1693,In_1624);
xnor U47 (N_47,In_1166,In_234);
nand U48 (N_48,In_1681,In_1644);
or U49 (N_49,In_270,In_336);
nand U50 (N_50,In_2341,In_589);
nor U51 (N_51,In_704,In_1984);
nor U52 (N_52,In_1750,In_1100);
nand U53 (N_53,In_1697,In_664);
or U54 (N_54,In_693,In_2117);
xor U55 (N_55,In_262,In_2407);
nor U56 (N_56,In_121,In_2427);
xor U57 (N_57,In_438,In_2032);
xor U58 (N_58,In_1805,In_1462);
nor U59 (N_59,In_97,In_1216);
or U60 (N_60,In_1142,In_577);
and U61 (N_61,In_1603,In_617);
and U62 (N_62,In_2350,In_1911);
and U63 (N_63,In_107,In_862);
nor U64 (N_64,In_1672,In_1245);
nand U65 (N_65,In_1885,In_827);
or U66 (N_66,In_235,In_1937);
and U67 (N_67,In_1281,In_314);
xor U68 (N_68,In_1808,In_945);
nor U69 (N_69,In_2413,In_1865);
nor U70 (N_70,In_908,In_1977);
or U71 (N_71,In_992,In_2466);
nand U72 (N_72,In_2257,In_498);
or U73 (N_73,In_1394,In_117);
nand U74 (N_74,In_685,In_404);
and U75 (N_75,In_130,In_910);
nor U76 (N_76,In_1860,In_1645);
or U77 (N_77,In_1222,In_2321);
nor U78 (N_78,In_228,In_317);
xor U79 (N_79,In_1706,In_924);
xnor U80 (N_80,In_1113,In_1218);
nand U81 (N_81,In_1756,In_1891);
nand U82 (N_82,In_2226,In_919);
and U83 (N_83,In_1555,In_1966);
and U84 (N_84,In_1533,In_89);
nor U85 (N_85,In_881,In_2189);
xnor U86 (N_86,In_1500,In_2326);
xor U87 (N_87,In_91,In_20);
nand U88 (N_88,In_853,In_2488);
or U89 (N_89,In_2459,In_1138);
xor U90 (N_90,In_713,In_2183);
nor U91 (N_91,In_2143,In_2303);
and U92 (N_92,In_35,In_534);
nor U93 (N_93,In_1813,In_973);
xor U94 (N_94,In_2178,In_1981);
nor U95 (N_95,In_2291,In_628);
nor U96 (N_96,In_918,In_1499);
and U97 (N_97,In_879,In_2288);
and U98 (N_98,In_1425,In_1414);
nor U99 (N_99,In_2154,In_1680);
or U100 (N_100,In_2273,In_576);
nor U101 (N_101,In_1006,In_640);
or U102 (N_102,In_1970,In_1411);
nand U103 (N_103,In_1579,In_1820);
nor U104 (N_104,In_1458,In_769);
nor U105 (N_105,In_1270,In_2147);
and U106 (N_106,In_750,In_1037);
nand U107 (N_107,In_118,In_1494);
nor U108 (N_108,In_2017,In_618);
and U109 (N_109,In_1530,In_29);
and U110 (N_110,In_2162,In_1392);
or U111 (N_111,In_2294,In_902);
or U112 (N_112,In_539,In_642);
xnor U113 (N_113,In_688,In_2403);
xnor U114 (N_114,In_140,In_1442);
or U115 (N_115,In_2258,In_2262);
or U116 (N_116,In_2027,In_649);
nand U117 (N_117,In_1171,In_653);
and U118 (N_118,In_1052,In_1360);
nand U119 (N_119,In_606,In_2112);
and U120 (N_120,In_559,In_1108);
nand U121 (N_121,In_321,In_209);
nand U122 (N_122,In_1557,In_570);
and U123 (N_123,In_1183,In_603);
and U124 (N_124,In_1935,In_626);
xor U125 (N_125,In_884,In_1542);
nand U126 (N_126,In_1091,In_1467);
nor U127 (N_127,In_1422,In_2149);
nor U128 (N_128,In_148,In_2345);
nor U129 (N_129,In_639,In_1673);
nand U130 (N_130,In_374,In_1141);
xnor U131 (N_131,In_1187,In_1651);
or U132 (N_132,In_1473,In_573);
nor U133 (N_133,In_981,In_2263);
nand U134 (N_134,In_761,In_877);
and U135 (N_135,In_1641,In_371);
and U136 (N_136,In_232,In_267);
or U137 (N_137,In_2397,In_2025);
xor U138 (N_138,In_1135,In_1015);
xor U139 (N_139,In_1883,In_2475);
nand U140 (N_140,In_939,In_2058);
and U141 (N_141,In_2365,In_2180);
or U142 (N_142,In_1548,In_697);
and U143 (N_143,In_656,In_825);
or U144 (N_144,In_2169,In_1861);
xnor U145 (N_145,In_1365,In_2153);
nor U146 (N_146,In_254,In_2040);
nand U147 (N_147,In_1965,In_289);
nand U148 (N_148,In_2405,In_178);
nor U149 (N_149,In_1927,In_1996);
and U150 (N_150,In_1878,In_201);
xor U151 (N_151,In_950,In_375);
and U152 (N_152,In_1544,In_857);
nor U153 (N_153,In_47,In_211);
or U154 (N_154,In_2177,In_2380);
nand U155 (N_155,In_1162,In_2465);
and U156 (N_156,In_1630,In_10);
or U157 (N_157,In_2088,In_2193);
nand U158 (N_158,In_2247,In_2196);
nand U159 (N_159,In_976,In_1549);
nor U160 (N_160,In_2367,In_1591);
or U161 (N_161,In_1249,In_2318);
xor U162 (N_162,In_968,In_1004);
and U163 (N_163,In_1008,In_1416);
and U164 (N_164,In_2469,In_1787);
and U165 (N_165,In_1482,In_1830);
nand U166 (N_166,In_2124,In_1749);
nand U167 (N_167,In_2444,In_2383);
and U168 (N_168,In_113,In_1423);
and U169 (N_169,In_2139,In_2270);
nor U170 (N_170,In_580,In_1944);
nor U171 (N_171,In_1429,In_2429);
or U172 (N_172,In_1527,In_350);
nand U173 (N_173,In_627,In_2389);
nand U174 (N_174,In_1933,In_789);
xnor U175 (N_175,In_1076,In_177);
nand U176 (N_176,In_666,In_1498);
nand U177 (N_177,In_2476,In_982);
or U178 (N_178,In_955,In_2387);
and U179 (N_179,In_93,In_548);
or U180 (N_180,In_775,In_949);
nand U181 (N_181,In_41,In_396);
and U182 (N_182,In_2198,In_830);
nor U183 (N_183,In_805,In_547);
nand U184 (N_184,In_2297,In_2472);
and U185 (N_185,In_2105,In_2379);
xor U186 (N_186,In_1248,In_2423);
xnor U187 (N_187,In_51,In_2101);
nor U188 (N_188,In_1192,In_2375);
nand U189 (N_189,In_1131,In_2075);
xnor U190 (N_190,In_1879,In_388);
nand U191 (N_191,In_528,In_2131);
nor U192 (N_192,In_2460,In_1957);
and U193 (N_193,In_1716,In_2213);
or U194 (N_194,In_736,In_1453);
and U195 (N_195,In_2235,In_979);
and U196 (N_196,In_181,In_711);
and U197 (N_197,In_1298,In_1842);
nand U198 (N_198,In_2349,In_1739);
or U199 (N_199,In_859,In_1760);
and U200 (N_200,In_2333,In_1190);
or U201 (N_201,In_1627,In_60);
or U202 (N_202,In_615,In_1753);
and U203 (N_203,In_788,In_1898);
nand U204 (N_204,In_1964,In_1892);
nand U205 (N_205,In_310,In_218);
nor U206 (N_206,In_871,In_325);
or U207 (N_207,In_832,In_75);
and U208 (N_208,In_1032,In_1287);
and U209 (N_209,In_2435,In_1198);
and U210 (N_210,In_2343,In_2185);
nor U211 (N_211,In_460,In_1304);
nor U212 (N_212,In_9,In_931);
or U213 (N_213,In_56,In_2285);
xnor U214 (N_214,In_1775,In_914);
or U215 (N_215,In_1819,In_1254);
nand U216 (N_216,In_2299,In_2142);
nand U217 (N_217,In_478,In_1844);
nand U218 (N_218,In_482,In_2448);
and U219 (N_219,In_1112,In_762);
xor U220 (N_220,In_1156,In_394);
nand U221 (N_221,In_744,In_1590);
and U222 (N_222,In_379,In_1825);
nor U223 (N_223,In_2061,In_929);
nor U224 (N_224,In_1828,In_1305);
or U225 (N_225,In_1691,In_2186);
nor U226 (N_226,In_1140,In_747);
xnor U227 (N_227,In_893,In_2481);
xor U228 (N_228,In_462,In_865);
and U229 (N_229,In_1746,In_1109);
nand U230 (N_230,In_322,In_182);
and U231 (N_231,In_475,In_70);
xor U232 (N_232,In_1235,In_105);
or U233 (N_233,In_1130,In_1435);
xnor U234 (N_234,In_1537,In_2480);
xnor U235 (N_235,In_204,In_2164);
or U236 (N_236,In_1649,In_2495);
xor U237 (N_237,In_2284,In_1168);
and U238 (N_238,In_1402,In_1488);
xnor U239 (N_239,In_1793,In_545);
and U240 (N_240,In_2406,In_1384);
nor U241 (N_241,In_2411,In_2228);
nand U242 (N_242,In_1573,In_2357);
and U243 (N_243,In_1761,In_508);
nor U244 (N_244,In_2311,In_2439);
xor U245 (N_245,In_619,In_1383);
nand U246 (N_246,In_2237,In_2359);
nand U247 (N_247,In_1072,In_1701);
and U248 (N_248,In_1239,In_1357);
nor U249 (N_249,In_1707,In_50);
nand U250 (N_250,In_2253,In_1652);
nor U251 (N_251,In_2047,In_1766);
or U252 (N_252,In_2430,In_1835);
xor U253 (N_253,In_1657,In_491);
nor U254 (N_254,In_2322,In_523);
or U255 (N_255,In_1577,In_894);
nor U256 (N_256,In_1090,In_916);
xnor U257 (N_257,In_263,In_1191);
nor U258 (N_258,In_956,In_1313);
or U259 (N_259,In_503,In_1559);
nor U260 (N_260,In_101,In_1181);
or U261 (N_261,In_1823,In_1928);
and U262 (N_262,In_1265,In_1475);
nor U263 (N_263,In_1042,In_889);
nor U264 (N_264,In_2374,In_2298);
nand U265 (N_265,In_1677,In_638);
nand U266 (N_266,In_367,In_2425);
nor U267 (N_267,In_2498,In_2064);
xnor U268 (N_268,In_2103,In_1926);
or U269 (N_269,In_695,In_2035);
or U270 (N_270,In_2358,In_726);
nand U271 (N_271,In_2006,In_1161);
nand U272 (N_272,In_464,In_1564);
nor U273 (N_273,In_2486,In_2012);
xnor U274 (N_274,In_376,In_2045);
nor U275 (N_275,In_868,In_2031);
or U276 (N_276,In_1864,In_1875);
nor U277 (N_277,In_1596,In_710);
nand U278 (N_278,In_696,In_1840);
or U279 (N_279,In_1080,In_1711);
and U280 (N_280,In_1476,In_1718);
nand U281 (N_281,In_1236,In_2130);
nand U282 (N_282,In_131,In_453);
and U283 (N_283,In_1800,In_2438);
and U284 (N_284,In_1920,In_813);
xor U285 (N_285,In_1754,In_1619);
and U286 (N_286,In_866,In_972);
xnor U287 (N_287,In_702,In_1744);
and U288 (N_288,In_1725,In_243);
xnor U289 (N_289,In_34,In_1356);
or U290 (N_290,In_2028,In_1049);
xor U291 (N_291,In_186,In_260);
and U292 (N_292,In_469,In_1889);
and U293 (N_293,In_252,In_890);
and U294 (N_294,In_153,In_1310);
xor U295 (N_295,In_2274,In_501);
or U296 (N_296,In_668,In_358);
or U297 (N_297,In_770,In_157);
xor U298 (N_298,In_1546,In_166);
and U299 (N_299,In_2420,In_585);
and U300 (N_300,In_1092,In_1443);
and U301 (N_301,In_454,In_551);
nor U302 (N_302,In_1373,In_978);
xor U303 (N_303,In_876,In_2323);
and U304 (N_304,In_1558,In_90);
nand U305 (N_305,In_2055,In_1811);
or U306 (N_306,In_299,In_1147);
xnor U307 (N_307,In_1240,In_2467);
nand U308 (N_308,In_2361,In_1803);
nor U309 (N_309,In_1084,In_2089);
xor U310 (N_310,In_1862,In_1382);
nor U311 (N_311,In_2458,In_215);
and U312 (N_312,In_1261,In_1556);
nand U313 (N_313,In_540,In_2083);
or U314 (N_314,In_1271,In_159);
and U315 (N_315,In_1269,In_116);
and U316 (N_316,In_936,In_2346);
nor U317 (N_317,In_1237,In_1719);
xnor U318 (N_318,In_1077,In_233);
nor U319 (N_319,In_212,In_1244);
or U320 (N_320,In_1780,In_84);
nand U321 (N_321,In_390,In_1116);
nor U322 (N_322,In_2450,In_1388);
xor U323 (N_323,In_386,In_730);
and U324 (N_324,In_941,In_856);
nand U325 (N_325,In_1541,In_944);
nand U326 (N_326,In_672,In_1592);
xnor U327 (N_327,In_1715,In_1782);
nand U328 (N_328,In_836,In_1315);
nor U329 (N_329,In_202,In_1250);
xor U330 (N_330,In_690,In_1943);
nand U331 (N_331,In_2229,In_354);
or U332 (N_332,In_2234,In_360);
and U333 (N_333,In_1428,In_784);
nor U334 (N_334,In_907,In_405);
xnor U335 (N_335,In_189,In_2194);
or U336 (N_336,In_1972,In_1005);
nand U337 (N_337,In_449,In_2119);
nor U338 (N_338,In_600,In_1783);
xnor U339 (N_339,In_899,In_2489);
nand U340 (N_340,In_807,In_1115);
or U341 (N_341,In_1751,In_999);
nand U342 (N_342,In_1931,In_1457);
nand U343 (N_343,In_2231,In_241);
or U344 (N_344,In_283,In_1111);
nor U345 (N_345,In_2307,In_1063);
or U346 (N_346,In_1387,In_1377);
xor U347 (N_347,In_909,In_732);
xor U348 (N_348,In_1769,In_1372);
or U349 (N_349,In_351,In_797);
nor U350 (N_350,In_2218,In_42);
nor U351 (N_351,In_984,In_1158);
or U352 (N_352,In_1125,In_2449);
nand U353 (N_353,In_1358,In_439);
nor U354 (N_354,In_95,In_757);
or U355 (N_355,In_1159,In_1616);
and U356 (N_356,In_1747,In_2204);
nand U357 (N_357,In_673,In_1913);
nand U358 (N_358,In_1188,In_2197);
and U359 (N_359,In_2026,In_538);
nor U360 (N_360,In_1132,In_607);
and U361 (N_361,In_1626,In_1709);
xnor U362 (N_362,In_81,In_318);
nand U363 (N_363,In_679,In_514);
nand U364 (N_364,In_524,In_417);
nand U365 (N_365,In_2004,In_2499);
and U366 (N_366,In_103,In_369);
nand U367 (N_367,In_1535,In_703);
nor U368 (N_368,In_1628,In_1955);
nor U369 (N_369,In_1604,In_1906);
nor U370 (N_370,In_1521,In_1771);
nor U371 (N_371,In_1038,In_1824);
xnor U372 (N_372,In_2109,In_300);
and U373 (N_373,In_1665,In_2426);
or U374 (N_374,In_1676,In_445);
and U375 (N_375,In_2399,In_2114);
xnor U376 (N_376,In_339,In_1389);
or U377 (N_377,In_1451,In_754);
xor U378 (N_378,In_122,In_219);
nor U379 (N_379,In_2474,In_2215);
xor U380 (N_380,In_1268,In_796);
nor U381 (N_381,In_1989,In_2351);
xnor U382 (N_382,In_112,In_1583);
xnor U383 (N_383,In_316,In_1799);
and U384 (N_384,In_2000,In_2071);
nor U385 (N_385,In_2201,In_1106);
xnor U386 (N_386,In_532,In_392);
nand U387 (N_387,In_1722,In_812);
nor U388 (N_388,In_399,In_352);
nand U389 (N_389,In_620,In_185);
and U390 (N_390,In_1774,In_1421);
nand U391 (N_391,In_330,In_2096);
nor U392 (N_392,In_2034,In_1636);
nor U393 (N_393,In_1914,In_1020);
and U394 (N_394,In_293,In_2144);
nor U395 (N_395,In_2111,In_1578);
xnor U396 (N_396,In_874,In_712);
xor U397 (N_397,In_142,In_922);
xnor U398 (N_398,In_194,In_2331);
nor U399 (N_399,In_1951,In_1485);
nand U400 (N_400,In_1735,In_2256);
and U401 (N_401,In_1638,In_2292);
nor U402 (N_402,In_748,In_1243);
nand U403 (N_403,In_1338,In_843);
nor U404 (N_404,In_1489,In_1888);
or U405 (N_405,In_2060,In_1678);
xor U406 (N_406,In_456,In_1266);
nor U407 (N_407,In_986,In_12);
and U408 (N_408,In_2052,In_1061);
nand U409 (N_409,In_311,In_1834);
nor U410 (N_410,In_1870,In_1000);
xor U411 (N_411,In_1566,In_1688);
xor U412 (N_412,In_845,In_1264);
xor U413 (N_413,In_2443,In_1973);
or U414 (N_414,In_1410,In_2009);
xnor U415 (N_415,In_1334,In_1798);
nor U416 (N_416,In_1520,In_605);
and U417 (N_417,In_237,In_1532);
or U418 (N_418,In_1481,In_1571);
xnor U419 (N_419,In_2330,In_735);
nor U420 (N_420,In_2038,In_2094);
and U421 (N_421,In_430,In_1880);
nand U422 (N_422,In_1364,In_2036);
and U423 (N_423,In_179,In_2222);
or U424 (N_424,In_477,In_217);
nand U425 (N_425,In_1136,In_1374);
nand U426 (N_426,In_362,In_1765);
or U427 (N_427,In_2095,In_1189);
nor U428 (N_428,In_173,In_226);
nand U429 (N_429,In_1703,In_952);
or U430 (N_430,In_2167,In_1855);
and U431 (N_431,In_435,In_1789);
xor U432 (N_432,In_1856,In_230);
nor U433 (N_433,In_1550,In_169);
xnor U434 (N_434,In_731,In_823);
xnor U435 (N_435,In_2492,In_2370);
or U436 (N_436,In_549,In_1668);
or U437 (N_437,In_1153,In_1595);
xnor U438 (N_438,In_895,In_1450);
or U439 (N_439,In_2457,In_323);
xnor U440 (N_440,In_2200,In_1796);
nor U441 (N_441,In_758,In_324);
xor U442 (N_442,In_443,In_1220);
nand U443 (N_443,In_2053,In_2352);
or U444 (N_444,In_1085,In_1991);
xnor U445 (N_445,In_1438,In_473);
xnor U446 (N_446,In_1110,In_2497);
nand U447 (N_447,In_1818,In_1529);
xnor U448 (N_448,In_455,In_2127);
and U449 (N_449,In_85,In_1105);
or U450 (N_450,In_378,In_2336);
nor U451 (N_451,In_1967,In_1954);
and U452 (N_452,In_1355,In_1200);
nand U453 (N_453,In_1759,In_776);
and U454 (N_454,In_2441,In_2240);
nor U455 (N_455,In_1023,In_1231);
or U456 (N_456,In_906,In_1225);
or U457 (N_457,In_338,In_2452);
nand U458 (N_458,In_657,In_2062);
xnor U459 (N_459,In_1867,In_517);
nor U460 (N_460,In_1427,In_2195);
nand U461 (N_461,In_1869,In_337);
xnor U462 (N_462,In_1143,In_1022);
or U463 (N_463,In_2199,In_782);
nor U464 (N_464,In_2072,In_347);
or U465 (N_465,In_1054,In_1371);
or U466 (N_466,In_340,In_709);
xor U467 (N_467,In_858,In_728);
xnor U468 (N_468,In_1790,In_2396);
nor U469 (N_469,In_1412,In_1838);
and U470 (N_470,In_1947,In_905);
nor U471 (N_471,In_1403,In_11);
xnor U472 (N_472,In_38,In_2168);
nand U473 (N_473,In_2417,In_1536);
xor U474 (N_474,In_581,In_2220);
nand U475 (N_475,In_250,In_586);
and U476 (N_476,In_2161,In_428);
and U477 (N_477,In_2020,In_2073);
and U478 (N_478,In_1210,In_389);
nor U479 (N_479,In_1924,In_319);
xor U480 (N_480,In_1922,In_564);
and U481 (N_481,In_1560,In_1363);
nand U482 (N_482,In_578,In_1202);
nand U483 (N_483,In_479,In_1601);
xnor U484 (N_484,In_1776,In_2015);
nor U485 (N_485,In_1728,In_493);
or U486 (N_486,In_1393,In_1272);
xor U487 (N_487,In_2451,In_214);
or U488 (N_488,In_2165,In_953);
nand U489 (N_489,In_958,In_32);
nor U490 (N_490,In_2157,In_719);
xor U491 (N_491,In_2163,In_1505);
or U492 (N_492,In_403,In_1609);
xnor U493 (N_493,In_1666,In_2041);
and U494 (N_494,In_1804,In_150);
nand U495 (N_495,In_2156,In_1826);
nor U496 (N_496,In_1993,In_74);
or U497 (N_497,In_402,In_2067);
nand U498 (N_498,In_1600,In_1515);
xor U499 (N_499,In_2140,In_1726);
nor U500 (N_500,In_1083,In_2381);
nand U501 (N_501,In_1217,In_2084);
or U502 (N_502,In_1945,In_1484);
nor U503 (N_503,In_921,In_763);
xnor U504 (N_504,In_1326,In_128);
and U505 (N_505,In_1321,In_82);
xnor U506 (N_506,In_1995,In_2356);
nor U507 (N_507,In_675,In_504);
and U508 (N_508,In_2246,In_1637);
and U509 (N_509,In_1490,In_1342);
nand U510 (N_510,In_651,In_1053);
nand U511 (N_511,In_888,In_499);
nand U512 (N_512,In_740,In_216);
nor U513 (N_513,In_655,In_974);
or U514 (N_514,In_1976,In_513);
and U515 (N_515,In_913,In_2102);
and U516 (N_516,In_2141,In_834);
xor U517 (N_517,In_2074,In_1695);
xor U518 (N_518,In_2049,In_1144);
nor U519 (N_519,In_2171,In_1399);
and U520 (N_520,In_1420,In_554);
xnor U521 (N_521,In_320,In_1608);
nor U522 (N_522,In_795,In_467);
xor U523 (N_523,In_370,In_298);
or U524 (N_524,In_2490,In_940);
or U525 (N_525,In_446,In_595);
nor U526 (N_526,In_44,In_1896);
or U527 (N_527,In_1858,In_425);
or U528 (N_528,In_1755,In_1460);
or U529 (N_529,In_1648,In_612);
xnor U530 (N_530,In_1308,In_154);
nand U531 (N_531,In_2445,In_1758);
nor U532 (N_532,In_512,In_2463);
xor U533 (N_533,In_2148,In_1850);
nand U534 (N_534,In_224,In_771);
and U535 (N_535,In_816,In_1417);
and U536 (N_536,In_33,In_1621);
or U537 (N_537,In_1713,In_1622);
and U538 (N_538,In_2134,In_745);
nor U539 (N_539,In_242,In_700);
nand U540 (N_540,In_132,In_515);
and U541 (N_541,In_1639,In_1857);
nor U542 (N_542,In_344,In_387);
xnor U543 (N_543,In_951,In_674);
nor U544 (N_544,In_2327,In_1884);
and U545 (N_545,In_1050,In_648);
xor U546 (N_546,In_2391,In_1743);
xnor U547 (N_547,In_2410,In_39);
or U548 (N_548,In_1814,In_1708);
or U549 (N_549,In_2176,In_808);
and U550 (N_550,In_2301,In_2118);
nand U551 (N_551,In_1679,In_1543);
or U552 (N_552,In_759,In_258);
or U553 (N_553,In_2278,In_1102);
nand U554 (N_554,In_1584,In_661);
or U555 (N_555,In_1224,In_1589);
nand U556 (N_556,In_2390,In_437);
xor U557 (N_557,In_1155,In_30);
xnor U558 (N_558,In_382,In_727);
xnor U559 (N_559,In_993,In_2302);
nand U560 (N_560,In_393,In_1444);
or U561 (N_561,In_76,In_518);
and U562 (N_562,In_1164,In_2408);
or U563 (N_563,In_329,In_36);
or U564 (N_564,In_2003,In_1684);
and U565 (N_565,In_1737,In_1432);
nor U566 (N_566,In_86,In_977);
nand U567 (N_567,In_1107,In_2360);
and U568 (N_568,In_487,In_1610);
nor U569 (N_569,In_2125,In_1282);
nand U570 (N_570,In_1229,In_848);
nor U571 (N_571,In_1230,In_1710);
xor U572 (N_572,In_1152,In_2279);
and U573 (N_573,In_1316,In_1859);
and U574 (N_574,In_1516,In_2428);
xnor U575 (N_575,In_1929,In_1545);
nor U576 (N_576,In_934,In_366);
or U577 (N_577,In_492,In_207);
nor U578 (N_578,In_1067,In_1199);
nor U579 (N_579,In_1470,In_2132);
xor U580 (N_580,In_1154,In_2209);
and U581 (N_581,In_765,In_1846);
nor U582 (N_582,In_2155,In_25);
and U583 (N_583,In_1285,In_303);
or U584 (N_584,In_544,In_1197);
xor U585 (N_585,In_629,In_1296);
and U586 (N_586,In_1522,In_1352);
xor U587 (N_587,In_1325,In_552);
and U588 (N_588,In_2479,In_134);
nor U589 (N_589,In_14,In_46);
xnor U590 (N_590,In_609,In_1643);
nand U591 (N_591,In_2092,In_1058);
or U592 (N_592,In_2233,In_1841);
nor U593 (N_593,In_457,In_463);
nor U594 (N_594,In_767,In_904);
or U595 (N_595,In_777,In_2376);
or U596 (N_596,In_383,In_1815);
and U597 (N_597,In_2151,In_1772);
and U598 (N_598,In_307,In_2377);
nor U599 (N_599,In_558,In_1930);
nor U600 (N_600,In_490,In_1670);
nand U601 (N_601,In_2080,In_1211);
nand U602 (N_602,In_1024,In_253);
nand U603 (N_603,In_1971,In_643);
xnor U604 (N_604,In_1398,In_1233);
or U605 (N_605,In_1007,In_898);
or U606 (N_606,In_1620,In_2100);
xor U607 (N_607,In_256,In_1501);
nor U608 (N_608,In_1816,In_659);
nand U609 (N_609,In_1887,In_541);
or U610 (N_610,In_1303,In_2238);
nor U611 (N_611,In_1478,In_1647);
or U612 (N_612,In_1319,In_1635);
nor U613 (N_613,In_1252,In_1606);
nor U614 (N_614,In_2315,In_149);
and U615 (N_615,In_1259,In_1041);
nand U616 (N_616,In_1445,In_297);
nor U617 (N_617,In_996,In_1661);
or U618 (N_618,In_1851,In_2310);
or U619 (N_619,In_1949,In_55);
xor U620 (N_620,In_1286,In_423);
and U621 (N_621,In_114,In_1277);
xnor U622 (N_622,In_275,In_384);
nor U623 (N_623,In_1406,In_2069);
or U624 (N_624,In_2289,In_1312);
nand U625 (N_625,In_535,In_1361);
or U626 (N_626,In_928,In_680);
or U627 (N_627,In_1987,In_1812);
or U628 (N_628,In_886,In_1340);
nor U629 (N_629,In_915,In_1201);
nand U630 (N_630,In_2473,In_630);
nand U631 (N_631,In_2388,In_175);
or U632 (N_632,In_1923,In_1035);
nor U633 (N_633,In_433,In_1221);
nor U634 (N_634,In_1045,In_1288);
xnor U635 (N_635,In_2251,In_1002);
and U636 (N_636,In_1863,In_2418);
nor U637 (N_637,In_421,In_1510);
nor U638 (N_638,In_1070,In_312);
and U639 (N_639,In_244,In_766);
nor U640 (N_640,In_125,In_1554);
and U641 (N_641,In_1205,In_669);
or U642 (N_642,In_1832,In_1509);
nor U643 (N_643,In_522,In_429);
and U644 (N_644,In_1974,In_192);
nor U645 (N_645,In_663,In_1390);
xor U646 (N_646,In_1784,In_2249);
nand U647 (N_647,In_1942,In_1873);
nor U648 (N_648,In_1263,In_2010);
xnor U649 (N_649,In_1299,In_1868);
xor U650 (N_650,In_1692,In_2271);
nand U651 (N_651,In_1184,In_183);
xnor U652 (N_652,In_1101,In_2470);
xnor U653 (N_653,In_1057,In_686);
xnor U654 (N_654,In_2395,In_264);
nand U655 (N_655,In_1436,In_1021);
and U656 (N_656,In_1741,In_530);
and U657 (N_657,In_171,In_24);
xor U658 (N_658,In_1997,In_2368);
or U659 (N_659,In_1448,In_1694);
xnor U660 (N_660,In_1587,In_1344);
nor U661 (N_661,In_923,In_332);
xor U662 (N_662,In_1646,In_1267);
or U663 (N_663,In_334,In_480);
nand U664 (N_664,In_2309,In_138);
and U665 (N_665,In_225,In_587);
xnor U666 (N_666,In_1588,In_1454);
or U667 (N_667,In_1433,In_760);
nor U668 (N_668,In_1311,In_333);
and U669 (N_669,In_1099,In_1905);
and U670 (N_670,In_1486,In_752);
or U671 (N_671,In_2099,In_1479);
xor U672 (N_672,In_2477,In_678);
nand U673 (N_673,In_2436,In_1497);
nor U674 (N_674,In_2264,In_1318);
nor U675 (N_675,In_660,In_1492);
or U676 (N_676,In_2366,In_2087);
nor U677 (N_677,In_1134,In_1214);
and U678 (N_678,In_1962,In_1336);
or U679 (N_679,In_963,In_779);
or U680 (N_680,In_1353,In_1001);
or U681 (N_681,In_883,In_1149);
and U682 (N_682,In_2355,In_1852);
nand U683 (N_683,In_1418,In_1513);
and U684 (N_684,In_1698,In_2421);
or U685 (N_685,In_287,In_100);
and U686 (N_686,In_281,In_2281);
nor U687 (N_687,In_2192,In_1585);
and U688 (N_688,In_1322,In_717);
nand U689 (N_689,In_184,In_826);
nand U690 (N_690,In_716,In_1208);
nor U691 (N_691,In_222,In_2243);
nand U692 (N_692,In_2014,In_2019);
nor U693 (N_693,In_1723,In_1104);
and U694 (N_694,In_451,In_1839);
or U695 (N_695,In_1031,In_1910);
and U696 (N_696,In_1345,In_2364);
nor U697 (N_697,In_2332,In_1011);
nor U698 (N_698,In_432,In_1094);
nor U699 (N_699,In_720,In_2483);
nor U700 (N_700,In_579,In_188);
nand U701 (N_701,In_601,In_13);
nor U702 (N_702,In_616,In_1017);
or U703 (N_703,In_1395,In_1999);
or U704 (N_704,In_2023,In_683);
nor U705 (N_705,In_1524,In_292);
or U706 (N_706,In_231,In_2097);
xor U707 (N_707,In_412,In_1682);
xor U708 (N_708,In_569,In_1491);
or U709 (N_709,In_444,In_635);
or U710 (N_710,In_1434,In_844);
xnor U711 (N_711,In_536,In_2063);
and U712 (N_712,In_1900,In_2022);
or U713 (N_713,In_1347,In_2236);
or U714 (N_714,In_1580,In_864);
nor U715 (N_715,In_2137,In_1483);
nor U716 (N_716,In_365,In_725);
nand U717 (N_717,In_2065,In_1717);
and U718 (N_718,In_1128,In_1385);
or U719 (N_719,In_1773,In_2033);
xnor U720 (N_720,In_1242,In_1300);
and U721 (N_721,In_2482,In_1258);
or U722 (N_722,In_21,In_1337);
xnor U723 (N_723,In_2224,In_556);
nand U724 (N_724,In_1466,In_500);
xor U725 (N_725,In_2037,In_1234);
and U726 (N_726,In_1854,In_917);
nand U727 (N_727,In_1948,In_2121);
nor U728 (N_728,In_1370,In_1934);
and U729 (N_729,In_1827,In_1256);
nand U730 (N_730,In_2227,In_1290);
and U731 (N_731,In_2042,In_1215);
or U732 (N_732,In_156,In_191);
and U733 (N_733,In_2329,In_2007);
xnor U734 (N_734,In_1990,In_567);
or U735 (N_735,In_1380,In_1633);
and U736 (N_736,In_2175,In_1291);
nand U737 (N_737,In_88,In_2393);
nand U738 (N_738,In_280,In_381);
or U739 (N_739,In_1602,In_468);
and U740 (N_740,In_1273,In_2335);
xnor U741 (N_741,In_634,In_1047);
or U742 (N_742,In_2082,In_7);
xor U743 (N_743,In_2440,In_1465);
xnor U744 (N_744,In_1551,In_261);
or U745 (N_745,In_1043,In_180);
and U746 (N_746,In_1821,In_2232);
xnor U747 (N_747,In_1354,In_1712);
nor U748 (N_748,In_355,In_793);
nor U749 (N_749,In_2265,In_1367);
xor U750 (N_750,In_436,In_2056);
or U751 (N_751,In_681,In_1686);
xnor U752 (N_752,In_519,In_1770);
or U753 (N_753,In_1969,In_2385);
and U754 (N_754,In_418,In_1103);
and U755 (N_755,In_1139,In_1219);
nand U756 (N_756,In_67,In_2431);
xor U757 (N_757,In_1607,In_165);
nor U758 (N_758,In_1368,In_2442);
nor U759 (N_759,In_64,In_1740);
or U760 (N_760,In_878,In_1343);
and U761 (N_761,In_819,In_1757);
nor U762 (N_762,In_2128,In_1179);
nand U763 (N_763,In_279,In_772);
or U764 (N_764,In_1196,In_2212);
xor U765 (N_765,In_2086,In_566);
and U766 (N_766,In_466,In_1391);
xnor U767 (N_767,In_2384,In_120);
or U768 (N_768,In_1320,In_2453);
and U769 (N_769,In_1659,In_1378);
and U770 (N_770,In_1980,In_1655);
or U771 (N_771,In_764,In_1807);
nand U772 (N_772,In_665,In_927);
or U773 (N_773,In_2485,In_1938);
and U774 (N_774,In_368,In_1611);
nor U775 (N_775,In_111,In_1597);
xor U776 (N_776,In_2098,In_521);
and U777 (N_777,In_516,In_1822);
or U778 (N_778,In_1040,In_2306);
nor U779 (N_779,In_2287,In_2290);
or U780 (N_780,In_1227,In_288);
nor U781 (N_781,In_1145,In_1939);
or U782 (N_782,In_2313,In_1386);
nand U783 (N_783,In_2314,In_37);
or U784 (N_784,In_1089,In_966);
nand U785 (N_785,In_1853,In_1182);
nor U786 (N_786,In_633,In_1014);
nor U787 (N_787,In_2454,In_525);
or U788 (N_788,In_1212,In_891);
nor U789 (N_789,In_108,In_1625);
or U790 (N_790,In_255,In_739);
and U791 (N_791,In_2210,In_1082);
or U792 (N_792,In_2402,In_141);
nor U793 (N_793,In_846,In_821);
and U794 (N_794,In_1632,In_1157);
nand U795 (N_795,In_2280,In_571);
or U796 (N_796,In_613,In_1642);
or U797 (N_797,In_593,In_452);
nor U798 (N_798,In_1472,In_1396);
nor U799 (N_799,In_127,In_604);
nor U800 (N_800,In_957,In_2382);
nand U801 (N_801,In_31,In_1120);
nor U802 (N_802,In_1916,In_2214);
and U803 (N_803,In_1463,In_1534);
nand U804 (N_804,In_542,In_1405);
or U805 (N_805,In_1565,In_484);
and U806 (N_806,In_1133,In_1193);
and U807 (N_807,In_1376,In_1160);
and U808 (N_808,In_2138,In_1705);
nand U809 (N_809,In_632,In_860);
nand U810 (N_810,In_597,In_869);
nor U811 (N_811,In_851,In_1685);
nor U812 (N_812,In_8,In_964);
nand U813 (N_813,In_1010,In_1866);
xnor U814 (N_814,In_818,In_1055);
and U815 (N_815,In_1151,In_1919);
and U816 (N_816,In_170,In_1294);
or U817 (N_817,In_1178,In_1302);
or U818 (N_818,In_792,In_136);
or U819 (N_819,In_1683,In_2085);
and U820 (N_820,In_472,In_2048);
nor U821 (N_821,In_975,In_1019);
nand U822 (N_822,In_248,In_251);
xor U823 (N_823,In_965,In_505);
nor U824 (N_824,In_266,In_2070);
or U825 (N_825,In_1618,In_2447);
nor U826 (N_826,In_2259,In_77);
or U827 (N_827,In_1561,In_133);
nand U828 (N_828,In_1833,In_863);
or U829 (N_829,In_1836,In_809);
xnor U830 (N_830,In_998,In_1333);
nand U831 (N_831,In_824,In_1039);
and U832 (N_832,In_980,In_2300);
or U833 (N_833,In_1605,In_221);
and U834 (N_834,In_1702,In_1806);
nor U835 (N_835,In_353,In_1902);
or U836 (N_836,In_229,In_2250);
nand U837 (N_837,In_2416,In_2252);
nand U838 (N_838,In_278,In_738);
and U839 (N_839,In_249,In_1582);
xnor U840 (N_840,In_2051,In_1401);
nor U841 (N_841,In_450,In_1480);
or U842 (N_842,In_1975,In_1046);
or U843 (N_843,In_1553,In_1570);
and U844 (N_844,In_1379,In_1690);
nand U845 (N_845,In_983,In_227);
and U846 (N_846,In_1956,In_948);
xor U847 (N_847,In_18,In_1764);
or U848 (N_848,In_1574,In_658);
nand U849 (N_849,In_2208,In_903);
or U850 (N_850,In_926,In_2276);
nor U851 (N_851,In_1687,In_2409);
xnor U852 (N_852,In_938,In_1502);
and U853 (N_853,In_290,In_502);
nand U854 (N_854,In_831,In_1495);
xnor U855 (N_855,In_377,In_1226);
xor U856 (N_856,In_1289,In_470);
nand U857 (N_857,In_271,In_1426);
or U858 (N_858,In_494,In_1952);
and U859 (N_859,In_2179,In_689);
nand U860 (N_860,In_1329,In_2437);
or U861 (N_861,In_59,In_692);
or U862 (N_862,In_1339,In_2296);
nor U863 (N_863,In_1207,In_427);
xor U864 (N_864,In_1194,In_733);
nand U865 (N_865,In_265,In_79);
nor U866 (N_866,In_2182,In_195);
or U867 (N_867,In_839,In_1893);
nand U868 (N_868,In_718,In_1915);
and U869 (N_869,In_327,In_572);
xnor U870 (N_870,In_220,In_239);
nor U871 (N_871,In_687,In_1081);
or U872 (N_872,In_1431,In_398);
nor U873 (N_873,In_2181,In_2225);
xnor U874 (N_874,In_1629,In_507);
nand U875 (N_875,In_161,In_822);
and U876 (N_876,In_19,In_2216);
xor U877 (N_877,In_1795,In_1148);
nor U878 (N_878,In_781,In_1381);
xnor U879 (N_879,In_442,In_2269);
xor U880 (N_880,In_2494,In_448);
nor U881 (N_881,In_1170,In_276);
nand U882 (N_882,In_1175,In_1843);
xor U883 (N_883,In_756,In_1714);
or U884 (N_884,In_2378,In_510);
nand U885 (N_885,In_2491,In_560);
or U886 (N_886,In_1631,In_441);
nor U887 (N_887,In_794,In_1729);
nor U888 (N_888,In_1349,In_2123);
nand U889 (N_889,In_2170,In_1247);
and U890 (N_890,In_1441,In_933);
nand U891 (N_891,In_2029,In_174);
nor U892 (N_892,In_647,In_1504);
and U893 (N_893,In_1903,In_2347);
nor U894 (N_894,In_746,In_842);
xnor U895 (N_895,In_2152,In_1786);
or U896 (N_896,In_1012,In_301);
nand U897 (N_897,In_1871,In_2115);
nor U898 (N_898,In_2184,In_1581);
and U899 (N_899,In_1051,In_424);
nand U900 (N_900,In_361,In_167);
and U901 (N_901,In_1172,In_1894);
nor U902 (N_902,In_1283,In_1118);
nand U903 (N_903,In_2305,In_1762);
xnor U904 (N_904,In_193,In_2211);
and U905 (N_905,In_671,In_1963);
nor U906 (N_906,In_96,In_854);
xor U907 (N_907,In_1552,In_69);
or U908 (N_908,In_2120,In_670);
or U909 (N_909,In_2219,In_1332);
or U910 (N_910,In_1531,In_1567);
and U911 (N_911,In_594,In_124);
xor U912 (N_912,In_1946,In_71);
and U913 (N_913,In_837,In_790);
and U914 (N_914,In_1959,In_1419);
nor U915 (N_915,In_734,In_92);
xnor U916 (N_916,In_359,In_1366);
xor U917 (N_917,In_447,In_1424);
nand U918 (N_918,In_583,In_1293);
nor U919 (N_919,In_1936,In_208);
and U920 (N_920,In_543,In_2424);
or U921 (N_921,In_401,In_1848);
nor U922 (N_922,In_1986,In_1872);
xor U923 (N_923,In_1309,In_486);
nor U924 (N_924,In_420,In_568);
and U925 (N_925,In_715,In_2);
nand U926 (N_926,In_1137,In_970);
or U927 (N_927,In_1468,In_1328);
xor U928 (N_928,In_1241,In_828);
or U929 (N_929,In_1526,In_465);
xor U930 (N_930,In_1059,In_414);
nand U931 (N_931,In_714,In_946);
nor U932 (N_932,In_1768,In_2362);
nor U933 (N_933,In_2001,In_306);
xnor U934 (N_934,In_1469,In_119);
or U935 (N_935,In_2013,In_611);
and U936 (N_936,In_1918,In_1674);
nor U937 (N_937,In_1881,In_1327);
nand U938 (N_938,In_2324,In_1439);
nand U939 (N_939,In_1062,In_991);
or U940 (N_940,In_553,In_644);
xnor U941 (N_941,In_45,In_2133);
or U942 (N_942,In_238,In_273);
nor U943 (N_943,In_22,In_698);
nand U944 (N_944,In_1362,In_1961);
and U945 (N_945,In_2398,In_1078);
nand U946 (N_946,In_2146,In_798);
nand U947 (N_947,In_422,In_1186);
and U948 (N_948,In_53,In_2093);
and U949 (N_949,In_63,In_1150);
nand U950 (N_950,In_855,In_2057);
or U951 (N_951,In_2091,In_1612);
nor U952 (N_952,In_815,In_2434);
nor U953 (N_953,In_1292,In_783);
and U954 (N_954,In_415,In_1279);
nand U955 (N_955,In_2239,In_110);
xor U956 (N_956,In_459,In_2016);
or U957 (N_957,In_691,In_531);
and U958 (N_958,In_2021,In_1452);
xor U959 (N_959,In_646,In_1792);
nand U960 (N_960,In_397,In_565);
and U961 (N_961,In_2011,In_1994);
and U962 (N_962,In_2317,In_840);
and U963 (N_963,In_1802,In_2328);
nand U964 (N_964,In_1788,In_814);
and U965 (N_965,In_925,In_641);
xor U966 (N_966,In_83,In_1228);
and U967 (N_967,In_395,In_335);
nor U968 (N_968,In_2478,In_546);
or U969 (N_969,In_363,In_3);
and U970 (N_970,In_526,In_631);
nand U971 (N_971,In_506,In_145);
nor U972 (N_972,In_190,In_1317);
nand U973 (N_973,In_1341,In_2493);
and U974 (N_974,In_1036,In_277);
xnor U975 (N_975,In_2188,In_48);
nand U976 (N_976,In_817,In_1968);
and U977 (N_977,In_342,In_1262);
nand U978 (N_978,In_2432,In_847);
xnor U979 (N_979,In_129,In_1528);
nor U980 (N_980,In_284,In_458);
xor U981 (N_981,In_1346,In_1568);
or U982 (N_982,In_806,In_489);
nor U983 (N_983,In_1696,In_1801);
or U984 (N_984,In_400,In_1506);
nor U985 (N_985,In_1278,In_1895);
nand U986 (N_986,In_1127,In_1314);
and U987 (N_987,In_1369,In_1079);
xnor U988 (N_988,In_373,In_213);
and U989 (N_989,In_410,In_1238);
or U990 (N_990,In_721,In_1016);
nor U991 (N_991,In_326,In_2261);
nand U992 (N_992,In_1123,In_885);
and U993 (N_993,In_54,In_1280);
nand U994 (N_994,In_2122,In_1904);
nor U995 (N_995,In_407,In_1066);
and U996 (N_996,In_408,In_176);
or U997 (N_997,In_1114,In_73);
nand U998 (N_998,In_625,In_1324);
nor U999 (N_999,In_2135,In_68);
nor U1000 (N_1000,In_385,In_1519);
nor U1001 (N_1001,In_1917,In_935);
and U1002 (N_1002,In_2187,In_172);
or U1003 (N_1003,In_1213,In_164);
and U1004 (N_1004,In_1060,In_667);
nand U1005 (N_1005,In_1594,In_2295);
xor U1006 (N_1006,In_1407,In_550);
and U1007 (N_1007,In_1662,In_1656);
xor U1008 (N_1008,In_1044,In_1932);
nand U1009 (N_1009,In_291,In_2206);
and U1010 (N_1010,In_1025,In_1496);
or U1011 (N_1011,In_223,In_803);
nor U1012 (N_1012,In_2160,In_2320);
nor U1013 (N_1013,In_662,In_820);
nand U1014 (N_1014,In_2205,In_2283);
xor U1015 (N_1015,In_1514,In_2078);
nor U1016 (N_1016,In_2446,In_155);
nand U1017 (N_1017,In_1983,In_1908);
nand U1018 (N_1018,In_1940,In_954);
nor U1019 (N_1019,In_247,In_802);
nand U1020 (N_1020,In_2268,In_1660);
nor U1021 (N_1021,In_1876,In_413);
and U1022 (N_1022,In_773,In_1253);
xnor U1023 (N_1023,In_2046,In_932);
or U1024 (N_1024,In_345,In_158);
nand U1025 (N_1025,In_575,In_1658);
or U1026 (N_1026,In_749,In_1847);
nand U1027 (N_1027,In_1809,In_1400);
xnor U1028 (N_1028,In_168,In_2277);
and U1029 (N_1029,In_751,In_356);
and U1030 (N_1030,In_562,In_811);
or U1031 (N_1031,In_126,In_624);
nor U1032 (N_1032,In_1295,In_1615);
nand U1033 (N_1033,In_1669,In_139);
nand U1034 (N_1034,In_1028,In_210);
or U1035 (N_1035,In_985,In_676);
xor U1036 (N_1036,In_240,In_1572);
nand U1037 (N_1037,In_799,In_1455);
xor U1038 (N_1038,In_1810,In_143);
xor U1039 (N_1039,In_1979,In_1960);
or U1040 (N_1040,In_1180,In_497);
xor U1041 (N_1041,In_236,In_61);
nand U1042 (N_1042,In_873,In_988);
and U1043 (N_1043,In_203,In_1525);
xnor U1044 (N_1044,In_2414,In_537);
nor U1045 (N_1045,In_1738,In_557);
or U1046 (N_1046,In_2316,In_364);
or U1047 (N_1047,In_200,In_1246);
and U1048 (N_1048,In_1540,In_1721);
and U1049 (N_1049,In_774,In_2005);
nand U1050 (N_1050,In_1617,In_1899);
nand U1051 (N_1051,In_2244,In_1121);
nand U1052 (N_1052,In_2159,In_87);
and U1053 (N_1053,In_2338,In_272);
nand U1054 (N_1054,In_2002,In_2223);
xnor U1055 (N_1055,In_722,In_28);
xor U1056 (N_1056,In_786,In_1064);
and U1057 (N_1057,In_2191,In_947);
or U1058 (N_1058,In_599,In_1165);
and U1059 (N_1059,In_146,In_778);
xnor U1060 (N_1060,In_1569,In_755);
or U1061 (N_1061,In_1177,In_1667);
xor U1062 (N_1062,In_677,In_708);
xnor U1063 (N_1063,In_1634,In_2337);
nand U1064 (N_1064,In_2325,In_1323);
nand U1065 (N_1065,In_1845,In_1727);
or U1066 (N_1066,In_1350,In_2339);
nor U1067 (N_1067,In_315,In_419);
xnor U1068 (N_1068,In_2024,In_1614);
nor U1069 (N_1069,In_206,In_2076);
and U1070 (N_1070,In_2293,In_1517);
or U1071 (N_1071,In_509,In_1331);
xor U1072 (N_1072,In_1518,In_533);
nor U1073 (N_1073,In_2400,In_1831);
xor U1074 (N_1074,In_1675,In_1056);
or U1075 (N_1075,In_2050,In_1117);
nor U1076 (N_1076,In_849,In_1071);
or U1077 (N_1077,In_1013,In_1732);
xnor U1078 (N_1078,In_2116,In_1095);
or U1079 (N_1079,In_440,In_98);
and U1080 (N_1080,In_596,In_94);
nand U1081 (N_1081,In_2304,In_309);
and U1082 (N_1082,In_2018,In_2203);
and U1083 (N_1083,In_78,In_1650);
nand U1084 (N_1084,In_431,In_4);
xnor U1085 (N_1085,In_2248,In_1767);
or U1086 (N_1086,In_529,In_989);
and U1087 (N_1087,In_2282,In_1988);
nand U1088 (N_1088,In_602,In_488);
and U1089 (N_1089,In_645,In_850);
or U1090 (N_1090,In_62,In_1511);
nand U1091 (N_1091,In_52,In_1752);
or U1092 (N_1092,In_829,In_1464);
nor U1093 (N_1093,In_2030,In_896);
and U1094 (N_1094,In_1330,In_1992);
xnor U1095 (N_1095,In_2319,In_187);
nor U1096 (N_1096,In_246,In_1446);
nor U1097 (N_1097,In_995,In_80);
or U1098 (N_1098,In_969,In_2166);
xnor U1099 (N_1099,In_1599,In_1477);
xor U1100 (N_1100,In_1576,In_684);
nor U1101 (N_1101,In_705,In_1018);
or U1102 (N_1102,In_2059,In_2275);
or U1103 (N_1103,In_1958,In_1003);
or U1104 (N_1104,In_2129,In_1174);
and U1105 (N_1105,In_2254,In_2104);
or U1106 (N_1106,In_520,In_987);
or U1107 (N_1107,In_729,In_852);
nand U1108 (N_1108,In_137,In_682);
or U1109 (N_1109,In_17,In_471);
nor U1110 (N_1110,In_2371,In_1030);
and U1111 (N_1111,In_787,In_937);
and U1112 (N_1112,In_5,In_1255);
nand U1113 (N_1113,In_2354,In_346);
and U1114 (N_1114,In_930,In_1663);
nand U1115 (N_1115,In_1547,In_123);
nand U1116 (N_1116,In_1742,In_1232);
nand U1117 (N_1117,In_282,In_1409);
and U1118 (N_1118,In_753,In_742);
and U1119 (N_1119,In_1523,In_341);
nor U1120 (N_1120,In_971,In_1953);
nand U1121 (N_1121,In_1791,In_2373);
nor U1122 (N_1122,In_2136,In_1415);
or U1123 (N_1123,In_2202,In_2372);
nor U1124 (N_1124,In_1129,In_2113);
xnor U1125 (N_1125,In_1173,In_1539);
or U1126 (N_1126,In_1777,In_496);
nand U1127 (N_1127,In_1474,In_1849);
nand U1128 (N_1128,In_16,In_1538);
and U1129 (N_1129,In_1404,In_2487);
nor U1130 (N_1130,In_1886,In_1297);
nor U1131 (N_1131,In_286,In_2267);
nor U1132 (N_1132,In_2044,In_706);
nand U1133 (N_1133,In_1941,In_1471);
nand U1134 (N_1134,In_2260,In_1689);
or U1135 (N_1135,In_527,In_2456);
or U1136 (N_1136,In_372,In_942);
nand U1137 (N_1137,In_308,In_1204);
nor U1138 (N_1138,In_621,In_1430);
and U1139 (N_1139,In_1459,In_650);
or U1140 (N_1140,In_741,In_962);
nor U1141 (N_1141,In_27,In_313);
xor U1142 (N_1142,In_1276,In_328);
or U1143 (N_1143,In_791,In_2496);
nor U1144 (N_1144,In_1034,In_707);
or U1145 (N_1145,In_2126,In_2342);
xor U1146 (N_1146,In_1206,In_2353);
or U1147 (N_1147,In_391,In_737);
and U1148 (N_1148,In_0,In_1284);
nand U1149 (N_1149,In_911,In_411);
or U1150 (N_1150,In_2081,In_2471);
and U1151 (N_1151,In_2108,In_994);
and U1152 (N_1152,In_810,In_875);
xor U1153 (N_1153,In_1440,In_416);
or U1154 (N_1154,In_1874,In_2348);
nand U1155 (N_1155,In_511,In_2054);
nand U1156 (N_1156,In_1306,In_2272);
nand U1157 (N_1157,In_897,In_838);
and U1158 (N_1158,In_867,In_1307);
and U1159 (N_1159,In_1260,In_2266);
and U1160 (N_1160,In_1575,In_1223);
or U1161 (N_1161,In_1781,In_1146);
or U1162 (N_1162,In_636,In_591);
nand U1163 (N_1163,In_1671,In_197);
nor U1164 (N_1164,In_296,In_1950);
xor U1165 (N_1165,In_1456,In_555);
xor U1166 (N_1166,In_476,In_622);
xor U1167 (N_1167,In_584,In_610);
nand U1168 (N_1168,In_2344,In_1048);
or U1169 (N_1169,In_2150,In_257);
nand U1170 (N_1170,In_1985,In_1209);
nand U1171 (N_1171,In_106,In_2255);
and U1172 (N_1172,In_598,In_2173);
xnor U1173 (N_1173,In_57,In_841);
nor U1174 (N_1174,In_768,In_1124);
nor U1175 (N_1175,In_343,In_109);
nand U1176 (N_1176,In_2464,In_66);
nor U1177 (N_1177,In_900,In_294);
or U1178 (N_1178,In_1664,In_960);
or U1179 (N_1179,In_2090,In_198);
nor U1180 (N_1180,In_1837,In_2340);
or U1181 (N_1181,In_1487,In_1026);
or U1182 (N_1182,In_409,In_561);
and U1183 (N_1183,In_1613,In_1512);
xor U1184 (N_1184,In_804,In_1075);
xor U1185 (N_1185,In_780,In_2369);
or U1186 (N_1186,In_1586,In_912);
nor U1187 (N_1187,In_2242,In_304);
nor U1188 (N_1188,In_1562,In_1251);
nand U1189 (N_1189,In_434,In_2462);
nor U1190 (N_1190,In_1720,In_1359);
xor U1191 (N_1191,In_1073,In_1699);
and U1192 (N_1192,In_2334,In_2404);
nor U1193 (N_1193,In_872,In_2422);
and U1194 (N_1194,In_2468,In_99);
nor U1195 (N_1195,In_1640,In_1);
nand U1196 (N_1196,In_724,In_1335);
or U1197 (N_1197,In_801,In_1274);
nor U1198 (N_1198,In_1449,In_2043);
or U1199 (N_1199,In_269,In_115);
xor U1200 (N_1200,In_887,In_1027);
nor U1201 (N_1201,In_1982,In_1724);
and U1202 (N_1202,In_1169,In_1375);
or U1203 (N_1203,In_861,In_1029);
nor U1204 (N_1204,In_1088,In_1033);
or U1205 (N_1205,In_2415,In_58);
and U1206 (N_1206,In_1447,In_2077);
nand U1207 (N_1207,In_833,In_349);
xnor U1208 (N_1208,In_1733,In_1009);
xnor U1209 (N_1209,In_892,In_1096);
and U1210 (N_1210,In_1351,In_2312);
nor U1211 (N_1211,In_15,In_1397);
and U1212 (N_1212,In_2107,In_23);
nor U1213 (N_1213,In_1097,In_6);
nor U1214 (N_1214,In_380,In_2066);
nor U1215 (N_1215,In_2401,In_1623);
or U1216 (N_1216,In_199,In_1503);
nand U1217 (N_1217,In_652,In_1901);
or U1218 (N_1218,In_1065,In_2008);
nor U1219 (N_1219,In_151,In_1126);
nand U1220 (N_1220,In_723,In_163);
nor U1221 (N_1221,In_205,In_2392);
and U1222 (N_1222,In_1176,In_1119);
xor U1223 (N_1223,In_1882,In_2484);
nor U1224 (N_1224,In_1700,In_147);
and U1225 (N_1225,In_623,In_943);
and U1226 (N_1226,In_1998,In_800);
or U1227 (N_1227,In_1074,In_1493);
xnor U1228 (N_1228,In_1068,In_608);
nand U1229 (N_1229,In_1797,In_102);
nand U1230 (N_1230,In_2386,In_582);
and U1231 (N_1231,In_592,In_2433);
and U1232 (N_1232,In_49,In_357);
nor U1233 (N_1233,In_26,In_1817);
and U1234 (N_1234,In_160,In_1779);
xnor U1235 (N_1235,In_1195,In_2394);
xor U1236 (N_1236,In_2068,In_2221);
nand U1237 (N_1237,In_40,In_882);
and U1238 (N_1238,In_2039,In_2106);
nand U1239 (N_1239,In_2158,In_2412);
nand U1240 (N_1240,In_135,In_302);
nor U1241 (N_1241,In_699,In_485);
nand U1242 (N_1242,In_997,In_1163);
nand U1243 (N_1243,In_1098,In_1413);
or U1244 (N_1244,In_588,In_65);
or U1245 (N_1245,In_2145,In_426);
or U1246 (N_1246,In_1829,In_901);
nand U1247 (N_1247,In_1348,In_694);
and U1248 (N_1248,In_2455,In_590);
nand U1249 (N_1249,In_2241,In_1301);
nor U1250 (N_1250,In_2438,In_2003);
and U1251 (N_1251,In_948,In_1103);
and U1252 (N_1252,In_2137,In_1975);
and U1253 (N_1253,In_2475,In_23);
or U1254 (N_1254,In_902,In_1660);
nor U1255 (N_1255,In_2159,In_860);
or U1256 (N_1256,In_1092,In_1013);
xor U1257 (N_1257,In_1771,In_110);
nor U1258 (N_1258,In_1296,In_406);
and U1259 (N_1259,In_1170,In_710);
and U1260 (N_1260,In_2378,In_905);
or U1261 (N_1261,In_699,In_983);
nand U1262 (N_1262,In_2495,In_36);
nand U1263 (N_1263,In_776,In_1320);
xor U1264 (N_1264,In_41,In_1490);
or U1265 (N_1265,In_2002,In_783);
and U1266 (N_1266,In_1150,In_826);
and U1267 (N_1267,In_2381,In_880);
or U1268 (N_1268,In_2241,In_2135);
xor U1269 (N_1269,In_136,In_676);
or U1270 (N_1270,In_294,In_1616);
nand U1271 (N_1271,In_1417,In_400);
and U1272 (N_1272,In_15,In_32);
nor U1273 (N_1273,In_2124,In_1737);
and U1274 (N_1274,In_2390,In_931);
xnor U1275 (N_1275,In_821,In_695);
xnor U1276 (N_1276,In_645,In_1194);
and U1277 (N_1277,In_2472,In_58);
xor U1278 (N_1278,In_1356,In_2310);
nand U1279 (N_1279,In_2187,In_239);
and U1280 (N_1280,In_1655,In_7);
and U1281 (N_1281,In_1336,In_1313);
xnor U1282 (N_1282,In_2040,In_2130);
or U1283 (N_1283,In_1199,In_575);
or U1284 (N_1284,In_1068,In_1761);
nor U1285 (N_1285,In_1501,In_2405);
xnor U1286 (N_1286,In_2480,In_548);
and U1287 (N_1287,In_1490,In_2027);
and U1288 (N_1288,In_1209,In_2486);
or U1289 (N_1289,In_1197,In_566);
nand U1290 (N_1290,In_102,In_42);
xnor U1291 (N_1291,In_2387,In_805);
xnor U1292 (N_1292,In_1691,In_26);
xnor U1293 (N_1293,In_2106,In_1421);
nor U1294 (N_1294,In_1647,In_2128);
nand U1295 (N_1295,In_1304,In_1931);
or U1296 (N_1296,In_136,In_1275);
and U1297 (N_1297,In_1421,In_341);
xnor U1298 (N_1298,In_2068,In_458);
and U1299 (N_1299,In_145,In_2086);
and U1300 (N_1300,In_1250,In_1197);
nand U1301 (N_1301,In_2079,In_1323);
or U1302 (N_1302,In_1575,In_2174);
xor U1303 (N_1303,In_1368,In_2088);
xor U1304 (N_1304,In_2220,In_1210);
xnor U1305 (N_1305,In_2185,In_1726);
and U1306 (N_1306,In_2396,In_1859);
xnor U1307 (N_1307,In_1718,In_882);
xnor U1308 (N_1308,In_765,In_990);
nor U1309 (N_1309,In_1125,In_2126);
nor U1310 (N_1310,In_2187,In_1773);
or U1311 (N_1311,In_897,In_1088);
or U1312 (N_1312,In_802,In_698);
nand U1313 (N_1313,In_1966,In_210);
xnor U1314 (N_1314,In_2440,In_2338);
xor U1315 (N_1315,In_669,In_1506);
nand U1316 (N_1316,In_1543,In_2097);
nor U1317 (N_1317,In_1165,In_1080);
xnor U1318 (N_1318,In_115,In_918);
or U1319 (N_1319,In_2165,In_2493);
or U1320 (N_1320,In_1907,In_630);
nor U1321 (N_1321,In_124,In_1795);
and U1322 (N_1322,In_1954,In_2062);
xor U1323 (N_1323,In_808,In_1115);
or U1324 (N_1324,In_1160,In_2102);
nand U1325 (N_1325,In_1747,In_692);
or U1326 (N_1326,In_137,In_355);
and U1327 (N_1327,In_2334,In_1395);
and U1328 (N_1328,In_2295,In_975);
nor U1329 (N_1329,In_1692,In_2141);
and U1330 (N_1330,In_780,In_401);
xnor U1331 (N_1331,In_1934,In_1919);
nor U1332 (N_1332,In_119,In_1498);
xor U1333 (N_1333,In_1499,In_2208);
and U1334 (N_1334,In_285,In_2444);
and U1335 (N_1335,In_740,In_1994);
nand U1336 (N_1336,In_2409,In_447);
xnor U1337 (N_1337,In_240,In_1007);
nand U1338 (N_1338,In_2437,In_2283);
nand U1339 (N_1339,In_557,In_1317);
xnor U1340 (N_1340,In_1044,In_711);
nand U1341 (N_1341,In_649,In_870);
and U1342 (N_1342,In_723,In_885);
nand U1343 (N_1343,In_1235,In_1759);
or U1344 (N_1344,In_1120,In_2219);
and U1345 (N_1345,In_1907,In_272);
xnor U1346 (N_1346,In_837,In_955);
and U1347 (N_1347,In_994,In_897);
or U1348 (N_1348,In_2303,In_2437);
or U1349 (N_1349,In_561,In_1235);
nor U1350 (N_1350,In_1208,In_1962);
or U1351 (N_1351,In_1174,In_1667);
nor U1352 (N_1352,In_1,In_1719);
and U1353 (N_1353,In_314,In_858);
nor U1354 (N_1354,In_1668,In_1165);
nand U1355 (N_1355,In_1189,In_434);
nor U1356 (N_1356,In_408,In_2202);
xor U1357 (N_1357,In_1097,In_2258);
nand U1358 (N_1358,In_1254,In_1153);
nor U1359 (N_1359,In_251,In_5);
and U1360 (N_1360,In_1371,In_1963);
xor U1361 (N_1361,In_822,In_2244);
xor U1362 (N_1362,In_1631,In_2365);
nor U1363 (N_1363,In_1231,In_2109);
nor U1364 (N_1364,In_1460,In_1484);
xnor U1365 (N_1365,In_1979,In_59);
and U1366 (N_1366,In_376,In_1469);
xor U1367 (N_1367,In_3,In_1315);
and U1368 (N_1368,In_1367,In_829);
and U1369 (N_1369,In_1563,In_1549);
nor U1370 (N_1370,In_484,In_1885);
or U1371 (N_1371,In_850,In_1131);
nor U1372 (N_1372,In_2045,In_294);
nor U1373 (N_1373,In_1885,In_2469);
xnor U1374 (N_1374,In_520,In_500);
nand U1375 (N_1375,In_753,In_1309);
nor U1376 (N_1376,In_895,In_1530);
xnor U1377 (N_1377,In_2033,In_254);
nor U1378 (N_1378,In_520,In_239);
or U1379 (N_1379,In_1554,In_2002);
and U1380 (N_1380,In_817,In_1402);
nor U1381 (N_1381,In_1194,In_1108);
xor U1382 (N_1382,In_1593,In_428);
and U1383 (N_1383,In_982,In_1979);
nor U1384 (N_1384,In_1815,In_1709);
xor U1385 (N_1385,In_481,In_1854);
nand U1386 (N_1386,In_1670,In_1551);
nor U1387 (N_1387,In_586,In_1550);
nor U1388 (N_1388,In_834,In_873);
or U1389 (N_1389,In_1137,In_1013);
nor U1390 (N_1390,In_1817,In_1948);
and U1391 (N_1391,In_346,In_2488);
or U1392 (N_1392,In_2277,In_158);
or U1393 (N_1393,In_2326,In_1793);
and U1394 (N_1394,In_1943,In_767);
nor U1395 (N_1395,In_227,In_2307);
or U1396 (N_1396,In_2015,In_1411);
xor U1397 (N_1397,In_1073,In_798);
nand U1398 (N_1398,In_2264,In_1604);
nor U1399 (N_1399,In_1096,In_1534);
nand U1400 (N_1400,In_1981,In_2352);
nand U1401 (N_1401,In_1327,In_121);
and U1402 (N_1402,In_2442,In_1201);
and U1403 (N_1403,In_1513,In_1145);
nand U1404 (N_1404,In_1336,In_1787);
nand U1405 (N_1405,In_497,In_57);
nor U1406 (N_1406,In_721,In_1746);
or U1407 (N_1407,In_1893,In_1305);
or U1408 (N_1408,In_1717,In_520);
nand U1409 (N_1409,In_1744,In_720);
and U1410 (N_1410,In_145,In_1323);
or U1411 (N_1411,In_737,In_1893);
or U1412 (N_1412,In_26,In_385);
or U1413 (N_1413,In_1213,In_475);
nor U1414 (N_1414,In_667,In_519);
nor U1415 (N_1415,In_237,In_1373);
nand U1416 (N_1416,In_2186,In_1798);
nor U1417 (N_1417,In_668,In_249);
and U1418 (N_1418,In_1323,In_2219);
or U1419 (N_1419,In_1361,In_444);
or U1420 (N_1420,In_1759,In_150);
xor U1421 (N_1421,In_1228,In_1162);
or U1422 (N_1422,In_2260,In_2209);
or U1423 (N_1423,In_1886,In_1001);
and U1424 (N_1424,In_766,In_1509);
or U1425 (N_1425,In_1461,In_564);
nor U1426 (N_1426,In_2295,In_381);
and U1427 (N_1427,In_2104,In_2325);
nor U1428 (N_1428,In_1412,In_499);
xnor U1429 (N_1429,In_1323,In_795);
nor U1430 (N_1430,In_435,In_1525);
xnor U1431 (N_1431,In_1960,In_512);
nand U1432 (N_1432,In_401,In_946);
nand U1433 (N_1433,In_1083,In_549);
xnor U1434 (N_1434,In_665,In_1736);
xnor U1435 (N_1435,In_2476,In_2210);
or U1436 (N_1436,In_201,In_1940);
and U1437 (N_1437,In_1435,In_1721);
nor U1438 (N_1438,In_217,In_1727);
xnor U1439 (N_1439,In_1758,In_89);
or U1440 (N_1440,In_2067,In_372);
and U1441 (N_1441,In_9,In_2403);
and U1442 (N_1442,In_1054,In_514);
or U1443 (N_1443,In_524,In_83);
xnor U1444 (N_1444,In_1114,In_2350);
nand U1445 (N_1445,In_2230,In_391);
xnor U1446 (N_1446,In_990,In_1301);
nand U1447 (N_1447,In_1099,In_2312);
xnor U1448 (N_1448,In_903,In_1196);
or U1449 (N_1449,In_681,In_1249);
xnor U1450 (N_1450,In_1086,In_1267);
or U1451 (N_1451,In_191,In_1953);
or U1452 (N_1452,In_2433,In_262);
and U1453 (N_1453,In_1964,In_2145);
nand U1454 (N_1454,In_1951,In_2087);
or U1455 (N_1455,In_1748,In_1224);
xor U1456 (N_1456,In_659,In_382);
or U1457 (N_1457,In_710,In_408);
or U1458 (N_1458,In_170,In_2390);
nand U1459 (N_1459,In_644,In_2065);
nor U1460 (N_1460,In_103,In_1541);
and U1461 (N_1461,In_167,In_1496);
nor U1462 (N_1462,In_694,In_1194);
and U1463 (N_1463,In_1799,In_2022);
or U1464 (N_1464,In_593,In_29);
nand U1465 (N_1465,In_2492,In_434);
or U1466 (N_1466,In_1506,In_2357);
nor U1467 (N_1467,In_1500,In_595);
or U1468 (N_1468,In_210,In_1545);
nor U1469 (N_1469,In_59,In_1023);
and U1470 (N_1470,In_1010,In_1235);
nor U1471 (N_1471,In_2296,In_1348);
and U1472 (N_1472,In_2347,In_577);
nor U1473 (N_1473,In_13,In_1684);
or U1474 (N_1474,In_1995,In_938);
nand U1475 (N_1475,In_1942,In_1226);
or U1476 (N_1476,In_2457,In_1560);
nor U1477 (N_1477,In_2020,In_1859);
nor U1478 (N_1478,In_825,In_1755);
nand U1479 (N_1479,In_1226,In_2014);
or U1480 (N_1480,In_1351,In_1558);
nand U1481 (N_1481,In_2240,In_2452);
or U1482 (N_1482,In_1310,In_2429);
or U1483 (N_1483,In_1458,In_854);
or U1484 (N_1484,In_1556,In_677);
or U1485 (N_1485,In_170,In_1272);
xor U1486 (N_1486,In_2378,In_2294);
or U1487 (N_1487,In_950,In_2097);
or U1488 (N_1488,In_833,In_375);
or U1489 (N_1489,In_1739,In_272);
and U1490 (N_1490,In_2138,In_54);
xor U1491 (N_1491,In_2397,In_464);
or U1492 (N_1492,In_1055,In_1331);
nor U1493 (N_1493,In_1051,In_87);
nor U1494 (N_1494,In_1660,In_365);
nor U1495 (N_1495,In_523,In_749);
and U1496 (N_1496,In_267,In_2234);
xor U1497 (N_1497,In_2092,In_1220);
xnor U1498 (N_1498,In_2128,In_294);
or U1499 (N_1499,In_1894,In_1212);
nor U1500 (N_1500,In_2300,In_236);
nand U1501 (N_1501,In_1436,In_2279);
or U1502 (N_1502,In_1900,In_1317);
nand U1503 (N_1503,In_486,In_2294);
and U1504 (N_1504,In_1737,In_583);
and U1505 (N_1505,In_552,In_1785);
xnor U1506 (N_1506,In_1619,In_618);
and U1507 (N_1507,In_1836,In_703);
and U1508 (N_1508,In_2041,In_1645);
nand U1509 (N_1509,In_1287,In_682);
or U1510 (N_1510,In_1323,In_2072);
nor U1511 (N_1511,In_2022,In_930);
nand U1512 (N_1512,In_1749,In_2448);
or U1513 (N_1513,In_30,In_2263);
nor U1514 (N_1514,In_437,In_2262);
nand U1515 (N_1515,In_2263,In_1050);
or U1516 (N_1516,In_2145,In_2301);
nand U1517 (N_1517,In_1339,In_1406);
and U1518 (N_1518,In_513,In_1403);
or U1519 (N_1519,In_41,In_274);
and U1520 (N_1520,In_536,In_1005);
or U1521 (N_1521,In_150,In_584);
or U1522 (N_1522,In_950,In_2379);
xor U1523 (N_1523,In_681,In_297);
and U1524 (N_1524,In_1577,In_1511);
xnor U1525 (N_1525,In_342,In_377);
xnor U1526 (N_1526,In_197,In_330);
nor U1527 (N_1527,In_328,In_1143);
and U1528 (N_1528,In_1785,In_2400);
and U1529 (N_1529,In_398,In_298);
and U1530 (N_1530,In_564,In_1541);
nand U1531 (N_1531,In_1613,In_1943);
xnor U1532 (N_1532,In_511,In_2455);
xor U1533 (N_1533,In_1333,In_826);
nand U1534 (N_1534,In_2138,In_1594);
and U1535 (N_1535,In_2321,In_1825);
and U1536 (N_1536,In_547,In_2103);
nor U1537 (N_1537,In_285,In_2322);
xnor U1538 (N_1538,In_681,In_1909);
nor U1539 (N_1539,In_571,In_888);
xnor U1540 (N_1540,In_2139,In_1747);
or U1541 (N_1541,In_1048,In_1945);
and U1542 (N_1542,In_1367,In_1670);
nor U1543 (N_1543,In_2388,In_1188);
nand U1544 (N_1544,In_1040,In_1568);
or U1545 (N_1545,In_2154,In_713);
or U1546 (N_1546,In_490,In_1036);
or U1547 (N_1547,In_1769,In_654);
or U1548 (N_1548,In_1098,In_438);
or U1549 (N_1549,In_2422,In_1544);
xor U1550 (N_1550,In_1903,In_2239);
and U1551 (N_1551,In_1467,In_1763);
and U1552 (N_1552,In_172,In_18);
or U1553 (N_1553,In_516,In_763);
nor U1554 (N_1554,In_722,In_1235);
or U1555 (N_1555,In_353,In_1367);
nor U1556 (N_1556,In_1112,In_2193);
xnor U1557 (N_1557,In_1872,In_711);
xnor U1558 (N_1558,In_539,In_1045);
or U1559 (N_1559,In_143,In_1212);
and U1560 (N_1560,In_1291,In_804);
nor U1561 (N_1561,In_1709,In_375);
and U1562 (N_1562,In_194,In_1688);
or U1563 (N_1563,In_1039,In_1523);
nor U1564 (N_1564,In_584,In_1482);
nand U1565 (N_1565,In_2454,In_2244);
or U1566 (N_1566,In_1790,In_274);
or U1567 (N_1567,In_1061,In_1525);
nand U1568 (N_1568,In_1875,In_65);
nand U1569 (N_1569,In_216,In_1662);
and U1570 (N_1570,In_594,In_2223);
nor U1571 (N_1571,In_1568,In_204);
nand U1572 (N_1572,In_845,In_1174);
nand U1573 (N_1573,In_1149,In_463);
and U1574 (N_1574,In_1341,In_1368);
and U1575 (N_1575,In_2279,In_1357);
or U1576 (N_1576,In_1072,In_1185);
nor U1577 (N_1577,In_1832,In_1222);
xor U1578 (N_1578,In_1899,In_1404);
or U1579 (N_1579,In_530,In_2369);
and U1580 (N_1580,In_2179,In_754);
nor U1581 (N_1581,In_1484,In_171);
or U1582 (N_1582,In_687,In_1598);
nand U1583 (N_1583,In_951,In_1569);
nor U1584 (N_1584,In_48,In_254);
nand U1585 (N_1585,In_1695,In_615);
xnor U1586 (N_1586,In_443,In_1635);
nand U1587 (N_1587,In_2440,In_371);
xnor U1588 (N_1588,In_2417,In_962);
or U1589 (N_1589,In_1679,In_1342);
xnor U1590 (N_1590,In_1459,In_617);
nand U1591 (N_1591,In_1398,In_1009);
nand U1592 (N_1592,In_532,In_465);
and U1593 (N_1593,In_1662,In_391);
nor U1594 (N_1594,In_139,In_1657);
or U1595 (N_1595,In_921,In_1373);
xor U1596 (N_1596,In_1570,In_1240);
or U1597 (N_1597,In_2292,In_1619);
nand U1598 (N_1598,In_1321,In_1479);
or U1599 (N_1599,In_1493,In_1822);
nand U1600 (N_1600,In_1738,In_1696);
nand U1601 (N_1601,In_224,In_938);
xor U1602 (N_1602,In_600,In_426);
xor U1603 (N_1603,In_1149,In_1466);
xnor U1604 (N_1604,In_1417,In_2292);
nor U1605 (N_1605,In_867,In_1056);
and U1606 (N_1606,In_510,In_1084);
nor U1607 (N_1607,In_1025,In_956);
nor U1608 (N_1608,In_2103,In_2287);
nand U1609 (N_1609,In_952,In_788);
and U1610 (N_1610,In_2058,In_48);
nor U1611 (N_1611,In_1517,In_2427);
or U1612 (N_1612,In_642,In_1655);
and U1613 (N_1613,In_554,In_2061);
and U1614 (N_1614,In_269,In_85);
nor U1615 (N_1615,In_1297,In_240);
xnor U1616 (N_1616,In_1856,In_2130);
xor U1617 (N_1617,In_249,In_1410);
or U1618 (N_1618,In_27,In_590);
xor U1619 (N_1619,In_2318,In_399);
or U1620 (N_1620,In_2424,In_1227);
xnor U1621 (N_1621,In_499,In_1227);
nand U1622 (N_1622,In_296,In_471);
and U1623 (N_1623,In_1589,In_1411);
or U1624 (N_1624,In_8,In_1566);
nand U1625 (N_1625,In_1666,In_48);
nand U1626 (N_1626,In_759,In_509);
or U1627 (N_1627,In_2011,In_26);
nor U1628 (N_1628,In_1516,In_210);
and U1629 (N_1629,In_697,In_1157);
nand U1630 (N_1630,In_1858,In_1185);
nor U1631 (N_1631,In_1873,In_1293);
or U1632 (N_1632,In_1697,In_2460);
or U1633 (N_1633,In_829,In_631);
nand U1634 (N_1634,In_1224,In_1985);
or U1635 (N_1635,In_2005,In_9);
xnor U1636 (N_1636,In_1710,In_1563);
nand U1637 (N_1637,In_1732,In_1491);
nand U1638 (N_1638,In_1076,In_2232);
nand U1639 (N_1639,In_331,In_157);
xor U1640 (N_1640,In_1333,In_859);
xnor U1641 (N_1641,In_2015,In_1056);
xor U1642 (N_1642,In_823,In_2210);
or U1643 (N_1643,In_33,In_1071);
or U1644 (N_1644,In_1559,In_1708);
xnor U1645 (N_1645,In_1614,In_356);
nand U1646 (N_1646,In_2154,In_788);
nand U1647 (N_1647,In_694,In_1111);
or U1648 (N_1648,In_1378,In_1441);
nor U1649 (N_1649,In_1892,In_66);
nor U1650 (N_1650,In_542,In_683);
and U1651 (N_1651,In_2130,In_2418);
nand U1652 (N_1652,In_1365,In_1619);
nand U1653 (N_1653,In_2463,In_763);
and U1654 (N_1654,In_2381,In_2211);
or U1655 (N_1655,In_1926,In_505);
or U1656 (N_1656,In_1034,In_198);
and U1657 (N_1657,In_611,In_1173);
nor U1658 (N_1658,In_1273,In_1141);
and U1659 (N_1659,In_404,In_289);
or U1660 (N_1660,In_1961,In_2462);
nor U1661 (N_1661,In_2082,In_1894);
nor U1662 (N_1662,In_318,In_203);
and U1663 (N_1663,In_2195,In_419);
xor U1664 (N_1664,In_1882,In_422);
xnor U1665 (N_1665,In_1625,In_2377);
nand U1666 (N_1666,In_2306,In_2316);
or U1667 (N_1667,In_1238,In_532);
or U1668 (N_1668,In_1561,In_237);
and U1669 (N_1669,In_2106,In_1422);
xnor U1670 (N_1670,In_2167,In_1988);
and U1671 (N_1671,In_1481,In_2072);
nand U1672 (N_1672,In_252,In_1483);
nor U1673 (N_1673,In_1030,In_583);
nor U1674 (N_1674,In_1458,In_2344);
and U1675 (N_1675,In_1046,In_1403);
nand U1676 (N_1676,In_2285,In_2302);
and U1677 (N_1677,In_1734,In_1324);
nor U1678 (N_1678,In_330,In_1456);
xnor U1679 (N_1679,In_428,In_856);
xor U1680 (N_1680,In_988,In_1289);
nor U1681 (N_1681,In_656,In_1721);
and U1682 (N_1682,In_634,In_2448);
and U1683 (N_1683,In_568,In_1529);
nand U1684 (N_1684,In_520,In_1058);
or U1685 (N_1685,In_37,In_996);
xnor U1686 (N_1686,In_976,In_2122);
and U1687 (N_1687,In_181,In_262);
nor U1688 (N_1688,In_1754,In_229);
nor U1689 (N_1689,In_2272,In_2394);
xor U1690 (N_1690,In_71,In_2176);
nor U1691 (N_1691,In_1035,In_199);
nor U1692 (N_1692,In_833,In_1987);
nand U1693 (N_1693,In_2147,In_1337);
nor U1694 (N_1694,In_616,In_667);
nor U1695 (N_1695,In_734,In_215);
or U1696 (N_1696,In_2393,In_584);
nand U1697 (N_1697,In_2366,In_719);
xnor U1698 (N_1698,In_647,In_560);
and U1699 (N_1699,In_706,In_2228);
nor U1700 (N_1700,In_2326,In_876);
xor U1701 (N_1701,In_1118,In_925);
and U1702 (N_1702,In_1680,In_403);
nand U1703 (N_1703,In_403,In_359);
nor U1704 (N_1704,In_1471,In_697);
xor U1705 (N_1705,In_1232,In_1283);
and U1706 (N_1706,In_94,In_1413);
nand U1707 (N_1707,In_363,In_380);
xor U1708 (N_1708,In_1989,In_1006);
xor U1709 (N_1709,In_1680,In_2069);
and U1710 (N_1710,In_1897,In_804);
and U1711 (N_1711,In_1924,In_1601);
or U1712 (N_1712,In_1189,In_1066);
nor U1713 (N_1713,In_1467,In_2364);
xnor U1714 (N_1714,In_650,In_423);
nand U1715 (N_1715,In_1065,In_2310);
nand U1716 (N_1716,In_2314,In_1620);
nand U1717 (N_1717,In_497,In_1370);
xor U1718 (N_1718,In_64,In_1186);
or U1719 (N_1719,In_743,In_1751);
or U1720 (N_1720,In_329,In_1311);
nand U1721 (N_1721,In_2496,In_2111);
xor U1722 (N_1722,In_898,In_1133);
nand U1723 (N_1723,In_1246,In_418);
nor U1724 (N_1724,In_2242,In_2421);
nor U1725 (N_1725,In_963,In_969);
nand U1726 (N_1726,In_1790,In_1039);
or U1727 (N_1727,In_453,In_1071);
and U1728 (N_1728,In_2243,In_502);
xnor U1729 (N_1729,In_504,In_1790);
and U1730 (N_1730,In_472,In_59);
or U1731 (N_1731,In_429,In_1920);
or U1732 (N_1732,In_928,In_692);
nor U1733 (N_1733,In_2053,In_80);
nand U1734 (N_1734,In_2145,In_2348);
nor U1735 (N_1735,In_70,In_177);
or U1736 (N_1736,In_1525,In_1780);
nand U1737 (N_1737,In_415,In_1700);
nand U1738 (N_1738,In_2222,In_370);
and U1739 (N_1739,In_1017,In_1250);
or U1740 (N_1740,In_1593,In_1405);
or U1741 (N_1741,In_1192,In_119);
xor U1742 (N_1742,In_1451,In_672);
and U1743 (N_1743,In_1903,In_2132);
or U1744 (N_1744,In_1736,In_1981);
and U1745 (N_1745,In_1509,In_813);
nand U1746 (N_1746,In_139,In_1381);
nand U1747 (N_1747,In_1562,In_860);
nor U1748 (N_1748,In_2058,In_474);
xor U1749 (N_1749,In_1187,In_1501);
or U1750 (N_1750,In_1575,In_2404);
nor U1751 (N_1751,In_1726,In_724);
and U1752 (N_1752,In_1305,In_12);
nand U1753 (N_1753,In_143,In_1931);
nor U1754 (N_1754,In_1867,In_1383);
and U1755 (N_1755,In_1431,In_2477);
and U1756 (N_1756,In_2383,In_748);
xor U1757 (N_1757,In_2022,In_1354);
nor U1758 (N_1758,In_341,In_1614);
nor U1759 (N_1759,In_1082,In_32);
xnor U1760 (N_1760,In_1388,In_270);
xnor U1761 (N_1761,In_2046,In_798);
or U1762 (N_1762,In_2059,In_868);
nor U1763 (N_1763,In_342,In_66);
nor U1764 (N_1764,In_1692,In_1091);
or U1765 (N_1765,In_2037,In_2027);
xor U1766 (N_1766,In_2268,In_2067);
nor U1767 (N_1767,In_1420,In_21);
and U1768 (N_1768,In_797,In_967);
and U1769 (N_1769,In_2404,In_2239);
xor U1770 (N_1770,In_707,In_1436);
and U1771 (N_1771,In_719,In_2102);
xnor U1772 (N_1772,In_324,In_2106);
nor U1773 (N_1773,In_1576,In_460);
xnor U1774 (N_1774,In_2155,In_807);
nand U1775 (N_1775,In_1934,In_1789);
or U1776 (N_1776,In_92,In_801);
nor U1777 (N_1777,In_2223,In_1374);
and U1778 (N_1778,In_1753,In_321);
xnor U1779 (N_1779,In_2291,In_2324);
xnor U1780 (N_1780,In_2290,In_1620);
nor U1781 (N_1781,In_1126,In_451);
nand U1782 (N_1782,In_2135,In_581);
nand U1783 (N_1783,In_1786,In_2404);
nand U1784 (N_1784,In_766,In_357);
and U1785 (N_1785,In_159,In_687);
and U1786 (N_1786,In_2111,In_547);
and U1787 (N_1787,In_76,In_857);
nand U1788 (N_1788,In_2320,In_9);
and U1789 (N_1789,In_356,In_2129);
xor U1790 (N_1790,In_1080,In_906);
nand U1791 (N_1791,In_1230,In_714);
nand U1792 (N_1792,In_112,In_2434);
nand U1793 (N_1793,In_1643,In_2308);
nand U1794 (N_1794,In_1826,In_1437);
or U1795 (N_1795,In_529,In_603);
nor U1796 (N_1796,In_1205,In_1455);
xnor U1797 (N_1797,In_1876,In_149);
or U1798 (N_1798,In_2261,In_2381);
or U1799 (N_1799,In_2446,In_1160);
xor U1800 (N_1800,In_527,In_943);
xor U1801 (N_1801,In_2241,In_484);
and U1802 (N_1802,In_1209,In_1212);
nand U1803 (N_1803,In_1744,In_2097);
or U1804 (N_1804,In_241,In_664);
nand U1805 (N_1805,In_1927,In_1612);
xor U1806 (N_1806,In_2373,In_1875);
xor U1807 (N_1807,In_445,In_689);
nand U1808 (N_1808,In_164,In_700);
and U1809 (N_1809,In_1602,In_1900);
or U1810 (N_1810,In_147,In_1124);
and U1811 (N_1811,In_339,In_223);
nor U1812 (N_1812,In_2279,In_710);
nor U1813 (N_1813,In_2020,In_584);
nor U1814 (N_1814,In_1544,In_347);
xnor U1815 (N_1815,In_2304,In_1527);
nand U1816 (N_1816,In_1017,In_328);
nand U1817 (N_1817,In_112,In_1784);
nand U1818 (N_1818,In_1479,In_1888);
nor U1819 (N_1819,In_1116,In_2015);
nand U1820 (N_1820,In_2182,In_281);
or U1821 (N_1821,In_391,In_1631);
nand U1822 (N_1822,In_1573,In_939);
nor U1823 (N_1823,In_2322,In_2145);
nand U1824 (N_1824,In_2390,In_2138);
nand U1825 (N_1825,In_657,In_2244);
xor U1826 (N_1826,In_27,In_2441);
nor U1827 (N_1827,In_904,In_2490);
and U1828 (N_1828,In_1279,In_2052);
or U1829 (N_1829,In_1940,In_896);
nor U1830 (N_1830,In_1880,In_1972);
xnor U1831 (N_1831,In_1982,In_2144);
nor U1832 (N_1832,In_800,In_1500);
and U1833 (N_1833,In_2315,In_2452);
or U1834 (N_1834,In_1484,In_370);
nand U1835 (N_1835,In_460,In_1606);
and U1836 (N_1836,In_2262,In_973);
or U1837 (N_1837,In_1564,In_625);
nor U1838 (N_1838,In_923,In_2195);
or U1839 (N_1839,In_1886,In_2387);
or U1840 (N_1840,In_2458,In_768);
nand U1841 (N_1841,In_2269,In_1932);
nor U1842 (N_1842,In_753,In_1157);
xor U1843 (N_1843,In_1305,In_2374);
nand U1844 (N_1844,In_429,In_1781);
and U1845 (N_1845,In_992,In_577);
nor U1846 (N_1846,In_1084,In_794);
and U1847 (N_1847,In_1910,In_55);
xor U1848 (N_1848,In_260,In_1276);
and U1849 (N_1849,In_103,In_2417);
and U1850 (N_1850,In_1143,In_168);
nor U1851 (N_1851,In_982,In_1845);
nor U1852 (N_1852,In_2110,In_242);
nand U1853 (N_1853,In_2302,In_1004);
nor U1854 (N_1854,In_261,In_977);
nand U1855 (N_1855,In_2009,In_1918);
or U1856 (N_1856,In_1729,In_709);
or U1857 (N_1857,In_1031,In_1879);
or U1858 (N_1858,In_1066,In_161);
or U1859 (N_1859,In_31,In_2115);
nor U1860 (N_1860,In_1969,In_984);
xnor U1861 (N_1861,In_655,In_1765);
nand U1862 (N_1862,In_962,In_1215);
xor U1863 (N_1863,In_294,In_1041);
nor U1864 (N_1864,In_149,In_1626);
nor U1865 (N_1865,In_1265,In_1998);
or U1866 (N_1866,In_139,In_303);
nor U1867 (N_1867,In_1030,In_856);
nor U1868 (N_1868,In_503,In_1783);
xnor U1869 (N_1869,In_1786,In_2043);
nand U1870 (N_1870,In_740,In_1033);
nor U1871 (N_1871,In_1282,In_1838);
nand U1872 (N_1872,In_1462,In_990);
and U1873 (N_1873,In_1021,In_725);
nand U1874 (N_1874,In_2247,In_2317);
xor U1875 (N_1875,In_2189,In_2493);
nand U1876 (N_1876,In_275,In_1791);
nor U1877 (N_1877,In_1442,In_616);
nand U1878 (N_1878,In_1442,In_646);
or U1879 (N_1879,In_1747,In_2170);
nand U1880 (N_1880,In_2401,In_2370);
and U1881 (N_1881,In_2020,In_2328);
nand U1882 (N_1882,In_1785,In_378);
nand U1883 (N_1883,In_914,In_2377);
xnor U1884 (N_1884,In_1246,In_1131);
xor U1885 (N_1885,In_141,In_1801);
and U1886 (N_1886,In_509,In_704);
and U1887 (N_1887,In_599,In_693);
nand U1888 (N_1888,In_916,In_2083);
xnor U1889 (N_1889,In_607,In_0);
and U1890 (N_1890,In_1782,In_143);
or U1891 (N_1891,In_1981,In_421);
or U1892 (N_1892,In_542,In_1343);
nor U1893 (N_1893,In_273,In_2048);
nand U1894 (N_1894,In_830,In_757);
nand U1895 (N_1895,In_2301,In_355);
and U1896 (N_1896,In_2205,In_1034);
or U1897 (N_1897,In_306,In_543);
and U1898 (N_1898,In_1489,In_1542);
and U1899 (N_1899,In_1548,In_183);
nand U1900 (N_1900,In_95,In_2011);
and U1901 (N_1901,In_1170,In_2128);
nand U1902 (N_1902,In_1076,In_1203);
xnor U1903 (N_1903,In_814,In_310);
xor U1904 (N_1904,In_100,In_1398);
and U1905 (N_1905,In_1216,In_134);
xnor U1906 (N_1906,In_1840,In_1270);
and U1907 (N_1907,In_1167,In_210);
and U1908 (N_1908,In_977,In_397);
nor U1909 (N_1909,In_335,In_1911);
xor U1910 (N_1910,In_217,In_106);
or U1911 (N_1911,In_1349,In_547);
and U1912 (N_1912,In_1087,In_2100);
or U1913 (N_1913,In_89,In_1448);
nand U1914 (N_1914,In_421,In_1764);
and U1915 (N_1915,In_488,In_2171);
xor U1916 (N_1916,In_1970,In_587);
nor U1917 (N_1917,In_215,In_627);
and U1918 (N_1918,In_1352,In_2409);
nor U1919 (N_1919,In_2421,In_1637);
nand U1920 (N_1920,In_2382,In_2250);
nor U1921 (N_1921,In_1915,In_1052);
or U1922 (N_1922,In_1359,In_2081);
or U1923 (N_1923,In_975,In_1261);
nor U1924 (N_1924,In_798,In_2499);
or U1925 (N_1925,In_1122,In_825);
nand U1926 (N_1926,In_984,In_2393);
nand U1927 (N_1927,In_1981,In_2229);
nand U1928 (N_1928,In_1881,In_217);
nor U1929 (N_1929,In_260,In_2361);
or U1930 (N_1930,In_485,In_1474);
and U1931 (N_1931,In_1874,In_219);
xor U1932 (N_1932,In_1702,In_898);
or U1933 (N_1933,In_1715,In_1942);
or U1934 (N_1934,In_1344,In_2321);
nand U1935 (N_1935,In_1779,In_1320);
nor U1936 (N_1936,In_287,In_1199);
nor U1937 (N_1937,In_1648,In_58);
or U1938 (N_1938,In_1956,In_1749);
or U1939 (N_1939,In_1630,In_706);
xnor U1940 (N_1940,In_759,In_2126);
xor U1941 (N_1941,In_2088,In_1874);
and U1942 (N_1942,In_456,In_1769);
nand U1943 (N_1943,In_205,In_542);
nand U1944 (N_1944,In_2222,In_583);
or U1945 (N_1945,In_1222,In_1912);
and U1946 (N_1946,In_553,In_1966);
xor U1947 (N_1947,In_465,In_184);
or U1948 (N_1948,In_1937,In_2459);
nor U1949 (N_1949,In_1602,In_1404);
nand U1950 (N_1950,In_268,In_1968);
or U1951 (N_1951,In_909,In_422);
or U1952 (N_1952,In_880,In_1984);
xnor U1953 (N_1953,In_92,In_880);
xor U1954 (N_1954,In_1451,In_1569);
or U1955 (N_1955,In_1871,In_1943);
or U1956 (N_1956,In_666,In_2140);
nand U1957 (N_1957,In_17,In_1846);
or U1958 (N_1958,In_837,In_70);
xnor U1959 (N_1959,In_1203,In_1972);
nor U1960 (N_1960,In_1105,In_1304);
and U1961 (N_1961,In_2041,In_598);
and U1962 (N_1962,In_1451,In_2065);
and U1963 (N_1963,In_618,In_116);
nand U1964 (N_1964,In_810,In_1564);
nor U1965 (N_1965,In_363,In_1572);
or U1966 (N_1966,In_76,In_1740);
or U1967 (N_1967,In_2399,In_1420);
and U1968 (N_1968,In_1206,In_271);
nor U1969 (N_1969,In_1950,In_763);
xnor U1970 (N_1970,In_2405,In_1683);
or U1971 (N_1971,In_911,In_1413);
xnor U1972 (N_1972,In_1357,In_2090);
xor U1973 (N_1973,In_944,In_321);
or U1974 (N_1974,In_603,In_2149);
and U1975 (N_1975,In_738,In_1093);
xor U1976 (N_1976,In_57,In_29);
nand U1977 (N_1977,In_1146,In_2216);
xor U1978 (N_1978,In_993,In_1393);
nand U1979 (N_1979,In_2058,In_11);
nor U1980 (N_1980,In_732,In_1774);
nor U1981 (N_1981,In_247,In_2417);
or U1982 (N_1982,In_2402,In_1752);
or U1983 (N_1983,In_922,In_679);
nand U1984 (N_1984,In_1765,In_1419);
and U1985 (N_1985,In_2009,In_2296);
or U1986 (N_1986,In_2211,In_105);
or U1987 (N_1987,In_1121,In_2034);
and U1988 (N_1988,In_830,In_255);
xnor U1989 (N_1989,In_257,In_1220);
nand U1990 (N_1990,In_135,In_1818);
xor U1991 (N_1991,In_495,In_1138);
nor U1992 (N_1992,In_1661,In_1413);
nor U1993 (N_1993,In_108,In_1825);
nand U1994 (N_1994,In_840,In_1996);
xnor U1995 (N_1995,In_1350,In_2236);
xor U1996 (N_1996,In_744,In_900);
or U1997 (N_1997,In_372,In_1439);
xor U1998 (N_1998,In_953,In_728);
nand U1999 (N_1999,In_1529,In_1657);
or U2000 (N_2000,In_1688,In_2403);
nor U2001 (N_2001,In_2447,In_1428);
nor U2002 (N_2002,In_65,In_2170);
and U2003 (N_2003,In_2303,In_1851);
nand U2004 (N_2004,In_911,In_1627);
xnor U2005 (N_2005,In_269,In_1313);
and U2006 (N_2006,In_988,In_1582);
nor U2007 (N_2007,In_2304,In_1644);
xor U2008 (N_2008,In_545,In_851);
nand U2009 (N_2009,In_321,In_230);
nand U2010 (N_2010,In_496,In_2211);
nor U2011 (N_2011,In_1429,In_448);
nand U2012 (N_2012,In_882,In_1896);
nor U2013 (N_2013,In_204,In_486);
or U2014 (N_2014,In_1821,In_2209);
nand U2015 (N_2015,In_827,In_2325);
nor U2016 (N_2016,In_1057,In_369);
nor U2017 (N_2017,In_1707,In_2066);
and U2018 (N_2018,In_1663,In_2012);
and U2019 (N_2019,In_481,In_1985);
or U2020 (N_2020,In_334,In_2227);
nand U2021 (N_2021,In_799,In_1231);
or U2022 (N_2022,In_2351,In_311);
nand U2023 (N_2023,In_1504,In_514);
or U2024 (N_2024,In_1871,In_2351);
nor U2025 (N_2025,In_905,In_756);
xor U2026 (N_2026,In_1349,In_1291);
or U2027 (N_2027,In_1793,In_799);
and U2028 (N_2028,In_1500,In_521);
nand U2029 (N_2029,In_1366,In_2151);
and U2030 (N_2030,In_707,In_1003);
nor U2031 (N_2031,In_81,In_2410);
or U2032 (N_2032,In_98,In_368);
and U2033 (N_2033,In_2059,In_2287);
nor U2034 (N_2034,In_1349,In_1849);
and U2035 (N_2035,In_1128,In_1051);
xnor U2036 (N_2036,In_1062,In_73);
nand U2037 (N_2037,In_502,In_1101);
and U2038 (N_2038,In_2466,In_1380);
xnor U2039 (N_2039,In_760,In_973);
or U2040 (N_2040,In_1928,In_785);
nand U2041 (N_2041,In_638,In_1789);
nor U2042 (N_2042,In_871,In_1238);
nor U2043 (N_2043,In_468,In_1456);
nor U2044 (N_2044,In_96,In_2018);
nand U2045 (N_2045,In_293,In_563);
xnor U2046 (N_2046,In_845,In_2394);
nand U2047 (N_2047,In_1618,In_1340);
nor U2048 (N_2048,In_1481,In_364);
or U2049 (N_2049,In_580,In_2270);
nor U2050 (N_2050,In_626,In_255);
xnor U2051 (N_2051,In_1484,In_1151);
nor U2052 (N_2052,In_669,In_51);
nor U2053 (N_2053,In_2147,In_1768);
and U2054 (N_2054,In_1710,In_1595);
nor U2055 (N_2055,In_740,In_2256);
nor U2056 (N_2056,In_1528,In_262);
or U2057 (N_2057,In_1095,In_2453);
or U2058 (N_2058,In_2393,In_2372);
nand U2059 (N_2059,In_1359,In_803);
xor U2060 (N_2060,In_1457,In_1453);
and U2061 (N_2061,In_1818,In_416);
or U2062 (N_2062,In_2457,In_1870);
nor U2063 (N_2063,In_1844,In_361);
xnor U2064 (N_2064,In_549,In_249);
and U2065 (N_2065,In_920,In_914);
xor U2066 (N_2066,In_1186,In_1848);
and U2067 (N_2067,In_543,In_2012);
xnor U2068 (N_2068,In_1116,In_514);
xnor U2069 (N_2069,In_2264,In_1995);
nand U2070 (N_2070,In_1197,In_543);
nor U2071 (N_2071,In_952,In_2106);
nand U2072 (N_2072,In_611,In_1767);
xnor U2073 (N_2073,In_284,In_1562);
nand U2074 (N_2074,In_2474,In_305);
nand U2075 (N_2075,In_553,In_1577);
nor U2076 (N_2076,In_284,In_2099);
nand U2077 (N_2077,In_1539,In_592);
and U2078 (N_2078,In_388,In_1471);
xor U2079 (N_2079,In_1159,In_758);
nand U2080 (N_2080,In_1371,In_297);
and U2081 (N_2081,In_2286,In_1110);
xnor U2082 (N_2082,In_1217,In_1959);
nand U2083 (N_2083,In_1972,In_472);
xor U2084 (N_2084,In_1973,In_749);
and U2085 (N_2085,In_1694,In_1053);
xnor U2086 (N_2086,In_1138,In_1438);
and U2087 (N_2087,In_2315,In_1427);
or U2088 (N_2088,In_670,In_330);
xor U2089 (N_2089,In_1249,In_2474);
xor U2090 (N_2090,In_2140,In_2173);
and U2091 (N_2091,In_962,In_820);
nand U2092 (N_2092,In_1646,In_595);
nand U2093 (N_2093,In_924,In_756);
and U2094 (N_2094,In_838,In_1718);
nor U2095 (N_2095,In_273,In_158);
xnor U2096 (N_2096,In_323,In_2261);
nor U2097 (N_2097,In_2382,In_2375);
and U2098 (N_2098,In_1994,In_867);
or U2099 (N_2099,In_183,In_2424);
xnor U2100 (N_2100,In_1336,In_1532);
or U2101 (N_2101,In_2435,In_1251);
or U2102 (N_2102,In_1347,In_2206);
and U2103 (N_2103,In_225,In_1461);
nor U2104 (N_2104,In_882,In_961);
or U2105 (N_2105,In_1296,In_1422);
nand U2106 (N_2106,In_75,In_2413);
and U2107 (N_2107,In_267,In_38);
xnor U2108 (N_2108,In_2009,In_2121);
xor U2109 (N_2109,In_410,In_675);
nand U2110 (N_2110,In_1917,In_186);
nand U2111 (N_2111,In_458,In_1189);
and U2112 (N_2112,In_310,In_749);
and U2113 (N_2113,In_1917,In_343);
nand U2114 (N_2114,In_2019,In_534);
nand U2115 (N_2115,In_2201,In_1925);
or U2116 (N_2116,In_2236,In_2389);
and U2117 (N_2117,In_1375,In_398);
xor U2118 (N_2118,In_605,In_1190);
xor U2119 (N_2119,In_1679,In_194);
xor U2120 (N_2120,In_1332,In_1133);
xor U2121 (N_2121,In_4,In_2043);
or U2122 (N_2122,In_472,In_1543);
and U2123 (N_2123,In_1082,In_732);
xnor U2124 (N_2124,In_150,In_1151);
or U2125 (N_2125,In_2026,In_135);
or U2126 (N_2126,In_1721,In_2471);
xor U2127 (N_2127,In_955,In_948);
and U2128 (N_2128,In_2056,In_2291);
xnor U2129 (N_2129,In_1848,In_2084);
nor U2130 (N_2130,In_2305,In_2257);
and U2131 (N_2131,In_740,In_1136);
and U2132 (N_2132,In_1587,In_2245);
nor U2133 (N_2133,In_2425,In_2146);
xnor U2134 (N_2134,In_1565,In_122);
or U2135 (N_2135,In_2372,In_258);
xor U2136 (N_2136,In_396,In_347);
nor U2137 (N_2137,In_2013,In_391);
or U2138 (N_2138,In_1776,In_355);
and U2139 (N_2139,In_2260,In_1433);
nor U2140 (N_2140,In_221,In_936);
nor U2141 (N_2141,In_2316,In_1685);
xor U2142 (N_2142,In_1779,In_336);
and U2143 (N_2143,In_1320,In_1576);
and U2144 (N_2144,In_723,In_897);
and U2145 (N_2145,In_2217,In_1025);
and U2146 (N_2146,In_1942,In_1315);
xor U2147 (N_2147,In_425,In_1916);
xnor U2148 (N_2148,In_1346,In_1998);
or U2149 (N_2149,In_1647,In_883);
nor U2150 (N_2150,In_682,In_1262);
xor U2151 (N_2151,In_1622,In_697);
nor U2152 (N_2152,In_2171,In_1301);
and U2153 (N_2153,In_1252,In_732);
or U2154 (N_2154,In_831,In_617);
nor U2155 (N_2155,In_399,In_2456);
nand U2156 (N_2156,In_286,In_926);
or U2157 (N_2157,In_639,In_459);
and U2158 (N_2158,In_2470,In_2051);
or U2159 (N_2159,In_1654,In_1102);
nand U2160 (N_2160,In_1241,In_524);
nand U2161 (N_2161,In_1422,In_2107);
xnor U2162 (N_2162,In_1886,In_1237);
nor U2163 (N_2163,In_452,In_1328);
or U2164 (N_2164,In_2430,In_1079);
and U2165 (N_2165,In_155,In_668);
xnor U2166 (N_2166,In_731,In_1755);
nor U2167 (N_2167,In_1423,In_572);
xnor U2168 (N_2168,In_426,In_1930);
xnor U2169 (N_2169,In_2325,In_1924);
nand U2170 (N_2170,In_1318,In_1726);
nor U2171 (N_2171,In_1186,In_1788);
or U2172 (N_2172,In_947,In_755);
or U2173 (N_2173,In_1011,In_898);
or U2174 (N_2174,In_2361,In_866);
and U2175 (N_2175,In_1092,In_513);
nand U2176 (N_2176,In_2142,In_912);
xor U2177 (N_2177,In_1565,In_2145);
and U2178 (N_2178,In_59,In_251);
nand U2179 (N_2179,In_690,In_2291);
xnor U2180 (N_2180,In_2385,In_1131);
or U2181 (N_2181,In_1122,In_309);
xnor U2182 (N_2182,In_118,In_2426);
nor U2183 (N_2183,In_797,In_672);
xor U2184 (N_2184,In_1205,In_959);
or U2185 (N_2185,In_2352,In_1642);
nand U2186 (N_2186,In_285,In_780);
and U2187 (N_2187,In_553,In_2225);
nor U2188 (N_2188,In_908,In_777);
nand U2189 (N_2189,In_1496,In_1026);
or U2190 (N_2190,In_570,In_1528);
or U2191 (N_2191,In_1492,In_680);
xnor U2192 (N_2192,In_2134,In_103);
nor U2193 (N_2193,In_1876,In_489);
or U2194 (N_2194,In_1527,In_1592);
nand U2195 (N_2195,In_1697,In_1534);
nor U2196 (N_2196,In_751,In_837);
and U2197 (N_2197,In_1826,In_2132);
nand U2198 (N_2198,In_24,In_2425);
nor U2199 (N_2199,In_767,In_1270);
or U2200 (N_2200,In_318,In_549);
or U2201 (N_2201,In_279,In_1352);
xnor U2202 (N_2202,In_29,In_134);
or U2203 (N_2203,In_2175,In_1145);
and U2204 (N_2204,In_215,In_4);
and U2205 (N_2205,In_1415,In_31);
nand U2206 (N_2206,In_1494,In_413);
and U2207 (N_2207,In_138,In_1906);
or U2208 (N_2208,In_753,In_1750);
and U2209 (N_2209,In_10,In_710);
nor U2210 (N_2210,In_584,In_691);
nand U2211 (N_2211,In_530,In_897);
nor U2212 (N_2212,In_1052,In_758);
xor U2213 (N_2213,In_131,In_2481);
nor U2214 (N_2214,In_1726,In_186);
xor U2215 (N_2215,In_490,In_1485);
nand U2216 (N_2216,In_241,In_1646);
nand U2217 (N_2217,In_1807,In_1472);
xnor U2218 (N_2218,In_51,In_2435);
xnor U2219 (N_2219,In_1623,In_2128);
and U2220 (N_2220,In_651,In_1637);
xnor U2221 (N_2221,In_2326,In_175);
nand U2222 (N_2222,In_2403,In_1270);
or U2223 (N_2223,In_1641,In_2094);
nor U2224 (N_2224,In_1974,In_2152);
nand U2225 (N_2225,In_1186,In_375);
nand U2226 (N_2226,In_249,In_157);
nor U2227 (N_2227,In_1579,In_2149);
or U2228 (N_2228,In_19,In_1620);
and U2229 (N_2229,In_1202,In_843);
and U2230 (N_2230,In_1879,In_534);
xnor U2231 (N_2231,In_1765,In_406);
and U2232 (N_2232,In_648,In_686);
nand U2233 (N_2233,In_1949,In_282);
nand U2234 (N_2234,In_767,In_2129);
or U2235 (N_2235,In_2062,In_813);
and U2236 (N_2236,In_1783,In_2280);
nor U2237 (N_2237,In_1403,In_621);
nor U2238 (N_2238,In_679,In_476);
nor U2239 (N_2239,In_294,In_483);
or U2240 (N_2240,In_843,In_846);
and U2241 (N_2241,In_1859,In_1523);
nand U2242 (N_2242,In_2358,In_1844);
or U2243 (N_2243,In_2198,In_2293);
nor U2244 (N_2244,In_201,In_1871);
and U2245 (N_2245,In_1505,In_280);
and U2246 (N_2246,In_2355,In_1871);
nand U2247 (N_2247,In_383,In_884);
nand U2248 (N_2248,In_2482,In_1410);
or U2249 (N_2249,In_404,In_666);
nand U2250 (N_2250,In_290,In_912);
and U2251 (N_2251,In_1823,In_347);
nand U2252 (N_2252,In_712,In_1496);
xor U2253 (N_2253,In_2430,In_1610);
and U2254 (N_2254,In_2154,In_667);
or U2255 (N_2255,In_1131,In_1722);
and U2256 (N_2256,In_400,In_305);
or U2257 (N_2257,In_375,In_1759);
and U2258 (N_2258,In_1460,In_822);
nor U2259 (N_2259,In_643,In_1726);
xnor U2260 (N_2260,In_1041,In_2151);
nor U2261 (N_2261,In_1909,In_582);
and U2262 (N_2262,In_1846,In_1999);
or U2263 (N_2263,In_1780,In_784);
nand U2264 (N_2264,In_179,In_892);
nor U2265 (N_2265,In_1777,In_788);
nand U2266 (N_2266,In_1091,In_738);
nor U2267 (N_2267,In_2213,In_2289);
nand U2268 (N_2268,In_237,In_1648);
nand U2269 (N_2269,In_1620,In_919);
nand U2270 (N_2270,In_595,In_34);
nand U2271 (N_2271,In_1866,In_2061);
and U2272 (N_2272,In_1432,In_1328);
or U2273 (N_2273,In_1226,In_1921);
nand U2274 (N_2274,In_924,In_451);
and U2275 (N_2275,In_724,In_1353);
nand U2276 (N_2276,In_1337,In_645);
xor U2277 (N_2277,In_367,In_1146);
xnor U2278 (N_2278,In_838,In_1087);
or U2279 (N_2279,In_887,In_1307);
and U2280 (N_2280,In_769,In_914);
and U2281 (N_2281,In_471,In_1454);
nand U2282 (N_2282,In_1492,In_2348);
or U2283 (N_2283,In_1927,In_645);
nand U2284 (N_2284,In_1418,In_916);
nor U2285 (N_2285,In_2225,In_1475);
nor U2286 (N_2286,In_1789,In_2250);
or U2287 (N_2287,In_93,In_1416);
or U2288 (N_2288,In_408,In_1309);
nand U2289 (N_2289,In_1306,In_633);
or U2290 (N_2290,In_1446,In_1309);
and U2291 (N_2291,In_1123,In_330);
and U2292 (N_2292,In_786,In_754);
nor U2293 (N_2293,In_260,In_2218);
nand U2294 (N_2294,In_503,In_2460);
xnor U2295 (N_2295,In_741,In_1525);
or U2296 (N_2296,In_2313,In_329);
nand U2297 (N_2297,In_2245,In_553);
nor U2298 (N_2298,In_1021,In_2071);
xnor U2299 (N_2299,In_1478,In_946);
nor U2300 (N_2300,In_464,In_1750);
nand U2301 (N_2301,In_1820,In_1650);
and U2302 (N_2302,In_294,In_257);
nor U2303 (N_2303,In_743,In_1294);
nor U2304 (N_2304,In_1695,In_2160);
and U2305 (N_2305,In_680,In_650);
nor U2306 (N_2306,In_1676,In_1335);
nand U2307 (N_2307,In_451,In_2222);
nor U2308 (N_2308,In_1483,In_1043);
nand U2309 (N_2309,In_2172,In_1361);
xnor U2310 (N_2310,In_2441,In_1067);
xnor U2311 (N_2311,In_1638,In_706);
xnor U2312 (N_2312,In_923,In_2080);
xnor U2313 (N_2313,In_782,In_1098);
nor U2314 (N_2314,In_2197,In_993);
nand U2315 (N_2315,In_1837,In_2158);
nand U2316 (N_2316,In_1650,In_1546);
nand U2317 (N_2317,In_744,In_177);
xnor U2318 (N_2318,In_1084,In_2417);
and U2319 (N_2319,In_1480,In_1277);
nand U2320 (N_2320,In_108,In_1750);
nand U2321 (N_2321,In_1697,In_2030);
xor U2322 (N_2322,In_806,In_335);
xnor U2323 (N_2323,In_2021,In_1599);
or U2324 (N_2324,In_747,In_477);
or U2325 (N_2325,In_1009,In_1253);
nor U2326 (N_2326,In_1366,In_987);
nand U2327 (N_2327,In_2445,In_2355);
nand U2328 (N_2328,In_1219,In_124);
nor U2329 (N_2329,In_1294,In_488);
or U2330 (N_2330,In_871,In_1692);
or U2331 (N_2331,In_145,In_2351);
nand U2332 (N_2332,In_852,In_1830);
nand U2333 (N_2333,In_684,In_1626);
nand U2334 (N_2334,In_322,In_1717);
nand U2335 (N_2335,In_2090,In_192);
or U2336 (N_2336,In_233,In_339);
xnor U2337 (N_2337,In_238,In_1141);
xor U2338 (N_2338,In_1480,In_581);
xnor U2339 (N_2339,In_234,In_1483);
nand U2340 (N_2340,In_833,In_598);
nand U2341 (N_2341,In_1061,In_285);
nor U2342 (N_2342,In_1261,In_619);
or U2343 (N_2343,In_1276,In_189);
and U2344 (N_2344,In_2003,In_531);
nand U2345 (N_2345,In_1290,In_1225);
xnor U2346 (N_2346,In_306,In_2221);
and U2347 (N_2347,In_1336,In_965);
or U2348 (N_2348,In_2138,In_618);
and U2349 (N_2349,In_1214,In_1949);
and U2350 (N_2350,In_1770,In_572);
nor U2351 (N_2351,In_875,In_1762);
nor U2352 (N_2352,In_2371,In_648);
nor U2353 (N_2353,In_1916,In_454);
and U2354 (N_2354,In_620,In_763);
or U2355 (N_2355,In_2424,In_11);
xnor U2356 (N_2356,In_2095,In_2288);
xnor U2357 (N_2357,In_43,In_2252);
and U2358 (N_2358,In_237,In_847);
or U2359 (N_2359,In_1661,In_1682);
and U2360 (N_2360,In_2150,In_594);
xnor U2361 (N_2361,In_1941,In_953);
nand U2362 (N_2362,In_637,In_136);
xnor U2363 (N_2363,In_1611,In_1229);
and U2364 (N_2364,In_2198,In_2179);
nor U2365 (N_2365,In_452,In_1694);
and U2366 (N_2366,In_1839,In_1661);
nand U2367 (N_2367,In_1103,In_398);
or U2368 (N_2368,In_2013,In_961);
and U2369 (N_2369,In_1534,In_2447);
xnor U2370 (N_2370,In_1181,In_341);
and U2371 (N_2371,In_1122,In_2441);
xor U2372 (N_2372,In_2038,In_1246);
or U2373 (N_2373,In_2103,In_2080);
and U2374 (N_2374,In_810,In_436);
nand U2375 (N_2375,In_43,In_1990);
nand U2376 (N_2376,In_1893,In_465);
xnor U2377 (N_2377,In_2023,In_1830);
and U2378 (N_2378,In_2340,In_1636);
nand U2379 (N_2379,In_543,In_938);
and U2380 (N_2380,In_527,In_1882);
and U2381 (N_2381,In_103,In_455);
nor U2382 (N_2382,In_1069,In_2301);
and U2383 (N_2383,In_680,In_17);
nand U2384 (N_2384,In_1887,In_2252);
xor U2385 (N_2385,In_953,In_49);
nand U2386 (N_2386,In_993,In_2279);
nand U2387 (N_2387,In_305,In_1572);
nand U2388 (N_2388,In_2087,In_510);
nor U2389 (N_2389,In_712,In_33);
and U2390 (N_2390,In_2130,In_1677);
nor U2391 (N_2391,In_1971,In_972);
or U2392 (N_2392,In_1535,In_1870);
nor U2393 (N_2393,In_1499,In_1220);
xor U2394 (N_2394,In_2013,In_1933);
xor U2395 (N_2395,In_1558,In_512);
nor U2396 (N_2396,In_2261,In_683);
or U2397 (N_2397,In_2060,In_1053);
or U2398 (N_2398,In_1899,In_2257);
nand U2399 (N_2399,In_54,In_642);
or U2400 (N_2400,In_198,In_2267);
xnor U2401 (N_2401,In_2198,In_1674);
nand U2402 (N_2402,In_549,In_1955);
nand U2403 (N_2403,In_740,In_858);
nand U2404 (N_2404,In_497,In_988);
or U2405 (N_2405,In_976,In_1330);
or U2406 (N_2406,In_1864,In_15);
nand U2407 (N_2407,In_218,In_5);
or U2408 (N_2408,In_497,In_2428);
nand U2409 (N_2409,In_1849,In_2355);
nor U2410 (N_2410,In_2380,In_684);
nor U2411 (N_2411,In_427,In_770);
nand U2412 (N_2412,In_1746,In_1186);
or U2413 (N_2413,In_2076,In_1851);
nor U2414 (N_2414,In_1536,In_1548);
and U2415 (N_2415,In_204,In_1186);
or U2416 (N_2416,In_404,In_417);
xor U2417 (N_2417,In_866,In_2113);
and U2418 (N_2418,In_524,In_672);
and U2419 (N_2419,In_1957,In_1981);
nor U2420 (N_2420,In_2010,In_756);
nor U2421 (N_2421,In_344,In_1721);
nand U2422 (N_2422,In_26,In_1828);
and U2423 (N_2423,In_1043,In_549);
and U2424 (N_2424,In_1979,In_1131);
and U2425 (N_2425,In_92,In_377);
xor U2426 (N_2426,In_1497,In_652);
nand U2427 (N_2427,In_864,In_2031);
nor U2428 (N_2428,In_2005,In_374);
and U2429 (N_2429,In_1804,In_1709);
nand U2430 (N_2430,In_949,In_2324);
nor U2431 (N_2431,In_1316,In_1802);
or U2432 (N_2432,In_1632,In_1174);
xor U2433 (N_2433,In_1802,In_89);
nor U2434 (N_2434,In_728,In_713);
or U2435 (N_2435,In_195,In_250);
and U2436 (N_2436,In_987,In_1064);
xor U2437 (N_2437,In_2137,In_2214);
or U2438 (N_2438,In_1068,In_2078);
nor U2439 (N_2439,In_1667,In_870);
and U2440 (N_2440,In_587,In_2322);
xnor U2441 (N_2441,In_290,In_571);
or U2442 (N_2442,In_1424,In_1955);
and U2443 (N_2443,In_1320,In_603);
xor U2444 (N_2444,In_2450,In_281);
nand U2445 (N_2445,In_2162,In_129);
nand U2446 (N_2446,In_1852,In_784);
and U2447 (N_2447,In_917,In_461);
and U2448 (N_2448,In_1633,In_1437);
xor U2449 (N_2449,In_1904,In_290);
xor U2450 (N_2450,In_1229,In_2178);
and U2451 (N_2451,In_706,In_520);
xnor U2452 (N_2452,In_1620,In_152);
nand U2453 (N_2453,In_2101,In_1825);
xor U2454 (N_2454,In_1418,In_338);
xnor U2455 (N_2455,In_158,In_824);
xnor U2456 (N_2456,In_676,In_738);
xor U2457 (N_2457,In_834,In_2394);
xnor U2458 (N_2458,In_1893,In_1004);
or U2459 (N_2459,In_872,In_1503);
nor U2460 (N_2460,In_1027,In_78);
nand U2461 (N_2461,In_214,In_1173);
xor U2462 (N_2462,In_2201,In_1033);
xnor U2463 (N_2463,In_2470,In_490);
or U2464 (N_2464,In_2091,In_1543);
nand U2465 (N_2465,In_1548,In_1104);
nand U2466 (N_2466,In_1979,In_362);
xor U2467 (N_2467,In_1485,In_1068);
xor U2468 (N_2468,In_2329,In_437);
xor U2469 (N_2469,In_1634,In_1245);
and U2470 (N_2470,In_2025,In_2347);
and U2471 (N_2471,In_2450,In_529);
and U2472 (N_2472,In_1739,In_1274);
or U2473 (N_2473,In_2211,In_525);
and U2474 (N_2474,In_1189,In_878);
and U2475 (N_2475,In_1477,In_2429);
xor U2476 (N_2476,In_584,In_2058);
and U2477 (N_2477,In_1637,In_1839);
nand U2478 (N_2478,In_472,In_298);
nand U2479 (N_2479,In_1266,In_1205);
nand U2480 (N_2480,In_756,In_2324);
xnor U2481 (N_2481,In_242,In_1033);
and U2482 (N_2482,In_1364,In_2196);
xnor U2483 (N_2483,In_1192,In_1579);
nor U2484 (N_2484,In_1694,In_496);
nand U2485 (N_2485,In_716,In_5);
or U2486 (N_2486,In_184,In_1613);
xnor U2487 (N_2487,In_277,In_1021);
and U2488 (N_2488,In_2356,In_517);
and U2489 (N_2489,In_1372,In_2039);
xnor U2490 (N_2490,In_1254,In_509);
nor U2491 (N_2491,In_1396,In_495);
or U2492 (N_2492,In_297,In_1867);
and U2493 (N_2493,In_1799,In_372);
and U2494 (N_2494,In_1144,In_946);
nand U2495 (N_2495,In_211,In_474);
or U2496 (N_2496,In_204,In_2294);
xnor U2497 (N_2497,In_496,In_1792);
and U2498 (N_2498,In_810,In_466);
and U2499 (N_2499,In_2311,In_2262);
nand U2500 (N_2500,In_1017,In_147);
or U2501 (N_2501,In_448,In_1135);
xnor U2502 (N_2502,In_2279,In_1112);
nor U2503 (N_2503,In_2401,In_1605);
or U2504 (N_2504,In_784,In_262);
nand U2505 (N_2505,In_1106,In_1297);
and U2506 (N_2506,In_334,In_1352);
xnor U2507 (N_2507,In_1436,In_1266);
xnor U2508 (N_2508,In_197,In_1916);
and U2509 (N_2509,In_443,In_538);
or U2510 (N_2510,In_340,In_179);
xnor U2511 (N_2511,In_2159,In_1456);
xnor U2512 (N_2512,In_2418,In_1047);
and U2513 (N_2513,In_2327,In_2127);
xnor U2514 (N_2514,In_2336,In_514);
nand U2515 (N_2515,In_837,In_1884);
nor U2516 (N_2516,In_1755,In_996);
and U2517 (N_2517,In_1004,In_1434);
nor U2518 (N_2518,In_2324,In_1823);
nand U2519 (N_2519,In_616,In_158);
or U2520 (N_2520,In_1919,In_1710);
xor U2521 (N_2521,In_2396,In_1600);
xnor U2522 (N_2522,In_1935,In_1527);
or U2523 (N_2523,In_505,In_774);
nand U2524 (N_2524,In_349,In_135);
and U2525 (N_2525,In_505,In_1872);
nand U2526 (N_2526,In_1899,In_2078);
or U2527 (N_2527,In_360,In_729);
nand U2528 (N_2528,In_103,In_1471);
or U2529 (N_2529,In_440,In_506);
nand U2530 (N_2530,In_401,In_1781);
nand U2531 (N_2531,In_1282,In_1391);
or U2532 (N_2532,In_1137,In_2000);
and U2533 (N_2533,In_347,In_1280);
xnor U2534 (N_2534,In_1558,In_664);
or U2535 (N_2535,In_1298,In_1702);
nand U2536 (N_2536,In_852,In_1836);
or U2537 (N_2537,In_723,In_905);
nor U2538 (N_2538,In_1105,In_978);
nor U2539 (N_2539,In_1881,In_1048);
and U2540 (N_2540,In_1748,In_2374);
and U2541 (N_2541,In_2235,In_1625);
and U2542 (N_2542,In_6,In_1436);
and U2543 (N_2543,In_1040,In_1675);
nor U2544 (N_2544,In_1264,In_372);
and U2545 (N_2545,In_1041,In_1888);
xor U2546 (N_2546,In_1535,In_2090);
nor U2547 (N_2547,In_13,In_1489);
nand U2548 (N_2548,In_989,In_2127);
nor U2549 (N_2549,In_2406,In_934);
nand U2550 (N_2550,In_1113,In_646);
xor U2551 (N_2551,In_1731,In_970);
nand U2552 (N_2552,In_1215,In_1844);
xnor U2553 (N_2553,In_2224,In_2216);
nand U2554 (N_2554,In_1973,In_1065);
nand U2555 (N_2555,In_2155,In_1204);
xnor U2556 (N_2556,In_503,In_626);
xor U2557 (N_2557,In_1510,In_1584);
or U2558 (N_2558,In_956,In_1065);
xnor U2559 (N_2559,In_475,In_1396);
nor U2560 (N_2560,In_2086,In_514);
xor U2561 (N_2561,In_1918,In_170);
xnor U2562 (N_2562,In_124,In_1948);
or U2563 (N_2563,In_749,In_384);
and U2564 (N_2564,In_1781,In_834);
nand U2565 (N_2565,In_290,In_927);
and U2566 (N_2566,In_795,In_1610);
and U2567 (N_2567,In_833,In_2034);
nor U2568 (N_2568,In_1730,In_2182);
nand U2569 (N_2569,In_917,In_1742);
nand U2570 (N_2570,In_1286,In_510);
and U2571 (N_2571,In_202,In_1304);
and U2572 (N_2572,In_2172,In_1906);
and U2573 (N_2573,In_1025,In_1709);
nor U2574 (N_2574,In_128,In_1991);
and U2575 (N_2575,In_775,In_2092);
and U2576 (N_2576,In_866,In_1626);
and U2577 (N_2577,In_1784,In_117);
and U2578 (N_2578,In_656,In_331);
or U2579 (N_2579,In_1996,In_1143);
xor U2580 (N_2580,In_2052,In_1484);
nor U2581 (N_2581,In_658,In_2114);
and U2582 (N_2582,In_1135,In_1862);
nor U2583 (N_2583,In_2245,In_1648);
nand U2584 (N_2584,In_611,In_320);
and U2585 (N_2585,In_279,In_2251);
nor U2586 (N_2586,In_1379,In_539);
nor U2587 (N_2587,In_2049,In_2050);
or U2588 (N_2588,In_2019,In_2008);
and U2589 (N_2589,In_890,In_17);
xor U2590 (N_2590,In_1677,In_1357);
xor U2591 (N_2591,In_814,In_1176);
or U2592 (N_2592,In_1876,In_1218);
xor U2593 (N_2593,In_290,In_2455);
xnor U2594 (N_2594,In_1586,In_2097);
xnor U2595 (N_2595,In_470,In_1366);
or U2596 (N_2596,In_1338,In_352);
xnor U2597 (N_2597,In_1026,In_731);
and U2598 (N_2598,In_70,In_2297);
or U2599 (N_2599,In_1005,In_716);
and U2600 (N_2600,In_407,In_1572);
nor U2601 (N_2601,In_892,In_2051);
or U2602 (N_2602,In_1589,In_734);
nor U2603 (N_2603,In_1526,In_187);
xnor U2604 (N_2604,In_1621,In_930);
and U2605 (N_2605,In_747,In_234);
or U2606 (N_2606,In_1781,In_1730);
or U2607 (N_2607,In_729,In_188);
and U2608 (N_2608,In_1777,In_1485);
nor U2609 (N_2609,In_177,In_851);
and U2610 (N_2610,In_1314,In_1829);
and U2611 (N_2611,In_2307,In_1793);
and U2612 (N_2612,In_696,In_570);
nand U2613 (N_2613,In_991,In_1492);
nand U2614 (N_2614,In_596,In_599);
nand U2615 (N_2615,In_1748,In_275);
nand U2616 (N_2616,In_318,In_1777);
or U2617 (N_2617,In_742,In_1380);
or U2618 (N_2618,In_1905,In_752);
xor U2619 (N_2619,In_1579,In_2469);
and U2620 (N_2620,In_2118,In_2190);
and U2621 (N_2621,In_2176,In_2262);
nand U2622 (N_2622,In_812,In_2279);
nand U2623 (N_2623,In_893,In_1185);
xnor U2624 (N_2624,In_1459,In_2189);
xnor U2625 (N_2625,In_351,In_2097);
xor U2626 (N_2626,In_1909,In_831);
and U2627 (N_2627,In_2048,In_1216);
xnor U2628 (N_2628,In_748,In_763);
or U2629 (N_2629,In_908,In_2087);
or U2630 (N_2630,In_817,In_1950);
or U2631 (N_2631,In_1961,In_1620);
xor U2632 (N_2632,In_1058,In_2304);
or U2633 (N_2633,In_1367,In_413);
or U2634 (N_2634,In_768,In_637);
or U2635 (N_2635,In_459,In_751);
and U2636 (N_2636,In_1725,In_1351);
or U2637 (N_2637,In_387,In_2230);
nor U2638 (N_2638,In_2420,In_1402);
nor U2639 (N_2639,In_1655,In_1628);
xnor U2640 (N_2640,In_1602,In_478);
and U2641 (N_2641,In_1091,In_2084);
nor U2642 (N_2642,In_863,In_2143);
or U2643 (N_2643,In_2136,In_435);
nor U2644 (N_2644,In_1885,In_1642);
nor U2645 (N_2645,In_1546,In_647);
or U2646 (N_2646,In_281,In_1810);
xor U2647 (N_2647,In_810,In_1677);
or U2648 (N_2648,In_1253,In_96);
or U2649 (N_2649,In_204,In_360);
xor U2650 (N_2650,In_46,In_141);
xor U2651 (N_2651,In_331,In_818);
nor U2652 (N_2652,In_202,In_2175);
or U2653 (N_2653,In_635,In_861);
or U2654 (N_2654,In_686,In_637);
or U2655 (N_2655,In_1591,In_1174);
and U2656 (N_2656,In_1598,In_1102);
or U2657 (N_2657,In_2466,In_1022);
nand U2658 (N_2658,In_1241,In_824);
or U2659 (N_2659,In_545,In_40);
nand U2660 (N_2660,In_1486,In_1952);
and U2661 (N_2661,In_2318,In_1542);
nor U2662 (N_2662,In_1479,In_1883);
or U2663 (N_2663,In_1038,In_2467);
nor U2664 (N_2664,In_1596,In_1083);
nor U2665 (N_2665,In_1000,In_866);
or U2666 (N_2666,In_1977,In_2466);
and U2667 (N_2667,In_840,In_351);
or U2668 (N_2668,In_1055,In_1642);
xnor U2669 (N_2669,In_2213,In_2263);
xnor U2670 (N_2670,In_1368,In_949);
nor U2671 (N_2671,In_336,In_266);
nor U2672 (N_2672,In_700,In_229);
and U2673 (N_2673,In_1330,In_1614);
or U2674 (N_2674,In_1549,In_114);
and U2675 (N_2675,In_496,In_814);
and U2676 (N_2676,In_2148,In_2128);
or U2677 (N_2677,In_895,In_2261);
nor U2678 (N_2678,In_2393,In_2112);
xor U2679 (N_2679,In_1861,In_1033);
xnor U2680 (N_2680,In_2171,In_1833);
nor U2681 (N_2681,In_1937,In_366);
xor U2682 (N_2682,In_563,In_626);
and U2683 (N_2683,In_304,In_2415);
and U2684 (N_2684,In_705,In_1408);
nor U2685 (N_2685,In_212,In_877);
nor U2686 (N_2686,In_144,In_782);
or U2687 (N_2687,In_1295,In_1425);
nor U2688 (N_2688,In_565,In_1703);
or U2689 (N_2689,In_140,In_2377);
nor U2690 (N_2690,In_927,In_1153);
and U2691 (N_2691,In_1991,In_1116);
nor U2692 (N_2692,In_1503,In_1969);
nor U2693 (N_2693,In_1258,In_937);
xor U2694 (N_2694,In_2282,In_478);
nand U2695 (N_2695,In_1245,In_201);
and U2696 (N_2696,In_1933,In_2192);
and U2697 (N_2697,In_2046,In_1609);
nand U2698 (N_2698,In_2481,In_1377);
and U2699 (N_2699,In_1120,In_2125);
nor U2700 (N_2700,In_1504,In_2239);
and U2701 (N_2701,In_809,In_950);
and U2702 (N_2702,In_2311,In_222);
or U2703 (N_2703,In_1732,In_1253);
xor U2704 (N_2704,In_1517,In_2234);
or U2705 (N_2705,In_374,In_1313);
or U2706 (N_2706,In_1785,In_184);
and U2707 (N_2707,In_893,In_2234);
and U2708 (N_2708,In_2251,In_1198);
xor U2709 (N_2709,In_2236,In_640);
nand U2710 (N_2710,In_281,In_243);
nand U2711 (N_2711,In_508,In_2021);
nor U2712 (N_2712,In_2092,In_2225);
nor U2713 (N_2713,In_1581,In_14);
or U2714 (N_2714,In_2281,In_808);
or U2715 (N_2715,In_693,In_2139);
or U2716 (N_2716,In_1706,In_435);
and U2717 (N_2717,In_2328,In_2482);
xnor U2718 (N_2718,In_1147,In_162);
and U2719 (N_2719,In_2398,In_2300);
nor U2720 (N_2720,In_18,In_229);
nand U2721 (N_2721,In_1258,In_525);
and U2722 (N_2722,In_2346,In_2044);
nand U2723 (N_2723,In_1466,In_895);
and U2724 (N_2724,In_792,In_2008);
xor U2725 (N_2725,In_1532,In_1401);
nand U2726 (N_2726,In_2399,In_8);
or U2727 (N_2727,In_32,In_909);
and U2728 (N_2728,In_2320,In_1174);
and U2729 (N_2729,In_765,In_1475);
nor U2730 (N_2730,In_2295,In_170);
nor U2731 (N_2731,In_1517,In_1788);
nand U2732 (N_2732,In_1368,In_2207);
xor U2733 (N_2733,In_2,In_1615);
nor U2734 (N_2734,In_636,In_927);
and U2735 (N_2735,In_1401,In_26);
or U2736 (N_2736,In_1965,In_1218);
nand U2737 (N_2737,In_2282,In_1560);
nand U2738 (N_2738,In_557,In_1749);
nor U2739 (N_2739,In_958,In_1243);
nor U2740 (N_2740,In_1066,In_1404);
and U2741 (N_2741,In_888,In_1861);
or U2742 (N_2742,In_1540,In_203);
nand U2743 (N_2743,In_79,In_2435);
or U2744 (N_2744,In_960,In_405);
xnor U2745 (N_2745,In_543,In_552);
nand U2746 (N_2746,In_674,In_421);
or U2747 (N_2747,In_187,In_1690);
or U2748 (N_2748,In_477,In_249);
nor U2749 (N_2749,In_95,In_295);
or U2750 (N_2750,In_612,In_2113);
xnor U2751 (N_2751,In_308,In_40);
nand U2752 (N_2752,In_551,In_162);
xor U2753 (N_2753,In_2473,In_1351);
and U2754 (N_2754,In_1535,In_1635);
nor U2755 (N_2755,In_1768,In_1863);
nor U2756 (N_2756,In_2054,In_2375);
nor U2757 (N_2757,In_1933,In_1798);
nand U2758 (N_2758,In_1466,In_2005);
xnor U2759 (N_2759,In_102,In_1662);
or U2760 (N_2760,In_348,In_30);
nor U2761 (N_2761,In_1428,In_1616);
xnor U2762 (N_2762,In_1360,In_1285);
or U2763 (N_2763,In_2301,In_1095);
or U2764 (N_2764,In_2208,In_1482);
xnor U2765 (N_2765,In_1718,In_1409);
nor U2766 (N_2766,In_1840,In_967);
nand U2767 (N_2767,In_61,In_1777);
nand U2768 (N_2768,In_763,In_1062);
and U2769 (N_2769,In_698,In_1502);
xor U2770 (N_2770,In_1245,In_517);
xnor U2771 (N_2771,In_1042,In_1451);
and U2772 (N_2772,In_1122,In_237);
xor U2773 (N_2773,In_2394,In_1591);
and U2774 (N_2774,In_2231,In_2209);
or U2775 (N_2775,In_270,In_1698);
nor U2776 (N_2776,In_1306,In_959);
nand U2777 (N_2777,In_1602,In_1525);
and U2778 (N_2778,In_1223,In_654);
nor U2779 (N_2779,In_1443,In_1163);
nor U2780 (N_2780,In_2103,In_473);
nor U2781 (N_2781,In_1053,In_1945);
and U2782 (N_2782,In_1319,In_1924);
nor U2783 (N_2783,In_2035,In_2354);
nand U2784 (N_2784,In_1108,In_204);
nand U2785 (N_2785,In_1529,In_860);
xor U2786 (N_2786,In_137,In_2452);
nand U2787 (N_2787,In_1050,In_2454);
and U2788 (N_2788,In_528,In_1422);
nand U2789 (N_2789,In_666,In_1640);
and U2790 (N_2790,In_374,In_1607);
and U2791 (N_2791,In_1279,In_328);
or U2792 (N_2792,In_1662,In_1215);
and U2793 (N_2793,In_2265,In_1521);
nor U2794 (N_2794,In_2354,In_18);
nor U2795 (N_2795,In_158,In_349);
or U2796 (N_2796,In_343,In_1912);
nor U2797 (N_2797,In_2405,In_2135);
nand U2798 (N_2798,In_2243,In_2075);
nand U2799 (N_2799,In_1365,In_734);
or U2800 (N_2800,In_450,In_632);
or U2801 (N_2801,In_1798,In_251);
xor U2802 (N_2802,In_1523,In_1433);
or U2803 (N_2803,In_2059,In_650);
nor U2804 (N_2804,In_2082,In_96);
nand U2805 (N_2805,In_2127,In_2139);
or U2806 (N_2806,In_1386,In_310);
nand U2807 (N_2807,In_298,In_1160);
nor U2808 (N_2808,In_1485,In_206);
or U2809 (N_2809,In_1005,In_2412);
nand U2810 (N_2810,In_2297,In_512);
nor U2811 (N_2811,In_1833,In_1486);
nor U2812 (N_2812,In_2395,In_781);
xnor U2813 (N_2813,In_1819,In_2354);
xnor U2814 (N_2814,In_85,In_1755);
xnor U2815 (N_2815,In_18,In_425);
and U2816 (N_2816,In_1139,In_737);
and U2817 (N_2817,In_501,In_989);
or U2818 (N_2818,In_205,In_2299);
nor U2819 (N_2819,In_398,In_115);
and U2820 (N_2820,In_711,In_1171);
nor U2821 (N_2821,In_2153,In_2399);
nor U2822 (N_2822,In_294,In_2096);
or U2823 (N_2823,In_2080,In_1856);
or U2824 (N_2824,In_151,In_1576);
nor U2825 (N_2825,In_994,In_1696);
nand U2826 (N_2826,In_1284,In_1975);
nor U2827 (N_2827,In_1097,In_1066);
nor U2828 (N_2828,In_1346,In_167);
nand U2829 (N_2829,In_1598,In_2465);
nand U2830 (N_2830,In_631,In_486);
or U2831 (N_2831,In_369,In_1355);
and U2832 (N_2832,In_1283,In_2296);
xor U2833 (N_2833,In_9,In_2177);
xnor U2834 (N_2834,In_2172,In_121);
or U2835 (N_2835,In_1914,In_1197);
and U2836 (N_2836,In_106,In_847);
or U2837 (N_2837,In_1370,In_2326);
nand U2838 (N_2838,In_1590,In_2193);
nand U2839 (N_2839,In_1527,In_1320);
and U2840 (N_2840,In_1739,In_1821);
xor U2841 (N_2841,In_462,In_399);
xor U2842 (N_2842,In_786,In_296);
xor U2843 (N_2843,In_2109,In_2227);
xnor U2844 (N_2844,In_1726,In_2363);
and U2845 (N_2845,In_201,In_1743);
xnor U2846 (N_2846,In_773,In_925);
nor U2847 (N_2847,In_5,In_360);
and U2848 (N_2848,In_817,In_457);
nor U2849 (N_2849,In_2465,In_1933);
and U2850 (N_2850,In_2023,In_1044);
or U2851 (N_2851,In_1635,In_1207);
nand U2852 (N_2852,In_248,In_738);
and U2853 (N_2853,In_119,In_1454);
nor U2854 (N_2854,In_1983,In_1794);
or U2855 (N_2855,In_2103,In_2438);
and U2856 (N_2856,In_315,In_1684);
or U2857 (N_2857,In_397,In_1587);
or U2858 (N_2858,In_0,In_1162);
xnor U2859 (N_2859,In_475,In_1995);
or U2860 (N_2860,In_1021,In_499);
or U2861 (N_2861,In_1846,In_1780);
xor U2862 (N_2862,In_1095,In_503);
xor U2863 (N_2863,In_2366,In_2015);
xor U2864 (N_2864,In_1981,In_985);
xor U2865 (N_2865,In_2109,In_1209);
nor U2866 (N_2866,In_1098,In_995);
and U2867 (N_2867,In_485,In_831);
nor U2868 (N_2868,In_10,In_863);
or U2869 (N_2869,In_1685,In_2126);
or U2870 (N_2870,In_727,In_910);
nor U2871 (N_2871,In_1354,In_2000);
and U2872 (N_2872,In_125,In_2360);
xnor U2873 (N_2873,In_338,In_1033);
or U2874 (N_2874,In_938,In_2086);
nor U2875 (N_2875,In_1756,In_543);
and U2876 (N_2876,In_1047,In_1048);
or U2877 (N_2877,In_1821,In_1043);
nand U2878 (N_2878,In_1196,In_925);
and U2879 (N_2879,In_1422,In_1614);
and U2880 (N_2880,In_728,In_2135);
xor U2881 (N_2881,In_2401,In_1130);
nand U2882 (N_2882,In_1078,In_1019);
nor U2883 (N_2883,In_999,In_2451);
nor U2884 (N_2884,In_1298,In_954);
nor U2885 (N_2885,In_305,In_1027);
xor U2886 (N_2886,In_1873,In_1182);
and U2887 (N_2887,In_651,In_363);
nand U2888 (N_2888,In_1192,In_2227);
nand U2889 (N_2889,In_1928,In_257);
nor U2890 (N_2890,In_592,In_1395);
and U2891 (N_2891,In_2167,In_905);
and U2892 (N_2892,In_635,In_139);
and U2893 (N_2893,In_298,In_1896);
and U2894 (N_2894,In_2148,In_2216);
and U2895 (N_2895,In_2217,In_1686);
nand U2896 (N_2896,In_1534,In_1871);
nor U2897 (N_2897,In_1141,In_490);
nand U2898 (N_2898,In_1897,In_662);
nor U2899 (N_2899,In_2308,In_1676);
and U2900 (N_2900,In_1699,In_2121);
and U2901 (N_2901,In_1879,In_2198);
xnor U2902 (N_2902,In_413,In_427);
and U2903 (N_2903,In_938,In_2351);
and U2904 (N_2904,In_1334,In_2294);
xnor U2905 (N_2905,In_342,In_1317);
and U2906 (N_2906,In_1952,In_1407);
xor U2907 (N_2907,In_788,In_2162);
and U2908 (N_2908,In_251,In_1885);
nand U2909 (N_2909,In_42,In_1305);
xor U2910 (N_2910,In_250,In_1044);
or U2911 (N_2911,In_1345,In_2084);
xor U2912 (N_2912,In_2361,In_1194);
and U2913 (N_2913,In_806,In_1784);
xor U2914 (N_2914,In_533,In_1767);
nand U2915 (N_2915,In_362,In_1935);
xor U2916 (N_2916,In_1019,In_1556);
nor U2917 (N_2917,In_1575,In_165);
xor U2918 (N_2918,In_827,In_1695);
nor U2919 (N_2919,In_540,In_939);
xor U2920 (N_2920,In_1773,In_101);
or U2921 (N_2921,In_2481,In_2343);
or U2922 (N_2922,In_1564,In_851);
nand U2923 (N_2923,In_1245,In_477);
xnor U2924 (N_2924,In_1224,In_1128);
nand U2925 (N_2925,In_708,In_84);
xnor U2926 (N_2926,In_336,In_2479);
and U2927 (N_2927,In_1646,In_2461);
xor U2928 (N_2928,In_1694,In_470);
nor U2929 (N_2929,In_2413,In_76);
xor U2930 (N_2930,In_56,In_464);
or U2931 (N_2931,In_2201,In_1871);
and U2932 (N_2932,In_502,In_965);
and U2933 (N_2933,In_490,In_1978);
nand U2934 (N_2934,In_2220,In_1513);
nand U2935 (N_2935,In_2383,In_1727);
nor U2936 (N_2936,In_2080,In_1109);
xnor U2937 (N_2937,In_1602,In_2434);
nand U2938 (N_2938,In_422,In_2171);
xor U2939 (N_2939,In_2469,In_258);
xor U2940 (N_2940,In_1555,In_544);
xor U2941 (N_2941,In_1324,In_1704);
or U2942 (N_2942,In_2043,In_1496);
nand U2943 (N_2943,In_727,In_831);
and U2944 (N_2944,In_427,In_2204);
or U2945 (N_2945,In_2262,In_2289);
or U2946 (N_2946,In_2127,In_512);
xnor U2947 (N_2947,In_1891,In_847);
nand U2948 (N_2948,In_1732,In_776);
and U2949 (N_2949,In_411,In_509);
xor U2950 (N_2950,In_887,In_1376);
nand U2951 (N_2951,In_78,In_1892);
and U2952 (N_2952,In_2318,In_2282);
and U2953 (N_2953,In_426,In_495);
or U2954 (N_2954,In_332,In_851);
and U2955 (N_2955,In_564,In_2244);
or U2956 (N_2956,In_1923,In_1913);
nand U2957 (N_2957,In_1796,In_1269);
nor U2958 (N_2958,In_900,In_1651);
nor U2959 (N_2959,In_681,In_2151);
xnor U2960 (N_2960,In_1630,In_2268);
or U2961 (N_2961,In_387,In_86);
and U2962 (N_2962,In_148,In_1937);
nand U2963 (N_2963,In_210,In_2308);
and U2964 (N_2964,In_176,In_1704);
nand U2965 (N_2965,In_591,In_2424);
and U2966 (N_2966,In_969,In_1211);
and U2967 (N_2967,In_937,In_1824);
or U2968 (N_2968,In_1339,In_608);
or U2969 (N_2969,In_1590,In_2454);
and U2970 (N_2970,In_241,In_359);
nor U2971 (N_2971,In_2428,In_594);
xnor U2972 (N_2972,In_2185,In_576);
nor U2973 (N_2973,In_1152,In_768);
nand U2974 (N_2974,In_1305,In_1892);
nor U2975 (N_2975,In_616,In_1718);
and U2976 (N_2976,In_427,In_1800);
nand U2977 (N_2977,In_862,In_171);
nor U2978 (N_2978,In_390,In_967);
or U2979 (N_2979,In_2311,In_1747);
and U2980 (N_2980,In_385,In_387);
nand U2981 (N_2981,In_1399,In_1011);
and U2982 (N_2982,In_1548,In_1643);
and U2983 (N_2983,In_149,In_1818);
nand U2984 (N_2984,In_1600,In_154);
xor U2985 (N_2985,In_2147,In_1902);
and U2986 (N_2986,In_433,In_1821);
xor U2987 (N_2987,In_1385,In_718);
nand U2988 (N_2988,In_981,In_72);
nand U2989 (N_2989,In_1637,In_81);
or U2990 (N_2990,In_389,In_1971);
and U2991 (N_2991,In_236,In_1256);
nor U2992 (N_2992,In_2065,In_530);
nand U2993 (N_2993,In_1257,In_1456);
or U2994 (N_2994,In_2373,In_2071);
nor U2995 (N_2995,In_1449,In_212);
nand U2996 (N_2996,In_2435,In_1061);
nand U2997 (N_2997,In_963,In_1136);
nor U2998 (N_2998,In_1867,In_827);
nand U2999 (N_2999,In_1411,In_728);
and U3000 (N_3000,In_1962,In_1475);
and U3001 (N_3001,In_2311,In_1187);
and U3002 (N_3002,In_100,In_83);
and U3003 (N_3003,In_970,In_1454);
nand U3004 (N_3004,In_948,In_221);
nand U3005 (N_3005,In_1375,In_961);
and U3006 (N_3006,In_1746,In_344);
or U3007 (N_3007,In_1084,In_987);
or U3008 (N_3008,In_1333,In_1477);
or U3009 (N_3009,In_382,In_1290);
xnor U3010 (N_3010,In_733,In_383);
or U3011 (N_3011,In_589,In_1543);
nor U3012 (N_3012,In_1976,In_2206);
and U3013 (N_3013,In_1401,In_568);
xnor U3014 (N_3014,In_1006,In_2078);
or U3015 (N_3015,In_906,In_2130);
and U3016 (N_3016,In_2411,In_670);
nand U3017 (N_3017,In_795,In_1418);
or U3018 (N_3018,In_904,In_1790);
nor U3019 (N_3019,In_19,In_1210);
and U3020 (N_3020,In_1637,In_138);
nor U3021 (N_3021,In_1352,In_2078);
nor U3022 (N_3022,In_370,In_2385);
nand U3023 (N_3023,In_659,In_623);
xor U3024 (N_3024,In_1931,In_990);
and U3025 (N_3025,In_2195,In_1611);
nor U3026 (N_3026,In_2376,In_2336);
xor U3027 (N_3027,In_1919,In_230);
nor U3028 (N_3028,In_2338,In_913);
nand U3029 (N_3029,In_1084,In_404);
nand U3030 (N_3030,In_905,In_1779);
or U3031 (N_3031,In_1786,In_32);
nand U3032 (N_3032,In_1971,In_383);
and U3033 (N_3033,In_122,In_2070);
xor U3034 (N_3034,In_1342,In_258);
or U3035 (N_3035,In_2350,In_241);
xor U3036 (N_3036,In_1116,In_451);
xnor U3037 (N_3037,In_603,In_482);
or U3038 (N_3038,In_880,In_1437);
or U3039 (N_3039,In_384,In_644);
xnor U3040 (N_3040,In_696,In_1896);
and U3041 (N_3041,In_1506,In_1733);
nand U3042 (N_3042,In_1640,In_241);
nor U3043 (N_3043,In_1497,In_1628);
or U3044 (N_3044,In_485,In_1469);
nor U3045 (N_3045,In_2244,In_548);
nor U3046 (N_3046,In_1577,In_1209);
or U3047 (N_3047,In_1747,In_1670);
nor U3048 (N_3048,In_1492,In_385);
and U3049 (N_3049,In_2248,In_2307);
and U3050 (N_3050,In_2160,In_1879);
nor U3051 (N_3051,In_2420,In_1683);
and U3052 (N_3052,In_1999,In_400);
xnor U3053 (N_3053,In_1680,In_1557);
nor U3054 (N_3054,In_1103,In_819);
or U3055 (N_3055,In_1276,In_1326);
xnor U3056 (N_3056,In_1066,In_965);
or U3057 (N_3057,In_1339,In_1758);
xnor U3058 (N_3058,In_2126,In_1655);
and U3059 (N_3059,In_688,In_2475);
xor U3060 (N_3060,In_2276,In_793);
xnor U3061 (N_3061,In_2037,In_1017);
and U3062 (N_3062,In_1825,In_1569);
or U3063 (N_3063,In_447,In_384);
nand U3064 (N_3064,In_227,In_14);
xnor U3065 (N_3065,In_542,In_342);
nand U3066 (N_3066,In_1788,In_2342);
and U3067 (N_3067,In_704,In_415);
nand U3068 (N_3068,In_639,In_1165);
nor U3069 (N_3069,In_1562,In_2321);
nand U3070 (N_3070,In_1243,In_1747);
nand U3071 (N_3071,In_2368,In_501);
and U3072 (N_3072,In_1297,In_1937);
nor U3073 (N_3073,In_682,In_150);
nand U3074 (N_3074,In_2172,In_1960);
and U3075 (N_3075,In_1567,In_1212);
nor U3076 (N_3076,In_836,In_2463);
nor U3077 (N_3077,In_290,In_1129);
xor U3078 (N_3078,In_2335,In_1977);
xnor U3079 (N_3079,In_252,In_2330);
nand U3080 (N_3080,In_1092,In_905);
nor U3081 (N_3081,In_828,In_1876);
nor U3082 (N_3082,In_102,In_1461);
nor U3083 (N_3083,In_125,In_1453);
xor U3084 (N_3084,In_865,In_2011);
nand U3085 (N_3085,In_1201,In_1830);
and U3086 (N_3086,In_53,In_1216);
and U3087 (N_3087,In_574,In_879);
xor U3088 (N_3088,In_1988,In_2382);
nor U3089 (N_3089,In_676,In_2008);
nor U3090 (N_3090,In_1678,In_2476);
nor U3091 (N_3091,In_133,In_452);
and U3092 (N_3092,In_2045,In_2059);
nor U3093 (N_3093,In_1756,In_974);
nand U3094 (N_3094,In_1782,In_1674);
nand U3095 (N_3095,In_1364,In_377);
and U3096 (N_3096,In_2130,In_2303);
nand U3097 (N_3097,In_1639,In_2352);
or U3098 (N_3098,In_1400,In_956);
and U3099 (N_3099,In_877,In_1173);
nor U3100 (N_3100,In_1159,In_314);
nor U3101 (N_3101,In_2119,In_2169);
and U3102 (N_3102,In_357,In_1264);
nand U3103 (N_3103,In_160,In_2045);
nand U3104 (N_3104,In_1696,In_798);
and U3105 (N_3105,In_2231,In_907);
or U3106 (N_3106,In_640,In_1875);
nor U3107 (N_3107,In_538,In_352);
xor U3108 (N_3108,In_944,In_2055);
or U3109 (N_3109,In_2067,In_110);
nor U3110 (N_3110,In_2227,In_39);
or U3111 (N_3111,In_2391,In_704);
or U3112 (N_3112,In_867,In_1806);
and U3113 (N_3113,In_1257,In_1721);
nand U3114 (N_3114,In_429,In_466);
or U3115 (N_3115,In_1624,In_236);
or U3116 (N_3116,In_810,In_1731);
nor U3117 (N_3117,In_1600,In_1749);
nor U3118 (N_3118,In_1229,In_1517);
and U3119 (N_3119,In_1455,In_2441);
and U3120 (N_3120,In_880,In_1694);
nand U3121 (N_3121,In_1294,In_2480);
and U3122 (N_3122,In_2474,In_1011);
nand U3123 (N_3123,In_2485,In_488);
nor U3124 (N_3124,In_1021,In_458);
and U3125 (N_3125,In_645,In_642);
and U3126 (N_3126,In_656,In_2228);
nor U3127 (N_3127,In_2239,In_1937);
nand U3128 (N_3128,In_655,In_313);
xor U3129 (N_3129,In_330,In_795);
or U3130 (N_3130,In_981,In_1686);
nand U3131 (N_3131,In_2208,In_2105);
nor U3132 (N_3132,In_1678,In_1854);
xnor U3133 (N_3133,In_346,In_975);
or U3134 (N_3134,In_64,In_906);
xnor U3135 (N_3135,In_482,In_245);
and U3136 (N_3136,In_864,In_322);
nor U3137 (N_3137,In_24,In_1108);
and U3138 (N_3138,In_2174,In_94);
xor U3139 (N_3139,In_2467,In_323);
or U3140 (N_3140,In_664,In_1979);
xor U3141 (N_3141,In_1013,In_337);
or U3142 (N_3142,In_2317,In_1961);
and U3143 (N_3143,In_792,In_644);
nand U3144 (N_3144,In_1207,In_1281);
nand U3145 (N_3145,In_649,In_1872);
xor U3146 (N_3146,In_1425,In_1756);
or U3147 (N_3147,In_1282,In_1495);
nor U3148 (N_3148,In_2399,In_566);
or U3149 (N_3149,In_732,In_2045);
nor U3150 (N_3150,In_1155,In_1542);
or U3151 (N_3151,In_534,In_198);
or U3152 (N_3152,In_1902,In_1167);
nand U3153 (N_3153,In_857,In_1138);
xor U3154 (N_3154,In_1986,In_771);
nand U3155 (N_3155,In_1018,In_949);
nand U3156 (N_3156,In_772,In_2426);
xor U3157 (N_3157,In_283,In_16);
nand U3158 (N_3158,In_1679,In_2168);
xnor U3159 (N_3159,In_718,In_1804);
and U3160 (N_3160,In_1038,In_326);
nor U3161 (N_3161,In_337,In_1898);
xnor U3162 (N_3162,In_1796,In_1551);
and U3163 (N_3163,In_947,In_1955);
nor U3164 (N_3164,In_1333,In_683);
or U3165 (N_3165,In_1423,In_2151);
xor U3166 (N_3166,In_1821,In_2357);
xnor U3167 (N_3167,In_2257,In_2327);
xnor U3168 (N_3168,In_264,In_2122);
nand U3169 (N_3169,In_279,In_1421);
and U3170 (N_3170,In_2239,In_1730);
nor U3171 (N_3171,In_1760,In_1539);
nand U3172 (N_3172,In_2126,In_1473);
nand U3173 (N_3173,In_1412,In_581);
nor U3174 (N_3174,In_2246,In_744);
nor U3175 (N_3175,In_1474,In_1478);
nand U3176 (N_3176,In_2182,In_155);
or U3177 (N_3177,In_2196,In_2018);
nand U3178 (N_3178,In_580,In_360);
nor U3179 (N_3179,In_2301,In_275);
and U3180 (N_3180,In_1056,In_641);
and U3181 (N_3181,In_1184,In_203);
xnor U3182 (N_3182,In_2165,In_1482);
nand U3183 (N_3183,In_237,In_151);
xor U3184 (N_3184,In_2165,In_1136);
or U3185 (N_3185,In_1289,In_1458);
nor U3186 (N_3186,In_1579,In_875);
or U3187 (N_3187,In_774,In_752);
nor U3188 (N_3188,In_424,In_2211);
xor U3189 (N_3189,In_676,In_1290);
and U3190 (N_3190,In_1270,In_1944);
or U3191 (N_3191,In_1691,In_278);
xnor U3192 (N_3192,In_1735,In_1128);
xor U3193 (N_3193,In_2379,In_1172);
xor U3194 (N_3194,In_1853,In_265);
xnor U3195 (N_3195,In_1098,In_2154);
nand U3196 (N_3196,In_1635,In_1448);
or U3197 (N_3197,In_897,In_1104);
nor U3198 (N_3198,In_338,In_1115);
nand U3199 (N_3199,In_882,In_1357);
nand U3200 (N_3200,In_23,In_637);
xor U3201 (N_3201,In_994,In_1028);
nor U3202 (N_3202,In_1164,In_1066);
or U3203 (N_3203,In_1200,In_1214);
or U3204 (N_3204,In_85,In_1560);
and U3205 (N_3205,In_1786,In_369);
and U3206 (N_3206,In_426,In_2032);
and U3207 (N_3207,In_76,In_2280);
or U3208 (N_3208,In_879,In_2214);
nand U3209 (N_3209,In_23,In_683);
or U3210 (N_3210,In_793,In_124);
and U3211 (N_3211,In_1482,In_649);
xor U3212 (N_3212,In_1277,In_8);
or U3213 (N_3213,In_1384,In_2203);
xor U3214 (N_3214,In_464,In_1169);
nand U3215 (N_3215,In_1994,In_1176);
or U3216 (N_3216,In_830,In_1830);
nor U3217 (N_3217,In_1836,In_1626);
xnor U3218 (N_3218,In_1297,In_781);
nand U3219 (N_3219,In_2251,In_1049);
nor U3220 (N_3220,In_16,In_1809);
nor U3221 (N_3221,In_1489,In_1773);
nand U3222 (N_3222,In_1194,In_757);
xor U3223 (N_3223,In_1954,In_825);
nor U3224 (N_3224,In_1961,In_2167);
nor U3225 (N_3225,In_1809,In_1950);
nand U3226 (N_3226,In_1199,In_1808);
xnor U3227 (N_3227,In_2143,In_1906);
or U3228 (N_3228,In_2394,In_1775);
or U3229 (N_3229,In_1688,In_1985);
or U3230 (N_3230,In_1223,In_1256);
or U3231 (N_3231,In_994,In_2129);
xor U3232 (N_3232,In_2022,In_2203);
nand U3233 (N_3233,In_277,In_1927);
nor U3234 (N_3234,In_1162,In_1499);
nand U3235 (N_3235,In_629,In_1158);
and U3236 (N_3236,In_2148,In_825);
xor U3237 (N_3237,In_2265,In_1513);
xor U3238 (N_3238,In_1005,In_1644);
nor U3239 (N_3239,In_1131,In_812);
and U3240 (N_3240,In_2434,In_1519);
nand U3241 (N_3241,In_325,In_2268);
or U3242 (N_3242,In_645,In_2439);
nor U3243 (N_3243,In_180,In_403);
xor U3244 (N_3244,In_1979,In_2302);
xor U3245 (N_3245,In_1813,In_180);
or U3246 (N_3246,In_1831,In_1815);
and U3247 (N_3247,In_392,In_1369);
nand U3248 (N_3248,In_1780,In_23);
nand U3249 (N_3249,In_1312,In_2296);
xor U3250 (N_3250,In_1676,In_553);
nand U3251 (N_3251,In_557,In_142);
and U3252 (N_3252,In_1050,In_507);
nand U3253 (N_3253,In_1240,In_2085);
or U3254 (N_3254,In_1234,In_2315);
nand U3255 (N_3255,In_566,In_75);
nor U3256 (N_3256,In_1387,In_879);
nand U3257 (N_3257,In_674,In_1036);
nand U3258 (N_3258,In_371,In_1935);
nand U3259 (N_3259,In_1716,In_1386);
or U3260 (N_3260,In_405,In_2450);
nor U3261 (N_3261,In_1877,In_2471);
xor U3262 (N_3262,In_739,In_165);
and U3263 (N_3263,In_107,In_1182);
nor U3264 (N_3264,In_1620,In_1263);
and U3265 (N_3265,In_2368,In_1205);
and U3266 (N_3266,In_2278,In_1482);
or U3267 (N_3267,In_2394,In_735);
nor U3268 (N_3268,In_1548,In_532);
xor U3269 (N_3269,In_1400,In_191);
and U3270 (N_3270,In_419,In_762);
and U3271 (N_3271,In_753,In_2084);
nor U3272 (N_3272,In_1166,In_1542);
nand U3273 (N_3273,In_2236,In_1339);
nand U3274 (N_3274,In_225,In_113);
nand U3275 (N_3275,In_753,In_2070);
and U3276 (N_3276,In_1624,In_1527);
or U3277 (N_3277,In_192,In_1167);
nand U3278 (N_3278,In_2186,In_1404);
xnor U3279 (N_3279,In_449,In_1322);
xnor U3280 (N_3280,In_2055,In_2008);
xor U3281 (N_3281,In_431,In_281);
nand U3282 (N_3282,In_1925,In_406);
or U3283 (N_3283,In_73,In_699);
nor U3284 (N_3284,In_415,In_760);
nand U3285 (N_3285,In_921,In_1891);
nand U3286 (N_3286,In_410,In_1438);
nand U3287 (N_3287,In_1242,In_1232);
xnor U3288 (N_3288,In_1003,In_2062);
nor U3289 (N_3289,In_2338,In_2121);
nor U3290 (N_3290,In_1495,In_476);
or U3291 (N_3291,In_1802,In_1548);
and U3292 (N_3292,In_2138,In_1295);
nor U3293 (N_3293,In_1383,In_2445);
nand U3294 (N_3294,In_1818,In_1319);
and U3295 (N_3295,In_1483,In_1347);
or U3296 (N_3296,In_287,In_2282);
xor U3297 (N_3297,In_1543,In_972);
nand U3298 (N_3298,In_1619,In_1683);
nor U3299 (N_3299,In_1115,In_644);
or U3300 (N_3300,In_27,In_1015);
xor U3301 (N_3301,In_2353,In_1676);
xor U3302 (N_3302,In_2031,In_2000);
nor U3303 (N_3303,In_1052,In_2126);
nand U3304 (N_3304,In_1693,In_81);
nand U3305 (N_3305,In_30,In_1959);
xnor U3306 (N_3306,In_2166,In_2404);
or U3307 (N_3307,In_433,In_1701);
nand U3308 (N_3308,In_99,In_2004);
nor U3309 (N_3309,In_1838,In_245);
nor U3310 (N_3310,In_2233,In_2478);
nand U3311 (N_3311,In_1196,In_1278);
and U3312 (N_3312,In_1142,In_1060);
nand U3313 (N_3313,In_2087,In_84);
and U3314 (N_3314,In_1801,In_1912);
and U3315 (N_3315,In_916,In_2162);
xnor U3316 (N_3316,In_2146,In_101);
nor U3317 (N_3317,In_306,In_1769);
nand U3318 (N_3318,In_1242,In_2459);
nand U3319 (N_3319,In_1060,In_922);
or U3320 (N_3320,In_433,In_2188);
xor U3321 (N_3321,In_989,In_2021);
nor U3322 (N_3322,In_1163,In_1415);
nor U3323 (N_3323,In_1551,In_389);
nand U3324 (N_3324,In_2433,In_1154);
and U3325 (N_3325,In_994,In_257);
nor U3326 (N_3326,In_48,In_1082);
or U3327 (N_3327,In_840,In_1107);
nor U3328 (N_3328,In_1882,In_16);
nand U3329 (N_3329,In_1497,In_259);
or U3330 (N_3330,In_831,In_1841);
nand U3331 (N_3331,In_1158,In_1930);
xor U3332 (N_3332,In_509,In_808);
and U3333 (N_3333,In_1048,In_2102);
or U3334 (N_3334,In_523,In_771);
and U3335 (N_3335,In_1917,In_2472);
or U3336 (N_3336,In_593,In_2081);
nor U3337 (N_3337,In_1261,In_2366);
and U3338 (N_3338,In_1911,In_664);
and U3339 (N_3339,In_202,In_1280);
xor U3340 (N_3340,In_962,In_765);
or U3341 (N_3341,In_1042,In_1226);
nor U3342 (N_3342,In_1127,In_978);
and U3343 (N_3343,In_2081,In_1537);
nor U3344 (N_3344,In_1747,In_947);
xor U3345 (N_3345,In_1376,In_1804);
nor U3346 (N_3346,In_2070,In_2315);
or U3347 (N_3347,In_1145,In_1252);
xor U3348 (N_3348,In_1860,In_2349);
or U3349 (N_3349,In_900,In_1526);
and U3350 (N_3350,In_932,In_945);
or U3351 (N_3351,In_638,In_1495);
or U3352 (N_3352,In_1633,In_857);
and U3353 (N_3353,In_2116,In_702);
nand U3354 (N_3354,In_196,In_1766);
or U3355 (N_3355,In_2042,In_315);
nor U3356 (N_3356,In_2227,In_1661);
nor U3357 (N_3357,In_2387,In_271);
nor U3358 (N_3358,In_1417,In_1952);
or U3359 (N_3359,In_2087,In_1572);
xor U3360 (N_3360,In_801,In_379);
xor U3361 (N_3361,In_14,In_176);
or U3362 (N_3362,In_1193,In_338);
and U3363 (N_3363,In_2470,In_1383);
nor U3364 (N_3364,In_835,In_990);
nand U3365 (N_3365,In_771,In_219);
or U3366 (N_3366,In_825,In_2414);
nand U3367 (N_3367,In_2079,In_2342);
and U3368 (N_3368,In_816,In_1421);
nor U3369 (N_3369,In_984,In_531);
or U3370 (N_3370,In_2362,In_224);
and U3371 (N_3371,In_1909,In_824);
or U3372 (N_3372,In_1838,In_1286);
xor U3373 (N_3373,In_579,In_2390);
nor U3374 (N_3374,In_534,In_1535);
and U3375 (N_3375,In_1812,In_839);
nor U3376 (N_3376,In_2159,In_162);
nand U3377 (N_3377,In_1950,In_494);
xor U3378 (N_3378,In_1310,In_1182);
and U3379 (N_3379,In_659,In_1889);
nand U3380 (N_3380,In_2414,In_1216);
xor U3381 (N_3381,In_1067,In_17);
and U3382 (N_3382,In_1192,In_1816);
or U3383 (N_3383,In_1356,In_144);
and U3384 (N_3384,In_8,In_529);
or U3385 (N_3385,In_1996,In_785);
nor U3386 (N_3386,In_306,In_1731);
nand U3387 (N_3387,In_1643,In_746);
or U3388 (N_3388,In_2429,In_346);
xnor U3389 (N_3389,In_506,In_1957);
nor U3390 (N_3390,In_772,In_672);
and U3391 (N_3391,In_349,In_2166);
and U3392 (N_3392,In_1177,In_25);
nor U3393 (N_3393,In_1088,In_1166);
or U3394 (N_3394,In_1134,In_52);
and U3395 (N_3395,In_1464,In_1166);
xnor U3396 (N_3396,In_895,In_2105);
or U3397 (N_3397,In_967,In_1881);
xor U3398 (N_3398,In_2461,In_2006);
or U3399 (N_3399,In_1283,In_1233);
xnor U3400 (N_3400,In_2135,In_75);
and U3401 (N_3401,In_1099,In_63);
nor U3402 (N_3402,In_2116,In_602);
xor U3403 (N_3403,In_1784,In_2086);
nand U3404 (N_3404,In_2029,In_2080);
xnor U3405 (N_3405,In_2223,In_799);
and U3406 (N_3406,In_272,In_1401);
xor U3407 (N_3407,In_294,In_2117);
xor U3408 (N_3408,In_2421,In_537);
nor U3409 (N_3409,In_2400,In_1140);
nor U3410 (N_3410,In_201,In_96);
xor U3411 (N_3411,In_372,In_2136);
nand U3412 (N_3412,In_409,In_2339);
nand U3413 (N_3413,In_1050,In_1919);
or U3414 (N_3414,In_1931,In_1410);
and U3415 (N_3415,In_2009,In_36);
nand U3416 (N_3416,In_526,In_252);
and U3417 (N_3417,In_2407,In_1430);
nand U3418 (N_3418,In_1368,In_881);
nand U3419 (N_3419,In_694,In_1878);
nor U3420 (N_3420,In_547,In_641);
nor U3421 (N_3421,In_1128,In_257);
nand U3422 (N_3422,In_1579,In_2006);
nand U3423 (N_3423,In_1195,In_2470);
or U3424 (N_3424,In_1103,In_1228);
or U3425 (N_3425,In_1880,In_2120);
nand U3426 (N_3426,In_417,In_1104);
and U3427 (N_3427,In_843,In_2392);
xor U3428 (N_3428,In_2451,In_2075);
xor U3429 (N_3429,In_1299,In_1809);
nand U3430 (N_3430,In_1935,In_2239);
nand U3431 (N_3431,In_1545,In_755);
or U3432 (N_3432,In_357,In_1726);
xnor U3433 (N_3433,In_893,In_831);
nand U3434 (N_3434,In_1120,In_1949);
nand U3435 (N_3435,In_1694,In_2100);
nand U3436 (N_3436,In_1503,In_2341);
and U3437 (N_3437,In_635,In_2391);
nor U3438 (N_3438,In_360,In_2034);
xor U3439 (N_3439,In_392,In_1816);
or U3440 (N_3440,In_790,In_1351);
xnor U3441 (N_3441,In_2240,In_1953);
nor U3442 (N_3442,In_484,In_1052);
and U3443 (N_3443,In_1331,In_2138);
and U3444 (N_3444,In_1205,In_370);
and U3445 (N_3445,In_2101,In_2244);
or U3446 (N_3446,In_278,In_1015);
and U3447 (N_3447,In_1350,In_2090);
nand U3448 (N_3448,In_2470,In_1334);
or U3449 (N_3449,In_2447,In_1280);
nand U3450 (N_3450,In_1092,In_1831);
nor U3451 (N_3451,In_2038,In_1045);
nand U3452 (N_3452,In_792,In_917);
nand U3453 (N_3453,In_2046,In_920);
nand U3454 (N_3454,In_2453,In_740);
nor U3455 (N_3455,In_548,In_1454);
and U3456 (N_3456,In_2012,In_1606);
nor U3457 (N_3457,In_246,In_925);
or U3458 (N_3458,In_245,In_1916);
and U3459 (N_3459,In_1101,In_2007);
nor U3460 (N_3460,In_63,In_150);
nor U3461 (N_3461,In_2266,In_1299);
xor U3462 (N_3462,In_1798,In_1994);
and U3463 (N_3463,In_997,In_1106);
nor U3464 (N_3464,In_666,In_1188);
or U3465 (N_3465,In_2466,In_2389);
nor U3466 (N_3466,In_347,In_1570);
xor U3467 (N_3467,In_1856,In_34);
and U3468 (N_3468,In_910,In_1562);
and U3469 (N_3469,In_1868,In_824);
and U3470 (N_3470,In_1800,In_377);
and U3471 (N_3471,In_1505,In_639);
xnor U3472 (N_3472,In_1759,In_1274);
or U3473 (N_3473,In_414,In_1388);
xnor U3474 (N_3474,In_721,In_760);
or U3475 (N_3475,In_212,In_2070);
nand U3476 (N_3476,In_1745,In_417);
nor U3477 (N_3477,In_134,In_1523);
and U3478 (N_3478,In_136,In_559);
and U3479 (N_3479,In_1747,In_713);
or U3480 (N_3480,In_1478,In_36);
xor U3481 (N_3481,In_1638,In_1907);
nand U3482 (N_3482,In_605,In_1358);
nand U3483 (N_3483,In_662,In_1174);
xnor U3484 (N_3484,In_2059,In_1092);
or U3485 (N_3485,In_2357,In_2401);
nand U3486 (N_3486,In_1484,In_1383);
nand U3487 (N_3487,In_1573,In_888);
nor U3488 (N_3488,In_253,In_381);
or U3489 (N_3489,In_329,In_1874);
or U3490 (N_3490,In_1101,In_2425);
xor U3491 (N_3491,In_2376,In_1090);
or U3492 (N_3492,In_919,In_490);
or U3493 (N_3493,In_193,In_970);
or U3494 (N_3494,In_362,In_2104);
nor U3495 (N_3495,In_268,In_82);
or U3496 (N_3496,In_326,In_1164);
or U3497 (N_3497,In_1507,In_668);
nor U3498 (N_3498,In_1211,In_1092);
or U3499 (N_3499,In_250,In_1223);
or U3500 (N_3500,In_796,In_777);
nand U3501 (N_3501,In_1783,In_2442);
nand U3502 (N_3502,In_235,In_2127);
and U3503 (N_3503,In_494,In_1130);
nand U3504 (N_3504,In_2303,In_310);
xnor U3505 (N_3505,In_1638,In_397);
nand U3506 (N_3506,In_1023,In_1912);
or U3507 (N_3507,In_1913,In_656);
and U3508 (N_3508,In_1085,In_970);
or U3509 (N_3509,In_2002,In_1806);
nor U3510 (N_3510,In_356,In_1490);
nor U3511 (N_3511,In_1769,In_1803);
or U3512 (N_3512,In_176,In_1776);
and U3513 (N_3513,In_1692,In_724);
nand U3514 (N_3514,In_1658,In_2008);
xor U3515 (N_3515,In_1150,In_2487);
nand U3516 (N_3516,In_882,In_768);
and U3517 (N_3517,In_329,In_318);
nor U3518 (N_3518,In_1110,In_2327);
nor U3519 (N_3519,In_1931,In_2148);
nor U3520 (N_3520,In_458,In_936);
xnor U3521 (N_3521,In_633,In_811);
and U3522 (N_3522,In_475,In_2109);
xnor U3523 (N_3523,In_1668,In_736);
xnor U3524 (N_3524,In_867,In_141);
or U3525 (N_3525,In_1392,In_2250);
xor U3526 (N_3526,In_398,In_389);
or U3527 (N_3527,In_1271,In_997);
nor U3528 (N_3528,In_677,In_1912);
nand U3529 (N_3529,In_2113,In_1554);
or U3530 (N_3530,In_1423,In_601);
and U3531 (N_3531,In_1312,In_1614);
or U3532 (N_3532,In_1039,In_270);
or U3533 (N_3533,In_673,In_404);
and U3534 (N_3534,In_1820,In_783);
xor U3535 (N_3535,In_1843,In_1710);
nor U3536 (N_3536,In_1284,In_1918);
nor U3537 (N_3537,In_2123,In_647);
or U3538 (N_3538,In_618,In_2233);
xor U3539 (N_3539,In_1093,In_787);
and U3540 (N_3540,In_2266,In_1502);
xor U3541 (N_3541,In_1964,In_688);
xor U3542 (N_3542,In_1699,In_1777);
xnor U3543 (N_3543,In_2042,In_1901);
or U3544 (N_3544,In_1153,In_1478);
or U3545 (N_3545,In_2113,In_766);
xor U3546 (N_3546,In_1725,In_843);
and U3547 (N_3547,In_628,In_891);
and U3548 (N_3548,In_489,In_375);
nor U3549 (N_3549,In_91,In_1407);
and U3550 (N_3550,In_606,In_1670);
nand U3551 (N_3551,In_59,In_1175);
or U3552 (N_3552,In_414,In_1597);
and U3553 (N_3553,In_561,In_1774);
and U3554 (N_3554,In_2444,In_1004);
nand U3555 (N_3555,In_1312,In_2326);
nand U3556 (N_3556,In_1856,In_64);
nand U3557 (N_3557,In_2200,In_1996);
nor U3558 (N_3558,In_1299,In_1357);
nor U3559 (N_3559,In_2308,In_1371);
nor U3560 (N_3560,In_2321,In_1667);
or U3561 (N_3561,In_1027,In_948);
nand U3562 (N_3562,In_1300,In_914);
xnor U3563 (N_3563,In_915,In_309);
nand U3564 (N_3564,In_1104,In_1625);
or U3565 (N_3565,In_411,In_1331);
and U3566 (N_3566,In_2193,In_506);
xor U3567 (N_3567,In_1012,In_2258);
xnor U3568 (N_3568,In_2339,In_2403);
nand U3569 (N_3569,In_1384,In_809);
or U3570 (N_3570,In_337,In_2079);
nor U3571 (N_3571,In_1694,In_1013);
nand U3572 (N_3572,In_773,In_2047);
or U3573 (N_3573,In_1072,In_962);
and U3574 (N_3574,In_175,In_2311);
and U3575 (N_3575,In_1886,In_313);
or U3576 (N_3576,In_848,In_262);
and U3577 (N_3577,In_1138,In_2278);
nand U3578 (N_3578,In_2208,In_2457);
nor U3579 (N_3579,In_274,In_1774);
and U3580 (N_3580,In_687,In_2077);
or U3581 (N_3581,In_963,In_1445);
nor U3582 (N_3582,In_1822,In_980);
nor U3583 (N_3583,In_1360,In_1346);
xnor U3584 (N_3584,In_1951,In_2444);
xnor U3585 (N_3585,In_1957,In_357);
xor U3586 (N_3586,In_2140,In_2053);
and U3587 (N_3587,In_1177,In_1978);
and U3588 (N_3588,In_101,In_529);
xnor U3589 (N_3589,In_5,In_2248);
nor U3590 (N_3590,In_1904,In_612);
nand U3591 (N_3591,In_1852,In_566);
xor U3592 (N_3592,In_746,In_1821);
nor U3593 (N_3593,In_574,In_1740);
or U3594 (N_3594,In_645,In_858);
nand U3595 (N_3595,In_1293,In_987);
nand U3596 (N_3596,In_2070,In_2403);
nor U3597 (N_3597,In_1214,In_2026);
nand U3598 (N_3598,In_361,In_1804);
or U3599 (N_3599,In_325,In_719);
nor U3600 (N_3600,In_2493,In_2342);
or U3601 (N_3601,In_1828,In_240);
and U3602 (N_3602,In_58,In_2427);
nor U3603 (N_3603,In_2134,In_541);
and U3604 (N_3604,In_133,In_166);
nand U3605 (N_3605,In_1067,In_1665);
nand U3606 (N_3606,In_1246,In_2238);
xnor U3607 (N_3607,In_1955,In_1487);
and U3608 (N_3608,In_829,In_483);
or U3609 (N_3609,In_1560,In_1190);
or U3610 (N_3610,In_813,In_213);
or U3611 (N_3611,In_698,In_1730);
nor U3612 (N_3612,In_2438,In_1604);
and U3613 (N_3613,In_2354,In_276);
nor U3614 (N_3614,In_3,In_1033);
nor U3615 (N_3615,In_1457,In_1487);
or U3616 (N_3616,In_638,In_1298);
xor U3617 (N_3617,In_1860,In_2269);
or U3618 (N_3618,In_1328,In_1363);
xor U3619 (N_3619,In_174,In_163);
nor U3620 (N_3620,In_749,In_1338);
nand U3621 (N_3621,In_771,In_447);
or U3622 (N_3622,In_1908,In_1662);
nand U3623 (N_3623,In_1885,In_819);
nor U3624 (N_3624,In_1844,In_1876);
nor U3625 (N_3625,In_1654,In_2141);
nor U3626 (N_3626,In_2465,In_846);
or U3627 (N_3627,In_1360,In_901);
nand U3628 (N_3628,In_1981,In_650);
nand U3629 (N_3629,In_1868,In_404);
xor U3630 (N_3630,In_1872,In_761);
xor U3631 (N_3631,In_1236,In_1369);
xor U3632 (N_3632,In_1487,In_1574);
xor U3633 (N_3633,In_1483,In_491);
and U3634 (N_3634,In_346,In_1049);
nand U3635 (N_3635,In_1030,In_2303);
or U3636 (N_3636,In_1801,In_553);
nand U3637 (N_3637,In_117,In_1237);
nor U3638 (N_3638,In_2327,In_14);
and U3639 (N_3639,In_2439,In_539);
or U3640 (N_3640,In_2430,In_979);
or U3641 (N_3641,In_1868,In_1975);
nand U3642 (N_3642,In_902,In_1089);
nand U3643 (N_3643,In_322,In_250);
nor U3644 (N_3644,In_1919,In_2444);
and U3645 (N_3645,In_36,In_2213);
and U3646 (N_3646,In_63,In_1461);
or U3647 (N_3647,In_2405,In_1728);
or U3648 (N_3648,In_759,In_2112);
and U3649 (N_3649,In_1833,In_2294);
and U3650 (N_3650,In_759,In_385);
nor U3651 (N_3651,In_1151,In_2175);
or U3652 (N_3652,In_92,In_1806);
or U3653 (N_3653,In_991,In_2061);
and U3654 (N_3654,In_384,In_1664);
nor U3655 (N_3655,In_1292,In_2173);
xor U3656 (N_3656,In_1382,In_1588);
and U3657 (N_3657,In_2344,In_2498);
xnor U3658 (N_3658,In_2003,In_994);
and U3659 (N_3659,In_2403,In_1548);
and U3660 (N_3660,In_1617,In_1278);
nor U3661 (N_3661,In_193,In_304);
xnor U3662 (N_3662,In_745,In_628);
or U3663 (N_3663,In_442,In_683);
nand U3664 (N_3664,In_409,In_983);
nor U3665 (N_3665,In_1971,In_1306);
and U3666 (N_3666,In_2154,In_1220);
nor U3667 (N_3667,In_627,In_490);
xor U3668 (N_3668,In_1848,In_124);
xor U3669 (N_3669,In_1674,In_2456);
nand U3670 (N_3670,In_298,In_1981);
xor U3671 (N_3671,In_1622,In_2054);
or U3672 (N_3672,In_858,In_1104);
nor U3673 (N_3673,In_2177,In_242);
nand U3674 (N_3674,In_148,In_1537);
and U3675 (N_3675,In_1032,In_542);
or U3676 (N_3676,In_99,In_821);
nor U3677 (N_3677,In_2320,In_1275);
xor U3678 (N_3678,In_1407,In_108);
and U3679 (N_3679,In_2013,In_1072);
and U3680 (N_3680,In_2413,In_2119);
nor U3681 (N_3681,In_1482,In_1494);
or U3682 (N_3682,In_982,In_2209);
and U3683 (N_3683,In_741,In_959);
nand U3684 (N_3684,In_512,In_1082);
and U3685 (N_3685,In_2119,In_272);
xor U3686 (N_3686,In_396,In_412);
nand U3687 (N_3687,In_134,In_2014);
nor U3688 (N_3688,In_2434,In_1293);
nor U3689 (N_3689,In_1010,In_68);
or U3690 (N_3690,In_592,In_1090);
or U3691 (N_3691,In_1748,In_2076);
or U3692 (N_3692,In_2417,In_239);
or U3693 (N_3693,In_449,In_1402);
and U3694 (N_3694,In_1496,In_953);
nand U3695 (N_3695,In_1908,In_1104);
or U3696 (N_3696,In_1571,In_6);
nor U3697 (N_3697,In_2199,In_2472);
nand U3698 (N_3698,In_545,In_1427);
nand U3699 (N_3699,In_2459,In_683);
and U3700 (N_3700,In_1896,In_2132);
and U3701 (N_3701,In_1500,In_550);
nand U3702 (N_3702,In_1074,In_1688);
and U3703 (N_3703,In_1713,In_358);
and U3704 (N_3704,In_1915,In_1822);
or U3705 (N_3705,In_1756,In_1104);
nand U3706 (N_3706,In_1918,In_1794);
or U3707 (N_3707,In_460,In_1986);
xnor U3708 (N_3708,In_1053,In_2364);
and U3709 (N_3709,In_1998,In_441);
and U3710 (N_3710,In_311,In_965);
and U3711 (N_3711,In_117,In_1952);
nand U3712 (N_3712,In_1150,In_1699);
xor U3713 (N_3713,In_166,In_982);
nand U3714 (N_3714,In_2274,In_648);
xnor U3715 (N_3715,In_2017,In_523);
nand U3716 (N_3716,In_163,In_261);
nand U3717 (N_3717,In_159,In_1829);
xnor U3718 (N_3718,In_302,In_1269);
and U3719 (N_3719,In_2135,In_2115);
and U3720 (N_3720,In_1608,In_1567);
xnor U3721 (N_3721,In_1097,In_785);
nor U3722 (N_3722,In_2462,In_203);
or U3723 (N_3723,In_1113,In_634);
xnor U3724 (N_3724,In_1388,In_1651);
nand U3725 (N_3725,In_2069,In_626);
nand U3726 (N_3726,In_275,In_945);
nand U3727 (N_3727,In_2416,In_647);
or U3728 (N_3728,In_1854,In_1944);
nor U3729 (N_3729,In_1311,In_2335);
or U3730 (N_3730,In_649,In_1791);
or U3731 (N_3731,In_721,In_757);
nand U3732 (N_3732,In_1640,In_1666);
and U3733 (N_3733,In_1030,In_88);
xor U3734 (N_3734,In_1355,In_1783);
and U3735 (N_3735,In_1700,In_836);
or U3736 (N_3736,In_1921,In_336);
or U3737 (N_3737,In_2429,In_253);
xor U3738 (N_3738,In_2370,In_1214);
or U3739 (N_3739,In_1598,In_1587);
xnor U3740 (N_3740,In_1980,In_915);
nand U3741 (N_3741,In_87,In_1721);
nand U3742 (N_3742,In_909,In_1263);
or U3743 (N_3743,In_439,In_2140);
and U3744 (N_3744,In_1249,In_1547);
nor U3745 (N_3745,In_1703,In_1714);
xnor U3746 (N_3746,In_195,In_1232);
and U3747 (N_3747,In_1340,In_1078);
nor U3748 (N_3748,In_776,In_215);
nand U3749 (N_3749,In_219,In_2007);
and U3750 (N_3750,In_2066,In_2104);
or U3751 (N_3751,In_1639,In_308);
nand U3752 (N_3752,In_1151,In_195);
or U3753 (N_3753,In_1942,In_318);
xnor U3754 (N_3754,In_1940,In_1925);
xnor U3755 (N_3755,In_1586,In_1168);
nor U3756 (N_3756,In_1403,In_897);
nand U3757 (N_3757,In_1372,In_2390);
nor U3758 (N_3758,In_343,In_280);
or U3759 (N_3759,In_2010,In_1915);
nand U3760 (N_3760,In_707,In_1799);
xor U3761 (N_3761,In_573,In_1728);
nand U3762 (N_3762,In_663,In_1879);
nand U3763 (N_3763,In_846,In_981);
or U3764 (N_3764,In_141,In_601);
or U3765 (N_3765,In_1700,In_1997);
and U3766 (N_3766,In_1708,In_664);
and U3767 (N_3767,In_1894,In_2489);
xnor U3768 (N_3768,In_101,In_2448);
or U3769 (N_3769,In_1621,In_888);
or U3770 (N_3770,In_1204,In_2440);
nor U3771 (N_3771,In_1286,In_339);
or U3772 (N_3772,In_1597,In_148);
xnor U3773 (N_3773,In_2440,In_2466);
xnor U3774 (N_3774,In_1543,In_1222);
or U3775 (N_3775,In_550,In_327);
xor U3776 (N_3776,In_540,In_1403);
xor U3777 (N_3777,In_646,In_1765);
xnor U3778 (N_3778,In_1936,In_1033);
nor U3779 (N_3779,In_1246,In_580);
and U3780 (N_3780,In_1190,In_1588);
and U3781 (N_3781,In_182,In_945);
xor U3782 (N_3782,In_1812,In_2279);
or U3783 (N_3783,In_747,In_1249);
or U3784 (N_3784,In_663,In_1128);
xnor U3785 (N_3785,In_1463,In_219);
and U3786 (N_3786,In_1970,In_2029);
nor U3787 (N_3787,In_32,In_1963);
or U3788 (N_3788,In_2046,In_2087);
and U3789 (N_3789,In_274,In_1864);
nand U3790 (N_3790,In_1572,In_491);
xor U3791 (N_3791,In_2179,In_1437);
xor U3792 (N_3792,In_1538,In_2302);
or U3793 (N_3793,In_1591,In_2187);
xnor U3794 (N_3794,In_1450,In_1134);
or U3795 (N_3795,In_1163,In_129);
and U3796 (N_3796,In_958,In_414);
nor U3797 (N_3797,In_2145,In_598);
and U3798 (N_3798,In_724,In_2085);
or U3799 (N_3799,In_453,In_564);
nor U3800 (N_3800,In_622,In_1882);
nor U3801 (N_3801,In_1458,In_815);
or U3802 (N_3802,In_1700,In_2459);
nand U3803 (N_3803,In_2417,In_1924);
or U3804 (N_3804,In_733,In_1362);
xor U3805 (N_3805,In_2221,In_1151);
nor U3806 (N_3806,In_1022,In_994);
nand U3807 (N_3807,In_972,In_888);
xor U3808 (N_3808,In_2243,In_36);
or U3809 (N_3809,In_1128,In_176);
and U3810 (N_3810,In_169,In_936);
nor U3811 (N_3811,In_1552,In_1347);
and U3812 (N_3812,In_2153,In_1789);
nand U3813 (N_3813,In_66,In_642);
nand U3814 (N_3814,In_272,In_1751);
xor U3815 (N_3815,In_682,In_692);
nand U3816 (N_3816,In_535,In_1194);
or U3817 (N_3817,In_311,In_805);
and U3818 (N_3818,In_2362,In_1222);
nor U3819 (N_3819,In_1692,In_1439);
nor U3820 (N_3820,In_1717,In_1938);
nand U3821 (N_3821,In_1073,In_1790);
nand U3822 (N_3822,In_1393,In_1568);
and U3823 (N_3823,In_1248,In_434);
nor U3824 (N_3824,In_746,In_2041);
nor U3825 (N_3825,In_621,In_1435);
and U3826 (N_3826,In_816,In_2428);
or U3827 (N_3827,In_2254,In_477);
xor U3828 (N_3828,In_378,In_417);
xor U3829 (N_3829,In_1716,In_2102);
xor U3830 (N_3830,In_1890,In_1273);
xnor U3831 (N_3831,In_843,In_1151);
xnor U3832 (N_3832,In_264,In_353);
or U3833 (N_3833,In_2075,In_2067);
and U3834 (N_3834,In_2034,In_260);
nor U3835 (N_3835,In_2345,In_1072);
and U3836 (N_3836,In_2023,In_918);
and U3837 (N_3837,In_2000,In_834);
or U3838 (N_3838,In_1432,In_2300);
xor U3839 (N_3839,In_2185,In_2286);
xnor U3840 (N_3840,In_2322,In_1767);
xor U3841 (N_3841,In_21,In_1685);
and U3842 (N_3842,In_193,In_2026);
nor U3843 (N_3843,In_132,In_131);
and U3844 (N_3844,In_898,In_2463);
nand U3845 (N_3845,In_1408,In_1350);
nand U3846 (N_3846,In_757,In_2109);
and U3847 (N_3847,In_2030,In_1450);
nor U3848 (N_3848,In_1235,In_563);
nor U3849 (N_3849,In_1948,In_1158);
or U3850 (N_3850,In_2269,In_2411);
or U3851 (N_3851,In_591,In_78);
nor U3852 (N_3852,In_96,In_1295);
and U3853 (N_3853,In_1486,In_1992);
nor U3854 (N_3854,In_386,In_2247);
xor U3855 (N_3855,In_424,In_314);
xor U3856 (N_3856,In_2177,In_981);
and U3857 (N_3857,In_460,In_1513);
nor U3858 (N_3858,In_1300,In_1198);
or U3859 (N_3859,In_881,In_1150);
xor U3860 (N_3860,In_820,In_1988);
nor U3861 (N_3861,In_114,In_1362);
and U3862 (N_3862,In_1294,In_1329);
nor U3863 (N_3863,In_333,In_2445);
or U3864 (N_3864,In_169,In_1077);
and U3865 (N_3865,In_2474,In_1182);
nor U3866 (N_3866,In_2363,In_396);
xor U3867 (N_3867,In_6,In_471);
xnor U3868 (N_3868,In_329,In_1209);
xor U3869 (N_3869,In_240,In_1023);
nor U3870 (N_3870,In_39,In_704);
and U3871 (N_3871,In_310,In_382);
or U3872 (N_3872,In_1096,In_121);
nor U3873 (N_3873,In_2344,In_563);
and U3874 (N_3874,In_1421,In_296);
nand U3875 (N_3875,In_1767,In_748);
nand U3876 (N_3876,In_2478,In_2030);
or U3877 (N_3877,In_1271,In_1452);
and U3878 (N_3878,In_2400,In_1889);
or U3879 (N_3879,In_2029,In_1860);
xnor U3880 (N_3880,In_1108,In_281);
and U3881 (N_3881,In_390,In_260);
nand U3882 (N_3882,In_382,In_1020);
and U3883 (N_3883,In_265,In_879);
nor U3884 (N_3884,In_916,In_1225);
or U3885 (N_3885,In_2335,In_1976);
xor U3886 (N_3886,In_756,In_1408);
nor U3887 (N_3887,In_965,In_2376);
and U3888 (N_3888,In_308,In_279);
or U3889 (N_3889,In_706,In_137);
and U3890 (N_3890,In_247,In_1336);
or U3891 (N_3891,In_2469,In_941);
and U3892 (N_3892,In_117,In_2231);
nor U3893 (N_3893,In_1793,In_1529);
nor U3894 (N_3894,In_899,In_696);
or U3895 (N_3895,In_1149,In_1971);
xnor U3896 (N_3896,In_671,In_829);
and U3897 (N_3897,In_764,In_834);
nand U3898 (N_3898,In_432,In_1616);
nor U3899 (N_3899,In_1485,In_1937);
nor U3900 (N_3900,In_1751,In_857);
xor U3901 (N_3901,In_2040,In_783);
nor U3902 (N_3902,In_1569,In_343);
nand U3903 (N_3903,In_1574,In_47);
or U3904 (N_3904,In_26,In_2412);
or U3905 (N_3905,In_2134,In_748);
nor U3906 (N_3906,In_1237,In_1987);
nor U3907 (N_3907,In_1621,In_309);
and U3908 (N_3908,In_1010,In_9);
and U3909 (N_3909,In_2242,In_77);
nand U3910 (N_3910,In_909,In_216);
nand U3911 (N_3911,In_417,In_1508);
and U3912 (N_3912,In_67,In_1267);
or U3913 (N_3913,In_1482,In_2161);
xor U3914 (N_3914,In_1819,In_1673);
or U3915 (N_3915,In_496,In_593);
xnor U3916 (N_3916,In_1834,In_2234);
and U3917 (N_3917,In_118,In_234);
and U3918 (N_3918,In_1783,In_1402);
and U3919 (N_3919,In_989,In_1652);
xnor U3920 (N_3920,In_828,In_1262);
and U3921 (N_3921,In_167,In_1741);
nor U3922 (N_3922,In_2454,In_1893);
or U3923 (N_3923,In_579,In_1380);
or U3924 (N_3924,In_2161,In_219);
and U3925 (N_3925,In_2365,In_1694);
or U3926 (N_3926,In_1652,In_553);
and U3927 (N_3927,In_2321,In_1994);
nor U3928 (N_3928,In_2230,In_812);
or U3929 (N_3929,In_1850,In_94);
nor U3930 (N_3930,In_1259,In_438);
or U3931 (N_3931,In_984,In_1402);
xor U3932 (N_3932,In_968,In_2366);
nor U3933 (N_3933,In_2391,In_1920);
and U3934 (N_3934,In_365,In_1429);
nor U3935 (N_3935,In_1929,In_288);
nand U3936 (N_3936,In_661,In_322);
nand U3937 (N_3937,In_27,In_791);
or U3938 (N_3938,In_908,In_1696);
xnor U3939 (N_3939,In_943,In_1307);
or U3940 (N_3940,In_2168,In_2336);
xnor U3941 (N_3941,In_1689,In_419);
xnor U3942 (N_3942,In_273,In_2051);
or U3943 (N_3943,In_2132,In_2468);
nand U3944 (N_3944,In_571,In_1923);
and U3945 (N_3945,In_981,In_1475);
xor U3946 (N_3946,In_168,In_1911);
xor U3947 (N_3947,In_1151,In_1353);
and U3948 (N_3948,In_2329,In_193);
and U3949 (N_3949,In_1993,In_1275);
or U3950 (N_3950,In_2137,In_1991);
or U3951 (N_3951,In_1479,In_1220);
nand U3952 (N_3952,In_910,In_1509);
or U3953 (N_3953,In_723,In_318);
or U3954 (N_3954,In_1107,In_1966);
and U3955 (N_3955,In_363,In_1816);
nor U3956 (N_3956,In_1807,In_794);
nand U3957 (N_3957,In_650,In_2236);
or U3958 (N_3958,In_1361,In_2465);
xnor U3959 (N_3959,In_1484,In_903);
nand U3960 (N_3960,In_1880,In_344);
xor U3961 (N_3961,In_2201,In_2064);
xnor U3962 (N_3962,In_2280,In_297);
and U3963 (N_3963,In_1500,In_1264);
nand U3964 (N_3964,In_2209,In_1005);
and U3965 (N_3965,In_439,In_2296);
nor U3966 (N_3966,In_696,In_1754);
nor U3967 (N_3967,In_780,In_280);
and U3968 (N_3968,In_1816,In_95);
xor U3969 (N_3969,In_918,In_494);
nor U3970 (N_3970,In_1611,In_847);
nor U3971 (N_3971,In_1258,In_1424);
or U3972 (N_3972,In_1251,In_1775);
and U3973 (N_3973,In_1813,In_744);
or U3974 (N_3974,In_878,In_173);
nor U3975 (N_3975,In_1983,In_698);
nor U3976 (N_3976,In_281,In_436);
nand U3977 (N_3977,In_2169,In_418);
nand U3978 (N_3978,In_36,In_1492);
or U3979 (N_3979,In_1114,In_1471);
nand U3980 (N_3980,In_2471,In_836);
xnor U3981 (N_3981,In_916,In_579);
nor U3982 (N_3982,In_1781,In_1592);
and U3983 (N_3983,In_1616,In_696);
xor U3984 (N_3984,In_1958,In_2182);
nand U3985 (N_3985,In_2416,In_845);
nor U3986 (N_3986,In_365,In_842);
nor U3987 (N_3987,In_1776,In_379);
and U3988 (N_3988,In_552,In_625);
and U3989 (N_3989,In_400,In_1032);
or U3990 (N_3990,In_2248,In_2188);
nor U3991 (N_3991,In_1688,In_2287);
xor U3992 (N_3992,In_1029,In_1425);
or U3993 (N_3993,In_1744,In_2106);
and U3994 (N_3994,In_1588,In_1724);
nand U3995 (N_3995,In_1197,In_969);
nor U3996 (N_3996,In_578,In_2262);
or U3997 (N_3997,In_1688,In_1317);
xor U3998 (N_3998,In_525,In_1608);
xnor U3999 (N_3999,In_2097,In_325);
and U4000 (N_4000,In_1712,In_2320);
or U4001 (N_4001,In_391,In_1764);
and U4002 (N_4002,In_1770,In_780);
nor U4003 (N_4003,In_1007,In_1784);
nand U4004 (N_4004,In_1818,In_2366);
nand U4005 (N_4005,In_1439,In_1191);
or U4006 (N_4006,In_842,In_1900);
and U4007 (N_4007,In_461,In_209);
and U4008 (N_4008,In_2258,In_777);
or U4009 (N_4009,In_1729,In_2479);
or U4010 (N_4010,In_2357,In_92);
nand U4011 (N_4011,In_479,In_1622);
nand U4012 (N_4012,In_697,In_2486);
xnor U4013 (N_4013,In_1289,In_2159);
or U4014 (N_4014,In_1587,In_1247);
xor U4015 (N_4015,In_11,In_333);
nand U4016 (N_4016,In_1665,In_260);
nand U4017 (N_4017,In_1780,In_314);
nand U4018 (N_4018,In_787,In_798);
nand U4019 (N_4019,In_1689,In_582);
nor U4020 (N_4020,In_969,In_1894);
and U4021 (N_4021,In_897,In_2163);
nand U4022 (N_4022,In_86,In_2435);
xor U4023 (N_4023,In_261,In_2203);
or U4024 (N_4024,In_446,In_2254);
nor U4025 (N_4025,In_1801,In_383);
and U4026 (N_4026,In_774,In_2419);
nand U4027 (N_4027,In_871,In_269);
xor U4028 (N_4028,In_1737,In_678);
nor U4029 (N_4029,In_131,In_2226);
xor U4030 (N_4030,In_1718,In_2167);
nor U4031 (N_4031,In_964,In_2036);
nand U4032 (N_4032,In_1942,In_771);
nor U4033 (N_4033,In_571,In_288);
nor U4034 (N_4034,In_283,In_1389);
nor U4035 (N_4035,In_887,In_9);
and U4036 (N_4036,In_1506,In_1307);
nor U4037 (N_4037,In_1883,In_1277);
or U4038 (N_4038,In_971,In_1017);
or U4039 (N_4039,In_2395,In_1457);
and U4040 (N_4040,In_2202,In_1483);
nor U4041 (N_4041,In_68,In_594);
or U4042 (N_4042,In_561,In_2462);
nand U4043 (N_4043,In_402,In_1095);
or U4044 (N_4044,In_192,In_648);
or U4045 (N_4045,In_388,In_731);
xor U4046 (N_4046,In_1880,In_2103);
nand U4047 (N_4047,In_517,In_1578);
and U4048 (N_4048,In_1454,In_1152);
nand U4049 (N_4049,In_657,In_2312);
and U4050 (N_4050,In_715,In_1781);
and U4051 (N_4051,In_1632,In_1066);
xor U4052 (N_4052,In_353,In_886);
nand U4053 (N_4053,In_1820,In_2409);
nand U4054 (N_4054,In_2014,In_1084);
and U4055 (N_4055,In_2265,In_1680);
nor U4056 (N_4056,In_1581,In_2029);
nand U4057 (N_4057,In_1987,In_2331);
or U4058 (N_4058,In_277,In_555);
nor U4059 (N_4059,In_1739,In_2046);
xnor U4060 (N_4060,In_751,In_1311);
nor U4061 (N_4061,In_699,In_319);
nor U4062 (N_4062,In_1575,In_235);
or U4063 (N_4063,In_1928,In_92);
nand U4064 (N_4064,In_1918,In_975);
nand U4065 (N_4065,In_228,In_478);
nor U4066 (N_4066,In_339,In_1576);
nor U4067 (N_4067,In_1745,In_948);
or U4068 (N_4068,In_1167,In_1298);
or U4069 (N_4069,In_2488,In_595);
nor U4070 (N_4070,In_2497,In_2247);
or U4071 (N_4071,In_795,In_1491);
or U4072 (N_4072,In_2107,In_2253);
or U4073 (N_4073,In_2466,In_2226);
nand U4074 (N_4074,In_875,In_1258);
and U4075 (N_4075,In_2443,In_2236);
and U4076 (N_4076,In_728,In_1062);
xor U4077 (N_4077,In_631,In_435);
or U4078 (N_4078,In_433,In_1295);
xnor U4079 (N_4079,In_2474,In_994);
xor U4080 (N_4080,In_154,In_399);
nand U4081 (N_4081,In_850,In_803);
or U4082 (N_4082,In_552,In_2363);
or U4083 (N_4083,In_1844,In_62);
or U4084 (N_4084,In_1694,In_678);
nand U4085 (N_4085,In_350,In_994);
nand U4086 (N_4086,In_1764,In_1766);
or U4087 (N_4087,In_457,In_1380);
nand U4088 (N_4088,In_2384,In_995);
nor U4089 (N_4089,In_325,In_1814);
xnor U4090 (N_4090,In_1121,In_1522);
nor U4091 (N_4091,In_894,In_932);
xor U4092 (N_4092,In_1528,In_40);
xnor U4093 (N_4093,In_1224,In_1668);
xnor U4094 (N_4094,In_2260,In_265);
and U4095 (N_4095,In_1382,In_2233);
and U4096 (N_4096,In_1753,In_1635);
and U4097 (N_4097,In_876,In_550);
and U4098 (N_4098,In_2490,In_2206);
xor U4099 (N_4099,In_382,In_1282);
and U4100 (N_4100,In_9,In_181);
nor U4101 (N_4101,In_390,In_2429);
nand U4102 (N_4102,In_1294,In_1142);
or U4103 (N_4103,In_636,In_1802);
nand U4104 (N_4104,In_1648,In_1988);
nand U4105 (N_4105,In_2082,In_70);
and U4106 (N_4106,In_91,In_259);
xor U4107 (N_4107,In_341,In_118);
xnor U4108 (N_4108,In_1771,In_1184);
or U4109 (N_4109,In_1892,In_2168);
nor U4110 (N_4110,In_1500,In_337);
and U4111 (N_4111,In_244,In_352);
and U4112 (N_4112,In_135,In_793);
nor U4113 (N_4113,In_2320,In_433);
xor U4114 (N_4114,In_2484,In_2252);
and U4115 (N_4115,In_1050,In_1140);
xnor U4116 (N_4116,In_1100,In_728);
nand U4117 (N_4117,In_1309,In_1488);
nand U4118 (N_4118,In_1516,In_1977);
and U4119 (N_4119,In_530,In_588);
and U4120 (N_4120,In_2116,In_191);
nand U4121 (N_4121,In_1554,In_2147);
and U4122 (N_4122,In_769,In_2398);
nor U4123 (N_4123,In_273,In_1409);
or U4124 (N_4124,In_1534,In_898);
or U4125 (N_4125,In_498,In_951);
nand U4126 (N_4126,In_949,In_1978);
and U4127 (N_4127,In_2183,In_554);
and U4128 (N_4128,In_678,In_1968);
and U4129 (N_4129,In_1835,In_842);
xor U4130 (N_4130,In_1100,In_1706);
nand U4131 (N_4131,In_1959,In_1191);
nand U4132 (N_4132,In_572,In_1300);
and U4133 (N_4133,In_1450,In_1513);
or U4134 (N_4134,In_1403,In_1857);
nor U4135 (N_4135,In_2003,In_1877);
or U4136 (N_4136,In_1785,In_147);
nand U4137 (N_4137,In_1950,In_181);
or U4138 (N_4138,In_1145,In_1792);
xnor U4139 (N_4139,In_559,In_1283);
or U4140 (N_4140,In_865,In_1250);
nand U4141 (N_4141,In_693,In_2243);
xnor U4142 (N_4142,In_868,In_1322);
nand U4143 (N_4143,In_2308,In_1410);
and U4144 (N_4144,In_1044,In_441);
nor U4145 (N_4145,In_401,In_1952);
nand U4146 (N_4146,In_612,In_1270);
and U4147 (N_4147,In_2213,In_1634);
and U4148 (N_4148,In_1149,In_1348);
and U4149 (N_4149,In_319,In_1943);
nor U4150 (N_4150,In_15,In_397);
or U4151 (N_4151,In_1521,In_1871);
nand U4152 (N_4152,In_808,In_711);
xor U4153 (N_4153,In_786,In_2075);
and U4154 (N_4154,In_1430,In_800);
nor U4155 (N_4155,In_967,In_203);
xnor U4156 (N_4156,In_1978,In_2222);
xnor U4157 (N_4157,In_1610,In_1698);
nand U4158 (N_4158,In_327,In_1998);
xnor U4159 (N_4159,In_2025,In_759);
nand U4160 (N_4160,In_1354,In_550);
or U4161 (N_4161,In_155,In_1143);
xnor U4162 (N_4162,In_65,In_660);
or U4163 (N_4163,In_1831,In_2093);
nor U4164 (N_4164,In_1083,In_709);
and U4165 (N_4165,In_1215,In_1899);
nand U4166 (N_4166,In_2248,In_1812);
nand U4167 (N_4167,In_1209,In_1828);
or U4168 (N_4168,In_1840,In_2002);
xnor U4169 (N_4169,In_1610,In_302);
xnor U4170 (N_4170,In_2414,In_552);
and U4171 (N_4171,In_986,In_1390);
nor U4172 (N_4172,In_1771,In_931);
or U4173 (N_4173,In_463,In_595);
nor U4174 (N_4174,In_2107,In_801);
nor U4175 (N_4175,In_577,In_2390);
nand U4176 (N_4176,In_2170,In_861);
xnor U4177 (N_4177,In_1944,In_1758);
and U4178 (N_4178,In_2477,In_2077);
nand U4179 (N_4179,In_1891,In_301);
or U4180 (N_4180,In_2257,In_2061);
or U4181 (N_4181,In_203,In_1791);
xnor U4182 (N_4182,In_1371,In_2117);
and U4183 (N_4183,In_1251,In_370);
or U4184 (N_4184,In_1792,In_1776);
nand U4185 (N_4185,In_1040,In_1298);
and U4186 (N_4186,In_1835,In_2067);
nand U4187 (N_4187,In_1853,In_278);
or U4188 (N_4188,In_1749,In_1144);
nand U4189 (N_4189,In_1720,In_739);
and U4190 (N_4190,In_2187,In_1907);
or U4191 (N_4191,In_332,In_2462);
or U4192 (N_4192,In_210,In_1378);
nor U4193 (N_4193,In_2179,In_903);
or U4194 (N_4194,In_707,In_2411);
nand U4195 (N_4195,In_2135,In_1083);
or U4196 (N_4196,In_1239,In_159);
xnor U4197 (N_4197,In_688,In_2248);
and U4198 (N_4198,In_97,In_1786);
or U4199 (N_4199,In_936,In_80);
nor U4200 (N_4200,In_2407,In_1285);
xnor U4201 (N_4201,In_541,In_1868);
or U4202 (N_4202,In_940,In_1850);
nand U4203 (N_4203,In_519,In_746);
xor U4204 (N_4204,In_1337,In_2165);
nor U4205 (N_4205,In_858,In_293);
nor U4206 (N_4206,In_1251,In_2407);
nand U4207 (N_4207,In_380,In_2294);
or U4208 (N_4208,In_149,In_1733);
xnor U4209 (N_4209,In_1831,In_2289);
nor U4210 (N_4210,In_1728,In_522);
xnor U4211 (N_4211,In_475,In_1091);
nor U4212 (N_4212,In_2077,In_182);
and U4213 (N_4213,In_1249,In_1581);
xnor U4214 (N_4214,In_564,In_884);
xor U4215 (N_4215,In_591,In_1006);
nor U4216 (N_4216,In_746,In_144);
nor U4217 (N_4217,In_1573,In_1251);
or U4218 (N_4218,In_1180,In_1971);
xor U4219 (N_4219,In_1238,In_1378);
and U4220 (N_4220,In_1990,In_1334);
nand U4221 (N_4221,In_2341,In_1479);
and U4222 (N_4222,In_1017,In_690);
nor U4223 (N_4223,In_1360,In_1900);
or U4224 (N_4224,In_1065,In_362);
xor U4225 (N_4225,In_2035,In_1123);
nor U4226 (N_4226,In_2093,In_1009);
nor U4227 (N_4227,In_2417,In_840);
nand U4228 (N_4228,In_1927,In_2090);
and U4229 (N_4229,In_2034,In_2193);
or U4230 (N_4230,In_1424,In_1782);
nor U4231 (N_4231,In_1175,In_1678);
xor U4232 (N_4232,In_696,In_354);
xor U4233 (N_4233,In_14,In_184);
nand U4234 (N_4234,In_2310,In_737);
nand U4235 (N_4235,In_153,In_15);
xor U4236 (N_4236,In_2227,In_2359);
or U4237 (N_4237,In_318,In_144);
or U4238 (N_4238,In_1917,In_1764);
and U4239 (N_4239,In_1170,In_1246);
nand U4240 (N_4240,In_1548,In_58);
or U4241 (N_4241,In_505,In_867);
xor U4242 (N_4242,In_1917,In_585);
and U4243 (N_4243,In_437,In_965);
nor U4244 (N_4244,In_2072,In_1709);
xor U4245 (N_4245,In_2130,In_2146);
xor U4246 (N_4246,In_511,In_2052);
or U4247 (N_4247,In_788,In_1675);
or U4248 (N_4248,In_962,In_1470);
xor U4249 (N_4249,In_406,In_1430);
nand U4250 (N_4250,In_1830,In_1613);
or U4251 (N_4251,In_622,In_2439);
xor U4252 (N_4252,In_1658,In_142);
nor U4253 (N_4253,In_2190,In_1966);
or U4254 (N_4254,In_1415,In_744);
and U4255 (N_4255,In_909,In_763);
and U4256 (N_4256,In_340,In_1227);
or U4257 (N_4257,In_155,In_1432);
or U4258 (N_4258,In_2329,In_512);
xnor U4259 (N_4259,In_1999,In_1264);
nand U4260 (N_4260,In_731,In_1964);
and U4261 (N_4261,In_1554,In_709);
nand U4262 (N_4262,In_1666,In_1174);
or U4263 (N_4263,In_2269,In_801);
nor U4264 (N_4264,In_688,In_2081);
and U4265 (N_4265,In_93,In_2226);
nand U4266 (N_4266,In_755,In_882);
nor U4267 (N_4267,In_1280,In_1998);
or U4268 (N_4268,In_2276,In_1053);
nand U4269 (N_4269,In_277,In_1811);
and U4270 (N_4270,In_531,In_1107);
nor U4271 (N_4271,In_1635,In_504);
xnor U4272 (N_4272,In_195,In_2122);
nand U4273 (N_4273,In_235,In_797);
xnor U4274 (N_4274,In_1327,In_1358);
xor U4275 (N_4275,In_1276,In_827);
and U4276 (N_4276,In_2265,In_1834);
and U4277 (N_4277,In_1665,In_1772);
or U4278 (N_4278,In_2373,In_1038);
nor U4279 (N_4279,In_1095,In_2335);
and U4280 (N_4280,In_562,In_1312);
xor U4281 (N_4281,In_1843,In_1551);
xor U4282 (N_4282,In_1968,In_551);
and U4283 (N_4283,In_280,In_1330);
and U4284 (N_4284,In_1769,In_614);
nor U4285 (N_4285,In_2071,In_1865);
xnor U4286 (N_4286,In_24,In_1559);
and U4287 (N_4287,In_1182,In_1916);
and U4288 (N_4288,In_1548,In_1711);
and U4289 (N_4289,In_1166,In_1899);
nor U4290 (N_4290,In_1846,In_2491);
or U4291 (N_4291,In_757,In_1019);
and U4292 (N_4292,In_2360,In_2211);
xor U4293 (N_4293,In_1610,In_378);
xnor U4294 (N_4294,In_243,In_1043);
nand U4295 (N_4295,In_2448,In_1980);
and U4296 (N_4296,In_1536,In_651);
or U4297 (N_4297,In_952,In_408);
nand U4298 (N_4298,In_306,In_612);
or U4299 (N_4299,In_901,In_1503);
nand U4300 (N_4300,In_85,In_2198);
xnor U4301 (N_4301,In_2488,In_905);
nor U4302 (N_4302,In_742,In_2182);
and U4303 (N_4303,In_1822,In_936);
xnor U4304 (N_4304,In_2314,In_1255);
and U4305 (N_4305,In_682,In_1703);
nand U4306 (N_4306,In_930,In_2362);
nand U4307 (N_4307,In_845,In_1118);
nor U4308 (N_4308,In_831,In_667);
nor U4309 (N_4309,In_1278,In_1921);
and U4310 (N_4310,In_2251,In_387);
or U4311 (N_4311,In_809,In_25);
nand U4312 (N_4312,In_184,In_1579);
nor U4313 (N_4313,In_692,In_1344);
nor U4314 (N_4314,In_1674,In_1051);
xor U4315 (N_4315,In_1994,In_353);
nor U4316 (N_4316,In_1911,In_399);
nand U4317 (N_4317,In_933,In_1590);
nor U4318 (N_4318,In_79,In_1369);
xnor U4319 (N_4319,In_1308,In_2130);
nor U4320 (N_4320,In_716,In_945);
or U4321 (N_4321,In_943,In_1157);
nand U4322 (N_4322,In_1674,In_525);
nor U4323 (N_4323,In_2161,In_390);
nor U4324 (N_4324,In_1579,In_2145);
and U4325 (N_4325,In_619,In_522);
and U4326 (N_4326,In_125,In_1329);
nand U4327 (N_4327,In_2228,In_89);
or U4328 (N_4328,In_1891,In_1224);
xor U4329 (N_4329,In_1980,In_2479);
or U4330 (N_4330,In_1133,In_2132);
xnor U4331 (N_4331,In_168,In_2015);
or U4332 (N_4332,In_1094,In_1141);
and U4333 (N_4333,In_117,In_2220);
nand U4334 (N_4334,In_1245,In_1292);
nand U4335 (N_4335,In_1505,In_2311);
nor U4336 (N_4336,In_153,In_746);
nand U4337 (N_4337,In_830,In_140);
or U4338 (N_4338,In_404,In_1052);
nand U4339 (N_4339,In_1989,In_1137);
and U4340 (N_4340,In_2401,In_210);
or U4341 (N_4341,In_121,In_870);
nand U4342 (N_4342,In_2349,In_1288);
or U4343 (N_4343,In_748,In_1038);
or U4344 (N_4344,In_1707,In_2470);
or U4345 (N_4345,In_1490,In_430);
nor U4346 (N_4346,In_792,In_1056);
or U4347 (N_4347,In_702,In_1026);
xor U4348 (N_4348,In_427,In_972);
and U4349 (N_4349,In_1526,In_2228);
nand U4350 (N_4350,In_1078,In_234);
nand U4351 (N_4351,In_917,In_815);
xor U4352 (N_4352,In_1768,In_1830);
nand U4353 (N_4353,In_764,In_2192);
nor U4354 (N_4354,In_1045,In_1486);
nor U4355 (N_4355,In_799,In_96);
xnor U4356 (N_4356,In_1025,In_1977);
nand U4357 (N_4357,In_1909,In_1239);
xor U4358 (N_4358,In_263,In_530);
nand U4359 (N_4359,In_90,In_658);
nor U4360 (N_4360,In_455,In_2327);
nand U4361 (N_4361,In_2467,In_2418);
nand U4362 (N_4362,In_234,In_279);
nand U4363 (N_4363,In_1662,In_2122);
nand U4364 (N_4364,In_1804,In_284);
or U4365 (N_4365,In_668,In_1732);
and U4366 (N_4366,In_1829,In_2057);
or U4367 (N_4367,In_91,In_76);
nand U4368 (N_4368,In_700,In_1114);
xor U4369 (N_4369,In_1369,In_1755);
and U4370 (N_4370,In_2097,In_2056);
and U4371 (N_4371,In_2442,In_682);
xor U4372 (N_4372,In_2327,In_1546);
nor U4373 (N_4373,In_1380,In_2015);
xor U4374 (N_4374,In_1202,In_930);
and U4375 (N_4375,In_459,In_581);
or U4376 (N_4376,In_344,In_383);
nor U4377 (N_4377,In_1192,In_213);
and U4378 (N_4378,In_1141,In_779);
or U4379 (N_4379,In_1293,In_844);
and U4380 (N_4380,In_1517,In_2116);
or U4381 (N_4381,In_1756,In_305);
nand U4382 (N_4382,In_432,In_2011);
xnor U4383 (N_4383,In_1340,In_1300);
or U4384 (N_4384,In_624,In_237);
or U4385 (N_4385,In_1307,In_2476);
nand U4386 (N_4386,In_1870,In_255);
and U4387 (N_4387,In_2037,In_179);
or U4388 (N_4388,In_2032,In_2461);
xnor U4389 (N_4389,In_2368,In_1751);
and U4390 (N_4390,In_1911,In_908);
nand U4391 (N_4391,In_2150,In_327);
nand U4392 (N_4392,In_2191,In_706);
or U4393 (N_4393,In_1715,In_1912);
xnor U4394 (N_4394,In_741,In_125);
nor U4395 (N_4395,In_2272,In_710);
nor U4396 (N_4396,In_663,In_1980);
nand U4397 (N_4397,In_2029,In_609);
and U4398 (N_4398,In_2170,In_1269);
nand U4399 (N_4399,In_223,In_1086);
nor U4400 (N_4400,In_992,In_959);
xnor U4401 (N_4401,In_34,In_684);
and U4402 (N_4402,In_2160,In_1108);
nor U4403 (N_4403,In_1191,In_954);
nand U4404 (N_4404,In_2188,In_123);
xnor U4405 (N_4405,In_640,In_543);
or U4406 (N_4406,In_554,In_1186);
xnor U4407 (N_4407,In_1398,In_419);
nand U4408 (N_4408,In_1294,In_385);
or U4409 (N_4409,In_435,In_2447);
nand U4410 (N_4410,In_784,In_857);
and U4411 (N_4411,In_1316,In_51);
nor U4412 (N_4412,In_304,In_2366);
nor U4413 (N_4413,In_857,In_1399);
and U4414 (N_4414,In_1385,In_1657);
nand U4415 (N_4415,In_876,In_399);
and U4416 (N_4416,In_468,In_1067);
or U4417 (N_4417,In_1271,In_2369);
nor U4418 (N_4418,In_519,In_2067);
nor U4419 (N_4419,In_613,In_865);
nand U4420 (N_4420,In_1672,In_1607);
or U4421 (N_4421,In_832,In_1615);
or U4422 (N_4422,In_1098,In_1107);
nor U4423 (N_4423,In_1929,In_661);
xor U4424 (N_4424,In_42,In_964);
nor U4425 (N_4425,In_2485,In_303);
xor U4426 (N_4426,In_2273,In_1214);
and U4427 (N_4427,In_203,In_2251);
and U4428 (N_4428,In_2114,In_1074);
nor U4429 (N_4429,In_1708,In_553);
nand U4430 (N_4430,In_31,In_574);
xnor U4431 (N_4431,In_558,In_1960);
nor U4432 (N_4432,In_2465,In_868);
xor U4433 (N_4433,In_1556,In_1998);
xnor U4434 (N_4434,In_902,In_1790);
or U4435 (N_4435,In_2436,In_985);
nor U4436 (N_4436,In_2214,In_1639);
or U4437 (N_4437,In_998,In_2064);
or U4438 (N_4438,In_674,In_962);
or U4439 (N_4439,In_437,In_1054);
and U4440 (N_4440,In_2474,In_1281);
nor U4441 (N_4441,In_776,In_85);
nand U4442 (N_4442,In_1693,In_221);
xor U4443 (N_4443,In_1314,In_1502);
or U4444 (N_4444,In_992,In_1795);
xnor U4445 (N_4445,In_2414,In_2212);
xor U4446 (N_4446,In_219,In_271);
and U4447 (N_4447,In_1356,In_2360);
xor U4448 (N_4448,In_1809,In_18);
or U4449 (N_4449,In_2173,In_1007);
xnor U4450 (N_4450,In_2225,In_1109);
nand U4451 (N_4451,In_437,In_2148);
nor U4452 (N_4452,In_257,In_1787);
or U4453 (N_4453,In_1515,In_100);
or U4454 (N_4454,In_1013,In_1537);
and U4455 (N_4455,In_2464,In_50);
nor U4456 (N_4456,In_2378,In_2276);
or U4457 (N_4457,In_2004,In_1242);
nor U4458 (N_4458,In_756,In_1776);
or U4459 (N_4459,In_118,In_1613);
nor U4460 (N_4460,In_2051,In_1902);
nand U4461 (N_4461,In_1845,In_1367);
nor U4462 (N_4462,In_14,In_1225);
and U4463 (N_4463,In_134,In_741);
nand U4464 (N_4464,In_2404,In_1687);
or U4465 (N_4465,In_271,In_679);
nand U4466 (N_4466,In_1931,In_125);
or U4467 (N_4467,In_1551,In_686);
nor U4468 (N_4468,In_42,In_2450);
xor U4469 (N_4469,In_409,In_1982);
nor U4470 (N_4470,In_431,In_1921);
or U4471 (N_4471,In_602,In_74);
nor U4472 (N_4472,In_1343,In_911);
xnor U4473 (N_4473,In_266,In_1667);
and U4474 (N_4474,In_905,In_1523);
nand U4475 (N_4475,In_715,In_2446);
or U4476 (N_4476,In_338,In_1256);
or U4477 (N_4477,In_627,In_2353);
and U4478 (N_4478,In_697,In_216);
or U4479 (N_4479,In_1612,In_229);
nor U4480 (N_4480,In_772,In_722);
nand U4481 (N_4481,In_886,In_1926);
and U4482 (N_4482,In_2437,In_2131);
and U4483 (N_4483,In_2488,In_107);
and U4484 (N_4484,In_1581,In_446);
nor U4485 (N_4485,In_132,In_889);
nor U4486 (N_4486,In_1247,In_99);
and U4487 (N_4487,In_882,In_495);
xnor U4488 (N_4488,In_900,In_2125);
nor U4489 (N_4489,In_931,In_2473);
xnor U4490 (N_4490,In_2196,In_1029);
nor U4491 (N_4491,In_2456,In_225);
nor U4492 (N_4492,In_432,In_1480);
and U4493 (N_4493,In_1257,In_1081);
nor U4494 (N_4494,In_850,In_2352);
nand U4495 (N_4495,In_1241,In_1534);
nor U4496 (N_4496,In_406,In_951);
and U4497 (N_4497,In_909,In_1715);
xnor U4498 (N_4498,In_777,In_1196);
nand U4499 (N_4499,In_387,In_1937);
or U4500 (N_4500,In_1290,In_299);
nor U4501 (N_4501,In_1014,In_752);
nand U4502 (N_4502,In_1824,In_1450);
or U4503 (N_4503,In_1586,In_1318);
nor U4504 (N_4504,In_681,In_833);
nand U4505 (N_4505,In_2319,In_1517);
nor U4506 (N_4506,In_900,In_1258);
nor U4507 (N_4507,In_166,In_2074);
or U4508 (N_4508,In_839,In_109);
xnor U4509 (N_4509,In_2184,In_1941);
nand U4510 (N_4510,In_1278,In_696);
and U4511 (N_4511,In_853,In_324);
xor U4512 (N_4512,In_2110,In_540);
or U4513 (N_4513,In_571,In_915);
and U4514 (N_4514,In_1392,In_527);
or U4515 (N_4515,In_1651,In_124);
xor U4516 (N_4516,In_1457,In_1725);
nand U4517 (N_4517,In_418,In_840);
and U4518 (N_4518,In_120,In_1880);
or U4519 (N_4519,In_2326,In_486);
and U4520 (N_4520,In_747,In_1458);
or U4521 (N_4521,In_1786,In_1935);
xnor U4522 (N_4522,In_1793,In_754);
and U4523 (N_4523,In_921,In_2043);
nor U4524 (N_4524,In_1414,In_2058);
and U4525 (N_4525,In_1769,In_839);
nor U4526 (N_4526,In_1104,In_554);
nor U4527 (N_4527,In_442,In_2346);
nor U4528 (N_4528,In_1309,In_2231);
or U4529 (N_4529,In_999,In_910);
nor U4530 (N_4530,In_362,In_1444);
and U4531 (N_4531,In_788,In_2023);
nand U4532 (N_4532,In_1498,In_286);
or U4533 (N_4533,In_2482,In_1260);
or U4534 (N_4534,In_83,In_1909);
or U4535 (N_4535,In_2393,In_502);
and U4536 (N_4536,In_1706,In_1035);
nor U4537 (N_4537,In_711,In_1818);
xnor U4538 (N_4538,In_1606,In_2023);
or U4539 (N_4539,In_75,In_578);
or U4540 (N_4540,In_1648,In_28);
nand U4541 (N_4541,In_1911,In_534);
nand U4542 (N_4542,In_871,In_1404);
and U4543 (N_4543,In_2352,In_1118);
xor U4544 (N_4544,In_1156,In_2115);
and U4545 (N_4545,In_107,In_2229);
nand U4546 (N_4546,In_2109,In_1327);
or U4547 (N_4547,In_1192,In_1253);
xor U4548 (N_4548,In_2202,In_1091);
nand U4549 (N_4549,In_2492,In_1272);
nor U4550 (N_4550,In_902,In_255);
xor U4551 (N_4551,In_2354,In_1032);
xor U4552 (N_4552,In_518,In_1665);
nor U4553 (N_4553,In_1420,In_1027);
or U4554 (N_4554,In_1469,In_2138);
nand U4555 (N_4555,In_404,In_27);
nand U4556 (N_4556,In_883,In_798);
nand U4557 (N_4557,In_257,In_370);
and U4558 (N_4558,In_1784,In_368);
nor U4559 (N_4559,In_2363,In_69);
and U4560 (N_4560,In_354,In_669);
and U4561 (N_4561,In_216,In_91);
xnor U4562 (N_4562,In_1245,In_2174);
or U4563 (N_4563,In_923,In_2274);
xor U4564 (N_4564,In_275,In_821);
nand U4565 (N_4565,In_2412,In_215);
nor U4566 (N_4566,In_938,In_2033);
xor U4567 (N_4567,In_1309,In_1496);
xor U4568 (N_4568,In_2177,In_68);
nand U4569 (N_4569,In_580,In_1859);
nand U4570 (N_4570,In_167,In_1308);
or U4571 (N_4571,In_807,In_904);
xor U4572 (N_4572,In_65,In_2460);
or U4573 (N_4573,In_928,In_2347);
nor U4574 (N_4574,In_166,In_314);
nand U4575 (N_4575,In_2215,In_1674);
nor U4576 (N_4576,In_1789,In_1503);
xnor U4577 (N_4577,In_1497,In_1271);
nor U4578 (N_4578,In_1510,In_2312);
nand U4579 (N_4579,In_890,In_367);
and U4580 (N_4580,In_544,In_2092);
or U4581 (N_4581,In_27,In_2356);
nand U4582 (N_4582,In_2486,In_1253);
xnor U4583 (N_4583,In_2129,In_1294);
nor U4584 (N_4584,In_309,In_1907);
xnor U4585 (N_4585,In_1177,In_18);
or U4586 (N_4586,In_1599,In_1320);
and U4587 (N_4587,In_4,In_178);
or U4588 (N_4588,In_2467,In_1142);
xor U4589 (N_4589,In_1166,In_210);
xnor U4590 (N_4590,In_1670,In_1015);
nor U4591 (N_4591,In_2193,In_646);
and U4592 (N_4592,In_574,In_1132);
nand U4593 (N_4593,In_1010,In_2073);
and U4594 (N_4594,In_1973,In_2165);
and U4595 (N_4595,In_1822,In_2109);
and U4596 (N_4596,In_1461,In_1744);
and U4597 (N_4597,In_1145,In_1826);
and U4598 (N_4598,In_2414,In_1382);
nand U4599 (N_4599,In_904,In_274);
or U4600 (N_4600,In_885,In_987);
nand U4601 (N_4601,In_115,In_878);
and U4602 (N_4602,In_1790,In_2305);
and U4603 (N_4603,In_2389,In_1484);
and U4604 (N_4604,In_1448,In_2346);
nand U4605 (N_4605,In_1003,In_2206);
and U4606 (N_4606,In_30,In_1439);
nor U4607 (N_4607,In_1073,In_2083);
or U4608 (N_4608,In_1850,In_566);
nor U4609 (N_4609,In_1977,In_2495);
nand U4610 (N_4610,In_1651,In_2440);
or U4611 (N_4611,In_2149,In_320);
nor U4612 (N_4612,In_2114,In_510);
nor U4613 (N_4613,In_892,In_1566);
nor U4614 (N_4614,In_2226,In_234);
and U4615 (N_4615,In_1188,In_1017);
nor U4616 (N_4616,In_2327,In_546);
nor U4617 (N_4617,In_754,In_412);
or U4618 (N_4618,In_2182,In_46);
nor U4619 (N_4619,In_344,In_1411);
nand U4620 (N_4620,In_2232,In_2384);
xor U4621 (N_4621,In_1272,In_2147);
and U4622 (N_4622,In_442,In_1591);
nor U4623 (N_4623,In_1617,In_903);
xnor U4624 (N_4624,In_1944,In_1261);
nand U4625 (N_4625,In_1909,In_2491);
and U4626 (N_4626,In_2482,In_1145);
and U4627 (N_4627,In_2011,In_2428);
or U4628 (N_4628,In_171,In_1380);
or U4629 (N_4629,In_1197,In_1039);
and U4630 (N_4630,In_1209,In_2053);
or U4631 (N_4631,In_677,In_2081);
xor U4632 (N_4632,In_777,In_715);
nand U4633 (N_4633,In_1063,In_1431);
and U4634 (N_4634,In_148,In_1599);
or U4635 (N_4635,In_1565,In_1475);
nor U4636 (N_4636,In_1409,In_1186);
and U4637 (N_4637,In_1707,In_1366);
or U4638 (N_4638,In_230,In_633);
nand U4639 (N_4639,In_2462,In_817);
nand U4640 (N_4640,In_1943,In_2076);
nor U4641 (N_4641,In_2283,In_355);
nor U4642 (N_4642,In_1997,In_36);
or U4643 (N_4643,In_944,In_1542);
nor U4644 (N_4644,In_1462,In_2259);
nand U4645 (N_4645,In_43,In_144);
nand U4646 (N_4646,In_861,In_1081);
or U4647 (N_4647,In_215,In_892);
and U4648 (N_4648,In_1040,In_2470);
nand U4649 (N_4649,In_121,In_748);
nand U4650 (N_4650,In_1328,In_1853);
or U4651 (N_4651,In_387,In_1660);
or U4652 (N_4652,In_842,In_671);
and U4653 (N_4653,In_1787,In_2498);
nand U4654 (N_4654,In_55,In_1695);
nor U4655 (N_4655,In_579,In_639);
nor U4656 (N_4656,In_1216,In_861);
or U4657 (N_4657,In_1608,In_2215);
nor U4658 (N_4658,In_664,In_894);
or U4659 (N_4659,In_969,In_1377);
xnor U4660 (N_4660,In_1801,In_554);
nand U4661 (N_4661,In_2382,In_1125);
xnor U4662 (N_4662,In_2267,In_1358);
xnor U4663 (N_4663,In_711,In_552);
and U4664 (N_4664,In_2396,In_2449);
xor U4665 (N_4665,In_1858,In_2305);
or U4666 (N_4666,In_159,In_2172);
and U4667 (N_4667,In_886,In_2187);
nand U4668 (N_4668,In_773,In_1002);
nor U4669 (N_4669,In_431,In_596);
and U4670 (N_4670,In_2094,In_1532);
or U4671 (N_4671,In_1226,In_680);
nor U4672 (N_4672,In_641,In_349);
nand U4673 (N_4673,In_1722,In_2196);
or U4674 (N_4674,In_65,In_2481);
nor U4675 (N_4675,In_97,In_2097);
nor U4676 (N_4676,In_1794,In_547);
and U4677 (N_4677,In_161,In_734);
or U4678 (N_4678,In_75,In_1367);
or U4679 (N_4679,In_699,In_1027);
or U4680 (N_4680,In_1161,In_1188);
nor U4681 (N_4681,In_1213,In_692);
xor U4682 (N_4682,In_19,In_646);
or U4683 (N_4683,In_1169,In_2303);
xor U4684 (N_4684,In_1617,In_340);
nor U4685 (N_4685,In_2465,In_1145);
xnor U4686 (N_4686,In_2226,In_362);
nand U4687 (N_4687,In_1211,In_1178);
nor U4688 (N_4688,In_556,In_128);
xor U4689 (N_4689,In_738,In_367);
and U4690 (N_4690,In_541,In_2386);
and U4691 (N_4691,In_1239,In_958);
xnor U4692 (N_4692,In_1279,In_2181);
nand U4693 (N_4693,In_223,In_1077);
xor U4694 (N_4694,In_2159,In_461);
or U4695 (N_4695,In_1152,In_1151);
nor U4696 (N_4696,In_865,In_79);
or U4697 (N_4697,In_1753,In_476);
nor U4698 (N_4698,In_633,In_144);
nor U4699 (N_4699,In_1731,In_290);
nand U4700 (N_4700,In_2236,In_1414);
nand U4701 (N_4701,In_1663,In_1941);
nor U4702 (N_4702,In_1791,In_1731);
and U4703 (N_4703,In_564,In_867);
or U4704 (N_4704,In_2212,In_1848);
nor U4705 (N_4705,In_1776,In_953);
xor U4706 (N_4706,In_2165,In_2492);
and U4707 (N_4707,In_204,In_987);
nor U4708 (N_4708,In_1116,In_1906);
nand U4709 (N_4709,In_1199,In_1168);
and U4710 (N_4710,In_39,In_1380);
nand U4711 (N_4711,In_821,In_1129);
nand U4712 (N_4712,In_1650,In_1462);
or U4713 (N_4713,In_1777,In_900);
nor U4714 (N_4714,In_415,In_995);
nor U4715 (N_4715,In_2080,In_904);
xnor U4716 (N_4716,In_2324,In_1079);
nor U4717 (N_4717,In_1076,In_2050);
xnor U4718 (N_4718,In_1553,In_283);
and U4719 (N_4719,In_1329,In_2051);
xnor U4720 (N_4720,In_571,In_1842);
nor U4721 (N_4721,In_2472,In_2313);
or U4722 (N_4722,In_1235,In_1222);
xor U4723 (N_4723,In_2039,In_1288);
nor U4724 (N_4724,In_430,In_1021);
or U4725 (N_4725,In_1765,In_1891);
and U4726 (N_4726,In_1987,In_1836);
and U4727 (N_4727,In_906,In_1239);
and U4728 (N_4728,In_195,In_1348);
xor U4729 (N_4729,In_1519,In_1624);
and U4730 (N_4730,In_1586,In_403);
and U4731 (N_4731,In_2424,In_929);
nor U4732 (N_4732,In_606,In_844);
xnor U4733 (N_4733,In_226,In_426);
and U4734 (N_4734,In_1962,In_326);
nor U4735 (N_4735,In_1378,In_543);
or U4736 (N_4736,In_2245,In_430);
nand U4737 (N_4737,In_1925,In_844);
nor U4738 (N_4738,In_1581,In_1646);
or U4739 (N_4739,In_189,In_589);
nand U4740 (N_4740,In_1912,In_1609);
and U4741 (N_4741,In_2133,In_1158);
or U4742 (N_4742,In_1882,In_2133);
nor U4743 (N_4743,In_999,In_1488);
and U4744 (N_4744,In_1643,In_2385);
or U4745 (N_4745,In_65,In_1775);
and U4746 (N_4746,In_2370,In_1871);
and U4747 (N_4747,In_1010,In_1906);
nor U4748 (N_4748,In_432,In_2227);
xnor U4749 (N_4749,In_1900,In_1818);
xor U4750 (N_4750,In_1738,In_1159);
nor U4751 (N_4751,In_2314,In_479);
and U4752 (N_4752,In_2110,In_457);
and U4753 (N_4753,In_1025,In_163);
xor U4754 (N_4754,In_1919,In_854);
and U4755 (N_4755,In_1789,In_199);
nand U4756 (N_4756,In_1456,In_537);
nor U4757 (N_4757,In_147,In_149);
nand U4758 (N_4758,In_778,In_2311);
nor U4759 (N_4759,In_1292,In_174);
nand U4760 (N_4760,In_836,In_1454);
xnor U4761 (N_4761,In_1443,In_1287);
xnor U4762 (N_4762,In_893,In_811);
or U4763 (N_4763,In_783,In_1979);
nor U4764 (N_4764,In_906,In_212);
xnor U4765 (N_4765,In_79,In_2378);
and U4766 (N_4766,In_1289,In_101);
nor U4767 (N_4767,In_1526,In_1988);
xor U4768 (N_4768,In_756,In_886);
and U4769 (N_4769,In_42,In_378);
nand U4770 (N_4770,In_795,In_517);
xor U4771 (N_4771,In_961,In_1341);
nand U4772 (N_4772,In_1564,In_298);
nand U4773 (N_4773,In_508,In_586);
nor U4774 (N_4774,In_2310,In_1848);
or U4775 (N_4775,In_1230,In_596);
xnor U4776 (N_4776,In_752,In_2034);
nand U4777 (N_4777,In_1068,In_684);
or U4778 (N_4778,In_1186,In_1925);
nand U4779 (N_4779,In_1470,In_2424);
and U4780 (N_4780,In_2011,In_984);
xnor U4781 (N_4781,In_1897,In_2270);
and U4782 (N_4782,In_130,In_27);
nor U4783 (N_4783,In_981,In_886);
nor U4784 (N_4784,In_682,In_794);
xor U4785 (N_4785,In_2306,In_2094);
nand U4786 (N_4786,In_2376,In_1134);
xor U4787 (N_4787,In_2499,In_1322);
nand U4788 (N_4788,In_445,In_654);
or U4789 (N_4789,In_2451,In_1666);
nand U4790 (N_4790,In_1834,In_605);
and U4791 (N_4791,In_63,In_1388);
or U4792 (N_4792,In_580,In_1316);
nor U4793 (N_4793,In_1536,In_482);
or U4794 (N_4794,In_400,In_161);
nor U4795 (N_4795,In_624,In_68);
and U4796 (N_4796,In_403,In_1822);
nor U4797 (N_4797,In_1475,In_2075);
and U4798 (N_4798,In_510,In_288);
xnor U4799 (N_4799,In_2142,In_120);
and U4800 (N_4800,In_886,In_622);
or U4801 (N_4801,In_891,In_700);
xor U4802 (N_4802,In_1968,In_6);
and U4803 (N_4803,In_1375,In_2351);
and U4804 (N_4804,In_1341,In_1255);
or U4805 (N_4805,In_818,In_1956);
nor U4806 (N_4806,In_64,In_214);
and U4807 (N_4807,In_1017,In_2410);
and U4808 (N_4808,In_450,In_1940);
nand U4809 (N_4809,In_1308,In_2271);
nor U4810 (N_4810,In_2491,In_2419);
nor U4811 (N_4811,In_1291,In_1860);
xor U4812 (N_4812,In_1335,In_1943);
and U4813 (N_4813,In_195,In_1715);
nor U4814 (N_4814,In_1106,In_2461);
and U4815 (N_4815,In_1637,In_1323);
and U4816 (N_4816,In_2393,In_1409);
nand U4817 (N_4817,In_1421,In_1162);
or U4818 (N_4818,In_2396,In_2085);
and U4819 (N_4819,In_1772,In_1054);
nor U4820 (N_4820,In_1713,In_1625);
nand U4821 (N_4821,In_806,In_2496);
nand U4822 (N_4822,In_21,In_626);
nor U4823 (N_4823,In_2323,In_2108);
and U4824 (N_4824,In_2254,In_1545);
nor U4825 (N_4825,In_1075,In_1646);
or U4826 (N_4826,In_1384,In_910);
and U4827 (N_4827,In_2309,In_799);
nand U4828 (N_4828,In_938,In_967);
and U4829 (N_4829,In_1400,In_692);
xnor U4830 (N_4830,In_1284,In_802);
xor U4831 (N_4831,In_1121,In_952);
nand U4832 (N_4832,In_1279,In_2451);
and U4833 (N_4833,In_1772,In_1055);
and U4834 (N_4834,In_2302,In_2244);
nand U4835 (N_4835,In_1348,In_480);
nor U4836 (N_4836,In_1572,In_318);
or U4837 (N_4837,In_1827,In_1315);
nor U4838 (N_4838,In_734,In_804);
xor U4839 (N_4839,In_489,In_1917);
xor U4840 (N_4840,In_80,In_665);
nor U4841 (N_4841,In_817,In_994);
or U4842 (N_4842,In_921,In_2206);
nand U4843 (N_4843,In_1807,In_353);
and U4844 (N_4844,In_1407,In_2023);
nor U4845 (N_4845,In_638,In_2064);
or U4846 (N_4846,In_552,In_327);
or U4847 (N_4847,In_2009,In_638);
xnor U4848 (N_4848,In_75,In_369);
and U4849 (N_4849,In_1565,In_365);
xor U4850 (N_4850,In_152,In_1084);
xnor U4851 (N_4851,In_1992,In_361);
xor U4852 (N_4852,In_110,In_1790);
xnor U4853 (N_4853,In_509,In_727);
xnor U4854 (N_4854,In_1469,In_2457);
and U4855 (N_4855,In_943,In_498);
nand U4856 (N_4856,In_2169,In_714);
or U4857 (N_4857,In_2168,In_2233);
or U4858 (N_4858,In_2404,In_402);
nor U4859 (N_4859,In_1441,In_881);
xnor U4860 (N_4860,In_1980,In_1925);
and U4861 (N_4861,In_1370,In_2214);
xor U4862 (N_4862,In_1840,In_430);
or U4863 (N_4863,In_239,In_2042);
nand U4864 (N_4864,In_931,In_992);
and U4865 (N_4865,In_570,In_2449);
xor U4866 (N_4866,In_572,In_2231);
and U4867 (N_4867,In_878,In_2240);
or U4868 (N_4868,In_1591,In_347);
nor U4869 (N_4869,In_984,In_291);
xor U4870 (N_4870,In_1429,In_624);
xor U4871 (N_4871,In_2340,In_267);
nor U4872 (N_4872,In_1108,In_2396);
or U4873 (N_4873,In_950,In_482);
nand U4874 (N_4874,In_1031,In_1852);
and U4875 (N_4875,In_2133,In_1736);
nor U4876 (N_4876,In_126,In_609);
xnor U4877 (N_4877,In_2145,In_1776);
and U4878 (N_4878,In_1680,In_1856);
xor U4879 (N_4879,In_177,In_2122);
and U4880 (N_4880,In_1685,In_362);
or U4881 (N_4881,In_1329,In_1906);
or U4882 (N_4882,In_1916,In_1117);
nor U4883 (N_4883,In_2333,In_851);
and U4884 (N_4884,In_1735,In_1354);
or U4885 (N_4885,In_1880,In_1788);
and U4886 (N_4886,In_1179,In_1596);
and U4887 (N_4887,In_287,In_1758);
and U4888 (N_4888,In_774,In_2489);
xnor U4889 (N_4889,In_2054,In_493);
or U4890 (N_4890,In_1902,In_340);
nor U4891 (N_4891,In_1469,In_579);
nand U4892 (N_4892,In_695,In_121);
nor U4893 (N_4893,In_1576,In_1443);
xnor U4894 (N_4894,In_1347,In_500);
or U4895 (N_4895,In_1484,In_1903);
and U4896 (N_4896,In_1778,In_1622);
and U4897 (N_4897,In_2314,In_373);
nand U4898 (N_4898,In_1911,In_1959);
or U4899 (N_4899,In_1356,In_1270);
or U4900 (N_4900,In_2201,In_1054);
and U4901 (N_4901,In_1323,In_2492);
and U4902 (N_4902,In_2366,In_694);
or U4903 (N_4903,In_1846,In_2295);
xor U4904 (N_4904,In_2266,In_248);
and U4905 (N_4905,In_1515,In_273);
and U4906 (N_4906,In_30,In_824);
nor U4907 (N_4907,In_87,In_822);
nor U4908 (N_4908,In_488,In_1714);
nor U4909 (N_4909,In_2317,In_1553);
nor U4910 (N_4910,In_2105,In_138);
xnor U4911 (N_4911,In_900,In_239);
and U4912 (N_4912,In_1354,In_2226);
and U4913 (N_4913,In_1563,In_2391);
xnor U4914 (N_4914,In_1729,In_394);
xor U4915 (N_4915,In_684,In_1620);
or U4916 (N_4916,In_844,In_341);
nand U4917 (N_4917,In_328,In_1478);
nor U4918 (N_4918,In_1195,In_2203);
or U4919 (N_4919,In_989,In_235);
or U4920 (N_4920,In_1141,In_31);
and U4921 (N_4921,In_10,In_111);
or U4922 (N_4922,In_670,In_1731);
and U4923 (N_4923,In_468,In_2377);
nor U4924 (N_4924,In_2335,In_780);
xor U4925 (N_4925,In_179,In_2094);
xnor U4926 (N_4926,In_1086,In_502);
nor U4927 (N_4927,In_1305,In_147);
or U4928 (N_4928,In_1608,In_751);
and U4929 (N_4929,In_1903,In_2416);
nor U4930 (N_4930,In_1832,In_721);
nor U4931 (N_4931,In_1543,In_73);
and U4932 (N_4932,In_800,In_2131);
nor U4933 (N_4933,In_2110,In_2452);
or U4934 (N_4934,In_1721,In_1004);
and U4935 (N_4935,In_828,In_691);
nor U4936 (N_4936,In_1393,In_253);
nor U4937 (N_4937,In_969,In_2022);
xnor U4938 (N_4938,In_2489,In_2184);
or U4939 (N_4939,In_936,In_2020);
and U4940 (N_4940,In_2407,In_1869);
nor U4941 (N_4941,In_1182,In_285);
nand U4942 (N_4942,In_1974,In_398);
xor U4943 (N_4943,In_1969,In_2261);
nand U4944 (N_4944,In_743,In_2168);
xnor U4945 (N_4945,In_1417,In_2449);
or U4946 (N_4946,In_138,In_42);
nor U4947 (N_4947,In_1504,In_1255);
xnor U4948 (N_4948,In_190,In_1424);
or U4949 (N_4949,In_1883,In_1331);
nand U4950 (N_4950,In_2205,In_532);
and U4951 (N_4951,In_2217,In_1276);
and U4952 (N_4952,In_1247,In_1866);
xor U4953 (N_4953,In_1490,In_366);
nor U4954 (N_4954,In_1420,In_168);
or U4955 (N_4955,In_2251,In_1232);
nand U4956 (N_4956,In_1032,In_366);
xor U4957 (N_4957,In_1467,In_1301);
or U4958 (N_4958,In_2208,In_1080);
nor U4959 (N_4959,In_1730,In_320);
nor U4960 (N_4960,In_2253,In_2081);
nor U4961 (N_4961,In_137,In_735);
and U4962 (N_4962,In_1330,In_1425);
nand U4963 (N_4963,In_904,In_442);
xnor U4964 (N_4964,In_1990,In_542);
nand U4965 (N_4965,In_786,In_1255);
nor U4966 (N_4966,In_2027,In_1882);
xor U4967 (N_4967,In_543,In_36);
or U4968 (N_4968,In_1728,In_2471);
nand U4969 (N_4969,In_549,In_1867);
and U4970 (N_4970,In_2109,In_492);
xnor U4971 (N_4971,In_1188,In_2238);
and U4972 (N_4972,In_66,In_2319);
or U4973 (N_4973,In_422,In_1539);
and U4974 (N_4974,In_51,In_1556);
and U4975 (N_4975,In_1738,In_1613);
nor U4976 (N_4976,In_770,In_433);
or U4977 (N_4977,In_1860,In_2177);
nor U4978 (N_4978,In_1994,In_279);
nand U4979 (N_4979,In_2099,In_1291);
and U4980 (N_4980,In_42,In_2313);
nand U4981 (N_4981,In_1101,In_1785);
or U4982 (N_4982,In_1782,In_2108);
xor U4983 (N_4983,In_1687,In_1596);
nand U4984 (N_4984,In_1468,In_642);
nor U4985 (N_4985,In_1188,In_1064);
xnor U4986 (N_4986,In_1409,In_2344);
nand U4987 (N_4987,In_2231,In_95);
nand U4988 (N_4988,In_1642,In_893);
xnor U4989 (N_4989,In_63,In_1886);
nor U4990 (N_4990,In_2362,In_2474);
and U4991 (N_4991,In_1741,In_1462);
or U4992 (N_4992,In_2470,In_234);
nor U4993 (N_4993,In_488,In_1519);
nor U4994 (N_4994,In_2215,In_828);
or U4995 (N_4995,In_2222,In_224);
xnor U4996 (N_4996,In_1477,In_2051);
nor U4997 (N_4997,In_243,In_279);
xnor U4998 (N_4998,In_625,In_1395);
nor U4999 (N_4999,In_2381,In_1895);
and U5000 (N_5000,In_167,In_1692);
nand U5001 (N_5001,In_2482,In_1964);
nand U5002 (N_5002,In_424,In_1136);
and U5003 (N_5003,In_819,In_69);
or U5004 (N_5004,In_739,In_719);
nand U5005 (N_5005,In_368,In_1817);
xor U5006 (N_5006,In_178,In_1767);
nand U5007 (N_5007,In_2043,In_1380);
or U5008 (N_5008,In_1395,In_312);
or U5009 (N_5009,In_2404,In_154);
xnor U5010 (N_5010,In_1157,In_979);
xnor U5011 (N_5011,In_159,In_2130);
or U5012 (N_5012,In_929,In_186);
and U5013 (N_5013,In_1927,In_799);
and U5014 (N_5014,In_1761,In_1081);
nor U5015 (N_5015,In_2354,In_1188);
nor U5016 (N_5016,In_1100,In_1219);
and U5017 (N_5017,In_954,In_1105);
nor U5018 (N_5018,In_1098,In_409);
nand U5019 (N_5019,In_1819,In_539);
nand U5020 (N_5020,In_2251,In_1476);
nor U5021 (N_5021,In_1351,In_755);
nand U5022 (N_5022,In_212,In_1099);
or U5023 (N_5023,In_1771,In_606);
xnor U5024 (N_5024,In_983,In_1300);
or U5025 (N_5025,In_401,In_1982);
nand U5026 (N_5026,In_13,In_1411);
or U5027 (N_5027,In_473,In_1093);
or U5028 (N_5028,In_62,In_15);
and U5029 (N_5029,In_1929,In_1935);
or U5030 (N_5030,In_690,In_450);
nor U5031 (N_5031,In_988,In_1942);
or U5032 (N_5032,In_966,In_489);
nor U5033 (N_5033,In_83,In_2334);
and U5034 (N_5034,In_102,In_1754);
or U5035 (N_5035,In_1817,In_215);
and U5036 (N_5036,In_1078,In_2023);
xor U5037 (N_5037,In_2202,In_1199);
nor U5038 (N_5038,In_2433,In_370);
or U5039 (N_5039,In_912,In_520);
xnor U5040 (N_5040,In_1123,In_1669);
nor U5041 (N_5041,In_1039,In_762);
xor U5042 (N_5042,In_513,In_491);
nor U5043 (N_5043,In_2179,In_829);
nor U5044 (N_5044,In_2447,In_820);
xnor U5045 (N_5045,In_0,In_877);
nand U5046 (N_5046,In_1222,In_477);
nor U5047 (N_5047,In_202,In_610);
xnor U5048 (N_5048,In_1123,In_1076);
and U5049 (N_5049,In_510,In_2213);
or U5050 (N_5050,In_2360,In_1285);
and U5051 (N_5051,In_2054,In_1047);
xor U5052 (N_5052,In_1369,In_1221);
or U5053 (N_5053,In_755,In_1561);
or U5054 (N_5054,In_2273,In_374);
nor U5055 (N_5055,In_1667,In_2368);
or U5056 (N_5056,In_1744,In_1812);
or U5057 (N_5057,In_1881,In_359);
and U5058 (N_5058,In_1674,In_16);
xnor U5059 (N_5059,In_2104,In_186);
xor U5060 (N_5060,In_336,In_1413);
nor U5061 (N_5061,In_1202,In_1443);
xor U5062 (N_5062,In_1724,In_334);
nor U5063 (N_5063,In_719,In_885);
nor U5064 (N_5064,In_893,In_707);
nor U5065 (N_5065,In_19,In_1640);
and U5066 (N_5066,In_1616,In_2372);
and U5067 (N_5067,In_1202,In_1130);
nand U5068 (N_5068,In_120,In_1568);
xnor U5069 (N_5069,In_1233,In_1200);
and U5070 (N_5070,In_1914,In_1245);
nand U5071 (N_5071,In_2045,In_2457);
nor U5072 (N_5072,In_12,In_617);
nor U5073 (N_5073,In_1675,In_246);
nand U5074 (N_5074,In_1048,In_2012);
or U5075 (N_5075,In_151,In_1408);
or U5076 (N_5076,In_2071,In_251);
nand U5077 (N_5077,In_284,In_1262);
or U5078 (N_5078,In_1509,In_1593);
and U5079 (N_5079,In_625,In_657);
and U5080 (N_5080,In_1303,In_451);
xor U5081 (N_5081,In_1006,In_576);
nand U5082 (N_5082,In_122,In_2492);
nor U5083 (N_5083,In_1432,In_348);
or U5084 (N_5084,In_1272,In_1069);
xor U5085 (N_5085,In_2097,In_479);
and U5086 (N_5086,In_841,In_1634);
or U5087 (N_5087,In_1691,In_1370);
nand U5088 (N_5088,In_1635,In_1719);
xnor U5089 (N_5089,In_243,In_810);
xor U5090 (N_5090,In_2140,In_1395);
or U5091 (N_5091,In_58,In_321);
nand U5092 (N_5092,In_1789,In_2357);
and U5093 (N_5093,In_2012,In_174);
and U5094 (N_5094,In_2164,In_2484);
and U5095 (N_5095,In_12,In_2125);
and U5096 (N_5096,In_919,In_640);
and U5097 (N_5097,In_1474,In_1312);
nand U5098 (N_5098,In_629,In_1142);
or U5099 (N_5099,In_1875,In_581);
nand U5100 (N_5100,In_1047,In_1492);
nor U5101 (N_5101,In_434,In_1285);
nand U5102 (N_5102,In_372,In_37);
and U5103 (N_5103,In_2359,In_1367);
xnor U5104 (N_5104,In_1877,In_377);
and U5105 (N_5105,In_793,In_1128);
or U5106 (N_5106,In_1110,In_1399);
xor U5107 (N_5107,In_256,In_2002);
nand U5108 (N_5108,In_2236,In_987);
nand U5109 (N_5109,In_1064,In_601);
xnor U5110 (N_5110,In_1125,In_1845);
and U5111 (N_5111,In_1875,In_150);
and U5112 (N_5112,In_379,In_1008);
nor U5113 (N_5113,In_1559,In_331);
nor U5114 (N_5114,In_1894,In_1236);
nand U5115 (N_5115,In_685,In_2218);
xor U5116 (N_5116,In_1060,In_1534);
or U5117 (N_5117,In_484,In_802);
or U5118 (N_5118,In_813,In_797);
xor U5119 (N_5119,In_941,In_1798);
or U5120 (N_5120,In_1386,In_1509);
nand U5121 (N_5121,In_48,In_884);
xnor U5122 (N_5122,In_2164,In_879);
nor U5123 (N_5123,In_2077,In_678);
nand U5124 (N_5124,In_1938,In_743);
or U5125 (N_5125,In_1953,In_1670);
and U5126 (N_5126,In_1001,In_1520);
and U5127 (N_5127,In_41,In_1962);
or U5128 (N_5128,In_947,In_775);
nor U5129 (N_5129,In_1767,In_1619);
nor U5130 (N_5130,In_1160,In_1035);
nor U5131 (N_5131,In_1828,In_647);
nor U5132 (N_5132,In_1118,In_160);
nand U5133 (N_5133,In_347,In_1139);
xnor U5134 (N_5134,In_184,In_1117);
xnor U5135 (N_5135,In_1626,In_560);
and U5136 (N_5136,In_1206,In_1459);
nor U5137 (N_5137,In_1944,In_796);
and U5138 (N_5138,In_92,In_1666);
and U5139 (N_5139,In_56,In_1550);
nor U5140 (N_5140,In_891,In_1969);
or U5141 (N_5141,In_2342,In_2221);
nand U5142 (N_5142,In_662,In_226);
or U5143 (N_5143,In_1624,In_1513);
nor U5144 (N_5144,In_2052,In_468);
and U5145 (N_5145,In_339,In_2038);
nor U5146 (N_5146,In_1968,In_2278);
and U5147 (N_5147,In_996,In_1858);
and U5148 (N_5148,In_509,In_1847);
and U5149 (N_5149,In_255,In_1087);
or U5150 (N_5150,In_1733,In_2037);
nor U5151 (N_5151,In_1312,In_2442);
nor U5152 (N_5152,In_1265,In_791);
xor U5153 (N_5153,In_2086,In_370);
and U5154 (N_5154,In_767,In_111);
nand U5155 (N_5155,In_1694,In_990);
or U5156 (N_5156,In_2123,In_1510);
nand U5157 (N_5157,In_980,In_2164);
xor U5158 (N_5158,In_1267,In_1633);
xor U5159 (N_5159,In_942,In_675);
and U5160 (N_5160,In_1396,In_18);
nor U5161 (N_5161,In_1521,In_2310);
xnor U5162 (N_5162,In_1249,In_1517);
xnor U5163 (N_5163,In_690,In_371);
and U5164 (N_5164,In_1650,In_2079);
and U5165 (N_5165,In_2293,In_1423);
nor U5166 (N_5166,In_1227,In_438);
or U5167 (N_5167,In_1681,In_845);
and U5168 (N_5168,In_897,In_846);
and U5169 (N_5169,In_645,In_1582);
and U5170 (N_5170,In_283,In_1625);
or U5171 (N_5171,In_2498,In_2475);
nor U5172 (N_5172,In_729,In_1875);
nand U5173 (N_5173,In_2396,In_2042);
nand U5174 (N_5174,In_952,In_1202);
xor U5175 (N_5175,In_17,In_2);
and U5176 (N_5176,In_1417,In_1447);
nor U5177 (N_5177,In_1789,In_1803);
or U5178 (N_5178,In_2413,In_1417);
nor U5179 (N_5179,In_1103,In_1273);
xor U5180 (N_5180,In_716,In_2146);
and U5181 (N_5181,In_2255,In_2043);
or U5182 (N_5182,In_2216,In_342);
xor U5183 (N_5183,In_1741,In_1598);
xor U5184 (N_5184,In_1245,In_1633);
nand U5185 (N_5185,In_2109,In_489);
and U5186 (N_5186,In_2129,In_589);
nand U5187 (N_5187,In_1843,In_1143);
xor U5188 (N_5188,In_838,In_1013);
nor U5189 (N_5189,In_2271,In_208);
nor U5190 (N_5190,In_1164,In_2131);
xor U5191 (N_5191,In_993,In_2454);
nor U5192 (N_5192,In_2373,In_2375);
nor U5193 (N_5193,In_1443,In_741);
xnor U5194 (N_5194,In_1521,In_935);
and U5195 (N_5195,In_660,In_2281);
and U5196 (N_5196,In_1518,In_2378);
xor U5197 (N_5197,In_692,In_397);
nor U5198 (N_5198,In_144,In_2386);
xnor U5199 (N_5199,In_879,In_1096);
nor U5200 (N_5200,In_955,In_2259);
nor U5201 (N_5201,In_921,In_1000);
xor U5202 (N_5202,In_13,In_2083);
nor U5203 (N_5203,In_120,In_1367);
nor U5204 (N_5204,In_158,In_712);
xor U5205 (N_5205,In_316,In_1938);
and U5206 (N_5206,In_1398,In_469);
or U5207 (N_5207,In_819,In_2085);
nand U5208 (N_5208,In_1906,In_2160);
or U5209 (N_5209,In_1746,In_1336);
nand U5210 (N_5210,In_1179,In_2378);
and U5211 (N_5211,In_435,In_382);
nand U5212 (N_5212,In_448,In_717);
nand U5213 (N_5213,In_1083,In_227);
xor U5214 (N_5214,In_105,In_1757);
xnor U5215 (N_5215,In_1172,In_2421);
xor U5216 (N_5216,In_60,In_2190);
nor U5217 (N_5217,In_2146,In_27);
nor U5218 (N_5218,In_2476,In_2081);
nand U5219 (N_5219,In_289,In_1386);
nor U5220 (N_5220,In_1718,In_794);
nand U5221 (N_5221,In_276,In_1234);
xnor U5222 (N_5222,In_1668,In_1660);
or U5223 (N_5223,In_418,In_79);
and U5224 (N_5224,In_2199,In_2063);
or U5225 (N_5225,In_1939,In_932);
or U5226 (N_5226,In_2480,In_2272);
or U5227 (N_5227,In_1379,In_1768);
and U5228 (N_5228,In_384,In_2023);
xnor U5229 (N_5229,In_753,In_503);
nor U5230 (N_5230,In_1703,In_81);
xnor U5231 (N_5231,In_879,In_842);
nand U5232 (N_5232,In_932,In_51);
or U5233 (N_5233,In_106,In_1038);
and U5234 (N_5234,In_2179,In_223);
nand U5235 (N_5235,In_1825,In_1963);
nor U5236 (N_5236,In_45,In_2306);
and U5237 (N_5237,In_715,In_1587);
or U5238 (N_5238,In_1274,In_779);
nand U5239 (N_5239,In_146,In_1877);
or U5240 (N_5240,In_2415,In_2086);
nor U5241 (N_5241,In_1130,In_1345);
nor U5242 (N_5242,In_2342,In_1808);
and U5243 (N_5243,In_1505,In_1864);
and U5244 (N_5244,In_721,In_1349);
xor U5245 (N_5245,In_2030,In_1186);
nand U5246 (N_5246,In_814,In_1122);
or U5247 (N_5247,In_840,In_456);
xor U5248 (N_5248,In_795,In_415);
nor U5249 (N_5249,In_2168,In_614);
nand U5250 (N_5250,In_471,In_2082);
nand U5251 (N_5251,In_2315,In_1557);
nor U5252 (N_5252,In_1601,In_1045);
xnor U5253 (N_5253,In_2000,In_2482);
xnor U5254 (N_5254,In_1093,In_524);
xor U5255 (N_5255,In_450,In_1280);
xnor U5256 (N_5256,In_1845,In_2408);
nand U5257 (N_5257,In_230,In_2306);
xor U5258 (N_5258,In_1161,In_14);
or U5259 (N_5259,In_1758,In_1016);
or U5260 (N_5260,In_2212,In_2343);
nand U5261 (N_5261,In_1850,In_446);
and U5262 (N_5262,In_1659,In_1801);
and U5263 (N_5263,In_838,In_2074);
nor U5264 (N_5264,In_1940,In_1141);
xnor U5265 (N_5265,In_1777,In_1233);
or U5266 (N_5266,In_1547,In_560);
or U5267 (N_5267,In_1023,In_1763);
and U5268 (N_5268,In_1277,In_841);
and U5269 (N_5269,In_1513,In_1366);
or U5270 (N_5270,In_2054,In_1654);
or U5271 (N_5271,In_619,In_1632);
xnor U5272 (N_5272,In_1204,In_2375);
nor U5273 (N_5273,In_1717,In_2092);
xor U5274 (N_5274,In_16,In_540);
or U5275 (N_5275,In_857,In_2421);
nor U5276 (N_5276,In_2031,In_1136);
nor U5277 (N_5277,In_1321,In_1701);
nand U5278 (N_5278,In_264,In_2068);
or U5279 (N_5279,In_483,In_1365);
or U5280 (N_5280,In_1033,In_277);
nor U5281 (N_5281,In_491,In_1652);
or U5282 (N_5282,In_574,In_76);
nor U5283 (N_5283,In_2146,In_2053);
nand U5284 (N_5284,In_1893,In_136);
nor U5285 (N_5285,In_1844,In_382);
and U5286 (N_5286,In_1497,In_524);
xnor U5287 (N_5287,In_1074,In_420);
xor U5288 (N_5288,In_293,In_461);
or U5289 (N_5289,In_1173,In_827);
nand U5290 (N_5290,In_2040,In_1631);
and U5291 (N_5291,In_665,In_1866);
nand U5292 (N_5292,In_1439,In_1711);
and U5293 (N_5293,In_536,In_2045);
and U5294 (N_5294,In_849,In_1443);
or U5295 (N_5295,In_2170,In_1410);
xor U5296 (N_5296,In_196,In_592);
and U5297 (N_5297,In_892,In_1160);
nor U5298 (N_5298,In_2011,In_1254);
or U5299 (N_5299,In_2338,In_212);
or U5300 (N_5300,In_855,In_831);
nor U5301 (N_5301,In_252,In_485);
and U5302 (N_5302,In_836,In_1105);
xnor U5303 (N_5303,In_122,In_1145);
xnor U5304 (N_5304,In_1537,In_1563);
nor U5305 (N_5305,In_474,In_1544);
nor U5306 (N_5306,In_747,In_1110);
and U5307 (N_5307,In_957,In_1743);
xor U5308 (N_5308,In_2181,In_2163);
xor U5309 (N_5309,In_238,In_2333);
nor U5310 (N_5310,In_1688,In_1282);
nor U5311 (N_5311,In_270,In_2359);
or U5312 (N_5312,In_47,In_2374);
and U5313 (N_5313,In_2342,In_336);
and U5314 (N_5314,In_489,In_397);
nor U5315 (N_5315,In_1638,In_1624);
or U5316 (N_5316,In_744,In_980);
and U5317 (N_5317,In_1032,In_1441);
and U5318 (N_5318,In_1127,In_767);
or U5319 (N_5319,In_1016,In_290);
and U5320 (N_5320,In_2343,In_1933);
or U5321 (N_5321,In_1613,In_926);
or U5322 (N_5322,In_238,In_369);
nor U5323 (N_5323,In_2320,In_1028);
or U5324 (N_5324,In_1120,In_1553);
nor U5325 (N_5325,In_79,In_567);
or U5326 (N_5326,In_1702,In_1052);
and U5327 (N_5327,In_174,In_2124);
or U5328 (N_5328,In_467,In_1796);
nor U5329 (N_5329,In_1666,In_383);
and U5330 (N_5330,In_385,In_2357);
and U5331 (N_5331,In_756,In_2189);
nor U5332 (N_5332,In_762,In_2030);
or U5333 (N_5333,In_200,In_1766);
and U5334 (N_5334,In_1572,In_1184);
xnor U5335 (N_5335,In_128,In_1762);
xor U5336 (N_5336,In_1503,In_686);
xor U5337 (N_5337,In_1454,In_2131);
nand U5338 (N_5338,In_855,In_1845);
nor U5339 (N_5339,In_1655,In_329);
or U5340 (N_5340,In_1123,In_2142);
nor U5341 (N_5341,In_1347,In_2490);
and U5342 (N_5342,In_432,In_1074);
and U5343 (N_5343,In_979,In_670);
or U5344 (N_5344,In_2159,In_337);
xor U5345 (N_5345,In_561,In_2059);
nor U5346 (N_5346,In_400,In_2025);
nor U5347 (N_5347,In_625,In_1590);
nor U5348 (N_5348,In_492,In_140);
nor U5349 (N_5349,In_1725,In_813);
or U5350 (N_5350,In_1483,In_782);
or U5351 (N_5351,In_2086,In_177);
nor U5352 (N_5352,In_1690,In_2096);
or U5353 (N_5353,In_341,In_522);
and U5354 (N_5354,In_161,In_1882);
nor U5355 (N_5355,In_1469,In_2438);
xnor U5356 (N_5356,In_2189,In_607);
and U5357 (N_5357,In_553,In_954);
nor U5358 (N_5358,In_578,In_70);
nand U5359 (N_5359,In_1943,In_1959);
nand U5360 (N_5360,In_1847,In_1580);
nand U5361 (N_5361,In_109,In_1405);
and U5362 (N_5362,In_60,In_1928);
and U5363 (N_5363,In_870,In_489);
and U5364 (N_5364,In_164,In_406);
nand U5365 (N_5365,In_615,In_1494);
nand U5366 (N_5366,In_944,In_638);
nand U5367 (N_5367,In_1212,In_1939);
nor U5368 (N_5368,In_2027,In_484);
nand U5369 (N_5369,In_1984,In_1250);
or U5370 (N_5370,In_1682,In_2133);
or U5371 (N_5371,In_853,In_589);
or U5372 (N_5372,In_1476,In_748);
and U5373 (N_5373,In_2116,In_682);
nor U5374 (N_5374,In_3,In_510);
or U5375 (N_5375,In_59,In_309);
nand U5376 (N_5376,In_2485,In_52);
nand U5377 (N_5377,In_250,In_1807);
or U5378 (N_5378,In_204,In_1643);
xor U5379 (N_5379,In_1780,In_1571);
nor U5380 (N_5380,In_904,In_1205);
xnor U5381 (N_5381,In_243,In_679);
nand U5382 (N_5382,In_606,In_1264);
nor U5383 (N_5383,In_885,In_1103);
and U5384 (N_5384,In_281,In_2484);
xnor U5385 (N_5385,In_384,In_216);
nand U5386 (N_5386,In_370,In_2475);
xnor U5387 (N_5387,In_950,In_2370);
and U5388 (N_5388,In_480,In_667);
xnor U5389 (N_5389,In_130,In_212);
nand U5390 (N_5390,In_1437,In_1243);
nand U5391 (N_5391,In_1238,In_171);
nor U5392 (N_5392,In_149,In_1628);
or U5393 (N_5393,In_371,In_1215);
or U5394 (N_5394,In_935,In_1628);
and U5395 (N_5395,In_634,In_86);
nor U5396 (N_5396,In_609,In_2045);
or U5397 (N_5397,In_1471,In_1334);
or U5398 (N_5398,In_1548,In_620);
nand U5399 (N_5399,In_488,In_15);
or U5400 (N_5400,In_318,In_1514);
xor U5401 (N_5401,In_1160,In_30);
nand U5402 (N_5402,In_2182,In_2204);
nand U5403 (N_5403,In_1358,In_1460);
nor U5404 (N_5404,In_1778,In_2381);
and U5405 (N_5405,In_1431,In_913);
nand U5406 (N_5406,In_893,In_1237);
nand U5407 (N_5407,In_1953,In_1559);
or U5408 (N_5408,In_138,In_999);
and U5409 (N_5409,In_1458,In_1603);
nor U5410 (N_5410,In_1935,In_370);
and U5411 (N_5411,In_1415,In_1371);
or U5412 (N_5412,In_1004,In_167);
xor U5413 (N_5413,In_1973,In_64);
xnor U5414 (N_5414,In_163,In_590);
nor U5415 (N_5415,In_2168,In_1631);
xor U5416 (N_5416,In_1421,In_1287);
nor U5417 (N_5417,In_378,In_1156);
nand U5418 (N_5418,In_404,In_600);
nor U5419 (N_5419,In_1706,In_1935);
xor U5420 (N_5420,In_52,In_2437);
and U5421 (N_5421,In_1594,In_2377);
and U5422 (N_5422,In_1201,In_1523);
xnor U5423 (N_5423,In_165,In_2185);
nand U5424 (N_5424,In_1968,In_2094);
nor U5425 (N_5425,In_1286,In_425);
or U5426 (N_5426,In_1509,In_436);
nor U5427 (N_5427,In_209,In_1628);
and U5428 (N_5428,In_818,In_2221);
or U5429 (N_5429,In_1054,In_1523);
xor U5430 (N_5430,In_373,In_191);
nand U5431 (N_5431,In_861,In_465);
nand U5432 (N_5432,In_1793,In_2378);
xnor U5433 (N_5433,In_70,In_1538);
and U5434 (N_5434,In_506,In_708);
nand U5435 (N_5435,In_1745,In_811);
nor U5436 (N_5436,In_2176,In_647);
and U5437 (N_5437,In_1916,In_2238);
or U5438 (N_5438,In_1342,In_569);
nand U5439 (N_5439,In_1515,In_2396);
nand U5440 (N_5440,In_2269,In_686);
nand U5441 (N_5441,In_2117,In_234);
nor U5442 (N_5442,In_335,In_2400);
xor U5443 (N_5443,In_1627,In_2275);
or U5444 (N_5444,In_357,In_349);
nor U5445 (N_5445,In_798,In_2464);
xnor U5446 (N_5446,In_2216,In_1158);
nor U5447 (N_5447,In_1420,In_658);
and U5448 (N_5448,In_2482,In_1566);
xnor U5449 (N_5449,In_2157,In_424);
or U5450 (N_5450,In_1698,In_1354);
nor U5451 (N_5451,In_1670,In_777);
nor U5452 (N_5452,In_825,In_1143);
or U5453 (N_5453,In_1728,In_1985);
or U5454 (N_5454,In_963,In_666);
nand U5455 (N_5455,In_1081,In_1468);
or U5456 (N_5456,In_2167,In_2150);
and U5457 (N_5457,In_2474,In_363);
nand U5458 (N_5458,In_2319,In_1126);
and U5459 (N_5459,In_566,In_459);
and U5460 (N_5460,In_1410,In_762);
nand U5461 (N_5461,In_78,In_994);
or U5462 (N_5462,In_2134,In_982);
and U5463 (N_5463,In_113,In_99);
nand U5464 (N_5464,In_1229,In_990);
nand U5465 (N_5465,In_489,In_540);
or U5466 (N_5466,In_2219,In_1052);
or U5467 (N_5467,In_1932,In_152);
xor U5468 (N_5468,In_1231,In_374);
xnor U5469 (N_5469,In_1685,In_1988);
or U5470 (N_5470,In_970,In_1398);
nand U5471 (N_5471,In_697,In_2037);
or U5472 (N_5472,In_2338,In_280);
nor U5473 (N_5473,In_50,In_2125);
and U5474 (N_5474,In_186,In_1333);
and U5475 (N_5475,In_1763,In_404);
or U5476 (N_5476,In_162,In_2062);
nand U5477 (N_5477,In_954,In_2106);
or U5478 (N_5478,In_1024,In_830);
or U5479 (N_5479,In_2422,In_369);
nor U5480 (N_5480,In_1482,In_1448);
xnor U5481 (N_5481,In_1514,In_2271);
nand U5482 (N_5482,In_2363,In_1849);
or U5483 (N_5483,In_763,In_2351);
or U5484 (N_5484,In_644,In_1989);
and U5485 (N_5485,In_1969,In_1998);
or U5486 (N_5486,In_2165,In_2083);
or U5487 (N_5487,In_141,In_931);
and U5488 (N_5488,In_2104,In_2209);
nor U5489 (N_5489,In_653,In_1355);
nand U5490 (N_5490,In_2137,In_1105);
nand U5491 (N_5491,In_1063,In_992);
or U5492 (N_5492,In_2344,In_1903);
nand U5493 (N_5493,In_2382,In_187);
nor U5494 (N_5494,In_1542,In_794);
and U5495 (N_5495,In_2153,In_1508);
nand U5496 (N_5496,In_2444,In_1505);
and U5497 (N_5497,In_442,In_298);
or U5498 (N_5498,In_1726,In_1331);
nand U5499 (N_5499,In_1870,In_701);
nor U5500 (N_5500,In_284,In_139);
and U5501 (N_5501,In_1885,In_542);
or U5502 (N_5502,In_620,In_1958);
and U5503 (N_5503,In_1988,In_2398);
and U5504 (N_5504,In_1478,In_363);
nor U5505 (N_5505,In_2418,In_988);
nand U5506 (N_5506,In_1804,In_1371);
and U5507 (N_5507,In_1171,In_946);
nor U5508 (N_5508,In_259,In_373);
xnor U5509 (N_5509,In_603,In_1311);
and U5510 (N_5510,In_66,In_71);
xnor U5511 (N_5511,In_1990,In_2351);
xnor U5512 (N_5512,In_1108,In_2100);
nand U5513 (N_5513,In_2260,In_2091);
and U5514 (N_5514,In_1681,In_688);
xnor U5515 (N_5515,In_167,In_520);
xor U5516 (N_5516,In_2113,In_616);
and U5517 (N_5517,In_1755,In_1174);
nand U5518 (N_5518,In_1174,In_2082);
nor U5519 (N_5519,In_938,In_940);
nor U5520 (N_5520,In_1252,In_2345);
nor U5521 (N_5521,In_2372,In_1977);
and U5522 (N_5522,In_2408,In_631);
nor U5523 (N_5523,In_1668,In_2063);
nor U5524 (N_5524,In_282,In_2421);
nand U5525 (N_5525,In_451,In_894);
or U5526 (N_5526,In_2072,In_2);
or U5527 (N_5527,In_392,In_1448);
nor U5528 (N_5528,In_2447,In_2302);
and U5529 (N_5529,In_1908,In_2322);
xor U5530 (N_5530,In_533,In_866);
and U5531 (N_5531,In_969,In_448);
nor U5532 (N_5532,In_2206,In_1480);
and U5533 (N_5533,In_2009,In_1189);
nand U5534 (N_5534,In_137,In_2465);
and U5535 (N_5535,In_968,In_1578);
nor U5536 (N_5536,In_1759,In_2249);
nand U5537 (N_5537,In_1902,In_1350);
and U5538 (N_5538,In_1493,In_1248);
nand U5539 (N_5539,In_73,In_1687);
nor U5540 (N_5540,In_822,In_635);
and U5541 (N_5541,In_1918,In_1871);
nor U5542 (N_5542,In_1128,In_133);
nor U5543 (N_5543,In_2195,In_692);
or U5544 (N_5544,In_2486,In_902);
or U5545 (N_5545,In_431,In_615);
nor U5546 (N_5546,In_63,In_718);
and U5547 (N_5547,In_1910,In_313);
or U5548 (N_5548,In_1014,In_1433);
xor U5549 (N_5549,In_267,In_1973);
nor U5550 (N_5550,In_686,In_1016);
and U5551 (N_5551,In_1873,In_1853);
or U5552 (N_5552,In_1912,In_2336);
or U5553 (N_5553,In_2115,In_1257);
and U5554 (N_5554,In_443,In_653);
nor U5555 (N_5555,In_1249,In_2168);
xnor U5556 (N_5556,In_1142,In_2254);
nor U5557 (N_5557,In_1551,In_1684);
or U5558 (N_5558,In_499,In_2056);
nor U5559 (N_5559,In_434,In_361);
xnor U5560 (N_5560,In_1701,In_2322);
and U5561 (N_5561,In_1389,In_412);
nor U5562 (N_5562,In_617,In_707);
xor U5563 (N_5563,In_492,In_1210);
nand U5564 (N_5564,In_1768,In_764);
or U5565 (N_5565,In_656,In_2268);
xor U5566 (N_5566,In_786,In_2093);
xor U5567 (N_5567,In_102,In_873);
or U5568 (N_5568,In_2284,In_854);
or U5569 (N_5569,In_2062,In_158);
xnor U5570 (N_5570,In_1844,In_1794);
or U5571 (N_5571,In_2166,In_1690);
or U5572 (N_5572,In_117,In_2011);
or U5573 (N_5573,In_1667,In_1980);
or U5574 (N_5574,In_1689,In_571);
nand U5575 (N_5575,In_1989,In_363);
xor U5576 (N_5576,In_1558,In_1971);
or U5577 (N_5577,In_585,In_1290);
nor U5578 (N_5578,In_1161,In_2479);
nor U5579 (N_5579,In_2303,In_759);
nand U5580 (N_5580,In_580,In_1581);
and U5581 (N_5581,In_2295,In_390);
nand U5582 (N_5582,In_804,In_1677);
nor U5583 (N_5583,In_956,In_1530);
nand U5584 (N_5584,In_2340,In_547);
nor U5585 (N_5585,In_1834,In_192);
or U5586 (N_5586,In_1811,In_990);
or U5587 (N_5587,In_1974,In_1715);
and U5588 (N_5588,In_695,In_200);
or U5589 (N_5589,In_2408,In_1048);
nand U5590 (N_5590,In_1035,In_1672);
xnor U5591 (N_5591,In_2153,In_962);
nand U5592 (N_5592,In_136,In_561);
nand U5593 (N_5593,In_60,In_2300);
nand U5594 (N_5594,In_1421,In_470);
nor U5595 (N_5595,In_55,In_1809);
xnor U5596 (N_5596,In_55,In_1612);
and U5597 (N_5597,In_2090,In_1511);
nor U5598 (N_5598,In_1004,In_1777);
xor U5599 (N_5599,In_99,In_1164);
and U5600 (N_5600,In_59,In_1281);
or U5601 (N_5601,In_1287,In_1769);
or U5602 (N_5602,In_64,In_982);
nand U5603 (N_5603,In_478,In_801);
or U5604 (N_5604,In_809,In_830);
nand U5605 (N_5605,In_1270,In_843);
nor U5606 (N_5606,In_1756,In_1576);
and U5607 (N_5607,In_699,In_2215);
xor U5608 (N_5608,In_575,In_227);
and U5609 (N_5609,In_491,In_7);
and U5610 (N_5610,In_1294,In_2221);
and U5611 (N_5611,In_1225,In_1459);
and U5612 (N_5612,In_844,In_1946);
or U5613 (N_5613,In_2129,In_1758);
or U5614 (N_5614,In_1080,In_1707);
or U5615 (N_5615,In_216,In_1917);
xor U5616 (N_5616,In_323,In_1780);
nor U5617 (N_5617,In_189,In_506);
nand U5618 (N_5618,In_356,In_2312);
and U5619 (N_5619,In_2269,In_326);
or U5620 (N_5620,In_1011,In_477);
or U5621 (N_5621,In_1427,In_1992);
or U5622 (N_5622,In_2130,In_917);
xor U5623 (N_5623,In_1169,In_850);
or U5624 (N_5624,In_2186,In_2286);
xor U5625 (N_5625,In_791,In_613);
xor U5626 (N_5626,In_1551,In_2097);
nor U5627 (N_5627,In_1601,In_1041);
or U5628 (N_5628,In_1502,In_406);
xor U5629 (N_5629,In_205,In_1386);
or U5630 (N_5630,In_1887,In_1405);
and U5631 (N_5631,In_540,In_557);
and U5632 (N_5632,In_1458,In_1641);
xor U5633 (N_5633,In_1856,In_166);
and U5634 (N_5634,In_2369,In_460);
xor U5635 (N_5635,In_289,In_42);
and U5636 (N_5636,In_2113,In_1954);
or U5637 (N_5637,In_352,In_749);
and U5638 (N_5638,In_1326,In_2051);
or U5639 (N_5639,In_1727,In_825);
or U5640 (N_5640,In_1721,In_1230);
xor U5641 (N_5641,In_98,In_871);
nand U5642 (N_5642,In_2439,In_328);
and U5643 (N_5643,In_839,In_1367);
xnor U5644 (N_5644,In_357,In_1120);
nor U5645 (N_5645,In_2033,In_2102);
xor U5646 (N_5646,In_1030,In_1592);
and U5647 (N_5647,In_1832,In_1240);
nand U5648 (N_5648,In_17,In_849);
nand U5649 (N_5649,In_2114,In_877);
and U5650 (N_5650,In_1699,In_1066);
and U5651 (N_5651,In_38,In_1814);
or U5652 (N_5652,In_404,In_1018);
or U5653 (N_5653,In_294,In_2371);
nand U5654 (N_5654,In_295,In_555);
nand U5655 (N_5655,In_1041,In_1132);
and U5656 (N_5656,In_716,In_158);
and U5657 (N_5657,In_2285,In_1826);
or U5658 (N_5658,In_635,In_1051);
nor U5659 (N_5659,In_277,In_1009);
and U5660 (N_5660,In_1668,In_648);
xor U5661 (N_5661,In_569,In_50);
or U5662 (N_5662,In_14,In_1546);
nor U5663 (N_5663,In_415,In_2177);
nor U5664 (N_5664,In_664,In_1184);
nand U5665 (N_5665,In_1730,In_503);
nor U5666 (N_5666,In_859,In_1064);
nand U5667 (N_5667,In_1973,In_2003);
xor U5668 (N_5668,In_2309,In_783);
xnor U5669 (N_5669,In_559,In_608);
nor U5670 (N_5670,In_1956,In_1130);
or U5671 (N_5671,In_490,In_1330);
nand U5672 (N_5672,In_433,In_527);
nand U5673 (N_5673,In_1491,In_1521);
nand U5674 (N_5674,In_683,In_1260);
nor U5675 (N_5675,In_330,In_1334);
nor U5676 (N_5676,In_1090,In_20);
and U5677 (N_5677,In_1923,In_91);
xnor U5678 (N_5678,In_2079,In_1339);
xnor U5679 (N_5679,In_1966,In_302);
or U5680 (N_5680,In_2248,In_1050);
nor U5681 (N_5681,In_1383,In_1691);
xor U5682 (N_5682,In_1311,In_1534);
and U5683 (N_5683,In_499,In_22);
nor U5684 (N_5684,In_0,In_2431);
nor U5685 (N_5685,In_515,In_187);
or U5686 (N_5686,In_795,In_2417);
or U5687 (N_5687,In_1366,In_720);
and U5688 (N_5688,In_1270,In_1292);
xnor U5689 (N_5689,In_47,In_1043);
and U5690 (N_5690,In_2068,In_2490);
nor U5691 (N_5691,In_823,In_1717);
or U5692 (N_5692,In_875,In_273);
and U5693 (N_5693,In_420,In_1421);
or U5694 (N_5694,In_2151,In_725);
nor U5695 (N_5695,In_1453,In_1218);
nor U5696 (N_5696,In_181,In_1258);
xnor U5697 (N_5697,In_2154,In_1894);
nor U5698 (N_5698,In_744,In_385);
and U5699 (N_5699,In_1620,In_282);
nor U5700 (N_5700,In_1142,In_1710);
xor U5701 (N_5701,In_2121,In_458);
and U5702 (N_5702,In_13,In_246);
or U5703 (N_5703,In_2342,In_478);
nand U5704 (N_5704,In_466,In_674);
and U5705 (N_5705,In_1002,In_1538);
or U5706 (N_5706,In_185,In_908);
xnor U5707 (N_5707,In_1722,In_2222);
nand U5708 (N_5708,In_1004,In_1997);
nor U5709 (N_5709,In_1036,In_2356);
and U5710 (N_5710,In_2106,In_1769);
and U5711 (N_5711,In_1785,In_594);
and U5712 (N_5712,In_241,In_1291);
nor U5713 (N_5713,In_228,In_2101);
nand U5714 (N_5714,In_1057,In_1319);
nor U5715 (N_5715,In_1071,In_2311);
nand U5716 (N_5716,In_1022,In_2193);
xnor U5717 (N_5717,In_5,In_1122);
and U5718 (N_5718,In_929,In_1876);
xnor U5719 (N_5719,In_158,In_497);
and U5720 (N_5720,In_501,In_277);
or U5721 (N_5721,In_2022,In_1570);
xor U5722 (N_5722,In_1358,In_2394);
or U5723 (N_5723,In_725,In_1481);
nand U5724 (N_5724,In_685,In_2374);
xor U5725 (N_5725,In_2318,In_434);
xor U5726 (N_5726,In_93,In_2019);
or U5727 (N_5727,In_2198,In_1594);
xnor U5728 (N_5728,In_1575,In_1422);
xnor U5729 (N_5729,In_536,In_312);
nor U5730 (N_5730,In_1785,In_895);
xnor U5731 (N_5731,In_2082,In_1818);
nor U5732 (N_5732,In_2401,In_370);
or U5733 (N_5733,In_1338,In_1065);
xnor U5734 (N_5734,In_2238,In_855);
nor U5735 (N_5735,In_1746,In_758);
and U5736 (N_5736,In_1910,In_923);
xor U5737 (N_5737,In_645,In_2303);
xor U5738 (N_5738,In_2221,In_727);
xor U5739 (N_5739,In_2439,In_598);
or U5740 (N_5740,In_1242,In_791);
xor U5741 (N_5741,In_646,In_529);
nor U5742 (N_5742,In_1996,In_999);
nand U5743 (N_5743,In_917,In_208);
or U5744 (N_5744,In_2430,In_2298);
xnor U5745 (N_5745,In_1612,In_1388);
nand U5746 (N_5746,In_1388,In_1307);
xnor U5747 (N_5747,In_2258,In_948);
and U5748 (N_5748,In_2406,In_1264);
nor U5749 (N_5749,In_1291,In_1910);
and U5750 (N_5750,In_1892,In_398);
and U5751 (N_5751,In_2313,In_1100);
or U5752 (N_5752,In_2283,In_465);
nor U5753 (N_5753,In_980,In_480);
nand U5754 (N_5754,In_64,In_146);
nand U5755 (N_5755,In_931,In_426);
nand U5756 (N_5756,In_1171,In_1199);
nand U5757 (N_5757,In_1480,In_116);
or U5758 (N_5758,In_671,In_1861);
xor U5759 (N_5759,In_2208,In_519);
nand U5760 (N_5760,In_720,In_2109);
xnor U5761 (N_5761,In_347,In_1128);
nand U5762 (N_5762,In_502,In_974);
xor U5763 (N_5763,In_2210,In_286);
or U5764 (N_5764,In_1509,In_2062);
nor U5765 (N_5765,In_145,In_2347);
nor U5766 (N_5766,In_1042,In_156);
and U5767 (N_5767,In_2169,In_2148);
and U5768 (N_5768,In_1582,In_2262);
and U5769 (N_5769,In_2336,In_2320);
nor U5770 (N_5770,In_2000,In_1056);
nand U5771 (N_5771,In_2114,In_1236);
nand U5772 (N_5772,In_1902,In_2031);
nor U5773 (N_5773,In_862,In_2230);
and U5774 (N_5774,In_861,In_1262);
nand U5775 (N_5775,In_2238,In_686);
nand U5776 (N_5776,In_1235,In_2312);
nor U5777 (N_5777,In_202,In_2085);
and U5778 (N_5778,In_1460,In_109);
nand U5779 (N_5779,In_2366,In_2013);
and U5780 (N_5780,In_472,In_1241);
nor U5781 (N_5781,In_337,In_2072);
or U5782 (N_5782,In_597,In_480);
nand U5783 (N_5783,In_802,In_2174);
nand U5784 (N_5784,In_313,In_2383);
and U5785 (N_5785,In_1888,In_2391);
or U5786 (N_5786,In_1611,In_393);
nand U5787 (N_5787,In_2066,In_2458);
nor U5788 (N_5788,In_1320,In_876);
or U5789 (N_5789,In_2190,In_1639);
xor U5790 (N_5790,In_1167,In_1388);
nand U5791 (N_5791,In_2112,In_997);
or U5792 (N_5792,In_949,In_1957);
xor U5793 (N_5793,In_2202,In_2346);
or U5794 (N_5794,In_76,In_715);
xor U5795 (N_5795,In_1481,In_39);
or U5796 (N_5796,In_934,In_235);
nor U5797 (N_5797,In_1366,In_1251);
nand U5798 (N_5798,In_249,In_1184);
and U5799 (N_5799,In_2314,In_883);
nor U5800 (N_5800,In_1335,In_1000);
nor U5801 (N_5801,In_2320,In_455);
xnor U5802 (N_5802,In_1039,In_950);
and U5803 (N_5803,In_1183,In_1456);
or U5804 (N_5804,In_286,In_469);
and U5805 (N_5805,In_1804,In_2475);
and U5806 (N_5806,In_1102,In_2363);
nand U5807 (N_5807,In_1053,In_1302);
and U5808 (N_5808,In_838,In_2359);
xor U5809 (N_5809,In_2104,In_2348);
or U5810 (N_5810,In_921,In_1323);
nand U5811 (N_5811,In_1332,In_786);
nand U5812 (N_5812,In_1214,In_1827);
and U5813 (N_5813,In_1751,In_2121);
nand U5814 (N_5814,In_1765,In_1802);
xor U5815 (N_5815,In_36,In_715);
and U5816 (N_5816,In_1681,In_1543);
nor U5817 (N_5817,In_329,In_986);
and U5818 (N_5818,In_1367,In_292);
and U5819 (N_5819,In_1661,In_1601);
and U5820 (N_5820,In_939,In_2392);
xor U5821 (N_5821,In_850,In_909);
xor U5822 (N_5822,In_1086,In_831);
and U5823 (N_5823,In_45,In_1892);
nor U5824 (N_5824,In_2143,In_571);
nand U5825 (N_5825,In_123,In_622);
and U5826 (N_5826,In_1050,In_712);
and U5827 (N_5827,In_178,In_496);
and U5828 (N_5828,In_974,In_900);
xor U5829 (N_5829,In_1827,In_1512);
nand U5830 (N_5830,In_242,In_1006);
or U5831 (N_5831,In_2167,In_1474);
nand U5832 (N_5832,In_1742,In_790);
and U5833 (N_5833,In_395,In_2315);
nor U5834 (N_5834,In_1278,In_2350);
and U5835 (N_5835,In_869,In_1246);
xor U5836 (N_5836,In_2449,In_1854);
and U5837 (N_5837,In_2077,In_314);
nor U5838 (N_5838,In_486,In_2196);
and U5839 (N_5839,In_21,In_2420);
nor U5840 (N_5840,In_363,In_1698);
and U5841 (N_5841,In_1523,In_1792);
nand U5842 (N_5842,In_605,In_505);
or U5843 (N_5843,In_2146,In_2084);
or U5844 (N_5844,In_1096,In_735);
or U5845 (N_5845,In_1292,In_973);
nor U5846 (N_5846,In_1872,In_668);
nor U5847 (N_5847,In_60,In_1918);
nand U5848 (N_5848,In_2056,In_143);
and U5849 (N_5849,In_259,In_516);
and U5850 (N_5850,In_967,In_312);
or U5851 (N_5851,In_656,In_2310);
and U5852 (N_5852,In_1361,In_1434);
xor U5853 (N_5853,In_777,In_266);
and U5854 (N_5854,In_282,In_132);
nor U5855 (N_5855,In_912,In_2467);
nand U5856 (N_5856,In_358,In_953);
nor U5857 (N_5857,In_2039,In_889);
nor U5858 (N_5858,In_631,In_2213);
and U5859 (N_5859,In_1337,In_1801);
and U5860 (N_5860,In_77,In_816);
nand U5861 (N_5861,In_1046,In_2354);
nand U5862 (N_5862,In_1844,In_864);
or U5863 (N_5863,In_1980,In_552);
or U5864 (N_5864,In_1773,In_1214);
nor U5865 (N_5865,In_1454,In_217);
nor U5866 (N_5866,In_1135,In_1793);
and U5867 (N_5867,In_642,In_679);
and U5868 (N_5868,In_134,In_942);
or U5869 (N_5869,In_1432,In_1062);
nand U5870 (N_5870,In_1245,In_2311);
nor U5871 (N_5871,In_909,In_300);
and U5872 (N_5872,In_2101,In_1689);
or U5873 (N_5873,In_2261,In_154);
and U5874 (N_5874,In_289,In_2016);
or U5875 (N_5875,In_1926,In_1227);
and U5876 (N_5876,In_1324,In_2333);
or U5877 (N_5877,In_78,In_2365);
nor U5878 (N_5878,In_189,In_690);
nand U5879 (N_5879,In_1857,In_1326);
or U5880 (N_5880,In_271,In_551);
and U5881 (N_5881,In_577,In_1085);
xor U5882 (N_5882,In_11,In_611);
and U5883 (N_5883,In_967,In_191);
and U5884 (N_5884,In_2050,In_2342);
nor U5885 (N_5885,In_2235,In_1622);
or U5886 (N_5886,In_832,In_2061);
xnor U5887 (N_5887,In_888,In_67);
or U5888 (N_5888,In_492,In_266);
xor U5889 (N_5889,In_311,In_313);
or U5890 (N_5890,In_677,In_1279);
and U5891 (N_5891,In_2172,In_1224);
nor U5892 (N_5892,In_1556,In_1095);
and U5893 (N_5893,In_1335,In_1346);
and U5894 (N_5894,In_1211,In_1744);
or U5895 (N_5895,In_1587,In_1381);
nor U5896 (N_5896,In_1902,In_1482);
nor U5897 (N_5897,In_1262,In_312);
nor U5898 (N_5898,In_2224,In_1493);
or U5899 (N_5899,In_719,In_893);
nand U5900 (N_5900,In_2121,In_2442);
and U5901 (N_5901,In_1838,In_1824);
and U5902 (N_5902,In_793,In_1159);
or U5903 (N_5903,In_2261,In_1453);
or U5904 (N_5904,In_1878,In_73);
xor U5905 (N_5905,In_1828,In_1835);
xnor U5906 (N_5906,In_1476,In_39);
nand U5907 (N_5907,In_1386,In_1870);
xor U5908 (N_5908,In_1946,In_1713);
nor U5909 (N_5909,In_939,In_1280);
nor U5910 (N_5910,In_1604,In_731);
nand U5911 (N_5911,In_1819,In_891);
or U5912 (N_5912,In_1708,In_847);
nand U5913 (N_5913,In_1717,In_2031);
or U5914 (N_5914,In_2250,In_371);
or U5915 (N_5915,In_1770,In_1434);
nor U5916 (N_5916,In_705,In_1234);
or U5917 (N_5917,In_1967,In_905);
or U5918 (N_5918,In_2104,In_2368);
and U5919 (N_5919,In_1359,In_525);
nor U5920 (N_5920,In_2112,In_279);
nor U5921 (N_5921,In_345,In_1277);
xor U5922 (N_5922,In_563,In_2474);
nor U5923 (N_5923,In_628,In_793);
nor U5924 (N_5924,In_2148,In_1051);
or U5925 (N_5925,In_1473,In_1417);
xor U5926 (N_5926,In_1445,In_1460);
nand U5927 (N_5927,In_1935,In_1063);
nor U5928 (N_5928,In_2128,In_197);
xnor U5929 (N_5929,In_1766,In_1986);
and U5930 (N_5930,In_293,In_1604);
and U5931 (N_5931,In_800,In_1521);
nand U5932 (N_5932,In_1436,In_1930);
nor U5933 (N_5933,In_2370,In_886);
nand U5934 (N_5934,In_1812,In_1614);
nor U5935 (N_5935,In_1012,In_649);
xor U5936 (N_5936,In_775,In_1367);
xnor U5937 (N_5937,In_47,In_55);
and U5938 (N_5938,In_1553,In_2031);
xnor U5939 (N_5939,In_1746,In_768);
xnor U5940 (N_5940,In_811,In_447);
nor U5941 (N_5941,In_121,In_573);
or U5942 (N_5942,In_2079,In_20);
nor U5943 (N_5943,In_488,In_2249);
nor U5944 (N_5944,In_742,In_1369);
nand U5945 (N_5945,In_2488,In_179);
nand U5946 (N_5946,In_1407,In_714);
or U5947 (N_5947,In_2014,In_1091);
xor U5948 (N_5948,In_2222,In_15);
xnor U5949 (N_5949,In_1860,In_330);
xor U5950 (N_5950,In_1741,In_917);
xor U5951 (N_5951,In_2408,In_1813);
or U5952 (N_5952,In_157,In_765);
nand U5953 (N_5953,In_1237,In_232);
xor U5954 (N_5954,In_245,In_2026);
nand U5955 (N_5955,In_1703,In_1362);
nand U5956 (N_5956,In_2279,In_1097);
nor U5957 (N_5957,In_1908,In_1135);
nand U5958 (N_5958,In_1754,In_2273);
xnor U5959 (N_5959,In_2377,In_152);
or U5960 (N_5960,In_1340,In_1262);
or U5961 (N_5961,In_814,In_1366);
xor U5962 (N_5962,In_1976,In_2124);
nand U5963 (N_5963,In_1965,In_1895);
and U5964 (N_5964,In_864,In_1375);
or U5965 (N_5965,In_30,In_1632);
nand U5966 (N_5966,In_1159,In_56);
and U5967 (N_5967,In_379,In_983);
or U5968 (N_5968,In_1518,In_12);
nand U5969 (N_5969,In_1141,In_1735);
nor U5970 (N_5970,In_1201,In_1644);
or U5971 (N_5971,In_407,In_801);
or U5972 (N_5972,In_1518,In_732);
and U5973 (N_5973,In_1292,In_628);
nand U5974 (N_5974,In_1718,In_2198);
and U5975 (N_5975,In_421,In_1750);
nor U5976 (N_5976,In_185,In_813);
and U5977 (N_5977,In_1796,In_468);
or U5978 (N_5978,In_1071,In_358);
nand U5979 (N_5979,In_1526,In_432);
and U5980 (N_5980,In_881,In_247);
nand U5981 (N_5981,In_2287,In_120);
xnor U5982 (N_5982,In_1709,In_133);
or U5983 (N_5983,In_2022,In_28);
or U5984 (N_5984,In_240,In_167);
and U5985 (N_5985,In_1962,In_2331);
xor U5986 (N_5986,In_444,In_166);
or U5987 (N_5987,In_558,In_2401);
and U5988 (N_5988,In_2477,In_603);
nor U5989 (N_5989,In_1462,In_768);
nor U5990 (N_5990,In_1679,In_659);
nand U5991 (N_5991,In_1712,In_1820);
nor U5992 (N_5992,In_1534,In_1007);
xor U5993 (N_5993,In_2017,In_1488);
nor U5994 (N_5994,In_1867,In_1039);
xnor U5995 (N_5995,In_20,In_1852);
nor U5996 (N_5996,In_1407,In_1726);
nor U5997 (N_5997,In_702,In_2338);
xor U5998 (N_5998,In_129,In_906);
xnor U5999 (N_5999,In_1841,In_1041);
nand U6000 (N_6000,In_1695,In_871);
and U6001 (N_6001,In_290,In_1983);
xnor U6002 (N_6002,In_261,In_1544);
xor U6003 (N_6003,In_156,In_581);
xor U6004 (N_6004,In_1612,In_1160);
xnor U6005 (N_6005,In_2403,In_2289);
or U6006 (N_6006,In_1807,In_1633);
nand U6007 (N_6007,In_35,In_1082);
and U6008 (N_6008,In_1475,In_897);
xnor U6009 (N_6009,In_768,In_701);
nor U6010 (N_6010,In_1899,In_123);
nand U6011 (N_6011,In_127,In_2301);
or U6012 (N_6012,In_434,In_223);
nand U6013 (N_6013,In_880,In_2361);
nor U6014 (N_6014,In_15,In_469);
and U6015 (N_6015,In_358,In_769);
nor U6016 (N_6016,In_431,In_1625);
xor U6017 (N_6017,In_2301,In_440);
nand U6018 (N_6018,In_1034,In_778);
and U6019 (N_6019,In_179,In_2278);
and U6020 (N_6020,In_82,In_1406);
or U6021 (N_6021,In_1166,In_628);
nor U6022 (N_6022,In_1307,In_1065);
or U6023 (N_6023,In_1172,In_1648);
xor U6024 (N_6024,In_2496,In_116);
nand U6025 (N_6025,In_55,In_2345);
and U6026 (N_6026,In_1273,In_110);
nor U6027 (N_6027,In_100,In_1942);
nor U6028 (N_6028,In_332,In_1368);
and U6029 (N_6029,In_1993,In_1733);
and U6030 (N_6030,In_1662,In_1308);
nand U6031 (N_6031,In_2337,In_2484);
nor U6032 (N_6032,In_1669,In_500);
and U6033 (N_6033,In_703,In_202);
and U6034 (N_6034,In_2217,In_2139);
nor U6035 (N_6035,In_872,In_840);
or U6036 (N_6036,In_254,In_154);
and U6037 (N_6037,In_2166,In_560);
and U6038 (N_6038,In_2280,In_34);
nor U6039 (N_6039,In_143,In_578);
and U6040 (N_6040,In_575,In_565);
nor U6041 (N_6041,In_2409,In_1242);
nand U6042 (N_6042,In_1450,In_1866);
nand U6043 (N_6043,In_260,In_789);
and U6044 (N_6044,In_1575,In_1559);
and U6045 (N_6045,In_1178,In_965);
nor U6046 (N_6046,In_2379,In_1297);
nor U6047 (N_6047,In_77,In_2252);
nand U6048 (N_6048,In_1640,In_2212);
xnor U6049 (N_6049,In_2331,In_379);
nor U6050 (N_6050,In_1928,In_1293);
nor U6051 (N_6051,In_1166,In_2403);
nor U6052 (N_6052,In_1716,In_462);
or U6053 (N_6053,In_2298,In_964);
nand U6054 (N_6054,In_111,In_945);
xor U6055 (N_6055,In_1714,In_1208);
and U6056 (N_6056,In_931,In_2086);
xnor U6057 (N_6057,In_1277,In_2191);
nand U6058 (N_6058,In_1195,In_1939);
nor U6059 (N_6059,In_2173,In_734);
xor U6060 (N_6060,In_724,In_2409);
nor U6061 (N_6061,In_699,In_1426);
nand U6062 (N_6062,In_1696,In_1541);
or U6063 (N_6063,In_1626,In_917);
or U6064 (N_6064,In_1276,In_1934);
and U6065 (N_6065,In_253,In_2123);
nand U6066 (N_6066,In_1243,In_2362);
and U6067 (N_6067,In_726,In_1318);
nand U6068 (N_6068,In_992,In_2301);
xor U6069 (N_6069,In_658,In_410);
and U6070 (N_6070,In_2476,In_1864);
nand U6071 (N_6071,In_2211,In_574);
nand U6072 (N_6072,In_2336,In_2366);
or U6073 (N_6073,In_250,In_1925);
nand U6074 (N_6074,In_903,In_2121);
nand U6075 (N_6075,In_1750,In_2195);
nand U6076 (N_6076,In_1622,In_1112);
xnor U6077 (N_6077,In_543,In_1758);
or U6078 (N_6078,In_1935,In_633);
xnor U6079 (N_6079,In_857,In_1574);
nor U6080 (N_6080,In_1703,In_1433);
or U6081 (N_6081,In_54,In_1877);
xor U6082 (N_6082,In_110,In_412);
and U6083 (N_6083,In_2221,In_2309);
and U6084 (N_6084,In_121,In_362);
xor U6085 (N_6085,In_2075,In_2289);
xor U6086 (N_6086,In_1561,In_2457);
xnor U6087 (N_6087,In_1598,In_2461);
nand U6088 (N_6088,In_448,In_2357);
or U6089 (N_6089,In_462,In_1513);
xnor U6090 (N_6090,In_2310,In_1589);
or U6091 (N_6091,In_1570,In_2488);
xor U6092 (N_6092,In_2142,In_2181);
or U6093 (N_6093,In_618,In_211);
nor U6094 (N_6094,In_1958,In_2149);
nor U6095 (N_6095,In_937,In_719);
nor U6096 (N_6096,In_583,In_1637);
nor U6097 (N_6097,In_1810,In_2138);
nand U6098 (N_6098,In_977,In_1255);
and U6099 (N_6099,In_1420,In_450);
or U6100 (N_6100,In_778,In_1411);
xor U6101 (N_6101,In_1070,In_117);
or U6102 (N_6102,In_118,In_847);
nand U6103 (N_6103,In_1130,In_196);
or U6104 (N_6104,In_1818,In_1280);
or U6105 (N_6105,In_623,In_1179);
nand U6106 (N_6106,In_2072,In_2402);
nor U6107 (N_6107,In_1213,In_1171);
nand U6108 (N_6108,In_120,In_899);
nor U6109 (N_6109,In_688,In_2164);
nand U6110 (N_6110,In_1927,In_929);
and U6111 (N_6111,In_863,In_1692);
xor U6112 (N_6112,In_1450,In_2210);
or U6113 (N_6113,In_1615,In_335);
nand U6114 (N_6114,In_941,In_1776);
nand U6115 (N_6115,In_2303,In_1439);
or U6116 (N_6116,In_1752,In_2139);
and U6117 (N_6117,In_1363,In_1909);
xnor U6118 (N_6118,In_1816,In_2392);
and U6119 (N_6119,In_1553,In_800);
and U6120 (N_6120,In_2074,In_248);
or U6121 (N_6121,In_1696,In_0);
and U6122 (N_6122,In_483,In_2095);
xnor U6123 (N_6123,In_1606,In_1272);
nand U6124 (N_6124,In_2448,In_1570);
nor U6125 (N_6125,In_613,In_61);
nand U6126 (N_6126,In_1167,In_1335);
nor U6127 (N_6127,In_632,In_1101);
or U6128 (N_6128,In_982,In_890);
xnor U6129 (N_6129,In_132,In_290);
xnor U6130 (N_6130,In_849,In_888);
xor U6131 (N_6131,In_625,In_2348);
xnor U6132 (N_6132,In_201,In_1223);
nor U6133 (N_6133,In_1527,In_1548);
or U6134 (N_6134,In_1216,In_2220);
and U6135 (N_6135,In_1026,In_1453);
nor U6136 (N_6136,In_2220,In_54);
or U6137 (N_6137,In_996,In_256);
or U6138 (N_6138,In_2251,In_1806);
xnor U6139 (N_6139,In_1509,In_413);
xnor U6140 (N_6140,In_1321,In_2064);
nand U6141 (N_6141,In_24,In_853);
and U6142 (N_6142,In_161,In_1993);
and U6143 (N_6143,In_286,In_1409);
and U6144 (N_6144,In_1501,In_1327);
and U6145 (N_6145,In_866,In_1164);
and U6146 (N_6146,In_1716,In_673);
nor U6147 (N_6147,In_1152,In_2094);
and U6148 (N_6148,In_1186,In_1915);
nand U6149 (N_6149,In_542,In_2289);
nor U6150 (N_6150,In_724,In_720);
or U6151 (N_6151,In_1611,In_623);
and U6152 (N_6152,In_265,In_146);
xnor U6153 (N_6153,In_1925,In_426);
nand U6154 (N_6154,In_938,In_1069);
xor U6155 (N_6155,In_2017,In_149);
nor U6156 (N_6156,In_759,In_1995);
and U6157 (N_6157,In_1449,In_1646);
and U6158 (N_6158,In_714,In_508);
xnor U6159 (N_6159,In_2202,In_1523);
nor U6160 (N_6160,In_180,In_2377);
or U6161 (N_6161,In_88,In_1646);
or U6162 (N_6162,In_2418,In_500);
xor U6163 (N_6163,In_2255,In_2269);
and U6164 (N_6164,In_133,In_2460);
nor U6165 (N_6165,In_758,In_479);
nor U6166 (N_6166,In_2274,In_2431);
xnor U6167 (N_6167,In_1162,In_1761);
or U6168 (N_6168,In_1366,In_671);
xor U6169 (N_6169,In_1445,In_16);
nand U6170 (N_6170,In_275,In_1648);
nand U6171 (N_6171,In_522,In_2169);
nor U6172 (N_6172,In_2115,In_1563);
and U6173 (N_6173,In_844,In_2433);
nor U6174 (N_6174,In_1277,In_892);
or U6175 (N_6175,In_798,In_1810);
nor U6176 (N_6176,In_1506,In_1719);
and U6177 (N_6177,In_1935,In_1579);
and U6178 (N_6178,In_494,In_2158);
and U6179 (N_6179,In_1875,In_576);
nand U6180 (N_6180,In_2366,In_2122);
or U6181 (N_6181,In_1762,In_441);
nand U6182 (N_6182,In_2070,In_2003);
and U6183 (N_6183,In_397,In_1813);
nor U6184 (N_6184,In_731,In_1212);
xnor U6185 (N_6185,In_9,In_1724);
or U6186 (N_6186,In_2457,In_1168);
or U6187 (N_6187,In_1148,In_1092);
nor U6188 (N_6188,In_986,In_2165);
nand U6189 (N_6189,In_1770,In_672);
xor U6190 (N_6190,In_2244,In_422);
or U6191 (N_6191,In_765,In_2488);
nand U6192 (N_6192,In_1935,In_664);
nand U6193 (N_6193,In_2015,In_2281);
xnor U6194 (N_6194,In_2247,In_1547);
xnor U6195 (N_6195,In_2033,In_184);
and U6196 (N_6196,In_2090,In_1032);
and U6197 (N_6197,In_604,In_235);
xnor U6198 (N_6198,In_1179,In_30);
nor U6199 (N_6199,In_579,In_2123);
and U6200 (N_6200,In_970,In_2490);
or U6201 (N_6201,In_2093,In_1941);
nor U6202 (N_6202,In_1354,In_1076);
xnor U6203 (N_6203,In_1150,In_1369);
nand U6204 (N_6204,In_1721,In_1242);
xnor U6205 (N_6205,In_797,In_127);
and U6206 (N_6206,In_1260,In_522);
and U6207 (N_6207,In_2027,In_2479);
xor U6208 (N_6208,In_2231,In_1349);
or U6209 (N_6209,In_386,In_1166);
nand U6210 (N_6210,In_142,In_683);
nor U6211 (N_6211,In_1746,In_1431);
xnor U6212 (N_6212,In_701,In_404);
and U6213 (N_6213,In_2481,In_1302);
xnor U6214 (N_6214,In_274,In_168);
nand U6215 (N_6215,In_1003,In_1225);
nor U6216 (N_6216,In_352,In_2400);
nor U6217 (N_6217,In_773,In_50);
and U6218 (N_6218,In_644,In_1113);
or U6219 (N_6219,In_2332,In_230);
nor U6220 (N_6220,In_1485,In_2127);
and U6221 (N_6221,In_629,In_1181);
xnor U6222 (N_6222,In_34,In_997);
xnor U6223 (N_6223,In_671,In_270);
or U6224 (N_6224,In_887,In_771);
or U6225 (N_6225,In_2077,In_1705);
xnor U6226 (N_6226,In_2164,In_2025);
and U6227 (N_6227,In_928,In_213);
and U6228 (N_6228,In_354,In_1224);
or U6229 (N_6229,In_592,In_2177);
nand U6230 (N_6230,In_1267,In_1165);
or U6231 (N_6231,In_1521,In_2371);
nor U6232 (N_6232,In_1787,In_2241);
nor U6233 (N_6233,In_418,In_391);
and U6234 (N_6234,In_1597,In_1900);
nor U6235 (N_6235,In_2494,In_1169);
or U6236 (N_6236,In_350,In_1601);
nor U6237 (N_6237,In_1503,In_498);
xor U6238 (N_6238,In_1330,In_675);
and U6239 (N_6239,In_687,In_2218);
nand U6240 (N_6240,In_764,In_2040);
nor U6241 (N_6241,In_1338,In_1094);
and U6242 (N_6242,In_2225,In_2218);
nor U6243 (N_6243,In_1473,In_1283);
or U6244 (N_6244,In_1880,In_933);
nor U6245 (N_6245,In_1461,In_660);
xor U6246 (N_6246,In_1175,In_1810);
xor U6247 (N_6247,In_1468,In_767);
or U6248 (N_6248,In_66,In_230);
nor U6249 (N_6249,In_1811,In_489);
nor U6250 (N_6250,N_933,N_3991);
and U6251 (N_6251,N_5545,N_3897);
and U6252 (N_6252,N_2773,N_2604);
and U6253 (N_6253,N_4812,N_1307);
nand U6254 (N_6254,N_5372,N_4560);
nor U6255 (N_6255,N_5185,N_6209);
and U6256 (N_6256,N_4109,N_451);
and U6257 (N_6257,N_4834,N_2362);
nand U6258 (N_6258,N_2164,N_516);
nand U6259 (N_6259,N_3162,N_5730);
nand U6260 (N_6260,N_1459,N_339);
or U6261 (N_6261,N_946,N_3782);
and U6262 (N_6262,N_4829,N_1063);
nand U6263 (N_6263,N_2612,N_1917);
or U6264 (N_6264,N_4489,N_4221);
or U6265 (N_6265,N_3003,N_4943);
and U6266 (N_6266,N_6108,N_2640);
nor U6267 (N_6267,N_1205,N_160);
xnor U6268 (N_6268,N_2494,N_5209);
and U6269 (N_6269,N_6167,N_4683);
nor U6270 (N_6270,N_932,N_5184);
nand U6271 (N_6271,N_142,N_1873);
or U6272 (N_6272,N_4995,N_4103);
xnor U6273 (N_6273,N_2405,N_4973);
nor U6274 (N_6274,N_2923,N_4934);
or U6275 (N_6275,N_2349,N_3879);
and U6276 (N_6276,N_1876,N_2653);
xnor U6277 (N_6277,N_2384,N_2308);
and U6278 (N_6278,N_4291,N_4009);
xnor U6279 (N_6279,N_4397,N_3772);
or U6280 (N_6280,N_1815,N_3519);
nand U6281 (N_6281,N_4106,N_1452);
xnor U6282 (N_6282,N_1090,N_5889);
xnor U6283 (N_6283,N_1145,N_11);
xnor U6284 (N_6284,N_880,N_1223);
nor U6285 (N_6285,N_1572,N_2326);
and U6286 (N_6286,N_4940,N_5325);
or U6287 (N_6287,N_5631,N_4907);
and U6288 (N_6288,N_1260,N_5382);
or U6289 (N_6289,N_4767,N_4749);
nor U6290 (N_6290,N_4609,N_742);
and U6291 (N_6291,N_3787,N_1637);
xor U6292 (N_6292,N_1927,N_518);
nor U6293 (N_6293,N_5276,N_5333);
or U6294 (N_6294,N_154,N_3270);
xor U6295 (N_6295,N_5704,N_2068);
xnor U6296 (N_6296,N_3946,N_5739);
nor U6297 (N_6297,N_1940,N_3129);
and U6298 (N_6298,N_2208,N_107);
nand U6299 (N_6299,N_302,N_2287);
nor U6300 (N_6300,N_3076,N_1949);
and U6301 (N_6301,N_0,N_216);
nand U6302 (N_6302,N_2944,N_4753);
nand U6303 (N_6303,N_924,N_4313);
nor U6304 (N_6304,N_508,N_3307);
or U6305 (N_6305,N_1044,N_5532);
nand U6306 (N_6306,N_822,N_5943);
nand U6307 (N_6307,N_4153,N_596);
or U6308 (N_6308,N_1505,N_200);
and U6309 (N_6309,N_140,N_6082);
or U6310 (N_6310,N_4408,N_1904);
xnor U6311 (N_6311,N_1237,N_4021);
nand U6312 (N_6312,N_1833,N_6064);
xnor U6313 (N_6313,N_3631,N_1339);
nor U6314 (N_6314,N_5831,N_4805);
or U6315 (N_6315,N_4688,N_3503);
or U6316 (N_6316,N_1640,N_105);
and U6317 (N_6317,N_873,N_2516);
or U6318 (N_6318,N_5025,N_4962);
or U6319 (N_6319,N_4233,N_796);
nand U6320 (N_6320,N_1476,N_453);
and U6321 (N_6321,N_953,N_5021);
nand U6322 (N_6322,N_2151,N_994);
or U6323 (N_6323,N_2966,N_43);
or U6324 (N_6324,N_5200,N_3878);
and U6325 (N_6325,N_3396,N_356);
nand U6326 (N_6326,N_492,N_5472);
or U6327 (N_6327,N_3889,N_3013);
or U6328 (N_6328,N_5969,N_1651);
nor U6329 (N_6329,N_1694,N_1606);
xor U6330 (N_6330,N_736,N_992);
or U6331 (N_6331,N_2450,N_4020);
or U6332 (N_6332,N_5544,N_3380);
nor U6333 (N_6333,N_5534,N_2753);
or U6334 (N_6334,N_4682,N_5525);
nor U6335 (N_6335,N_6141,N_6109);
xnor U6336 (N_6336,N_4541,N_4900);
xnor U6337 (N_6337,N_4949,N_1207);
nand U6338 (N_6338,N_2144,N_252);
nor U6339 (N_6339,N_3045,N_5024);
and U6340 (N_6340,N_2254,N_1338);
xnor U6341 (N_6341,N_5441,N_2314);
or U6342 (N_6342,N_3639,N_909);
xor U6343 (N_6343,N_3952,N_6044);
xor U6344 (N_6344,N_4612,N_3979);
and U6345 (N_6345,N_4809,N_5772);
nor U6346 (N_6346,N_340,N_3750);
and U6347 (N_6347,N_4290,N_2150);
and U6348 (N_6348,N_983,N_5416);
or U6349 (N_6349,N_1231,N_2203);
or U6350 (N_6350,N_4051,N_1422);
xor U6351 (N_6351,N_1152,N_1678);
nor U6352 (N_6352,N_4214,N_5787);
and U6353 (N_6353,N_1209,N_979);
xor U6354 (N_6354,N_1866,N_4244);
xnor U6355 (N_6355,N_5082,N_2005);
or U6356 (N_6356,N_1586,N_5947);
nor U6357 (N_6357,N_361,N_2272);
nor U6358 (N_6358,N_127,N_4019);
xor U6359 (N_6359,N_3723,N_772);
nand U6360 (N_6360,N_4968,N_2479);
nor U6361 (N_6361,N_2976,N_632);
xor U6362 (N_6362,N_5454,N_4909);
or U6363 (N_6363,N_807,N_5320);
xor U6364 (N_6364,N_5049,N_929);
and U6365 (N_6365,N_2820,N_3858);
or U6366 (N_6366,N_5809,N_2665);
nand U6367 (N_6367,N_4737,N_4704);
xnor U6368 (N_6368,N_3106,N_259);
nor U6369 (N_6369,N_834,N_3704);
nor U6370 (N_6370,N_5361,N_2410);
and U6371 (N_6371,N_5196,N_4887);
nand U6372 (N_6372,N_6084,N_5229);
nor U6373 (N_6373,N_5150,N_2477);
or U6374 (N_6374,N_3993,N_1334);
or U6375 (N_6375,N_902,N_1082);
and U6376 (N_6376,N_2674,N_1031);
and U6377 (N_6377,N_5503,N_2236);
or U6378 (N_6378,N_2731,N_1448);
xnor U6379 (N_6379,N_5285,N_4288);
xor U6380 (N_6380,N_3887,N_5955);
and U6381 (N_6381,N_4360,N_3105);
xor U6382 (N_6382,N_5788,N_5425);
xor U6383 (N_6383,N_1493,N_5379);
nor U6384 (N_6384,N_1652,N_4450);
nor U6385 (N_6385,N_4657,N_3851);
nor U6386 (N_6386,N_5204,N_3699);
xor U6387 (N_6387,N_5565,N_4321);
and U6388 (N_6388,N_3786,N_3619);
or U6389 (N_6389,N_4403,N_274);
nor U6390 (N_6390,N_6124,N_2412);
nor U6391 (N_6391,N_2109,N_2040);
or U6392 (N_6392,N_3612,N_237);
xnor U6393 (N_6393,N_6101,N_2488);
xnor U6394 (N_6394,N_1976,N_5006);
xor U6395 (N_6395,N_3660,N_5849);
xnor U6396 (N_6396,N_912,N_4026);
nor U6397 (N_6397,N_229,N_1633);
or U6398 (N_6398,N_3967,N_2163);
nor U6399 (N_6399,N_2324,N_6138);
nor U6400 (N_6400,N_6061,N_2469);
xor U6401 (N_6401,N_757,N_592);
and U6402 (N_6402,N_1988,N_1955);
nor U6403 (N_6403,N_5804,N_2235);
xor U6404 (N_6404,N_4857,N_2948);
and U6405 (N_6405,N_2610,N_2845);
nand U6406 (N_6406,N_472,N_3199);
and U6407 (N_6407,N_3232,N_3022);
xor U6408 (N_6408,N_5368,N_2293);
xor U6409 (N_6409,N_1696,N_3789);
nand U6410 (N_6410,N_5376,N_1043);
or U6411 (N_6411,N_218,N_3100);
nand U6412 (N_6412,N_2379,N_5658);
or U6413 (N_6413,N_1605,N_3385);
nand U6414 (N_6414,N_4952,N_735);
nand U6415 (N_6415,N_2505,N_2213);
nor U6416 (N_6416,N_3138,N_3605);
or U6417 (N_6417,N_6234,N_4782);
nor U6418 (N_6418,N_2438,N_609);
or U6419 (N_6419,N_1925,N_2698);
nand U6420 (N_6420,N_1120,N_5836);
xor U6421 (N_6421,N_3883,N_1329);
xnor U6422 (N_6422,N_6146,N_4309);
nand U6423 (N_6423,N_4084,N_5973);
nand U6424 (N_6424,N_1982,N_145);
xor U6425 (N_6425,N_3743,N_5106);
and U6426 (N_6426,N_1822,N_5666);
and U6427 (N_6427,N_3513,N_4517);
or U6428 (N_6428,N_3689,N_5300);
nand U6429 (N_6429,N_2912,N_4792);
nor U6430 (N_6430,N_1810,N_2840);
or U6431 (N_6431,N_5263,N_5046);
and U6432 (N_6432,N_5426,N_146);
xor U6433 (N_6433,N_1749,N_5984);
nand U6434 (N_6434,N_3779,N_5612);
xnor U6435 (N_6435,N_1746,N_2296);
or U6436 (N_6436,N_3661,N_1932);
or U6437 (N_6437,N_6112,N_6071);
nor U6438 (N_6438,N_5220,N_3831);
and U6439 (N_6439,N_2004,N_3222);
and U6440 (N_6440,N_1861,N_4908);
and U6441 (N_6441,N_1534,N_852);
and U6442 (N_6442,N_1497,N_5863);
nor U6443 (N_6443,N_3215,N_2320);
nor U6444 (N_6444,N_799,N_1164);
nor U6445 (N_6445,N_2327,N_840);
xor U6446 (N_6446,N_6107,N_5340);
or U6447 (N_6447,N_4384,N_3367);
and U6448 (N_6448,N_4929,N_493);
nand U6449 (N_6449,N_1217,N_185);
or U6450 (N_6450,N_3680,N_5564);
or U6451 (N_6451,N_2549,N_3525);
or U6452 (N_6452,N_5607,N_3566);
or U6453 (N_6453,N_4405,N_2202);
xnor U6454 (N_6454,N_6191,N_2560);
xor U6455 (N_6455,N_4735,N_3522);
or U6456 (N_6456,N_4811,N_5594);
and U6457 (N_6457,N_4056,N_1563);
nor U6458 (N_6458,N_2078,N_5750);
and U6459 (N_6459,N_5711,N_5897);
or U6460 (N_6460,N_484,N_608);
nand U6461 (N_6461,N_2413,N_5855);
xor U6462 (N_6462,N_5164,N_2493);
nor U6463 (N_6463,N_925,N_877);
or U6464 (N_6464,N_2016,N_3854);
or U6465 (N_6465,N_2717,N_1972);
and U6466 (N_6466,N_6157,N_897);
nand U6467 (N_6467,N_684,N_4236);
nand U6468 (N_6468,N_5362,N_3590);
nand U6469 (N_6469,N_2597,N_6090);
and U6470 (N_6470,N_5946,N_5131);
nand U6471 (N_6471,N_4827,N_3486);
and U6472 (N_6472,N_4326,N_2533);
and U6473 (N_6473,N_2222,N_4184);
xnor U6474 (N_6474,N_3456,N_4761);
xor U6475 (N_6475,N_3824,N_3810);
and U6476 (N_6476,N_588,N_1681);
or U6477 (N_6477,N_1764,N_4891);
nand U6478 (N_6478,N_1475,N_4849);
and U6479 (N_6479,N_2969,N_3527);
and U6480 (N_6480,N_1403,N_4577);
xor U6481 (N_6481,N_995,N_827);
or U6482 (N_6482,N_5094,N_5850);
and U6483 (N_6483,N_404,N_4462);
or U6484 (N_6484,N_293,N_2748);
xor U6485 (N_6485,N_253,N_2161);
nor U6486 (N_6486,N_6104,N_67);
nand U6487 (N_6487,N_5347,N_3769);
and U6488 (N_6488,N_2357,N_2981);
xnor U6489 (N_6489,N_2908,N_4672);
or U6490 (N_6490,N_4766,N_2531);
or U6491 (N_6491,N_2485,N_1585);
nand U6492 (N_6492,N_1745,N_3707);
and U6493 (N_6493,N_3646,N_3412);
or U6494 (N_6494,N_1113,N_5640);
and U6495 (N_6495,N_1457,N_247);
and U6496 (N_6496,N_558,N_6135);
nand U6497 (N_6497,N_6202,N_2134);
xor U6498 (N_6498,N_4378,N_3264);
and U6499 (N_6499,N_5352,N_4629);
and U6500 (N_6500,N_4882,N_1786);
and U6501 (N_6501,N_872,N_878);
nand U6502 (N_6502,N_5488,N_4063);
nor U6503 (N_6503,N_5490,N_5538);
and U6504 (N_6504,N_4961,N_4198);
nor U6505 (N_6505,N_2782,N_582);
nand U6506 (N_6506,N_5696,N_2375);
and U6507 (N_6507,N_5090,N_3033);
xor U6508 (N_6508,N_956,N_3895);
nor U6509 (N_6509,N_4215,N_1716);
and U6510 (N_6510,N_1358,N_4796);
nand U6511 (N_6511,N_3599,N_307);
nand U6512 (N_6512,N_5899,N_5625);
xor U6513 (N_6513,N_4711,N_5098);
nor U6514 (N_6514,N_4387,N_2309);
nor U6515 (N_6515,N_2921,N_3450);
xnor U6516 (N_6516,N_2386,N_5950);
xor U6517 (N_6517,N_6119,N_2081);
nor U6518 (N_6518,N_4391,N_1996);
nor U6519 (N_6519,N_2775,N_1446);
nand U6520 (N_6520,N_480,N_5664);
nor U6521 (N_6521,N_1395,N_1084);
and U6522 (N_6522,N_3829,N_3682);
nor U6523 (N_6523,N_5790,N_3475);
or U6524 (N_6524,N_2749,N_1426);
nor U6525 (N_6525,N_4700,N_2591);
or U6526 (N_6526,N_4052,N_3694);
and U6527 (N_6527,N_1985,N_5732);
or U6528 (N_6528,N_347,N_4365);
nor U6529 (N_6529,N_4947,N_5695);
nand U6530 (N_6530,N_387,N_1445);
and U6531 (N_6531,N_5143,N_3179);
nand U6532 (N_6532,N_5092,N_4859);
and U6533 (N_6533,N_6125,N_3103);
nor U6534 (N_6534,N_6024,N_208);
and U6535 (N_6535,N_4126,N_4837);
and U6536 (N_6536,N_261,N_5309);
nor U6537 (N_6537,N_3902,N_4108);
and U6538 (N_6538,N_1235,N_667);
nor U6539 (N_6539,N_2300,N_2816);
or U6540 (N_6540,N_3067,N_2274);
nand U6541 (N_6541,N_1901,N_2524);
xnor U6542 (N_6542,N_4987,N_3280);
nor U6543 (N_6543,N_4062,N_2183);
nand U6544 (N_6544,N_5477,N_618);
xnor U6545 (N_6545,N_3257,N_2044);
xor U6546 (N_6546,N_1142,N_5223);
nor U6547 (N_6547,N_5822,N_1523);
and U6548 (N_6548,N_1492,N_943);
or U6549 (N_6549,N_6099,N_4427);
and U6550 (N_6550,N_4006,N_6201);
xor U6551 (N_6551,N_1343,N_3039);
and U6552 (N_6552,N_2012,N_3400);
nor U6553 (N_6553,N_5518,N_560);
nand U6554 (N_6554,N_600,N_3524);
nor U6555 (N_6555,N_5939,N_3693);
nor U6556 (N_6556,N_1874,N_2434);
or U6557 (N_6557,N_1021,N_189);
nor U6558 (N_6558,N_1653,N_867);
nand U6559 (N_6559,N_5255,N_3742);
xnor U6560 (N_6560,N_2294,N_2862);
nand U6561 (N_6561,N_2866,N_1539);
or U6562 (N_6562,N_4698,N_3186);
or U6563 (N_6563,N_2529,N_3271);
nor U6564 (N_6564,N_3384,N_2657);
xor U6565 (N_6565,N_616,N_2446);
and U6566 (N_6566,N_370,N_539);
nor U6567 (N_6567,N_821,N_1923);
or U6568 (N_6568,N_407,N_2846);
nand U6569 (N_6569,N_4640,N_732);
and U6570 (N_6570,N_963,N_198);
or U6571 (N_6571,N_441,N_1624);
and U6572 (N_6572,N_5685,N_694);
nand U6573 (N_6573,N_298,N_405);
nand U6574 (N_6574,N_4188,N_5608);
or U6575 (N_6575,N_5630,N_1070);
and U6576 (N_6576,N_5166,N_3021);
or U6577 (N_6577,N_1373,N_5869);
nand U6578 (N_6578,N_5222,N_512);
or U6579 (N_6579,N_5174,N_1228);
xor U6580 (N_6580,N_433,N_5231);
or U6581 (N_6581,N_5641,N_883);
xor U6582 (N_6582,N_2869,N_1051);
xnor U6583 (N_6583,N_2280,N_4129);
or U6584 (N_6584,N_3868,N_4658);
or U6585 (N_6585,N_1608,N_915);
xnor U6586 (N_6586,N_4912,N_6227);
or U6587 (N_6587,N_4027,N_2718);
and U6588 (N_6588,N_393,N_6106);
nor U6589 (N_6589,N_5590,N_2942);
or U6590 (N_6590,N_4663,N_2933);
nand U6591 (N_6591,N_678,N_3618);
or U6592 (N_6592,N_106,N_4162);
nor U6593 (N_6593,N_2204,N_5703);
xnor U6594 (N_6594,N_683,N_1361);
and U6595 (N_6595,N_5448,N_2961);
and U6596 (N_6596,N_5643,N_4773);
or U6597 (N_6597,N_213,N_3261);
and U6598 (N_6598,N_5107,N_1580);
or U6599 (N_6599,N_1530,N_5815);
nor U6600 (N_6600,N_4446,N_431);
nor U6601 (N_6601,N_335,N_529);
nor U6602 (N_6602,N_171,N_5951);
nand U6603 (N_6603,N_301,N_227);
nand U6604 (N_6604,N_1919,N_969);
or U6605 (N_6605,N_2681,N_3212);
and U6606 (N_6606,N_5919,N_5306);
nor U6607 (N_6607,N_4016,N_5183);
nand U6608 (N_6608,N_4581,N_1524);
nor U6609 (N_6609,N_2655,N_4477);
or U6610 (N_6610,N_6,N_6034);
and U6611 (N_6611,N_4150,N_2009);
and U6612 (N_6612,N_841,N_2960);
xor U6613 (N_6613,N_156,N_3720);
xnor U6614 (N_6614,N_5879,N_5660);
xnor U6615 (N_6615,N_2979,N_4259);
nand U6616 (N_6616,N_1480,N_2700);
xnor U6617 (N_6617,N_6028,N_6088);
nor U6618 (N_6618,N_6115,N_1303);
xor U6619 (N_6619,N_1515,N_3511);
or U6620 (N_6620,N_3908,N_3019);
xor U6621 (N_6621,N_1751,N_1087);
nor U6622 (N_6622,N_2066,N_1258);
nand U6623 (N_6623,N_4240,N_465);
xor U6624 (N_6624,N_6154,N_428);
and U6625 (N_6625,N_5635,N_3101);
xnor U6626 (N_6626,N_4183,N_3551);
nor U6627 (N_6627,N_3855,N_4636);
xor U6628 (N_6628,N_3393,N_1748);
nand U6629 (N_6629,N_4161,N_5410);
and U6630 (N_6630,N_4239,N_4127);
and U6631 (N_6631,N_4249,N_2790);
nor U6632 (N_6632,N_2715,N_3095);
and U6633 (N_6633,N_1269,N_2685);
nor U6634 (N_6634,N_2833,N_763);
and U6635 (N_6635,N_3500,N_222);
nand U6636 (N_6636,N_3625,N_4421);
nor U6637 (N_6637,N_2891,N_6226);
xor U6638 (N_6638,N_3184,N_4538);
or U6639 (N_6639,N_1545,N_5875);
and U6640 (N_6640,N_4706,N_5508);
or U6641 (N_6641,N_766,N_4209);
and U6642 (N_6642,N_1892,N_4713);
nand U6643 (N_6643,N_3477,N_1865);
or U6644 (N_6644,N_1970,N_3240);
xor U6645 (N_6645,N_3172,N_1879);
xnor U6646 (N_6646,N_1344,N_1083);
xnor U6647 (N_6647,N_3165,N_5818);
xor U6648 (N_6648,N_95,N_1841);
nor U6649 (N_6649,N_4960,N_3637);
or U6650 (N_6650,N_4025,N_5672);
and U6651 (N_6651,N_217,N_6233);
or U6652 (N_6652,N_4145,N_5353);
or U6653 (N_6653,N_916,N_3131);
xnor U6654 (N_6654,N_5398,N_993);
xnor U6655 (N_6655,N_2950,N_934);
or U6656 (N_6656,N_4347,N_6188);
xnor U6657 (N_6657,N_5535,N_2954);
nand U6658 (N_6658,N_5171,N_906);
or U6659 (N_6659,N_1806,N_291);
or U6660 (N_6660,N_3490,N_4433);
and U6661 (N_6661,N_3430,N_2802);
nand U6662 (N_6662,N_378,N_3096);
nor U6663 (N_6663,N_1360,N_1491);
or U6664 (N_6664,N_5527,N_4953);
and U6665 (N_6665,N_2171,N_5032);
xnor U6666 (N_6666,N_3239,N_186);
nor U6667 (N_6667,N_2528,N_3840);
or U6668 (N_6668,N_6019,N_1671);
and U6669 (N_6669,N_3933,N_5087);
nor U6670 (N_6670,N_334,N_5820);
nand U6671 (N_6671,N_2955,N_1770);
and U6672 (N_6672,N_3320,N_5470);
and U6673 (N_6673,N_6147,N_811);
xor U6674 (N_6674,N_3959,N_455);
xnor U6675 (N_6675,N_1897,N_5045);
and U6676 (N_6676,N_2087,N_874);
or U6677 (N_6677,N_4603,N_3091);
nor U6678 (N_6678,N_4457,N_295);
or U6679 (N_6679,N_3536,N_1193);
and U6680 (N_6680,N_52,N_1049);
nor U6681 (N_6681,N_411,N_4554);
nor U6682 (N_6682,N_2812,N_6070);
xnor U6683 (N_6683,N_2116,N_2936);
and U6684 (N_6684,N_1001,N_1836);
xor U6685 (N_6685,N_2145,N_4583);
or U6686 (N_6686,N_3960,N_3417);
xor U6687 (N_6687,N_5668,N_1827);
or U6688 (N_6688,N_3009,N_1868);
nor U6689 (N_6689,N_3964,N_2750);
or U6690 (N_6690,N_4734,N_2378);
xnor U6691 (N_6691,N_1712,N_865);
nand U6692 (N_6692,N_3148,N_3717);
xor U6693 (N_6693,N_5186,N_4675);
or U6694 (N_6694,N_3808,N_5001);
nand U6695 (N_6695,N_2433,N_5233);
xor U6696 (N_6696,N_3079,N_6100);
or U6697 (N_6697,N_4567,N_4911);
nor U6698 (N_6698,N_5253,N_2777);
nor U6699 (N_6699,N_6048,N_2152);
nand U6700 (N_6700,N_3837,N_94);
and U6701 (N_6701,N_4558,N_5011);
nand U6702 (N_6702,N_964,N_5840);
nor U6703 (N_6703,N_1462,N_2886);
or U6704 (N_6704,N_3956,N_5782);
xor U6705 (N_6705,N_2607,N_5550);
xor U6706 (N_6706,N_6152,N_886);
xor U6707 (N_6707,N_2588,N_6161);
or U6708 (N_6708,N_5471,N_1644);
nand U6709 (N_6709,N_4097,N_2818);
nand U6710 (N_6710,N_354,N_4177);
and U6711 (N_6711,N_1076,N_5676);
nor U6712 (N_6712,N_2805,N_634);
xnor U6713 (N_6713,N_6089,N_172);
nor U6714 (N_6714,N_5418,N_4059);
nand U6715 (N_6715,N_3201,N_5278);
and U6716 (N_6716,N_1799,N_2423);
or U6717 (N_6717,N_3112,N_2959);
nand U6718 (N_6718,N_3474,N_1754);
or U6719 (N_6719,N_3405,N_5059);
nor U6720 (N_6720,N_1857,N_1625);
xnor U6721 (N_6721,N_1790,N_3501);
xor U6722 (N_6722,N_5043,N_5913);
xnor U6723 (N_6723,N_6130,N_2963);
and U6724 (N_6724,N_1573,N_507);
nand U6725 (N_6725,N_5719,N_5111);
nor U6726 (N_6726,N_464,N_743);
nand U6727 (N_6727,N_5742,N_1397);
or U6728 (N_6728,N_4057,N_2015);
or U6729 (N_6729,N_2053,N_124);
nand U6730 (N_6730,N_3623,N_6229);
xnor U6731 (N_6731,N_2489,N_4394);
xnor U6732 (N_6732,N_4996,N_1283);
xor U6733 (N_6733,N_4200,N_2964);
or U6734 (N_6734,N_648,N_2683);
nor U6735 (N_6735,N_1595,N_479);
and U6736 (N_6736,N_5243,N_3411);
xor U6737 (N_6737,N_2023,N_2870);
or U6738 (N_6738,N_1276,N_5316);
xor U6739 (N_6739,N_4740,N_6219);
nor U6740 (N_6740,N_2579,N_5561);
nand U6741 (N_6741,N_39,N_2508);
nor U6742 (N_6742,N_3074,N_5293);
nor U6743 (N_6743,N_4265,N_3927);
xnor U6744 (N_6744,N_402,N_2216);
and U6745 (N_6745,N_1944,N_1202);
or U6746 (N_6746,N_4725,N_5069);
xor U6747 (N_6747,N_5462,N_3903);
nor U6748 (N_6748,N_344,N_4122);
nor U6749 (N_6749,N_483,N_4283);
and U6750 (N_6750,N_1842,N_3616);
xnor U6751 (N_6751,N_2074,N_3622);
or U6752 (N_6752,N_1778,N_1248);
and U6753 (N_6753,N_3802,N_372);
nor U6754 (N_6754,N_1060,N_3912);
xnor U6755 (N_6755,N_3277,N_1359);
nand U6756 (N_6756,N_1460,N_242);
and U6757 (N_6757,N_2894,N_1085);
xor U6758 (N_6758,N_5778,N_5883);
xor U6759 (N_6759,N_6001,N_5030);
and U6760 (N_6760,N_2571,N_1992);
nor U6761 (N_6761,N_2435,N_5530);
xnor U6762 (N_6762,N_5281,N_5560);
and U6763 (N_6763,N_3735,N_2352);
nor U6764 (N_6764,N_5400,N_3173);
nor U6765 (N_6765,N_1025,N_2514);
and U6766 (N_6766,N_5351,N_4373);
or U6767 (N_6767,N_3738,N_2615);
and U6768 (N_6768,N_4219,N_1702);
nand U6769 (N_6769,N_670,N_2828);
xor U6770 (N_6770,N_314,N_3109);
nand U6771 (N_6771,N_4595,N_3149);
and U6772 (N_6772,N_2772,N_4223);
and U6773 (N_6773,N_3005,N_1823);
xor U6774 (N_6774,N_4342,N_4945);
xor U6775 (N_6775,N_571,N_3630);
nor U6776 (N_6776,N_4647,N_996);
nor U6777 (N_6777,N_2257,N_5851);
nor U6778 (N_6778,N_1381,N_3754);
nand U6779 (N_6779,N_1969,N_1829);
nor U6780 (N_6780,N_4398,N_790);
nand U6781 (N_6781,N_4825,N_4042);
nor U6782 (N_6782,N_2882,N_603);
nand U6783 (N_6783,N_1700,N_6006);
nand U6784 (N_6784,N_1869,N_36);
xnor U6785 (N_6785,N_4176,N_3957);
and U6786 (N_6786,N_6065,N_526);
or U6787 (N_6787,N_5121,N_764);
xor U6788 (N_6788,N_1870,N_5865);
xnor U6789 (N_6789,N_273,N_21);
or U6790 (N_6790,N_5414,N_3128);
nand U6791 (N_6791,N_2737,N_1533);
or U6792 (N_6792,N_3992,N_2819);
xnor U6793 (N_6793,N_1386,N_1902);
and U6794 (N_6794,N_3805,N_5232);
and U6795 (N_6795,N_2224,N_1814);
nand U6796 (N_6796,N_5866,N_550);
and U6797 (N_6797,N_2086,N_5598);
or U6798 (N_6798,N_2629,N_803);
or U6799 (N_6799,N_2659,N_1638);
nand U6800 (N_6800,N_4546,N_3285);
and U6801 (N_6801,N_3675,N_158);
nor U6802 (N_6802,N_4328,N_6214);
xor U6803 (N_6803,N_1721,N_674);
and U6804 (N_6804,N_817,N_692);
nand U6805 (N_6805,N_5413,N_720);
nor U6806 (N_6806,N_1377,N_1909);
or U6807 (N_6807,N_3935,N_6046);
nand U6808 (N_6808,N_3546,N_926);
xnor U6809 (N_6809,N_209,N_4959);
or U6810 (N_6810,N_2481,N_1635);
or U6811 (N_6811,N_1320,N_3666);
or U6812 (N_6812,N_1185,N_624);
nor U6813 (N_6813,N_860,N_4550);
and U6814 (N_6814,N_5235,N_5674);
nor U6815 (N_6815,N_5614,N_3235);
xor U6816 (N_6816,N_1527,N_4717);
or U6817 (N_6817,N_3247,N_5095);
nand U6818 (N_6818,N_4821,N_4090);
nand U6819 (N_6819,N_1903,N_6045);
nor U6820 (N_6820,N_1672,N_1456);
nand U6821 (N_6821,N_1163,N_1830);
and U6822 (N_6822,N_896,N_5596);
and U6823 (N_6823,N_446,N_4190);
xor U6824 (N_6824,N_4083,N_3617);
and U6825 (N_6825,N_5944,N_5816);
and U6826 (N_6826,N_1081,N_966);
nor U6827 (N_6827,N_5738,N_96);
and U6828 (N_6828,N_5086,N_4765);
nand U6829 (N_6829,N_2745,N_535);
xnor U6830 (N_6830,N_704,N_5593);
nand U6831 (N_6831,N_2578,N_3340);
nor U6832 (N_6832,N_323,N_3026);
nand U6833 (N_6833,N_1102,N_2428);
xnor U6834 (N_6834,N_2317,N_3073);
and U6835 (N_6835,N_5331,N_305);
nand U6836 (N_6836,N_776,N_2095);
nand U6837 (N_6837,N_4637,N_3634);
or U6838 (N_6838,N_2470,N_4362);
and U6839 (N_6839,N_330,N_4716);
nand U6840 (N_6840,N_1689,N_6230);
xor U6841 (N_6841,N_3465,N_4061);
or U6842 (N_6842,N_3489,N_1654);
xor U6843 (N_6843,N_972,N_1659);
or U6844 (N_6844,N_4802,N_4482);
nor U6845 (N_6845,N_269,N_3414);
nor U6846 (N_6846,N_1126,N_1285);
or U6847 (N_6847,N_3462,N_325);
nor U6848 (N_6848,N_2266,N_656);
nor U6849 (N_6849,N_4091,N_28);
nand U6850 (N_6850,N_3234,N_1756);
or U6851 (N_6851,N_6132,N_4493);
nor U6852 (N_6852,N_3081,N_1943);
nor U6853 (N_6853,N_133,N_2118);
or U6854 (N_6854,N_4522,N_4422);
nand U6855 (N_6855,N_5582,N_5305);
and U6856 (N_6856,N_4588,N_57);
or U6857 (N_6857,N_3934,N_1738);
or U6858 (N_6858,N_5050,N_3667);
xor U6859 (N_6859,N_6078,N_2584);
nand U6860 (N_6860,N_4054,N_4497);
nor U6861 (N_6861,N_4179,N_3379);
and U6862 (N_6862,N_2207,N_833);
nor U6863 (N_6863,N_4768,N_6123);
nor U6864 (N_6864,N_3007,N_1680);
nand U6865 (N_6865,N_5431,N_3410);
nand U6866 (N_6866,N_3950,N_1407);
and U6867 (N_6867,N_3092,N_3585);
nand U6868 (N_6868,N_1559,N_4628);
nor U6869 (N_6869,N_3523,N_3495);
nor U6870 (N_6870,N_5245,N_3867);
nor U6871 (N_6871,N_5862,N_3594);
nor U6872 (N_6872,N_4844,N_5385);
nand U6873 (N_6873,N_2030,N_4838);
or U6874 (N_6874,N_1350,N_3482);
xnor U6875 (N_6875,N_4831,N_4438);
or U6876 (N_6876,N_745,N_42);
and U6877 (N_6877,N_4339,N_3632);
and U6878 (N_6878,N_4424,N_5447);
nand U6879 (N_6879,N_1785,N_5803);
and U6880 (N_6880,N_3722,N_3183);
or U6881 (N_6881,N_1157,N_2611);
nor U6882 (N_6882,N_6043,N_6022);
nand U6883 (N_6883,N_3168,N_780);
or U6884 (N_6884,N_5290,N_6190);
nand U6885 (N_6885,N_3161,N_2227);
nand U6886 (N_6886,N_6185,N_5452);
nor U6887 (N_6887,N_3088,N_6240);
xnor U6888 (N_6888,N_5683,N_3804);
and U6889 (N_6889,N_1747,N_1349);
and U6890 (N_6890,N_3355,N_1977);
nor U6891 (N_6891,N_738,N_4490);
nand U6892 (N_6892,N_197,N_4687);
nor U6893 (N_6893,N_238,N_2103);
and U6894 (N_6894,N_3378,N_4324);
nand U6895 (N_6895,N_6239,N_2376);
nor U6896 (N_6896,N_271,N_2896);
nand U6897 (N_6897,N_102,N_4079);
nand U6898 (N_6898,N_1424,N_5084);
xnor U6899 (N_6899,N_2543,N_4876);
xnor U6900 (N_6900,N_2632,N_5230);
xor U6901 (N_6901,N_6086,N_3304);
and U6902 (N_6902,N_1341,N_1845);
nor U6903 (N_6903,N_3955,N_727);
or U6904 (N_6904,N_1722,N_1012);
and U6905 (N_6905,N_5602,N_5387);
nand U6906 (N_6906,N_1108,N_2860);
nor U6907 (N_6907,N_2407,N_2922);
nand U6908 (N_6908,N_5236,N_3494);
and U6909 (N_6909,N_2836,N_2644);
or U6910 (N_6910,N_3374,N_1317);
or U6911 (N_6911,N_1301,N_5964);
xor U6912 (N_6912,N_4860,N_3930);
nand U6913 (N_6913,N_4207,N_3873);
nand U6914 (N_6914,N_5187,N_279);
or U6915 (N_6915,N_2011,N_4262);
nand U6916 (N_6916,N_2603,N_6140);
or U6917 (N_6917,N_4074,N_3588);
and U6918 (N_6918,N_6150,N_617);
or U6919 (N_6919,N_1675,N_4923);
and U6920 (N_6920,N_496,N_6018);
or U6921 (N_6921,N_1136,N_3251);
nor U6922 (N_6922,N_4044,N_3770);
or U6923 (N_6923,N_3901,N_3206);
or U6924 (N_6924,N_3517,N_5348);
nand U6925 (N_6925,N_4224,N_581);
nor U6926 (N_6926,N_1905,N_108);
nand U6927 (N_6927,N_1732,N_2186);
or U6928 (N_6928,N_4480,N_1332);
nor U6929 (N_6929,N_5918,N_1168);
nand U6930 (N_6930,N_3455,N_205);
and U6931 (N_6931,N_3958,N_3446);
and U6932 (N_6932,N_957,N_2598);
and U6933 (N_6933,N_4479,N_2451);
and U6934 (N_6934,N_2071,N_5128);
nand U6935 (N_6935,N_1111,N_2523);
nand U6936 (N_6936,N_664,N_406);
nand U6937 (N_6937,N_3066,N_5694);
or U6938 (N_6938,N_686,N_3461);
and U6939 (N_6939,N_3552,N_3300);
and U6940 (N_6940,N_3228,N_3645);
xnor U6941 (N_6941,N_1280,N_3702);
xor U6942 (N_6942,N_338,N_3187);
xnor U6943 (N_6943,N_5770,N_5456);
nand U6944 (N_6944,N_519,N_2721);
nand U6945 (N_6945,N_2953,N_3424);
or U6946 (N_6946,N_5224,N_3975);
and U6947 (N_6947,N_3048,N_1396);
and U6948 (N_6948,N_1392,N_6095);
xor U6949 (N_6949,N_1498,N_5479);
xor U6950 (N_6950,N_310,N_3783);
nand U6951 (N_6951,N_2429,N_33);
nor U6952 (N_6952,N_644,N_4516);
or U6953 (N_6953,N_1391,N_2929);
and U6954 (N_6954,N_5386,N_1007);
or U6955 (N_6955,N_3940,N_3180);
nand U6956 (N_6956,N_2594,N_5894);
xnor U6957 (N_6957,N_3124,N_5146);
xnor U6958 (N_6958,N_2388,N_3529);
nor U6959 (N_6959,N_1400,N_5838);
and U6960 (N_6960,N_3850,N_4251);
xnor U6961 (N_6961,N_2399,N_2425);
and U6962 (N_6962,N_2858,N_3740);
nor U6963 (N_6963,N_3954,N_4757);
and U6964 (N_6964,N_1047,N_4864);
xor U6965 (N_6965,N_4915,N_895);
and U6966 (N_6966,N_4978,N_3174);
nand U6967 (N_6967,N_3929,N_215);
xor U6968 (N_6968,N_698,N_3828);
and U6969 (N_6969,N_1667,N_437);
nor U6970 (N_6970,N_2783,N_4899);
xor U6971 (N_6971,N_2347,N_3611);
and U6972 (N_6972,N_2643,N_2853);
or U6973 (N_6973,N_4335,N_540);
and U6974 (N_6974,N_882,N_777);
xnor U6975 (N_6975,N_6091,N_2634);
xor U6976 (N_6976,N_53,N_2967);
or U6977 (N_6977,N_5466,N_1528);
and U6978 (N_6978,N_4664,N_5284);
or U6979 (N_6979,N_2082,N_4211);
and U6980 (N_6980,N_3163,N_4715);
nand U6981 (N_6981,N_4846,N_2689);
xor U6982 (N_6982,N_4692,N_1466);
nand U6983 (N_6983,N_977,N_5036);
nor U6984 (N_6984,N_2895,N_5731);
and U6985 (N_6985,N_5942,N_1881);
nand U6986 (N_6986,N_5832,N_2199);
nor U6987 (N_6987,N_2465,N_6092);
or U6988 (N_6988,N_1146,N_4893);
nor U6989 (N_6989,N_1851,N_5007);
xor U6990 (N_6990,N_3139,N_4178);
xnor U6991 (N_6991,N_4801,N_4948);
and U6992 (N_6992,N_2427,N_3914);
or U6993 (N_6993,N_921,N_4295);
nand U6994 (N_6994,N_2613,N_3063);
or U6995 (N_6995,N_5190,N_1619);
xnor U6996 (N_6996,N_4002,N_1251);
or U6997 (N_6997,N_2888,N_5747);
nor U6998 (N_6998,N_4730,N_506);
or U6999 (N_6999,N_2218,N_5632);
and U7000 (N_7000,N_181,N_5321);
xnor U7001 (N_7001,N_5211,N_3592);
nor U7002 (N_7002,N_5902,N_6128);
and U7003 (N_7003,N_5307,N_5475);
nor U7004 (N_7004,N_4884,N_5626);
xnor U7005 (N_7005,N_1180,N_3922);
xor U7006 (N_7006,N_575,N_767);
xor U7007 (N_7007,N_1556,N_4505);
nor U7008 (N_7008,N_4304,N_2080);
xnor U7009 (N_7009,N_2740,N_3428);
xor U7010 (N_7010,N_5012,N_2455);
or U7011 (N_7011,N_202,N_1924);
and U7012 (N_7012,N_3980,N_3921);
nor U7013 (N_7013,N_2400,N_1346);
and U7014 (N_7014,N_4048,N_5142);
nor U7015 (N_7015,N_3575,N_4333);
nand U7016 (N_7016,N_2621,N_169);
nand U7017 (N_7017,N_2867,N_4856);
xor U7018 (N_7018,N_1929,N_1907);
or U7019 (N_7019,N_5935,N_1225);
xor U7020 (N_7020,N_315,N_1128);
xor U7021 (N_7021,N_832,N_3947);
and U7022 (N_7022,N_542,N_1692);
xnor U7023 (N_7023,N_153,N_1981);
nand U7024 (N_7024,N_4684,N_1388);
nor U7025 (N_7025,N_3532,N_1368);
nor U7026 (N_7026,N_5713,N_4545);
xor U7027 (N_7027,N_4447,N_5239);
xnor U7028 (N_7028,N_1316,N_6002);
nand U7029 (N_7029,N_3464,N_5286);
nor U7030 (N_7030,N_3539,N_3449);
or U7031 (N_7031,N_2055,N_4889);
nand U7032 (N_7032,N_1479,N_4524);
nor U7033 (N_7033,N_4358,N_6156);
or U7034 (N_7034,N_4419,N_2297);
or U7035 (N_7035,N_2492,N_6011);
xor U7036 (N_7036,N_5769,N_2211);
nand U7037 (N_7037,N_2911,N_5078);
and U7038 (N_7038,N_5210,N_5161);
nor U7039 (N_7039,N_4954,N_196);
or U7040 (N_7040,N_1171,N_2822);
nand U7041 (N_7041,N_5112,N_1995);
nand U7042 (N_7042,N_2447,N_3057);
and U7043 (N_7043,N_3994,N_5274);
and U7044 (N_7044,N_791,N_1568);
nand U7045 (N_7045,N_5776,N_1883);
nor U7046 (N_7046,N_2977,N_3028);
and U7047 (N_7047,N_2147,N_751);
xnor U7048 (N_7048,N_1987,N_1310);
and U7049 (N_7049,N_5374,N_4785);
or U7050 (N_7050,N_2075,N_5749);
nor U7051 (N_7051,N_1971,N_1313);
xnor U7052 (N_7052,N_5657,N_2471);
nor U7053 (N_7053,N_3973,N_5445);
nand U7054 (N_7054,N_2160,N_3020);
or U7055 (N_7055,N_1399,N_2335);
or U7056 (N_7056,N_5578,N_311);
nor U7057 (N_7057,N_4372,N_4096);
xnor U7058 (N_7058,N_1779,N_2099);
xnor U7059 (N_7059,N_3181,N_4067);
xnor U7060 (N_7060,N_4736,N_4494);
nand U7061 (N_7061,N_6080,N_3422);
xor U7062 (N_7062,N_2061,N_1352);
xnor U7063 (N_7063,N_4351,N_1551);
nor U7064 (N_7064,N_798,N_2337);
nand U7065 (N_7065,N_3190,N_4064);
xor U7066 (N_7066,N_5597,N_2623);
and U7067 (N_7067,N_5117,N_1464);
and U7068 (N_7068,N_3319,N_5123);
xor U7069 (N_7069,N_5960,N_3915);
nor U7070 (N_7070,N_5589,N_3778);
and U7071 (N_7071,N_5442,N_1305);
nand U7072 (N_7072,N_318,N_653);
and U7073 (N_7073,N_1941,N_5624);
nand U7074 (N_7074,N_3357,N_2017);
nor U7075 (N_7075,N_3999,N_231);
nor U7076 (N_7076,N_3170,N_2766);
and U7077 (N_7077,N_2270,N_392);
and U7078 (N_7078,N_7,N_4518);
or U7079 (N_7079,N_1507,N_3712);
xor U7080 (N_7080,N_5698,N_4449);
and U7081 (N_7081,N_3093,N_1335);
xor U7082 (N_7082,N_3258,N_2008);
and U7083 (N_7083,N_337,N_594);
nor U7084 (N_7084,N_5267,N_1284);
or U7085 (N_7085,N_3542,N_3528);
and U7086 (N_7086,N_2664,N_5020);
nand U7087 (N_7087,N_2628,N_2641);
or U7088 (N_7088,N_1516,N_4793);
nand U7089 (N_7089,N_2617,N_4902);
nor U7090 (N_7090,N_3535,N_1817);
nor U7091 (N_7091,N_3753,N_111);
and U7092 (N_7092,N_848,N_520);
xor U7093 (N_7093,N_3880,N_2563);
xor U7094 (N_7094,N_1394,N_2687);
or U7095 (N_7095,N_2032,N_666);
or U7096 (N_7096,N_5439,N_221);
xor U7097 (N_7097,N_4140,N_4294);
or U7098 (N_7098,N_5812,N_3147);
nand U7099 (N_7099,N_4468,N_2305);
nand U7100 (N_7100,N_5162,N_5740);
nor U7101 (N_7101,N_3077,N_374);
and U7102 (N_7102,N_3273,N_4344);
and U7103 (N_7103,N_1300,N_697);
or U7104 (N_7104,N_6212,N_3852);
nor U7105 (N_7105,N_5487,N_4514);
or U7106 (N_7106,N_4620,N_117);
and U7107 (N_7107,N_2581,N_6160);
nand U7108 (N_7108,N_1591,N_5420);
and U7109 (N_7109,N_4944,N_4147);
and U7110 (N_7110,N_4903,N_869);
and U7111 (N_7111,N_5659,N_403);
nand U7112 (N_7112,N_4511,N_4038);
or U7113 (N_7113,N_4937,N_3118);
and U7114 (N_7114,N_3122,N_3766);
or U7115 (N_7115,N_627,N_5334);
nor U7116 (N_7116,N_2024,N_2467);
nor U7117 (N_7117,N_6241,N_2339);
nor U7118 (N_7118,N_4787,N_1383);
or U7119 (N_7119,N_5254,N_3196);
nand U7120 (N_7120,N_889,N_6208);
xnor U7121 (N_7121,N_5982,N_32);
and U7122 (N_7122,N_1765,N_2177);
nor U7123 (N_7123,N_3084,N_1803);
and U7124 (N_7124,N_3870,N_3031);
xor U7125 (N_7125,N_6013,N_2088);
or U7126 (N_7126,N_2938,N_5921);
nand U7127 (N_7127,N_5934,N_482);
nand U7128 (N_7128,N_2408,N_5514);
xor U7129 (N_7129,N_2825,N_5541);
nand U7130 (N_7130,N_1115,N_225);
or U7131 (N_7131,N_5781,N_4374);
nor U7132 (N_7132,N_4616,N_2031);
or U7133 (N_7133,N_1072,N_4203);
nor U7134 (N_7134,N_6008,N_3387);
and U7135 (N_7135,N_6204,N_1192);
xnor U7136 (N_7136,N_2215,N_3705);
or U7137 (N_7137,N_5102,N_839);
and U7138 (N_7138,N_5500,N_4041);
and U7139 (N_7139,N_155,N_3158);
nor U7140 (N_7140,N_368,N_23);
or U7141 (N_7141,N_1942,N_4602);
or U7142 (N_7142,N_4544,N_249);
nor U7143 (N_7143,N_1615,N_2230);
and U7144 (N_7144,N_3860,N_4369);
or U7145 (N_7145,N_2616,N_5081);
nor U7146 (N_7146,N_4395,N_4182);
nand U7147 (N_7147,N_8,N_650);
or U7148 (N_7148,N_6038,N_6131);
xor U7149 (N_7149,N_1038,N_1106);
and U7150 (N_7150,N_5355,N_4642);
or U7151 (N_7151,N_4705,N_2139);
nor U7152 (N_7152,N_5129,N_4037);
nor U7153 (N_7153,N_2431,N_5194);
nand U7154 (N_7154,N_5868,N_6096);
or U7155 (N_7155,N_1206,N_3688);
and U7156 (N_7156,N_2101,N_4904);
nand U7157 (N_7157,N_3364,N_3359);
or U7158 (N_7158,N_5465,N_4828);
or U7159 (N_7159,N_2680,N_3288);
nand U7160 (N_7160,N_4573,N_5342);
xor U7161 (N_7161,N_3569,N_6228);
or U7162 (N_7162,N_5890,N_3407);
xnor U7163 (N_7163,N_6235,N_6232);
nand U7164 (N_7164,N_705,N_2338);
nor U7165 (N_7165,N_187,N_2196);
and U7166 (N_7166,N_2136,N_5800);
or U7167 (N_7167,N_5570,N_1893);
nor U7168 (N_7168,N_1447,N_4361);
or U7169 (N_7169,N_4824,N_938);
nor U7170 (N_7170,N_4301,N_5330);
nand U7171 (N_7171,N_173,N_724);
xor U7172 (N_7172,N_1241,N_4587);
nand U7173 (N_7173,N_1630,N_1097);
or U7174 (N_7174,N_2444,N_4241);
nor U7175 (N_7175,N_5707,N_3035);
and U7176 (N_7176,N_5228,N_3709);
xor U7177 (N_7177,N_4777,N_4731);
and U7178 (N_7178,N_4257,N_1831);
and U7179 (N_7179,N_5743,N_5833);
or U7180 (N_7180,N_2541,N_468);
and U7181 (N_7181,N_1835,N_2618);
nand U7182 (N_7182,N_557,N_219);
and U7183 (N_7183,N_2776,N_6073);
and U7184 (N_7184,N_1268,N_3182);
nand U7185 (N_7185,N_2110,N_1244);
and U7186 (N_7186,N_3869,N_3938);
nand U7187 (N_7187,N_5345,N_2752);
xor U7188 (N_7188,N_2809,N_2374);
or U7189 (N_7189,N_800,N_1724);
nand U7190 (N_7190,N_5088,N_3730);
nand U7191 (N_7191,N_1061,N_5018);
or U7192 (N_7192,N_962,N_348);
xnor U7193 (N_7193,N_2569,N_207);
or U7194 (N_7194,N_191,N_4414);
xnor U7195 (N_7195,N_1046,N_4383);
and U7196 (N_7196,N_3441,N_4112);
nor U7197 (N_7197,N_3208,N_2231);
and U7198 (N_7198,N_2878,N_645);
and U7199 (N_7199,N_1939,N_3784);
and U7200 (N_7200,N_3269,N_5691);
nor U7201 (N_7201,N_4467,N_2237);
xor U7202 (N_7202,N_4268,N_22);
or U7203 (N_7203,N_6111,N_1683);
nand U7204 (N_7204,N_1900,N_5559);
and U7205 (N_7205,N_4121,N_3607);
or U7206 (N_7206,N_528,N_2544);
xor U7207 (N_7207,N_4982,N_3972);
nand U7208 (N_7208,N_3540,N_3537);
and U7209 (N_7209,N_5134,N_974);
or U7210 (N_7210,N_4445,N_3445);
nand U7211 (N_7211,N_4537,N_1431);
nor U7212 (N_7212,N_1908,N_2759);
and U7213 (N_7213,N_5678,N_3715);
nand U7214 (N_7214,N_5110,N_2518);
nand U7215 (N_7215,N_3732,N_3610);
nor U7216 (N_7216,N_2767,N_3691);
or U7217 (N_7217,N_5613,N_2299);
or U7218 (N_7218,N_4630,N_1933);
or U7219 (N_7219,N_1846,N_1401);
or U7220 (N_7220,N_1643,N_1503);
nand U7221 (N_7221,N_2058,N_355);
or U7222 (N_7222,N_5268,N_2456);
xor U7223 (N_7223,N_3315,N_4928);
or U7224 (N_7224,N_4810,N_5605);
and U7225 (N_7225,N_3328,N_637);
nand U7226 (N_7226,N_2262,N_611);
xor U7227 (N_7227,N_5144,N_5389);
nor U7228 (N_7228,N_24,N_1353);
xor U7229 (N_7229,N_5983,N_4312);
xor U7230 (N_7230,N_2496,N_511);
nand U7231 (N_7231,N_3308,N_809);
and U7232 (N_7232,N_2038,N_927);
nand U7233 (N_7233,N_5715,N_3254);
or U7234 (N_7234,N_3739,N_5537);
and U7235 (N_7235,N_3818,N_2645);
and U7236 (N_7236,N_2688,N_4515);
xnor U7237 (N_7237,N_1661,N_4453);
nor U7238 (N_7238,N_4417,N_2561);
and U7239 (N_7239,N_4769,N_1840);
and U7240 (N_7240,N_1686,N_88);
and U7241 (N_7241,N_4501,N_4858);
xor U7242 (N_7242,N_1254,N_3443);
nand U7243 (N_7243,N_4869,N_746);
nor U7244 (N_7244,N_1159,N_1960);
or U7245 (N_7245,N_631,N_1682);
or U7246 (N_7246,N_3626,N_2385);
and U7247 (N_7247,N_5356,N_1123);
nor U7248 (N_7248,N_1252,N_761);
and U7249 (N_7249,N_2049,N_5299);
xnor U7250 (N_7250,N_1194,N_2857);
and U7251 (N_7251,N_265,N_5350);
or U7252 (N_7252,N_4938,N_1796);
nand U7253 (N_7253,N_3352,N_2247);
xor U7254 (N_7254,N_903,N_5057);
or U7255 (N_7255,N_5887,N_2794);
nor U7256 (N_7256,N_818,N_4714);
or U7257 (N_7257,N_1406,N_2567);
and U7258 (N_7258,N_4932,N_4941);
xnor U7259 (N_7259,N_3674,N_3323);
and U7260 (N_7260,N_1918,N_4406);
nor U7261 (N_7261,N_4280,N_1805);
or U7262 (N_7262,N_395,N_4985);
xor U7263 (N_7263,N_4316,N_4261);
nand U7264 (N_7264,N_2527,N_5315);
nand U7265 (N_7265,N_949,N_435);
xor U7266 (N_7266,N_500,N_1141);
xor U7267 (N_7267,N_6184,N_4691);
and U7268 (N_7268,N_6210,N_652);
and U7269 (N_7269,N_4033,N_3483);
or U7270 (N_7270,N_3219,N_2690);
nor U7271 (N_7271,N_1578,N_3591);
nor U7272 (N_7272,N_1213,N_1058);
xnor U7273 (N_7273,N_1191,N_195);
xor U7274 (N_7274,N_2808,N_1139);
or U7275 (N_7275,N_5941,N_3899);
nand U7276 (N_7276,N_5138,N_965);
xnor U7277 (N_7277,N_2486,N_1628);
or U7278 (N_7278,N_4906,N_5981);
xor U7279 (N_7279,N_4286,N_2525);
and U7280 (N_7280,N_5422,N_1467);
or U7281 (N_7281,N_3925,N_2734);
or U7282 (N_7282,N_4113,N_3052);
and U7283 (N_7283,N_1419,N_2515);
xnor U7284 (N_7284,N_139,N_1066);
xnor U7285 (N_7285,N_5746,N_3953);
or U7286 (N_7286,N_5019,N_1609);
nor U7287 (N_7287,N_3849,N_4300);
nand U7288 (N_7288,N_2736,N_4080);
xnor U7289 (N_7289,N_959,N_1239);
or U7290 (N_7290,N_3797,N_255);
xnor U7291 (N_7291,N_3885,N_6074);
or U7292 (N_7292,N_4788,N_2072);
xor U7293 (N_7293,N_4055,N_3476);
or U7294 (N_7294,N_711,N_5893);
nand U7295 (N_7295,N_4878,N_786);
xor U7296 (N_7296,N_5002,N_3227);
or U7297 (N_7297,N_2319,N_352);
and U7298 (N_7298,N_3481,N_4274);
nor U7299 (N_7299,N_513,N_4341);
xnor U7300 (N_7300,N_3864,N_4470);
or U7301 (N_7301,N_861,N_3046);
nor U7302 (N_7302,N_3800,N_5835);
xor U7303 (N_7303,N_4246,N_1211);
nor U7304 (N_7304,N_2383,N_2306);
xor U7305 (N_7305,N_2506,N_3538);
nand U7306 (N_7306,N_264,N_5845);
xor U7307 (N_7307,N_4014,N_4918);
xor U7308 (N_7308,N_5575,N_744);
nor U7309 (N_7309,N_3238,N_2475);
nor U7310 (N_7310,N_2201,N_6197);
nor U7311 (N_7311,N_254,N_263);
nor U7312 (N_7312,N_4348,N_6016);
nor U7313 (N_7313,N_3884,N_6085);
and U7314 (N_7314,N_3724,N_3893);
and U7315 (N_7315,N_2754,N_4786);
xor U7316 (N_7316,N_6127,N_2510);
nor U7317 (N_7317,N_4591,N_3339);
nor U7318 (N_7318,N_5040,N_855);
nor U7319 (N_7319,N_3658,N_3041);
nand U7320 (N_7320,N_3404,N_1333);
nor U7321 (N_7321,N_4282,N_1602);
nand U7322 (N_7322,N_5072,N_1375);
nand U7323 (N_7323,N_695,N_1374);
nor U7324 (N_7324,N_2003,N_1465);
and U7325 (N_7325,N_819,N_5606);
nand U7326 (N_7326,N_4029,N_4181);
xor U7327 (N_7327,N_2130,N_2725);
nor U7328 (N_7328,N_1797,N_5473);
xor U7329 (N_7329,N_2893,N_1882);
xor U7330 (N_7330,N_1483,N_6189);
or U7331 (N_7331,N_4694,N_2059);
xor U7332 (N_7332,N_3189,N_4499);
nand U7333 (N_7333,N_388,N_1916);
or U7334 (N_7334,N_748,N_3518);
or U7335 (N_7335,N_1687,N_5667);
xor U7336 (N_7336,N_3656,N_911);
nand U7337 (N_7337,N_3541,N_1576);
nor U7338 (N_7338,N_4139,N_2351);
or U7339 (N_7339,N_3613,N_4305);
or U7340 (N_7340,N_2279,N_2554);
xor U7341 (N_7341,N_2387,N_2189);
xor U7342 (N_7342,N_2415,N_3296);
xor U7343 (N_7343,N_5858,N_4738);
or U7344 (N_7344,N_5857,N_2182);
nor U7345 (N_7345,N_163,N_4371);
nand U7346 (N_7346,N_5055,N_4865);
nor U7347 (N_7347,N_3792,N_2179);
nor U7348 (N_7348,N_1297,N_4748);
nor U7349 (N_7349,N_1034,N_5975);
nor U7350 (N_7350,N_409,N_17);
xor U7351 (N_7351,N_1143,N_4458);
or U7352 (N_7352,N_3002,N_1246);
nand U7353 (N_7353,N_4702,N_3624);
and U7354 (N_7354,N_2115,N_5126);
nor U7355 (N_7355,N_6081,N_2587);
xor U7356 (N_7356,N_5617,N_1623);
and U7357 (N_7357,N_241,N_975);
and U7358 (N_7358,N_6010,N_2934);
nor U7359 (N_7359,N_3497,N_3961);
and U7360 (N_7360,N_2988,N_2153);
nand U7361 (N_7361,N_5047,N_4874);
or U7362 (N_7362,N_5328,N_703);
or U7363 (N_7363,N_3628,N_3621);
xnor U7364 (N_7364,N_1453,N_1860);
nor U7365 (N_7365,N_3847,N_2865);
and U7366 (N_7366,N_2791,N_5073);
nor U7367 (N_7367,N_2765,N_2990);
or U7368 (N_7368,N_843,N_427);
or U7369 (N_7369,N_5974,N_3358);
nand U7370 (N_7370,N_5048,N_4195);
or U7371 (N_7371,N_6143,N_1760);
nor U7372 (N_7372,N_4942,N_2803);
nor U7373 (N_7373,N_1795,N_1330);
nor U7374 (N_7374,N_2982,N_3399);
nor U7375 (N_7375,N_1472,N_5871);
and U7376 (N_7376,N_3655,N_3719);
or U7377 (N_7377,N_3875,N_3721);
xor U7378 (N_7378,N_3906,N_5175);
nand U7379 (N_7379,N_5203,N_4659);
nand U7380 (N_7380,N_1685,N_2991);
xor U7381 (N_7381,N_2225,N_6216);
xor U7382 (N_7382,N_920,N_2651);
and U7383 (N_7383,N_1039,N_2155);
xnor U7384 (N_7384,N_831,N_5924);
xnor U7385 (N_7385,N_4771,N_5637);
nor U7386 (N_7386,N_1272,N_4732);
and U7387 (N_7387,N_3836,N_716);
or U7388 (N_7388,N_3447,N_2996);
or U7389 (N_7389,N_5880,N_1203);
nor U7390 (N_7390,N_5940,N_5114);
nor U7391 (N_7391,N_1501,N_2849);
xor U7392 (N_7392,N_2166,N_3633);
and U7393 (N_7393,N_914,N_870);
or U7394 (N_7394,N_753,N_5587);
or U7395 (N_7395,N_1729,N_2480);
xor U7396 (N_7396,N_3563,N_4431);
and U7397 (N_7397,N_5972,N_5802);
nand U7398 (N_7398,N_5074,N_1558);
xor U7399 (N_7399,N_3326,N_2756);
nand U7400 (N_7400,N_3318,N_1165);
or U7401 (N_7401,N_1372,N_2329);
xnor U7402 (N_7402,N_3872,N_1014);
nor U7403 (N_7403,N_3652,N_3650);
nor U7404 (N_7404,N_5977,N_4440);
nand U7405 (N_7405,N_1617,N_5282);
xnor U7406 (N_7406,N_1502,N_5931);
nor U7407 (N_7407,N_4622,N_3882);
xnor U7408 (N_7408,N_3911,N_4709);
xnor U7409 (N_7409,N_1286,N_2473);
or U7410 (N_7410,N_366,N_3086);
nor U7411 (N_7411,N_3214,N_5795);
nor U7412 (N_7412,N_1037,N_4352);
nor U7413 (N_7413,N_6062,N_5936);
and U7414 (N_7414,N_5319,N_3886);
or U7415 (N_7415,N_1234,N_3791);
nor U7416 (N_7416,N_5105,N_3714);
nand U7417 (N_7417,N_51,N_3926);
and U7418 (N_7418,N_3102,N_5681);
and U7419 (N_7419,N_2125,N_3132);
nor U7420 (N_7420,N_662,N_3821);
nand U7421 (N_7421,N_6168,N_1632);
and U7422 (N_7422,N_4726,N_5434);
xor U7423 (N_7423,N_4755,N_5828);
xor U7424 (N_7424,N_4644,N_551);
nor U7425 (N_7425,N_210,N_2797);
nor U7426 (N_7426,N_5958,N_147);
or U7427 (N_7427,N_3602,N_2345);
and U7428 (N_7428,N_3796,N_4165);
or U7429 (N_7429,N_5633,N_5008);
xor U7430 (N_7430,N_6164,N_2361);
or U7431 (N_7431,N_5044,N_2986);
nand U7432 (N_7432,N_72,N_1022);
or U7433 (N_7433,N_5039,N_3001);
nor U7434 (N_7434,N_2596,N_3143);
nand U7435 (N_7435,N_910,N_4266);
and U7436 (N_7436,N_4886,N_4879);
nor U7437 (N_7437,N_2484,N_2804);
and U7438 (N_7438,N_68,N_2916);
and U7439 (N_7439,N_408,N_3309);
nor U7440 (N_7440,N_568,N_4046);
nor U7441 (N_7441,N_1348,N_4235);
nand U7442 (N_7442,N_4230,N_922);
nand U7443 (N_7443,N_4024,N_3008);
xor U7444 (N_7444,N_5159,N_5751);
xor U7445 (N_7445,N_1574,N_4665);
xnor U7446 (N_7446,N_991,N_3265);
nand U7447 (N_7447,N_3,N_415);
nor U7448 (N_7448,N_1253,N_723);
nand U7449 (N_7449,N_5783,N_6151);
nand U7450 (N_7450,N_2835,N_4509);
or U7451 (N_7451,N_3983,N_5509);
or U7452 (N_7452,N_802,N_2924);
xnor U7453 (N_7453,N_4432,N_4132);
xnor U7454 (N_7454,N_2132,N_2951);
nor U7455 (N_7455,N_2260,N_4349);
nand U7456 (N_7456,N_6114,N_5557);
nor U7457 (N_7457,N_1931,N_1440);
nor U7458 (N_7458,N_2897,N_4851);
or U7459 (N_7459,N_421,N_1816);
xor U7460 (N_7460,N_591,N_1910);
nand U7461 (N_7461,N_3762,N_1198);
and U7462 (N_7462,N_5415,N_6247);
and U7463 (N_7463,N_4739,N_2646);
or U7464 (N_7464,N_2122,N_103);
and U7465 (N_7465,N_369,N_1218);
or U7466 (N_7466,N_19,N_4654);
xnor U7467 (N_7467,N_585,N_167);
nor U7468 (N_7468,N_986,N_5392);
xnor U7469 (N_7469,N_3635,N_1557);
nor U7470 (N_7470,N_5085,N_4625);
and U7471 (N_7471,N_534,N_121);
or U7472 (N_7472,N_3493,N_351);
and U7473 (N_7473,N_722,N_2649);
and U7474 (N_7474,N_3337,N_1922);
xnor U7475 (N_7475,N_3609,N_2000);
and U7476 (N_7476,N_1912,N_2318);
nand U7477 (N_7477,N_300,N_5834);
or U7478 (N_7478,N_707,N_2601);
and U7479 (N_7479,N_2089,N_2768);
xor U7480 (N_7480,N_6198,N_34);
and U7481 (N_7481,N_466,N_4100);
and U7482 (N_7482,N_6116,N_5218);
nand U7483 (N_7483,N_6103,N_5004);
xnor U7484 (N_7484,N_3436,N_5761);
or U7485 (N_7485,N_4334,N_5177);
xnor U7486 (N_7486,N_3888,N_935);
xor U7487 (N_7487,N_691,N_3344);
and U7488 (N_7488,N_5189,N_3568);
and U7489 (N_7489,N_2441,N_3543);
nand U7490 (N_7490,N_178,N_4407);
and U7491 (N_7491,N_4293,N_2255);
xnor U7492 (N_7492,N_289,N_143);
and U7493 (N_7493,N_3900,N_5895);
and U7494 (N_7494,N_980,N_6003);
and U7495 (N_7495,N_2709,N_1915);
xnor U7496 (N_7496,N_3917,N_5796);
nand U7497 (N_7497,N_4319,N_4222);
nand U7498 (N_7498,N_1616,N_5735);
nor U7499 (N_7499,N_5584,N_6098);
nor U7500 (N_7500,N_6137,N_1802);
and U7501 (N_7501,N_1130,N_5406);
xnor U7502 (N_7502,N_1232,N_1701);
nor U7503 (N_7503,N_5149,N_3460);
nand U7504 (N_7504,N_1104,N_1676);
or U7505 (N_7505,N_5642,N_5373);
xor U7506 (N_7506,N_3050,N_3734);
nand U7507 (N_7507,N_3844,N_2704);
nand U7508 (N_7508,N_4970,N_1322);
and U7509 (N_7509,N_2392,N_6047);
and U7510 (N_7510,N_981,N_5764);
nand U7511 (N_7511,N_1532,N_3297);
and U7512 (N_7512,N_6030,N_1148);
xor U7513 (N_7513,N_1362,N_3562);
or U7514 (N_7514,N_2807,N_5497);
or U7515 (N_7515,N_5327,N_5480);
nor U7516 (N_7516,N_5493,N_1782);
xor U7517 (N_7517,N_5517,N_1825);
xnor U7518 (N_7518,N_2701,N_1318);
nor U7519 (N_7519,N_3094,N_1994);
and U7520 (N_7520,N_1065,N_2786);
and U7521 (N_7521,N_5157,N_2310);
xnor U7522 (N_7522,N_4572,N_235);
and U7523 (N_7523,N_4066,N_4604);
and U7524 (N_7524,N_623,N_4728);
nor U7525 (N_7525,N_1511,N_654);
and U7526 (N_7526,N_5793,N_5992);
xnor U7527 (N_7527,N_5013,N_3759);
nor U7528 (N_7528,N_1596,N_5917);
nand U7529 (N_7529,N_2770,N_5369);
nor U7530 (N_7530,N_1314,N_2285);
nand U7531 (N_7531,N_4491,N_236);
nand U7532 (N_7532,N_3386,N_4094);
or U7533 (N_7533,N_1030,N_434);
xor U7534 (N_7534,N_1668,N_2298);
or U7535 (N_7535,N_700,N_2682);
and U7536 (N_7536,N_2522,N_4689);
nand U7537 (N_7537,N_567,N_2393);
xor U7538 (N_7538,N_3224,N_3974);
and U7539 (N_7539,N_5450,N_1116);
or U7540 (N_7540,N_1024,N_577);
nand U7541 (N_7541,N_5338,N_308);
nor U7542 (N_7542,N_5063,N_4166);
xnor U7543 (N_7543,N_5219,N_982);
or U7544 (N_7544,N_2624,N_3905);
or U7545 (N_7545,N_2273,N_5847);
xnor U7546 (N_7546,N_5912,N_5152);
and U7547 (N_7547,N_5484,N_3423);
nand U7548 (N_7548,N_5725,N_3371);
nand U7549 (N_7549,N_2968,N_3069);
or U7550 (N_7550,N_1016,N_1517);
nor U7551 (N_7551,N_774,N_3098);
xnor U7552 (N_7552,N_714,N_1020);
nor U7553 (N_7553,N_680,N_5677);
xnor U7554 (N_7554,N_2271,N_4790);
nor U7555 (N_7555,N_2238,N_256);
or U7556 (N_7556,N_6170,N_967);
nor U7557 (N_7557,N_4783,N_4813);
and U7558 (N_7558,N_2158,N_1017);
or U7559 (N_7559,N_1581,N_4443);
xor U7560 (N_7560,N_5404,N_3761);
nand U7561 (N_7561,N_1514,N_4815);
nor U7562 (N_7562,N_1062,N_2033);
and U7563 (N_7563,N_3089,N_1250);
xnor U7564 (N_7564,N_5600,N_416);
or U7565 (N_7565,N_240,N_2021);
nand U7566 (N_7566,N_4245,N_3571);
and U7567 (N_7567,N_3703,N_2970);
nand U7568 (N_7568,N_625,N_4561);
or U7569 (N_7569,N_5323,N_2478);
nand U7570 (N_7570,N_923,N_3341);
or U7571 (N_7571,N_1990,N_2937);
or U7572 (N_7572,N_5501,N_968);
nor U7573 (N_7573,N_1366,N_2432);
or U7574 (N_7574,N_5581,N_4566);
and U7575 (N_7575,N_3383,N_287);
or U7576 (N_7576,N_4191,N_4131);
or U7577 (N_7577,N_3256,N_2291);
and U7578 (N_7578,N_6223,N_134);
xor U7579 (N_7579,N_3194,N_3644);
xor U7580 (N_7580,N_3560,N_988);
xnor U7581 (N_7581,N_2173,N_1914);
nor U7582 (N_7582,N_2864,N_2143);
xnor U7583 (N_7583,N_2422,N_3727);
or U7584 (N_7584,N_3241,N_4719);
nand U7585 (N_7585,N_1811,N_4680);
nor U7586 (N_7586,N_4742,N_5915);
and U7587 (N_7587,N_5486,N_3555);
nand U7588 (N_7588,N_635,N_1854);
nor U7589 (N_7589,N_2394,N_816);
or U7590 (N_7590,N_4791,N_2788);
and U7591 (N_7591,N_4306,N_1801);
nor U7592 (N_7592,N_812,N_1565);
nor U7593 (N_7593,N_5033,N_6049);
xor U7594 (N_7594,N_6040,N_4120);
and U7595 (N_7595,N_3225,N_1147);
xor U7596 (N_7596,N_4969,N_1880);
xnor U7597 (N_7597,N_5837,N_866);
xor U7598 (N_7598,N_1812,N_485);
and U7599 (N_7599,N_3231,N_3894);
or U7600 (N_7600,N_5799,N_1490);
nand U7601 (N_7601,N_3576,N_1621);
or U7602 (N_7602,N_4510,N_6148);
nand U7603 (N_7603,N_2779,N_3207);
xnor U7604 (N_7604,N_4086,N_2250);
nor U7605 (N_7605,N_3113,N_5773);
xnor U7606 (N_7606,N_3395,N_1720);
xnor U7607 (N_7607,N_4413,N_1266);
nand U7608 (N_7608,N_2699,N_476);
or U7609 (N_7609,N_5539,N_1962);
xor U7610 (N_7610,N_3205,N_503);
and U7611 (N_7611,N_5930,N_1056);
nor U7612 (N_7612,N_4641,N_2693);
nand U7613 (N_7613,N_2253,N_2219);
or U7614 (N_7614,N_423,N_1278);
or U7615 (N_7615,N_4476,N_5080);
nor U7616 (N_7616,N_2176,N_10);
nand U7617 (N_7617,N_5549,N_984);
and U7618 (N_7618,N_5402,N_3037);
xor U7619 (N_7619,N_829,N_3292);
xnor U7620 (N_7620,N_2212,N_595);
and U7621 (N_7621,N_3303,N_2630);
or U7622 (N_7622,N_5669,N_4368);
or U7623 (N_7623,N_2875,N_3369);
or U7624 (N_7624,N_4703,N_3790);
xnor U7625 (N_7625,N_2558,N_607);
nand U7626 (N_7626,N_2915,N_3653);
nor U7627 (N_7627,N_1839,N_4451);
and U7628 (N_7628,N_157,N_2763);
nor U7629 (N_7629,N_1363,N_2719);
nor U7630 (N_7630,N_5714,N_3279);
and U7631 (N_7631,N_4474,N_258);
and U7632 (N_7632,N_3141,N_2856);
nand U7633 (N_7633,N_5118,N_4154);
nand U7634 (N_7634,N_1040,N_3565);
nand U7635 (N_7635,N_379,N_5882);
or U7636 (N_7636,N_5824,N_1947);
nand U7637 (N_7637,N_5929,N_3487);
xor U7638 (N_7638,N_3289,N_3556);
nor U7639 (N_7639,N_2036,N_2842);
xnor U7640 (N_7640,N_5444,N_1529);
nor U7641 (N_7641,N_3171,N_1601);
nor U7642 (N_7642,N_1098,N_4610);
and U7643 (N_7643,N_367,N_3090);
nand U7644 (N_7644,N_725,N_1184);
xnor U7645 (N_7645,N_4946,N_1264);
nand U7646 (N_7646,N_1665,N_2168);
and U7647 (N_7647,N_808,N_3659);
xnor U7648 (N_7648,N_952,N_2495);
xor U7649 (N_7649,N_3636,N_4818);
nand U7650 (N_7650,N_665,N_1646);
and U7651 (N_7651,N_3806,N_92);
xor U7652 (N_7652,N_4930,N_4194);
nor U7653 (N_7653,N_4201,N_6200);
xor U7654 (N_7654,N_6207,N_2787);
nor U7655 (N_7655,N_2054,N_1315);
nor U7656 (N_7656,N_5364,N_2542);
and U7657 (N_7657,N_3731,N_3117);
nand U7658 (N_7658,N_212,N_5234);
and U7659 (N_7659,N_3321,N_4584);
xor U7660 (N_7660,N_2589,N_5566);
and U7661 (N_7661,N_5645,N_6113);
or U7662 (N_7662,N_5060,N_5458);
or U7663 (N_7663,N_4576,N_5756);
or U7664 (N_7664,N_5303,N_306);
and U7665 (N_7665,N_2686,N_5188);
or U7666 (N_7666,N_2877,N_1135);
nor U7667 (N_7667,N_5226,N_4830);
and U7668 (N_7668,N_2281,N_363);
xor U7669 (N_7669,N_5363,N_190);
or U7670 (N_7670,N_1292,N_5628);
and U7671 (N_7671,N_2198,N_1834);
nand U7672 (N_7672,N_2952,N_5344);
nand U7673 (N_7673,N_1398,N_5846);
nand U7674 (N_7674,N_5215,N_45);
and U7675 (N_7675,N_2974,N_5221);
and U7676 (N_7676,N_5572,N_5979);
and U7677 (N_7677,N_4107,N_2192);
xor U7678 (N_7678,N_2365,N_4173);
and U7679 (N_7679,N_2321,N_4314);
xnor U7680 (N_7680,N_2824,N_5670);
and U7681 (N_7681,N_1849,N_844);
or U7682 (N_7682,N_2830,N_1221);
nor U7683 (N_7683,N_1186,N_5180);
or U7684 (N_7684,N_2586,N_3586);
and U7685 (N_7685,N_2743,N_730);
xor U7686 (N_7686,N_4998,N_5817);
or U7687 (N_7687,N_1520,N_1734);
or U7688 (N_7688,N_1858,N_4243);
nand U7689 (N_7689,N_2184,N_1666);
or U7690 (N_7690,N_3177,N_1004);
nor U7691 (N_7691,N_3942,N_1064);
nand U7692 (N_7692,N_6177,N_223);
and U7693 (N_7693,N_789,N_5213);
nand U7694 (N_7694,N_184,N_412);
nand U7695 (N_7695,N_2670,N_3040);
xnor U7696 (N_7696,N_1864,N_239);
and U7697 (N_7697,N_729,N_1800);
nand U7698 (N_7698,N_4163,N_2993);
or U7699 (N_7699,N_4034,N_4285);
and U7700 (N_7700,N_4017,N_2056);
xnor U7701 (N_7701,N_4187,N_2667);
and U7702 (N_7702,N_1593,N_3425);
or U7703 (N_7703,N_3943,N_5101);
xnor U7704 (N_7704,N_3298,N_1259);
nand U7705 (N_7705,N_3266,N_100);
and U7706 (N_7706,N_2156,N_2512);
nor U7707 (N_7707,N_2232,N_48);
nor U7708 (N_7708,N_4039,N_5901);
xor U7709 (N_7709,N_2574,N_6035);
nor U7710 (N_7710,N_5591,N_1478);
xnor U7711 (N_7711,N_4327,N_1416);
nand U7712 (N_7712,N_1414,N_2368);
and U7713 (N_7713,N_3043,N_971);
xnor U7714 (N_7714,N_3603,N_2943);
xnor U7715 (N_7715,N_4833,N_4852);
xor U7716 (N_7716,N_6169,N_2223);
or U7717 (N_7717,N_1302,N_159);
nand U7718 (N_7718,N_3924,N_319);
nand U7719 (N_7719,N_5580,N_4278);
nand U7720 (N_7720,N_4208,N_3463);
nor U7721 (N_7721,N_4011,N_4600);
and U7722 (N_7722,N_6077,N_5135);
nor U7723 (N_7723,N_2367,N_4758);
and U7724 (N_7724,N_5247,N_754);
nor U7725 (N_7725,N_782,N_30);
xor U7726 (N_7726,N_2724,N_5432);
and U7727 (N_7727,N_5653,N_1005);
or U7728 (N_7728,N_3584,N_5038);
xnor U7729 (N_7729,N_4030,N_4141);
and U7730 (N_7730,N_1088,N_2798);
or U7731 (N_7731,N_1587,N_739);
or U7732 (N_7732,N_4648,N_4137);
nand U7733 (N_7733,N_112,N_876);
or U7734 (N_7734,N_5665,N_1634);
or U7735 (N_7735,N_1052,N_2248);
nand U7736 (N_7736,N_4745,N_593);
or U7737 (N_7737,N_1449,N_1983);
or U7738 (N_7738,N_5712,N_792);
nor U7739 (N_7739,N_1336,N_2532);
nand U7740 (N_7740,N_1890,N_1347);
and U7741 (N_7741,N_1019,N_4498);
xnor U7742 (N_7742,N_5481,N_2047);
nor U7743 (N_7743,N_6211,N_4853);
or U7744 (N_7744,N_1277,N_2648);
nor U7745 (N_7745,N_1236,N_4124);
or U7746 (N_7746,N_950,N_1639);
xor U7747 (N_7747,N_5051,N_220);
nor U7748 (N_7748,N_3302,N_3572);
nor U7749 (N_7749,N_4527,N_639);
or U7750 (N_7750,N_135,N_2133);
nand U7751 (N_7751,N_4881,N_4085);
or U7752 (N_7752,N_572,N_543);
xnor U7753 (N_7753,N_1265,N_4710);
and U7754 (N_7754,N_1118,N_713);
nand U7755 (N_7755,N_2552,N_3785);
nor U7756 (N_7756,N_6105,N_3392);
or U7757 (N_7757,N_2593,N_5014);
and U7758 (N_7758,N_3944,N_5568);
or U7759 (N_7759,N_675,N_2424);
nor U7760 (N_7760,N_50,N_3920);
xor U7761 (N_7761,N_2771,N_3409);
and U7762 (N_7762,N_3382,N_2973);
xnor U7763 (N_7763,N_5016,N_2246);
nor U7764 (N_7764,N_5652,N_4143);
and U7765 (N_7765,N_4416,N_2276);
xor U7766 (N_7766,N_779,N_5562);
xor U7767 (N_7767,N_5806,N_4475);
or U7768 (N_7768,N_1086,N_286);
and U7769 (N_7769,N_1153,N_2927);
nor U7770 (N_7770,N_2572,N_233);
and U7771 (N_7771,N_2355,N_5805);
nand U7772 (N_7772,N_3757,N_3025);
nand U7773 (N_7773,N_5962,N_2102);
nand U7774 (N_7774,N_6187,N_3745);
xnor U7775 (N_7775,N_3135,N_4808);
and U7776 (N_7776,N_5546,N_4643);
nand U7777 (N_7777,N_2373,N_681);
and U7778 (N_7778,N_5577,N_3375);
and U7779 (N_7779,N_1768,N_3771);
xnor U7780 (N_7780,N_3554,N_2372);
and U7781 (N_7781,N_290,N_570);
nand U7782 (N_7782,N_5965,N_1312);
nor U7783 (N_7783,N_1345,N_4553);
nand U7784 (N_7784,N_4256,N_4117);
nand U7785 (N_7785,N_3333,N_2174);
and U7786 (N_7786,N_3547,N_18);
nand U7787 (N_7787,N_4456,N_2288);
nand U7788 (N_7788,N_4152,N_6017);
and U7789 (N_7789,N_4258,N_6026);
and U7790 (N_7790,N_244,N_785);
nor U7791 (N_7791,N_5298,N_2501);
nand U7792 (N_7792,N_1095,N_610);
or U7793 (N_7793,N_3415,N_5611);
nor U7794 (N_7794,N_4585,N_3406);
nand U7795 (N_7795,N_4855,N_4382);
or U7796 (N_7796,N_4345,N_4635);
nand U7797 (N_7797,N_4718,N_4646);
or U7798 (N_7798,N_1409,N_2001);
xor U7799 (N_7799,N_1555,N_5798);
nand U7800 (N_7800,N_2636,N_4322);
nand U7801 (N_7801,N_2014,N_4379);
xor U7802 (N_7802,N_5780,N_1546);
and U7803 (N_7803,N_1337,N_5914);
or U7804 (N_7804,N_2555,N_3881);
nor U7805 (N_7805,N_5070,N_91);
and U7806 (N_7806,N_3803,N_3051);
nand U7807 (N_7807,N_4212,N_3338);
and U7808 (N_7808,N_2170,N_4060);
xnor U7809 (N_7809,N_204,N_5744);
xnor U7810 (N_7810,N_3014,N_1385);
xor U7811 (N_7811,N_2006,N_4800);
nand U7812 (N_7812,N_1129,N_797);
xor U7813 (N_7813,N_2025,N_1607);
nor U7814 (N_7814,N_3642,N_6094);
nor U7815 (N_7815,N_2573,N_278);
or U7816 (N_7816,N_862,N_4400);
nand U7817 (N_7817,N_2098,N_1122);
and U7818 (N_7818,N_4933,N_4747);
nor U7819 (N_7819,N_4170,N_4817);
xor U7820 (N_7820,N_5396,N_69);
and U7821 (N_7821,N_4135,N_1100);
xnor U7822 (N_7822,N_2726,N_4264);
and U7823 (N_7823,N_4781,N_5852);
xor U7824 (N_7824,N_2738,N_5599);
nand U7825 (N_7825,N_5052,N_4155);
nor U7826 (N_7826,N_4377,N_2608);
nand U7827 (N_7827,N_1597,N_3434);
nor U7828 (N_7828,N_6012,N_3070);
and U7829 (N_7829,N_4905,N_740);
and U7830 (N_7830,N_4963,N_4423);
and U7831 (N_7831,N_3573,N_141);
and U7832 (N_7832,N_4965,N_1522);
or U7833 (N_7833,N_2366,N_1934);
nand U7834 (N_7834,N_4077,N_2275);
xnor U7835 (N_7835,N_3752,N_2769);
nor U7836 (N_7836,N_1699,N_3676);
xor U7837 (N_7837,N_3949,N_2411);
or U7838 (N_7838,N_4180,N_947);
and U7839 (N_7839,N_4888,N_856);
xnor U7840 (N_7840,N_804,N_3368);
and U7841 (N_7841,N_4464,N_5216);
or U7842 (N_7842,N_3916,N_297);
nand U7843 (N_7843,N_525,N_4272);
nand U7844 (N_7844,N_2380,N_2987);
nor U7845 (N_7845,N_3919,N_4712);
nand U7846 (N_7846,N_4875,N_2395);
or U7847 (N_7847,N_1189,N_1526);
nand U7848 (N_7848,N_4172,N_3939);
nand U7849 (N_7849,N_2913,N_1412);
and U7850 (N_7850,N_5341,N_376);
and U7851 (N_7851,N_5317,N_3408);
or U7852 (N_7852,N_4028,N_4854);
xnor U7853 (N_7853,N_2464,N_5009);
nand U7854 (N_7854,N_2221,N_620);
nor U7855 (N_7855,N_4069,N_2582);
xnor U7856 (N_7856,N_3853,N_385);
nand U7857 (N_7857,N_2048,N_3838);
xnor U7858 (N_7858,N_1281,N_29);
nand U7859 (N_7859,N_2590,N_44);
and U7860 (N_7860,N_4220,N_837);
or U7861 (N_7861,N_898,N_893);
xor U7862 (N_7862,N_3984,N_1282);
or U7863 (N_7863,N_597,N_1660);
nand U7864 (N_7864,N_1197,N_1663);
nand U7865 (N_7865,N_1382,N_2834);
and U7866 (N_7866,N_2764,N_5768);
nand U7867 (N_7867,N_267,N_1980);
or U7868 (N_7868,N_4255,N_2868);
nor U7869 (N_7869,N_5104,N_5989);
nor U7870 (N_7870,N_4913,N_5966);
xnor U7871 (N_7871,N_3389,N_762);
nand U7872 (N_7872,N_2466,N_628);
xor U7873 (N_7873,N_1693,N_2245);
nor U7874 (N_7874,N_4999,N_3696);
xor U7875 (N_7875,N_537,N_5745);
and U7876 (N_7876,N_1781,N_353);
xnor U7877 (N_7877,N_4530,N_806);
and U7878 (N_7878,N_5757,N_2120);
xor U7879 (N_7879,N_2920,N_74);
or U7880 (N_7880,N_2565,N_5132);
nor U7881 (N_7881,N_2369,N_5521);
xor U7882 (N_7882,N_4650,N_3698);
nand U7883 (N_7883,N_4975,N_5904);
nand U7884 (N_7884,N_1603,N_2713);
and U7885 (N_7885,N_5644,N_2165);
xnor U7886 (N_7886,N_2268,N_5766);
nand U7887 (N_7887,N_1270,N_148);
and U7888 (N_7888,N_2312,N_2242);
nor U7889 (N_7889,N_6173,N_5523);
and U7890 (N_7890,N_5403,N_1319);
nor U7891 (N_7891,N_661,N_3505);
and U7892 (N_7892,N_4478,N_4863);
and U7893 (N_7893,N_5097,N_3629);
and U7894 (N_7894,N_342,N_5179);
nor U7895 (N_7895,N_4317,N_132);
nor U7896 (N_7896,N_4428,N_3498);
and U7897 (N_7897,N_773,N_5794);
nor U7898 (N_7898,N_1561,N_475);
nor U7899 (N_7899,N_1378,N_6126);
xnor U7900 (N_7900,N_5156,N_2334);
or U7901 (N_7901,N_3848,N_3192);
nand U7902 (N_7902,N_6155,N_1787);
and U7903 (N_7903,N_5524,N_590);
or U7904 (N_7904,N_246,N_2546);
or U7905 (N_7905,N_1261,N_4273);
nor U7906 (N_7906,N_2507,N_4723);
or U7907 (N_7907,N_4820,N_5827);
xnor U7908 (N_7908,N_3941,N_6242);
nand U7909 (N_7909,N_2917,N_2070);
nor U7910 (N_7910,N_1509,N_1131);
xnor U7911 (N_7911,N_2259,N_5841);
xnor U7912 (N_7912,N_4441,N_1626);
nor U7913 (N_7913,N_5467,N_4979);
nand U7914 (N_7914,N_1604,N_2839);
and U7915 (N_7915,N_2633,N_5304);
nor U7916 (N_7916,N_3558,N_5010);
and U7917 (N_7917,N_3988,N_1504);
nand U7918 (N_7918,N_214,N_1288);
nor U7919 (N_7919,N_5585,N_3032);
and U7920 (N_7920,N_288,N_5716);
xnor U7921 (N_7921,N_997,N_3055);
nor U7922 (N_7922,N_90,N_3433);
or U7923 (N_7923,N_1564,N_2437);
nand U7924 (N_7924,N_2978,N_2416);
or U7925 (N_7925,N_1216,N_2902);
and U7926 (N_7926,N_4359,N_1589);
nand U7927 (N_7927,N_3865,N_1852);
and U7928 (N_7928,N_5656,N_1736);
or U7929 (N_7929,N_5358,N_5830);
nand U7930 (N_7930,N_3751,N_6029);
nor U7931 (N_7931,N_2551,N_4981);
and U7932 (N_7932,N_5158,N_2382);
nand U7933 (N_7933,N_2,N_1190);
nand U7934 (N_7934,N_3728,N_4536);
nor U7935 (N_7935,N_1963,N_1519);
or U7936 (N_7936,N_2703,N_6181);
or U7937 (N_7937,N_3670,N_4232);
or U7938 (N_7938,N_4671,N_1175);
and U7939 (N_7939,N_1499,N_3388);
nor U7940 (N_7940,N_718,N_6192);
nor U7941 (N_7941,N_2758,N_3923);
nor U7942 (N_7942,N_5029,N_3018);
nand U7943 (N_7943,N_3833,N_3664);
nor U7944 (N_7944,N_4593,N_1997);
and U7945 (N_7945,N_1620,N_2723);
nand U7946 (N_7946,N_4539,N_4690);
and U7947 (N_7947,N_6180,N_5571);
and U7948 (N_7948,N_2483,N_2562);
and U7949 (N_7949,N_3776,N_4872);
nand U7950 (N_7950,N_1758,N_383);
xnor U7951 (N_7951,N_1521,N_6183);
xor U7952 (N_7952,N_4804,N_79);
and U7953 (N_7953,N_2851,N_1859);
or U7954 (N_7954,N_3470,N_4110);
nand U7955 (N_7955,N_3643,N_4608);
nor U7956 (N_7956,N_4778,N_5031);
nand U7957 (N_7957,N_2998,N_3647);
or U7958 (N_7958,N_4645,N_1821);
or U7959 (N_7959,N_1158,N_3978);
xnor U7960 (N_7960,N_3510,N_365);
nand U7961 (N_7961,N_2290,N_5482);
xnor U7962 (N_7962,N_5198,N_2557);
and U7963 (N_7963,N_5242,N_4897);
xnor U7964 (N_7964,N_401,N_2909);
nand U7965 (N_7965,N_3741,N_2945);
xnor U7966 (N_7966,N_1733,N_1124);
xnor U7967 (N_7967,N_1964,N_2022);
nand U7968 (N_7968,N_333,N_1068);
xor U7969 (N_7969,N_4098,N_54);
and U7970 (N_7970,N_6060,N_2396);
nand U7971 (N_7971,N_2679,N_4101);
xnor U7972 (N_7972,N_2043,N_4556);
or U7973 (N_7973,N_5370,N_2696);
or U7974 (N_7974,N_2890,N_3342);
and U7975 (N_7975,N_4254,N_2575);
nand U7976 (N_7976,N_2702,N_1886);
nand U7977 (N_7977,N_2111,N_1263);
nor U7978 (N_7978,N_4633,N_2121);
nor U7979 (N_7979,N_5133,N_2370);
and U7980 (N_7980,N_5429,N_1788);
nor U7981 (N_7981,N_1953,N_2210);
nor U7982 (N_7982,N_2537,N_630);
xnor U7983 (N_7983,N_1848,N_2999);
nand U7984 (N_7984,N_3155,N_3780);
nand U7985 (N_7985,N_177,N_1850);
nand U7986 (N_7986,N_602,N_545);
or U7987 (N_7987,N_4528,N_633);
xor U7988 (N_7988,N_4502,N_4448);
nand U7989 (N_7989,N_4507,N_3058);
and U7990 (N_7990,N_6149,N_3286);
nor U7991 (N_7991,N_5054,N_5784);
or U7992 (N_7992,N_6020,N_1862);
xor U7993 (N_7993,N_989,N_5108);
and U7994 (N_7994,N_614,N_1599);
nor U7995 (N_7995,N_850,N_2185);
nor U7996 (N_7996,N_4575,N_626);
xor U7997 (N_7997,N_5701,N_1759);
or U7998 (N_7998,N_4632,N_1295);
or U7999 (N_7999,N_3439,N_1488);
and U8000 (N_8000,N_3123,N_3281);
xnor U8001 (N_8001,N_2606,N_1002);
and U8002 (N_8002,N_643,N_5765);
nand U8003 (N_8003,N_2874,N_1641);
nor U8004 (N_8004,N_1240,N_4997);
xor U8005 (N_8005,N_1461,N_1899);
or U8006 (N_8006,N_1956,N_3663);
xor U8007 (N_8007,N_4569,N_4435);
xnor U8008 (N_8008,N_4533,N_3697);
or U8009 (N_8009,N_1196,N_4631);
nor U8010 (N_8010,N_3985,N_494);
nor U8011 (N_8011,N_1618,N_3249);
nand U8012 (N_8012,N_5615,N_4053);
nor U8013 (N_8013,N_343,N_908);
xnor U8014 (N_8014,N_3313,N_2057);
nand U8015 (N_8015,N_4621,N_2691);
xor U8016 (N_8016,N_4367,N_5343);
nor U8017 (N_8017,N_768,N_262);
and U8018 (N_8018,N_881,N_4425);
nor U8019 (N_8019,N_6178,N_3990);
or U8020 (N_8020,N_5423,N_4678);
nand U8021 (N_8021,N_1073,N_5302);
xor U8022 (N_8022,N_4862,N_4564);
nand U8023 (N_8023,N_2258,N_120);
and U8024 (N_8024,N_5250,N_1222);
xor U8025 (N_8025,N_2430,N_1508);
and U8026 (N_8026,N_2550,N_2013);
or U8027 (N_8027,N_4275,N_851);
or U8028 (N_8028,N_2880,N_1071);
and U8029 (N_8029,N_5212,N_3348);
and U8030 (N_8030,N_5191,N_5154);
and U8031 (N_8031,N_1948,N_1717);
nor U8032 (N_8032,N_3250,N_459);
and U8033 (N_8033,N_1878,N_410);
and U8034 (N_8034,N_1000,N_3114);
and U8035 (N_8035,N_1370,N_5925);
xnor U8036 (N_8036,N_5737,N_2398);
nor U8037 (N_8037,N_1967,N_2035);
xnor U8038 (N_8038,N_4115,N_1415);
or U8039 (N_8039,N_1707,N_3726);
or U8040 (N_8040,N_6014,N_2639);
xnor U8041 (N_8041,N_489,N_5823);
xnor U8042 (N_8042,N_1256,N_1818);
xor U8043 (N_8043,N_5504,N_891);
nor U8044 (N_8044,N_5860,N_765);
xor U8045 (N_8045,N_4350,N_4238);
nor U8046 (N_8046,N_1421,N_549);
nor U8047 (N_8047,N_2873,N_3976);
nand U8048 (N_8048,N_4890,N_1772);
xnor U8049 (N_8049,N_2060,N_1107);
and U8050 (N_8050,N_3151,N_4901);
nor U8051 (N_8051,N_3822,N_5542);
xnor U8052 (N_8052,N_1710,N_5137);
and U8053 (N_8053,N_1027,N_4551);
nor U8054 (N_8054,N_2553,N_3904);
or U8055 (N_8055,N_6066,N_6033);
xor U8056 (N_8056,N_2513,N_3082);
nand U8057 (N_8057,N_4794,N_449);
nor U8058 (N_8058,N_5753,N_586);
nand U8059 (N_8059,N_5311,N_5459);
nand U8060 (N_8060,N_4189,N_13);
nor U8061 (N_8061,N_2117,N_2958);
or U8062 (N_8062,N_3193,N_122);
nor U8063 (N_8063,N_3577,N_3963);
or U8064 (N_8064,N_6243,N_3064);
and U8065 (N_8065,N_71,N_1588);
nor U8066 (N_8066,N_726,N_25);
nor U8067 (N_8067,N_676,N_5246);
or U8068 (N_8068,N_4916,N_3898);
nor U8069 (N_8069,N_149,N_5264);
and U8070 (N_8070,N_3042,N_5988);
nand U8071 (N_8071,N_1935,N_5586);
and U8072 (N_8072,N_4229,N_2114);
nor U8073 (N_8073,N_4409,N_4035);
or U8074 (N_8074,N_6245,N_4218);
and U8075 (N_8075,N_1149,N_4136);
nor U8076 (N_8076,N_1592,N_4701);
and U8077 (N_8077,N_5854,N_5103);
nor U8078 (N_8078,N_2585,N_3545);
nor U8079 (N_8079,N_61,N_5603);
xor U8080 (N_8080,N_5623,N_3866);
or U8081 (N_8081,N_5214,N_35);
nor U8082 (N_8082,N_3452,N_1807);
and U8083 (N_8083,N_2975,N_649);
nor U8084 (N_8084,N_4542,N_5872);
nand U8085 (N_8085,N_5881,N_5408);
xor U8086 (N_8086,N_2661,N_749);
nand U8087 (N_8087,N_4297,N_5829);
nand U8088 (N_8088,N_2732,N_3133);
and U8089 (N_8089,N_3756,N_2785);
and U8090 (N_8090,N_605,N_4660);
nor U8091 (N_8091,N_70,N_5821);
and U8092 (N_8092,N_894,N_2064);
nor U8093 (N_8093,N_4205,N_3420);
nand U8094 (N_8094,N_5693,N_5205);
nand U8095 (N_8095,N_3951,N_4670);
nor U8096 (N_8096,N_1622,N_2461);
and U8097 (N_8097,N_5271,N_1371);
nand U8098 (N_8098,N_5067,N_1518);
and U8099 (N_8099,N_2251,N_2694);
nor U8100 (N_8100,N_2796,N_2391);
nor U8101 (N_8101,N_199,N_4779);
or U8102 (N_8102,N_180,N_4439);
nand U8103 (N_8103,N_2925,N_5443);
xnor U8104 (N_8104,N_4994,N_2137);
or U8105 (N_8105,N_2240,N_5015);
or U8106 (N_8106,N_2482,N_4204);
nor U8107 (N_8107,N_1776,N_5967);
nand U8108 (N_8108,N_2445,N_3421);
and U8109 (N_8109,N_1425,N_4430);
xor U8110 (N_8110,N_6134,N_4914);
nor U8111 (N_8111,N_2919,N_5124);
nand U8112 (N_8112,N_2930,N_4452);
nand U8113 (N_8113,N_3130,N_5533);
or U8114 (N_8114,N_3627,N_2898);
and U8115 (N_8115,N_75,N_556);
nor U8116 (N_8116,N_2307,N_2556);
nand U8117 (N_8117,N_6027,N_2879);
nor U8118 (N_8118,N_3157,N_4164);
xnor U8119 (N_8119,N_2154,N_272);
nand U8120 (N_8120,N_2311,N_3295);
nand U8121 (N_8121,N_5147,N_394);
xor U8122 (N_8122,N_3351,N_4227);
and U8123 (N_8123,N_3678,N_2371);
nor U8124 (N_8124,N_5217,N_701);
and U8125 (N_8125,N_2353,N_5028);
xnor U8126 (N_8126,N_26,N_4520);
xnor U8127 (N_8127,N_1204,N_2096);
nand U8128 (N_8128,N_6224,N_709);
nor U8129 (N_8129,N_5427,N_5998);
nor U8130 (N_8130,N_3801,N_3530);
nor U8131 (N_8131,N_5053,N_3773);
nor U8132 (N_8132,N_4866,N_5864);
nor U8133 (N_8133,N_2625,N_2965);
xnor U8134 (N_8134,N_3968,N_270);
nor U8135 (N_8135,N_3024,N_3457);
nor U8136 (N_8136,N_4925,N_3468);
nor U8137 (N_8137,N_2286,N_6244);
xnor U8138 (N_8138,N_5758,N_5906);
nand U8139 (N_8139,N_1958,N_5968);
xor U8140 (N_8140,N_4105,N_3595);
xnor U8141 (N_8141,N_5826,N_4772);
xnor U8142 (N_8142,N_2077,N_5954);
nor U8143 (N_8143,N_436,N_5380);
nor U8144 (N_8144,N_430,N_6248);
nand U8145 (N_8145,N_4148,N_2847);
or U8146 (N_8146,N_4455,N_4870);
nor U8147 (N_8147,N_3507,N_2097);
xor U8148 (N_8148,N_3725,N_2390);
nor U8149 (N_8149,N_4311,N_4807);
nand U8150 (N_8150,N_1670,N_2810);
or U8151 (N_8151,N_810,N_6087);
nand U8152 (N_8152,N_3060,N_835);
or U8153 (N_8153,N_3559,N_3809);
and U8154 (N_8154,N_4565,N_2330);
or U8155 (N_8155,N_4093,N_5383);
nand U8156 (N_8156,N_2580,N_5748);
nor U8157 (N_8157,N_4525,N_5148);
nor U8158 (N_8158,N_775,N_569);
or U8159 (N_8159,N_2148,N_6196);
nor U8160 (N_8160,N_2226,N_3294);
nor U8161 (N_8161,N_4036,N_1188);
and U8162 (N_8162,N_5706,N_5424);
xnor U8163 (N_8163,N_2397,N_3306);
nand U8164 (N_8164,N_5945,N_2159);
and U8165 (N_8165,N_3549,N_3226);
and U8166 (N_8166,N_1655,N_3651);
and U8167 (N_8167,N_486,N_1629);
or U8168 (N_8168,N_97,N_5898);
xor U8169 (N_8169,N_4308,N_6238);
xnor U8170 (N_8170,N_6021,N_2863);
nand U8171 (N_8171,N_2442,N_2459);
or U8172 (N_8172,N_281,N_5916);
and U8173 (N_8173,N_3349,N_2046);
or U8174 (N_8174,N_2304,N_671);
xor U8175 (N_8175,N_5262,N_1757);
nand U8176 (N_8176,N_2233,N_4578);
or U8177 (N_8177,N_41,N_5686);
xnor U8178 (N_8178,N_4535,N_3080);
xor U8179 (N_8179,N_4072,N_3910);
xnor U8180 (N_8180,N_5963,N_6220);
or U8181 (N_8181,N_2045,N_3310);
nand U8182 (N_8182,N_741,N_2458);
nor U8183 (N_8183,N_6072,N_4202);
xnor U8184 (N_8184,N_5310,N_3534);
nor U8185 (N_8185,N_973,N_5167);
and U8186 (N_8186,N_5792,N_783);
or U8187 (N_8187,N_2949,N_83);
or U8188 (N_8188,N_884,N_2535);
xnor U8189 (N_8189,N_76,N_4082);
and U8190 (N_8190,N_5193,N_1853);
and U8191 (N_8191,N_442,N_1950);
or U8192 (N_8192,N_5089,N_4638);
nor U8193 (N_8193,N_1959,N_380);
or U8194 (N_8194,N_3597,N_2277);
nor U8195 (N_8195,N_4896,N_1470);
nor U8196 (N_8196,N_6165,N_4986);
or U8197 (N_8197,N_2106,N_4780);
and U8198 (N_8198,N_5061,N_6194);
nor U8199 (N_8199,N_5269,N_4375);
or U8200 (N_8200,N_3499,N_398);
or U8201 (N_8201,N_6031,N_3767);
nand U8202 (N_8202,N_2503,N_6225);
nand U8203 (N_8203,N_1214,N_2671);
and U8204 (N_8204,N_3440,N_2105);
nand U8205 (N_8205,N_3185,N_4267);
nand U8206 (N_8206,N_4242,N_136);
and U8207 (N_8207,N_760,N_5388);
nand U8208 (N_8208,N_46,N_4673);
nand U8209 (N_8209,N_2806,N_5723);
nand U8210 (N_8210,N_2730,N_6076);
nand U8211 (N_8211,N_5451,N_497);
nand U8212 (N_8212,N_5516,N_3402);
or U8213 (N_8213,N_5522,N_2972);
or U8214 (N_8214,N_1809,N_2568);
nor U8215 (N_8215,N_5023,N_346);
and U8216 (N_8216,N_4465,N_5688);
nand U8217 (N_8217,N_561,N_2729);
or U8218 (N_8218,N_192,N_3178);
nand U8219 (N_8219,N_1013,N_885);
or U8220 (N_8220,N_2928,N_5397);
xnor U8221 (N_8221,N_477,N_4225);
xor U8222 (N_8222,N_470,N_329);
or U8223 (N_8223,N_2914,N_1092);
nor U8224 (N_8224,N_548,N_2795);
and U8225 (N_8225,N_3166,N_2520);
nand U8226 (N_8226,N_3246,N_5116);
nor U8227 (N_8227,N_1989,N_2107);
nand U8228 (N_8228,N_2234,N_450);
xor U8229 (N_8229,N_2162,N_4649);
and U8230 (N_8230,N_4958,N_1898);
nand U8231 (N_8231,N_3936,N_3115);
nor U8232 (N_8232,N_928,N_5843);
nor U8233 (N_8233,N_5876,N_4213);
and U8234 (N_8234,N_6221,N_4500);
xnor U8235 (N_8235,N_2521,N_2052);
nand U8236 (N_8236,N_5911,N_5700);
xor U8237 (N_8237,N_5099,N_3451);
xnor U8238 (N_8238,N_606,N_3426);
or U8239 (N_8239,N_1547,N_942);
nand U8240 (N_8240,N_2751,N_2564);
or U8241 (N_8241,N_2206,N_2595);
nor U8242 (N_8242,N_5990,N_2660);
and U8243 (N_8243,N_1719,N_5435);
nor U8244 (N_8244,N_341,N_4018);
xor U8245 (N_8245,N_3931,N_4296);
nor U8246 (N_8246,N_4662,N_5949);
and U8247 (N_8247,N_382,N_3479);
and U8248 (N_8248,N_2980,N_5093);
or U8249 (N_8249,N_4032,N_1174);
nand U8250 (N_8250,N_3071,N_4168);
nor U8251 (N_8251,N_2517,N_3354);
or U8252 (N_8252,N_5460,N_424);
nor U8253 (N_8253,N_1598,N_1627);
nand U8254 (N_8254,N_3345,N_4617);
or U8255 (N_8255,N_2076,N_1871);
nand U8256 (N_8256,N_1114,N_3472);
nand U8257 (N_8257,N_4967,N_663);
nor U8258 (N_8258,N_3000,N_5000);
and U8259 (N_8259,N_1274,N_2941);
nor U8260 (N_8260,N_5547,N_4504);
nand U8261 (N_8261,N_5928,N_1455);
or U8262 (N_8262,N_260,N_2409);
xor U8263 (N_8263,N_1121,N_2956);
and U8264 (N_8264,N_4526,N_3649);
xor U8265 (N_8265,N_1575,N_5690);
or U8266 (N_8266,N_951,N_2739);
and U8267 (N_8267,N_3107,N_4984);
and U8268 (N_8268,N_84,N_266);
nor U8269 (N_8269,N_3928,N_4924);
or U8270 (N_8270,N_116,N_390);
or U8271 (N_8271,N_824,N_1045);
nand U8272 (N_8272,N_2190,N_3807);
nand U8273 (N_8273,N_5176,N_5884);
xor U8274 (N_8274,N_1298,N_5937);
nor U8275 (N_8275,N_2420,N_4402);
or U8276 (N_8276,N_1074,N_1525);
nand U8277 (N_8277,N_317,N_5237);
nor U8278 (N_8278,N_3969,N_3514);
nor U8279 (N_8279,N_5957,N_1201);
or U8280 (N_8280,N_4484,N_636);
nand U8281 (N_8281,N_2539,N_1450);
and U8282 (N_8282,N_4128,N_4832);
and U8283 (N_8283,N_5588,N_1708);
nand U8284 (N_8284,N_5797,N_3049);
nand U8285 (N_8285,N_3890,N_3736);
and U8286 (N_8286,N_3669,N_4111);
or U8287 (N_8287,N_1794,N_5948);
nor U8288 (N_8288,N_615,N_3706);
nor U8289 (N_8289,N_900,N_4078);
nor U8290 (N_8290,N_4814,N_5421);
nor U8291 (N_8291,N_541,N_1755);
xnor U8292 (N_8292,N_1895,N_4156);
xnor U8293 (N_8293,N_3274,N_3365);
nor U8294 (N_8294,N_201,N_879);
nor U8295 (N_8295,N_4666,N_5139);
or U8296 (N_8296,N_3012,N_5058);
nor U8297 (N_8297,N_1187,N_3373);
nand U8298 (N_8298,N_784,N_3121);
nand U8299 (N_8299,N_2939,N_166);
nor U8300 (N_8300,N_3671,N_4894);
or U8301 (N_8301,N_3480,N_3574);
nor U8302 (N_8302,N_1713,N_2620);
nor U8303 (N_8303,N_2364,N_1735);
nor U8304 (N_8304,N_1245,N_1730);
or U8305 (N_8305,N_1015,N_2079);
nor U8306 (N_8306,N_5721,N_5556);
xnor U8307 (N_8307,N_2252,N_2781);
nand U8308 (N_8308,N_3331,N_2626);
nor U8309 (N_8309,N_3317,N_138);
nor U8310 (N_8310,N_6117,N_5734);
nand U8311 (N_8311,N_1792,N_4043);
nand U8312 (N_8312,N_6142,N_2313);
xnor U8313 (N_8313,N_2181,N_3413);
nor U8314 (N_8314,N_5366,N_3301);
nor U8315 (N_8315,N_5390,N_4729);
or U8316 (N_8316,N_5616,N_1356);
or U8317 (N_8317,N_4485,N_1091);
nand U8318 (N_8318,N_6236,N_5249);
and U8319 (N_8319,N_4789,N_2534);
xor U8320 (N_8320,N_3859,N_1405);
nor U8321 (N_8321,N_721,N_4763);
or U8322 (N_8322,N_4574,N_234);
or U8323 (N_8323,N_2289,N_2910);
or U8324 (N_8324,N_2838,N_1752);
xor U8325 (N_8325,N_3398,N_99);
and U8326 (N_8326,N_875,N_3216);
and U8327 (N_8327,N_5375,N_5359);
nor U8328 (N_8328,N_2265,N_6050);
xnor U8329 (N_8329,N_1137,N_1227);
and U8330 (N_8330,N_4547,N_3203);
nand U8331 (N_8331,N_5679,N_5367);
nor U8332 (N_8332,N_3363,N_1321);
xor U8333 (N_8333,N_2800,N_1548);
or U8334 (N_8334,N_1059,N_4356);
and U8335 (N_8335,N_3746,N_327);
nor U8336 (N_8336,N_5634,N_1891);
or U8337 (N_8337,N_5754,N_1067);
xnor U8338 (N_8338,N_2209,N_5907);
or U8339 (N_8339,N_1896,N_1946);
nor U8340 (N_8340,N_5842,N_5438);
nand U8341 (N_8341,N_3713,N_1789);
or U8342 (N_8342,N_1427,N_3335);
and U8343 (N_8343,N_460,N_1340);
and U8344 (N_8344,N_5708,N_3965);
or U8345 (N_8345,N_1309,N_5324);
or U8346 (N_8346,N_1242,N_5573);
nor U8347 (N_8347,N_5755,N_4031);
and U8348 (N_8348,N_1885,N_5256);
xnor U8349 (N_8349,N_4508,N_5440);
nand U8350 (N_8350,N_1326,N_2146);
nand U8351 (N_8351,N_5042,N_5558);
or U8352 (N_8352,N_2341,N_6166);
xor U8353 (N_8353,N_4354,N_2599);
or U8354 (N_8354,N_27,N_4803);
xor U8355 (N_8355,N_2962,N_1631);
nand U8356 (N_8356,N_5294,N_3608);
or U8357 (N_8357,N_4355,N_5505);
nand U8358 (N_8358,N_2141,N_12);
and U8359 (N_8359,N_1402,N_1042);
or U8360 (N_8360,N_3749,N_1436);
nand U8361 (N_8361,N_4895,N_2837);
xor U8362 (N_8362,N_6052,N_2935);
xor U8363 (N_8363,N_5401,N_6179);
nand U8364 (N_8364,N_3347,N_3126);
xor U8365 (N_8365,N_4559,N_846);
nand U8366 (N_8366,N_422,N_4420);
nor U8367 (N_8367,N_659,N_4277);
xnor U8368 (N_8368,N_913,N_5601);
or U8369 (N_8369,N_3362,N_3583);
nor U8370 (N_8370,N_5621,N_5292);
or U8371 (N_8371,N_359,N_1828);
and U8372 (N_8372,N_349,N_641);
nand U8373 (N_8373,N_4353,N_1162);
nor U8374 (N_8374,N_3909,N_4592);
and U8375 (N_8375,N_3614,N_598);
and U8376 (N_8376,N_4197,N_2439);
nand U8377 (N_8377,N_533,N_858);
nor U8378 (N_8378,N_5938,N_3567);
xor U8379 (N_8379,N_1554,N_4935);
nor U8380 (N_8380,N_438,N_2029);
or U8381 (N_8381,N_4919,N_563);
or U8382 (N_8382,N_457,N_3578);
or U8383 (N_8383,N_2316,N_5192);
nand U8384 (N_8384,N_4606,N_4653);
nand U8385 (N_8385,N_321,N_3097);
and U8386 (N_8386,N_182,N_386);
xor U8387 (N_8387,N_4217,N_565);
nand U8388 (N_8388,N_931,N_820);
nand U8389 (N_8389,N_657,N_3962);
nand U8390 (N_8390,N_3134,N_3356);
and U8391 (N_8391,N_2755,N_5077);
and U8392 (N_8392,N_251,N_3977);
xor U8393 (N_8393,N_4503,N_5275);
or U8394 (N_8394,N_3305,N_2499);
nand U8395 (N_8395,N_4186,N_2315);
xnor U8396 (N_8396,N_4964,N_2619);
nor U8397 (N_8397,N_1279,N_292);
or U8398 (N_8398,N_4436,N_312);
nand U8399 (N_8399,N_3520,N_3827);
xor U8400 (N_8400,N_3108,N_1094);
nand U8401 (N_8401,N_604,N_4582);
nor U8402 (N_8402,N_3531,N_2903);
and U8403 (N_8403,N_3116,N_5540);
nor U8404 (N_8404,N_1023,N_3325);
nand U8405 (N_8405,N_530,N_3291);
nor U8406 (N_8406,N_4050,N_296);
or U8407 (N_8407,N_4228,N_6057);
nand U8408 (N_8408,N_4676,N_945);
nor U8409 (N_8409,N_3376,N_5779);
nor U8410 (N_8410,N_377,N_3029);
and U8411 (N_8411,N_5483,N_1048);
xnor U8412 (N_8412,N_5910,N_5595);
and U8413 (N_8413,N_4532,N_5391);
nand U8414 (N_8414,N_3062,N_1369);
or U8415 (N_8415,N_2167,N_5461);
xnor U8416 (N_8416,N_2852,N_3823);
or U8417 (N_8417,N_2757,N_14);
nand U8418 (N_8418,N_3996,N_4330);
and U8419 (N_8419,N_3981,N_2576);
and U8420 (N_8420,N_5555,N_3544);
or U8421 (N_8421,N_3948,N_5277);
and U8422 (N_8422,N_702,N_4957);
or U8423 (N_8423,N_1647,N_5027);
or U8424 (N_8424,N_2401,N_4939);
xnor U8425 (N_8425,N_5520,N_2647);
nor U8426 (N_8426,N_5127,N_5337);
nand U8427 (N_8427,N_1229,N_2092);
nand U8428 (N_8428,N_3145,N_456);
nor U8429 (N_8429,N_2843,N_179);
xnor U8430 (N_8430,N_677,N_6000);
nor U8431 (N_8431,N_4065,N_1938);
and U8432 (N_8432,N_836,N_5908);
or U8433 (N_8433,N_1649,N_414);
and U8434 (N_8434,N_523,N_6058);
nand U8435 (N_8435,N_3397,N_5961);
nor U8436 (N_8436,N_5741,N_2710);
nand U8437 (N_8437,N_4004,N_1112);
xnor U8438 (N_8438,N_2815,N_1167);
nand U8439 (N_8439,N_4668,N_4624);
nor U8440 (N_8440,N_5181,N_5786);
xor U8441 (N_8441,N_5900,N_1740);
or U8442 (N_8442,N_1636,N_788);
nor U8443 (N_8443,N_3469,N_2093);
nor U8444 (N_8444,N_4138,N_4656);
nand U8445 (N_8445,N_1393,N_1212);
xnor U8446 (N_8446,N_2342,N_4390);
and U8447 (N_8447,N_3444,N_1856);
or U8448 (N_8448,N_5151,N_2491);
xor U8449 (N_8449,N_1008,N_1423);
xor U8450 (N_8450,N_1099,N_5339);
xnor U8451 (N_8451,N_1079,N_3582);
nand U8452 (N_8452,N_4898,N_651);
nor U8453 (N_8453,N_1709,N_6206);
xor U8454 (N_8454,N_5349,N_3533);
and U8455 (N_8455,N_1384,N_203);
and U8456 (N_8456,N_5811,N_3695);
nand U8457 (N_8457,N_5702,N_6097);
nand U8458 (N_8458,N_1296,N_693);
nor U8459 (N_8459,N_2197,N_752);
and U8460 (N_8460,N_6159,N_1029);
and U8461 (N_8461,N_1562,N_6118);
and U8462 (N_8462,N_4776,N_4798);
and U8463 (N_8463,N_487,N_1473);
and U8464 (N_8464,N_3681,N_547);
and U8465 (N_8465,N_4325,N_3237);
nand U8466 (N_8466,N_2421,N_3377);
nor U8467 (N_8467,N_248,N_4357);
xnor U8468 (N_8468,N_5682,N_1054);
nand U8469 (N_8469,N_1688,N_4303);
and U8470 (N_8470,N_554,N_2861);
and U8471 (N_8471,N_6056,N_5720);
xnor U8472 (N_8472,N_5814,N_781);
or U8473 (N_8473,N_5075,N_3561);
or U8474 (N_8474,N_5909,N_2906);
or U8475 (N_8475,N_87,N_587);
or U8476 (N_8476,N_1156,N_3876);
xnor U8477 (N_8477,N_2241,N_4921);
xor U8478 (N_8478,N_1798,N_3600);
nor U8479 (N_8479,N_1454,N_4013);
and U8480 (N_8480,N_5553,N_1494);
xnor U8481 (N_8481,N_4364,N_6079);
nor U8482 (N_8482,N_5332,N_4861);
nand U8483 (N_8483,N_2509,N_2971);
and U8484 (N_8484,N_619,N_845);
nand U8485 (N_8485,N_4696,N_813);
and U8486 (N_8486,N_717,N_4167);
xor U8487 (N_8487,N_1482,N_708);
and U8488 (N_8488,N_2995,N_2028);
nand U8489 (N_8489,N_2650,N_5314);
nand U8490 (N_8490,N_2609,N_939);
nor U8491 (N_8491,N_6055,N_2854);
and U8492 (N_8492,N_397,N_2140);
nor U8493 (N_8493,N_1430,N_345);
or U8494 (N_8494,N_613,N_5638);
and U8495 (N_8495,N_960,N_3419);
nand U8496 (N_8496,N_4823,N_566);
or U8497 (N_8497,N_4579,N_467);
and U8498 (N_8498,N_2269,N_4263);
nand U8499 (N_8499,N_4460,N_391);
xnor U8500 (N_8500,N_978,N_2742);
nand U8501 (N_8501,N_1642,N_815);
nor U8502 (N_8502,N_6122,N_3593);
or U8503 (N_8503,N_1417,N_161);
nor U8504 (N_8504,N_4580,N_1863);
or U8505 (N_8505,N_4956,N_1872);
and U8506 (N_8506,N_5970,N_2476);
nand U8507 (N_8507,N_1109,N_5474);
and U8508 (N_8508,N_331,N_1433);
and U8509 (N_8509,N_1199,N_1936);
nand U8510 (N_8510,N_3816,N_5825);
xor U8511 (N_8511,N_756,N_3160);
xnor U8512 (N_8512,N_904,N_793);
nor U8513 (N_8513,N_250,N_5265);
nand U8514 (N_8514,N_6075,N_3255);
nor U8515 (N_8515,N_5609,N_1697);
or U8516 (N_8516,N_4917,N_2301);
nand U8517 (N_8517,N_5646,N_2712);
nand U8518 (N_8518,N_2214,N_2666);
xnor U8519 (N_8519,N_5412,N_2067);
or U8520 (N_8520,N_2722,N_440);
and U8521 (N_8521,N_3120,N_4605);
xor U8522 (N_8522,N_4775,N_3438);
or U8523 (N_8523,N_1926,N_2545);
and U8524 (N_8524,N_5971,N_3711);
or U8525 (N_8525,N_4442,N_6025);
nor U8526 (N_8526,N_5141,N_2811);
xnor U8527 (N_8527,N_2083,N_2457);
xor U8528 (N_8528,N_4469,N_360);
nand U8529 (N_8529,N_1177,N_3010);
nor U8530 (N_8530,N_2692,N_2789);
nor U8531 (N_8531,N_3755,N_2112);
or U8532 (N_8532,N_2548,N_4481);
xnor U8533 (N_8533,N_1567,N_1271);
nand U8534 (N_8534,N_1703,N_5636);
nor U8535 (N_8535,N_3557,N_2195);
nor U8536 (N_8536,N_5789,N_2708);
or U8537 (N_8537,N_1813,N_1117);
xor U8538 (N_8538,N_5810,N_1495);
xnor U8539 (N_8539,N_3023,N_4883);
nand U8540 (N_8540,N_3502,N_1691);
and U8541 (N_8541,N_1484,N_1249);
nor U8542 (N_8542,N_3521,N_183);
and U8543 (N_8543,N_1306,N_2926);
nand U8544 (N_8544,N_3729,N_1351);
nand U8545 (N_8545,N_1715,N_5499);
nand U8546 (N_8546,N_3606,N_4693);
or U8547 (N_8547,N_5248,N_2654);
nor U8548 (N_8548,N_2220,N_2239);
xnor U8549 (N_8549,N_1463,N_4607);
xnor U8550 (N_8550,N_5241,N_3775);
and U8551 (N_8551,N_1968,N_2490);
nor U8552 (N_8552,N_3164,N_1767);
xor U8553 (N_8553,N_4289,N_4206);
xnor U8554 (N_8554,N_55,N_5959);
or U8555 (N_8555,N_2026,N_2462);
xor U8556 (N_8556,N_5100,N_1826);
or U8557 (N_8557,N_2500,N_3458);
xor U8558 (N_8558,N_1364,N_690);
and U8559 (N_8559,N_4543,N_2989);
and U8560 (N_8560,N_5371,N_1552);
and U8561 (N_8561,N_2994,N_4679);
xor U8562 (N_8562,N_110,N_4169);
xor U8563 (N_8563,N_3350,N_6036);
xnor U8564 (N_8564,N_1161,N_3843);
nor U8565 (N_8565,N_49,N_936);
xor U8566 (N_8566,N_1154,N_5130);
xor U8567 (N_8567,N_4068,N_2997);
or U8568 (N_8568,N_2675,N_4618);
xor U8569 (N_8569,N_3692,N_176);
and U8570 (N_8570,N_3401,N_2526);
xor U8571 (N_8571,N_144,N_3564);
and U8572 (N_8572,N_206,N_4774);
nor U8573 (N_8573,N_3550,N_2855);
or U8574 (N_8574,N_1182,N_5710);
and U8575 (N_8575,N_3431,N_1210);
or U8576 (N_8576,N_2684,N_4001);
nand U8577 (N_8577,N_3243,N_1571);
and U8578 (N_8578,N_151,N_573);
xor U8579 (N_8579,N_4459,N_3986);
nand U8580 (N_8580,N_1773,N_868);
and U8581 (N_8581,N_1684,N_2498);
and U8582 (N_8582,N_6037,N_5722);
xnor U8583 (N_8583,N_277,N_119);
and U8584 (N_8584,N_98,N_6172);
or U8585 (N_8585,N_445,N_4599);
and U8586 (N_8586,N_3159,N_4385);
xor U8587 (N_8587,N_2344,N_1877);
xor U8588 (N_8588,N_5987,N_5394);
and U8589 (N_8589,N_5287,N_3263);
nor U8590 (N_8590,N_4411,N_1966);
nand U8591 (N_8591,N_1127,N_1952);
nand U8592 (N_8592,N_2283,N_944);
nor U8593 (N_8593,N_1342,N_1727);
nand U8594 (N_8594,N_3799,N_2263);
or U8595 (N_8595,N_2343,N_1506);
nand U8596 (N_8596,N_2418,N_3846);
nor U8597 (N_8597,N_918,N_1390);
nand U8598 (N_8598,N_1238,N_4989);
xor U8599 (N_8599,N_2652,N_5724);
nand U8600 (N_8600,N_5844,N_3813);
nand U8601 (N_8601,N_4320,N_4634);
xnor U8602 (N_8602,N_59,N_917);
nor U8603 (N_8603,N_1355,N_4253);
or U8604 (N_8604,N_3768,N_1774);
nor U8605 (N_8605,N_4114,N_5026);
or U8606 (N_8606,N_1404,N_5492);
xnor U8607 (N_8607,N_4412,N_3104);
and U8608 (N_8608,N_5207,N_1181);
nor U8609 (N_8609,N_1053,N_4226);
and U8610 (N_8610,N_1974,N_1195);
xnor U8611 (N_8611,N_4410,N_232);
xor U8612 (N_8612,N_4826,N_5991);
xnor U8613 (N_8613,N_5718,N_3748);
and U8614 (N_8614,N_5079,N_3471);
nor U8615 (N_8615,N_4843,N_2073);
nor U8616 (N_8616,N_4071,N_672);
nand U8617 (N_8617,N_4130,N_3512);
nand U8618 (N_8618,N_1714,N_128);
nand U8619 (N_8619,N_5125,N_1331);
nand U8620 (N_8620,N_2228,N_5076);
or U8621 (N_8621,N_2635,N_2538);
and U8622 (N_8622,N_5096,N_1233);
or U8623 (N_8623,N_5259,N_1763);
xor U8624 (N_8624,N_3299,N_5853);
nor U8625 (N_8625,N_6015,N_4871);
and U8626 (N_8626,N_463,N_3276);
or U8627 (N_8627,N_2104,N_4597);
nand U8628 (N_8628,N_2784,N_5003);
nor U8629 (N_8629,N_3332,N_5885);
nand U8630 (N_8630,N_532,N_1741);
nor U8631 (N_8631,N_1920,N_328);
nand U8632 (N_8632,N_4795,N_4133);
or U8633 (N_8633,N_2992,N_1544);
and U8634 (N_8634,N_646,N_6171);
and U8635 (N_8635,N_3774,N_3360);
and U8636 (N_8636,N_3034,N_2883);
or U8637 (N_8637,N_510,N_524);
nor U8638 (N_8638,N_658,N_4473);
or U8639 (N_8639,N_1230,N_2792);
and U8640 (N_8640,N_621,N_2452);
xor U8641 (N_8641,N_5297,N_5512);
and U8642 (N_8642,N_4087,N_990);
and U8643 (N_8643,N_2069,N_4549);
nand U8644 (N_8644,N_4483,N_3892);
or U8645 (N_8645,N_3812,N_4799);
xor U8646 (N_8646,N_20,N_4116);
nor U8647 (N_8647,N_188,N_109);
or U8648 (N_8648,N_1262,N_1010);
and U8649 (N_8649,N_4980,N_1793);
or U8650 (N_8650,N_1906,N_3083);
and U8651 (N_8651,N_830,N_5569);
or U8652 (N_8652,N_5629,N_3662);
nand U8653 (N_8653,N_4835,N_755);
and U8654 (N_8654,N_3987,N_4623);
or U8655 (N_8655,N_4396,N_4877);
xor U8656 (N_8656,N_1200,N_1645);
and U8657 (N_8657,N_5650,N_1614);
xnor U8658 (N_8658,N_5727,N_5037);
nor U8659 (N_8659,N_1411,N_857);
or U8660 (N_8660,N_5160,N_2780);
nor U8661 (N_8661,N_5976,N_1033);
xor U8662 (N_8662,N_4880,N_5283);
nor U8663 (N_8663,N_4196,N_1441);
or U8664 (N_8664,N_1183,N_3085);
nand U8665 (N_8665,N_5655,N_2193);
or U8666 (N_8666,N_2826,N_425);
and U8667 (N_8667,N_4839,N_985);
and U8668 (N_8668,N_3038,N_384);
and U8669 (N_8669,N_137,N_3191);
or U8670 (N_8670,N_1583,N_5346);
nand U8671 (N_8671,N_283,N_4531);
or U8672 (N_8672,N_5022,N_1328);
xor U8673 (N_8673,N_5197,N_400);
and U8674 (N_8674,N_673,N_3202);
nor U8675 (N_8675,N_2892,N_175);
or U8676 (N_8676,N_5801,N_1357);
or U8677 (N_8677,N_4434,N_1376);
or U8678 (N_8678,N_2695,N_4529);
or U8679 (N_8679,N_6182,N_4323);
or U8680 (N_8680,N_3011,N_759);
nand U8681 (N_8681,N_4655,N_899);
or U8682 (N_8682,N_1847,N_5291);
xor U8683 (N_8683,N_1324,N_1489);
or U8684 (N_8684,N_1468,N_4298);
or U8685 (N_8685,N_1075,N_2187);
or U8686 (N_8686,N_3937,N_1132);
nand U8687 (N_8687,N_2817,N_1705);
and U8688 (N_8688,N_4281,N_1537);
xor U8689 (N_8689,N_3760,N_3087);
nand U8690 (N_8690,N_640,N_3672);
nor U8691 (N_8691,N_3737,N_4076);
nor U8692 (N_8692,N_1951,N_5381);
nor U8693 (N_8693,N_3372,N_230);
nor U8694 (N_8694,N_5759,N_1170);
nor U8695 (N_8695,N_1739,N_2504);
xor U8696 (N_8696,N_5610,N_5848);
xor U8697 (N_8697,N_3056,N_5767);
nand U8698 (N_8698,N_280,N_5436);
nand U8699 (N_8699,N_2303,N_3744);
and U8700 (N_8700,N_3006,N_2360);
or U8701 (N_8701,N_847,N_5322);
nand U8702 (N_8702,N_842,N_1679);
or U8703 (N_8703,N_4598,N_6213);
xnor U8704 (N_8704,N_4310,N_5170);
nor U8705 (N_8705,N_1742,N_439);
and U8706 (N_8706,N_5622,N_1887);
nand U8707 (N_8707,N_6110,N_4966);
xnor U8708 (N_8708,N_3874,N_2907);
and U8709 (N_8709,N_2714,N_5579);
xor U8710 (N_8710,N_4471,N_2744);
or U8711 (N_8711,N_3429,N_3654);
or U8712 (N_8712,N_1612,N_2727);
nor U8713 (N_8713,N_505,N_2436);
and U8714 (N_8714,N_1208,N_2264);
nand U8715 (N_8715,N_38,N_2841);
nand U8716 (N_8716,N_4594,N_3275);
nand U8717 (N_8717,N_612,N_2829);
and U8718 (N_8718,N_4007,N_2350);
and U8719 (N_8719,N_1662,N_4487);
nor U8720 (N_8720,N_3466,N_1226);
nand U8721 (N_8721,N_417,N_1018);
nor U8722 (N_8722,N_5115,N_2728);
nand U8723 (N_8723,N_429,N_2261);
nor U8724 (N_8724,N_4512,N_1287);
or U8725 (N_8725,N_389,N_958);
xor U8726 (N_8726,N_6222,N_1500);
nand U8727 (N_8727,N_1469,N_299);
nand U8728 (N_8728,N_174,N_3078);
and U8729 (N_8729,N_2760,N_3427);
nand U8730 (N_8730,N_1323,N_3110);
nand U8731 (N_8731,N_419,N_4697);
xor U8732 (N_8732,N_5252,N_5478);
xnor U8733 (N_8733,N_3334,N_4381);
xnor U8734 (N_8734,N_1050,N_5457);
nand U8735 (N_8735,N_4370,N_1698);
xnor U8736 (N_8736,N_3416,N_6042);
nand U8737 (N_8737,N_1677,N_1179);
and U8738 (N_8738,N_5671,N_6195);
or U8739 (N_8739,N_919,N_5752);
nor U8740 (N_8740,N_4418,N_5433);
xor U8741 (N_8741,N_1134,N_3278);
nor U8742 (N_8742,N_4784,N_77);
xnor U8743 (N_8743,N_4157,N_418);
xor U8744 (N_8744,N_4506,N_1535);
and U8745 (N_8745,N_4750,N_444);
nor U8746 (N_8746,N_795,N_2502);
or U8747 (N_8747,N_3244,N_5357);
nand U8748 (N_8748,N_58,N_1884);
xnor U8749 (N_8749,N_3144,N_3229);
and U8750 (N_8750,N_871,N_130);
nor U8751 (N_8751,N_3579,N_1474);
or U8752 (N_8752,N_4174,N_131);
xor U8753 (N_8753,N_1674,N_5867);
nor U8754 (N_8754,N_4983,N_5225);
xor U8755 (N_8755,N_275,N_5202);
nor U8756 (N_8756,N_3581,N_3793);
nor U8757 (N_8757,N_1650,N_5329);
xor U8758 (N_8758,N_2778,N_1753);
nand U8759 (N_8759,N_5510,N_1078);
and U8760 (N_8760,N_3845,N_4399);
nor U8761 (N_8761,N_509,N_1485);
nor U8762 (N_8762,N_2774,N_5335);
nand U8763 (N_8763,N_2559,N_3684);
or U8764 (N_8764,N_1577,N_1613);
xnor U8765 (N_8765,N_3509,N_2884);
nor U8766 (N_8766,N_499,N_2094);
nor U8767 (N_8767,N_1133,N_324);
nor U8768 (N_8768,N_4415,N_5922);
xor U8769 (N_8769,N_1327,N_5926);
nand U8770 (N_8770,N_4392,N_1291);
nor U8771 (N_8771,N_907,N_5288);
and U8772 (N_8772,N_4751,N_5199);
nor U8773 (N_8773,N_4376,N_2876);
nand U8774 (N_8774,N_3065,N_1325);
and U8775 (N_8775,N_1664,N_1176);
xnor U8776 (N_8776,N_3233,N_5273);
xnor U8777 (N_8777,N_1543,N_515);
or U8778 (N_8778,N_284,N_3777);
xor U8779 (N_8779,N_2844,N_5378);
nand U8780 (N_8780,N_481,N_3798);
xnor U8781 (N_8781,N_5903,N_1695);
nor U8782 (N_8782,N_3459,N_2631);
and U8783 (N_8783,N_1820,N_3508);
nor U8784 (N_8784,N_313,N_4389);
nand U8785 (N_8785,N_4741,N_1560);
or U8786 (N_8786,N_4160,N_276);
or U8787 (N_8787,N_1894,N_4548);
nand U8788 (N_8788,N_5697,N_5182);
nand U8789 (N_8789,N_3781,N_5468);
nand U8790 (N_8790,N_3198,N_3146);
nand U8791 (N_8791,N_114,N_4822);
nor U8792 (N_8792,N_5377,N_2761);
nand U8793 (N_8793,N_1718,N_2123);
or U8794 (N_8794,N_6237,N_5195);
or U8795 (N_8795,N_4519,N_3282);
nand U8796 (N_8796,N_1486,N_1824);
or U8797 (N_8797,N_2381,N_3832);
xnor U8798 (N_8798,N_4720,N_1838);
nand U8799 (N_8799,N_2129,N_2175);
xor U8800 (N_8800,N_2918,N_2346);
and U8801 (N_8801,N_4332,N_5905);
or U8802 (N_8802,N_1510,N_3072);
xnor U8803 (N_8803,N_2229,N_2985);
nand U8804 (N_8804,N_3099,N_5113);
or U8805 (N_8805,N_1690,N_3366);
and U8806 (N_8806,N_5326,N_4492);
nor U8807 (N_8807,N_2363,N_6217);
nor U8808 (N_8808,N_4521,N_2832);
and U8809 (N_8809,N_3167,N_601);
xnor U8810 (N_8810,N_4045,N_5494);
nand U8811 (N_8811,N_1553,N_823);
nor U8812 (N_8812,N_3142,N_696);
or U8813 (N_8813,N_5178,N_3036);
nor U8814 (N_8814,N_113,N_5430);
or U8815 (N_8815,N_6163,N_1855);
or U8816 (N_8816,N_3015,N_1928);
or U8817 (N_8817,N_3188,N_1993);
xor U8818 (N_8818,N_3700,N_471);
and U8819 (N_8819,N_987,N_2108);
nor U8820 (N_8820,N_1656,N_1215);
nor U8821 (N_8821,N_15,N_517);
or U8822 (N_8822,N_309,N_2359);
xor U8823 (N_8823,N_2801,N_6120);
or U8824 (N_8824,N_3213,N_5498);
and U8825 (N_8825,N_660,N_1178);
xor U8826 (N_8826,N_3127,N_5260);
xor U8827 (N_8827,N_4555,N_4023);
or U8828 (N_8828,N_5145,N_4613);
and U8829 (N_8829,N_2205,N_4927);
xor U8830 (N_8830,N_1294,N_2282);
nor U8831 (N_8831,N_458,N_770);
or U8832 (N_8832,N_1961,N_5201);
nand U8833 (N_8833,N_5861,N_478);
or U8834 (N_8834,N_1155,N_4250);
and U8835 (N_8835,N_853,N_9);
or U8836 (N_8836,N_4331,N_115);
nor U8837 (N_8837,N_2614,N_747);
xor U8838 (N_8838,N_941,N_1975);
nor U8839 (N_8839,N_2859,N_2440);
nand U8840 (N_8840,N_3068,N_778);
and U8841 (N_8841,N_1784,N_5891);
xor U8842 (N_8842,N_6174,N_5469);
xor U8843 (N_8843,N_2540,N_2302);
nand U8844 (N_8844,N_961,N_488);
xnor U8845 (N_8845,N_3209,N_4806);
or U8846 (N_8846,N_3601,N_4488);
xor U8847 (N_8847,N_3210,N_1921);
nand U8848 (N_8848,N_4840,N_3262);
xnor U8849 (N_8849,N_2249,N_5301);
and U8850 (N_8850,N_6203,N_4047);
and U8851 (N_8851,N_2417,N_888);
and U8852 (N_8852,N_3329,N_5923);
nand U8853 (N_8853,N_4000,N_638);
and U8854 (N_8854,N_1584,N_1432);
nor U8855 (N_8855,N_1978,N_5258);
xor U8856 (N_8856,N_4463,N_1428);
or U8857 (N_8857,N_4552,N_4102);
and U8858 (N_8858,N_3027,N_4707);
or U8859 (N_8859,N_864,N_1611);
and U8860 (N_8860,N_5673,N_5208);
or U8861 (N_8861,N_4842,N_357);
and U8862 (N_8862,N_2124,N_4652);
xor U8863 (N_8863,N_3017,N_6136);
or U8864 (N_8864,N_4234,N_2642);
nand U8865 (N_8865,N_6051,N_474);
nor U8866 (N_8866,N_854,N_5165);
and U8867 (N_8867,N_1036,N_5771);
or U8868 (N_8868,N_3283,N_2142);
nor U8869 (N_8869,N_5155,N_3640);
or U8870 (N_8870,N_371,N_2871);
nor U8871 (N_8871,N_1420,N_5661);
nand U8872 (N_8872,N_4119,N_5062);
nand U8873 (N_8873,N_5312,N_381);
nand U8874 (N_8874,N_6218,N_4010);
xor U8875 (N_8875,N_5153,N_1743);
xnor U8876 (N_8876,N_2284,N_4075);
or U8877 (N_8877,N_4733,N_4746);
xnor U8878 (N_8878,N_4049,N_5980);
xor U8879 (N_8879,N_4237,N_2126);
or U8880 (N_8880,N_1408,N_521);
nand U8881 (N_8881,N_3435,N_118);
nand U8882 (N_8882,N_4756,N_5651);
nor U8883 (N_8883,N_2323,N_123);
or U8884 (N_8884,N_3998,N_2463);
or U8885 (N_8885,N_6023,N_527);
and U8886 (N_8886,N_4991,N_2414);
nor U8887 (N_8887,N_4922,N_555);
nand U8888 (N_8888,N_4845,N_4722);
xnor U8889 (N_8889,N_1769,N_4279);
or U8890 (N_8890,N_3856,N_5280);
and U8891 (N_8891,N_2474,N_5485);
or U8892 (N_8892,N_2328,N_4343);
nor U8893 (N_8893,N_712,N_2454);
or U8894 (N_8894,N_332,N_3211);
or U8895 (N_8895,N_3403,N_443);
nand U8896 (N_8896,N_4639,N_1032);
nor U8897 (N_8897,N_4744,N_3394);
nor U8898 (N_8898,N_5295,N_6005);
xnor U8899 (N_8899,N_125,N_1041);
xnor U8900 (N_8900,N_1451,N_2511);
nor U8901 (N_8901,N_1138,N_1435);
or U8902 (N_8902,N_5886,N_6004);
xnor U8903 (N_8903,N_1169,N_4674);
xnor U8904 (N_8904,N_2295,N_4426);
nor U8905 (N_8905,N_432,N_1875);
nor U8906 (N_8906,N_3140,N_3252);
xor U8907 (N_8907,N_3353,N_3484);
xor U8908 (N_8908,N_5017,N_2403);
or U8909 (N_8909,N_5620,N_170);
and U8910 (N_8910,N_583,N_552);
or U8911 (N_8911,N_2358,N_3053);
nand U8912 (N_8912,N_4466,N_3268);
nand U8913 (N_8913,N_1429,N_3496);
nand U8914 (N_8914,N_4873,N_5680);
nand U8915 (N_8915,N_3195,N_4092);
and U8916 (N_8916,N_3817,N_3150);
nand U8917 (N_8917,N_2677,N_5411);
nand U8918 (N_8918,N_211,N_4762);
nor U8919 (N_8919,N_1224,N_2157);
xnor U8920 (N_8920,N_589,N_5005);
xnor U8921 (N_8921,N_3391,N_4770);
nor U8922 (N_8922,N_3217,N_2821);
nand U8923 (N_8923,N_4146,N_5506);
and U8924 (N_8924,N_5417,N_452);
or U8925 (N_8925,N_2453,N_5856);
nand U8926 (N_8926,N_3913,N_5318);
nor U8927 (N_8927,N_3330,N_1648);
xor U8928 (N_8928,N_3156,N_226);
and U8929 (N_8929,N_1737,N_4850);
nor U8930 (N_8930,N_5985,N_5238);
nor U8931 (N_8931,N_3125,N_358);
and U8932 (N_8932,N_5227,N_4977);
or U8933 (N_8933,N_5996,N_1954);
or U8934 (N_8934,N_1711,N_3442);
xnor U8935 (N_8935,N_1150,N_5995);
nand U8936 (N_8936,N_2872,N_5563);
nand U8937 (N_8937,N_531,N_4681);
or U8938 (N_8938,N_5687,N_6193);
nand U8939 (N_8939,N_5791,N_6176);
or U8940 (N_8940,N_682,N_1035);
or U8941 (N_8941,N_2256,N_801);
and U8942 (N_8942,N_1844,N_2547);
nand U8943 (N_8943,N_6083,N_706);
and U8944 (N_8944,N_4486,N_2762);
and U8945 (N_8945,N_426,N_901);
and U8946 (N_8946,N_3437,N_4276);
and U8947 (N_8947,N_4210,N_1477);
and U8948 (N_8948,N_3834,N_375);
nor U8949 (N_8949,N_4104,N_473);
nor U8950 (N_8950,N_89,N_5536);
or U8951 (N_8951,N_1089,N_80);
or U8952 (N_8952,N_4216,N_3665);
or U8953 (N_8953,N_3473,N_66);
and U8954 (N_8954,N_1443,N_4454);
nand U8955 (N_8955,N_3825,N_3153);
or U8956 (N_8956,N_1160,N_2449);
xor U8957 (N_8957,N_2707,N_4158);
nor U8958 (N_8958,N_4885,N_2243);
nand U8959 (N_8959,N_5531,N_3260);
and U8960 (N_8960,N_3641,N_1783);
and U8961 (N_8961,N_3136,N_2577);
and U8962 (N_8962,N_2267,N_73);
and U8963 (N_8963,N_814,N_5035);
or U8964 (N_8964,N_1594,N_5122);
xor U8965 (N_8965,N_81,N_4337);
and U8966 (N_8966,N_5999,N_1669);
nand U8967 (N_8967,N_4340,N_892);
or U8968 (N_8968,N_1512,N_3685);
xor U8969 (N_8969,N_60,N_3044);
or U8970 (N_8970,N_2904,N_976);
nor U8971 (N_8971,N_5618,N_5068);
nand U8972 (N_8972,N_85,N_6068);
or U8973 (N_8973,N_4661,N_536);
or U8974 (N_8974,N_3891,N_2519);
and U8975 (N_8975,N_1998,N_162);
or U8976 (N_8976,N_2172,N_2244);
and U8977 (N_8977,N_4601,N_1536);
or U8978 (N_8978,N_5065,N_1055);
nand U8979 (N_8979,N_1600,N_5997);
nand U8980 (N_8980,N_1937,N_2885);
xnor U8981 (N_8981,N_3324,N_1103);
nand U8982 (N_8982,N_3814,N_4142);
and U8983 (N_8983,N_5639,N_63);
and U8984 (N_8984,N_1275,N_1439);
or U8985 (N_8985,N_2497,N_1804);
or U8986 (N_8986,N_1,N_3432);
nand U8987 (N_8987,N_3970,N_5034);
nor U8988 (N_8988,N_3598,N_4346);
nand U8989 (N_8989,N_4568,N_3454);
nor U8990 (N_8990,N_734,N_6205);
nand U8991 (N_8991,N_1365,N_3862);
nand U8992 (N_8992,N_5463,N_413);
and U8993 (N_8993,N_5760,N_5511);
xor U8994 (N_8994,N_6063,N_3716);
nor U8995 (N_8995,N_6041,N_4847);
and U8996 (N_8996,N_2472,N_4307);
nor U8997 (N_8997,N_3708,N_47);
xnor U8998 (N_8998,N_316,N_584);
nand U8999 (N_8999,N_3491,N_5120);
xor U9000 (N_9000,N_1819,N_2487);
xor U9001 (N_9001,N_3826,N_4318);
or U9002 (N_9002,N_64,N_2113);
or U9003 (N_9003,N_514,N_2813);
xor U9004 (N_9004,N_2678,N_2034);
and U9005 (N_9005,N_3242,N_3492);
xnor U9006 (N_9006,N_3657,N_93);
or U9007 (N_9007,N_4727,N_5813);
nor U9008 (N_9008,N_1442,N_3548);
nand U9009 (N_9009,N_4764,N_6158);
and U9010 (N_9010,N_5109,N_5507);
nor U9011 (N_9011,N_4724,N_3673);
and U9012 (N_9012,N_1766,N_5496);
nor U9013 (N_9013,N_5870,N_3259);
nor U9014 (N_9014,N_1731,N_4910);
nor U9015 (N_9015,N_3620,N_5733);
xnor U9016 (N_9016,N_3230,N_3204);
or U9017 (N_9017,N_4444,N_1531);
nand U9018 (N_9018,N_5762,N_4686);
nand U9019 (N_9019,N_2188,N_574);
nand U9020 (N_9020,N_5437,N_642);
and U9021 (N_9021,N_56,N_1257);
xnor U9022 (N_9022,N_4299,N_1538);
or U9023 (N_9023,N_689,N_3370);
nand U9024 (N_9024,N_5528,N_2905);
nand U9025 (N_9025,N_2946,N_4159);
nor U9026 (N_9026,N_2128,N_5649);
nor U9027 (N_9027,N_3677,N_5272);
and U9028 (N_9028,N_3989,N_2020);
nand U9029 (N_9029,N_794,N_5654);
or U9030 (N_9030,N_4496,N_2622);
nor U9031 (N_9031,N_4743,N_2669);
nand U9032 (N_9032,N_6067,N_5513);
nand U9033 (N_9033,N_3418,N_3154);
or U9034 (N_9034,N_787,N_5453);
nor U9035 (N_9035,N_3322,N_538);
and U9036 (N_9036,N_1582,N_3075);
and U9037 (N_9037,N_2084,N_3982);
or U9038 (N_9038,N_5567,N_825);
xor U9039 (N_9039,N_5819,N_4540);
and U9040 (N_9040,N_3788,N_3004);
nand U9041 (N_9041,N_3248,N_4144);
and U9042 (N_9042,N_930,N_1471);
xnor U9043 (N_9043,N_1267,N_955);
nor U9044 (N_9044,N_4955,N_1247);
nand U9045 (N_9045,N_5777,N_6186);
nand U9046 (N_9046,N_5395,N_5526);
nor U9047 (N_9047,N_3765,N_4619);
or U9048 (N_9048,N_1570,N_336);
xor U9049 (N_9049,N_4836,N_2637);
nor U9050 (N_9050,N_6093,N_2658);
or U9051 (N_9051,N_1913,N_3137);
nor U9052 (N_9052,N_6121,N_4563);
nand U9053 (N_9053,N_3811,N_2354);
and U9054 (N_9054,N_863,N_4099);
and U9055 (N_9055,N_362,N_448);
xor U9056 (N_9056,N_3795,N_491);
nor U9057 (N_9057,N_1513,N_3175);
or U9058 (N_9058,N_2389,N_396);
or U9059 (N_9059,N_469,N_3287);
nor U9060 (N_9060,N_948,N_1379);
nor U9061 (N_9061,N_461,N_1367);
xor U9062 (N_9062,N_40,N_1867);
nor U9063 (N_9063,N_5684,N_3683);
and U9064 (N_9064,N_3343,N_4950);
and U9065 (N_9065,N_4095,N_1105);
xor U9066 (N_9066,N_4992,N_2747);
nand U9067 (N_9067,N_5163,N_1569);
nor U9068 (N_9068,N_5041,N_2932);
nor U9069 (N_9069,N_6129,N_522);
nor U9070 (N_9070,N_715,N_2931);
nor U9071 (N_9071,N_4685,N_2814);
or U9072 (N_9072,N_3236,N_3686);
nand U9073 (N_9073,N_6059,N_364);
nand U9074 (N_9074,N_1984,N_3861);
nor U9075 (N_9075,N_2356,N_5663);
and U9076 (N_9076,N_4123,N_4951);
nor U9077 (N_9077,N_3485,N_3648);
nand U9078 (N_9078,N_2050,N_3030);
nand U9079 (N_9079,N_3758,N_2668);
nand U9080 (N_9080,N_322,N_3111);
or U9081 (N_9081,N_6175,N_5554);
nor U9082 (N_9082,N_3971,N_2705);
nand U9083 (N_9083,N_669,N_495);
or U9084 (N_9084,N_257,N_4185);
nand U9085 (N_9085,N_194,N_5675);
and U9086 (N_9086,N_5279,N_5717);
and U9087 (N_9087,N_5808,N_5839);
nor U9088 (N_9088,N_1991,N_4022);
or U9089 (N_9089,N_2402,N_4892);
or U9090 (N_9090,N_3918,N_4193);
nand U9091 (N_9091,N_4125,N_3570);
nand U9092 (N_9092,N_3679,N_5091);
or U9093 (N_9093,N_399,N_687);
xnor U9094 (N_9094,N_1777,N_5583);
or U9095 (N_9095,N_5446,N_2325);
xnor U9096 (N_9096,N_2831,N_688);
nand U9097 (N_9097,N_5736,N_699);
nand U9098 (N_9098,N_3820,N_3361);
nor U9099 (N_9099,N_1704,N_4708);
nand U9100 (N_9100,N_4557,N_5336);
xnor U9101 (N_9101,N_1590,N_5775);
xor U9102 (N_9102,N_2138,N_2947);
xnor U9103 (N_9103,N_6199,N_326);
xor U9104 (N_9104,N_2336,N_498);
nand U9105 (N_9105,N_2900,N_5240);
nor U9106 (N_9106,N_1761,N_4231);
xor U9107 (N_9107,N_4615,N_559);
or U9108 (N_9108,N_5648,N_2018);
and U9109 (N_9109,N_5920,N_5244);
nand U9110 (N_9110,N_4089,N_4461);
or U9111 (N_9111,N_4292,N_5169);
nor U9112 (N_9112,N_1541,N_3966);
nor U9113 (N_9113,N_2278,N_3290);
xnor U9114 (N_9114,N_1957,N_1889);
or U9115 (N_9115,N_4752,N_5266);
and U9116 (N_9116,N_224,N_3169);
and U9117 (N_9117,N_954,N_4012);
xor U9118 (N_9118,N_373,N_5956);
xnor U9119 (N_9119,N_6246,N_6102);
nor U9120 (N_9120,N_1762,N_849);
nor U9121 (N_9121,N_1673,N_5662);
or U9122 (N_9122,N_5172,N_4252);
or U9123 (N_9123,N_4248,N_3877);
xnor U9124 (N_9124,N_859,N_1658);
nor U9125 (N_9125,N_2720,N_5257);
or U9126 (N_9126,N_3448,N_4302);
xnor U9127 (N_9127,N_3311,N_3016);
nand U9128 (N_9128,N_3997,N_2735);
nand U9129 (N_9129,N_6249,N_2065);
xor U9130 (N_9130,N_3668,N_4401);
nor U9131 (N_9131,N_5994,N_1151);
nand U9132 (N_9132,N_3839,N_905);
and U9133 (N_9133,N_2042,N_3835);
and U9134 (N_9134,N_3152,N_622);
xnor U9135 (N_9135,N_4003,N_5774);
nand U9136 (N_9136,N_5726,N_2406);
and U9137 (N_9137,N_2530,N_5529);
and U9138 (N_9138,N_5261,N_2673);
nor U9139 (N_9139,N_4523,N_5548);
xnor U9140 (N_9140,N_2085,N_3221);
or U9141 (N_9141,N_1780,N_2889);
nand U9142 (N_9142,N_4677,N_2746);
nand U9143 (N_9143,N_4972,N_2899);
nor U9144 (N_9144,N_4926,N_5206);
xor U9145 (N_9145,N_5574,N_3119);
xnor U9146 (N_9146,N_599,N_5952);
and U9147 (N_9147,N_728,N_940);
xnor U9148 (N_9148,N_2443,N_1808);
and U9149 (N_9149,N_999,N_3526);
nor U9150 (N_9150,N_2149,N_5140);
and U9151 (N_9151,N_1706,N_1725);
and U9152 (N_9152,N_2823,N_1542);
xor U9153 (N_9153,N_5689,N_2983);
nand U9154 (N_9154,N_6069,N_168);
xnor U9155 (N_9155,N_3267,N_2062);
or U9156 (N_9156,N_1389,N_1610);
nor U9157 (N_9157,N_2827,N_579);
or U9158 (N_9158,N_3589,N_668);
xor U9159 (N_9159,N_4841,N_3516);
and U9160 (N_9160,N_3945,N_5877);
nor U9161 (N_9161,N_1566,N_3794);
nor U9162 (N_9162,N_2627,N_2672);
or U9163 (N_9163,N_5705,N_887);
xnor U9164 (N_9164,N_5289,N_5409);
nor U9165 (N_9165,N_3054,N_2799);
xnor U9166 (N_9166,N_1069,N_3220);
and U9167 (N_9167,N_3467,N_3553);
or U9168 (N_9168,N_5859,N_193);
nand U9169 (N_9169,N_4976,N_2697);
nand U9170 (N_9170,N_1657,N_3830);
nand U9171 (N_9171,N_5576,N_2178);
and U9172 (N_9172,N_769,N_1243);
and U9173 (N_9173,N_4721,N_4669);
xor U9174 (N_9174,N_2340,N_4393);
nor U9175 (N_9175,N_5308,N_5619);
nand U9176 (N_9176,N_2063,N_5489);
xnor U9177 (N_9177,N_3284,N_2039);
nor U9178 (N_9178,N_6009,N_420);
and U9179 (N_9179,N_4589,N_1172);
and U9180 (N_9180,N_4614,N_2940);
or U9181 (N_9181,N_2676,N_1771);
or U9182 (N_9182,N_1979,N_5168);
xor U9183 (N_9183,N_2041,N_129);
or U9184 (N_9184,N_1481,N_3478);
nand U9185 (N_9185,N_1458,N_4495);
nor U9186 (N_9186,N_1550,N_2716);
xnor U9187 (N_9187,N_6039,N_3815);
nand U9188 (N_9188,N_2322,N_4570);
xor U9189 (N_9189,N_2468,N_4627);
and U9190 (N_9190,N_4386,N_2733);
nand U9191 (N_9191,N_2566,N_5119);
nand U9192 (N_9192,N_4199,N_501);
xnor U9193 (N_9193,N_2881,N_4586);
or U9194 (N_9194,N_2027,N_282);
xnor U9195 (N_9195,N_1911,N_2957);
xnor U9196 (N_9196,N_4380,N_4848);
nand U9197 (N_9197,N_294,N_4971);
xor U9198 (N_9198,N_679,N_2333);
and U9199 (N_9199,N_5552,N_4287);
and U9200 (N_9200,N_3312,N_2850);
and U9201 (N_9201,N_4429,N_4867);
nor U9202 (N_9202,N_1273,N_4437);
and U9203 (N_9203,N_1387,N_5313);
nand U9204 (N_9204,N_5495,N_1096);
nand U9205 (N_9205,N_16,N_82);
or U9206 (N_9206,N_5270,N_2460);
xor U9207 (N_9207,N_3596,N_1750);
xor U9208 (N_9208,N_4015,N_578);
xnor U9209 (N_9209,N_1026,N_2600);
nand U9210 (N_9210,N_1354,N_685);
xor U9211 (N_9211,N_1843,N_1125);
and U9212 (N_9212,N_3907,N_3176);
and U9213 (N_9213,N_4040,N_3272);
nor U9214 (N_9214,N_5932,N_6144);
or U9215 (N_9215,N_5384,N_3763);
or U9216 (N_9216,N_2583,N_6231);
xor U9217 (N_9217,N_1444,N_629);
nor U9218 (N_9218,N_2002,N_6007);
nand U9219 (N_9219,N_1304,N_4590);
nor U9220 (N_9220,N_1009,N_6133);
xor U9221 (N_9221,N_3687,N_4284);
nand U9222 (N_9222,N_4171,N_37);
or U9223 (N_9223,N_1173,N_5807);
or U9224 (N_9224,N_1888,N_3314);
xor U9225 (N_9225,N_2605,N_4993);
and U9226 (N_9226,N_285,N_5592);
nand U9227 (N_9227,N_2332,N_3506);
and U9228 (N_9228,N_3253,N_3245);
nor U9229 (N_9229,N_2404,N_3995);
or U9230 (N_9230,N_2292,N_3764);
xor U9231 (N_9231,N_6053,N_4363);
xor U9232 (N_9232,N_2180,N_655);
xor U9233 (N_9233,N_5604,N_3504);
or U9234 (N_9234,N_3842,N_3747);
nor U9235 (N_9235,N_2135,N_1410);
xnor U9236 (N_9236,N_5354,N_6215);
nand U9237 (N_9237,N_5692,N_2662);
or U9238 (N_9238,N_5173,N_1437);
and U9239 (N_9239,N_3218,N_1006);
and U9240 (N_9240,N_243,N_5056);
xor U9241 (N_9241,N_805,N_1973);
nor U9242 (N_9242,N_6162,N_1945);
xnor U9243 (N_9243,N_2887,N_3327);
or U9244 (N_9244,N_4149,N_719);
xor U9245 (N_9245,N_5873,N_4868);
and U9246 (N_9246,N_5551,N_1728);
and U9247 (N_9247,N_2741,N_3580);
and U9248 (N_9248,N_4936,N_1723);
nand U9249 (N_9249,N_2131,N_5878);
nand U9250 (N_9250,N_2638,N_502);
xor U9251 (N_9251,N_1965,N_1832);
xor U9252 (N_9252,N_5874,N_164);
nor U9253 (N_9253,N_2536,N_3059);
and U9254 (N_9254,N_3587,N_5728);
xnor U9255 (N_9255,N_970,N_1380);
xnor U9256 (N_9256,N_1003,N_2602);
or U9257 (N_9257,N_647,N_1434);
and U9258 (N_9258,N_1119,N_1930);
xnor U9259 (N_9259,N_3390,N_3701);
nand U9260 (N_9260,N_1496,N_490);
nand U9261 (N_9261,N_5464,N_1791);
xor U9262 (N_9262,N_4611,N_838);
and U9263 (N_9263,N_3819,N_447);
xnor U9264 (N_9264,N_5,N_3733);
xor U9265 (N_9265,N_4797,N_4931);
and U9266 (N_9266,N_4695,N_562);
and U9267 (N_9267,N_4134,N_1299);
nand U9268 (N_9268,N_5763,N_4269);
nand U9269 (N_9269,N_4175,N_3718);
nand U9270 (N_9270,N_5136,N_5953);
nor U9271 (N_9271,N_62,N_4699);
nand U9272 (N_9272,N_5888,N_4562);
nor U9273 (N_9273,N_1438,N_5428);
nand U9274 (N_9274,N_5491,N_3336);
nand U9275 (N_9275,N_5399,N_4754);
and U9276 (N_9276,N_4651,N_2706);
or U9277 (N_9277,N_2019,N_5360);
and U9278 (N_9278,N_2793,N_3047);
nand U9279 (N_9279,N_4270,N_737);
nand U9280 (N_9280,N_5543,N_2331);
xor U9281 (N_9281,N_1540,N_5365);
nand U9282 (N_9282,N_1289,N_5407);
nor U9283 (N_9283,N_2007,N_4472);
and U9284 (N_9284,N_4,N_2984);
and U9285 (N_9285,N_5083,N_4819);
or U9286 (N_9286,N_4008,N_4816);
nand U9287 (N_9287,N_2901,N_3863);
or U9288 (N_9288,N_2426,N_4088);
nand U9289 (N_9289,N_4005,N_3346);
xnor U9290 (N_9290,N_5502,N_1166);
nand U9291 (N_9291,N_4388,N_3488);
and U9292 (N_9292,N_2377,N_104);
or U9293 (N_9293,N_5419,N_2127);
and U9294 (N_9294,N_3515,N_1140);
xnor U9295 (N_9295,N_2119,N_5993);
xnor U9296 (N_9296,N_2169,N_454);
xor U9297 (N_9297,N_890,N_5066);
nand U9298 (N_9298,N_350,N_1413);
and U9299 (N_9299,N_1220,N_2051);
nor U9300 (N_9300,N_4404,N_1219);
nand U9301 (N_9301,N_4336,N_4070);
nand U9302 (N_9302,N_4192,N_3857);
or U9303 (N_9303,N_3061,N_303);
nand U9304 (N_9304,N_4988,N_5627);
and U9305 (N_9305,N_3615,N_5892);
nand U9306 (N_9306,N_4513,N_1837);
nand U9307 (N_9307,N_2191,N_304);
or U9308 (N_9308,N_3896,N_126);
nor U9309 (N_9309,N_1080,N_462);
nand U9310 (N_9310,N_3690,N_2217);
xnor U9311 (N_9311,N_2348,N_6139);
and U9312 (N_9312,N_3841,N_4247);
nand U9313 (N_9313,N_553,N_5476);
nand U9314 (N_9314,N_1077,N_245);
xor U9315 (N_9315,N_150,N_152);
nor U9316 (N_9316,N_4974,N_2037);
and U9317 (N_9317,N_2656,N_268);
nor U9318 (N_9318,N_998,N_3871);
or U9319 (N_9319,N_3604,N_4271);
or U9320 (N_9320,N_4151,N_5709);
or U9321 (N_9321,N_1418,N_4260);
or U9322 (N_9322,N_4667,N_576);
and U9323 (N_9323,N_4990,N_5519);
nor U9324 (N_9324,N_6054,N_2419);
xor U9325 (N_9325,N_4081,N_2010);
nor U9326 (N_9326,N_2200,N_771);
or U9327 (N_9327,N_5986,N_101);
or U9328 (N_9328,N_1028,N_2570);
xnor U9329 (N_9329,N_5978,N_78);
and U9330 (N_9330,N_228,N_4329);
nor U9331 (N_9331,N_5515,N_4118);
or U9332 (N_9332,N_1093,N_2448);
and U9333 (N_9333,N_1775,N_4626);
xor U9334 (N_9334,N_4759,N_4571);
and U9335 (N_9335,N_5896,N_3197);
nor U9336 (N_9336,N_710,N_3223);
nand U9337 (N_9337,N_6145,N_733);
or U9338 (N_9338,N_2194,N_564);
nand U9339 (N_9339,N_3200,N_320);
and U9340 (N_9340,N_1011,N_2711);
nand U9341 (N_9341,N_2090,N_1110);
nor U9342 (N_9342,N_5455,N_546);
nor U9343 (N_9343,N_5064,N_5405);
and U9344 (N_9344,N_1290,N_828);
xnor U9345 (N_9345,N_5393,N_4596);
nor U9346 (N_9346,N_1579,N_1549);
nor U9347 (N_9347,N_1144,N_1999);
nor U9348 (N_9348,N_1255,N_4315);
xnor U9349 (N_9349,N_5699,N_2592);
or U9350 (N_9350,N_3710,N_937);
nand U9351 (N_9351,N_1308,N_5933);
nand U9352 (N_9352,N_5449,N_1487);
or U9353 (N_9353,N_2100,N_1986);
nand U9354 (N_9354,N_6153,N_5647);
or U9355 (N_9355,N_1311,N_5785);
nand U9356 (N_9356,N_1057,N_2848);
nor U9357 (N_9357,N_4366,N_1101);
and U9358 (N_9358,N_4920,N_1293);
and U9359 (N_9359,N_731,N_4760);
nand U9360 (N_9360,N_5071,N_3293);
and U9361 (N_9361,N_5251,N_544);
xnor U9362 (N_9362,N_3932,N_86);
and U9363 (N_9363,N_4338,N_758);
nand U9364 (N_9364,N_580,N_31);
nand U9365 (N_9365,N_3316,N_504);
or U9366 (N_9366,N_4534,N_5729);
nor U9367 (N_9367,N_750,N_3638);
and U9368 (N_9368,N_3453,N_4058);
nor U9369 (N_9369,N_4073,N_5296);
nor U9370 (N_9370,N_65,N_2091);
and U9371 (N_9371,N_2663,N_1726);
and U9372 (N_9372,N_3381,N_826);
and U9373 (N_9373,N_165,N_5927);
nand U9374 (N_9374,N_1744,N_6032);
xnor U9375 (N_9375,N_1858,N_2087);
nand U9376 (N_9376,N_6093,N_4779);
and U9377 (N_9377,N_5076,N_3174);
or U9378 (N_9378,N_3298,N_6131);
and U9379 (N_9379,N_4711,N_6174);
and U9380 (N_9380,N_2961,N_334);
nor U9381 (N_9381,N_4748,N_282);
or U9382 (N_9382,N_4106,N_2444);
or U9383 (N_9383,N_2944,N_5868);
nor U9384 (N_9384,N_4765,N_286);
and U9385 (N_9385,N_1949,N_5346);
or U9386 (N_9386,N_4706,N_5586);
xor U9387 (N_9387,N_1636,N_207);
or U9388 (N_9388,N_3638,N_1587);
nand U9389 (N_9389,N_749,N_4852);
nand U9390 (N_9390,N_5573,N_4636);
xor U9391 (N_9391,N_4332,N_5475);
nor U9392 (N_9392,N_814,N_3552);
or U9393 (N_9393,N_3038,N_3792);
xor U9394 (N_9394,N_2960,N_200);
and U9395 (N_9395,N_2529,N_6224);
nand U9396 (N_9396,N_436,N_5863);
xnor U9397 (N_9397,N_2262,N_5522);
nor U9398 (N_9398,N_320,N_3113);
or U9399 (N_9399,N_4704,N_5572);
nand U9400 (N_9400,N_4061,N_5847);
nor U9401 (N_9401,N_3773,N_706);
or U9402 (N_9402,N_1025,N_1451);
and U9403 (N_9403,N_1401,N_4095);
nor U9404 (N_9404,N_414,N_2772);
or U9405 (N_9405,N_4067,N_4174);
or U9406 (N_9406,N_796,N_704);
nand U9407 (N_9407,N_3777,N_4556);
and U9408 (N_9408,N_4118,N_4578);
nor U9409 (N_9409,N_2859,N_3348);
nor U9410 (N_9410,N_179,N_2861);
or U9411 (N_9411,N_4227,N_5738);
or U9412 (N_9412,N_1546,N_2063);
or U9413 (N_9413,N_1425,N_2388);
and U9414 (N_9414,N_1967,N_1493);
and U9415 (N_9415,N_5834,N_4805);
and U9416 (N_9416,N_5178,N_3418);
nand U9417 (N_9417,N_929,N_83);
nand U9418 (N_9418,N_721,N_1888);
nand U9419 (N_9419,N_5303,N_5965);
xnor U9420 (N_9420,N_35,N_5965);
xnor U9421 (N_9421,N_1471,N_795);
nand U9422 (N_9422,N_4711,N_3579);
xnor U9423 (N_9423,N_3910,N_5499);
or U9424 (N_9424,N_2991,N_93);
nor U9425 (N_9425,N_3608,N_517);
and U9426 (N_9426,N_2345,N_2933);
nor U9427 (N_9427,N_4536,N_4928);
nand U9428 (N_9428,N_4402,N_4659);
nor U9429 (N_9429,N_3428,N_4773);
nor U9430 (N_9430,N_1786,N_3784);
nand U9431 (N_9431,N_5639,N_2840);
nor U9432 (N_9432,N_322,N_4137);
nand U9433 (N_9433,N_1710,N_1224);
nand U9434 (N_9434,N_2586,N_2730);
nand U9435 (N_9435,N_2436,N_248);
nor U9436 (N_9436,N_2404,N_2002);
and U9437 (N_9437,N_517,N_2371);
or U9438 (N_9438,N_3285,N_2897);
or U9439 (N_9439,N_664,N_559);
xnor U9440 (N_9440,N_4658,N_3740);
nand U9441 (N_9441,N_4794,N_3539);
nor U9442 (N_9442,N_1062,N_482);
nand U9443 (N_9443,N_5975,N_2076);
and U9444 (N_9444,N_3966,N_2693);
or U9445 (N_9445,N_2547,N_546);
or U9446 (N_9446,N_1725,N_4940);
xor U9447 (N_9447,N_5995,N_1374);
nand U9448 (N_9448,N_2798,N_6091);
xor U9449 (N_9449,N_145,N_5527);
and U9450 (N_9450,N_517,N_4854);
xor U9451 (N_9451,N_4011,N_615);
nor U9452 (N_9452,N_5751,N_2394);
or U9453 (N_9453,N_5688,N_2611);
nand U9454 (N_9454,N_1566,N_2768);
nand U9455 (N_9455,N_4993,N_5447);
or U9456 (N_9456,N_3599,N_27);
nor U9457 (N_9457,N_1861,N_1095);
xor U9458 (N_9458,N_2634,N_2368);
and U9459 (N_9459,N_5667,N_1439);
xnor U9460 (N_9460,N_2210,N_1851);
xnor U9461 (N_9461,N_5551,N_985);
nand U9462 (N_9462,N_4319,N_4375);
xnor U9463 (N_9463,N_4886,N_5691);
nand U9464 (N_9464,N_2748,N_460);
nand U9465 (N_9465,N_5944,N_4479);
nor U9466 (N_9466,N_824,N_3998);
and U9467 (N_9467,N_2610,N_4557);
or U9468 (N_9468,N_5909,N_1021);
or U9469 (N_9469,N_3957,N_1947);
or U9470 (N_9470,N_4480,N_2734);
and U9471 (N_9471,N_5204,N_2126);
or U9472 (N_9472,N_209,N_1936);
xnor U9473 (N_9473,N_3102,N_4491);
xnor U9474 (N_9474,N_1030,N_456);
nor U9475 (N_9475,N_3249,N_3856);
or U9476 (N_9476,N_3108,N_4772);
xnor U9477 (N_9477,N_755,N_3911);
or U9478 (N_9478,N_3064,N_2230);
xnor U9479 (N_9479,N_5283,N_5697);
nand U9480 (N_9480,N_2082,N_5880);
xor U9481 (N_9481,N_27,N_3627);
xor U9482 (N_9482,N_1820,N_3452);
and U9483 (N_9483,N_3989,N_1932);
xnor U9484 (N_9484,N_3268,N_4493);
nand U9485 (N_9485,N_5913,N_5353);
or U9486 (N_9486,N_6125,N_4541);
or U9487 (N_9487,N_2226,N_4666);
nand U9488 (N_9488,N_4549,N_2949);
xnor U9489 (N_9489,N_3671,N_1699);
or U9490 (N_9490,N_2549,N_5461);
nor U9491 (N_9491,N_3211,N_2560);
nand U9492 (N_9492,N_3588,N_828);
nand U9493 (N_9493,N_1826,N_4568);
and U9494 (N_9494,N_1163,N_1126);
nand U9495 (N_9495,N_1110,N_3091);
nor U9496 (N_9496,N_4466,N_1263);
nand U9497 (N_9497,N_1209,N_1823);
or U9498 (N_9498,N_5965,N_1120);
xor U9499 (N_9499,N_3550,N_345);
and U9500 (N_9500,N_5344,N_6186);
nor U9501 (N_9501,N_4725,N_5581);
nand U9502 (N_9502,N_4098,N_1966);
and U9503 (N_9503,N_3981,N_929);
nor U9504 (N_9504,N_5009,N_3060);
nand U9505 (N_9505,N_2764,N_190);
or U9506 (N_9506,N_841,N_4478);
xnor U9507 (N_9507,N_2438,N_2879);
xor U9508 (N_9508,N_970,N_809);
or U9509 (N_9509,N_3465,N_3421);
xnor U9510 (N_9510,N_1053,N_6097);
nand U9511 (N_9511,N_2830,N_267);
nor U9512 (N_9512,N_446,N_3256);
nand U9513 (N_9513,N_4499,N_1178);
or U9514 (N_9514,N_2315,N_2151);
nor U9515 (N_9515,N_4287,N_6048);
xor U9516 (N_9516,N_3352,N_1447);
nand U9517 (N_9517,N_5905,N_4923);
and U9518 (N_9518,N_4054,N_912);
xor U9519 (N_9519,N_4976,N_2036);
nand U9520 (N_9520,N_3778,N_3262);
xor U9521 (N_9521,N_2853,N_3308);
or U9522 (N_9522,N_2065,N_5112);
nor U9523 (N_9523,N_5338,N_5741);
xor U9524 (N_9524,N_5323,N_4791);
nor U9525 (N_9525,N_3686,N_1021);
or U9526 (N_9526,N_176,N_3280);
or U9527 (N_9527,N_5171,N_2430);
nor U9528 (N_9528,N_3853,N_2935);
nand U9529 (N_9529,N_3317,N_1457);
xor U9530 (N_9530,N_3173,N_3502);
nor U9531 (N_9531,N_1085,N_4997);
or U9532 (N_9532,N_3134,N_6219);
xor U9533 (N_9533,N_2123,N_786);
or U9534 (N_9534,N_237,N_4832);
nand U9535 (N_9535,N_1836,N_6203);
xnor U9536 (N_9536,N_4002,N_4839);
or U9537 (N_9537,N_263,N_5269);
and U9538 (N_9538,N_3695,N_1975);
and U9539 (N_9539,N_5877,N_2767);
nand U9540 (N_9540,N_1317,N_2181);
xnor U9541 (N_9541,N_2120,N_759);
nand U9542 (N_9542,N_5307,N_6061);
and U9543 (N_9543,N_1179,N_5040);
nor U9544 (N_9544,N_5756,N_1748);
nand U9545 (N_9545,N_2507,N_4654);
nand U9546 (N_9546,N_2886,N_2537);
nor U9547 (N_9547,N_4489,N_1448);
nor U9548 (N_9548,N_3294,N_2383);
xor U9549 (N_9549,N_2705,N_5462);
nand U9550 (N_9550,N_3270,N_5298);
and U9551 (N_9551,N_4880,N_3271);
and U9552 (N_9552,N_5613,N_4737);
nand U9553 (N_9553,N_820,N_375);
or U9554 (N_9554,N_3609,N_4293);
and U9555 (N_9555,N_4364,N_3203);
and U9556 (N_9556,N_167,N_5967);
or U9557 (N_9557,N_1721,N_873);
or U9558 (N_9558,N_5144,N_4529);
and U9559 (N_9559,N_3750,N_405);
nor U9560 (N_9560,N_473,N_1103);
or U9561 (N_9561,N_2549,N_3453);
xor U9562 (N_9562,N_5532,N_3292);
and U9563 (N_9563,N_4909,N_2623);
nand U9564 (N_9564,N_3894,N_3379);
nand U9565 (N_9565,N_2109,N_5181);
xnor U9566 (N_9566,N_4622,N_5212);
nand U9567 (N_9567,N_5468,N_5821);
and U9568 (N_9568,N_3529,N_4463);
or U9569 (N_9569,N_2493,N_5074);
nor U9570 (N_9570,N_4195,N_4861);
and U9571 (N_9571,N_511,N_30);
nor U9572 (N_9572,N_3365,N_2520);
and U9573 (N_9573,N_1054,N_5941);
xnor U9574 (N_9574,N_2494,N_5953);
xnor U9575 (N_9575,N_1020,N_4750);
nor U9576 (N_9576,N_4178,N_1672);
nor U9577 (N_9577,N_5645,N_392);
nor U9578 (N_9578,N_4033,N_2332);
and U9579 (N_9579,N_795,N_2212);
nor U9580 (N_9580,N_3643,N_2872);
or U9581 (N_9581,N_2758,N_5301);
xnor U9582 (N_9582,N_5011,N_5349);
xor U9583 (N_9583,N_621,N_2853);
nor U9584 (N_9584,N_35,N_5897);
or U9585 (N_9585,N_1270,N_1021);
or U9586 (N_9586,N_5737,N_5258);
nor U9587 (N_9587,N_5433,N_945);
xnor U9588 (N_9588,N_3026,N_5901);
or U9589 (N_9589,N_4529,N_1363);
and U9590 (N_9590,N_810,N_3344);
nor U9591 (N_9591,N_3626,N_535);
or U9592 (N_9592,N_5528,N_618);
nand U9593 (N_9593,N_2103,N_1191);
or U9594 (N_9594,N_2056,N_484);
nand U9595 (N_9595,N_5199,N_5261);
or U9596 (N_9596,N_3261,N_2815);
and U9597 (N_9597,N_2212,N_5473);
nor U9598 (N_9598,N_1763,N_4778);
or U9599 (N_9599,N_5971,N_5248);
or U9600 (N_9600,N_4765,N_796);
nor U9601 (N_9601,N_2387,N_5165);
xnor U9602 (N_9602,N_4936,N_1241);
nor U9603 (N_9603,N_4400,N_3687);
nand U9604 (N_9604,N_5240,N_105);
nand U9605 (N_9605,N_2507,N_3864);
and U9606 (N_9606,N_2022,N_3654);
and U9607 (N_9607,N_2114,N_4727);
and U9608 (N_9608,N_5791,N_1796);
and U9609 (N_9609,N_5669,N_5154);
nand U9610 (N_9610,N_2745,N_1678);
nor U9611 (N_9611,N_5549,N_1715);
xor U9612 (N_9612,N_2429,N_5775);
xor U9613 (N_9613,N_657,N_5645);
xor U9614 (N_9614,N_4864,N_565);
xor U9615 (N_9615,N_4529,N_1574);
and U9616 (N_9616,N_3838,N_1722);
nand U9617 (N_9617,N_5041,N_82);
nand U9618 (N_9618,N_4414,N_2440);
or U9619 (N_9619,N_2489,N_1978);
xor U9620 (N_9620,N_1868,N_429);
and U9621 (N_9621,N_646,N_2073);
or U9622 (N_9622,N_5949,N_5235);
nor U9623 (N_9623,N_4441,N_2313);
nor U9624 (N_9624,N_534,N_5747);
and U9625 (N_9625,N_4857,N_187);
nand U9626 (N_9626,N_513,N_4727);
and U9627 (N_9627,N_5371,N_5508);
xnor U9628 (N_9628,N_5631,N_3286);
xor U9629 (N_9629,N_1441,N_4887);
or U9630 (N_9630,N_3290,N_4767);
and U9631 (N_9631,N_309,N_5212);
xnor U9632 (N_9632,N_3076,N_3015);
nand U9633 (N_9633,N_2851,N_5491);
or U9634 (N_9634,N_204,N_2806);
xnor U9635 (N_9635,N_5009,N_4519);
and U9636 (N_9636,N_4246,N_283);
and U9637 (N_9637,N_3332,N_3871);
nor U9638 (N_9638,N_1237,N_1083);
or U9639 (N_9639,N_4663,N_3901);
or U9640 (N_9640,N_4709,N_3620);
and U9641 (N_9641,N_2856,N_4398);
or U9642 (N_9642,N_1917,N_835);
and U9643 (N_9643,N_5164,N_3024);
or U9644 (N_9644,N_5675,N_2852);
nand U9645 (N_9645,N_2706,N_3269);
and U9646 (N_9646,N_2374,N_5609);
or U9647 (N_9647,N_4090,N_5504);
or U9648 (N_9648,N_6063,N_4668);
xnor U9649 (N_9649,N_3500,N_2493);
or U9650 (N_9650,N_3973,N_4230);
xor U9651 (N_9651,N_5893,N_2187);
and U9652 (N_9652,N_3864,N_3829);
and U9653 (N_9653,N_1337,N_319);
nand U9654 (N_9654,N_3056,N_1410);
nor U9655 (N_9655,N_2360,N_2928);
xnor U9656 (N_9656,N_1646,N_4492);
nand U9657 (N_9657,N_4503,N_5781);
and U9658 (N_9658,N_5363,N_4390);
nand U9659 (N_9659,N_3315,N_4630);
xnor U9660 (N_9660,N_5209,N_4161);
and U9661 (N_9661,N_5608,N_3784);
nor U9662 (N_9662,N_3443,N_2179);
nor U9663 (N_9663,N_5082,N_2372);
nor U9664 (N_9664,N_2732,N_1265);
and U9665 (N_9665,N_5737,N_876);
xor U9666 (N_9666,N_1570,N_3479);
and U9667 (N_9667,N_1916,N_5056);
and U9668 (N_9668,N_3288,N_2557);
or U9669 (N_9669,N_2030,N_652);
xor U9670 (N_9670,N_968,N_5334);
xor U9671 (N_9671,N_3326,N_2856);
nand U9672 (N_9672,N_367,N_369);
nor U9673 (N_9673,N_5592,N_5719);
nor U9674 (N_9674,N_2385,N_1694);
and U9675 (N_9675,N_4943,N_50);
and U9676 (N_9676,N_5318,N_1211);
nand U9677 (N_9677,N_521,N_2753);
nor U9678 (N_9678,N_2856,N_3702);
or U9679 (N_9679,N_5853,N_3211);
nor U9680 (N_9680,N_3010,N_4436);
nor U9681 (N_9681,N_3394,N_2491);
nand U9682 (N_9682,N_605,N_3831);
or U9683 (N_9683,N_609,N_1177);
and U9684 (N_9684,N_998,N_4880);
nor U9685 (N_9685,N_3771,N_3840);
nand U9686 (N_9686,N_118,N_4695);
and U9687 (N_9687,N_2134,N_1043);
nor U9688 (N_9688,N_1428,N_5612);
xor U9689 (N_9689,N_5021,N_2);
nand U9690 (N_9690,N_3486,N_2692);
xnor U9691 (N_9691,N_1233,N_867);
and U9692 (N_9692,N_5156,N_5541);
and U9693 (N_9693,N_3392,N_4698);
nor U9694 (N_9694,N_4335,N_1284);
xnor U9695 (N_9695,N_249,N_3510);
and U9696 (N_9696,N_3874,N_1119);
or U9697 (N_9697,N_2917,N_973);
or U9698 (N_9698,N_4341,N_2928);
or U9699 (N_9699,N_741,N_161);
or U9700 (N_9700,N_4868,N_4458);
nand U9701 (N_9701,N_1002,N_442);
or U9702 (N_9702,N_4946,N_2811);
nand U9703 (N_9703,N_4686,N_443);
nor U9704 (N_9704,N_1417,N_2682);
xnor U9705 (N_9705,N_324,N_4497);
and U9706 (N_9706,N_2752,N_2486);
xnor U9707 (N_9707,N_4157,N_5898);
and U9708 (N_9708,N_3602,N_2311);
and U9709 (N_9709,N_5744,N_5605);
xor U9710 (N_9710,N_5790,N_99);
nand U9711 (N_9711,N_4401,N_296);
nor U9712 (N_9712,N_6003,N_5378);
nand U9713 (N_9713,N_5756,N_5833);
and U9714 (N_9714,N_1949,N_4557);
and U9715 (N_9715,N_1931,N_3792);
and U9716 (N_9716,N_2408,N_4661);
nor U9717 (N_9717,N_4992,N_5107);
and U9718 (N_9718,N_2676,N_3304);
xor U9719 (N_9719,N_3840,N_4420);
xor U9720 (N_9720,N_4026,N_1863);
and U9721 (N_9721,N_985,N_882);
and U9722 (N_9722,N_2341,N_4875);
nand U9723 (N_9723,N_3383,N_1118);
and U9724 (N_9724,N_112,N_13);
xnor U9725 (N_9725,N_1588,N_2531);
nor U9726 (N_9726,N_4442,N_4606);
and U9727 (N_9727,N_2893,N_5233);
or U9728 (N_9728,N_4315,N_4401);
xnor U9729 (N_9729,N_5876,N_4668);
and U9730 (N_9730,N_2678,N_613);
nor U9731 (N_9731,N_5303,N_5778);
and U9732 (N_9732,N_1260,N_3549);
and U9733 (N_9733,N_5018,N_3421);
nor U9734 (N_9734,N_2942,N_546);
or U9735 (N_9735,N_848,N_2842);
and U9736 (N_9736,N_1978,N_2167);
xnor U9737 (N_9737,N_966,N_5747);
xnor U9738 (N_9738,N_2984,N_3471);
nand U9739 (N_9739,N_726,N_2662);
or U9740 (N_9740,N_5114,N_792);
nor U9741 (N_9741,N_2750,N_6109);
or U9742 (N_9742,N_1597,N_4125);
or U9743 (N_9743,N_1531,N_430);
and U9744 (N_9744,N_265,N_3648);
or U9745 (N_9745,N_4249,N_3761);
xnor U9746 (N_9746,N_897,N_4720);
nand U9747 (N_9747,N_5309,N_5059);
xnor U9748 (N_9748,N_4150,N_1237);
nor U9749 (N_9749,N_3775,N_4292);
or U9750 (N_9750,N_1135,N_1389);
and U9751 (N_9751,N_65,N_851);
nand U9752 (N_9752,N_2542,N_1971);
or U9753 (N_9753,N_5171,N_2936);
and U9754 (N_9754,N_5349,N_4543);
or U9755 (N_9755,N_5071,N_3459);
nand U9756 (N_9756,N_2405,N_3576);
nand U9757 (N_9757,N_1265,N_91);
and U9758 (N_9758,N_5740,N_2572);
nor U9759 (N_9759,N_1976,N_5557);
and U9760 (N_9760,N_188,N_4574);
xnor U9761 (N_9761,N_1484,N_2114);
and U9762 (N_9762,N_3724,N_563);
nand U9763 (N_9763,N_3959,N_6214);
nand U9764 (N_9764,N_3853,N_1652);
or U9765 (N_9765,N_5722,N_986);
and U9766 (N_9766,N_4499,N_5124);
nor U9767 (N_9767,N_1138,N_5647);
xor U9768 (N_9768,N_5463,N_5903);
xor U9769 (N_9769,N_1248,N_2062);
or U9770 (N_9770,N_5862,N_2462);
xor U9771 (N_9771,N_956,N_3390);
and U9772 (N_9772,N_2714,N_75);
nand U9773 (N_9773,N_6124,N_1618);
nor U9774 (N_9774,N_3876,N_5756);
xnor U9775 (N_9775,N_2806,N_5662);
or U9776 (N_9776,N_2000,N_520);
nor U9777 (N_9777,N_551,N_5569);
nand U9778 (N_9778,N_876,N_2344);
and U9779 (N_9779,N_3972,N_1304);
or U9780 (N_9780,N_701,N_2934);
nor U9781 (N_9781,N_2650,N_4730);
or U9782 (N_9782,N_1544,N_4134);
nor U9783 (N_9783,N_2750,N_3759);
or U9784 (N_9784,N_1663,N_5336);
nor U9785 (N_9785,N_469,N_2003);
or U9786 (N_9786,N_88,N_4200);
or U9787 (N_9787,N_3289,N_4164);
nand U9788 (N_9788,N_967,N_5342);
nor U9789 (N_9789,N_6000,N_3958);
and U9790 (N_9790,N_3776,N_2922);
or U9791 (N_9791,N_3497,N_1264);
and U9792 (N_9792,N_17,N_330);
xnor U9793 (N_9793,N_4342,N_6236);
nand U9794 (N_9794,N_2754,N_2151);
and U9795 (N_9795,N_4361,N_2443);
and U9796 (N_9796,N_2532,N_6164);
nor U9797 (N_9797,N_3000,N_3750);
nand U9798 (N_9798,N_3321,N_4931);
nand U9799 (N_9799,N_5590,N_221);
nor U9800 (N_9800,N_4146,N_4785);
xor U9801 (N_9801,N_5639,N_660);
xor U9802 (N_9802,N_6087,N_3679);
nand U9803 (N_9803,N_928,N_3407);
or U9804 (N_9804,N_3190,N_153);
nor U9805 (N_9805,N_3491,N_1769);
or U9806 (N_9806,N_5313,N_2610);
nand U9807 (N_9807,N_1602,N_676);
xor U9808 (N_9808,N_197,N_3908);
nor U9809 (N_9809,N_4633,N_2068);
nor U9810 (N_9810,N_5983,N_546);
nand U9811 (N_9811,N_475,N_1644);
or U9812 (N_9812,N_2161,N_2721);
and U9813 (N_9813,N_4526,N_3750);
nor U9814 (N_9814,N_1434,N_537);
xor U9815 (N_9815,N_2967,N_6127);
and U9816 (N_9816,N_345,N_4166);
and U9817 (N_9817,N_5392,N_5965);
nor U9818 (N_9818,N_2989,N_2033);
nor U9819 (N_9819,N_2200,N_3550);
and U9820 (N_9820,N_117,N_953);
or U9821 (N_9821,N_2646,N_4533);
and U9822 (N_9822,N_3081,N_2272);
and U9823 (N_9823,N_111,N_2486);
nor U9824 (N_9824,N_5904,N_3826);
nor U9825 (N_9825,N_1697,N_5572);
or U9826 (N_9826,N_5099,N_743);
nand U9827 (N_9827,N_3212,N_3872);
nor U9828 (N_9828,N_4316,N_1222);
nand U9829 (N_9829,N_459,N_1971);
nand U9830 (N_9830,N_6001,N_4571);
nor U9831 (N_9831,N_5950,N_2013);
nor U9832 (N_9832,N_5002,N_5665);
nor U9833 (N_9833,N_2768,N_673);
nand U9834 (N_9834,N_497,N_4391);
or U9835 (N_9835,N_5310,N_207);
and U9836 (N_9836,N_4070,N_4770);
nor U9837 (N_9837,N_5716,N_3285);
xnor U9838 (N_9838,N_3526,N_3800);
xor U9839 (N_9839,N_860,N_4209);
and U9840 (N_9840,N_295,N_3971);
nand U9841 (N_9841,N_6230,N_5958);
nor U9842 (N_9842,N_1574,N_1959);
nor U9843 (N_9843,N_1298,N_4549);
nor U9844 (N_9844,N_3491,N_338);
xor U9845 (N_9845,N_1045,N_1300);
nand U9846 (N_9846,N_3126,N_379);
nor U9847 (N_9847,N_4880,N_2134);
nand U9848 (N_9848,N_2613,N_5836);
nand U9849 (N_9849,N_809,N_4646);
nor U9850 (N_9850,N_151,N_3201);
nor U9851 (N_9851,N_397,N_5531);
xnor U9852 (N_9852,N_1940,N_6060);
and U9853 (N_9853,N_769,N_5444);
nand U9854 (N_9854,N_1018,N_5935);
nand U9855 (N_9855,N_3825,N_0);
xor U9856 (N_9856,N_666,N_263);
and U9857 (N_9857,N_4676,N_849);
nand U9858 (N_9858,N_5512,N_2795);
xor U9859 (N_9859,N_4458,N_292);
and U9860 (N_9860,N_780,N_3831);
or U9861 (N_9861,N_4222,N_905);
or U9862 (N_9862,N_4043,N_878);
or U9863 (N_9863,N_536,N_4349);
nand U9864 (N_9864,N_210,N_2622);
and U9865 (N_9865,N_4291,N_3454);
and U9866 (N_9866,N_756,N_1849);
nand U9867 (N_9867,N_2183,N_740);
and U9868 (N_9868,N_4202,N_3505);
or U9869 (N_9869,N_4442,N_322);
nand U9870 (N_9870,N_540,N_4624);
nor U9871 (N_9871,N_1596,N_4574);
or U9872 (N_9872,N_5317,N_5309);
nor U9873 (N_9873,N_5230,N_4104);
and U9874 (N_9874,N_4849,N_47);
and U9875 (N_9875,N_1168,N_4038);
nor U9876 (N_9876,N_1078,N_5941);
and U9877 (N_9877,N_5276,N_4017);
nand U9878 (N_9878,N_4054,N_16);
and U9879 (N_9879,N_1061,N_1613);
or U9880 (N_9880,N_2409,N_5038);
nor U9881 (N_9881,N_4511,N_1536);
nor U9882 (N_9882,N_3267,N_5216);
and U9883 (N_9883,N_5153,N_418);
nand U9884 (N_9884,N_538,N_5192);
nand U9885 (N_9885,N_667,N_27);
nor U9886 (N_9886,N_1894,N_524);
or U9887 (N_9887,N_5253,N_6124);
xor U9888 (N_9888,N_54,N_3138);
and U9889 (N_9889,N_2069,N_959);
xnor U9890 (N_9890,N_3969,N_5142);
or U9891 (N_9891,N_1953,N_979);
nor U9892 (N_9892,N_3025,N_6176);
nor U9893 (N_9893,N_2565,N_4346);
and U9894 (N_9894,N_4631,N_193);
nand U9895 (N_9895,N_3991,N_4393);
or U9896 (N_9896,N_444,N_6165);
and U9897 (N_9897,N_53,N_3748);
or U9898 (N_9898,N_3401,N_1254);
and U9899 (N_9899,N_5141,N_2770);
nand U9900 (N_9900,N_2735,N_6205);
or U9901 (N_9901,N_1440,N_4070);
nand U9902 (N_9902,N_4783,N_3893);
nor U9903 (N_9903,N_2235,N_3621);
nor U9904 (N_9904,N_1166,N_2671);
and U9905 (N_9905,N_1647,N_2247);
nor U9906 (N_9906,N_3055,N_1867);
nor U9907 (N_9907,N_781,N_4702);
nand U9908 (N_9908,N_4898,N_2257);
xnor U9909 (N_9909,N_6042,N_5380);
or U9910 (N_9910,N_1663,N_937);
nor U9911 (N_9911,N_1602,N_5329);
xnor U9912 (N_9912,N_4294,N_3367);
and U9913 (N_9913,N_3309,N_1972);
nor U9914 (N_9914,N_2123,N_4518);
and U9915 (N_9915,N_4786,N_5400);
or U9916 (N_9916,N_2209,N_2022);
and U9917 (N_9917,N_4232,N_2959);
xor U9918 (N_9918,N_3921,N_5304);
nor U9919 (N_9919,N_107,N_367);
nand U9920 (N_9920,N_2886,N_5567);
nand U9921 (N_9921,N_3755,N_2885);
nand U9922 (N_9922,N_4950,N_1188);
and U9923 (N_9923,N_5644,N_958);
xnor U9924 (N_9924,N_2053,N_4227);
xor U9925 (N_9925,N_4032,N_360);
and U9926 (N_9926,N_6069,N_2436);
nor U9927 (N_9927,N_2461,N_4006);
xnor U9928 (N_9928,N_974,N_159);
or U9929 (N_9929,N_4903,N_2494);
nand U9930 (N_9930,N_5649,N_5753);
xor U9931 (N_9931,N_3189,N_1908);
nand U9932 (N_9932,N_2887,N_1147);
and U9933 (N_9933,N_1713,N_2616);
nand U9934 (N_9934,N_5577,N_1687);
and U9935 (N_9935,N_2291,N_6049);
and U9936 (N_9936,N_2998,N_1173);
nor U9937 (N_9937,N_2295,N_42);
nand U9938 (N_9938,N_2625,N_4060);
and U9939 (N_9939,N_2757,N_4340);
nor U9940 (N_9940,N_5443,N_2139);
nand U9941 (N_9941,N_2400,N_155);
nor U9942 (N_9942,N_5021,N_395);
or U9943 (N_9943,N_515,N_5988);
nand U9944 (N_9944,N_2471,N_2239);
nand U9945 (N_9945,N_537,N_2141);
xor U9946 (N_9946,N_4309,N_2747);
and U9947 (N_9947,N_872,N_1826);
nand U9948 (N_9948,N_3106,N_2670);
xor U9949 (N_9949,N_1754,N_2260);
nand U9950 (N_9950,N_4312,N_2599);
nand U9951 (N_9951,N_4756,N_5193);
nor U9952 (N_9952,N_5747,N_485);
xor U9953 (N_9953,N_3444,N_3944);
xnor U9954 (N_9954,N_157,N_636);
xnor U9955 (N_9955,N_5036,N_6059);
xnor U9956 (N_9956,N_2505,N_214);
nand U9957 (N_9957,N_892,N_5907);
nor U9958 (N_9958,N_1945,N_4006);
and U9959 (N_9959,N_3548,N_1486);
xor U9960 (N_9960,N_2924,N_2813);
xnor U9961 (N_9961,N_18,N_3005);
xor U9962 (N_9962,N_5621,N_5841);
and U9963 (N_9963,N_3036,N_29);
or U9964 (N_9964,N_4087,N_2068);
nand U9965 (N_9965,N_4229,N_566);
nor U9966 (N_9966,N_736,N_2563);
or U9967 (N_9967,N_3420,N_2872);
nand U9968 (N_9968,N_95,N_2840);
xor U9969 (N_9969,N_124,N_5921);
and U9970 (N_9970,N_710,N_4302);
xnor U9971 (N_9971,N_4919,N_2236);
nor U9972 (N_9972,N_3059,N_3328);
xnor U9973 (N_9973,N_797,N_4515);
xnor U9974 (N_9974,N_3957,N_4678);
nor U9975 (N_9975,N_70,N_5502);
xnor U9976 (N_9976,N_6040,N_5180);
or U9977 (N_9977,N_5492,N_3219);
nor U9978 (N_9978,N_4678,N_2582);
nor U9979 (N_9979,N_421,N_337);
nand U9980 (N_9980,N_3315,N_4972);
nand U9981 (N_9981,N_4296,N_5652);
or U9982 (N_9982,N_1340,N_2682);
nand U9983 (N_9983,N_3787,N_5176);
nand U9984 (N_9984,N_414,N_942);
and U9985 (N_9985,N_5573,N_5771);
and U9986 (N_9986,N_1814,N_4123);
and U9987 (N_9987,N_3857,N_5103);
xnor U9988 (N_9988,N_5380,N_1042);
and U9989 (N_9989,N_4202,N_1270);
or U9990 (N_9990,N_476,N_3919);
and U9991 (N_9991,N_4491,N_1736);
nand U9992 (N_9992,N_3527,N_1046);
nand U9993 (N_9993,N_6078,N_4085);
or U9994 (N_9994,N_3606,N_3009);
nand U9995 (N_9995,N_5295,N_4794);
nor U9996 (N_9996,N_1762,N_2806);
nor U9997 (N_9997,N_4533,N_2876);
nand U9998 (N_9998,N_1390,N_2042);
nor U9999 (N_9999,N_5983,N_3955);
or U10000 (N_10000,N_25,N_3985);
and U10001 (N_10001,N_3705,N_1283);
xnor U10002 (N_10002,N_1711,N_4030);
xnor U10003 (N_10003,N_1880,N_4832);
nor U10004 (N_10004,N_3088,N_3069);
or U10005 (N_10005,N_2808,N_1014);
or U10006 (N_10006,N_1031,N_4588);
or U10007 (N_10007,N_5500,N_3546);
or U10008 (N_10008,N_466,N_372);
nor U10009 (N_10009,N_5843,N_5071);
nand U10010 (N_10010,N_4359,N_1986);
nor U10011 (N_10011,N_5263,N_97);
xor U10012 (N_10012,N_2261,N_4877);
xnor U10013 (N_10013,N_3843,N_4551);
and U10014 (N_10014,N_3903,N_397);
nand U10015 (N_10015,N_5473,N_3505);
nor U10016 (N_10016,N_930,N_3391);
nand U10017 (N_10017,N_717,N_2894);
and U10018 (N_10018,N_3131,N_4315);
nand U10019 (N_10019,N_5443,N_699);
xor U10020 (N_10020,N_1094,N_4633);
and U10021 (N_10021,N_4170,N_882);
or U10022 (N_10022,N_6240,N_3918);
and U10023 (N_10023,N_3541,N_3971);
nor U10024 (N_10024,N_4174,N_3645);
or U10025 (N_10025,N_1152,N_2096);
or U10026 (N_10026,N_221,N_4570);
and U10027 (N_10027,N_1415,N_4219);
and U10028 (N_10028,N_2928,N_2648);
nand U10029 (N_10029,N_2353,N_3522);
nor U10030 (N_10030,N_2213,N_2966);
xor U10031 (N_10031,N_4148,N_1573);
or U10032 (N_10032,N_2456,N_5786);
and U10033 (N_10033,N_5372,N_3285);
or U10034 (N_10034,N_2749,N_4447);
and U10035 (N_10035,N_1782,N_3051);
nand U10036 (N_10036,N_4613,N_2695);
or U10037 (N_10037,N_2824,N_3516);
nand U10038 (N_10038,N_1215,N_2979);
and U10039 (N_10039,N_62,N_91);
nand U10040 (N_10040,N_211,N_4113);
xor U10041 (N_10041,N_3946,N_160);
or U10042 (N_10042,N_588,N_6231);
or U10043 (N_10043,N_4457,N_3761);
nand U10044 (N_10044,N_3139,N_1109);
nand U10045 (N_10045,N_4880,N_2286);
nor U10046 (N_10046,N_308,N_1393);
and U10047 (N_10047,N_5998,N_35);
xnor U10048 (N_10048,N_3207,N_3195);
and U10049 (N_10049,N_4600,N_2842);
or U10050 (N_10050,N_1753,N_3773);
or U10051 (N_10051,N_2789,N_1926);
nand U10052 (N_10052,N_1326,N_2284);
nand U10053 (N_10053,N_1080,N_3042);
nand U10054 (N_10054,N_657,N_2341);
nor U10055 (N_10055,N_759,N_3654);
nand U10056 (N_10056,N_2427,N_747);
or U10057 (N_10057,N_1030,N_1031);
and U10058 (N_10058,N_3592,N_2696);
nand U10059 (N_10059,N_2926,N_5008);
and U10060 (N_10060,N_3012,N_4445);
or U10061 (N_10061,N_274,N_4423);
nor U10062 (N_10062,N_1925,N_2479);
nand U10063 (N_10063,N_2513,N_510);
xor U10064 (N_10064,N_2684,N_3504);
or U10065 (N_10065,N_2805,N_3563);
nor U10066 (N_10066,N_2406,N_501);
nor U10067 (N_10067,N_4107,N_2497);
xnor U10068 (N_10068,N_3462,N_5479);
and U10069 (N_10069,N_3049,N_4287);
and U10070 (N_10070,N_4307,N_5787);
nor U10071 (N_10071,N_5831,N_1264);
xnor U10072 (N_10072,N_4140,N_5367);
or U10073 (N_10073,N_1020,N_4240);
nand U10074 (N_10074,N_2451,N_3466);
nor U10075 (N_10075,N_4154,N_5761);
nand U10076 (N_10076,N_505,N_929);
nand U10077 (N_10077,N_4449,N_4863);
and U10078 (N_10078,N_3554,N_3471);
and U10079 (N_10079,N_3029,N_3252);
nand U10080 (N_10080,N_1812,N_66);
nand U10081 (N_10081,N_1760,N_5202);
and U10082 (N_10082,N_6230,N_737);
xnor U10083 (N_10083,N_648,N_2708);
nor U10084 (N_10084,N_1060,N_5231);
nand U10085 (N_10085,N_4410,N_1081);
nand U10086 (N_10086,N_4823,N_3924);
and U10087 (N_10087,N_1514,N_1908);
or U10088 (N_10088,N_3668,N_5825);
nor U10089 (N_10089,N_5502,N_4646);
nor U10090 (N_10090,N_2674,N_3447);
and U10091 (N_10091,N_4721,N_2538);
nor U10092 (N_10092,N_5142,N_2801);
nand U10093 (N_10093,N_4142,N_2961);
or U10094 (N_10094,N_2365,N_5289);
xor U10095 (N_10095,N_4316,N_4924);
nor U10096 (N_10096,N_4323,N_1268);
xnor U10097 (N_10097,N_486,N_1338);
and U10098 (N_10098,N_2820,N_5059);
xnor U10099 (N_10099,N_4577,N_480);
nand U10100 (N_10100,N_3021,N_360);
nor U10101 (N_10101,N_1606,N_1680);
and U10102 (N_10102,N_3483,N_3564);
nor U10103 (N_10103,N_472,N_92);
and U10104 (N_10104,N_5505,N_3936);
nand U10105 (N_10105,N_660,N_4229);
xnor U10106 (N_10106,N_5535,N_157);
xor U10107 (N_10107,N_3156,N_169);
or U10108 (N_10108,N_1458,N_5346);
or U10109 (N_10109,N_3734,N_101);
nor U10110 (N_10110,N_6217,N_1189);
and U10111 (N_10111,N_1572,N_4269);
or U10112 (N_10112,N_6003,N_4994);
or U10113 (N_10113,N_6008,N_1896);
nor U10114 (N_10114,N_3411,N_3815);
xor U10115 (N_10115,N_423,N_2534);
or U10116 (N_10116,N_5205,N_1441);
xor U10117 (N_10117,N_820,N_476);
or U10118 (N_10118,N_6047,N_174);
nor U10119 (N_10119,N_590,N_3264);
or U10120 (N_10120,N_3590,N_2942);
or U10121 (N_10121,N_4979,N_5028);
nand U10122 (N_10122,N_4140,N_4635);
and U10123 (N_10123,N_4816,N_3453);
xnor U10124 (N_10124,N_2485,N_2814);
or U10125 (N_10125,N_5434,N_726);
nand U10126 (N_10126,N_1586,N_3208);
and U10127 (N_10127,N_4170,N_4627);
nor U10128 (N_10128,N_799,N_5381);
xor U10129 (N_10129,N_84,N_5878);
nand U10130 (N_10130,N_1370,N_3887);
nor U10131 (N_10131,N_2586,N_5576);
xnor U10132 (N_10132,N_914,N_4341);
xor U10133 (N_10133,N_1943,N_2101);
or U10134 (N_10134,N_4090,N_2342);
nor U10135 (N_10135,N_5526,N_1847);
or U10136 (N_10136,N_3849,N_3715);
and U10137 (N_10137,N_1153,N_1359);
nor U10138 (N_10138,N_819,N_3721);
nor U10139 (N_10139,N_3132,N_1530);
or U10140 (N_10140,N_4126,N_1661);
nand U10141 (N_10141,N_6121,N_5375);
nor U10142 (N_10142,N_2289,N_456);
or U10143 (N_10143,N_5745,N_349);
xnor U10144 (N_10144,N_48,N_4275);
or U10145 (N_10145,N_3735,N_4965);
and U10146 (N_10146,N_5404,N_1369);
nand U10147 (N_10147,N_2304,N_3740);
nand U10148 (N_10148,N_2150,N_5119);
or U10149 (N_10149,N_1788,N_2565);
nor U10150 (N_10150,N_863,N_2762);
nor U10151 (N_10151,N_1469,N_3469);
nand U10152 (N_10152,N_5714,N_4121);
and U10153 (N_10153,N_1460,N_878);
nor U10154 (N_10154,N_5711,N_2271);
xnor U10155 (N_10155,N_4087,N_4468);
xor U10156 (N_10156,N_784,N_102);
or U10157 (N_10157,N_1018,N_450);
and U10158 (N_10158,N_1750,N_2266);
nor U10159 (N_10159,N_1249,N_3872);
xor U10160 (N_10160,N_2071,N_5792);
or U10161 (N_10161,N_4005,N_591);
xor U10162 (N_10162,N_4858,N_6061);
xnor U10163 (N_10163,N_5089,N_604);
and U10164 (N_10164,N_181,N_4087);
nor U10165 (N_10165,N_5314,N_3465);
and U10166 (N_10166,N_6134,N_4923);
or U10167 (N_10167,N_4560,N_2717);
xor U10168 (N_10168,N_3709,N_2704);
nand U10169 (N_10169,N_1242,N_5931);
nand U10170 (N_10170,N_5377,N_5614);
xnor U10171 (N_10171,N_5299,N_1390);
nor U10172 (N_10172,N_4686,N_2737);
or U10173 (N_10173,N_71,N_4219);
nand U10174 (N_10174,N_5866,N_2150);
nor U10175 (N_10175,N_3912,N_5591);
or U10176 (N_10176,N_1579,N_5524);
and U10177 (N_10177,N_5215,N_1233);
and U10178 (N_10178,N_1477,N_3916);
nand U10179 (N_10179,N_2664,N_37);
nand U10180 (N_10180,N_5917,N_2113);
and U10181 (N_10181,N_3078,N_31);
or U10182 (N_10182,N_1976,N_1126);
nand U10183 (N_10183,N_1199,N_2359);
and U10184 (N_10184,N_2931,N_4504);
xnor U10185 (N_10185,N_4127,N_916);
nand U10186 (N_10186,N_867,N_4665);
and U10187 (N_10187,N_2582,N_2180);
and U10188 (N_10188,N_6245,N_1350);
and U10189 (N_10189,N_969,N_4271);
xor U10190 (N_10190,N_2074,N_783);
or U10191 (N_10191,N_4110,N_6230);
and U10192 (N_10192,N_3244,N_6208);
and U10193 (N_10193,N_6123,N_2634);
xor U10194 (N_10194,N_939,N_3546);
and U10195 (N_10195,N_2911,N_3559);
xnor U10196 (N_10196,N_3822,N_2315);
xor U10197 (N_10197,N_210,N_3507);
nor U10198 (N_10198,N_1900,N_219);
xor U10199 (N_10199,N_2021,N_3851);
nor U10200 (N_10200,N_969,N_632);
nor U10201 (N_10201,N_1709,N_4417);
nor U10202 (N_10202,N_2256,N_5386);
nand U10203 (N_10203,N_3480,N_861);
nand U10204 (N_10204,N_65,N_3900);
or U10205 (N_10205,N_2362,N_5605);
nand U10206 (N_10206,N_4922,N_1819);
or U10207 (N_10207,N_1257,N_5343);
and U10208 (N_10208,N_1030,N_1882);
xor U10209 (N_10209,N_1063,N_1330);
and U10210 (N_10210,N_2297,N_2372);
nand U10211 (N_10211,N_6121,N_199);
xor U10212 (N_10212,N_891,N_410);
or U10213 (N_10213,N_5467,N_1035);
nor U10214 (N_10214,N_5054,N_223);
nand U10215 (N_10215,N_3504,N_5681);
nand U10216 (N_10216,N_6078,N_4511);
xor U10217 (N_10217,N_910,N_2979);
or U10218 (N_10218,N_6170,N_4849);
and U10219 (N_10219,N_886,N_3718);
nor U10220 (N_10220,N_3446,N_2352);
or U10221 (N_10221,N_2396,N_5388);
nand U10222 (N_10222,N_65,N_3183);
xnor U10223 (N_10223,N_5721,N_1635);
or U10224 (N_10224,N_5459,N_1278);
nand U10225 (N_10225,N_939,N_1766);
xor U10226 (N_10226,N_1783,N_1935);
or U10227 (N_10227,N_2028,N_368);
nor U10228 (N_10228,N_4875,N_6221);
nand U10229 (N_10229,N_3519,N_4567);
or U10230 (N_10230,N_3664,N_3806);
nand U10231 (N_10231,N_3212,N_2623);
nor U10232 (N_10232,N_514,N_4467);
and U10233 (N_10233,N_5247,N_3437);
nor U10234 (N_10234,N_3404,N_5041);
xor U10235 (N_10235,N_5592,N_1802);
and U10236 (N_10236,N_5235,N_6077);
and U10237 (N_10237,N_1835,N_2062);
nor U10238 (N_10238,N_1985,N_3243);
or U10239 (N_10239,N_3578,N_1914);
or U10240 (N_10240,N_3051,N_2166);
and U10241 (N_10241,N_1428,N_4226);
xnor U10242 (N_10242,N_6136,N_4823);
or U10243 (N_10243,N_4155,N_252);
nor U10244 (N_10244,N_1210,N_3740);
and U10245 (N_10245,N_5737,N_4337);
and U10246 (N_10246,N_2468,N_5890);
nand U10247 (N_10247,N_2375,N_3668);
nor U10248 (N_10248,N_348,N_225);
or U10249 (N_10249,N_2078,N_3675);
nor U10250 (N_10250,N_355,N_2900);
or U10251 (N_10251,N_4602,N_1187);
nor U10252 (N_10252,N_4819,N_2675);
xnor U10253 (N_10253,N_3379,N_1405);
nor U10254 (N_10254,N_6169,N_3580);
or U10255 (N_10255,N_3524,N_107);
nor U10256 (N_10256,N_5070,N_4214);
or U10257 (N_10257,N_1948,N_5852);
nor U10258 (N_10258,N_1662,N_571);
nor U10259 (N_10259,N_2149,N_5923);
nor U10260 (N_10260,N_72,N_1495);
and U10261 (N_10261,N_2309,N_5226);
and U10262 (N_10262,N_3459,N_3309);
nand U10263 (N_10263,N_4374,N_5773);
and U10264 (N_10264,N_2543,N_3742);
and U10265 (N_10265,N_847,N_55);
nor U10266 (N_10266,N_2475,N_4093);
and U10267 (N_10267,N_6202,N_6061);
and U10268 (N_10268,N_714,N_5786);
and U10269 (N_10269,N_2843,N_5610);
or U10270 (N_10270,N_2849,N_3611);
nand U10271 (N_10271,N_6142,N_3915);
xor U10272 (N_10272,N_4636,N_2639);
or U10273 (N_10273,N_3818,N_1575);
and U10274 (N_10274,N_177,N_4980);
and U10275 (N_10275,N_2918,N_195);
or U10276 (N_10276,N_3495,N_5533);
or U10277 (N_10277,N_2585,N_559);
nor U10278 (N_10278,N_3733,N_2710);
nor U10279 (N_10279,N_3329,N_2537);
nand U10280 (N_10280,N_3147,N_2276);
nand U10281 (N_10281,N_491,N_495);
and U10282 (N_10282,N_958,N_2709);
nor U10283 (N_10283,N_5799,N_510);
xnor U10284 (N_10284,N_4829,N_5131);
and U10285 (N_10285,N_179,N_4753);
and U10286 (N_10286,N_2679,N_5071);
nor U10287 (N_10287,N_6235,N_5247);
nor U10288 (N_10288,N_3700,N_5565);
nor U10289 (N_10289,N_2515,N_4394);
nand U10290 (N_10290,N_754,N_5615);
or U10291 (N_10291,N_3872,N_4412);
or U10292 (N_10292,N_6096,N_4231);
nand U10293 (N_10293,N_2880,N_5913);
nand U10294 (N_10294,N_5503,N_140);
nand U10295 (N_10295,N_5706,N_4989);
xnor U10296 (N_10296,N_3938,N_2433);
xnor U10297 (N_10297,N_3538,N_5229);
and U10298 (N_10298,N_447,N_3678);
xor U10299 (N_10299,N_5951,N_3117);
or U10300 (N_10300,N_2665,N_6099);
xnor U10301 (N_10301,N_5960,N_302);
nand U10302 (N_10302,N_2581,N_4743);
nand U10303 (N_10303,N_5222,N_5917);
xor U10304 (N_10304,N_2269,N_5170);
and U10305 (N_10305,N_2188,N_4810);
nor U10306 (N_10306,N_4618,N_1156);
xnor U10307 (N_10307,N_1136,N_2886);
nor U10308 (N_10308,N_699,N_2118);
xor U10309 (N_10309,N_3037,N_2407);
xnor U10310 (N_10310,N_3332,N_5666);
and U10311 (N_10311,N_519,N_6052);
nor U10312 (N_10312,N_4457,N_2762);
xnor U10313 (N_10313,N_1605,N_3888);
and U10314 (N_10314,N_1411,N_2402);
and U10315 (N_10315,N_2295,N_5710);
and U10316 (N_10316,N_4758,N_2967);
nand U10317 (N_10317,N_5944,N_590);
xor U10318 (N_10318,N_3075,N_4248);
and U10319 (N_10319,N_2537,N_4802);
and U10320 (N_10320,N_2798,N_3423);
xor U10321 (N_10321,N_4768,N_743);
nand U10322 (N_10322,N_3349,N_2968);
and U10323 (N_10323,N_2930,N_6182);
and U10324 (N_10324,N_2835,N_2139);
xnor U10325 (N_10325,N_3716,N_5657);
nand U10326 (N_10326,N_3233,N_3720);
and U10327 (N_10327,N_4751,N_4591);
nor U10328 (N_10328,N_4993,N_5448);
nand U10329 (N_10329,N_1348,N_6011);
or U10330 (N_10330,N_4804,N_4655);
nor U10331 (N_10331,N_135,N_3969);
or U10332 (N_10332,N_3324,N_6095);
xnor U10333 (N_10333,N_1348,N_3765);
or U10334 (N_10334,N_3532,N_2685);
or U10335 (N_10335,N_5060,N_3668);
and U10336 (N_10336,N_4921,N_4603);
xnor U10337 (N_10337,N_3204,N_338);
and U10338 (N_10338,N_297,N_4964);
and U10339 (N_10339,N_4439,N_181);
nor U10340 (N_10340,N_1150,N_895);
nor U10341 (N_10341,N_916,N_3710);
and U10342 (N_10342,N_2113,N_5504);
nand U10343 (N_10343,N_5034,N_3786);
nor U10344 (N_10344,N_5511,N_5958);
nand U10345 (N_10345,N_1606,N_4495);
nor U10346 (N_10346,N_3670,N_5828);
and U10347 (N_10347,N_3813,N_121);
nor U10348 (N_10348,N_5055,N_1083);
xor U10349 (N_10349,N_5684,N_5084);
and U10350 (N_10350,N_3607,N_534);
nor U10351 (N_10351,N_2913,N_1065);
nor U10352 (N_10352,N_1927,N_905);
nand U10353 (N_10353,N_3056,N_2224);
or U10354 (N_10354,N_6070,N_3997);
nor U10355 (N_10355,N_4806,N_753);
nand U10356 (N_10356,N_5945,N_52);
nor U10357 (N_10357,N_3866,N_5215);
nor U10358 (N_10358,N_4391,N_4646);
nand U10359 (N_10359,N_4592,N_1484);
xor U10360 (N_10360,N_1834,N_2836);
xor U10361 (N_10361,N_5477,N_6088);
xor U10362 (N_10362,N_6240,N_398);
and U10363 (N_10363,N_2657,N_829);
nor U10364 (N_10364,N_5917,N_4486);
or U10365 (N_10365,N_1910,N_5043);
nand U10366 (N_10366,N_4228,N_5138);
and U10367 (N_10367,N_4209,N_15);
xnor U10368 (N_10368,N_4903,N_2868);
nand U10369 (N_10369,N_4526,N_3597);
nor U10370 (N_10370,N_4363,N_4170);
or U10371 (N_10371,N_3823,N_3898);
and U10372 (N_10372,N_4070,N_2800);
nor U10373 (N_10373,N_6087,N_1458);
nor U10374 (N_10374,N_5093,N_5380);
or U10375 (N_10375,N_3246,N_2998);
and U10376 (N_10376,N_6002,N_5276);
nor U10377 (N_10377,N_1821,N_2770);
or U10378 (N_10378,N_1345,N_152);
nand U10379 (N_10379,N_2240,N_624);
nand U10380 (N_10380,N_3388,N_3769);
xnor U10381 (N_10381,N_2793,N_4646);
or U10382 (N_10382,N_3178,N_2047);
nand U10383 (N_10383,N_2482,N_5342);
xnor U10384 (N_10384,N_5727,N_892);
xor U10385 (N_10385,N_4818,N_313);
nand U10386 (N_10386,N_2661,N_4921);
and U10387 (N_10387,N_3564,N_3435);
and U10388 (N_10388,N_3722,N_5326);
xnor U10389 (N_10389,N_3042,N_4335);
nor U10390 (N_10390,N_5766,N_5549);
or U10391 (N_10391,N_6148,N_2105);
or U10392 (N_10392,N_4507,N_4285);
or U10393 (N_10393,N_1961,N_5126);
nand U10394 (N_10394,N_3753,N_3528);
and U10395 (N_10395,N_2236,N_969);
nand U10396 (N_10396,N_4543,N_215);
xnor U10397 (N_10397,N_1979,N_5093);
nand U10398 (N_10398,N_5947,N_1334);
and U10399 (N_10399,N_5181,N_2670);
or U10400 (N_10400,N_5081,N_4637);
and U10401 (N_10401,N_2369,N_426);
or U10402 (N_10402,N_3372,N_2953);
or U10403 (N_10403,N_2518,N_2916);
nand U10404 (N_10404,N_305,N_5380);
or U10405 (N_10405,N_2873,N_3751);
or U10406 (N_10406,N_1382,N_3493);
nor U10407 (N_10407,N_6220,N_5925);
or U10408 (N_10408,N_4083,N_5896);
or U10409 (N_10409,N_1594,N_1964);
nor U10410 (N_10410,N_3480,N_4819);
nor U10411 (N_10411,N_4125,N_2377);
and U10412 (N_10412,N_149,N_2321);
nor U10413 (N_10413,N_2165,N_2769);
or U10414 (N_10414,N_4392,N_5527);
nor U10415 (N_10415,N_6135,N_4811);
nor U10416 (N_10416,N_3779,N_3177);
or U10417 (N_10417,N_4321,N_4757);
and U10418 (N_10418,N_2432,N_396);
nand U10419 (N_10419,N_2368,N_5740);
nand U10420 (N_10420,N_187,N_5990);
or U10421 (N_10421,N_1269,N_6120);
xor U10422 (N_10422,N_2419,N_6035);
xor U10423 (N_10423,N_664,N_392);
nor U10424 (N_10424,N_5062,N_4602);
and U10425 (N_10425,N_5077,N_1765);
nand U10426 (N_10426,N_4807,N_5779);
or U10427 (N_10427,N_1251,N_2052);
or U10428 (N_10428,N_4667,N_4680);
xnor U10429 (N_10429,N_3364,N_5706);
nand U10430 (N_10430,N_6168,N_118);
nor U10431 (N_10431,N_193,N_4210);
nor U10432 (N_10432,N_304,N_2226);
or U10433 (N_10433,N_744,N_155);
nor U10434 (N_10434,N_472,N_1569);
nor U10435 (N_10435,N_1256,N_5784);
or U10436 (N_10436,N_5329,N_6098);
nor U10437 (N_10437,N_5812,N_2838);
xor U10438 (N_10438,N_886,N_3000);
or U10439 (N_10439,N_5803,N_5655);
or U10440 (N_10440,N_1714,N_2877);
nand U10441 (N_10441,N_4934,N_4397);
xnor U10442 (N_10442,N_441,N_1658);
nor U10443 (N_10443,N_1153,N_1785);
or U10444 (N_10444,N_3744,N_448);
or U10445 (N_10445,N_2412,N_356);
or U10446 (N_10446,N_2504,N_4552);
nor U10447 (N_10447,N_1692,N_47);
nor U10448 (N_10448,N_107,N_728);
nor U10449 (N_10449,N_4669,N_1812);
xor U10450 (N_10450,N_817,N_1599);
nor U10451 (N_10451,N_1997,N_2438);
and U10452 (N_10452,N_3124,N_2032);
xor U10453 (N_10453,N_5920,N_1966);
nand U10454 (N_10454,N_1012,N_1374);
xnor U10455 (N_10455,N_1133,N_3753);
nor U10456 (N_10456,N_4335,N_470);
xor U10457 (N_10457,N_2081,N_470);
or U10458 (N_10458,N_383,N_6059);
nor U10459 (N_10459,N_777,N_2391);
nor U10460 (N_10460,N_2586,N_1347);
nor U10461 (N_10461,N_1921,N_1547);
nor U10462 (N_10462,N_5534,N_3458);
xnor U10463 (N_10463,N_2509,N_257);
or U10464 (N_10464,N_1782,N_2890);
and U10465 (N_10465,N_5022,N_5832);
or U10466 (N_10466,N_3714,N_4661);
or U10467 (N_10467,N_1539,N_4762);
and U10468 (N_10468,N_2019,N_3654);
nand U10469 (N_10469,N_3599,N_2996);
nor U10470 (N_10470,N_538,N_1383);
nor U10471 (N_10471,N_790,N_5014);
nand U10472 (N_10472,N_2003,N_826);
nor U10473 (N_10473,N_2567,N_4897);
and U10474 (N_10474,N_6139,N_297);
and U10475 (N_10475,N_669,N_960);
nand U10476 (N_10476,N_3154,N_4580);
or U10477 (N_10477,N_3136,N_960);
xnor U10478 (N_10478,N_580,N_1229);
and U10479 (N_10479,N_4046,N_3081);
and U10480 (N_10480,N_3931,N_2006);
xor U10481 (N_10481,N_119,N_2154);
nor U10482 (N_10482,N_6017,N_2428);
and U10483 (N_10483,N_3708,N_3285);
xor U10484 (N_10484,N_1844,N_3066);
xnor U10485 (N_10485,N_1548,N_3598);
xor U10486 (N_10486,N_4545,N_3661);
xnor U10487 (N_10487,N_1331,N_4405);
xnor U10488 (N_10488,N_4912,N_5626);
nor U10489 (N_10489,N_2439,N_1170);
and U10490 (N_10490,N_1230,N_3769);
and U10491 (N_10491,N_5230,N_2708);
nand U10492 (N_10492,N_3508,N_2500);
nor U10493 (N_10493,N_761,N_2607);
nor U10494 (N_10494,N_2110,N_5295);
or U10495 (N_10495,N_4030,N_753);
xor U10496 (N_10496,N_1106,N_4506);
or U10497 (N_10497,N_6073,N_5607);
and U10498 (N_10498,N_2387,N_4256);
and U10499 (N_10499,N_2257,N_2027);
or U10500 (N_10500,N_2767,N_5736);
xnor U10501 (N_10501,N_5498,N_1313);
and U10502 (N_10502,N_538,N_300);
and U10503 (N_10503,N_3112,N_5875);
or U10504 (N_10504,N_5605,N_2954);
nor U10505 (N_10505,N_2961,N_771);
or U10506 (N_10506,N_2831,N_4973);
xnor U10507 (N_10507,N_893,N_2663);
nand U10508 (N_10508,N_4888,N_1236);
and U10509 (N_10509,N_2904,N_2789);
xor U10510 (N_10510,N_5403,N_5075);
nor U10511 (N_10511,N_3184,N_374);
nand U10512 (N_10512,N_2134,N_3055);
nor U10513 (N_10513,N_4309,N_2388);
and U10514 (N_10514,N_1555,N_3961);
xnor U10515 (N_10515,N_4731,N_5928);
or U10516 (N_10516,N_4095,N_4829);
nand U10517 (N_10517,N_5145,N_5415);
nand U10518 (N_10518,N_6113,N_1835);
nand U10519 (N_10519,N_2197,N_6186);
nand U10520 (N_10520,N_4182,N_3315);
nor U10521 (N_10521,N_215,N_457);
or U10522 (N_10522,N_4542,N_5756);
and U10523 (N_10523,N_3052,N_3945);
and U10524 (N_10524,N_4834,N_1857);
and U10525 (N_10525,N_3179,N_0);
xnor U10526 (N_10526,N_3138,N_1233);
xor U10527 (N_10527,N_4277,N_4630);
nor U10528 (N_10528,N_1094,N_5530);
xnor U10529 (N_10529,N_3980,N_6170);
or U10530 (N_10530,N_4588,N_957);
and U10531 (N_10531,N_4820,N_2577);
or U10532 (N_10532,N_5034,N_5716);
nand U10533 (N_10533,N_1368,N_2121);
or U10534 (N_10534,N_1877,N_4527);
or U10535 (N_10535,N_2508,N_4827);
xor U10536 (N_10536,N_2871,N_2110);
nand U10537 (N_10537,N_139,N_3531);
or U10538 (N_10538,N_3028,N_264);
or U10539 (N_10539,N_4345,N_4690);
nand U10540 (N_10540,N_2591,N_761);
or U10541 (N_10541,N_3273,N_1368);
xor U10542 (N_10542,N_5325,N_4310);
xnor U10543 (N_10543,N_562,N_836);
xnor U10544 (N_10544,N_640,N_5714);
nand U10545 (N_10545,N_4099,N_207);
nor U10546 (N_10546,N_4547,N_2137);
nor U10547 (N_10547,N_3314,N_1148);
nor U10548 (N_10548,N_2888,N_2716);
or U10549 (N_10549,N_291,N_548);
and U10550 (N_10550,N_2840,N_4972);
or U10551 (N_10551,N_4026,N_4893);
or U10552 (N_10552,N_5909,N_194);
nand U10553 (N_10553,N_1826,N_3186);
and U10554 (N_10554,N_4596,N_5357);
nand U10555 (N_10555,N_2697,N_6000);
or U10556 (N_10556,N_4816,N_1187);
and U10557 (N_10557,N_3429,N_3448);
nor U10558 (N_10558,N_3531,N_4444);
and U10559 (N_10559,N_5371,N_1250);
nand U10560 (N_10560,N_2605,N_2632);
or U10561 (N_10561,N_5219,N_4419);
nand U10562 (N_10562,N_293,N_5383);
and U10563 (N_10563,N_5540,N_4609);
or U10564 (N_10564,N_2013,N_25);
and U10565 (N_10565,N_3074,N_5441);
and U10566 (N_10566,N_406,N_2632);
xnor U10567 (N_10567,N_4256,N_4128);
xor U10568 (N_10568,N_4001,N_804);
nand U10569 (N_10569,N_350,N_104);
nand U10570 (N_10570,N_946,N_4450);
and U10571 (N_10571,N_360,N_5422);
nand U10572 (N_10572,N_3720,N_3056);
nor U10573 (N_10573,N_6187,N_4216);
nand U10574 (N_10574,N_2193,N_757);
nor U10575 (N_10575,N_4792,N_6161);
and U10576 (N_10576,N_4433,N_2643);
nand U10577 (N_10577,N_1213,N_4859);
and U10578 (N_10578,N_2604,N_2222);
nand U10579 (N_10579,N_4968,N_5586);
and U10580 (N_10580,N_3173,N_1230);
and U10581 (N_10581,N_1348,N_21);
nor U10582 (N_10582,N_3001,N_217);
or U10583 (N_10583,N_6030,N_226);
nand U10584 (N_10584,N_3147,N_1767);
and U10585 (N_10585,N_539,N_4685);
and U10586 (N_10586,N_2954,N_4337);
nor U10587 (N_10587,N_4727,N_561);
nor U10588 (N_10588,N_1591,N_3752);
xor U10589 (N_10589,N_4521,N_2973);
nor U10590 (N_10590,N_3115,N_5322);
and U10591 (N_10591,N_3657,N_3490);
xor U10592 (N_10592,N_4311,N_995);
nor U10593 (N_10593,N_4413,N_3685);
nand U10594 (N_10594,N_2543,N_4914);
nand U10595 (N_10595,N_2902,N_6235);
or U10596 (N_10596,N_5125,N_3813);
or U10597 (N_10597,N_4449,N_3866);
nand U10598 (N_10598,N_4546,N_4802);
xnor U10599 (N_10599,N_203,N_3584);
nand U10600 (N_10600,N_4221,N_4053);
nand U10601 (N_10601,N_1461,N_3759);
nor U10602 (N_10602,N_1077,N_4096);
nand U10603 (N_10603,N_938,N_4137);
nor U10604 (N_10604,N_4682,N_463);
nor U10605 (N_10605,N_3008,N_5796);
xnor U10606 (N_10606,N_4536,N_3573);
nor U10607 (N_10607,N_3014,N_5602);
and U10608 (N_10608,N_3043,N_321);
nor U10609 (N_10609,N_3266,N_5521);
and U10610 (N_10610,N_1727,N_2083);
or U10611 (N_10611,N_2754,N_897);
nand U10612 (N_10612,N_719,N_1257);
nor U10613 (N_10613,N_1173,N_3972);
nand U10614 (N_10614,N_6116,N_1509);
or U10615 (N_10615,N_5662,N_5763);
and U10616 (N_10616,N_3705,N_3001);
xnor U10617 (N_10617,N_3899,N_5734);
xor U10618 (N_10618,N_640,N_5098);
xor U10619 (N_10619,N_2417,N_1119);
xor U10620 (N_10620,N_6131,N_4933);
nand U10621 (N_10621,N_5159,N_6162);
nor U10622 (N_10622,N_3116,N_4469);
nor U10623 (N_10623,N_346,N_4864);
or U10624 (N_10624,N_5134,N_3558);
and U10625 (N_10625,N_3214,N_3659);
or U10626 (N_10626,N_2293,N_3810);
nand U10627 (N_10627,N_1016,N_2901);
or U10628 (N_10628,N_4221,N_1336);
xor U10629 (N_10629,N_2669,N_1226);
nor U10630 (N_10630,N_3169,N_3716);
nand U10631 (N_10631,N_5447,N_5547);
xor U10632 (N_10632,N_4249,N_425);
nor U10633 (N_10633,N_3747,N_4012);
and U10634 (N_10634,N_934,N_1963);
nand U10635 (N_10635,N_5076,N_5826);
nand U10636 (N_10636,N_1446,N_6105);
xor U10637 (N_10637,N_134,N_5305);
xor U10638 (N_10638,N_4014,N_3514);
nand U10639 (N_10639,N_3767,N_2141);
and U10640 (N_10640,N_5729,N_4060);
nand U10641 (N_10641,N_2019,N_1433);
xnor U10642 (N_10642,N_426,N_3062);
and U10643 (N_10643,N_2688,N_3256);
nand U10644 (N_10644,N_2744,N_4252);
nor U10645 (N_10645,N_2645,N_5819);
xor U10646 (N_10646,N_2178,N_808);
xnor U10647 (N_10647,N_3079,N_5690);
nor U10648 (N_10648,N_1523,N_5262);
or U10649 (N_10649,N_1293,N_5661);
and U10650 (N_10650,N_1743,N_4840);
xnor U10651 (N_10651,N_4969,N_270);
nand U10652 (N_10652,N_2875,N_2235);
nand U10653 (N_10653,N_3025,N_2361);
nor U10654 (N_10654,N_3879,N_2341);
xnor U10655 (N_10655,N_356,N_2169);
nor U10656 (N_10656,N_2014,N_1134);
nand U10657 (N_10657,N_8,N_3586);
xnor U10658 (N_10658,N_1703,N_3800);
nand U10659 (N_10659,N_5407,N_2192);
nor U10660 (N_10660,N_4452,N_2098);
xor U10661 (N_10661,N_2563,N_2938);
and U10662 (N_10662,N_337,N_5193);
nor U10663 (N_10663,N_853,N_2640);
xnor U10664 (N_10664,N_975,N_3550);
xnor U10665 (N_10665,N_2728,N_511);
or U10666 (N_10666,N_2601,N_4068);
nand U10667 (N_10667,N_2393,N_788);
and U10668 (N_10668,N_6027,N_2277);
xor U10669 (N_10669,N_2552,N_3297);
and U10670 (N_10670,N_907,N_4204);
nor U10671 (N_10671,N_2179,N_6207);
and U10672 (N_10672,N_1937,N_5135);
and U10673 (N_10673,N_2799,N_4765);
and U10674 (N_10674,N_81,N_658);
and U10675 (N_10675,N_576,N_6111);
or U10676 (N_10676,N_1800,N_5327);
xnor U10677 (N_10677,N_1854,N_3967);
or U10678 (N_10678,N_702,N_2915);
or U10679 (N_10679,N_3557,N_2523);
nand U10680 (N_10680,N_5726,N_5611);
and U10681 (N_10681,N_1070,N_222);
nor U10682 (N_10682,N_393,N_5066);
xor U10683 (N_10683,N_5823,N_5521);
or U10684 (N_10684,N_2520,N_3428);
nand U10685 (N_10685,N_2300,N_5153);
nor U10686 (N_10686,N_4491,N_6165);
and U10687 (N_10687,N_3544,N_116);
and U10688 (N_10688,N_4602,N_6090);
nor U10689 (N_10689,N_1324,N_3123);
or U10690 (N_10690,N_3334,N_1826);
nor U10691 (N_10691,N_3049,N_2758);
and U10692 (N_10692,N_5167,N_2563);
or U10693 (N_10693,N_5389,N_3924);
and U10694 (N_10694,N_4191,N_1327);
xor U10695 (N_10695,N_5044,N_3642);
nor U10696 (N_10696,N_5998,N_3236);
or U10697 (N_10697,N_4620,N_896);
nor U10698 (N_10698,N_1302,N_3286);
nand U10699 (N_10699,N_3190,N_69);
or U10700 (N_10700,N_4766,N_1832);
nand U10701 (N_10701,N_1739,N_5204);
xnor U10702 (N_10702,N_3256,N_2045);
or U10703 (N_10703,N_5123,N_1230);
nor U10704 (N_10704,N_5458,N_2213);
or U10705 (N_10705,N_6106,N_5115);
xnor U10706 (N_10706,N_4195,N_5852);
or U10707 (N_10707,N_5295,N_4437);
nor U10708 (N_10708,N_579,N_2251);
xor U10709 (N_10709,N_381,N_4674);
nor U10710 (N_10710,N_2397,N_328);
nand U10711 (N_10711,N_1886,N_354);
nand U10712 (N_10712,N_2531,N_907);
xor U10713 (N_10713,N_3217,N_3858);
nor U10714 (N_10714,N_3469,N_535);
nor U10715 (N_10715,N_162,N_3441);
and U10716 (N_10716,N_1756,N_155);
nor U10717 (N_10717,N_25,N_3921);
and U10718 (N_10718,N_4339,N_3942);
nor U10719 (N_10719,N_125,N_2858);
or U10720 (N_10720,N_4789,N_4237);
nand U10721 (N_10721,N_4299,N_2484);
or U10722 (N_10722,N_5464,N_654);
xnor U10723 (N_10723,N_2424,N_1765);
nand U10724 (N_10724,N_4782,N_1165);
xor U10725 (N_10725,N_425,N_2616);
nor U10726 (N_10726,N_4207,N_3481);
and U10727 (N_10727,N_1733,N_1479);
and U10728 (N_10728,N_624,N_4211);
nor U10729 (N_10729,N_1960,N_1809);
xnor U10730 (N_10730,N_2231,N_4143);
and U10731 (N_10731,N_2140,N_4183);
or U10732 (N_10732,N_2157,N_2819);
or U10733 (N_10733,N_5553,N_2897);
nor U10734 (N_10734,N_3683,N_229);
nor U10735 (N_10735,N_374,N_884);
and U10736 (N_10736,N_2864,N_2348);
nor U10737 (N_10737,N_394,N_863);
or U10738 (N_10738,N_896,N_1127);
xor U10739 (N_10739,N_2395,N_3511);
nor U10740 (N_10740,N_79,N_4464);
nor U10741 (N_10741,N_4011,N_720);
and U10742 (N_10742,N_4380,N_1322);
nand U10743 (N_10743,N_2323,N_4667);
xnor U10744 (N_10744,N_5996,N_4440);
xnor U10745 (N_10745,N_2382,N_1231);
nand U10746 (N_10746,N_4449,N_3155);
and U10747 (N_10747,N_990,N_3685);
nand U10748 (N_10748,N_5781,N_3187);
and U10749 (N_10749,N_6187,N_3676);
nor U10750 (N_10750,N_5620,N_1706);
nand U10751 (N_10751,N_3893,N_650);
xnor U10752 (N_10752,N_657,N_4315);
xor U10753 (N_10753,N_2794,N_5967);
nor U10754 (N_10754,N_2332,N_5286);
and U10755 (N_10755,N_3248,N_331);
or U10756 (N_10756,N_3690,N_2191);
nor U10757 (N_10757,N_884,N_4613);
and U10758 (N_10758,N_3502,N_5688);
or U10759 (N_10759,N_5682,N_4986);
nand U10760 (N_10760,N_3930,N_183);
nor U10761 (N_10761,N_3952,N_3694);
nor U10762 (N_10762,N_3127,N_1658);
or U10763 (N_10763,N_46,N_2194);
nor U10764 (N_10764,N_4758,N_2078);
or U10765 (N_10765,N_102,N_3594);
xnor U10766 (N_10766,N_2129,N_728);
and U10767 (N_10767,N_4520,N_3624);
nand U10768 (N_10768,N_2822,N_676);
or U10769 (N_10769,N_3006,N_741);
nor U10770 (N_10770,N_3289,N_1442);
nor U10771 (N_10771,N_3339,N_2955);
nor U10772 (N_10772,N_498,N_5004);
and U10773 (N_10773,N_266,N_746);
xnor U10774 (N_10774,N_2304,N_5571);
nor U10775 (N_10775,N_1783,N_3583);
and U10776 (N_10776,N_3355,N_3161);
or U10777 (N_10777,N_79,N_1642);
xor U10778 (N_10778,N_3440,N_4053);
and U10779 (N_10779,N_5486,N_4607);
nor U10780 (N_10780,N_4190,N_3767);
xnor U10781 (N_10781,N_2080,N_415);
nand U10782 (N_10782,N_1536,N_4203);
xor U10783 (N_10783,N_5866,N_2456);
nand U10784 (N_10784,N_1353,N_144);
nand U10785 (N_10785,N_3477,N_4503);
xnor U10786 (N_10786,N_5465,N_206);
nor U10787 (N_10787,N_522,N_1656);
nand U10788 (N_10788,N_4905,N_2355);
nor U10789 (N_10789,N_1928,N_13);
and U10790 (N_10790,N_995,N_1318);
or U10791 (N_10791,N_4383,N_939);
or U10792 (N_10792,N_474,N_4547);
nor U10793 (N_10793,N_4622,N_2181);
or U10794 (N_10794,N_2319,N_5213);
nand U10795 (N_10795,N_2216,N_6210);
or U10796 (N_10796,N_2717,N_3290);
and U10797 (N_10797,N_4153,N_4536);
or U10798 (N_10798,N_4840,N_1593);
or U10799 (N_10799,N_984,N_3060);
xnor U10800 (N_10800,N_5991,N_6176);
nand U10801 (N_10801,N_2118,N_429);
nor U10802 (N_10802,N_4391,N_2889);
nor U10803 (N_10803,N_4456,N_1002);
and U10804 (N_10804,N_4174,N_5507);
xnor U10805 (N_10805,N_5201,N_5260);
and U10806 (N_10806,N_3136,N_860);
nor U10807 (N_10807,N_2954,N_4554);
nor U10808 (N_10808,N_3645,N_4178);
or U10809 (N_10809,N_2947,N_4385);
xnor U10810 (N_10810,N_87,N_2547);
and U10811 (N_10811,N_3179,N_419);
or U10812 (N_10812,N_1695,N_5669);
nor U10813 (N_10813,N_823,N_668);
xor U10814 (N_10814,N_2811,N_1350);
nor U10815 (N_10815,N_711,N_5705);
or U10816 (N_10816,N_462,N_4263);
and U10817 (N_10817,N_824,N_693);
and U10818 (N_10818,N_5567,N_871);
xnor U10819 (N_10819,N_4848,N_5796);
nand U10820 (N_10820,N_4772,N_1668);
or U10821 (N_10821,N_1957,N_3993);
nor U10822 (N_10822,N_3571,N_4651);
xnor U10823 (N_10823,N_902,N_2233);
or U10824 (N_10824,N_4983,N_3023);
nor U10825 (N_10825,N_4809,N_3939);
or U10826 (N_10826,N_4832,N_653);
nor U10827 (N_10827,N_2626,N_3652);
nor U10828 (N_10828,N_3337,N_1786);
xnor U10829 (N_10829,N_1713,N_4033);
and U10830 (N_10830,N_4324,N_2010);
xnor U10831 (N_10831,N_5068,N_4422);
or U10832 (N_10832,N_2011,N_2101);
and U10833 (N_10833,N_4973,N_928);
nand U10834 (N_10834,N_4959,N_4311);
xor U10835 (N_10835,N_5803,N_6012);
xnor U10836 (N_10836,N_2574,N_2624);
nand U10837 (N_10837,N_5322,N_3474);
nand U10838 (N_10838,N_6132,N_3086);
or U10839 (N_10839,N_1684,N_1568);
nor U10840 (N_10840,N_5157,N_3140);
xor U10841 (N_10841,N_4649,N_1615);
xnor U10842 (N_10842,N_2993,N_4930);
xnor U10843 (N_10843,N_1848,N_3928);
nand U10844 (N_10844,N_187,N_636);
nor U10845 (N_10845,N_4157,N_5897);
and U10846 (N_10846,N_5169,N_5976);
or U10847 (N_10847,N_730,N_1300);
or U10848 (N_10848,N_3466,N_5880);
nor U10849 (N_10849,N_4910,N_1451);
nand U10850 (N_10850,N_1538,N_1063);
nand U10851 (N_10851,N_5955,N_2603);
and U10852 (N_10852,N_1687,N_4412);
and U10853 (N_10853,N_2830,N_1104);
xor U10854 (N_10854,N_3110,N_2428);
or U10855 (N_10855,N_6141,N_4126);
and U10856 (N_10856,N_5846,N_2980);
xnor U10857 (N_10857,N_4030,N_338);
and U10858 (N_10858,N_6141,N_1184);
and U10859 (N_10859,N_259,N_5014);
nor U10860 (N_10860,N_4886,N_4336);
and U10861 (N_10861,N_4916,N_2357);
xnor U10862 (N_10862,N_2711,N_6067);
nor U10863 (N_10863,N_73,N_1689);
and U10864 (N_10864,N_4115,N_5160);
or U10865 (N_10865,N_5050,N_1191);
or U10866 (N_10866,N_227,N_2446);
nand U10867 (N_10867,N_2981,N_3960);
or U10868 (N_10868,N_3573,N_1991);
nand U10869 (N_10869,N_5329,N_2110);
xnor U10870 (N_10870,N_4281,N_2703);
and U10871 (N_10871,N_3517,N_4677);
and U10872 (N_10872,N_5229,N_2889);
or U10873 (N_10873,N_5532,N_787);
and U10874 (N_10874,N_3754,N_3632);
nor U10875 (N_10875,N_1150,N_2402);
and U10876 (N_10876,N_1227,N_1596);
xnor U10877 (N_10877,N_4715,N_5083);
nor U10878 (N_10878,N_2101,N_3466);
and U10879 (N_10879,N_2493,N_3222);
nor U10880 (N_10880,N_549,N_5215);
nand U10881 (N_10881,N_3601,N_2567);
or U10882 (N_10882,N_1286,N_4808);
and U10883 (N_10883,N_5415,N_4684);
and U10884 (N_10884,N_4495,N_2529);
or U10885 (N_10885,N_5312,N_4397);
xnor U10886 (N_10886,N_5079,N_1412);
nand U10887 (N_10887,N_2468,N_5185);
nand U10888 (N_10888,N_1208,N_2386);
xor U10889 (N_10889,N_625,N_494);
and U10890 (N_10890,N_3023,N_5285);
nand U10891 (N_10891,N_2763,N_4036);
xor U10892 (N_10892,N_2733,N_4118);
and U10893 (N_10893,N_2738,N_5769);
nand U10894 (N_10894,N_5355,N_1705);
or U10895 (N_10895,N_548,N_76);
and U10896 (N_10896,N_5261,N_3981);
nor U10897 (N_10897,N_3775,N_4017);
nand U10898 (N_10898,N_3143,N_6189);
xor U10899 (N_10899,N_2241,N_2731);
and U10900 (N_10900,N_3461,N_2292);
and U10901 (N_10901,N_6117,N_2804);
xor U10902 (N_10902,N_2113,N_2660);
or U10903 (N_10903,N_5744,N_4293);
nor U10904 (N_10904,N_908,N_1846);
and U10905 (N_10905,N_3666,N_6029);
nand U10906 (N_10906,N_5251,N_5201);
and U10907 (N_10907,N_5558,N_305);
nand U10908 (N_10908,N_5040,N_389);
xor U10909 (N_10909,N_5080,N_5825);
nor U10910 (N_10910,N_1337,N_5040);
and U10911 (N_10911,N_4716,N_5768);
and U10912 (N_10912,N_2083,N_3990);
xor U10913 (N_10913,N_2491,N_942);
nor U10914 (N_10914,N_2525,N_2828);
nand U10915 (N_10915,N_1966,N_5855);
xnor U10916 (N_10916,N_4636,N_3839);
nand U10917 (N_10917,N_5448,N_5980);
nand U10918 (N_10918,N_5823,N_5736);
xnor U10919 (N_10919,N_2189,N_5636);
nand U10920 (N_10920,N_3800,N_6004);
or U10921 (N_10921,N_3746,N_4200);
xor U10922 (N_10922,N_2640,N_6168);
xor U10923 (N_10923,N_5618,N_5638);
nand U10924 (N_10924,N_3572,N_290);
nor U10925 (N_10925,N_2621,N_2145);
nand U10926 (N_10926,N_1807,N_6096);
and U10927 (N_10927,N_1643,N_4450);
and U10928 (N_10928,N_3866,N_1973);
or U10929 (N_10929,N_6234,N_2181);
and U10930 (N_10930,N_598,N_2243);
nor U10931 (N_10931,N_664,N_4302);
or U10932 (N_10932,N_3470,N_1683);
nor U10933 (N_10933,N_3091,N_3659);
nor U10934 (N_10934,N_1458,N_5739);
xor U10935 (N_10935,N_6030,N_2894);
nand U10936 (N_10936,N_1129,N_1935);
nor U10937 (N_10937,N_846,N_3333);
nand U10938 (N_10938,N_1045,N_2464);
xnor U10939 (N_10939,N_1344,N_5259);
or U10940 (N_10940,N_4700,N_2732);
nand U10941 (N_10941,N_1011,N_1196);
nor U10942 (N_10942,N_3981,N_6227);
and U10943 (N_10943,N_556,N_2117);
nand U10944 (N_10944,N_2504,N_6034);
or U10945 (N_10945,N_1105,N_4979);
xnor U10946 (N_10946,N_2532,N_5108);
nand U10947 (N_10947,N_582,N_2352);
nor U10948 (N_10948,N_5230,N_5022);
nor U10949 (N_10949,N_2140,N_4832);
and U10950 (N_10950,N_1010,N_4639);
nor U10951 (N_10951,N_3923,N_4225);
and U10952 (N_10952,N_5094,N_2242);
nor U10953 (N_10953,N_4367,N_4914);
nand U10954 (N_10954,N_3304,N_5798);
nand U10955 (N_10955,N_4497,N_2346);
or U10956 (N_10956,N_5575,N_1936);
xor U10957 (N_10957,N_1647,N_1984);
xor U10958 (N_10958,N_1060,N_5076);
xnor U10959 (N_10959,N_2352,N_1707);
or U10960 (N_10960,N_3961,N_5127);
or U10961 (N_10961,N_4034,N_5525);
or U10962 (N_10962,N_4457,N_5220);
nand U10963 (N_10963,N_988,N_1656);
xor U10964 (N_10964,N_1189,N_546);
xor U10965 (N_10965,N_2033,N_3308);
and U10966 (N_10966,N_579,N_2736);
and U10967 (N_10967,N_2510,N_3509);
nor U10968 (N_10968,N_2741,N_2169);
xor U10969 (N_10969,N_4975,N_5509);
and U10970 (N_10970,N_4847,N_2185);
or U10971 (N_10971,N_2654,N_751);
xor U10972 (N_10972,N_5791,N_5914);
nand U10973 (N_10973,N_1470,N_5005);
xor U10974 (N_10974,N_496,N_5893);
nand U10975 (N_10975,N_4440,N_1368);
or U10976 (N_10976,N_5242,N_1654);
nor U10977 (N_10977,N_4590,N_1183);
and U10978 (N_10978,N_4864,N_4779);
xnor U10979 (N_10979,N_5220,N_1051);
nor U10980 (N_10980,N_2240,N_2963);
nand U10981 (N_10981,N_1931,N_978);
or U10982 (N_10982,N_884,N_2997);
xor U10983 (N_10983,N_5402,N_5970);
xor U10984 (N_10984,N_3269,N_6173);
xnor U10985 (N_10985,N_2851,N_6071);
nand U10986 (N_10986,N_466,N_2637);
nor U10987 (N_10987,N_3064,N_2419);
xnor U10988 (N_10988,N_4874,N_85);
nor U10989 (N_10989,N_2548,N_5821);
or U10990 (N_10990,N_4060,N_4622);
xnor U10991 (N_10991,N_1715,N_889);
or U10992 (N_10992,N_5963,N_5525);
xor U10993 (N_10993,N_4266,N_940);
xnor U10994 (N_10994,N_6031,N_199);
and U10995 (N_10995,N_4398,N_6064);
nor U10996 (N_10996,N_1121,N_1391);
and U10997 (N_10997,N_3410,N_1867);
or U10998 (N_10998,N_2697,N_3602);
nor U10999 (N_10999,N_1702,N_2593);
nor U11000 (N_11000,N_5510,N_2487);
and U11001 (N_11001,N_2098,N_1068);
nand U11002 (N_11002,N_3927,N_1160);
and U11003 (N_11003,N_1521,N_994);
or U11004 (N_11004,N_6247,N_2567);
xnor U11005 (N_11005,N_461,N_5519);
and U11006 (N_11006,N_3324,N_3684);
nand U11007 (N_11007,N_4179,N_3082);
or U11008 (N_11008,N_130,N_350);
and U11009 (N_11009,N_2872,N_3139);
and U11010 (N_11010,N_2068,N_1453);
and U11011 (N_11011,N_2765,N_5855);
xor U11012 (N_11012,N_5796,N_3749);
nor U11013 (N_11013,N_2788,N_1114);
nor U11014 (N_11014,N_2818,N_5284);
nor U11015 (N_11015,N_3502,N_4861);
or U11016 (N_11016,N_873,N_4268);
xor U11017 (N_11017,N_4583,N_5685);
or U11018 (N_11018,N_2230,N_1256);
or U11019 (N_11019,N_6219,N_1367);
and U11020 (N_11020,N_1999,N_1800);
xor U11021 (N_11021,N_2224,N_85);
or U11022 (N_11022,N_6168,N_220);
nor U11023 (N_11023,N_870,N_6150);
or U11024 (N_11024,N_4805,N_5472);
nor U11025 (N_11025,N_1756,N_4876);
or U11026 (N_11026,N_275,N_4841);
xnor U11027 (N_11027,N_5734,N_1001);
nor U11028 (N_11028,N_3114,N_2457);
nor U11029 (N_11029,N_146,N_1252);
xnor U11030 (N_11030,N_437,N_939);
xnor U11031 (N_11031,N_4471,N_2837);
nor U11032 (N_11032,N_2658,N_1302);
nor U11033 (N_11033,N_2058,N_807);
or U11034 (N_11034,N_16,N_6228);
or U11035 (N_11035,N_5880,N_337);
xnor U11036 (N_11036,N_76,N_4066);
xnor U11037 (N_11037,N_5394,N_2857);
nor U11038 (N_11038,N_4403,N_6232);
and U11039 (N_11039,N_1215,N_2622);
nor U11040 (N_11040,N_5101,N_4802);
and U11041 (N_11041,N_4458,N_4394);
nand U11042 (N_11042,N_3783,N_5227);
nor U11043 (N_11043,N_5750,N_5562);
xor U11044 (N_11044,N_3771,N_1951);
nor U11045 (N_11045,N_5409,N_3630);
nor U11046 (N_11046,N_2689,N_3787);
nor U11047 (N_11047,N_4147,N_1353);
nand U11048 (N_11048,N_1274,N_5343);
or U11049 (N_11049,N_5208,N_1993);
or U11050 (N_11050,N_1159,N_2467);
and U11051 (N_11051,N_3840,N_531);
or U11052 (N_11052,N_1421,N_5892);
xnor U11053 (N_11053,N_141,N_1767);
and U11054 (N_11054,N_2078,N_5982);
nand U11055 (N_11055,N_5630,N_5290);
nand U11056 (N_11056,N_2622,N_4114);
or U11057 (N_11057,N_4142,N_4837);
nor U11058 (N_11058,N_6016,N_2838);
or U11059 (N_11059,N_3438,N_2112);
xnor U11060 (N_11060,N_3925,N_6003);
or U11061 (N_11061,N_3417,N_2742);
nor U11062 (N_11062,N_2485,N_3970);
or U11063 (N_11063,N_5021,N_2395);
nor U11064 (N_11064,N_6187,N_5161);
xnor U11065 (N_11065,N_17,N_2550);
xnor U11066 (N_11066,N_2196,N_655);
or U11067 (N_11067,N_5847,N_5254);
nor U11068 (N_11068,N_2448,N_4455);
nand U11069 (N_11069,N_3687,N_97);
or U11070 (N_11070,N_6078,N_6049);
nor U11071 (N_11071,N_3393,N_5394);
or U11072 (N_11072,N_643,N_5117);
and U11073 (N_11073,N_3553,N_628);
or U11074 (N_11074,N_3850,N_281);
nand U11075 (N_11075,N_3994,N_2740);
nor U11076 (N_11076,N_5817,N_4604);
or U11077 (N_11077,N_1634,N_3257);
or U11078 (N_11078,N_4795,N_2904);
or U11079 (N_11079,N_428,N_4153);
xnor U11080 (N_11080,N_2739,N_1021);
nor U11081 (N_11081,N_1926,N_1737);
and U11082 (N_11082,N_5823,N_94);
nor U11083 (N_11083,N_2446,N_5318);
and U11084 (N_11084,N_1226,N_2544);
nor U11085 (N_11085,N_2105,N_3429);
nor U11086 (N_11086,N_5519,N_858);
and U11087 (N_11087,N_4060,N_3222);
and U11088 (N_11088,N_1442,N_535);
nand U11089 (N_11089,N_3461,N_232);
nor U11090 (N_11090,N_4445,N_2955);
and U11091 (N_11091,N_3995,N_2276);
and U11092 (N_11092,N_2587,N_1947);
or U11093 (N_11093,N_6228,N_5594);
xnor U11094 (N_11094,N_495,N_5758);
or U11095 (N_11095,N_2009,N_2632);
or U11096 (N_11096,N_6032,N_4366);
or U11097 (N_11097,N_3388,N_1762);
and U11098 (N_11098,N_1017,N_5357);
nor U11099 (N_11099,N_5877,N_1139);
or U11100 (N_11100,N_2215,N_1371);
xnor U11101 (N_11101,N_6143,N_140);
xor U11102 (N_11102,N_3033,N_273);
and U11103 (N_11103,N_4332,N_1932);
xnor U11104 (N_11104,N_5360,N_3667);
and U11105 (N_11105,N_1612,N_4820);
nand U11106 (N_11106,N_414,N_4596);
nor U11107 (N_11107,N_1868,N_4279);
or U11108 (N_11108,N_874,N_5981);
xnor U11109 (N_11109,N_5941,N_857);
nor U11110 (N_11110,N_657,N_5256);
nor U11111 (N_11111,N_656,N_1341);
or U11112 (N_11112,N_3007,N_5942);
or U11113 (N_11113,N_4748,N_4477);
or U11114 (N_11114,N_5978,N_2595);
and U11115 (N_11115,N_2181,N_5713);
nand U11116 (N_11116,N_2247,N_1925);
nand U11117 (N_11117,N_1823,N_3901);
xor U11118 (N_11118,N_3639,N_478);
xnor U11119 (N_11119,N_1236,N_5851);
nor U11120 (N_11120,N_1773,N_4233);
nand U11121 (N_11121,N_6188,N_1742);
xnor U11122 (N_11122,N_4812,N_4977);
and U11123 (N_11123,N_3158,N_6047);
or U11124 (N_11124,N_289,N_3019);
nor U11125 (N_11125,N_371,N_249);
or U11126 (N_11126,N_4102,N_1090);
and U11127 (N_11127,N_6197,N_2816);
nor U11128 (N_11128,N_3776,N_5347);
or U11129 (N_11129,N_4203,N_2604);
and U11130 (N_11130,N_4866,N_3734);
xor U11131 (N_11131,N_613,N_5526);
or U11132 (N_11132,N_3378,N_2845);
or U11133 (N_11133,N_5576,N_5603);
xnor U11134 (N_11134,N_5844,N_3889);
and U11135 (N_11135,N_2644,N_438);
and U11136 (N_11136,N_2553,N_4380);
nor U11137 (N_11137,N_2377,N_629);
nand U11138 (N_11138,N_2139,N_6182);
xor U11139 (N_11139,N_2983,N_5971);
nand U11140 (N_11140,N_3721,N_5522);
xor U11141 (N_11141,N_5588,N_962);
or U11142 (N_11142,N_3100,N_4670);
nand U11143 (N_11143,N_30,N_4992);
or U11144 (N_11144,N_3815,N_6176);
xnor U11145 (N_11145,N_4977,N_2570);
nand U11146 (N_11146,N_4365,N_6187);
and U11147 (N_11147,N_1866,N_356);
nand U11148 (N_11148,N_1112,N_2499);
nand U11149 (N_11149,N_635,N_5814);
nand U11150 (N_11150,N_223,N_2130);
nor U11151 (N_11151,N_2799,N_4944);
nor U11152 (N_11152,N_5181,N_5799);
nand U11153 (N_11153,N_3821,N_2574);
and U11154 (N_11154,N_5264,N_2453);
nand U11155 (N_11155,N_6060,N_2786);
xnor U11156 (N_11156,N_2062,N_465);
nand U11157 (N_11157,N_555,N_2990);
or U11158 (N_11158,N_4571,N_2079);
xnor U11159 (N_11159,N_5476,N_5964);
nand U11160 (N_11160,N_4919,N_5571);
or U11161 (N_11161,N_4967,N_6039);
xnor U11162 (N_11162,N_3438,N_5630);
nand U11163 (N_11163,N_3761,N_1092);
xnor U11164 (N_11164,N_4855,N_3505);
nand U11165 (N_11165,N_5005,N_5992);
nand U11166 (N_11166,N_5118,N_5816);
or U11167 (N_11167,N_934,N_4654);
nand U11168 (N_11168,N_1176,N_2515);
nand U11169 (N_11169,N_1391,N_1734);
or U11170 (N_11170,N_5186,N_3272);
or U11171 (N_11171,N_3986,N_941);
xnor U11172 (N_11172,N_838,N_3886);
nor U11173 (N_11173,N_4221,N_1813);
and U11174 (N_11174,N_6156,N_245);
nor U11175 (N_11175,N_2152,N_4763);
and U11176 (N_11176,N_5040,N_1141);
xor U11177 (N_11177,N_2939,N_3401);
and U11178 (N_11178,N_4981,N_3613);
xnor U11179 (N_11179,N_2807,N_2383);
or U11180 (N_11180,N_4552,N_6097);
xnor U11181 (N_11181,N_859,N_5319);
nand U11182 (N_11182,N_67,N_3069);
or U11183 (N_11183,N_27,N_5397);
nand U11184 (N_11184,N_6189,N_4803);
or U11185 (N_11185,N_1792,N_2235);
nor U11186 (N_11186,N_4617,N_4269);
xor U11187 (N_11187,N_152,N_5489);
and U11188 (N_11188,N_2941,N_2523);
and U11189 (N_11189,N_2145,N_5356);
nand U11190 (N_11190,N_5536,N_3722);
nand U11191 (N_11191,N_3612,N_1257);
and U11192 (N_11192,N_378,N_2805);
nand U11193 (N_11193,N_167,N_3841);
and U11194 (N_11194,N_2136,N_3252);
xor U11195 (N_11195,N_2386,N_1498);
nor U11196 (N_11196,N_3367,N_3282);
nand U11197 (N_11197,N_297,N_3416);
nor U11198 (N_11198,N_678,N_3340);
nor U11199 (N_11199,N_2091,N_4780);
xor U11200 (N_11200,N_3969,N_1684);
and U11201 (N_11201,N_5328,N_5677);
xnor U11202 (N_11202,N_4082,N_3236);
xnor U11203 (N_11203,N_3121,N_5693);
and U11204 (N_11204,N_5656,N_1570);
and U11205 (N_11205,N_4043,N_2544);
xnor U11206 (N_11206,N_5568,N_4116);
xor U11207 (N_11207,N_2971,N_2476);
nand U11208 (N_11208,N_1391,N_796);
nor U11209 (N_11209,N_1069,N_3939);
xor U11210 (N_11210,N_3177,N_4975);
nor U11211 (N_11211,N_2474,N_3896);
or U11212 (N_11212,N_1763,N_3743);
nand U11213 (N_11213,N_1977,N_1069);
and U11214 (N_11214,N_2578,N_2115);
and U11215 (N_11215,N_2583,N_2683);
nor U11216 (N_11216,N_3842,N_3094);
or U11217 (N_11217,N_4948,N_142);
xnor U11218 (N_11218,N_5326,N_776);
nand U11219 (N_11219,N_3799,N_1162);
nand U11220 (N_11220,N_2910,N_2352);
xnor U11221 (N_11221,N_2278,N_3959);
xor U11222 (N_11222,N_3110,N_4640);
nand U11223 (N_11223,N_5576,N_2785);
or U11224 (N_11224,N_2021,N_2810);
nand U11225 (N_11225,N_3743,N_3865);
nand U11226 (N_11226,N_6054,N_5809);
nor U11227 (N_11227,N_1871,N_67);
or U11228 (N_11228,N_5548,N_6072);
or U11229 (N_11229,N_2644,N_3375);
xnor U11230 (N_11230,N_1234,N_4512);
nand U11231 (N_11231,N_2559,N_1781);
xor U11232 (N_11232,N_1353,N_5981);
xor U11233 (N_11233,N_4405,N_1109);
and U11234 (N_11234,N_1085,N_3769);
nor U11235 (N_11235,N_4644,N_5571);
and U11236 (N_11236,N_1077,N_4425);
nor U11237 (N_11237,N_2692,N_2316);
nand U11238 (N_11238,N_1854,N_298);
xor U11239 (N_11239,N_911,N_5466);
xor U11240 (N_11240,N_2793,N_1385);
nor U11241 (N_11241,N_5844,N_2033);
xor U11242 (N_11242,N_3267,N_4433);
nand U11243 (N_11243,N_5967,N_563);
xor U11244 (N_11244,N_5342,N_5473);
and U11245 (N_11245,N_616,N_4945);
nand U11246 (N_11246,N_4452,N_3126);
xnor U11247 (N_11247,N_2240,N_1993);
nand U11248 (N_11248,N_3156,N_1540);
xnor U11249 (N_11249,N_3739,N_1214);
nor U11250 (N_11250,N_1207,N_4417);
and U11251 (N_11251,N_2542,N_1319);
nor U11252 (N_11252,N_297,N_6034);
or U11253 (N_11253,N_1025,N_1083);
xor U11254 (N_11254,N_2938,N_1774);
nand U11255 (N_11255,N_962,N_5289);
or U11256 (N_11256,N_3450,N_4819);
xor U11257 (N_11257,N_5318,N_5188);
and U11258 (N_11258,N_834,N_5924);
or U11259 (N_11259,N_3916,N_1390);
nand U11260 (N_11260,N_4890,N_519);
and U11261 (N_11261,N_4992,N_241);
and U11262 (N_11262,N_3385,N_1355);
xor U11263 (N_11263,N_3537,N_4182);
xor U11264 (N_11264,N_4192,N_1681);
nor U11265 (N_11265,N_5590,N_4338);
or U11266 (N_11266,N_2276,N_2459);
or U11267 (N_11267,N_1471,N_5690);
nand U11268 (N_11268,N_1924,N_1912);
nand U11269 (N_11269,N_5222,N_1297);
and U11270 (N_11270,N_221,N_729);
and U11271 (N_11271,N_6148,N_222);
nor U11272 (N_11272,N_4464,N_1420);
and U11273 (N_11273,N_830,N_6149);
nor U11274 (N_11274,N_4875,N_2728);
or U11275 (N_11275,N_1285,N_3581);
and U11276 (N_11276,N_1509,N_5230);
nand U11277 (N_11277,N_2221,N_5012);
xor U11278 (N_11278,N_3701,N_5545);
xor U11279 (N_11279,N_363,N_2576);
xnor U11280 (N_11280,N_5212,N_4601);
or U11281 (N_11281,N_643,N_4033);
xor U11282 (N_11282,N_4864,N_4434);
or U11283 (N_11283,N_4118,N_2751);
or U11284 (N_11284,N_5066,N_2849);
xnor U11285 (N_11285,N_4680,N_3385);
xor U11286 (N_11286,N_2382,N_1161);
xor U11287 (N_11287,N_236,N_5857);
xnor U11288 (N_11288,N_695,N_3165);
nor U11289 (N_11289,N_4062,N_2681);
xnor U11290 (N_11290,N_4015,N_1188);
and U11291 (N_11291,N_4577,N_185);
xnor U11292 (N_11292,N_5532,N_3521);
nand U11293 (N_11293,N_6104,N_5713);
nand U11294 (N_11294,N_4690,N_1335);
nand U11295 (N_11295,N_5224,N_3047);
nor U11296 (N_11296,N_5992,N_2444);
and U11297 (N_11297,N_1222,N_291);
nor U11298 (N_11298,N_5799,N_5619);
and U11299 (N_11299,N_2840,N_3318);
nor U11300 (N_11300,N_2704,N_1716);
nor U11301 (N_11301,N_2931,N_2734);
or U11302 (N_11302,N_3090,N_3206);
or U11303 (N_11303,N_1694,N_5141);
nor U11304 (N_11304,N_1611,N_6176);
or U11305 (N_11305,N_2071,N_717);
nor U11306 (N_11306,N_2908,N_2139);
nand U11307 (N_11307,N_4008,N_4766);
nor U11308 (N_11308,N_5288,N_2946);
xor U11309 (N_11309,N_4159,N_5026);
xnor U11310 (N_11310,N_2563,N_1649);
xor U11311 (N_11311,N_1448,N_316);
and U11312 (N_11312,N_1592,N_1227);
and U11313 (N_11313,N_2531,N_1632);
or U11314 (N_11314,N_867,N_5801);
nand U11315 (N_11315,N_4465,N_4195);
nor U11316 (N_11316,N_2560,N_6114);
and U11317 (N_11317,N_1456,N_1776);
nand U11318 (N_11318,N_2779,N_2108);
and U11319 (N_11319,N_3317,N_2636);
nand U11320 (N_11320,N_3543,N_163);
and U11321 (N_11321,N_1712,N_5792);
and U11322 (N_11322,N_2112,N_1079);
nand U11323 (N_11323,N_6185,N_3828);
xor U11324 (N_11324,N_623,N_5373);
or U11325 (N_11325,N_4153,N_1686);
nor U11326 (N_11326,N_683,N_1449);
nor U11327 (N_11327,N_37,N_2680);
nand U11328 (N_11328,N_2634,N_4550);
nor U11329 (N_11329,N_353,N_5001);
xnor U11330 (N_11330,N_2808,N_2268);
and U11331 (N_11331,N_2915,N_418);
or U11332 (N_11332,N_2290,N_3052);
or U11333 (N_11333,N_3323,N_4189);
and U11334 (N_11334,N_5664,N_2080);
and U11335 (N_11335,N_3089,N_6172);
nor U11336 (N_11336,N_2449,N_3586);
or U11337 (N_11337,N_4375,N_5803);
or U11338 (N_11338,N_1897,N_3711);
and U11339 (N_11339,N_4449,N_3497);
nor U11340 (N_11340,N_3363,N_2864);
nor U11341 (N_11341,N_3346,N_1300);
and U11342 (N_11342,N_5208,N_3387);
nor U11343 (N_11343,N_2235,N_3978);
nand U11344 (N_11344,N_766,N_5946);
or U11345 (N_11345,N_4485,N_1562);
and U11346 (N_11346,N_3773,N_4190);
and U11347 (N_11347,N_2229,N_2537);
xor U11348 (N_11348,N_993,N_3709);
nand U11349 (N_11349,N_5893,N_3911);
nand U11350 (N_11350,N_3279,N_2635);
and U11351 (N_11351,N_448,N_3210);
xor U11352 (N_11352,N_3898,N_3593);
xor U11353 (N_11353,N_3937,N_2967);
or U11354 (N_11354,N_2259,N_3746);
and U11355 (N_11355,N_1834,N_4996);
xnor U11356 (N_11356,N_4679,N_4967);
nand U11357 (N_11357,N_2228,N_2357);
nor U11358 (N_11358,N_337,N_900);
nor U11359 (N_11359,N_3830,N_71);
nand U11360 (N_11360,N_4278,N_2755);
and U11361 (N_11361,N_1052,N_5060);
or U11362 (N_11362,N_837,N_4633);
or U11363 (N_11363,N_4102,N_1844);
or U11364 (N_11364,N_2821,N_3378);
nor U11365 (N_11365,N_5973,N_4054);
xnor U11366 (N_11366,N_1577,N_160);
xor U11367 (N_11367,N_754,N_5307);
or U11368 (N_11368,N_2053,N_671);
and U11369 (N_11369,N_2960,N_1980);
or U11370 (N_11370,N_1050,N_4867);
nand U11371 (N_11371,N_4731,N_2816);
nand U11372 (N_11372,N_6201,N_488);
nand U11373 (N_11373,N_2785,N_4302);
xor U11374 (N_11374,N_3339,N_2932);
xor U11375 (N_11375,N_5509,N_3593);
nor U11376 (N_11376,N_3205,N_2186);
nand U11377 (N_11377,N_5068,N_1943);
nor U11378 (N_11378,N_1911,N_1270);
nor U11379 (N_11379,N_4397,N_699);
nand U11380 (N_11380,N_6088,N_1302);
or U11381 (N_11381,N_2061,N_1610);
xor U11382 (N_11382,N_330,N_5860);
and U11383 (N_11383,N_1369,N_2365);
or U11384 (N_11384,N_2034,N_3764);
or U11385 (N_11385,N_4917,N_274);
nor U11386 (N_11386,N_5959,N_1589);
xnor U11387 (N_11387,N_5463,N_1409);
or U11388 (N_11388,N_888,N_3698);
xnor U11389 (N_11389,N_2440,N_3062);
nor U11390 (N_11390,N_3826,N_1673);
nor U11391 (N_11391,N_93,N_3466);
and U11392 (N_11392,N_2522,N_402);
xor U11393 (N_11393,N_6015,N_2589);
nor U11394 (N_11394,N_4047,N_1237);
nand U11395 (N_11395,N_4220,N_4003);
xnor U11396 (N_11396,N_3559,N_5084);
and U11397 (N_11397,N_3218,N_5246);
nand U11398 (N_11398,N_3033,N_5750);
xnor U11399 (N_11399,N_1477,N_1191);
xnor U11400 (N_11400,N_2668,N_3356);
or U11401 (N_11401,N_5105,N_2970);
xnor U11402 (N_11402,N_2929,N_2044);
nor U11403 (N_11403,N_1781,N_1713);
nand U11404 (N_11404,N_1926,N_288);
nor U11405 (N_11405,N_6246,N_3412);
xor U11406 (N_11406,N_3401,N_5810);
and U11407 (N_11407,N_4530,N_1553);
or U11408 (N_11408,N_4208,N_446);
and U11409 (N_11409,N_225,N_3487);
nor U11410 (N_11410,N_4939,N_5094);
or U11411 (N_11411,N_2700,N_4619);
nand U11412 (N_11412,N_2380,N_476);
or U11413 (N_11413,N_6035,N_368);
nor U11414 (N_11414,N_5106,N_3485);
and U11415 (N_11415,N_4322,N_4734);
xor U11416 (N_11416,N_3234,N_821);
nor U11417 (N_11417,N_1166,N_975);
or U11418 (N_11418,N_5624,N_502);
xnor U11419 (N_11419,N_5792,N_5427);
xor U11420 (N_11420,N_3040,N_3353);
and U11421 (N_11421,N_4189,N_713);
nand U11422 (N_11422,N_1861,N_5198);
nand U11423 (N_11423,N_3297,N_3865);
and U11424 (N_11424,N_812,N_2953);
xnor U11425 (N_11425,N_3095,N_5179);
or U11426 (N_11426,N_5301,N_1002);
nor U11427 (N_11427,N_1988,N_471);
and U11428 (N_11428,N_3334,N_5499);
nand U11429 (N_11429,N_102,N_3266);
and U11430 (N_11430,N_5016,N_5404);
xnor U11431 (N_11431,N_5407,N_3188);
xor U11432 (N_11432,N_3540,N_2572);
xor U11433 (N_11433,N_1756,N_2481);
and U11434 (N_11434,N_1535,N_1281);
nor U11435 (N_11435,N_2060,N_1091);
or U11436 (N_11436,N_5786,N_701);
or U11437 (N_11437,N_3664,N_2952);
nand U11438 (N_11438,N_4332,N_4927);
xnor U11439 (N_11439,N_2966,N_5142);
nand U11440 (N_11440,N_2950,N_4129);
nand U11441 (N_11441,N_2607,N_917);
nand U11442 (N_11442,N_3667,N_3605);
or U11443 (N_11443,N_4009,N_425);
nor U11444 (N_11444,N_1264,N_1761);
or U11445 (N_11445,N_3854,N_4841);
xnor U11446 (N_11446,N_3461,N_1424);
xnor U11447 (N_11447,N_5840,N_663);
nor U11448 (N_11448,N_6075,N_5997);
or U11449 (N_11449,N_2844,N_5057);
xor U11450 (N_11450,N_429,N_6075);
xnor U11451 (N_11451,N_557,N_5025);
xnor U11452 (N_11452,N_5246,N_2481);
or U11453 (N_11453,N_2729,N_141);
xor U11454 (N_11454,N_5367,N_935);
xor U11455 (N_11455,N_2245,N_2913);
or U11456 (N_11456,N_1168,N_119);
nand U11457 (N_11457,N_1861,N_3416);
or U11458 (N_11458,N_4723,N_491);
or U11459 (N_11459,N_3017,N_5152);
or U11460 (N_11460,N_1842,N_2235);
xnor U11461 (N_11461,N_5341,N_3617);
nor U11462 (N_11462,N_3961,N_4402);
nor U11463 (N_11463,N_5708,N_3230);
nor U11464 (N_11464,N_4105,N_892);
nor U11465 (N_11465,N_5296,N_3514);
or U11466 (N_11466,N_859,N_3030);
and U11467 (N_11467,N_1011,N_4097);
xor U11468 (N_11468,N_5403,N_3785);
nor U11469 (N_11469,N_5407,N_134);
nor U11470 (N_11470,N_4918,N_1273);
and U11471 (N_11471,N_4274,N_3021);
nand U11472 (N_11472,N_3152,N_3055);
xor U11473 (N_11473,N_3305,N_3308);
xor U11474 (N_11474,N_4909,N_5020);
and U11475 (N_11475,N_2407,N_4193);
nor U11476 (N_11476,N_1634,N_2560);
nand U11477 (N_11477,N_463,N_625);
or U11478 (N_11478,N_218,N_2340);
nor U11479 (N_11479,N_713,N_4029);
nand U11480 (N_11480,N_39,N_4448);
xor U11481 (N_11481,N_4790,N_6109);
nor U11482 (N_11482,N_6218,N_2626);
nor U11483 (N_11483,N_2670,N_569);
and U11484 (N_11484,N_1354,N_3057);
nand U11485 (N_11485,N_2318,N_632);
and U11486 (N_11486,N_1855,N_1951);
and U11487 (N_11487,N_6214,N_5656);
nand U11488 (N_11488,N_2404,N_5300);
nand U11489 (N_11489,N_935,N_2843);
or U11490 (N_11490,N_72,N_3472);
nand U11491 (N_11491,N_1293,N_3747);
or U11492 (N_11492,N_804,N_5160);
or U11493 (N_11493,N_2288,N_3051);
xor U11494 (N_11494,N_5510,N_3174);
xor U11495 (N_11495,N_437,N_5386);
or U11496 (N_11496,N_4859,N_2534);
or U11497 (N_11497,N_354,N_1367);
xor U11498 (N_11498,N_1941,N_706);
xnor U11499 (N_11499,N_5270,N_4366);
or U11500 (N_11500,N_3214,N_140);
and U11501 (N_11501,N_2248,N_1392);
or U11502 (N_11502,N_3901,N_3856);
nor U11503 (N_11503,N_320,N_1069);
xnor U11504 (N_11504,N_4416,N_2825);
or U11505 (N_11505,N_388,N_2100);
nand U11506 (N_11506,N_1150,N_2293);
and U11507 (N_11507,N_2877,N_5101);
and U11508 (N_11508,N_1176,N_3668);
or U11509 (N_11509,N_10,N_5586);
nand U11510 (N_11510,N_1697,N_1222);
nand U11511 (N_11511,N_142,N_969);
or U11512 (N_11512,N_3585,N_4314);
nor U11513 (N_11513,N_5788,N_1551);
nand U11514 (N_11514,N_794,N_31);
nand U11515 (N_11515,N_1105,N_3951);
and U11516 (N_11516,N_5362,N_5914);
or U11517 (N_11517,N_138,N_6047);
and U11518 (N_11518,N_1990,N_4037);
nor U11519 (N_11519,N_5035,N_6097);
nor U11520 (N_11520,N_5636,N_2691);
or U11521 (N_11521,N_1228,N_3092);
nand U11522 (N_11522,N_3531,N_4457);
or U11523 (N_11523,N_4235,N_5554);
nand U11524 (N_11524,N_3055,N_4405);
nor U11525 (N_11525,N_3481,N_6194);
or U11526 (N_11526,N_1065,N_3819);
nand U11527 (N_11527,N_3546,N_3708);
nand U11528 (N_11528,N_2398,N_5694);
and U11529 (N_11529,N_2199,N_4847);
and U11530 (N_11530,N_3093,N_4349);
and U11531 (N_11531,N_5210,N_3016);
nand U11532 (N_11532,N_3980,N_428);
xnor U11533 (N_11533,N_3428,N_1853);
xor U11534 (N_11534,N_1536,N_1127);
nand U11535 (N_11535,N_5232,N_5957);
nor U11536 (N_11536,N_1264,N_2076);
and U11537 (N_11537,N_2766,N_3445);
or U11538 (N_11538,N_4367,N_1630);
or U11539 (N_11539,N_150,N_4856);
nand U11540 (N_11540,N_6210,N_2339);
and U11541 (N_11541,N_5089,N_2341);
or U11542 (N_11542,N_5226,N_4742);
xnor U11543 (N_11543,N_4913,N_1468);
or U11544 (N_11544,N_3220,N_3141);
or U11545 (N_11545,N_3516,N_1297);
or U11546 (N_11546,N_4892,N_3528);
nand U11547 (N_11547,N_5935,N_2761);
or U11548 (N_11548,N_755,N_2849);
or U11549 (N_11549,N_5767,N_3912);
nand U11550 (N_11550,N_3994,N_4734);
nand U11551 (N_11551,N_5605,N_208);
and U11552 (N_11552,N_1,N_1617);
nor U11553 (N_11553,N_5622,N_6088);
or U11554 (N_11554,N_3654,N_1481);
and U11555 (N_11555,N_244,N_2406);
or U11556 (N_11556,N_2069,N_4313);
xor U11557 (N_11557,N_4326,N_2905);
nor U11558 (N_11558,N_5579,N_48);
and U11559 (N_11559,N_4584,N_3165);
nand U11560 (N_11560,N_730,N_1136);
or U11561 (N_11561,N_3473,N_4041);
xor U11562 (N_11562,N_776,N_1099);
nand U11563 (N_11563,N_5489,N_4096);
xnor U11564 (N_11564,N_128,N_5659);
xor U11565 (N_11565,N_3765,N_2608);
or U11566 (N_11566,N_2747,N_4044);
or U11567 (N_11567,N_5006,N_1806);
xor U11568 (N_11568,N_323,N_1350);
xnor U11569 (N_11569,N_1619,N_976);
nand U11570 (N_11570,N_2801,N_757);
xor U11571 (N_11571,N_142,N_2977);
or U11572 (N_11572,N_141,N_5896);
nand U11573 (N_11573,N_5410,N_5266);
or U11574 (N_11574,N_898,N_3134);
nor U11575 (N_11575,N_5986,N_3318);
nor U11576 (N_11576,N_4459,N_5836);
nand U11577 (N_11577,N_3865,N_5819);
nand U11578 (N_11578,N_4080,N_4230);
and U11579 (N_11579,N_1380,N_2832);
or U11580 (N_11580,N_5194,N_4800);
nor U11581 (N_11581,N_2443,N_4411);
and U11582 (N_11582,N_5302,N_3047);
or U11583 (N_11583,N_1595,N_3452);
or U11584 (N_11584,N_5744,N_2750);
and U11585 (N_11585,N_3347,N_707);
nor U11586 (N_11586,N_227,N_2437);
or U11587 (N_11587,N_6200,N_6144);
nor U11588 (N_11588,N_5795,N_4666);
nand U11589 (N_11589,N_6120,N_2751);
and U11590 (N_11590,N_4079,N_1983);
nor U11591 (N_11591,N_4825,N_1461);
and U11592 (N_11592,N_998,N_6006);
and U11593 (N_11593,N_6013,N_2602);
xnor U11594 (N_11594,N_904,N_4066);
or U11595 (N_11595,N_5722,N_3575);
and U11596 (N_11596,N_383,N_5811);
and U11597 (N_11597,N_5461,N_2114);
xor U11598 (N_11598,N_3796,N_3749);
xor U11599 (N_11599,N_3425,N_15);
nand U11600 (N_11600,N_3665,N_1070);
and U11601 (N_11601,N_5897,N_5123);
nor U11602 (N_11602,N_1324,N_4584);
xor U11603 (N_11603,N_3874,N_3165);
or U11604 (N_11604,N_5138,N_2843);
xor U11605 (N_11605,N_1983,N_5436);
nor U11606 (N_11606,N_5022,N_5853);
xor U11607 (N_11607,N_5919,N_4563);
xnor U11608 (N_11608,N_225,N_3950);
nor U11609 (N_11609,N_2163,N_1499);
or U11610 (N_11610,N_5318,N_5669);
nand U11611 (N_11611,N_2073,N_531);
nand U11612 (N_11612,N_4648,N_2719);
nor U11613 (N_11613,N_4463,N_1957);
nor U11614 (N_11614,N_5183,N_6197);
xor U11615 (N_11615,N_2590,N_1353);
xnor U11616 (N_11616,N_4170,N_1358);
or U11617 (N_11617,N_5861,N_1373);
nand U11618 (N_11618,N_4768,N_2198);
or U11619 (N_11619,N_475,N_5515);
and U11620 (N_11620,N_4887,N_2090);
nor U11621 (N_11621,N_1216,N_2496);
nor U11622 (N_11622,N_2063,N_1427);
or U11623 (N_11623,N_4493,N_5900);
nor U11624 (N_11624,N_1129,N_3573);
xnor U11625 (N_11625,N_5982,N_2359);
xor U11626 (N_11626,N_6006,N_6047);
xor U11627 (N_11627,N_499,N_3052);
and U11628 (N_11628,N_5099,N_2860);
nand U11629 (N_11629,N_1538,N_1489);
nor U11630 (N_11630,N_826,N_1659);
nor U11631 (N_11631,N_3721,N_4856);
and U11632 (N_11632,N_1012,N_513);
and U11633 (N_11633,N_3958,N_3852);
nor U11634 (N_11634,N_1918,N_2445);
nor U11635 (N_11635,N_3114,N_2407);
xnor U11636 (N_11636,N_3101,N_3414);
xor U11637 (N_11637,N_1840,N_3203);
nand U11638 (N_11638,N_1917,N_2104);
nor U11639 (N_11639,N_4141,N_345);
nand U11640 (N_11640,N_3792,N_3398);
nor U11641 (N_11641,N_5754,N_632);
or U11642 (N_11642,N_1640,N_3495);
or U11643 (N_11643,N_5326,N_5475);
xor U11644 (N_11644,N_250,N_4330);
nor U11645 (N_11645,N_4938,N_5498);
or U11646 (N_11646,N_1281,N_5093);
or U11647 (N_11647,N_835,N_129);
nor U11648 (N_11648,N_1740,N_511);
or U11649 (N_11649,N_1412,N_4750);
nand U11650 (N_11650,N_2683,N_2670);
nor U11651 (N_11651,N_4290,N_4798);
nand U11652 (N_11652,N_5839,N_5936);
and U11653 (N_11653,N_5275,N_2162);
xor U11654 (N_11654,N_2369,N_4772);
and U11655 (N_11655,N_2877,N_2712);
and U11656 (N_11656,N_1425,N_520);
nor U11657 (N_11657,N_6068,N_6069);
nor U11658 (N_11658,N_445,N_6128);
nor U11659 (N_11659,N_5803,N_701);
xnor U11660 (N_11660,N_1208,N_2519);
nand U11661 (N_11661,N_5945,N_149);
xnor U11662 (N_11662,N_1687,N_4161);
nor U11663 (N_11663,N_61,N_5092);
nor U11664 (N_11664,N_3794,N_6128);
nand U11665 (N_11665,N_4424,N_543);
nand U11666 (N_11666,N_4549,N_3498);
or U11667 (N_11667,N_5195,N_1711);
nor U11668 (N_11668,N_3,N_2632);
and U11669 (N_11669,N_3816,N_5313);
nor U11670 (N_11670,N_4645,N_3937);
nand U11671 (N_11671,N_4811,N_4526);
and U11672 (N_11672,N_4393,N_1420);
nand U11673 (N_11673,N_2331,N_2572);
or U11674 (N_11674,N_5892,N_4814);
xnor U11675 (N_11675,N_1685,N_1619);
nand U11676 (N_11676,N_3588,N_6229);
xor U11677 (N_11677,N_4309,N_3042);
or U11678 (N_11678,N_2499,N_3398);
nand U11679 (N_11679,N_5651,N_4403);
xor U11680 (N_11680,N_5585,N_4106);
nand U11681 (N_11681,N_787,N_1831);
xor U11682 (N_11682,N_2309,N_837);
xnor U11683 (N_11683,N_3523,N_3269);
nor U11684 (N_11684,N_240,N_5035);
nor U11685 (N_11685,N_5241,N_2379);
xnor U11686 (N_11686,N_1866,N_5984);
and U11687 (N_11687,N_2847,N_4117);
nor U11688 (N_11688,N_4382,N_948);
nor U11689 (N_11689,N_5974,N_3049);
nor U11690 (N_11690,N_3052,N_3661);
xor U11691 (N_11691,N_2514,N_2856);
or U11692 (N_11692,N_902,N_1392);
and U11693 (N_11693,N_743,N_99);
and U11694 (N_11694,N_5093,N_6045);
nor U11695 (N_11695,N_2773,N_360);
nand U11696 (N_11696,N_4255,N_224);
or U11697 (N_11697,N_736,N_5680);
nor U11698 (N_11698,N_3882,N_5877);
xor U11699 (N_11699,N_3755,N_3005);
or U11700 (N_11700,N_935,N_6243);
and U11701 (N_11701,N_4773,N_4318);
nor U11702 (N_11702,N_2613,N_3387);
nor U11703 (N_11703,N_2110,N_3266);
xnor U11704 (N_11704,N_2388,N_5799);
nor U11705 (N_11705,N_783,N_588);
and U11706 (N_11706,N_4172,N_947);
nand U11707 (N_11707,N_5213,N_2325);
nor U11708 (N_11708,N_5867,N_440);
xnor U11709 (N_11709,N_5947,N_3416);
nor U11710 (N_11710,N_5117,N_6229);
or U11711 (N_11711,N_3720,N_546);
xnor U11712 (N_11712,N_2729,N_3831);
and U11713 (N_11713,N_3537,N_2687);
nand U11714 (N_11714,N_4897,N_39);
nor U11715 (N_11715,N_4214,N_5187);
nor U11716 (N_11716,N_5270,N_1913);
and U11717 (N_11717,N_3855,N_132);
nor U11718 (N_11718,N_4788,N_1381);
nand U11719 (N_11719,N_6232,N_5542);
nor U11720 (N_11720,N_5263,N_896);
xnor U11721 (N_11721,N_4286,N_1583);
nor U11722 (N_11722,N_122,N_82);
and U11723 (N_11723,N_4165,N_5427);
and U11724 (N_11724,N_4574,N_4363);
or U11725 (N_11725,N_4295,N_6188);
xor U11726 (N_11726,N_1183,N_1570);
and U11727 (N_11727,N_1539,N_1882);
xor U11728 (N_11728,N_2561,N_4317);
and U11729 (N_11729,N_4178,N_5248);
and U11730 (N_11730,N_3044,N_2509);
nand U11731 (N_11731,N_5513,N_6132);
xor U11732 (N_11732,N_5786,N_420);
xor U11733 (N_11733,N_1239,N_2924);
nor U11734 (N_11734,N_5825,N_4468);
and U11735 (N_11735,N_1,N_3040);
nand U11736 (N_11736,N_6018,N_367);
and U11737 (N_11737,N_1561,N_3336);
xor U11738 (N_11738,N_685,N_3297);
and U11739 (N_11739,N_5535,N_3402);
nand U11740 (N_11740,N_2053,N_5928);
and U11741 (N_11741,N_93,N_958);
and U11742 (N_11742,N_4077,N_5689);
or U11743 (N_11743,N_5791,N_3242);
nor U11744 (N_11744,N_1306,N_5596);
nand U11745 (N_11745,N_5704,N_1298);
nor U11746 (N_11746,N_2013,N_2046);
nor U11747 (N_11747,N_5698,N_1963);
nor U11748 (N_11748,N_1056,N_3790);
xnor U11749 (N_11749,N_3303,N_1149);
and U11750 (N_11750,N_3958,N_3241);
and U11751 (N_11751,N_4921,N_1962);
or U11752 (N_11752,N_3051,N_3639);
nand U11753 (N_11753,N_832,N_3787);
or U11754 (N_11754,N_2234,N_4051);
or U11755 (N_11755,N_201,N_5482);
nand U11756 (N_11756,N_346,N_2111);
nor U11757 (N_11757,N_497,N_1112);
nor U11758 (N_11758,N_5476,N_3629);
xor U11759 (N_11759,N_4447,N_5948);
nor U11760 (N_11760,N_2350,N_279);
nand U11761 (N_11761,N_4560,N_4432);
nor U11762 (N_11762,N_1856,N_6007);
xnor U11763 (N_11763,N_491,N_3036);
or U11764 (N_11764,N_4232,N_3505);
nand U11765 (N_11765,N_5892,N_575);
nand U11766 (N_11766,N_2123,N_4243);
and U11767 (N_11767,N_685,N_3689);
xor U11768 (N_11768,N_5605,N_2968);
nand U11769 (N_11769,N_199,N_5233);
and U11770 (N_11770,N_4526,N_5875);
nor U11771 (N_11771,N_4084,N_741);
nor U11772 (N_11772,N_4329,N_5223);
and U11773 (N_11773,N_3709,N_3266);
nand U11774 (N_11774,N_3012,N_149);
or U11775 (N_11775,N_3845,N_2092);
or U11776 (N_11776,N_10,N_4104);
nor U11777 (N_11777,N_2299,N_2872);
or U11778 (N_11778,N_1448,N_3597);
xnor U11779 (N_11779,N_4537,N_5799);
or U11780 (N_11780,N_1220,N_1539);
and U11781 (N_11781,N_3768,N_1911);
nor U11782 (N_11782,N_365,N_2872);
nor U11783 (N_11783,N_3269,N_1972);
or U11784 (N_11784,N_4070,N_4751);
and U11785 (N_11785,N_3352,N_2410);
and U11786 (N_11786,N_2467,N_2414);
xnor U11787 (N_11787,N_3724,N_4215);
nand U11788 (N_11788,N_3154,N_2752);
xnor U11789 (N_11789,N_3557,N_4113);
nand U11790 (N_11790,N_4040,N_55);
and U11791 (N_11791,N_3586,N_862);
xor U11792 (N_11792,N_3321,N_1860);
nor U11793 (N_11793,N_3211,N_5422);
and U11794 (N_11794,N_125,N_1511);
nand U11795 (N_11795,N_790,N_50);
or U11796 (N_11796,N_2055,N_2104);
and U11797 (N_11797,N_5375,N_2724);
and U11798 (N_11798,N_585,N_3365);
nand U11799 (N_11799,N_725,N_554);
and U11800 (N_11800,N_1920,N_94);
xor U11801 (N_11801,N_682,N_5835);
nor U11802 (N_11802,N_4432,N_636);
and U11803 (N_11803,N_167,N_3296);
nor U11804 (N_11804,N_842,N_3584);
or U11805 (N_11805,N_836,N_3192);
xor U11806 (N_11806,N_1758,N_2686);
nor U11807 (N_11807,N_474,N_1426);
and U11808 (N_11808,N_3401,N_6095);
nand U11809 (N_11809,N_4299,N_1190);
and U11810 (N_11810,N_2448,N_4206);
xnor U11811 (N_11811,N_6139,N_2578);
nand U11812 (N_11812,N_5193,N_2575);
or U11813 (N_11813,N_5657,N_5566);
nand U11814 (N_11814,N_1666,N_1155);
xor U11815 (N_11815,N_2735,N_5218);
or U11816 (N_11816,N_1612,N_296);
and U11817 (N_11817,N_6016,N_5476);
nand U11818 (N_11818,N_5372,N_4837);
or U11819 (N_11819,N_4214,N_2230);
or U11820 (N_11820,N_3213,N_1448);
nor U11821 (N_11821,N_6213,N_2609);
and U11822 (N_11822,N_3520,N_6000);
and U11823 (N_11823,N_5240,N_743);
xnor U11824 (N_11824,N_3198,N_6127);
or U11825 (N_11825,N_331,N_5485);
and U11826 (N_11826,N_74,N_2425);
nor U11827 (N_11827,N_4017,N_2220);
nor U11828 (N_11828,N_5805,N_3648);
nor U11829 (N_11829,N_3770,N_115);
nor U11830 (N_11830,N_3848,N_5897);
nand U11831 (N_11831,N_5544,N_5613);
nor U11832 (N_11832,N_6125,N_812);
or U11833 (N_11833,N_3920,N_68);
nor U11834 (N_11834,N_5303,N_538);
xnor U11835 (N_11835,N_5724,N_5920);
and U11836 (N_11836,N_944,N_5753);
nor U11837 (N_11837,N_288,N_5427);
and U11838 (N_11838,N_557,N_5807);
nor U11839 (N_11839,N_1937,N_6114);
or U11840 (N_11840,N_6066,N_2816);
xor U11841 (N_11841,N_4974,N_3804);
nor U11842 (N_11842,N_3786,N_5116);
nor U11843 (N_11843,N_3481,N_4178);
and U11844 (N_11844,N_5449,N_1741);
or U11845 (N_11845,N_358,N_3488);
nand U11846 (N_11846,N_3693,N_2548);
nor U11847 (N_11847,N_2615,N_4377);
and U11848 (N_11848,N_658,N_5585);
nand U11849 (N_11849,N_2849,N_1761);
xor U11850 (N_11850,N_3083,N_3595);
and U11851 (N_11851,N_2111,N_6104);
nand U11852 (N_11852,N_1187,N_1471);
xor U11853 (N_11853,N_3365,N_5955);
nor U11854 (N_11854,N_5464,N_3827);
and U11855 (N_11855,N_71,N_2325);
nand U11856 (N_11856,N_1136,N_3614);
nor U11857 (N_11857,N_4331,N_6117);
or U11858 (N_11858,N_4807,N_1566);
and U11859 (N_11859,N_611,N_3945);
or U11860 (N_11860,N_3689,N_4770);
nand U11861 (N_11861,N_696,N_3946);
or U11862 (N_11862,N_356,N_6170);
xnor U11863 (N_11863,N_4598,N_3239);
xor U11864 (N_11864,N_5481,N_6199);
or U11865 (N_11865,N_3117,N_815);
and U11866 (N_11866,N_3570,N_2703);
and U11867 (N_11867,N_2768,N_45);
or U11868 (N_11868,N_1134,N_834);
nand U11869 (N_11869,N_1327,N_2861);
and U11870 (N_11870,N_2003,N_1930);
xnor U11871 (N_11871,N_5458,N_5811);
or U11872 (N_11872,N_3270,N_2423);
xor U11873 (N_11873,N_985,N_4183);
xor U11874 (N_11874,N_3639,N_5655);
or U11875 (N_11875,N_1580,N_6005);
xor U11876 (N_11876,N_3292,N_3201);
nor U11877 (N_11877,N_3984,N_6043);
and U11878 (N_11878,N_4178,N_787);
or U11879 (N_11879,N_228,N_2552);
nor U11880 (N_11880,N_1045,N_694);
and U11881 (N_11881,N_5344,N_6231);
xor U11882 (N_11882,N_4370,N_5334);
and U11883 (N_11883,N_5194,N_3894);
xor U11884 (N_11884,N_3473,N_482);
nand U11885 (N_11885,N_1678,N_2777);
xnor U11886 (N_11886,N_465,N_4053);
or U11887 (N_11887,N_326,N_3737);
xnor U11888 (N_11888,N_1549,N_5737);
xor U11889 (N_11889,N_1261,N_593);
or U11890 (N_11890,N_4625,N_2382);
or U11891 (N_11891,N_957,N_5658);
or U11892 (N_11892,N_3126,N_4651);
and U11893 (N_11893,N_1359,N_505);
and U11894 (N_11894,N_1500,N_4921);
or U11895 (N_11895,N_2769,N_4136);
or U11896 (N_11896,N_1592,N_3428);
nor U11897 (N_11897,N_5115,N_346);
xor U11898 (N_11898,N_276,N_2099);
and U11899 (N_11899,N_3617,N_2110);
or U11900 (N_11900,N_1874,N_5920);
xnor U11901 (N_11901,N_2433,N_4973);
nand U11902 (N_11902,N_5850,N_4008);
xnor U11903 (N_11903,N_5424,N_1802);
nor U11904 (N_11904,N_5210,N_4960);
or U11905 (N_11905,N_1669,N_4297);
and U11906 (N_11906,N_6098,N_2728);
and U11907 (N_11907,N_5913,N_4806);
nor U11908 (N_11908,N_1713,N_4083);
nand U11909 (N_11909,N_4326,N_1373);
nor U11910 (N_11910,N_2256,N_1566);
or U11911 (N_11911,N_5624,N_626);
and U11912 (N_11912,N_367,N_6232);
nor U11913 (N_11913,N_5680,N_268);
nand U11914 (N_11914,N_87,N_2214);
or U11915 (N_11915,N_151,N_1293);
nor U11916 (N_11916,N_2910,N_489);
nand U11917 (N_11917,N_5004,N_3784);
and U11918 (N_11918,N_2318,N_4796);
and U11919 (N_11919,N_1111,N_6055);
xor U11920 (N_11920,N_277,N_608);
nand U11921 (N_11921,N_4143,N_416);
or U11922 (N_11922,N_3705,N_4759);
xor U11923 (N_11923,N_539,N_4771);
nand U11924 (N_11924,N_2082,N_4578);
or U11925 (N_11925,N_1843,N_1157);
nand U11926 (N_11926,N_154,N_577);
xnor U11927 (N_11927,N_1804,N_1259);
nand U11928 (N_11928,N_779,N_1483);
nand U11929 (N_11929,N_4132,N_5183);
and U11930 (N_11930,N_657,N_2817);
nor U11931 (N_11931,N_269,N_6207);
xor U11932 (N_11932,N_4458,N_2585);
and U11933 (N_11933,N_1789,N_6014);
nor U11934 (N_11934,N_5085,N_724);
nand U11935 (N_11935,N_294,N_5764);
and U11936 (N_11936,N_2330,N_727);
xor U11937 (N_11937,N_2455,N_2474);
or U11938 (N_11938,N_2059,N_5084);
xnor U11939 (N_11939,N_2158,N_2350);
nand U11940 (N_11940,N_4864,N_3300);
nand U11941 (N_11941,N_2086,N_4512);
and U11942 (N_11942,N_371,N_5554);
nor U11943 (N_11943,N_4832,N_1359);
or U11944 (N_11944,N_6007,N_1909);
nand U11945 (N_11945,N_4593,N_238);
and U11946 (N_11946,N_3139,N_2206);
nor U11947 (N_11947,N_5022,N_1710);
nor U11948 (N_11948,N_1468,N_4637);
nor U11949 (N_11949,N_527,N_3176);
xor U11950 (N_11950,N_2643,N_5003);
nor U11951 (N_11951,N_4055,N_327);
xnor U11952 (N_11952,N_4552,N_250);
xnor U11953 (N_11953,N_2420,N_1574);
and U11954 (N_11954,N_5987,N_371);
xor U11955 (N_11955,N_4623,N_5530);
and U11956 (N_11956,N_1864,N_5148);
nor U11957 (N_11957,N_3248,N_4267);
nor U11958 (N_11958,N_5850,N_2618);
nor U11959 (N_11959,N_1768,N_1097);
nand U11960 (N_11960,N_1156,N_2169);
nor U11961 (N_11961,N_5547,N_1302);
nand U11962 (N_11962,N_717,N_1978);
and U11963 (N_11963,N_3558,N_5771);
nand U11964 (N_11964,N_4667,N_1066);
and U11965 (N_11965,N_3130,N_5020);
and U11966 (N_11966,N_1231,N_5096);
nand U11967 (N_11967,N_141,N_4083);
and U11968 (N_11968,N_5284,N_1079);
xor U11969 (N_11969,N_5393,N_3076);
and U11970 (N_11970,N_1229,N_2173);
nand U11971 (N_11971,N_4495,N_1693);
and U11972 (N_11972,N_2231,N_4164);
nor U11973 (N_11973,N_3120,N_5782);
xnor U11974 (N_11974,N_2534,N_4814);
or U11975 (N_11975,N_1934,N_4264);
nor U11976 (N_11976,N_3878,N_4876);
or U11977 (N_11977,N_4368,N_3334);
nand U11978 (N_11978,N_5405,N_1773);
nand U11979 (N_11979,N_773,N_3453);
or U11980 (N_11980,N_6012,N_6246);
xor U11981 (N_11981,N_4736,N_3239);
xor U11982 (N_11982,N_1920,N_2387);
or U11983 (N_11983,N_2514,N_3539);
or U11984 (N_11984,N_344,N_3152);
or U11985 (N_11985,N_4331,N_5216);
and U11986 (N_11986,N_2254,N_5474);
and U11987 (N_11987,N_1981,N_5791);
and U11988 (N_11988,N_5447,N_3983);
xor U11989 (N_11989,N_1039,N_5642);
and U11990 (N_11990,N_5624,N_3820);
xor U11991 (N_11991,N_5396,N_4959);
nor U11992 (N_11992,N_2457,N_1088);
xor U11993 (N_11993,N_5716,N_2617);
nor U11994 (N_11994,N_1183,N_5473);
nand U11995 (N_11995,N_5963,N_4801);
or U11996 (N_11996,N_3420,N_1978);
nand U11997 (N_11997,N_5261,N_478);
nand U11998 (N_11998,N_3271,N_1789);
nand U11999 (N_11999,N_766,N_2206);
or U12000 (N_12000,N_3707,N_269);
nand U12001 (N_12001,N_5208,N_1173);
nor U12002 (N_12002,N_1431,N_5656);
nor U12003 (N_12003,N_5413,N_4037);
xnor U12004 (N_12004,N_340,N_880);
nand U12005 (N_12005,N_1442,N_1780);
xor U12006 (N_12006,N_5690,N_340);
xnor U12007 (N_12007,N_4689,N_4067);
and U12008 (N_12008,N_4527,N_3497);
and U12009 (N_12009,N_3931,N_4975);
or U12010 (N_12010,N_458,N_2553);
nand U12011 (N_12011,N_3801,N_1180);
and U12012 (N_12012,N_2189,N_2527);
and U12013 (N_12013,N_6155,N_5573);
and U12014 (N_12014,N_6126,N_355);
nand U12015 (N_12015,N_6142,N_4783);
and U12016 (N_12016,N_4674,N_3756);
xor U12017 (N_12017,N_3262,N_4057);
nor U12018 (N_12018,N_1043,N_756);
and U12019 (N_12019,N_5163,N_3157);
nor U12020 (N_12020,N_2689,N_3904);
or U12021 (N_12021,N_4381,N_1525);
nand U12022 (N_12022,N_5165,N_1595);
nor U12023 (N_12023,N_214,N_1999);
nor U12024 (N_12024,N_5661,N_1309);
and U12025 (N_12025,N_5488,N_4269);
and U12026 (N_12026,N_2182,N_3997);
xnor U12027 (N_12027,N_1328,N_2948);
nand U12028 (N_12028,N_2755,N_1831);
xnor U12029 (N_12029,N_6044,N_2988);
and U12030 (N_12030,N_3245,N_1277);
and U12031 (N_12031,N_2566,N_1784);
nand U12032 (N_12032,N_2810,N_3996);
and U12033 (N_12033,N_1038,N_4474);
nand U12034 (N_12034,N_2468,N_1741);
and U12035 (N_12035,N_3337,N_4239);
nand U12036 (N_12036,N_3532,N_5194);
nor U12037 (N_12037,N_3244,N_1613);
or U12038 (N_12038,N_5707,N_4364);
xnor U12039 (N_12039,N_980,N_2872);
or U12040 (N_12040,N_3691,N_368);
nor U12041 (N_12041,N_5254,N_3245);
and U12042 (N_12042,N_1125,N_5230);
or U12043 (N_12043,N_5274,N_4373);
nand U12044 (N_12044,N_1615,N_580);
xor U12045 (N_12045,N_477,N_3491);
nand U12046 (N_12046,N_1251,N_5796);
and U12047 (N_12047,N_6048,N_3900);
nor U12048 (N_12048,N_4994,N_4863);
nand U12049 (N_12049,N_1100,N_5148);
nand U12050 (N_12050,N_3512,N_3587);
xor U12051 (N_12051,N_517,N_2926);
xor U12052 (N_12052,N_756,N_3049);
xor U12053 (N_12053,N_2742,N_3692);
and U12054 (N_12054,N_5045,N_6197);
or U12055 (N_12055,N_5807,N_5269);
or U12056 (N_12056,N_5580,N_4149);
nor U12057 (N_12057,N_3979,N_232);
nor U12058 (N_12058,N_492,N_5505);
and U12059 (N_12059,N_5568,N_4789);
or U12060 (N_12060,N_1971,N_5146);
nand U12061 (N_12061,N_2878,N_5464);
or U12062 (N_12062,N_6114,N_754);
and U12063 (N_12063,N_4861,N_446);
and U12064 (N_12064,N_5744,N_3755);
or U12065 (N_12065,N_4914,N_381);
xnor U12066 (N_12066,N_3367,N_2832);
xnor U12067 (N_12067,N_2595,N_5450);
or U12068 (N_12068,N_2281,N_589);
and U12069 (N_12069,N_3163,N_4654);
nand U12070 (N_12070,N_1494,N_1031);
xor U12071 (N_12071,N_5468,N_1457);
and U12072 (N_12072,N_2374,N_3782);
xnor U12073 (N_12073,N_399,N_2877);
or U12074 (N_12074,N_4763,N_3556);
and U12075 (N_12075,N_1113,N_2436);
or U12076 (N_12076,N_2908,N_4370);
nand U12077 (N_12077,N_457,N_5311);
or U12078 (N_12078,N_1676,N_2431);
and U12079 (N_12079,N_1272,N_4846);
or U12080 (N_12080,N_2333,N_797);
or U12081 (N_12081,N_4002,N_5040);
and U12082 (N_12082,N_5880,N_326);
nand U12083 (N_12083,N_4951,N_1903);
or U12084 (N_12084,N_1948,N_4283);
or U12085 (N_12085,N_4157,N_262);
xnor U12086 (N_12086,N_6160,N_1938);
nor U12087 (N_12087,N_2679,N_557);
or U12088 (N_12088,N_1602,N_4350);
xor U12089 (N_12089,N_2815,N_2284);
and U12090 (N_12090,N_6048,N_648);
xnor U12091 (N_12091,N_3675,N_4161);
or U12092 (N_12092,N_5634,N_613);
and U12093 (N_12093,N_2226,N_3372);
xor U12094 (N_12094,N_4157,N_6177);
and U12095 (N_12095,N_6162,N_938);
nor U12096 (N_12096,N_3278,N_5482);
xnor U12097 (N_12097,N_4564,N_1143);
or U12098 (N_12098,N_1219,N_2090);
xnor U12099 (N_12099,N_4723,N_1339);
xnor U12100 (N_12100,N_4725,N_1362);
and U12101 (N_12101,N_1974,N_2660);
nor U12102 (N_12102,N_2143,N_5809);
and U12103 (N_12103,N_3855,N_2321);
or U12104 (N_12104,N_3789,N_5301);
and U12105 (N_12105,N_4527,N_2684);
and U12106 (N_12106,N_4427,N_5906);
nor U12107 (N_12107,N_358,N_1229);
or U12108 (N_12108,N_1474,N_2893);
and U12109 (N_12109,N_3233,N_4386);
or U12110 (N_12110,N_4188,N_6175);
nand U12111 (N_12111,N_4217,N_5366);
nand U12112 (N_12112,N_5550,N_950);
xnor U12113 (N_12113,N_2849,N_704);
nand U12114 (N_12114,N_382,N_957);
and U12115 (N_12115,N_1634,N_5161);
or U12116 (N_12116,N_2059,N_1129);
xor U12117 (N_12117,N_1911,N_4512);
nand U12118 (N_12118,N_4056,N_5739);
and U12119 (N_12119,N_3574,N_3516);
and U12120 (N_12120,N_2842,N_5655);
xnor U12121 (N_12121,N_2668,N_2546);
nor U12122 (N_12122,N_3777,N_3279);
xnor U12123 (N_12123,N_1454,N_4429);
nor U12124 (N_12124,N_4357,N_4981);
nand U12125 (N_12125,N_5760,N_1995);
or U12126 (N_12126,N_2929,N_2725);
xnor U12127 (N_12127,N_55,N_1963);
and U12128 (N_12128,N_2784,N_5401);
nor U12129 (N_12129,N_2499,N_2032);
nand U12130 (N_12130,N_4001,N_2129);
xor U12131 (N_12131,N_5370,N_2581);
nand U12132 (N_12132,N_2638,N_4203);
nand U12133 (N_12133,N_2468,N_4279);
nand U12134 (N_12134,N_2498,N_4111);
and U12135 (N_12135,N_5742,N_3792);
and U12136 (N_12136,N_1612,N_3991);
and U12137 (N_12137,N_1329,N_6062);
nor U12138 (N_12138,N_1893,N_1213);
xnor U12139 (N_12139,N_5525,N_5318);
or U12140 (N_12140,N_5431,N_3124);
nor U12141 (N_12141,N_1016,N_4119);
xnor U12142 (N_12142,N_1818,N_640);
and U12143 (N_12143,N_3807,N_3738);
xnor U12144 (N_12144,N_3501,N_364);
and U12145 (N_12145,N_3208,N_6096);
and U12146 (N_12146,N_285,N_5019);
and U12147 (N_12147,N_5596,N_4530);
xnor U12148 (N_12148,N_4774,N_3370);
xor U12149 (N_12149,N_2929,N_4143);
xor U12150 (N_12150,N_3376,N_6184);
nand U12151 (N_12151,N_2578,N_2226);
xor U12152 (N_12152,N_286,N_4006);
nand U12153 (N_12153,N_895,N_607);
or U12154 (N_12154,N_2130,N_4781);
nor U12155 (N_12155,N_1065,N_2461);
nand U12156 (N_12156,N_3224,N_1898);
xor U12157 (N_12157,N_16,N_1921);
or U12158 (N_12158,N_2551,N_2964);
or U12159 (N_12159,N_5536,N_2478);
nor U12160 (N_12160,N_4875,N_290);
nor U12161 (N_12161,N_4644,N_5633);
nor U12162 (N_12162,N_4673,N_4595);
and U12163 (N_12163,N_680,N_3626);
nand U12164 (N_12164,N_3323,N_2458);
and U12165 (N_12165,N_4297,N_2046);
xnor U12166 (N_12166,N_5005,N_1961);
nor U12167 (N_12167,N_2331,N_5188);
xor U12168 (N_12168,N_3850,N_799);
nand U12169 (N_12169,N_1418,N_6104);
nand U12170 (N_12170,N_1391,N_4044);
xor U12171 (N_12171,N_2711,N_597);
or U12172 (N_12172,N_3106,N_1764);
or U12173 (N_12173,N_1496,N_2721);
nor U12174 (N_12174,N_41,N_784);
xor U12175 (N_12175,N_4743,N_3724);
nand U12176 (N_12176,N_2244,N_5058);
xor U12177 (N_12177,N_5466,N_918);
or U12178 (N_12178,N_3327,N_2217);
or U12179 (N_12179,N_3131,N_1898);
or U12180 (N_12180,N_194,N_713);
or U12181 (N_12181,N_2969,N_3777);
nand U12182 (N_12182,N_4514,N_2092);
nor U12183 (N_12183,N_553,N_561);
nor U12184 (N_12184,N_280,N_2661);
nor U12185 (N_12185,N_1656,N_6107);
and U12186 (N_12186,N_2229,N_3918);
xnor U12187 (N_12187,N_6238,N_626);
or U12188 (N_12188,N_3009,N_3894);
xor U12189 (N_12189,N_3636,N_6214);
and U12190 (N_12190,N_4452,N_6125);
nand U12191 (N_12191,N_3488,N_1213);
or U12192 (N_12192,N_3298,N_4203);
nand U12193 (N_12193,N_1204,N_5529);
and U12194 (N_12194,N_2830,N_3441);
nand U12195 (N_12195,N_2786,N_3745);
nand U12196 (N_12196,N_6124,N_3588);
nor U12197 (N_12197,N_3485,N_1535);
nand U12198 (N_12198,N_3875,N_1354);
nor U12199 (N_12199,N_5088,N_918);
and U12200 (N_12200,N_5324,N_1477);
xor U12201 (N_12201,N_4941,N_1380);
or U12202 (N_12202,N_1366,N_4253);
xnor U12203 (N_12203,N_1589,N_3947);
xnor U12204 (N_12204,N_1599,N_4107);
and U12205 (N_12205,N_425,N_1163);
nand U12206 (N_12206,N_2786,N_2243);
and U12207 (N_12207,N_5654,N_393);
or U12208 (N_12208,N_5780,N_866);
and U12209 (N_12209,N_3315,N_3481);
xor U12210 (N_12210,N_4573,N_3436);
or U12211 (N_12211,N_3586,N_3197);
nor U12212 (N_12212,N_172,N_169);
nor U12213 (N_12213,N_1928,N_804);
nand U12214 (N_12214,N_5851,N_3434);
xnor U12215 (N_12215,N_5028,N_2875);
nand U12216 (N_12216,N_3211,N_699);
or U12217 (N_12217,N_1589,N_5605);
nand U12218 (N_12218,N_2006,N_5260);
nor U12219 (N_12219,N_5941,N_5134);
or U12220 (N_12220,N_2713,N_1084);
xnor U12221 (N_12221,N_3511,N_2800);
nand U12222 (N_12222,N_1000,N_1888);
or U12223 (N_12223,N_6092,N_935);
nand U12224 (N_12224,N_5857,N_2212);
or U12225 (N_12225,N_4615,N_5995);
nand U12226 (N_12226,N_1093,N_5589);
nand U12227 (N_12227,N_3603,N_3773);
or U12228 (N_12228,N_5372,N_569);
nor U12229 (N_12229,N_1440,N_1735);
and U12230 (N_12230,N_4231,N_243);
nor U12231 (N_12231,N_2631,N_1996);
xor U12232 (N_12232,N_1194,N_3319);
xnor U12233 (N_12233,N_594,N_2699);
nand U12234 (N_12234,N_4471,N_5742);
or U12235 (N_12235,N_4141,N_3952);
or U12236 (N_12236,N_291,N_4176);
and U12237 (N_12237,N_3631,N_2113);
nand U12238 (N_12238,N_3714,N_5204);
nand U12239 (N_12239,N_2127,N_262);
or U12240 (N_12240,N_5866,N_1533);
xor U12241 (N_12241,N_4896,N_3374);
nor U12242 (N_12242,N_5627,N_3505);
nor U12243 (N_12243,N_5653,N_2401);
xor U12244 (N_12244,N_1270,N_2789);
or U12245 (N_12245,N_2928,N_3664);
nor U12246 (N_12246,N_3870,N_2757);
nand U12247 (N_12247,N_3823,N_1780);
or U12248 (N_12248,N_405,N_5323);
or U12249 (N_12249,N_384,N_6108);
and U12250 (N_12250,N_3228,N_2538);
or U12251 (N_12251,N_2366,N_493);
xnor U12252 (N_12252,N_5085,N_3357);
xor U12253 (N_12253,N_4753,N_150);
xnor U12254 (N_12254,N_3363,N_4472);
or U12255 (N_12255,N_2991,N_1120);
xnor U12256 (N_12256,N_1727,N_4335);
or U12257 (N_12257,N_1013,N_3287);
and U12258 (N_12258,N_398,N_1769);
and U12259 (N_12259,N_3146,N_4228);
nand U12260 (N_12260,N_2852,N_869);
nor U12261 (N_12261,N_1999,N_4348);
nor U12262 (N_12262,N_5450,N_4706);
and U12263 (N_12263,N_771,N_5213);
nor U12264 (N_12264,N_5164,N_5404);
nand U12265 (N_12265,N_1706,N_2106);
xor U12266 (N_12266,N_3526,N_845);
xor U12267 (N_12267,N_5366,N_1609);
nand U12268 (N_12268,N_3049,N_1850);
nand U12269 (N_12269,N_727,N_1389);
or U12270 (N_12270,N_6060,N_3998);
or U12271 (N_12271,N_5507,N_1519);
nor U12272 (N_12272,N_2529,N_5486);
and U12273 (N_12273,N_2957,N_2202);
and U12274 (N_12274,N_3680,N_4327);
xnor U12275 (N_12275,N_2032,N_10);
and U12276 (N_12276,N_5811,N_5810);
or U12277 (N_12277,N_1581,N_3887);
nor U12278 (N_12278,N_4011,N_1279);
nand U12279 (N_12279,N_5271,N_1428);
and U12280 (N_12280,N_5706,N_1163);
nand U12281 (N_12281,N_5399,N_3723);
xnor U12282 (N_12282,N_4809,N_112);
nand U12283 (N_12283,N_4463,N_1378);
nand U12284 (N_12284,N_4242,N_2540);
nand U12285 (N_12285,N_184,N_1889);
xor U12286 (N_12286,N_3723,N_5408);
nand U12287 (N_12287,N_1868,N_4803);
xor U12288 (N_12288,N_3500,N_6222);
nor U12289 (N_12289,N_3286,N_555);
nand U12290 (N_12290,N_4429,N_2538);
and U12291 (N_12291,N_3924,N_5317);
and U12292 (N_12292,N_1995,N_2897);
and U12293 (N_12293,N_1004,N_5932);
or U12294 (N_12294,N_3885,N_3379);
nand U12295 (N_12295,N_2592,N_1879);
xor U12296 (N_12296,N_5230,N_3080);
and U12297 (N_12297,N_3903,N_5354);
xor U12298 (N_12298,N_1581,N_1791);
and U12299 (N_12299,N_730,N_1900);
nand U12300 (N_12300,N_2033,N_2322);
or U12301 (N_12301,N_3369,N_471);
nand U12302 (N_12302,N_3379,N_4311);
xor U12303 (N_12303,N_1988,N_6062);
xor U12304 (N_12304,N_1176,N_1883);
nor U12305 (N_12305,N_4656,N_3472);
nand U12306 (N_12306,N_2854,N_594);
or U12307 (N_12307,N_5850,N_6227);
or U12308 (N_12308,N_2136,N_1888);
xnor U12309 (N_12309,N_5504,N_558);
xor U12310 (N_12310,N_5559,N_2833);
nor U12311 (N_12311,N_1514,N_460);
nor U12312 (N_12312,N_236,N_5452);
nor U12313 (N_12313,N_267,N_708);
and U12314 (N_12314,N_5394,N_3813);
and U12315 (N_12315,N_5578,N_5777);
or U12316 (N_12316,N_4578,N_1963);
xnor U12317 (N_12317,N_1932,N_663);
or U12318 (N_12318,N_3164,N_5512);
and U12319 (N_12319,N_5164,N_4968);
nor U12320 (N_12320,N_5695,N_5737);
nand U12321 (N_12321,N_5590,N_3018);
and U12322 (N_12322,N_5543,N_5330);
or U12323 (N_12323,N_2841,N_1924);
nand U12324 (N_12324,N_3672,N_5089);
nor U12325 (N_12325,N_4727,N_6016);
xor U12326 (N_12326,N_5440,N_4102);
and U12327 (N_12327,N_2135,N_1082);
or U12328 (N_12328,N_3452,N_1304);
nand U12329 (N_12329,N_1446,N_5325);
xor U12330 (N_12330,N_5396,N_4805);
nand U12331 (N_12331,N_459,N_4505);
xnor U12332 (N_12332,N_2268,N_2494);
or U12333 (N_12333,N_6197,N_1508);
nor U12334 (N_12334,N_5956,N_3028);
nor U12335 (N_12335,N_792,N_481);
xor U12336 (N_12336,N_5467,N_4844);
nand U12337 (N_12337,N_626,N_2340);
xor U12338 (N_12338,N_4750,N_4661);
and U12339 (N_12339,N_1860,N_1400);
nand U12340 (N_12340,N_2070,N_3374);
nand U12341 (N_12341,N_1662,N_5528);
xor U12342 (N_12342,N_4377,N_584);
nand U12343 (N_12343,N_2308,N_3469);
nor U12344 (N_12344,N_5953,N_3011);
and U12345 (N_12345,N_2922,N_4021);
nand U12346 (N_12346,N_1533,N_4782);
and U12347 (N_12347,N_700,N_965);
or U12348 (N_12348,N_5496,N_6002);
nor U12349 (N_12349,N_3035,N_2480);
nor U12350 (N_12350,N_4414,N_5853);
and U12351 (N_12351,N_1651,N_963);
nand U12352 (N_12352,N_431,N_2035);
nor U12353 (N_12353,N_4160,N_5956);
and U12354 (N_12354,N_2391,N_1339);
nor U12355 (N_12355,N_1930,N_2641);
or U12356 (N_12356,N_836,N_3409);
or U12357 (N_12357,N_79,N_1873);
nand U12358 (N_12358,N_1305,N_1815);
or U12359 (N_12359,N_4386,N_1865);
xor U12360 (N_12360,N_1858,N_653);
xor U12361 (N_12361,N_1970,N_6014);
nor U12362 (N_12362,N_3923,N_4723);
nand U12363 (N_12363,N_4487,N_511);
or U12364 (N_12364,N_872,N_307);
nor U12365 (N_12365,N_5198,N_1185);
and U12366 (N_12366,N_3819,N_2648);
nand U12367 (N_12367,N_2045,N_3656);
or U12368 (N_12368,N_4072,N_3223);
and U12369 (N_12369,N_4768,N_6099);
and U12370 (N_12370,N_4041,N_76);
or U12371 (N_12371,N_4139,N_828);
nand U12372 (N_12372,N_633,N_420);
and U12373 (N_12373,N_5156,N_3413);
and U12374 (N_12374,N_4181,N_4553);
nand U12375 (N_12375,N_5963,N_11);
nand U12376 (N_12376,N_5631,N_4183);
xor U12377 (N_12377,N_4667,N_5233);
and U12378 (N_12378,N_5461,N_3966);
nand U12379 (N_12379,N_95,N_5626);
xnor U12380 (N_12380,N_715,N_1806);
nand U12381 (N_12381,N_3114,N_1939);
xor U12382 (N_12382,N_1058,N_5484);
nor U12383 (N_12383,N_4794,N_711);
nor U12384 (N_12384,N_3259,N_3009);
nand U12385 (N_12385,N_5799,N_2606);
nand U12386 (N_12386,N_690,N_2586);
nor U12387 (N_12387,N_3257,N_3404);
or U12388 (N_12388,N_1898,N_3048);
and U12389 (N_12389,N_4546,N_2955);
nor U12390 (N_12390,N_2841,N_2520);
xnor U12391 (N_12391,N_4023,N_1411);
xnor U12392 (N_12392,N_5298,N_1964);
or U12393 (N_12393,N_3527,N_874);
xor U12394 (N_12394,N_2295,N_1466);
nand U12395 (N_12395,N_4723,N_3593);
or U12396 (N_12396,N_101,N_1270);
or U12397 (N_12397,N_6160,N_2371);
nand U12398 (N_12398,N_3237,N_1555);
and U12399 (N_12399,N_4187,N_5639);
or U12400 (N_12400,N_4131,N_1893);
nand U12401 (N_12401,N_1801,N_6049);
and U12402 (N_12402,N_3013,N_3643);
or U12403 (N_12403,N_5490,N_1111);
xor U12404 (N_12404,N_5853,N_5947);
nor U12405 (N_12405,N_4029,N_4831);
nand U12406 (N_12406,N_5904,N_2309);
nor U12407 (N_12407,N_2287,N_3314);
nand U12408 (N_12408,N_2607,N_196);
or U12409 (N_12409,N_3248,N_3278);
or U12410 (N_12410,N_3873,N_167);
xnor U12411 (N_12411,N_2897,N_5192);
or U12412 (N_12412,N_5118,N_941);
nand U12413 (N_12413,N_5707,N_526);
and U12414 (N_12414,N_1114,N_1417);
nor U12415 (N_12415,N_4813,N_3486);
xor U12416 (N_12416,N_5516,N_2706);
nand U12417 (N_12417,N_1920,N_1428);
nor U12418 (N_12418,N_3120,N_4643);
nand U12419 (N_12419,N_6086,N_735);
and U12420 (N_12420,N_6113,N_4944);
nor U12421 (N_12421,N_4342,N_2179);
and U12422 (N_12422,N_853,N_3029);
xor U12423 (N_12423,N_3648,N_1753);
nand U12424 (N_12424,N_2351,N_1048);
xnor U12425 (N_12425,N_2182,N_205);
and U12426 (N_12426,N_3816,N_878);
nor U12427 (N_12427,N_5992,N_3032);
and U12428 (N_12428,N_1903,N_3906);
nor U12429 (N_12429,N_4131,N_4506);
nor U12430 (N_12430,N_5768,N_1277);
xor U12431 (N_12431,N_1411,N_2753);
nand U12432 (N_12432,N_3796,N_4892);
and U12433 (N_12433,N_4013,N_3388);
or U12434 (N_12434,N_5068,N_988);
nor U12435 (N_12435,N_6179,N_2505);
and U12436 (N_12436,N_2299,N_3362);
and U12437 (N_12437,N_2959,N_2396);
xor U12438 (N_12438,N_1118,N_4678);
and U12439 (N_12439,N_1527,N_4288);
or U12440 (N_12440,N_139,N_1144);
xor U12441 (N_12441,N_4469,N_5305);
and U12442 (N_12442,N_3982,N_4669);
or U12443 (N_12443,N_1752,N_4330);
nand U12444 (N_12444,N_5071,N_3325);
and U12445 (N_12445,N_3478,N_1945);
or U12446 (N_12446,N_1842,N_5701);
xnor U12447 (N_12447,N_3649,N_542);
nand U12448 (N_12448,N_2022,N_5997);
xnor U12449 (N_12449,N_4773,N_4735);
and U12450 (N_12450,N_2578,N_1706);
nor U12451 (N_12451,N_2259,N_4780);
xnor U12452 (N_12452,N_2241,N_932);
or U12453 (N_12453,N_5734,N_4498);
xor U12454 (N_12454,N_4662,N_6192);
nor U12455 (N_12455,N_5907,N_1375);
or U12456 (N_12456,N_699,N_6164);
xor U12457 (N_12457,N_1570,N_2535);
nand U12458 (N_12458,N_5468,N_228);
nand U12459 (N_12459,N_5967,N_3527);
nor U12460 (N_12460,N_3762,N_3313);
or U12461 (N_12461,N_2455,N_4649);
nand U12462 (N_12462,N_6167,N_2757);
nand U12463 (N_12463,N_4420,N_3273);
and U12464 (N_12464,N_672,N_2397);
and U12465 (N_12465,N_2810,N_461);
and U12466 (N_12466,N_606,N_2833);
or U12467 (N_12467,N_5886,N_2561);
and U12468 (N_12468,N_4843,N_5257);
nand U12469 (N_12469,N_4801,N_871);
or U12470 (N_12470,N_5342,N_5840);
xor U12471 (N_12471,N_5311,N_217);
xnor U12472 (N_12472,N_6243,N_4646);
or U12473 (N_12473,N_3490,N_1736);
nand U12474 (N_12474,N_5979,N_4382);
and U12475 (N_12475,N_4682,N_2485);
or U12476 (N_12476,N_904,N_1356);
nand U12477 (N_12477,N_1050,N_4274);
nor U12478 (N_12478,N_1140,N_3570);
xor U12479 (N_12479,N_121,N_5170);
and U12480 (N_12480,N_3324,N_207);
xnor U12481 (N_12481,N_1598,N_2407);
nor U12482 (N_12482,N_4157,N_4374);
nand U12483 (N_12483,N_2363,N_924);
and U12484 (N_12484,N_5627,N_4609);
xor U12485 (N_12485,N_1799,N_6230);
nand U12486 (N_12486,N_3862,N_2401);
or U12487 (N_12487,N_5816,N_4151);
nor U12488 (N_12488,N_3229,N_1553);
xor U12489 (N_12489,N_552,N_1230);
nand U12490 (N_12490,N_2673,N_4262);
xor U12491 (N_12491,N_237,N_4982);
or U12492 (N_12492,N_130,N_1404);
nand U12493 (N_12493,N_20,N_6006);
xnor U12494 (N_12494,N_4888,N_1132);
or U12495 (N_12495,N_968,N_2409);
or U12496 (N_12496,N_3100,N_1552);
nor U12497 (N_12497,N_574,N_1300);
nor U12498 (N_12498,N_3592,N_6115);
xnor U12499 (N_12499,N_3840,N_4897);
xor U12500 (N_12500,N_9686,N_10676);
nand U12501 (N_12501,N_12425,N_9018);
or U12502 (N_12502,N_9043,N_8832);
nor U12503 (N_12503,N_11246,N_8263);
and U12504 (N_12504,N_6982,N_7162);
and U12505 (N_12505,N_9115,N_10421);
nand U12506 (N_12506,N_10732,N_7021);
and U12507 (N_12507,N_8445,N_9007);
nor U12508 (N_12508,N_6908,N_11829);
or U12509 (N_12509,N_11183,N_9544);
nor U12510 (N_12510,N_8635,N_10583);
or U12511 (N_12511,N_9768,N_12335);
nand U12512 (N_12512,N_8498,N_11136);
or U12513 (N_12513,N_8567,N_7845);
and U12514 (N_12514,N_10498,N_11629);
xor U12515 (N_12515,N_10920,N_8184);
nand U12516 (N_12516,N_6509,N_9934);
nand U12517 (N_12517,N_9222,N_12178);
xnor U12518 (N_12518,N_9969,N_12442);
or U12519 (N_12519,N_10212,N_11395);
or U12520 (N_12520,N_12007,N_9141);
xnor U12521 (N_12521,N_8869,N_10288);
nor U12522 (N_12522,N_12189,N_8109);
nand U12523 (N_12523,N_12325,N_6406);
and U12524 (N_12524,N_7847,N_7894);
nor U12525 (N_12525,N_10655,N_7812);
and U12526 (N_12526,N_10472,N_6827);
nor U12527 (N_12527,N_11817,N_7155);
nor U12528 (N_12528,N_10411,N_8349);
xor U12529 (N_12529,N_6878,N_12200);
nand U12530 (N_12530,N_6881,N_6634);
xnor U12531 (N_12531,N_12220,N_8959);
nor U12532 (N_12532,N_8291,N_9269);
nand U12533 (N_12533,N_10821,N_10519);
and U12534 (N_12534,N_8745,N_11156);
xor U12535 (N_12535,N_6670,N_11804);
or U12536 (N_12536,N_10773,N_6429);
xnor U12537 (N_12537,N_10559,N_12395);
nand U12538 (N_12538,N_6582,N_9539);
and U12539 (N_12539,N_11244,N_6741);
nand U12540 (N_12540,N_8592,N_6272);
or U12541 (N_12541,N_8446,N_8827);
or U12542 (N_12542,N_6382,N_9663);
or U12543 (N_12543,N_11847,N_8720);
xor U12544 (N_12544,N_7405,N_8862);
nand U12545 (N_12545,N_9498,N_10639);
and U12546 (N_12546,N_9487,N_10038);
xor U12547 (N_12547,N_6698,N_7854);
nand U12548 (N_12548,N_9084,N_12107);
nand U12549 (N_12549,N_7904,N_8489);
or U12550 (N_12550,N_7294,N_7185);
nand U12551 (N_12551,N_11686,N_9267);
nand U12552 (N_12552,N_6836,N_7417);
and U12553 (N_12553,N_6365,N_11736);
xnor U12554 (N_12554,N_7580,N_9714);
or U12555 (N_12555,N_10573,N_9514);
or U12556 (N_12556,N_7932,N_7948);
xor U12557 (N_12557,N_7280,N_9294);
nor U12558 (N_12558,N_12260,N_10343);
nor U12559 (N_12559,N_8835,N_6478);
nor U12560 (N_12560,N_8633,N_6375);
xor U12561 (N_12561,N_11441,N_11398);
nand U12562 (N_12562,N_6685,N_8554);
nand U12563 (N_12563,N_7484,N_6469);
nand U12564 (N_12564,N_11692,N_10048);
nor U12565 (N_12565,N_10495,N_9656);
nand U12566 (N_12566,N_6867,N_10911);
nor U12567 (N_12567,N_7397,N_10678);
xor U12568 (N_12568,N_7382,N_8629);
and U12569 (N_12569,N_9235,N_10935);
xor U12570 (N_12570,N_8262,N_11981);
and U12571 (N_12571,N_7131,N_12142);
nor U12572 (N_12572,N_8158,N_9467);
or U12573 (N_12573,N_6734,N_10784);
nand U12574 (N_12574,N_7446,N_6435);
or U12575 (N_12575,N_8575,N_7342);
nor U12576 (N_12576,N_6477,N_9098);
or U12577 (N_12577,N_10051,N_12330);
xor U12578 (N_12578,N_9622,N_9310);
nor U12579 (N_12579,N_7698,N_10005);
nor U12580 (N_12580,N_11864,N_7217);
nor U12581 (N_12581,N_10841,N_8630);
nand U12582 (N_12582,N_7331,N_11207);
xor U12583 (N_12583,N_7369,N_9633);
nand U12584 (N_12584,N_6453,N_7514);
or U12585 (N_12585,N_8686,N_6749);
nor U12586 (N_12586,N_6797,N_6804);
and U12587 (N_12587,N_11260,N_10582);
or U12588 (N_12588,N_6377,N_8218);
xor U12589 (N_12589,N_9326,N_11780);
xor U12590 (N_12590,N_7154,N_12285);
nor U12591 (N_12591,N_9315,N_7090);
nor U12592 (N_12592,N_11234,N_8643);
nand U12593 (N_12593,N_7093,N_6779);
or U12594 (N_12594,N_11946,N_8607);
or U12595 (N_12595,N_8905,N_9480);
xor U12596 (N_12596,N_10645,N_12493);
or U12597 (N_12597,N_6679,N_7241);
or U12598 (N_12598,N_7588,N_11514);
and U12599 (N_12599,N_7936,N_8766);
nand U12600 (N_12600,N_7767,N_11184);
or U12601 (N_12601,N_10646,N_10301);
nand U12602 (N_12602,N_8357,N_6673);
xnor U12603 (N_12603,N_11676,N_10396);
nand U12604 (N_12604,N_9057,N_11811);
and U12605 (N_12605,N_8809,N_8235);
and U12606 (N_12606,N_7960,N_10834);
xnor U12607 (N_12607,N_12246,N_10752);
and U12608 (N_12608,N_6364,N_11525);
or U12609 (N_12609,N_9575,N_10529);
nand U12610 (N_12610,N_7994,N_12129);
and U12611 (N_12611,N_9028,N_12472);
or U12612 (N_12612,N_8776,N_11285);
nand U12613 (N_12613,N_8361,N_10838);
nand U12614 (N_12614,N_9702,N_9876);
and U12615 (N_12615,N_6960,N_11650);
nand U12616 (N_12616,N_8781,N_10158);
nand U12617 (N_12617,N_6636,N_10159);
and U12618 (N_12618,N_9767,N_8464);
nand U12619 (N_12619,N_10137,N_10316);
or U12620 (N_12620,N_10563,N_7365);
or U12621 (N_12621,N_9662,N_8042);
nor U12622 (N_12622,N_10609,N_7554);
xnor U12623 (N_12623,N_11769,N_9674);
and U12624 (N_12624,N_7631,N_7308);
or U12625 (N_12625,N_8564,N_8694);
and U12626 (N_12626,N_8719,N_8267);
or U12627 (N_12627,N_6274,N_8674);
xnor U12628 (N_12628,N_8988,N_11017);
nand U12629 (N_12629,N_12413,N_10749);
nor U12630 (N_12630,N_7489,N_10807);
nand U12631 (N_12631,N_11434,N_7575);
and U12632 (N_12632,N_12070,N_8196);
xnor U12633 (N_12633,N_11296,N_11595);
nand U12634 (N_12634,N_7065,N_10763);
nand U12635 (N_12635,N_10263,N_8849);
or U12636 (N_12636,N_8825,N_11520);
nor U12637 (N_12637,N_11265,N_6403);
nor U12638 (N_12638,N_10871,N_11245);
nand U12639 (N_12639,N_7597,N_9274);
or U12640 (N_12640,N_12205,N_8691);
and U12641 (N_12641,N_10647,N_9629);
or U12642 (N_12642,N_7766,N_10085);
nand U12643 (N_12643,N_8769,N_9220);
nand U12644 (N_12644,N_10877,N_9064);
or U12645 (N_12645,N_11367,N_8282);
or U12646 (N_12646,N_11497,N_11490);
and U12647 (N_12647,N_9855,N_8363);
xnor U12648 (N_12648,N_9446,N_12323);
nor U12649 (N_12649,N_9939,N_9229);
nand U12650 (N_12650,N_7047,N_10750);
or U12651 (N_12651,N_8797,N_10248);
and U12652 (N_12652,N_11733,N_9857);
and U12653 (N_12653,N_7205,N_7800);
nand U12654 (N_12654,N_11097,N_12296);
or U12655 (N_12655,N_12455,N_6830);
xnor U12656 (N_12656,N_7385,N_9762);
nor U12657 (N_12657,N_6424,N_10754);
nor U12658 (N_12658,N_9021,N_9212);
nor U12659 (N_12659,N_9973,N_10814);
nand U12660 (N_12660,N_10412,N_8442);
nor U12661 (N_12661,N_10228,N_12033);
and U12662 (N_12662,N_8568,N_11799);
nor U12663 (N_12663,N_9193,N_9343);
xor U12664 (N_12664,N_7106,N_6610);
nand U12665 (N_12665,N_8022,N_11626);
and U12666 (N_12666,N_11500,N_10990);
and U12667 (N_12667,N_10889,N_7248);
xor U12668 (N_12668,N_9036,N_12376);
and U12669 (N_12669,N_9799,N_10103);
or U12670 (N_12670,N_12418,N_10059);
xor U12671 (N_12671,N_10695,N_11982);
xnor U12672 (N_12672,N_10973,N_9053);
or U12673 (N_12673,N_7692,N_11222);
nand U12674 (N_12674,N_9887,N_8013);
or U12675 (N_12675,N_11341,N_11975);
nand U12676 (N_12676,N_12240,N_10507);
and U12677 (N_12677,N_11945,N_11484);
or U12678 (N_12678,N_12417,N_9667);
or U12679 (N_12679,N_12021,N_9779);
nand U12680 (N_12680,N_11415,N_7873);
nand U12681 (N_12681,N_10648,N_12406);
nand U12682 (N_12682,N_9199,N_9351);
nor U12683 (N_12683,N_9687,N_8093);
nand U12684 (N_12684,N_10312,N_7105);
or U12685 (N_12685,N_6680,N_8283);
nand U12686 (N_12686,N_8049,N_11916);
xor U12687 (N_12687,N_10672,N_6397);
nand U12688 (N_12688,N_8402,N_12256);
or U12689 (N_12689,N_8947,N_8579);
or U12690 (N_12690,N_6566,N_7302);
nand U12691 (N_12691,N_9417,N_6289);
xnor U12692 (N_12692,N_7718,N_7410);
xnor U12693 (N_12693,N_7978,N_8495);
nand U12694 (N_12694,N_9037,N_11448);
nand U12695 (N_12695,N_6853,N_8838);
nor U12696 (N_12696,N_7035,N_7350);
or U12697 (N_12697,N_8562,N_9150);
xor U12698 (N_12698,N_7899,N_7291);
nor U12699 (N_12699,N_8886,N_10456);
or U12700 (N_12700,N_10400,N_10196);
and U12701 (N_12701,N_9104,N_7952);
or U12702 (N_12702,N_10241,N_6912);
nand U12703 (N_12703,N_10951,N_7616);
nand U12704 (N_12704,N_9706,N_9119);
nor U12705 (N_12705,N_11897,N_8191);
nand U12706 (N_12706,N_6690,N_9995);
or U12707 (N_12707,N_9355,N_10413);
nor U12708 (N_12708,N_11475,N_12036);
or U12709 (N_12709,N_10977,N_7149);
nand U12710 (N_12710,N_8364,N_12268);
nor U12711 (N_12711,N_12227,N_11647);
xor U12712 (N_12712,N_6941,N_6413);
and U12713 (N_12713,N_10824,N_10466);
nor U12714 (N_12714,N_6884,N_12232);
xnor U12715 (N_12715,N_6258,N_10922);
and U12716 (N_12716,N_9012,N_8255);
nand U12717 (N_12717,N_11277,N_7166);
nor U12718 (N_12718,N_9170,N_6452);
xor U12719 (N_12719,N_7088,N_6824);
nor U12720 (N_12720,N_8619,N_12423);
xor U12721 (N_12721,N_9410,N_10937);
nor U12722 (N_12722,N_10178,N_10450);
or U12723 (N_12723,N_6931,N_8612);
or U12724 (N_12724,N_8517,N_11027);
xor U12725 (N_12725,N_9972,N_7303);
xor U12726 (N_12726,N_11024,N_6711);
nand U12727 (N_12727,N_10641,N_7051);
nand U12728 (N_12728,N_11710,N_6611);
nor U12729 (N_12729,N_12103,N_6992);
nor U12730 (N_12730,N_12080,N_10964);
and U12731 (N_12731,N_7375,N_8974);
nand U12732 (N_12732,N_7234,N_7925);
nand U12733 (N_12733,N_6745,N_8165);
nand U12734 (N_12734,N_10933,N_6727);
or U12735 (N_12735,N_11918,N_6456);
nor U12736 (N_12736,N_7829,N_7057);
nand U12737 (N_12737,N_7286,N_10029);
nand U12738 (N_12738,N_10697,N_6756);
and U12739 (N_12739,N_9694,N_8439);
or U12740 (N_12740,N_8006,N_10723);
xor U12741 (N_12741,N_10293,N_8840);
or U12742 (N_12742,N_9591,N_10362);
and U12743 (N_12743,N_7409,N_10168);
nor U12744 (N_12744,N_11549,N_12102);
xnor U12745 (N_12745,N_9904,N_9808);
nor U12746 (N_12746,N_7190,N_6539);
and U12747 (N_12747,N_9769,N_8546);
or U12748 (N_12748,N_11917,N_8377);
xor U12749 (N_12749,N_6526,N_9834);
xnor U12750 (N_12750,N_12464,N_6291);
and U12751 (N_12751,N_9618,N_11488);
xor U12752 (N_12752,N_9962,N_8750);
or U12753 (N_12753,N_11262,N_8278);
nor U12754 (N_12754,N_7493,N_8395);
and U12755 (N_12755,N_8756,N_7858);
nand U12756 (N_12756,N_8707,N_10200);
nor U12757 (N_12757,N_11194,N_11286);
nand U12758 (N_12758,N_9565,N_10332);
or U12759 (N_12759,N_8659,N_11288);
nor U12760 (N_12760,N_9283,N_6313);
xnor U12761 (N_12761,N_11414,N_6296);
xor U12762 (N_12762,N_6772,N_7170);
xnor U12763 (N_12763,N_12286,N_8984);
nor U12764 (N_12764,N_11450,N_8742);
xnor U12765 (N_12765,N_8167,N_11170);
nor U12766 (N_12766,N_9951,N_10128);
or U12767 (N_12767,N_8520,N_10260);
nand U12768 (N_12768,N_12072,N_11826);
xnor U12769 (N_12769,N_8468,N_11088);
xnor U12770 (N_12770,N_10356,N_11747);
or U12771 (N_12771,N_6370,N_11369);
xnor U12772 (N_12772,N_10094,N_10330);
and U12773 (N_12773,N_7797,N_10976);
nand U12774 (N_12774,N_8941,N_7662);
nand U12775 (N_12775,N_11028,N_10170);
nor U12776 (N_12776,N_7485,N_10827);
or U12777 (N_12777,N_11612,N_9206);
xnor U12778 (N_12778,N_9987,N_10189);
xnor U12779 (N_12779,N_9583,N_10165);
xnor U12780 (N_12780,N_9158,N_11791);
and U12781 (N_12781,N_11540,N_9493);
nand U12782 (N_12782,N_8189,N_7212);
and U12783 (N_12783,N_9841,N_9554);
xor U12784 (N_12784,N_10437,N_9682);
nand U12785 (N_12785,N_11870,N_6668);
or U12786 (N_12786,N_10809,N_8640);
nor U12787 (N_12787,N_6737,N_8116);
nor U12788 (N_12788,N_7715,N_11765);
nor U12789 (N_12789,N_7956,N_12393);
xor U12790 (N_12790,N_9318,N_11180);
nor U12791 (N_12791,N_7523,N_8038);
xnor U12792 (N_12792,N_8256,N_7543);
nand U12793 (N_12793,N_8565,N_10138);
or U12794 (N_12794,N_7884,N_8356);
xnor U12795 (N_12795,N_10032,N_7566);
and U12796 (N_12796,N_11951,N_11345);
nand U12797 (N_12797,N_6683,N_6973);
xor U12798 (N_12798,N_10016,N_6844);
nand U12799 (N_12799,N_9996,N_9704);
nor U12800 (N_12800,N_10524,N_9536);
nand U12801 (N_12801,N_8807,N_12125);
and U12802 (N_12802,N_9932,N_7230);
xnor U12803 (N_12803,N_12071,N_12404);
nand U12804 (N_12804,N_10984,N_9558);
xnor U12805 (N_12805,N_11397,N_8681);
xor U12806 (N_12806,N_11958,N_10543);
nor U12807 (N_12807,N_10436,N_8700);
nand U12808 (N_12808,N_6788,N_10802);
or U12809 (N_12809,N_7657,N_9162);
or U12810 (N_12810,N_9907,N_6280);
and U12811 (N_12811,N_11904,N_8104);
or U12812 (N_12812,N_9650,N_7279);
or U12813 (N_12813,N_7137,N_11760);
and U12814 (N_12814,N_12462,N_6856);
xor U12815 (N_12815,N_11637,N_8508);
and U12816 (N_12816,N_6691,N_11089);
nand U12817 (N_12817,N_9407,N_9336);
and U12818 (N_12818,N_8340,N_11995);
or U12819 (N_12819,N_11730,N_8272);
or U12820 (N_12820,N_8563,N_6650);
nand U12821 (N_12821,N_9548,N_6495);
xnor U12822 (N_12822,N_10477,N_10216);
and U12823 (N_12823,N_10021,N_8025);
and U12824 (N_12824,N_8952,N_6874);
and U12825 (N_12825,N_9872,N_7503);
xor U12826 (N_12826,N_11485,N_10186);
nand U12827 (N_12827,N_11299,N_8755);
xor U12828 (N_12828,N_6842,N_11197);
nor U12829 (N_12829,N_10699,N_9709);
xnor U12830 (N_12830,N_7240,N_8246);
nand U12831 (N_12831,N_9450,N_10596);
nand U12832 (N_12832,N_9810,N_8779);
xnor U12833 (N_12833,N_11346,N_7272);
nand U12834 (N_12834,N_9495,N_10464);
or U12835 (N_12835,N_9384,N_6502);
nor U12836 (N_12836,N_9088,N_7896);
or U12837 (N_12837,N_9676,N_10360);
and U12838 (N_12838,N_7686,N_8066);
and U12839 (N_12839,N_9496,N_9572);
nand U12840 (N_12840,N_11214,N_10331);
xnor U12841 (N_12841,N_12274,N_10694);
and U12842 (N_12842,N_6340,N_9010);
and U12843 (N_12843,N_7706,N_6308);
xnor U12844 (N_12844,N_12495,N_11573);
and U12845 (N_12845,N_11060,N_12075);
or U12846 (N_12846,N_11147,N_11304);
or U12847 (N_12847,N_9794,N_10275);
xnor U12848 (N_12848,N_8033,N_6773);
and U12849 (N_12849,N_6480,N_12380);
and U12850 (N_12850,N_7680,N_7578);
or U12851 (N_12851,N_8185,N_7096);
nand U12852 (N_12852,N_6883,N_6927);
nor U12853 (N_12853,N_12491,N_10551);
and U12854 (N_12854,N_8726,N_11314);
xnor U12855 (N_12855,N_9047,N_6431);
and U12856 (N_12856,N_8311,N_12115);
nor U12857 (N_12857,N_6288,N_8505);
or U12858 (N_12858,N_12299,N_10446);
or U12859 (N_12859,N_9713,N_9801);
nor U12860 (N_12860,N_9268,N_12241);
or U12861 (N_12861,N_8928,N_7512);
or U12862 (N_12862,N_11396,N_7458);
xnor U12863 (N_12863,N_7796,N_10790);
and U12864 (N_12864,N_12447,N_10082);
and U12865 (N_12865,N_6360,N_7132);
nor U12866 (N_12866,N_11287,N_8581);
nor U12867 (N_12867,N_9105,N_8039);
nand U12868 (N_12868,N_11332,N_8799);
nand U12869 (N_12869,N_10409,N_10358);
and U12870 (N_12870,N_8011,N_8697);
or U12871 (N_12871,N_10395,N_7322);
nor U12872 (N_12872,N_7822,N_11495);
or U12873 (N_12873,N_8456,N_9491);
or U12874 (N_12874,N_8626,N_8310);
or U12875 (N_12875,N_6472,N_10355);
nor U12876 (N_12876,N_10095,N_8326);
or U12877 (N_12877,N_7231,N_12377);
or U12878 (N_12878,N_7102,N_9559);
nand U12879 (N_12879,N_7262,N_10506);
nor U12880 (N_12880,N_10910,N_8435);
xor U12881 (N_12881,N_8761,N_9231);
xor U12882 (N_12882,N_11627,N_7610);
or U12883 (N_12883,N_11057,N_6279);
and U12884 (N_12884,N_9168,N_9254);
nor U12885 (N_12885,N_10879,N_9439);
or U12886 (N_12886,N_8919,N_6860);
nand U12887 (N_12887,N_7659,N_7592);
nor U12888 (N_12888,N_8739,N_11825);
xor U12889 (N_12889,N_10187,N_12186);
xnor U12890 (N_12890,N_11135,N_6765);
and U12891 (N_12891,N_12153,N_12093);
nor U12892 (N_12892,N_9014,N_6389);
or U12893 (N_12893,N_11546,N_12052);
xor U12894 (N_12894,N_11478,N_7050);
and U12895 (N_12895,N_10420,N_9073);
nand U12896 (N_12896,N_7844,N_12426);
xnor U12897 (N_12897,N_10020,N_10025);
and U12898 (N_12898,N_11401,N_9649);
and U12899 (N_12899,N_7900,N_6644);
nor U12900 (N_12900,N_8767,N_9066);
xor U12901 (N_12901,N_6770,N_10220);
xnor U12902 (N_12902,N_8161,N_11023);
nor U12903 (N_12903,N_11357,N_9230);
xor U12904 (N_12904,N_9752,N_12421);
and U12905 (N_12905,N_6961,N_10885);
and U12906 (N_12906,N_7219,N_8083);
or U12907 (N_12907,N_10592,N_6843);
nand U12908 (N_12908,N_6705,N_12044);
or U12909 (N_12909,N_11376,N_6387);
and U12910 (N_12910,N_10338,N_8155);
or U12911 (N_12911,N_8031,N_8589);
nand U12912 (N_12912,N_9325,N_8091);
xnor U12913 (N_12913,N_8450,N_12234);
or U12914 (N_12914,N_7196,N_12130);
xnor U12915 (N_12915,N_6421,N_11402);
and U12916 (N_12916,N_7573,N_9870);
nor U12917 (N_12917,N_11782,N_8064);
nor U12918 (N_12918,N_7368,N_8077);
nor U12919 (N_12919,N_6731,N_10649);
xnor U12920 (N_12920,N_9469,N_9606);
and U12921 (N_12921,N_9822,N_11935);
xor U12922 (N_12922,N_8899,N_7762);
and U12923 (N_12923,N_9525,N_11235);
nand U12924 (N_12924,N_7653,N_6868);
nor U12925 (N_12925,N_7336,N_9090);
nor U12926 (N_12926,N_12489,N_11436);
xnor U12927 (N_12927,N_7747,N_10224);
or U12928 (N_12928,N_9929,N_12144);
xnor U12929 (N_12929,N_6753,N_10387);
xor U12930 (N_12930,N_9397,N_8693);
xnor U12931 (N_12931,N_7491,N_11099);
xor U12932 (N_12932,N_10971,N_7957);
nand U12933 (N_12933,N_8534,N_10927);
and U12934 (N_12934,N_8647,N_8580);
and U12935 (N_12935,N_6807,N_9152);
nor U12936 (N_12936,N_12438,N_8156);
and U12937 (N_12937,N_12067,N_8783);
and U12938 (N_12938,N_7235,N_10550);
xnor U12939 (N_12939,N_10939,N_12212);
nand U12940 (N_12940,N_6969,N_7816);
xnor U12941 (N_12941,N_11077,N_7069);
nor U12942 (N_12942,N_6800,N_6740);
nor U12943 (N_12943,N_12336,N_9427);
nand U12944 (N_12944,N_11542,N_10193);
nand U12945 (N_12945,N_11326,N_7676);
nor U12946 (N_12946,N_7346,N_9197);
nor U12947 (N_12947,N_11474,N_10003);
and U12948 (N_12948,N_11157,N_9052);
and U12949 (N_12949,N_8405,N_6864);
nand U12950 (N_12950,N_8611,N_10126);
or U12951 (N_12951,N_7656,N_12313);
and U12952 (N_12952,N_6544,N_10535);
nor U12953 (N_12953,N_10418,N_10610);
or U12954 (N_12954,N_8614,N_7700);
nor U12955 (N_12955,N_7638,N_9700);
nand U12956 (N_12956,N_8316,N_11698);
or U12957 (N_12957,N_7769,N_11822);
and U12958 (N_12958,N_7674,N_11081);
nand U12959 (N_12959,N_10390,N_9748);
or U12960 (N_12960,N_7856,N_8142);
or U12961 (N_12961,N_10426,N_10523);
xnor U12962 (N_12962,N_8012,N_7004);
nand U12963 (N_12963,N_10903,N_9499);
nand U12964 (N_12964,N_9905,N_10268);
and U12965 (N_12965,N_7753,N_8058);
and U12966 (N_12966,N_6651,N_8902);
nor U12967 (N_12967,N_6767,N_7483);
xor U12968 (N_12968,N_9476,N_11227);
or U12969 (N_12969,N_9941,N_9344);
or U12970 (N_12970,N_8560,N_9042);
xor U12971 (N_12971,N_10736,N_6825);
and U12972 (N_12972,N_8199,N_8863);
nand U12973 (N_12973,N_6932,N_9542);
or U12974 (N_12974,N_10876,N_11554);
xor U12975 (N_12975,N_7617,N_11164);
and U12976 (N_12976,N_11226,N_10063);
nand U12977 (N_12977,N_6338,N_10629);
or U12978 (N_12978,N_8458,N_6632);
xor U12979 (N_12979,N_8063,N_6260);
nor U12980 (N_12980,N_7545,N_10148);
nand U12981 (N_12981,N_6631,N_7049);
and U12982 (N_12982,N_7252,N_7064);
nor U12983 (N_12983,N_6505,N_9011);
xnor U12984 (N_12984,N_10467,N_9204);
xnor U12985 (N_12985,N_6870,N_12085);
or U12986 (N_12986,N_10375,N_7407);
nand U12987 (N_12987,N_9298,N_10452);
or U12988 (N_12988,N_9160,N_9695);
or U12989 (N_12989,N_9297,N_11219);
and U12990 (N_12990,N_8639,N_10757);
nor U12991 (N_12991,N_10869,N_10053);
xor U12992 (N_12992,N_8574,N_7508);
or U12993 (N_12993,N_10227,N_10213);
or U12994 (N_12994,N_10240,N_8129);
xor U12995 (N_12995,N_10846,N_12430);
or U12996 (N_12996,N_8714,N_11842);
nand U12997 (N_12997,N_10547,N_9167);
and U12998 (N_12998,N_9711,N_8898);
xnor U12999 (N_12999,N_9081,N_12182);
nand U13000 (N_13000,N_10961,N_9359);
and U13001 (N_13001,N_9054,N_11877);
xnor U13002 (N_13002,N_10104,N_11863);
xor U13003 (N_13003,N_11741,N_11026);
or U13004 (N_13004,N_7323,N_10010);
and U13005 (N_13005,N_12100,N_6709);
nor U13006 (N_13006,N_6263,N_6445);
and U13007 (N_13007,N_12319,N_11766);
nor U13008 (N_13008,N_11708,N_11608);
and U13009 (N_13009,N_6298,N_9085);
xor U13010 (N_13010,N_12089,N_11233);
nor U13011 (N_13011,N_8906,N_10576);
nand U13012 (N_13012,N_9665,N_10001);
and U13013 (N_13013,N_11014,N_11320);
or U13014 (N_13014,N_11854,N_7371);
xnor U13015 (N_13015,N_8771,N_7157);
nand U13016 (N_13016,N_11310,N_11015);
or U13017 (N_13017,N_12190,N_7129);
nor U13018 (N_13018,N_8623,N_10662);
nand U13019 (N_13019,N_9993,N_10236);
nand U13020 (N_13020,N_11137,N_6750);
nand U13021 (N_13021,N_10110,N_11366);
nand U13022 (N_13022,N_8644,N_6593);
nor U13023 (N_13023,N_10781,N_8017);
and U13024 (N_13024,N_7220,N_11643);
nand U13025 (N_13025,N_7445,N_9418);
xor U13026 (N_13026,N_6427,N_10665);
nand U13027 (N_13027,N_7953,N_6527);
nand U13028 (N_13028,N_8523,N_11211);
and U13029 (N_13029,N_6717,N_9096);
nand U13030 (N_13030,N_9648,N_7029);
or U13031 (N_13031,N_11289,N_8319);
or U13032 (N_13032,N_12357,N_6774);
and U13033 (N_13033,N_10287,N_9845);
or U13034 (N_13034,N_9002,N_9940);
nand U13035 (N_13035,N_12217,N_6682);
and U13036 (N_13036,N_10011,N_7919);
nand U13037 (N_13037,N_8106,N_11221);
nand U13038 (N_13038,N_11171,N_11681);
or U13039 (N_13039,N_8350,N_8015);
xor U13040 (N_13040,N_7224,N_7255);
xor U13041 (N_13041,N_8500,N_7831);
and U13042 (N_13042,N_10344,N_9025);
and U13043 (N_13043,N_11303,N_10735);
nor U13044 (N_13044,N_7040,N_10518);
xnor U13045 (N_13045,N_7067,N_9376);
nand U13046 (N_13046,N_7347,N_11002);
nor U13047 (N_13047,N_10217,N_12134);
or U13048 (N_13048,N_10677,N_9227);
or U13049 (N_13049,N_9116,N_10620);
xor U13050 (N_13050,N_11128,N_10710);
and U13051 (N_13051,N_10232,N_10147);
xnor U13052 (N_13052,N_6879,N_11054);
and U13053 (N_13053,N_12219,N_7383);
and U13054 (N_13054,N_8774,N_8194);
nand U13055 (N_13055,N_9597,N_11921);
nor U13056 (N_13056,N_11667,N_7533);
or U13057 (N_13057,N_7703,N_11740);
or U13058 (N_13058,N_7713,N_10096);
nand U13059 (N_13059,N_8415,N_8335);
or U13060 (N_13060,N_12174,N_12229);
xor U13061 (N_13061,N_10372,N_8951);
or U13062 (N_13062,N_9412,N_6620);
nor U13063 (N_13063,N_7879,N_9251);
and U13064 (N_13064,N_7540,N_11115);
xor U13065 (N_13065,N_8045,N_6760);
xnor U13066 (N_13066,N_7661,N_10720);
nor U13067 (N_13067,N_7734,N_9612);
nor U13068 (N_13068,N_11756,N_9807);
nand U13069 (N_13069,N_10404,N_11984);
nor U13070 (N_13070,N_7804,N_10759);
and U13071 (N_13071,N_6963,N_12370);
or U13072 (N_13072,N_9209,N_11548);
nor U13073 (N_13073,N_11122,N_7835);
nand U13074 (N_13074,N_10009,N_10278);
and U13075 (N_13075,N_7848,N_7202);
and U13076 (N_13076,N_8741,N_10361);
xnor U13077 (N_13077,N_9576,N_7513);
or U13078 (N_13078,N_7920,N_7292);
xor U13079 (N_13079,N_11291,N_9272);
or U13080 (N_13080,N_6589,N_7825);
nand U13081 (N_13081,N_10603,N_8309);
xnor U13082 (N_13082,N_10658,N_9839);
and U13083 (N_13083,N_12249,N_8971);
xor U13084 (N_13084,N_7889,N_8469);
or U13085 (N_13085,N_8108,N_11899);
and U13086 (N_13086,N_12356,N_12046);
and U13087 (N_13087,N_10786,N_11487);
nand U13088 (N_13088,N_7515,N_10965);
or U13089 (N_13089,N_10915,N_11315);
and U13090 (N_13090,N_8847,N_7477);
or U13091 (N_13091,N_7501,N_10865);
xor U13092 (N_13092,N_9239,N_7167);
or U13093 (N_13093,N_8918,N_9208);
nor U13094 (N_13094,N_8699,N_6766);
or U13095 (N_13095,N_6599,N_7642);
nand U13096 (N_13096,N_8670,N_10496);
and U13097 (N_13097,N_9317,N_11579);
nand U13098 (N_13098,N_6901,N_8656);
or U13099 (N_13099,N_9745,N_7949);
xnor U13100 (N_13100,N_11435,N_11693);
xnor U13101 (N_13101,N_12269,N_10040);
or U13102 (N_13102,N_6575,N_9477);
and U13103 (N_13103,N_9999,N_7435);
nand U13104 (N_13104,N_8385,N_10812);
xor U13105 (N_13105,N_6396,N_11439);
nor U13106 (N_13106,N_9411,N_7263);
and U13107 (N_13107,N_9792,N_8970);
and U13108 (N_13108,N_8355,N_7763);
nand U13109 (N_13109,N_10042,N_11584);
nand U13110 (N_13110,N_9092,N_9615);
xnor U13111 (N_13111,N_8099,N_7095);
or U13112 (N_13112,N_11205,N_9257);
and U13113 (N_13113,N_8880,N_11449);
xnor U13114 (N_13114,N_9500,N_11634);
nand U13115 (N_13115,N_11068,N_7637);
nor U13116 (N_13116,N_10948,N_7118);
and U13117 (N_13117,N_7386,N_7901);
or U13118 (N_13118,N_9775,N_7670);
xnor U13119 (N_13119,N_10315,N_6987);
nor U13120 (N_13120,N_10666,N_11848);
xor U13121 (N_13121,N_6646,N_10851);
and U13122 (N_13122,N_10221,N_11592);
xnor U13123 (N_13123,N_10870,N_10605);
nor U13124 (N_13124,N_11102,N_7681);
nand U13125 (N_13125,N_10257,N_6565);
or U13126 (N_13126,N_10602,N_12231);
nand U13127 (N_13127,N_6314,N_11350);
xnor U13128 (N_13128,N_10256,N_12277);
nand U13129 (N_13129,N_7549,N_8328);
xnor U13130 (N_13130,N_12222,N_9849);
xnor U13131 (N_13131,N_8958,N_9144);
nor U13132 (N_13132,N_6633,N_7984);
or U13133 (N_13133,N_9858,N_8048);
nor U13134 (N_13134,N_11890,N_10680);
or U13135 (N_13135,N_10223,N_6557);
xnor U13136 (N_13136,N_10124,N_8926);
or U13137 (N_13137,N_6508,N_9473);
or U13138 (N_13138,N_11901,N_8532);
nor U13139 (N_13139,N_12402,N_10843);
nor U13140 (N_13140,N_8453,N_7687);
nor U13141 (N_13141,N_12443,N_6306);
nor U13142 (N_13142,N_8922,N_8678);
xnor U13143 (N_13143,N_11294,N_7787);
xor U13144 (N_13144,N_11787,N_9866);
xor U13145 (N_13145,N_7705,N_8923);
or U13146 (N_13146,N_7227,N_11888);
xor U13147 (N_13147,N_9584,N_11220);
nand U13148 (N_13148,N_8181,N_7551);
and U13149 (N_13149,N_6483,N_8945);
or U13150 (N_13150,N_10785,N_7062);
and U13151 (N_13151,N_10743,N_10219);
xnor U13152 (N_13152,N_8131,N_9482);
or U13153 (N_13153,N_9820,N_12312);
or U13154 (N_13154,N_9520,N_9225);
and U13155 (N_13155,N_8482,N_12251);
nand U13156 (N_13156,N_7644,N_11114);
xor U13157 (N_13157,N_6820,N_7720);
and U13158 (N_13158,N_8519,N_10584);
nor U13159 (N_13159,N_11202,N_11508);
and U13160 (N_13160,N_9369,N_10341);
xor U13161 (N_13161,N_8462,N_11705);
xor U13162 (N_13162,N_7817,N_7649);
or U13163 (N_13163,N_9830,N_7208);
nand U13164 (N_13164,N_12106,N_8228);
xor U13165 (N_13165,N_7296,N_10099);
and U13166 (N_13166,N_11132,N_8541);
xor U13167 (N_13167,N_10511,N_6922);
and U13168 (N_13168,N_9139,N_7404);
nand U13169 (N_13169,N_11695,N_9620);
or U13170 (N_13170,N_9955,N_8530);
and U13171 (N_13171,N_11066,N_7834);
xnor U13172 (N_13172,N_7793,N_7140);
xor U13173 (N_13173,N_11506,N_9579);
xnor U13174 (N_13174,N_10631,N_7909);
or U13175 (N_13175,N_7906,N_8891);
nor U13176 (N_13176,N_6335,N_9644);
or U13177 (N_13177,N_11044,N_11639);
and U13178 (N_13178,N_8288,N_11714);
or U13179 (N_13179,N_9488,N_8730);
nand U13180 (N_13180,N_6798,N_11313);
nand U13181 (N_13181,N_6547,N_8577);
xnor U13182 (N_13182,N_10914,N_6341);
xnor U13183 (N_13183,N_10345,N_10816);
or U13184 (N_13184,N_8230,N_6639);
and U13185 (N_13185,N_6905,N_8538);
or U13186 (N_13186,N_8831,N_6748);
or U13187 (N_13187,N_6970,N_6357);
xnor U13188 (N_13188,N_9937,N_11581);
xor U13189 (N_13189,N_10703,N_10724);
or U13190 (N_13190,N_12487,N_9363);
nor U13191 (N_13191,N_7063,N_9191);
or U13192 (N_13192,N_8650,N_8392);
and U13193 (N_13193,N_7560,N_10210);
or U13194 (N_13194,N_6533,N_11290);
and U13195 (N_13195,N_6819,N_12304);
and U13196 (N_13196,N_9848,N_12478);
and U13197 (N_13197,N_7288,N_12169);
or U13198 (N_13198,N_12209,N_7012);
nor U13199 (N_13199,N_7546,N_7223);
nand U13200 (N_13200,N_12154,N_6408);
and U13201 (N_13201,N_8298,N_11726);
nand U13202 (N_13202,N_7784,N_10726);
or U13203 (N_13203,N_8821,N_8005);
nor U13204 (N_13204,N_9432,N_12162);
nand U13205 (N_13205,N_6513,N_10394);
and U13206 (N_13206,N_11091,N_6626);
or U13207 (N_13207,N_9390,N_8695);
or U13208 (N_13208,N_9724,N_8372);
and U13209 (N_13209,N_7635,N_6346);
xor U13210 (N_13210,N_9192,N_6716);
xnor U13211 (N_13211,N_10117,N_6956);
or U13212 (N_13212,N_10064,N_12244);
nand U13213 (N_13213,N_11431,N_9282);
xor U13214 (N_13214,N_6928,N_11344);
nor U13215 (N_13215,N_7811,N_12081);
and U13216 (N_13216,N_7039,N_11472);
xor U13217 (N_13217,N_7997,N_11539);
and U13218 (N_13218,N_10424,N_8127);
and U13219 (N_13219,N_8599,N_10753);
nor U13220 (N_13220,N_11481,N_6838);
and U13221 (N_13221,N_8086,N_9688);
nand U13222 (N_13222,N_8909,N_10987);
and U13223 (N_13223,N_10577,N_10708);
nor U13224 (N_13224,N_10149,N_10253);
nand U13225 (N_13225,N_11104,N_11513);
nor U13226 (N_13226,N_7995,N_8222);
or U13227 (N_13227,N_11352,N_7916);
nor U13228 (N_13228,N_12345,N_10113);
nor U13229 (N_13229,N_9114,N_9234);
or U13230 (N_13230,N_11618,N_11820);
nand U13231 (N_13231,N_9502,N_8657);
nand U13232 (N_13232,N_8864,N_9639);
xor U13233 (N_13233,N_9302,N_6738);
or U13234 (N_13234,N_10866,N_11343);
and U13235 (N_13235,N_12090,N_11691);
nor U13236 (N_13236,N_11809,N_7521);
xor U13237 (N_13237,N_11492,N_10244);
xnor U13238 (N_13238,N_8729,N_9777);
nand U13239 (N_13239,N_12032,N_6271);
and U13240 (N_13240,N_8164,N_12394);
nor U13241 (N_13241,N_9421,N_7466);
and U13242 (N_13242,N_8930,N_10060);
and U13243 (N_13243,N_9529,N_7277);
nor U13244 (N_13244,N_11893,N_7524);
nand U13245 (N_13245,N_7749,N_9782);
nand U13246 (N_13246,N_9638,N_9957);
and U13247 (N_13247,N_10326,N_8646);
and U13248 (N_13248,N_6890,N_9788);
or U13249 (N_13249,N_8303,N_7542);
xor U13250 (N_13250,N_11688,N_7374);
nand U13251 (N_13251,N_11039,N_12029);
or U13252 (N_13252,N_9567,N_9136);
xnor U13253 (N_13253,N_6909,N_8590);
or U13254 (N_13254,N_6997,N_6577);
or U13255 (N_13255,N_12119,N_11138);
xnor U13256 (N_13256,N_9903,N_11266);
nor U13257 (N_13257,N_12168,N_6697);
xor U13258 (N_13258,N_7141,N_12164);
or U13259 (N_13259,N_7178,N_11225);
or U13260 (N_13260,N_8248,N_9331);
or U13261 (N_13261,N_12140,N_10504);
xnor U13262 (N_13262,N_6447,N_9958);
nor U13263 (N_13263,N_12113,N_7393);
xnor U13264 (N_13264,N_7194,N_9623);
nand U13265 (N_13265,N_9610,N_8252);
xnor U13266 (N_13266,N_10906,N_8747);
nand U13267 (N_13267,N_6552,N_12397);
or U13268 (N_13268,N_7697,N_11228);
xor U13269 (N_13269,N_8219,N_9835);
nor U13270 (N_13270,N_10651,N_10758);
nor U13271 (N_13271,N_10856,N_11161);
xnor U13272 (N_13272,N_9747,N_7730);
nor U13273 (N_13273,N_7297,N_6990);
nand U13274 (N_13274,N_10991,N_8786);
or U13275 (N_13275,N_9960,N_10923);
and U13276 (N_13276,N_7647,N_7574);
or U13277 (N_13277,N_10106,N_6792);
nor U13278 (N_13278,N_9535,N_6906);
nand U13279 (N_13279,N_7092,N_8894);
nand U13280 (N_13280,N_11757,N_8859);
or U13281 (N_13281,N_12054,N_11036);
xor U13282 (N_13282,N_8065,N_10934);
xor U13283 (N_13283,N_6479,N_7450);
xnor U13284 (N_13284,N_7396,N_12185);
nor U13285 (N_13285,N_9774,N_10416);
nand U13286 (N_13286,N_6768,N_7434);
and U13287 (N_13287,N_11407,N_8452);
xnor U13288 (N_13288,N_10630,N_8874);
xor U13289 (N_13289,N_12308,N_10070);
or U13290 (N_13290,N_8290,N_7152);
nand U13291 (N_13291,N_11469,N_7400);
or U13292 (N_13292,N_10633,N_9602);
nor U13293 (N_13293,N_8374,N_9795);
and U13294 (N_13294,N_7363,N_9526);
and U13295 (N_13295,N_10988,N_8603);
or U13296 (N_13296,N_10438,N_10304);
or U13297 (N_13297,N_8790,N_7711);
xnor U13298 (N_13298,N_9925,N_11276);
or U13299 (N_13299,N_10015,N_7465);
nor U13300 (N_13300,N_11365,N_10346);
xnor U13301 (N_13301,N_11124,N_7394);
nor U13302 (N_13302,N_8531,N_6543);
and U13303 (N_13303,N_9123,N_9323);
or U13304 (N_13304,N_8060,N_10858);
and U13305 (N_13305,N_12365,N_6563);
or U13306 (N_13306,N_11617,N_8329);
or U13307 (N_13307,N_8884,N_10859);
xor U13308 (N_13308,N_8428,N_6865);
nand U13309 (N_13309,N_9812,N_10151);
nor U13310 (N_13310,N_9264,N_10225);
nand U13311 (N_13311,N_11072,N_6281);
or U13312 (N_13312,N_10700,N_11354);
or U13313 (N_13313,N_11552,N_6733);
or U13314 (N_13314,N_6422,N_9394);
xor U13315 (N_13315,N_12041,N_8705);
xnor U13316 (N_13316,N_9276,N_8417);
nand U13317 (N_13317,N_7613,N_9321);
and U13318 (N_13318,N_7742,N_10174);
nand U13319 (N_13319,N_6914,N_9214);
xor U13320 (N_13320,N_7603,N_6486);
xnor U13321 (N_13321,N_9106,N_8661);
and U13322 (N_13322,N_8760,N_7174);
nand U13323 (N_13323,N_8911,N_9306);
nand U13324 (N_13324,N_7479,N_10449);
or U13325 (N_13325,N_7918,N_11964);
or U13326 (N_13326,N_12123,N_7682);
and U13327 (N_13327,N_8964,N_10545);
or U13328 (N_13328,N_9444,N_10526);
or U13329 (N_13329,N_6643,N_11867);
and U13330 (N_13330,N_10185,N_12034);
xnor U13331 (N_13331,N_10854,N_7030);
nand U13332 (N_13332,N_12255,N_10623);
nor U13333 (N_13333,N_10201,N_9385);
or U13334 (N_13334,N_6945,N_9614);
nor U13335 (N_13335,N_10528,N_10388);
nor U13336 (N_13336,N_7717,N_11839);
xnor U13337 (N_13337,N_7517,N_10549);
and U13338 (N_13338,N_6304,N_10890);
nand U13339 (N_13339,N_10881,N_6470);
nor U13340 (N_13340,N_9327,N_9669);
or U13341 (N_13341,N_11498,N_12416);
and U13342 (N_13342,N_10382,N_9426);
xor U13343 (N_13343,N_9802,N_10269);
and U13344 (N_13344,N_6746,N_7614);
nor U13345 (N_13345,N_7403,N_10572);
or U13346 (N_13346,N_9356,N_11375);
xnor U13347 (N_13347,N_7373,N_8673);
nand U13348 (N_13348,N_11849,N_7824);
nand U13349 (N_13349,N_8459,N_10475);
nand U13350 (N_13350,N_11181,N_12152);
or U13351 (N_13351,N_11165,N_7419);
and U13352 (N_13352,N_8535,N_11674);
xnor U13353 (N_13353,N_10340,N_10281);
xor U13354 (N_13354,N_11527,N_12305);
nand U13355 (N_13355,N_7462,N_12450);
and U13356 (N_13356,N_11464,N_11781);
and U13357 (N_13357,N_9821,N_8654);
xnor U13358 (N_13358,N_9734,N_8994);
xor U13359 (N_13359,N_10019,N_11465);
or U13360 (N_13360,N_6278,N_8808);
nor U13361 (N_13361,N_8188,N_11866);
or U13362 (N_13362,N_7748,N_11467);
xor U13363 (N_13363,N_10482,N_7182);
xnor U13364 (N_13364,N_9683,N_6307);
nor U13365 (N_13365,N_7760,N_10428);
xnor U13366 (N_13366,N_10043,N_8387);
nor U13367 (N_13367,N_12114,N_11198);
or U13368 (N_13368,N_10455,N_7530);
nor U13369 (N_13369,N_11744,N_11943);
nand U13370 (N_13370,N_8791,N_8289);
xor U13371 (N_13371,N_10779,N_8461);
and U13372 (N_13372,N_7343,N_11096);
nand U13373 (N_13373,N_12180,N_11522);
xor U13374 (N_13374,N_7773,N_11339);
and U13375 (N_13375,N_10502,N_9005);
or U13376 (N_13376,N_9055,N_7963);
and U13377 (N_13377,N_11961,N_9013);
xor U13378 (N_13378,N_8944,N_6926);
and U13379 (N_13379,N_6978,N_9422);
nand U13380 (N_13380,N_7699,N_8432);
and U13381 (N_13381,N_7669,N_9443);
and U13382 (N_13382,N_10905,N_11144);
and U13383 (N_13383,N_7239,N_10832);
or U13384 (N_13384,N_12431,N_8878);
xor U13385 (N_13385,N_11447,N_9374);
nand U13386 (N_13386,N_9330,N_8621);
and U13387 (N_13387,N_11727,N_7199);
and U13388 (N_13388,N_7265,N_7037);
or U13389 (N_13389,N_7482,N_7945);
xor U13390 (N_13390,N_9530,N_12475);
nor U13391 (N_13391,N_11622,N_11869);
and U13392 (N_13392,N_8845,N_6940);
nor U13393 (N_13393,N_10747,N_9051);
xor U13394 (N_13394,N_11020,N_7077);
nand U13395 (N_13395,N_6324,N_9641);
xor U13396 (N_13396,N_10963,N_8245);
or U13397 (N_13397,N_9402,N_11636);
xor U13398 (N_13398,N_11004,N_7036);
nor U13399 (N_13399,N_12139,N_7430);
nor U13400 (N_13400,N_6292,N_6568);
xnor U13401 (N_13401,N_6315,N_10661);
nand U13402 (N_13402,N_11322,N_11966);
and U13403 (N_13403,N_9408,N_6763);
nor U13404 (N_13404,N_8497,N_6754);
nor U13405 (N_13405,N_9708,N_9864);
xor U13406 (N_13406,N_6739,N_11923);
and U13407 (N_13407,N_11589,N_10501);
xor U13408 (N_13408,N_6423,N_6345);
xor U13409 (N_13409,N_9468,N_10246);
nor U13410 (N_13410,N_11594,N_6411);
and U13411 (N_13411,N_11007,N_9949);
and U13412 (N_13412,N_8551,N_11420);
nand U13413 (N_13413,N_9608,N_8286);
and U13414 (N_13414,N_10194,N_10872);
or U13415 (N_13415,N_10483,N_9675);
xor U13416 (N_13416,N_6833,N_11256);
xnor U13417 (N_13417,N_6885,N_7218);
nand U13418 (N_13418,N_11437,N_10062);
nor U13419 (N_13419,N_9865,N_8602);
xnor U13420 (N_13420,N_7066,N_6596);
xnor U13421 (N_13421,N_11535,N_7256);
and U13422 (N_13422,N_7284,N_10270);
or U13423 (N_13423,N_10026,N_7320);
xor U13424 (N_13424,N_7869,N_7852);
nand U13425 (N_13425,N_6621,N_11715);
or U13426 (N_13426,N_9205,N_11788);
nor U13427 (N_13427,N_9833,N_12398);
nand U13428 (N_13428,N_10539,N_8113);
or U13429 (N_13429,N_9375,N_11312);
or U13430 (N_13430,N_10722,N_7572);
xnor U13431 (N_13431,N_8737,N_9642);
nor U13432 (N_13432,N_10597,N_8888);
or U13433 (N_13433,N_6251,N_11048);
nor U13434 (N_13434,N_9185,N_9977);
and U13435 (N_13435,N_8526,N_12147);
nand U13436 (N_13436,N_7142,N_6572);
or U13437 (N_13437,N_6531,N_6608);
xor U13438 (N_13438,N_10339,N_7646);
nor U13439 (N_13439,N_9059,N_6999);
nand U13440 (N_13440,N_7875,N_6268);
xnor U13441 (N_13441,N_10267,N_9147);
or U13442 (N_13442,N_10588,N_12451);
xnor U13443 (N_13443,N_11706,N_6813);
nor U13444 (N_13444,N_6492,N_11340);
and U13445 (N_13445,N_7553,N_7388);
nand U13446 (N_13446,N_11925,N_12181);
nand U13447 (N_13447,N_10264,N_6635);
and U13448 (N_13448,N_8496,N_10701);
nor U13449 (N_13449,N_11587,N_11406);
xor U13450 (N_13450,N_6564,N_11019);
and U13451 (N_13451,N_12373,N_11307);
xnor U13452 (N_13452,N_11536,N_10627);
and U13453 (N_13453,N_11547,N_11179);
nor U13454 (N_13454,N_6585,N_7569);
or U13455 (N_13455,N_11253,N_11275);
xor U13456 (N_13456,N_7708,N_11005);
nor U13457 (N_13457,N_7108,N_8118);
nand U13458 (N_13458,N_7321,N_11336);
and U13459 (N_13459,N_8376,N_7685);
xnor U13460 (N_13460,N_10571,N_10897);
and U13461 (N_13461,N_7565,N_7878);
or U13462 (N_13462,N_10744,N_8215);
nand U13463 (N_13463,N_10992,N_8907);
or U13464 (N_13464,N_8391,N_8990);
or U13465 (N_13465,N_9717,N_6250);
and U13466 (N_13466,N_6446,N_10983);
and U13467 (N_13467,N_11209,N_12328);
and U13468 (N_13468,N_12124,N_7144);
and U13469 (N_13469,N_7716,N_9441);
nand U13470 (N_13470,N_12307,N_10883);
and U13471 (N_13471,N_11793,N_7444);
and U13472 (N_13472,N_12051,N_11251);
nor U13473 (N_13473,N_7478,N_7008);
and U13474 (N_13474,N_12165,N_10080);
and U13475 (N_13475,N_8631,N_9431);
xor U13476 (N_13476,N_12342,N_10969);
or U13477 (N_13477,N_11106,N_11590);
nor U13478 (N_13478,N_10668,N_6416);
and U13479 (N_13479,N_7738,N_8570);
xor U13480 (N_13480,N_11259,N_6327);
nand U13481 (N_13481,N_10391,N_11950);
nand U13482 (N_13482,N_11565,N_6262);
xor U13483 (N_13483,N_7534,N_6448);
or U13484 (N_13484,N_12013,N_10163);
or U13485 (N_13485,N_8846,N_9780);
xor U13486 (N_13486,N_10849,N_9182);
or U13487 (N_13487,N_11169,N_12436);
and U13488 (N_13488,N_11654,N_9854);
nor U13489 (N_13489,N_10537,N_8867);
nand U13490 (N_13490,N_12267,N_11655);
and U13491 (N_13491,N_10564,N_8024);
and U13492 (N_13492,N_7305,N_7378);
nand U13493 (N_13493,N_11720,N_6913);
xor U13494 (N_13494,N_6920,N_8466);
nor U13495 (N_13495,N_10172,N_6933);
nor U13496 (N_13496,N_11558,N_8186);
and U13497 (N_13497,N_8916,N_9716);
xor U13498 (N_13498,N_6812,N_9825);
nor U13499 (N_13499,N_10797,N_7652);
xnor U13500 (N_13500,N_9449,N_9731);
nor U13501 (N_13501,N_10073,N_6886);
or U13502 (N_13502,N_10465,N_8679);
or U13503 (N_13503,N_11968,N_10857);
nand U13504 (N_13504,N_9244,N_11620);
nor U13505 (N_13505,N_7833,N_12145);
and U13506 (N_13506,N_7516,N_12327);
nand U13507 (N_13507,N_10478,N_9003);
xnor U13508 (N_13508,N_8692,N_8636);
nor U13509 (N_13509,N_10458,N_6265);
and U13510 (N_13510,N_8306,N_11379);
xnor U13511 (N_13511,N_10393,N_11377);
nor U13512 (N_13512,N_12482,N_11109);
and U13513 (N_13513,N_8125,N_10235);
nand U13514 (N_13514,N_6269,N_8668);
xnor U13515 (N_13515,N_11580,N_7275);
nand U13516 (N_13516,N_9837,N_7251);
nand U13517 (N_13517,N_9346,N_12193);
and U13518 (N_13518,N_10739,N_11427);
nor U13519 (N_13519,N_12435,N_9367);
or U13520 (N_13520,N_11734,N_11373);
nor U13521 (N_13521,N_6255,N_6309);
xnor U13522 (N_13522,N_12132,N_8287);
xnor U13523 (N_13523,N_10132,N_7887);
nor U13524 (N_13524,N_12494,N_11659);
nand U13525 (N_13525,N_7001,N_9122);
nand U13526 (N_13526,N_8318,N_9741);
nand U13527 (N_13527,N_11583,N_8824);
xor U13528 (N_13528,N_8793,N_12049);
xor U13529 (N_13529,N_9846,N_6852);
nor U13530 (N_13530,N_10308,N_7032);
and U13531 (N_13531,N_10941,N_6829);
xnor U13532 (N_13532,N_11922,N_11926);
nor U13533 (N_13533,N_11268,N_7317);
nor U13534 (N_13534,N_11333,N_10893);
nand U13535 (N_13535,N_7010,N_11502);
and U13536 (N_13536,N_7238,N_7808);
xor U13537 (N_13537,N_9388,N_9513);
nor U13538 (N_13538,N_8998,N_12480);
or U13539 (N_13539,N_6282,N_12091);
and U13540 (N_13540,N_6550,N_7476);
or U13541 (N_13541,N_8198,N_6579);
nand U13542 (N_13542,N_6876,N_6594);
and U13543 (N_13543,N_7552,N_9031);
nand U13544 (N_13544,N_11021,N_9738);
nand U13545 (N_13545,N_7645,N_7274);
nand U13546 (N_13546,N_10924,N_9759);
xor U13547 (N_13547,N_12074,N_9308);
xnor U13548 (N_13548,N_9891,N_8547);
nand U13549 (N_13549,N_11153,N_7024);
nor U13550 (N_13550,N_9436,N_10290);
xor U13551 (N_13551,N_11784,N_11016);
or U13552 (N_13552,N_10685,N_12216);
nor U13553 (N_13553,N_8424,N_6671);
nand U13554 (N_13554,N_9655,N_6723);
nand U13555 (N_13555,N_11742,N_9009);
and U13556 (N_13556,N_8953,N_7098);
or U13557 (N_13557,N_11466,N_6628);
nand U13558 (N_13558,N_6712,N_11082);
or U13559 (N_13559,N_9291,N_8067);
nor U13560 (N_13560,N_8162,N_7151);
nor U13561 (N_13561,N_7683,N_9755);
or U13562 (N_13562,N_7821,N_10364);
nand U13563 (N_13563,N_7861,N_8128);
and U13564 (N_13564,N_7589,N_9393);
nand U13565 (N_13565,N_8383,N_12350);
and U13566 (N_13566,N_11669,N_9151);
xnor U13567 (N_13567,N_7060,N_7913);
nand U13568 (N_13568,N_12338,N_6323);
xor U13569 (N_13569,N_8961,N_7600);
nand U13570 (N_13570,N_7632,N_9172);
xor U13571 (N_13571,N_7663,N_9240);
xnor U13572 (N_13572,N_9624,N_7469);
nor U13573 (N_13573,N_9404,N_7921);
and U13574 (N_13574,N_10493,N_9859);
and U13575 (N_13575,N_12389,N_11624);
xor U13576 (N_13576,N_11559,N_11962);
nand U13577 (N_13577,N_11399,N_12437);
or U13578 (N_13578,N_10861,N_10255);
nand U13579 (N_13579,N_8231,N_11403);
or U13580 (N_13580,N_9149,N_7086);
and U13581 (N_13581,N_11728,N_8332);
and U13582 (N_13582,N_8569,N_8875);
nor U13583 (N_13583,N_7420,N_11683);
nor U13584 (N_13584,N_11131,N_7495);
or U13585 (N_13585,N_7402,N_10191);
xor U13586 (N_13586,N_8315,N_8573);
nor U13587 (N_13587,N_8001,N_10118);
nand U13588 (N_13588,N_10863,N_9761);
or U13589 (N_13589,N_12384,N_7888);
or U13590 (N_13590,N_10245,N_10454);
and U13591 (N_13591,N_11480,N_9187);
nand U13592 (N_13592,N_12331,N_8365);
and U13593 (N_13593,N_6858,N_7160);
and U13594 (N_13594,N_6337,N_6376);
xor U13595 (N_13595,N_11711,N_11121);
nand U13596 (N_13596,N_6540,N_9869);
or U13597 (N_13597,N_6818,N_10632);
or U13598 (N_13598,N_11871,N_11063);
nor U13599 (N_13599,N_10028,N_8708);
nand U13600 (N_13600,N_8177,N_8016);
nor U13601 (N_13601,N_10313,N_7702);
nor U13602 (N_13602,N_8400,N_6808);
xnor U13603 (N_13603,N_7246,N_9146);
nand U13604 (N_13604,N_12473,N_9657);
nor U13605 (N_13605,N_11670,N_9601);
or U13606 (N_13606,N_11947,N_11600);
xnor U13607 (N_13607,N_8240,N_8075);
nor U13608 (N_13608,N_6958,N_10777);
xor U13609 (N_13609,N_6828,N_8279);
or U13610 (N_13610,N_12223,N_7237);
nor U13611 (N_13611,N_11772,N_7528);
nand U13612 (N_13612,N_8773,N_11666);
and U13613 (N_13613,N_8314,N_9603);
or U13614 (N_13614,N_10643,N_6320);
xnor U13615 (N_13615,N_11006,N_10972);
and U13616 (N_13616,N_7633,N_10745);
or U13617 (N_13617,N_6514,N_9178);
and U13618 (N_13618,N_10262,N_8743);
and U13619 (N_13619,N_11318,N_7688);
xnor U13620 (N_13620,N_11578,N_7176);
xor U13621 (N_13621,N_7384,N_10143);
nand U13622 (N_13622,N_10134,N_11737);
xnor U13623 (N_13623,N_9161,N_8900);
or U13624 (N_13624,N_11660,N_9188);
nand U13625 (N_13625,N_12422,N_8035);
nor U13626 (N_13626,N_12022,N_11111);
xor U13627 (N_13627,N_11810,N_6379);
or U13628 (N_13628,N_7538,N_8023);
or U13629 (N_13629,N_10022,N_12433);
and U13630 (N_13630,N_7865,N_11806);
nand U13631 (N_13631,N_7707,N_11151);
nor U13632 (N_13632,N_9678,N_6457);
nor U13633 (N_13633,N_6264,N_9198);
xnor U13634 (N_13634,N_6331,N_9726);
or U13635 (N_13635,N_11671,N_9357);
and U13636 (N_13636,N_11507,N_6399);
nand U13637 (N_13637,N_11886,N_7245);
and U13638 (N_13638,N_10226,N_7003);
or U13639 (N_13639,N_12010,N_9409);
or U13640 (N_13640,N_7768,N_7965);
xnor U13641 (N_13641,N_9983,N_6353);
nand U13642 (N_13642,N_9077,N_6647);
nor U13643 (N_13643,N_12470,N_8557);
nor U13644 (N_13644,N_6802,N_10908);
nor U13645 (N_13645,N_12306,N_9360);
or U13646 (N_13646,N_11148,N_7436);
nor U13647 (N_13647,N_9501,N_9528);
xnor U13648 (N_13648,N_7867,N_6742);
and U13649 (N_13649,N_9625,N_10309);
nor U13650 (N_13650,N_11394,N_10089);
xnor U13651 (N_13651,N_8802,N_7853);
nand U13652 (N_13652,N_7007,N_11646);
xnor U13653 (N_13653,N_9645,N_11176);
nor U13654 (N_13654,N_9459,N_8598);
xnor U13655 (N_13655,N_9403,N_9398);
nand U13656 (N_13656,N_9253,N_8932);
and U13657 (N_13657,N_8073,N_8652);
xor U13658 (N_13658,N_9811,N_6570);
and U13659 (N_13659,N_7153,N_6782);
or U13660 (N_13660,N_8143,N_6725);
or U13661 (N_13661,N_9428,N_11022);
nand U13662 (N_13662,N_10788,N_11582);
xor U13663 (N_13663,N_9851,N_11911);
nand U13664 (N_13664,N_10139,N_10684);
nand U13665 (N_13665,N_9710,N_10591);
or U13666 (N_13666,N_7745,N_7548);
xor U13667 (N_13667,N_11883,N_7339);
xor U13668 (N_13668,N_12188,N_6747);
xnor U13669 (N_13669,N_7882,N_10692);
nand U13670 (N_13670,N_7802,N_11349);
or U13671 (N_13671,N_6276,N_12272);
nor U13672 (N_13672,N_8973,N_8816);
nor U13673 (N_13673,N_12339,N_11974);
nor U13674 (N_13674,N_9580,N_8053);
or U13675 (N_13675,N_7046,N_12059);
xnor U13676 (N_13676,N_11640,N_10617);
xnor U13677 (N_13677,N_10613,N_8558);
and U13678 (N_13678,N_7100,N_8715);
xnor U13679 (N_13679,N_11887,N_9108);
nor U13680 (N_13680,N_7527,N_9391);
nand U13681 (N_13681,N_12265,N_7537);
xnor U13682 (N_13682,N_10589,N_6977);
xnor U13683 (N_13683,N_11504,N_10957);
or U13684 (N_13684,N_9515,N_9350);
xor U13685 (N_13685,N_6880,N_7555);
and U13686 (N_13686,N_8307,N_10540);
nor U13687 (N_13687,N_11986,N_8622);
nand U13688 (N_13688,N_6902,N_7915);
xor U13689 (N_13689,N_7969,N_7353);
xor U13690 (N_13690,N_9883,N_7658);
and U13691 (N_13691,N_12340,N_9165);
nand U13692 (N_13692,N_7883,N_9101);
and U13693 (N_13693,N_8087,N_6266);
nor U13694 (N_13694,N_6944,N_9176);
nor U13695 (N_13695,N_9594,N_12354);
and U13696 (N_13696,N_8667,N_7992);
xnor U13697 (N_13697,N_10055,N_7832);
or U13698 (N_13698,N_7038,N_7620);
and U13699 (N_13699,N_9707,N_8339);
or U13700 (N_13700,N_9994,N_7287);
nor U13701 (N_13701,N_8410,N_10955);
nor U13702 (N_13702,N_10183,N_12420);
and U13703 (N_13703,N_12024,N_7186);
and U13704 (N_13704,N_9034,N_11284);
xnor U13705 (N_13705,N_10173,N_8672);
xor U13706 (N_13706,N_12198,N_6762);
xnor U13707 (N_13707,N_9091,N_8320);
or U13708 (N_13708,N_11010,N_11252);
nor U13709 (N_13709,N_10782,N_11572);
nor U13710 (N_13710,N_11300,N_6487);
nor U13711 (N_13711,N_7986,N_8920);
xnor U13712 (N_13712,N_6706,N_8059);
and U13713 (N_13713,N_11000,N_9998);
nand U13714 (N_13714,N_10471,N_12449);
nor U13715 (N_13715,N_6546,N_11800);
nand U13716 (N_13716,N_11012,N_6924);
xnor U13717 (N_13717,N_6925,N_11913);
xor U13718 (N_13718,N_7872,N_8817);
or U13719 (N_13719,N_8960,N_10792);
nor U13720 (N_13720,N_6664,N_8226);
xnor U13721 (N_13721,N_11551,N_10989);
and U13722 (N_13722,N_11593,N_6504);
nand U13723 (N_13723,N_12073,N_11001);
and U13724 (N_13724,N_9793,N_10261);
nand U13725 (N_13725,N_6846,N_7236);
xor U13726 (N_13726,N_7249,N_10215);
or U13727 (N_13727,N_11040,N_7313);
or U13728 (N_13728,N_9832,N_11071);
xor U13729 (N_13729,N_12008,N_7944);
and U13730 (N_13730,N_10670,N_11459);
and U13731 (N_13731,N_6722,N_9666);
or U13732 (N_13732,N_7054,N_12221);
nand U13733 (N_13733,N_8360,N_11758);
or U13734 (N_13734,N_11486,N_7765);
and U13735 (N_13735,N_10958,N_10979);
nand U13736 (N_13736,N_11410,N_9540);
nand U13737 (N_13737,N_7031,N_9236);
nor U13738 (N_13738,N_12247,N_11566);
xor U13739 (N_13739,N_8536,N_6573);
xnor U13740 (N_13740,N_11383,N_10659);
or U13741 (N_13741,N_6653,N_7452);
and U13742 (N_13742,N_8966,N_10853);
xnor U13743 (N_13743,N_11139,N_6708);
and U13744 (N_13744,N_11224,N_12228);
xor U13745 (N_13745,N_11729,N_10835);
or U13746 (N_13746,N_7367,N_11802);
xor U13747 (N_13747,N_9027,N_9751);
and U13748 (N_13748,N_9494,N_8511);
nor U13749 (N_13749,N_7529,N_10121);
nand U13750 (N_13750,N_6300,N_10329);
nand U13751 (N_13751,N_11993,N_12427);
or U13752 (N_13752,N_12276,N_10938);
or U13753 (N_13753,N_12486,N_11368);
nor U13754 (N_13754,N_11528,N_7226);
nand U13755 (N_13755,N_7789,N_7609);
or U13756 (N_13756,N_10044,N_9089);
or U13757 (N_13757,N_10921,N_7950);
or U13758 (N_13758,N_7191,N_8733);
nand U13759 (N_13759,N_11631,N_10442);
or U13760 (N_13760,N_8019,N_7437);
nor U13761 (N_13761,N_12009,N_7618);
xnor U13762 (N_13762,N_11295,N_10615);
nor U13763 (N_13763,N_8239,N_10956);
and U13764 (N_13764,N_8342,N_11783);
xnor U13765 (N_13765,N_8036,N_6385);
xnor U13766 (N_13766,N_11451,N_11607);
and U13767 (N_13767,N_7594,N_9511);
or U13768 (N_13768,N_8595,N_10381);
xnor U13769 (N_13769,N_8403,N_7931);
or U13770 (N_13770,N_11997,N_9690);
or U13771 (N_13771,N_6771,N_10399);
xor U13772 (N_13772,N_8380,N_9523);
nand U13773 (N_13773,N_9029,N_11041);
or U13774 (N_13774,N_11055,N_12468);
or U13775 (N_13775,N_10491,N_12105);
xnor U13776 (N_13776,N_8985,N_12127);
nand U13777 (N_13777,N_8115,N_7356);
nand U13778 (N_13778,N_9035,N_12088);
and U13779 (N_13779,N_8593,N_7803);
and U13780 (N_13780,N_8642,N_12361);
and U13781 (N_13781,N_11083,N_7070);
and U13782 (N_13782,N_8576,N_9143);
and U13783 (N_13783,N_11404,N_9312);
xnor U13784 (N_13784,N_9270,N_8304);
or U13785 (N_13785,N_6918,N_6616);
and U13786 (N_13786,N_12448,N_8524);
nand U13787 (N_13787,N_9130,N_7340);
or U13788 (N_13788,N_11818,N_9458);
nor U13789 (N_13789,N_7729,N_9933);
or U13790 (N_13790,N_10199,N_7972);
nand U13791 (N_13791,N_6951,N_7344);
xnor U13792 (N_13792,N_6518,N_8375);
nor U13793 (N_13793,N_12314,N_10558);
xnor U13794 (N_13794,N_7128,N_8718);
or U13795 (N_13795,N_7312,N_12458);
nand U13796 (N_13796,N_11080,N_8166);
nor U13797 (N_13797,N_9736,N_7431);
nand U13798 (N_13798,N_7366,N_12390);
nand U13799 (N_13799,N_6799,N_6655);
or U13800 (N_13800,N_10587,N_11653);
nor U13801 (N_13801,N_9348,N_10033);
xnor U13802 (N_13802,N_11489,N_11790);
or U13803 (N_13803,N_10544,N_8996);
nand U13804 (N_13804,N_9527,N_8470);
or U13805 (N_13805,N_7897,N_8632);
and U13806 (N_13806,N_6984,N_8353);
xor U13807 (N_13807,N_10488,N_7447);
nor U13808 (N_13808,N_9097,N_6648);
and U13809 (N_13809,N_9266,N_6783);
and U13810 (N_13810,N_12359,N_11725);
nor U13811 (N_13811,N_6775,N_9924);
nor U13812 (N_13812,N_10947,N_11215);
nor U13813 (N_13813,N_7282,N_7161);
and U13814 (N_13814,N_9661,N_9471);
nand U13815 (N_13815,N_10122,N_11694);
nand U13816 (N_13816,N_11476,N_7243);
or U13817 (N_13817,N_7467,N_6310);
or U13818 (N_13818,N_8149,N_12412);
or U13819 (N_13819,N_10310,N_12239);
nand U13820 (N_13820,N_8082,N_9261);
nand U13821 (N_13821,N_10886,N_12157);
nor U13822 (N_13822,N_7983,N_10017);
and U13823 (N_13823,N_9879,N_11807);
nand U13824 (N_13824,N_8914,N_7820);
nor U13825 (N_13825,N_9918,N_8484);
or U13826 (N_13826,N_12419,N_8095);
nor U13827 (N_13827,N_7694,N_11358);
xnor U13828 (N_13828,N_11411,N_10030);
or U13829 (N_13829,N_9434,N_9750);
xnor U13830 (N_13830,N_9466,N_10336);
and U13831 (N_13831,N_7541,N_10681);
and U13832 (N_13832,N_8805,N_9772);
nor U13833 (N_13833,N_7571,N_8748);
or U13834 (N_13834,N_11696,N_6826);
nand U13835 (N_13835,N_10850,N_8114);
or U13836 (N_13836,N_6989,N_9293);
and U13837 (N_13837,N_10414,N_12367);
nor U13838 (N_13838,N_6554,N_10741);
and U13839 (N_13839,N_8704,N_12461);
nor U13840 (N_13840,N_9982,N_8251);
nand U13841 (N_13841,N_9339,N_6784);
nor U13842 (N_13842,N_11677,N_7125);
or U13843 (N_13843,N_8983,N_6454);
or U13844 (N_13844,N_11743,N_8801);
nand U13845 (N_13845,N_6869,N_7561);
and U13846 (N_13846,N_12061,N_12136);
nor U13847 (N_13847,N_11133,N_8987);
or U13848 (N_13848,N_10004,N_6394);
and U13849 (N_13849,N_10833,N_10202);
and U13850 (N_13850,N_8946,N_10405);
nand U13851 (N_13851,N_6581,N_7025);
nor U13852 (N_13852,N_9016,N_12343);
and U13853 (N_13853,N_7838,N_10283);
xnor U13854 (N_13854,N_10621,N_11845);
nor U13855 (N_13855,N_11330,N_8214);
nand U13856 (N_13856,N_9598,N_6507);
or U13857 (N_13857,N_8811,N_7457);
nor U13858 (N_13858,N_8412,N_9474);
xnor U13859 (N_13859,N_9423,N_7071);
or U13860 (N_13860,N_6270,N_9280);
xnor U13861 (N_13861,N_10660,N_12194);
nor U13862 (N_13862,N_6556,N_7490);
nand U13863 (N_13863,N_9971,N_10461);
nor U13864 (N_13864,N_9786,N_6700);
or U13865 (N_13865,N_9224,N_9353);
or U13866 (N_13866,N_10230,N_9691);
nand U13867 (N_13867,N_10878,N_7472);
or U13868 (N_13868,N_12254,N_8351);
and U13869 (N_13869,N_8195,N_7778);
nor U13870 (N_13870,N_6284,N_7641);
and U13871 (N_13871,N_7018,N_8675);
or U13872 (N_13872,N_12457,N_9930);
nor U13873 (N_13873,N_10415,N_8119);
xnor U13874 (N_13874,N_12315,N_7612);
nand U13875 (N_13875,N_6414,N_8433);
or U13876 (N_13876,N_7968,N_10508);
xnor U13877 (N_13877,N_9067,N_10974);
nor U13878 (N_13878,N_12362,N_8890);
xnor U13879 (N_13879,N_6850,N_6432);
nand U13880 (N_13880,N_12016,N_11855);
and U13881 (N_13881,N_11709,N_8749);
or U13882 (N_13882,N_12490,N_7424);
nand U13883 (N_13883,N_6371,N_7774);
or U13884 (N_13884,N_8187,N_12082);
and U13885 (N_13885,N_8393,N_9945);
or U13886 (N_13886,N_12171,N_7330);
nand U13887 (N_13887,N_8430,N_7043);
nor U13888 (N_13888,N_8716,N_6499);
nor U13889 (N_13889,N_11537,N_12014);
nor U13890 (N_13890,N_7422,N_9680);
xor U13891 (N_13891,N_7315,N_8152);
nor U13892 (N_13892,N_9770,N_11717);
and U13893 (N_13893,N_9928,N_12400);
or U13894 (N_13894,N_6857,N_8662);
xor U13895 (N_13895,N_7926,N_10468);
or U13896 (N_13896,N_11217,N_10565);
nor U13897 (N_13897,N_8873,N_6855);
nor U13898 (N_13898,N_11994,N_10925);
and U13899 (N_13899,N_10954,N_11047);
or U13900 (N_13900,N_7679,N_12439);
and U13901 (N_13901,N_11107,N_7962);
xnor U13902 (N_13902,N_9562,N_6328);
or U13903 (N_13903,N_7016,N_11281);
and U13904 (N_13904,N_7372,N_11526);
nand U13905 (N_13905,N_11178,N_12062);
xor U13906 (N_13906,N_10484,N_11533);
or U13907 (N_13907,N_8211,N_8897);
nor U13908 (N_13908,N_10774,N_11110);
or U13909 (N_13909,N_10600,N_8157);
or U13910 (N_13910,N_7998,N_6393);
xor U13911 (N_13911,N_8788,N_10322);
and U13912 (N_13912,N_9311,N_9364);
xnor U13913 (N_13913,N_12309,N_9950);
nor U13914 (N_13914,N_6458,N_6392);
nand U13915 (N_13915,N_10536,N_10373);
nor U13916 (N_13916,N_11374,N_7136);
nor U13917 (N_13917,N_10368,N_11473);
and U13918 (N_13918,N_11596,N_10731);
nand U13919 (N_13919,N_11908,N_7982);
xnor U13920 (N_13920,N_9505,N_6391);
and U13921 (N_13921,N_9279,N_8549);
nor U13922 (N_13922,N_10490,N_8510);
or U13923 (N_13923,N_10998,N_11503);
nand U13924 (N_13924,N_6465,N_11761);
nor U13925 (N_13925,N_9347,N_7135);
or U13926 (N_13926,N_12184,N_8302);
nor U13927 (N_13927,N_6624,N_7890);
nor U13928 (N_13928,N_10377,N_9342);
and U13929 (N_13929,N_7354,N_9069);
or U13930 (N_13930,N_6503,N_7213);
or U13931 (N_13931,N_8834,N_6366);
or U13932 (N_13932,N_12236,N_10291);
and U13933 (N_13933,N_8056,N_8578);
xor U13934 (N_13934,N_11561,N_11453);
and U13935 (N_13935,N_7500,N_11909);
nand U13936 (N_13936,N_6724,N_8883);
nor U13937 (N_13937,N_7481,N_10907);
or U13938 (N_13938,N_12363,N_11013);
and U13939 (N_13939,N_8641,N_10614);
nand U13940 (N_13940,N_12324,N_6451);
or U13941 (N_13941,N_6380,N_9201);
nand U13942 (N_13942,N_9537,N_6571);
or U13943 (N_13943,N_7361,N_7819);
or U13944 (N_13944,N_7788,N_6815);
nor U13945 (N_13945,N_6654,N_6966);
nand U13946 (N_13946,N_6814,N_8266);
or U13947 (N_13947,N_6823,N_6330);
and U13948 (N_13948,N_6859,N_11363);
and U13949 (N_13949,N_6811,N_7744);
nand U13950 (N_13950,N_7451,N_9600);
nand U13951 (N_13951,N_10803,N_9181);
nor U13952 (N_13952,N_7843,N_7268);
nor U13953 (N_13953,N_10894,N_8192);
and U13954 (N_13954,N_11668,N_7116);
nor U13955 (N_13955,N_9796,N_11978);
nand U13956 (N_13956,N_8627,N_9836);
and U13957 (N_13957,N_7643,N_8746);
nand U13958 (N_13958,N_7961,N_9215);
or U13959 (N_13959,N_6591,N_9878);
and U13960 (N_13960,N_9804,N_7922);
or U13961 (N_13961,N_6523,N_7453);
nor U13962 (N_13962,N_6805,N_12006);
or U13963 (N_13963,N_8420,N_6981);
nand U13964 (N_13964,N_8921,N_12261);
xnor U13965 (N_13965,N_8481,N_10930);
nor U13966 (N_13966,N_6840,N_11098);
nor U13967 (N_13967,N_11884,N_8995);
and U13968 (N_13968,N_6420,N_11146);
nor U13969 (N_13969,N_10767,N_6261);
and U13970 (N_13970,N_11282,N_11501);
and U13971 (N_13971,N_8993,N_9281);
nor U13972 (N_13972,N_8709,N_7939);
and U13973 (N_13973,N_8227,N_10593);
or U13974 (N_13974,N_9936,N_8096);
or U13975 (N_13975,N_10822,N_7229);
xor U13976 (N_13976,N_12083,N_12108);
or U13977 (N_13977,N_7193,N_11249);
nand U13978 (N_13978,N_9948,N_9287);
nand U13979 (N_13979,N_11872,N_12318);
and U13980 (N_13980,N_9684,N_6605);
and U13981 (N_13981,N_11018,N_7973);
nor U13982 (N_13982,N_9301,N_9171);
or U13983 (N_13983,N_10100,N_12474);
and U13984 (N_13984,N_8582,N_10075);
and U13985 (N_13985,N_9232,N_7740);
xnor U13986 (N_13986,N_8744,N_7775);
nand U13987 (N_13987,N_9889,N_11610);
or U13988 (N_13988,N_11534,N_6301);
nor U13989 (N_13989,N_8438,N_7408);
xor U13990 (N_13990,N_8525,N_7473);
xnor U13991 (N_13991,N_11416,N_10534);
nor U13992 (N_13992,N_8029,N_8244);
xor U13993 (N_13993,N_8620,N_8346);
nand U13994 (N_13994,N_9138,N_8431);
and U13995 (N_13995,N_6693,N_7002);
xnor U13996 (N_13996,N_7441,N_8358);
or U13997 (N_13997,N_8490,N_10771);
or U13998 (N_13998,N_7188,N_10242);
or U13999 (N_13999,N_7562,N_7876);
nand U14000 (N_14000,N_6780,N_6629);
or U14001 (N_14001,N_8506,N_11664);
nand U14002 (N_14002,N_10909,N_10825);
or U14003 (N_14003,N_8903,N_10601);
nor U14004 (N_14004,N_6972,N_11857);
nand U14005 (N_14005,N_11910,N_7072);
nand U14006 (N_14006,N_9030,N_6267);
nand U14007 (N_14007,N_10799,N_10860);
or U14008 (N_14008,N_11087,N_10274);
or U14009 (N_14009,N_10560,N_8132);
nor U14010 (N_14010,N_11835,N_7133);
nand U14011 (N_14011,N_10901,N_12415);
nor U14012 (N_14012,N_10775,N_11306);
nor U14013 (N_14013,N_11247,N_10806);
and U14014 (N_14014,N_12484,N_8325);
or U14015 (N_14015,N_10386,N_9732);
nor U14016 (N_14016,N_9566,N_12146);
or U14017 (N_14017,N_9448,N_6911);
nand U14018 (N_14018,N_6888,N_9345);
or U14019 (N_14019,N_8070,N_7818);
xor U14020 (N_14020,N_8111,N_11933);
or U14021 (N_14021,N_8421,N_9076);
xnor U14022 (N_14022,N_6450,N_9715);
nand U14023 (N_14023,N_7608,N_7958);
nand U14024 (N_14024,N_7085,N_10679);
nand U14025 (N_14025,N_11134,N_10530);
nor U14026 (N_14026,N_9959,N_11038);
or U14027 (N_14027,N_9453,N_11651);
and U14028 (N_14028,N_9368,N_7326);
nor U14029 (N_14029,N_11370,N_7651);
xor U14030 (N_14030,N_9479,N_10120);
nand U14031 (N_14031,N_8028,N_9743);
and U14032 (N_14032,N_7917,N_7406);
nor U14033 (N_14033,N_12056,N_6936);
nor U14034 (N_14034,N_7439,N_7341);
and U14035 (N_14035,N_10847,N_11362);
nor U14036 (N_14036,N_12432,N_12063);
nor U14037 (N_14037,N_11609,N_11239);
nand U14038 (N_14038,N_9733,N_10234);
or U14039 (N_14039,N_11093,N_9195);
or U14040 (N_14040,N_12031,N_8594);
xor U14041 (N_14041,N_12326,N_7985);
nor U14042 (N_14042,N_12133,N_10705);
xnor U14043 (N_14043,N_6785,N_8021);
or U14044 (N_14044,N_12273,N_6462);
xnor U14045 (N_14045,N_8172,N_7905);
xnor U14046 (N_14046,N_6506,N_12405);
or U14047 (N_14047,N_7519,N_11763);
xor U14048 (N_14048,N_11230,N_9145);
nand U14049 (N_14049,N_8819,N_8676);
nor U14050 (N_14050,N_11567,N_12179);
and U14051 (N_14051,N_7840,N_6674);
nor U14052 (N_14052,N_7044,N_9712);
and U14053 (N_14053,N_11979,N_10801);
or U14054 (N_14054,N_7139,N_9626);
and U14055 (N_14055,N_6368,N_10505);
or U14056 (N_14056,N_11903,N_8542);
or U14057 (N_14057,N_7741,N_10725);
nor U14058 (N_14058,N_12456,N_11254);
nor U14059 (N_14059,N_11920,N_8308);
nand U14060 (N_14060,N_11934,N_7673);
and U14061 (N_14061,N_11808,N_9475);
or U14062 (N_14062,N_6362,N_10622);
xor U14063 (N_14063,N_11679,N_11130);
nand U14064 (N_14064,N_10892,N_6437);
and U14065 (N_14065,N_7604,N_11894);
nor U14066 (N_14066,N_11364,N_8980);
xnor U14067 (N_14067,N_12068,N_9366);
and U14068 (N_14068,N_9895,N_7866);
nor U14069 (N_14069,N_10815,N_7987);
and U14070 (N_14070,N_11129,N_11174);
nor U14071 (N_14071,N_12320,N_8258);
xor U14072 (N_14072,N_6959,N_10181);
xor U14073 (N_14073,N_6743,N_10864);
xor U14074 (N_14074,N_11987,N_9309);
nor U14075 (N_14075,N_11585,N_9210);
nor U14076 (N_14076,N_9503,N_8955);
nor U14077 (N_14077,N_7189,N_8559);
nand U14078 (N_14078,N_9329,N_6485);
nand U14079 (N_14079,N_6532,N_9863);
or U14080 (N_14080,N_8653,N_11270);
xor U14081 (N_14081,N_7207,N_9543);
and U14082 (N_14082,N_12101,N_8588);
nand U14083 (N_14083,N_9843,N_9131);
nor U14084 (N_14084,N_7159,N_10116);
or U14085 (N_14085,N_9730,N_6968);
nor U14086 (N_14086,N_9980,N_11035);
xnor U14087 (N_14087,N_10772,N_12492);
nand U14088 (N_14088,N_11977,N_10728);
nand U14089 (N_14089,N_11778,N_8293);
or U14090 (N_14090,N_6400,N_8610);
nand U14091 (N_14091,N_10770,N_6976);
xor U14092 (N_14092,N_8703,N_9723);
xnor U14093 (N_14093,N_6293,N_7991);
xnor U14094 (N_14094,N_7398,N_6349);
nand U14095 (N_14095,N_9532,N_12224);
nor U14096 (N_14096,N_11927,N_7880);
nand U14097 (N_14097,N_9551,N_7929);
xnor U14098 (N_14098,N_11972,N_11338);
xnor U14099 (N_14099,N_10556,N_11794);
and U14100 (N_14100,N_8002,N_11095);
xor U14101 (N_14101,N_6363,N_9378);
xor U14102 (N_14102,N_7841,N_8806);
xor U14103 (N_14103,N_7772,N_12283);
nand U14104 (N_14104,N_12156,N_10546);
and U14105 (N_14105,N_9372,N_7752);
nand U14106 (N_14106,N_10469,N_8472);
or U14107 (N_14107,N_11834,N_8370);
xor U14108 (N_14108,N_9966,N_11424);
nand U14109 (N_14109,N_11269,N_6898);
xnor U14110 (N_14110,N_7380,N_8242);
or U14111 (N_14111,N_10327,N_10047);
nand U14112 (N_14112,N_6923,N_7668);
nor U14113 (N_14113,N_8270,N_8711);
or U14114 (N_14114,N_10606,N_7094);
and U14115 (N_14115,N_9154,N_9590);
nand U14116 (N_14116,N_9132,N_8381);
nor U14117 (N_14117,N_6388,N_11853);
nand U14118 (N_14118,N_9668,N_10975);
xor U14119 (N_14119,N_6736,N_7449);
nor U14120 (N_14120,N_6849,N_11983);
nor U14121 (N_14121,N_11774,N_12128);
or U14122 (N_14122,N_10018,N_7650);
and U14123 (N_14123,N_12000,N_12383);
or U14124 (N_14124,N_8216,N_11103);
nand U14125 (N_14125,N_11658,N_7827);
xnor U14126 (N_14126,N_10704,N_11575);
nand U14127 (N_14127,N_8865,N_6952);
or U14128 (N_14128,N_12043,N_6560);
and U14129 (N_14129,N_8305,N_6287);
or U14130 (N_14130,N_11892,N_9478);
nand U14131 (N_14131,N_7910,N_11673);
and U14132 (N_14132,N_11078,N_12199);
or U14133 (N_14133,N_7411,N_12414);
or U14134 (N_14134,N_12048,N_11602);
or U14135 (N_14135,N_8727,N_9646);
or U14136 (N_14136,N_7850,N_12317);
xnor U14137 (N_14137,N_7976,N_8780);
nand U14138 (N_14138,N_9517,N_11837);
xnor U14139 (N_14139,N_11672,N_12017);
nor U14140 (N_14140,N_10348,N_7907);
nand U14141 (N_14141,N_11545,N_8555);
or U14142 (N_14142,N_12284,N_11874);
or U14143 (N_14143,N_8655,N_10578);
and U14144 (N_14144,N_11801,N_9103);
and U14145 (N_14145,N_9063,N_10978);
nor U14146 (N_14146,N_7497,N_11381);
nor U14147 (N_14147,N_11271,N_6520);
nand U14148 (N_14148,N_11828,N_7935);
xnor U14149 (N_14149,N_11657,N_8584);
nor U14150 (N_14150,N_10780,N_6549);
and U14151 (N_14151,N_12004,N_6537);
nand U14152 (N_14152,N_7630,N_11944);
or U14153 (N_14153,N_6796,N_6915);
xnor U14154 (N_14154,N_8830,N_8209);
nor U14155 (N_14155,N_7349,N_9926);
and U14156 (N_14156,N_7648,N_8537);
nor U14157 (N_14157,N_9056,N_11588);
nor U14158 (N_14158,N_11405,N_7701);
nand U14159 (N_14159,N_10366,N_10206);
or U14160 (N_14160,N_11159,N_10823);
and U14161 (N_14161,N_8072,N_7558);
xor U14162 (N_14162,N_11076,N_12386);
and U14163 (N_14163,N_8702,N_10000);
xor U14164 (N_14164,N_7805,N_10581);
or U14165 (N_14165,N_10334,N_6882);
nor U14166 (N_14166,N_12278,N_6358);
xor U14167 (N_14167,N_11380,N_6916);
nand U14168 (N_14168,N_7332,N_10940);
nor U14169 (N_14169,N_8160,N_7795);
nor U14170 (N_14170,N_11680,N_10127);
xnor U14171 (N_14171,N_8866,N_9290);
xnor U14172 (N_14172,N_6887,N_11428);
xor U14173 (N_14173,N_10298,N_6464);
xnor U14174 (N_14174,N_8137,N_10325);
nor U14175 (N_14175,N_7893,N_6930);
nor U14176 (N_14176,N_6657,N_11142);
nor U14177 (N_14177,N_10252,N_7045);
nor U14178 (N_14178,N_11937,N_8409);
nand U14179 (N_14179,N_6894,N_8193);
and U14180 (N_14180,N_8102,N_9722);
nand U14181 (N_14181,N_11621,N_10521);
xor U14182 (N_14182,N_11928,N_11242);
and U14183 (N_14183,N_10203,N_10755);
or U14184 (N_14184,N_8276,N_7079);
and U14185 (N_14185,N_11232,N_8717);
nor U14186 (N_14186,N_10765,N_9574);
xor U14187 (N_14187,N_11764,N_9039);
xnor U14188 (N_14188,N_8855,N_11557);
nand U14189 (N_14189,N_7525,N_10024);
nor U14190 (N_14190,N_11830,N_11438);
nor U14191 (N_14191,N_6484,N_6369);
nand U14192 (N_14192,N_11560,N_8701);
and U14193 (N_14193,N_7253,N_9538);
and U14194 (N_14194,N_6979,N_6695);
and U14195 (N_14195,N_11597,N_6381);
nand U14196 (N_14196,N_10422,N_9760);
xor U14197 (N_14197,N_10756,N_12375);
nand U14198 (N_14198,N_11347,N_11391);
nor U14199 (N_14199,N_11840,N_8117);
nand U14200 (N_14200,N_9899,N_11750);
nand U14201 (N_14201,N_11860,N_7389);
and U14202 (N_14202,N_6386,N_8969);
or U14203 (N_14203,N_7980,N_12329);
xnor U14204 (N_14204,N_9640,N_7023);
and U14205 (N_14205,N_7233,N_9976);
and U14206 (N_14206,N_12408,N_7337);
nor U14207 (N_14207,N_6600,N_12262);
nand U14208 (N_14208,N_6669,N_11518);
nor U14209 (N_14209,N_10081,N_6415);
nand U14210 (N_14210,N_12399,N_11703);
and U14211 (N_14211,N_9510,N_6517);
nand U14212 (N_14212,N_7593,N_10766);
xnor U14213 (N_14213,N_7776,N_8734);
nand U14214 (N_14214,N_7055,N_9789);
nor U14215 (N_14215,N_6316,N_7020);
or U14216 (N_14216,N_11999,N_7785);
xor U14217 (N_14217,N_6617,N_6623);
xor U14218 (N_14218,N_8148,N_8406);
and U14219 (N_14219,N_10917,N_10328);
xnor U14220 (N_14220,N_10486,N_6524);
or U14221 (N_14221,N_12275,N_8413);
nor U14222 (N_14222,N_6692,N_11297);
or U14223 (N_14223,N_10076,N_6832);
xor U14224 (N_14224,N_12242,N_6355);
and U14225 (N_14225,N_7859,N_9358);
xor U14226 (N_14226,N_6339,N_11160);
nand U14227 (N_14227,N_10192,N_6954);
xnor U14228 (N_14228,N_7172,N_6917);
xor U14229 (N_14229,N_10532,N_8881);
xor U14230 (N_14230,N_10145,N_8671);
and U14231 (N_14231,N_6398,N_7598);
nand U14232 (N_14232,N_8936,N_8268);
or U14233 (N_14233,N_11494,N_8604);
xnor U14234 (N_14234,N_10993,N_8770);
and U14235 (N_14235,N_8948,N_10205);
xor U14236 (N_14236,N_8475,N_8853);
nand U14237 (N_14237,N_7126,N_8680);
nor U14238 (N_14238,N_9140,N_7304);
or U14239 (N_14239,N_11210,N_9773);
or U14240 (N_14240,N_10636,N_8366);
or U14241 (N_14241,N_11616,N_8956);
nor U14242 (N_14242,N_6603,N_11779);
or U14243 (N_14243,N_10397,N_8870);
xnor U14244 (N_14244,N_10027,N_7664);
nand U14245 (N_14245,N_8499,N_12045);
and U14246 (N_14246,N_12467,N_12215);
nand U14247 (N_14247,N_12117,N_9975);
and U14248 (N_14248,N_12481,N_9183);
or U14249 (N_14249,N_6481,N_8369);
xor U14250 (N_14250,N_10258,N_7556);
and U14251 (N_14251,N_6500,N_8933);
or U14252 (N_14252,N_8217,N_10068);
xor U14253 (N_14253,N_10097,N_9681);
and U14254 (N_14254,N_7761,N_6607);
or U14255 (N_14255,N_10259,N_11989);
nand U14256 (N_14256,N_7934,N_11969);
nor U14257 (N_14257,N_8051,N_7532);
nor U14258 (N_14258,N_6795,N_6612);
nand U14259 (N_14259,N_11154,N_6277);
xor U14260 (N_14260,N_11685,N_8130);
nor U14261 (N_14261,N_8254,N_12202);
nor U14262 (N_14262,N_8076,N_7550);
nor U14263 (N_14263,N_7416,N_8061);
nand U14264 (N_14264,N_9242,N_11400);
or U14265 (N_14265,N_9978,N_9023);
or U14266 (N_14266,N_10083,N_7619);
and U14267 (N_14267,N_8271,N_11493);
or U14268 (N_14268,N_7022,N_10487);
and U14269 (N_14269,N_12225,N_10875);
or U14270 (N_14270,N_6551,N_11432);
nand U14271 (N_14271,N_6735,N_8813);
and U14272 (N_14272,N_10156,N_6329);
and U14273 (N_14273,N_11117,N_9072);
and U14274 (N_14274,N_12208,N_7146);
nand U14275 (N_14275,N_8379,N_7625);
nand U14276 (N_14276,N_12349,N_11280);
nand U14277 (N_14277,N_8388,N_11896);
xnor U14278 (N_14278,N_6350,N_6597);
and U14279 (N_14279,N_8637,N_6656);
or U14280 (N_14280,N_9155,N_11905);
and U14281 (N_14281,N_9586,N_7590);
or U14282 (N_14282,N_11912,N_8485);
or U14283 (N_14283,N_11050,N_6254);
or U14284 (N_14284,N_9506,N_8856);
and U14285 (N_14285,N_8529,N_8301);
nor U14286 (N_14286,N_6548,N_11754);
nor U14287 (N_14287,N_11675,N_10664);
nand U14288 (N_14288,N_8828,N_11317);
xor U14289 (N_14289,N_12161,N_8330);
nor U14290 (N_14290,N_7081,N_7970);
nand U14291 (N_14291,N_7830,N_9392);
and U14292 (N_14292,N_8787,N_9207);
and U14293 (N_14293,N_9296,N_9275);
and U14294 (N_14294,N_11327,N_9703);
or U14295 (N_14295,N_9370,N_10367);
nand U14296 (N_14296,N_6974,N_10794);
xnor U14297 (N_14297,N_6322,N_12104);
nor U14298 (N_14298,N_11663,N_6252);
or U14299 (N_14299,N_12211,N_8826);
nor U14300 (N_14300,N_6640,N_10319);
and U14301 (N_14301,N_11628,N_8018);
nor U14302 (N_14302,N_6718,N_9082);
xor U14303 (N_14303,N_7143,N_12271);
nor U14304 (N_14304,N_7727,N_10459);
nor U14305 (N_14305,N_8852,N_11712);
or U14306 (N_14306,N_11851,N_11043);
and U14307 (N_14307,N_8871,N_9701);
or U14308 (N_14308,N_6459,N_9927);
nand U14309 (N_14309,N_7257,N_8601);
or U14310 (N_14310,N_7184,N_6538);
nor U14311 (N_14311,N_10764,N_10154);
or U14312 (N_14312,N_9284,N_11101);
nand U14313 (N_14313,N_11092,N_12094);
nor U14314 (N_14314,N_7943,N_6900);
or U14315 (N_14315,N_10696,N_9452);
and U14316 (N_14316,N_11963,N_10429);
nand U14317 (N_14317,N_9017,N_7892);
xor U14318 (N_14318,N_10276,N_11348);
nand U14319 (N_14319,N_11516,N_11113);
xnor U14320 (N_14320,N_10112,N_7266);
nand U14321 (N_14321,N_10007,N_7206);
and U14322 (N_14322,N_7298,N_12387);
or U14323 (N_14323,N_9430,N_8685);
xnor U14324 (N_14324,N_9256,N_8896);
nor U14325 (N_14325,N_7197,N_6574);
xnor U14326 (N_14326,N_6604,N_7954);
xnor U14327 (N_14327,N_6696,N_9902);
and U14328 (N_14328,N_12264,N_8201);
nand U14329 (N_14329,N_12371,N_12253);
xor U14330 (N_14330,N_6993,N_7871);
nor U14331 (N_14331,N_7042,N_10485);
nand U14332 (N_14332,N_7942,N_11591);
nand U14333 (N_14333,N_8938,N_9785);
and U14334 (N_14334,N_7183,N_12195);
nor U14335 (N_14335,N_11445,N_7123);
or U14336 (N_14336,N_10798,N_8378);
nor U14337 (N_14337,N_8123,N_8146);
nor U14338 (N_14338,N_8197,N_8617);
nand U14339 (N_14339,N_12243,N_8836);
nand U14340 (N_14340,N_10607,N_12453);
or U14341 (N_14341,N_8940,N_9965);
and U14342 (N_14342,N_11815,N_9382);
nor U14343 (N_14343,N_12381,N_7690);
xnor U14344 (N_14344,N_9881,N_8493);
or U14345 (N_14345,N_7335,N_11273);
xor U14346 (N_14346,N_12311,N_12445);
or U14347 (N_14347,N_9961,N_10265);
nand U14348 (N_14348,N_9333,N_11325);
and U14349 (N_14349,N_11751,N_9026);
and U14350 (N_14350,N_9061,N_7672);
or U14351 (N_14351,N_6789,N_11510);
xnor U14352 (N_14352,N_10638,N_7413);
nand U14353 (N_14353,N_8465,N_8243);
or U14354 (N_14354,N_11722,N_8474);
and U14355 (N_14355,N_12079,N_8151);
nand U14356 (N_14356,N_12060,N_11541);
nand U14357 (N_14357,N_8422,N_8407);
nand U14358 (N_14358,N_9577,N_12353);
and U14359 (N_14359,N_11898,N_9129);
and U14360 (N_14360,N_10453,N_11455);
nor U14361 (N_14361,N_9373,N_10479);
nor U14362 (N_14362,N_11067,N_8352);
or U14363 (N_14363,N_7864,N_6835);
nand U14364 (N_14364,N_8912,N_10962);
or U14365 (N_14365,N_7026,N_6342);
xor U14366 (N_14366,N_7504,N_7017);
and U14367 (N_14367,N_11656,N_7732);
nand U14368 (N_14368,N_8367,N_11795);
or U14369 (N_14369,N_11827,N_8225);
nand U14370 (N_14370,N_10489,N_8503);
or U14371 (N_14371,N_11070,N_7602);
nand U14372 (N_14372,N_11195,N_8120);
or U14373 (N_14373,N_7480,N_10719);
and U14374 (N_14374,N_9038,N_8608);
and U14375 (N_14375,N_7862,N_8026);
or U14376 (N_14376,N_6305,N_9218);
nor U14377 (N_14377,N_7427,N_7498);
or U14378 (N_14378,N_10380,N_6991);
xnor U14379 (N_14379,N_11531,N_11199);
or U14380 (N_14380,N_8397,N_10912);
nor U14381 (N_14381,N_8234,N_8238);
xnor U14382 (N_14382,N_8848,N_10144);
or U14383 (N_14383,N_9856,N_10590);
and U14384 (N_14384,N_9387,N_10433);
or U14385 (N_14385,N_11084,N_7874);
nor U14386 (N_14386,N_6964,N_9341);
or U14387 (N_14387,N_7736,N_11949);
and U14388 (N_14388,N_7163,N_10960);
and U14389 (N_14389,N_12429,N_10474);
nand U14390 (N_14390,N_8908,N_11193);
and U14391 (N_14391,N_9159,N_10553);
or U14392 (N_14392,N_9541,N_12149);
or U14393 (N_14393,N_11568,N_9589);
and U14394 (N_14394,N_12459,N_9578);
xor U14395 (N_14395,N_10286,N_11702);
nor U14396 (N_14396,N_6935,N_7714);
or U14397 (N_14397,N_7120,N_11037);
nor U14398 (N_14398,N_9989,N_7228);
xnor U14399 (N_14399,N_10575,N_10566);
nor U14400 (N_14400,N_6689,N_9621);
xnor U14401 (N_14401,N_11841,N_8925);
or U14402 (N_14402,N_8447,N_8850);
nor U14403 (N_14403,N_9265,N_11571);
nor U14404 (N_14404,N_10966,N_12407);
xor U14405 (N_14405,N_11889,N_10098);
nand U14406 (N_14406,N_6790,N_9689);
nand U14407 (N_14407,N_9720,N_9637);
xnor U14408 (N_14408,N_10088,N_6934);
nor U14409 (N_14409,N_6728,N_11615);
or U14410 (N_14410,N_11505,N_12230);
xor U14411 (N_14411,N_8299,N_10828);
and U14412 (N_14412,N_11461,N_6253);
or U14413 (N_14413,N_8613,N_11483);
nor U14414 (N_14414,N_11328,N_10347);
nand U14415 (N_14415,N_9819,N_7173);
or U14416 (N_14416,N_8333,N_7443);
and U14417 (N_14417,N_7712,N_8074);
nand U14418 (N_14418,N_12410,N_11086);
nor U14419 (N_14419,N_8728,N_6946);
and U14420 (N_14420,N_6545,N_11371);
and U14421 (N_14421,N_11172,N_11468);
and U14422 (N_14422,N_6875,N_7911);
nor U14423 (N_14423,N_12050,N_9954);
or U14424 (N_14424,N_9416,N_6259);
and U14425 (N_14425,N_9163,N_10445);
and U14426 (N_14426,N_11360,N_6980);
nor U14427 (N_14427,N_11970,N_7739);
and U14428 (N_14428,N_11470,N_11633);
or U14429 (N_14429,N_11924,N_7494);
nor U14430 (N_14430,N_8999,N_6417);
nand U14431 (N_14431,N_11491,N_11635);
or U14432 (N_14432,N_9922,N_10131);
nor U14433 (N_14433,N_7496,N_8414);
or U14434 (N_14434,N_7471,N_11538);
and U14435 (N_14435,N_9613,N_6809);
and U14436 (N_14436,N_9083,N_8735);
and U14437 (N_14437,N_9000,N_9705);
xor U14438 (N_14438,N_7019,N_10599);
nor U14439 (N_14439,N_6311,N_7790);
nor U14440 (N_14440,N_8477,N_7232);
xnor U14441 (N_14441,N_7977,N_11419);
nand U14442 (N_14442,N_7655,N_7671);
or U14443 (N_14443,N_11796,N_12294);
and U14444 (N_14444,N_10946,N_7791);
nor U14445 (N_14445,N_12411,N_10342);
or U14446 (N_14446,N_10527,N_10829);
and U14447 (N_14447,N_10180,N_12187);
nor U14448 (N_14448,N_10497,N_10155);
nor U14449 (N_14449,N_8292,N_6430);
and U14450 (N_14450,N_7175,N_7052);
xor U14451 (N_14451,N_11885,N_7786);
nor U14452 (N_14452,N_7933,N_9277);
nor U14453 (N_14453,N_11274,N_12039);
nand U14454 (N_14454,N_9219,N_10787);
nor U14455 (N_14455,N_6390,N_9243);
nand U14456 (N_14456,N_8764,N_12018);
or U14457 (N_14457,N_10078,N_7723);
and U14458 (N_14458,N_8963,N_11661);
nor U14459 (N_14459,N_8738,N_7547);
nor U14460 (N_14460,N_6761,N_8753);
nor U14461 (N_14461,N_6702,N_8649);
and U14462 (N_14462,N_9174,N_9588);
nand U14463 (N_14463,N_8020,N_10204);
nand U14464 (N_14464,N_8223,N_11598);
or U14465 (N_14465,N_11206,N_6434);
and U14466 (N_14466,N_7492,N_11511);
or U14467 (N_14467,N_6719,N_8950);
or U14468 (N_14468,N_8986,N_6787);
and U14469 (N_14469,N_12047,N_9463);
nor U14470 (N_14470,N_6466,N_11329);
or U14471 (N_14471,N_9508,N_8982);
xnor U14472 (N_14472,N_9058,N_9921);
nor U14473 (N_14473,N_10307,N_9217);
and U14474 (N_14474,N_11838,N_11011);
xnor U14475 (N_14475,N_9125,N_11752);
nor U14476 (N_14476,N_11614,N_6333);
nand U14477 (N_14477,N_8625,N_7605);
xor U14478 (N_14478,N_7470,N_11267);
nor U14479 (N_14479,N_6995,N_9758);
nand U14480 (N_14480,N_11008,N_10311);
and U14481 (N_14481,N_12001,N_7870);
or U14482 (N_14482,N_7951,N_9180);
and U14483 (N_14483,N_8634,N_8844);
xor U14484 (N_14484,N_7158,N_11843);
nand U14485 (N_14485,N_10130,N_7311);
nand U14486 (N_14486,N_10233,N_10050);
and U14487 (N_14487,N_9923,N_9213);
xnor U14488 (N_14488,N_6553,N_9803);
and U14489 (N_14489,N_8937,N_11189);
nor U14490 (N_14490,N_8540,N_8803);
and U14491 (N_14491,N_6521,N_12037);
xor U14492 (N_14492,N_9592,N_7329);
and U14493 (N_14493,N_6361,N_9867);
or U14494 (N_14494,N_8487,N_6374);
xnor U14495 (N_14495,N_8822,N_10229);
and U14496 (N_14496,N_11250,N_7247);
nand U14497 (N_14497,N_7187,N_8513);
xor U14498 (N_14498,N_8591,N_6907);
xnor U14499 (N_14499,N_8528,N_8600);
nor U14500 (N_14500,N_9888,N_10997);
nand U14501 (N_14501,N_9157,N_7535);
or U14502 (N_14502,N_6955,N_12409);
and U14503 (N_14503,N_11361,N_7990);
nand U14504 (N_14504,N_8411,N_10594);
nand U14505 (N_14505,N_8122,N_9124);
and U14506 (N_14506,N_8147,N_7842);
xor U14507 (N_14507,N_9286,N_10729);
and U14508 (N_14508,N_10066,N_10818);
and U14509 (N_14509,N_12042,N_7710);
nor U14510 (N_14510,N_10141,N_10830);
xnor U14511 (N_14511,N_9756,N_7113);
and U14512 (N_14512,N_9727,N_11704);
and U14513 (N_14513,N_8854,N_7087);
nor U14514 (N_14514,N_9946,N_7048);
xor U14515 (N_14515,N_7782,N_8176);
xor U14516 (N_14516,N_10652,N_7810);
or U14517 (N_14517,N_10884,N_11045);
or U14518 (N_14518,N_10845,N_9117);
or U14519 (N_14519,N_11515,N_10107);
nor U14520 (N_14520,N_7209,N_7743);
or U14521 (N_14521,N_9285,N_11409);
xnor U14522 (N_14522,N_8052,N_6460);
nand U14523 (N_14523,N_8795,N_10657);
nand U14524 (N_14524,N_11223,N_10280);
or U14525 (N_14525,N_8260,N_10443);
nor U14526 (N_14526,N_10435,N_8079);
or U14527 (N_14527,N_10888,N_10690);
nor U14528 (N_14528,N_10354,N_9917);
nand U14529 (N_14529,N_11971,N_11316);
nor U14530 (N_14530,N_12364,N_7783);
nand U14531 (N_14531,N_6343,N_7722);
and U14532 (N_14532,N_11423,N_7179);
nand U14533 (N_14533,N_11553,N_7080);
nor U14534 (N_14534,N_7168,N_7813);
xor U14535 (N_14535,N_11649,N_11768);
nand U14536 (N_14536,N_7316,N_6384);
and U14537 (N_14537,N_12122,N_7258);
nor U14538 (N_14538,N_11141,N_10284);
nand U14539 (N_14539,N_10351,N_12030);
nand U14540 (N_14540,N_7180,N_8521);
xor U14541 (N_14541,N_11384,N_7583);
and U14542 (N_14542,N_8389,N_8706);
nand U14543 (N_14543,N_6871,N_9413);
xor U14544 (N_14544,N_8514,N_7041);
or U14545 (N_14545,N_7860,N_11059);
and U14546 (N_14546,N_12300,N_10303);
nor U14547 (N_14547,N_10604,N_9685);
nand U14548 (N_14548,N_7164,N_12351);
nand U14549 (N_14549,N_9555,N_10463);
and U14550 (N_14550,N_8841,N_6562);
xor U14551 (N_14551,N_10716,N_8014);
or U14552 (N_14552,N_11305,N_7755);
nor U14553 (N_14553,N_9271,N_12379);
or U14554 (N_14554,N_8887,N_8092);
nor U14555 (N_14555,N_7567,N_6602);
nand U14556 (N_14556,N_11960,N_10039);
xor U14557 (N_14557,N_7377,N_8502);
nand U14558 (N_14558,N_11865,N_8669);
and U14559 (N_14559,N_11418,N_9556);
xor U14560 (N_14560,N_12238,N_8972);
or U14561 (N_14561,N_11208,N_11052);
nand U14562 (N_14562,N_10115,N_7557);
xnor U14563 (N_14563,N_9766,N_9447);
xnor U14564 (N_14564,N_9102,N_8232);
nor U14565 (N_14565,N_9070,N_10153);
nand U14566 (N_14566,N_9844,N_7442);
or U14567 (N_14567,N_8250,N_9964);
nor U14568 (N_14568,N_9587,N_10222);
nor U14569 (N_14569,N_11061,N_7940);
and U14570 (N_14570,N_6713,N_7076);
nand U14571 (N_14571,N_7966,N_7399);
nor U14572 (N_14572,N_8280,N_10928);
nor U14573 (N_14573,N_10585,N_10706);
nand U14574 (N_14574,N_8606,N_9041);
or U14575 (N_14575,N_9963,N_6356);
nor U14576 (N_14576,N_8434,N_11177);
or U14577 (N_14577,N_6578,N_9068);
and U14578 (N_14578,N_11162,N_10509);
and U14579 (N_14579,N_10162,N_9349);
and U14580 (N_14580,N_6662,N_8991);
xnor U14581 (N_14581,N_8071,N_9828);
nor U14582 (N_14582,N_6412,N_8296);
or U14583 (N_14583,N_7930,N_10333);
nand U14584 (N_14584,N_10207,N_10119);
nor U14585 (N_14585,N_9861,N_10392);
or U14586 (N_14586,N_7728,N_10295);
or U14587 (N_14587,N_9048,N_10142);
nor U14588 (N_14588,N_11053,N_8721);
and U14589 (N_14589,N_7107,N_8597);
xor U14590 (N_14590,N_6863,N_7314);
nor U14591 (N_14591,N_10037,N_11771);
nor U14592 (N_14592,N_11648,N_7211);
nor U14593 (N_14593,N_7014,N_6471);
and U14594 (N_14594,N_8893,N_6794);
xor U14595 (N_14595,N_11462,N_7809);
nand U14596 (N_14596,N_12002,N_7364);
or U14597 (N_14597,N_10305,N_9938);
nand U14598 (N_14598,N_7563,N_11150);
xnor U14599 (N_14599,N_11880,N_7006);
and U14600 (N_14600,N_11953,N_10045);
or U14601 (N_14601,N_11090,N_9652);
or U14602 (N_14602,N_7771,N_8173);
nand U14603 (N_14603,N_10552,N_12466);
nor U14604 (N_14604,N_10434,N_7928);
nand U14605 (N_14605,N_11248,N_11604);
nand U14606 (N_14606,N_10231,N_8664);
and U14607 (N_14607,N_10642,N_10052);
nand U14608 (N_14608,N_9617,N_7271);
nor U14609 (N_14609,N_10574,N_11678);
nor U14610 (N_14610,N_11645,N_7474);
or U14611 (N_14611,N_8473,N_9420);
nor U14612 (N_14612,N_6686,N_9764);
xnor U14613 (N_14613,N_6786,N_10175);
nor U14614 (N_14614,N_10239,N_11623);
and U14615 (N_14615,N_12358,N_12166);
nand U14616 (N_14616,N_10714,N_7737);
xor U14617 (N_14617,N_7709,N_10439);
nor U14618 (N_14618,N_9278,N_8220);
and U14619 (N_14619,N_7596,N_6744);
and U14620 (N_14620,N_12058,N_12237);
or U14621 (N_14621,N_7564,N_12175);
or U14622 (N_14622,N_8785,N_10669);
or U14623 (N_14623,N_6704,N_10012);
xor U14624 (N_14624,N_11046,N_8460);
nor U14625 (N_14625,N_10949,N_7414);
xnor U14626 (N_14626,N_10738,N_9322);
and U14627 (N_14627,N_8437,N_6630);
or U14628 (N_14628,N_6938,N_11948);
nor U14629 (N_14629,N_10237,N_11562);
nand U14630 (N_14630,N_7130,N_9470);
and U14631 (N_14631,N_9569,N_8687);
or U14632 (N_14632,N_10492,N_10751);
nand U14633 (N_14633,N_8810,N_12463);
or U14634 (N_14634,N_11731,N_10383);
nor U14635 (N_14635,N_11203,N_8324);
nand U14636 (N_14636,N_7599,N_12163);
nand U14637 (N_14637,N_7454,N_11833);
and U14638 (N_14638,N_7836,N_10448);
nand U14639 (N_14639,N_7801,N_8275);
or U14640 (N_14640,N_8443,N_6528);
or U14641 (N_14641,N_12226,N_11577);
and U14642 (N_14642,N_6529,N_10999);
and U14643 (N_14643,N_9783,N_6555);
nor U14644 (N_14644,N_7568,N_6559);
xor U14645 (N_14645,N_10899,N_12204);
and U14646 (N_14646,N_11051,N_6519);
nand U14647 (N_14647,N_7611,N_9512);
and U14648 (N_14648,N_7101,N_6418);
or U14649 (N_14649,N_10084,N_7828);
xnor U14650 (N_14650,N_12158,N_7750);
nor U14651 (N_14651,N_7204,N_10136);
nand U14652 (N_14652,N_6996,N_7487);
or U14653 (N_14653,N_9659,N_10711);
and U14654 (N_14654,N_6541,N_6892);
or U14655 (N_14655,N_12151,N_7124);
nor U14656 (N_14656,N_6985,N_6468);
and U14657 (N_14657,N_8483,N_9435);
nor U14658 (N_14658,N_7348,N_10440);
and U14659 (N_14659,N_6511,N_9735);
xor U14660 (N_14660,N_8451,N_6821);
or U14661 (N_14661,N_10819,N_6439);
or U14662 (N_14662,N_7122,N_9616);
and U14663 (N_14663,N_11665,N_12137);
nand U14664 (N_14664,N_10152,N_10795);
or U14665 (N_14665,N_11429,N_8404);
xor U14666 (N_14666,N_6778,N_11932);
nand U14667 (N_14667,N_9992,N_8322);
and U14668 (N_14668,N_9252,N_9062);
xnor U14669 (N_14669,N_8784,N_12392);
nor U14670 (N_14670,N_6663,N_12120);
nand U14671 (N_14671,N_10123,N_11990);
xnor U14672 (N_14672,N_8440,N_9313);
nor U14673 (N_14673,N_8829,N_7756);
nor U14674 (N_14674,N_8112,N_9518);
nand U14675 (N_14675,N_8486,N_9415);
and U14676 (N_14676,N_9223,N_8949);
nor U14677 (N_14677,N_10164,N_8182);
nand U14678 (N_14678,N_9340,N_7624);
and U14679 (N_14679,N_8976,N_10644);
or U14680 (N_14680,N_9386,N_6325);
nor U14681 (N_14681,N_7780,N_10451);
xnor U14682 (N_14682,N_9221,N_7615);
xnor U14683 (N_14683,N_8030,N_7486);
or U14684 (N_14684,N_6525,N_8494);
and U14685 (N_14685,N_6442,N_11697);
nand U14686 (N_14686,N_8934,N_6845);
nor U14687 (N_14687,N_11524,N_8552);
or U14688 (N_14688,N_10177,N_10994);
nand U14689 (N_14689,N_7370,N_12170);
and U14690 (N_14690,N_7351,N_8757);
nor U14691 (N_14691,N_8740,N_10580);
nor U14692 (N_14692,N_9248,N_9303);
nand U14693 (N_14693,N_11619,N_7506);
xnor U14694 (N_14694,N_12069,N_11029);
nor U14695 (N_14695,N_10531,N_7660);
nor U14696 (N_14696,N_8507,N_9634);
nand U14697 (N_14697,N_12476,N_11512);
nand U14698 (N_14698,N_6793,N_9489);
nor U14699 (N_14699,N_11532,N_9693);
nand U14700 (N_14700,N_11606,N_9153);
nand U14701 (N_14701,N_10243,N_9886);
and U14702 (N_14702,N_8000,N_8003);
xor U14703 (N_14703,N_8624,N_11716);
or U14704 (N_14704,N_8394,N_6401);
nor U14705 (N_14705,N_8688,N_10430);
nand U14706 (N_14706,N_7210,N_8103);
xor U14707 (N_14707,N_10209,N_12206);
xor U14708 (N_14708,N_9399,N_7171);
nand U14709 (N_14709,N_9547,N_9485);
nor U14710 (N_14710,N_9568,N_9815);
nand U14711 (N_14711,N_8977,N_7387);
nand U14712 (N_14712,N_6586,N_6489);
or U14713 (N_14713,N_7293,N_10904);
xor U14714 (N_14714,N_9246,N_10717);
nor U14715 (N_14715,N_8777,N_9086);
and U14716 (N_14716,N_11564,N_8585);
and U14717 (N_14717,N_6687,N_8794);
xnor U14718 (N_14718,N_8253,N_11576);
or U14719 (N_14719,N_8978,N_8203);
nor U14720 (N_14720,N_11319,N_9596);
nor U14721 (N_14721,N_6667,N_8068);
or U14722 (N_14722,N_9245,N_10034);
nand U14723 (N_14723,N_9778,N_11302);
and U14724 (N_14724,N_10087,N_10374);
or U14725 (N_14725,N_10916,N_12401);
xor U14726 (N_14726,N_11243,N_9429);
nor U14727 (N_14727,N_9238,N_8943);
xnor U14728 (N_14728,N_12086,N_6677);
nand U14729 (N_14729,N_11175,N_9241);
nand U14730 (N_14730,N_12259,N_8206);
or U14731 (N_14731,N_8088,N_10848);
and U14732 (N_14732,N_6383,N_8723);
nor U14733 (N_14733,N_12289,N_11955);
xnor U14734 (N_14734,N_9189,N_9631);
and U14735 (N_14735,N_7324,N_7895);
or U14736 (N_14736,N_7779,N_10654);
or U14737 (N_14737,N_7587,N_6776);
or U14738 (N_14738,N_11723,N_9442);
and U14739 (N_14739,N_11283,N_6587);
xor U14740 (N_14740,N_8512,N_11759);
or U14741 (N_14741,N_9046,N_11145);
nand U14742 (N_14742,N_9203,N_9643);
nor U14743 (N_14743,N_10182,N_8539);
xnor U14744 (N_14744,N_10013,N_10520);
nand U14745 (N_14745,N_8050,N_10279);
nand U14746 (N_14746,N_12391,N_11372);
nor U14747 (N_14747,N_12203,N_9753);
or U14748 (N_14748,N_12477,N_8889);
xnor U14749 (N_14749,N_6473,N_11687);
nand U14750 (N_14750,N_8009,N_10031);
nand U14751 (N_14751,N_10090,N_10985);
nor U14752 (N_14752,N_8183,N_11200);
xnor U14753 (N_14753,N_7849,N_11954);
or U14754 (N_14754,N_11856,N_7576);
and U14755 (N_14755,N_6347,N_8772);
and U14756 (N_14756,N_9490,N_9604);
and U14757 (N_14757,N_6684,N_10114);
nor U14758 (N_14758,N_10318,N_6676);
nor U14759 (N_14759,N_10789,N_6542);
and U14760 (N_14760,N_9651,N_7448);
xnor U14761 (N_14761,N_8100,N_11938);
nor U14762 (N_14762,N_9460,N_12138);
nor U14763 (N_14763,N_7695,N_10111);
nor U14764 (N_14764,N_7974,N_10320);
nand U14765 (N_14765,N_11237,N_9328);
or U14766 (N_14766,N_10944,N_8548);
and U14767 (N_14767,N_9893,N_9920);
or U14768 (N_14768,N_10653,N_7015);
nor U14769 (N_14769,N_10673,N_7117);
xnor U14770 (N_14770,N_11721,N_8789);
nor U14771 (N_14771,N_10323,N_8628);
and U14772 (N_14772,N_8895,N_9095);
nand U14773 (N_14773,N_8782,N_8180);
nor U14774 (N_14774,N_6841,N_6791);
nand U14775 (N_14775,N_8725,N_7759);
and U14776 (N_14776,N_11042,N_9184);
nand U14777 (N_14777,N_7623,N_8975);
or U14778 (N_14778,N_6939,N_9324);
or U14779 (N_14779,N_8796,N_10800);
or U14780 (N_14780,N_10254,N_11064);
nand U14781 (N_14781,N_8800,N_10811);
nand U14782 (N_14782,N_10918,N_6975);
nor U14783 (N_14783,N_11699,N_11967);
or U14784 (N_14784,N_11033,N_9437);
and U14785 (N_14785,N_9827,N_11976);
or U14786 (N_14786,N_10238,N_10968);
or U14787 (N_14787,N_9906,N_12488);
nor U14788 (N_14788,N_9582,N_7078);
or U14789 (N_14789,N_10514,N_8269);
nor U14790 (N_14790,N_8273,N_11814);
nand U14791 (N_14791,N_7379,N_11331);
nand U14792 (N_14792,N_8010,N_11859);
xnor U14793 (N_14793,N_6474,N_8313);
or U14794 (N_14794,N_12279,N_8818);
or U14795 (N_14795,N_9024,N_11603);
and U14796 (N_14796,N_12403,N_10586);
or U14797 (N_14797,N_6910,N_6714);
nand U14798 (N_14798,N_9194,N_7301);
or U14799 (N_14799,N_8081,N_11939);
xnor U14800 (N_14800,N_11386,N_8992);
xnor U14801 (N_14801,N_7988,N_8927);
or U14802 (N_14802,N_7147,N_11770);
nand U14803 (N_14803,N_7327,N_7511);
nand U14804 (N_14804,N_10500,N_12038);
xor U14805 (N_14805,N_7857,N_9456);
nand U14806 (N_14806,N_10611,N_9110);
xor U14807 (N_14807,N_7358,N_12385);
xnor U14808 (N_14808,N_11030,N_8689);
xnor U14809 (N_14809,N_11112,N_7927);
nor U14810 (N_14810,N_8327,N_8345);
and U14811 (N_14811,N_10470,N_9564);
nand U14812 (N_14812,N_9121,N_9740);
nor U14813 (N_14813,N_11191,N_6757);
and U14814 (N_14814,N_7868,N_10077);
and U14815 (N_14815,N_8441,N_6561);
nand U14816 (N_14816,N_11140,N_8362);
nor U14817 (N_14817,N_7333,N_7798);
nand U14818 (N_14818,N_8684,N_11069);
xnor U14819 (N_14819,N_8586,N_9135);
xor U14820 (N_14820,N_9560,N_10852);
nor U14821 (N_14821,N_11426,N_6681);
nor U14822 (N_14822,N_7391,N_12297);
or U14823 (N_14823,N_11718,N_7083);
and U14824 (N_14824,N_6351,N_7754);
nor U14825 (N_14825,N_11187,N_7903);
xnor U14826 (N_14826,N_12496,N_10337);
nand U14827 (N_14827,N_6512,N_8426);
nand U14828 (N_14828,N_6326,N_8261);
or U14829 (N_14829,N_6962,N_8915);
or U14830 (N_14830,N_11773,N_8265);
or U14831 (N_14831,N_11878,N_7746);
and U14832 (N_14832,N_6409,N_7148);
or U14833 (N_14833,N_10855,N_10980);
nor U14834 (N_14834,N_11929,N_10650);
or U14835 (N_14835,N_11523,N_8094);
or U14836 (N_14836,N_7704,N_9381);
or U14837 (N_14837,N_10515,N_10982);
nand U14838 (N_14838,N_10862,N_11126);
nor U14839 (N_14839,N_10092,N_8153);
and U14840 (N_14840,N_10285,N_9557);
nand U14841 (N_14841,N_10562,N_8416);
xnor U14842 (N_14842,N_11707,N_9826);
xor U14843 (N_14843,N_8264,N_8663);
nand U14844 (N_14844,N_7119,N_11965);
xor U14845 (N_14845,N_8150,N_6348);
or U14846 (N_14846,N_8815,N_7601);
xnor U14847 (N_14847,N_8935,N_10568);
or U14848 (N_14848,N_6891,N_7639);
and U14849 (N_14849,N_9099,N_8427);
or U14850 (N_14850,N_10481,N_11652);
and U14851 (N_14851,N_8204,N_6803);
or U14852 (N_14852,N_12471,N_12116);
and U14853 (N_14853,N_6283,N_8775);
xor U14854 (N_14854,N_8210,N_7777);
nor U14855 (N_14855,N_9632,N_9425);
and U14856 (N_14856,N_6515,N_7626);
nand U14857 (N_14857,N_11062,N_8962);
xor U14858 (N_14858,N_12291,N_9383);
and U14859 (N_14859,N_10072,N_8323);
or U14860 (N_14860,N_12369,N_9860);
nor U14861 (N_14861,N_7826,N_9300);
nor U14862 (N_14862,N_9997,N_10926);
nand U14863 (N_14863,N_9424,N_10689);
or U14864 (N_14864,N_9800,N_8098);
nor U14865 (N_14865,N_9045,N_8241);
xor U14866 (N_14866,N_6652,N_9094);
nand U14867 (N_14867,N_7510,N_6615);
xnor U14868 (N_14868,N_11543,N_8208);
nand U14869 (N_14869,N_9250,N_10836);
xnor U14870 (N_14870,N_8904,N_9289);
and U14871 (N_14871,N_9004,N_10715);
nand U14872 (N_14872,N_8476,N_10734);
and U14873 (N_14873,N_8467,N_7027);
or U14874 (N_14874,N_11264,N_8931);
nand U14875 (N_14875,N_8257,N_12196);
nand U14876 (N_14876,N_9850,N_11032);
xor U14877 (N_14877,N_9970,N_7053);
xor U14878 (N_14878,N_8159,N_7426);
nand U14879 (N_14879,N_10880,N_11255);
nand U14880 (N_14880,N_10065,N_8168);
xor U14881 (N_14881,N_9986,N_6929);
or U14882 (N_14882,N_8154,N_6257);
xor U14883 (N_14883,N_8041,N_11471);
nor U14884 (N_14884,N_12160,N_12235);
or U14885 (N_14885,N_9877,N_11638);
nor U14886 (N_14886,N_7005,N_9305);
nand U14887 (N_14887,N_10996,N_7570);
or U14888 (N_14888,N_8924,N_10208);
and U14889 (N_14889,N_9433,N_9044);
or U14890 (N_14890,N_10762,N_8336);
xnor U14891 (N_14891,N_6732,N_8399);
or U14892 (N_14892,N_7959,N_8516);
nand U14893 (N_14893,N_7815,N_11985);
or U14894 (N_14894,N_6588,N_7846);
or U14895 (N_14895,N_11998,N_8876);
and U14896 (N_14896,N_9233,N_10567);
nand U14897 (N_14897,N_9916,N_7254);
and U14898 (N_14898,N_8044,N_10618);
and U14899 (N_14899,N_9692,N_7198);
and U14900 (N_14900,N_11108,N_8759);
and U14901 (N_14901,N_7306,N_11496);
nor U14902 (N_14902,N_9299,N_9791);
nand U14903 (N_14903,N_9545,N_9352);
and U14904 (N_14904,N_7579,N_12173);
nand U14905 (N_14905,N_8583,N_8731);
or U14906 (N_14906,N_7996,N_6275);
or U14907 (N_14907,N_9365,N_10057);
or U14908 (N_14908,N_12290,N_8382);
nand U14909 (N_14909,N_11858,N_7807);
and U14910 (N_14910,N_11301,N_11942);
nor U14911 (N_14911,N_11105,N_7855);
xnor U14912 (N_14912,N_9901,N_10006);
nor U14913 (N_14913,N_7073,N_10271);
nor U14914 (N_14914,N_11425,N_10160);
or U14915 (N_14915,N_11311,N_8851);
and U14916 (N_14916,N_8034,N_9338);
and U14917 (N_14917,N_8139,N_7423);
xnor U14918 (N_14918,N_10169,N_10813);
nand U14919 (N_14919,N_7967,N_9818);
nor U14920 (N_14920,N_7941,N_9627);
or U14921 (N_14921,N_8645,N_12465);
nand U14922 (N_14922,N_12172,N_10663);
or U14923 (N_14923,N_11996,N_11213);
nor U14924 (N_14924,N_11238,N_7285);
nand U14925 (N_14925,N_8054,N_11413);
or U14926 (N_14926,N_12483,N_11956);
xnor U14927 (N_14927,N_8101,N_11463);
nor U14928 (N_14928,N_7781,N_10682);
and U14929 (N_14929,N_10093,N_12281);
nand U14930 (N_14930,N_7201,N_6516);
or U14931 (N_14931,N_10403,N_7428);
and U14932 (N_14932,N_6606,N_8205);
and U14933 (N_14933,N_7667,N_10349);
xnor U14934 (N_14934,N_6294,N_9078);
nand U14935 (N_14935,N_7536,N_10049);
or U14936 (N_14936,N_10778,N_8221);
nand U14937 (N_14937,N_9438,N_10176);
nor U14938 (N_14938,N_7091,N_11873);
and U14939 (N_14939,N_9784,N_11821);
nand U14940 (N_14940,N_9910,N_7216);
nor U14941 (N_14941,N_9304,N_12121);
xor U14942 (N_14942,N_12266,N_8989);
xnor U14943 (N_14943,N_12293,N_7595);
nor U14944 (N_14944,N_11569,N_10959);
and U14945 (N_14945,N_9561,N_8069);
nand U14946 (N_14946,N_9137,N_8212);
and U14947 (N_14947,N_6759,N_6467);
nand U14948 (N_14948,N_8615,N_6425);
or U14949 (N_14949,N_6694,N_9454);
nor U14950 (N_14950,N_12485,N_6497);
xnor U14951 (N_14951,N_6755,N_10913);
nor U14952 (N_14952,N_7923,N_10900);
and U14953 (N_14953,N_6872,N_9660);
nor U14954 (N_14954,N_12197,N_11421);
nand U14955 (N_14955,N_9112,N_11798);
and U14956 (N_14956,N_12065,N_10266);
nor U14957 (N_14957,N_9546,N_9472);
and U14958 (N_14958,N_9019,N_7138);
xnor U14959 (N_14959,N_10675,N_7993);
or U14960 (N_14960,N_7863,N_8455);
xnor U14961 (N_14961,N_10598,N_9120);
xnor U14962 (N_14962,N_8861,N_11422);
xnor U14963 (N_14963,N_11058,N_11278);
or U14964 (N_14964,N_8418,N_8179);
nor U14965 (N_14965,N_8343,N_11003);
nand U14966 (N_14966,N_12064,N_10282);
and U14967 (N_14967,N_8007,N_6440);
or U14968 (N_14968,N_6319,N_10067);
nand U14969 (N_14969,N_7877,N_9465);
nor U14970 (N_14970,N_8174,N_12026);
and U14971 (N_14971,N_12148,N_8492);
nor U14972 (N_14972,N_12444,N_7691);
xnor U14973 (N_14973,N_9445,N_11477);
xor U14974 (N_14974,N_11355,N_11846);
or U14975 (N_14975,N_11075,N_9862);
xnor U14976 (N_14976,N_9990,N_6367);
nor U14977 (N_14977,N_9396,N_11777);
nor U14978 (N_14978,N_11085,N_11844);
or U14979 (N_14979,N_7975,N_9295);
nor U14980 (N_14980,N_6441,N_9173);
xor U14981 (N_14981,N_10188,N_11196);
nand U14982 (N_14982,N_8722,N_10376);
nand U14983 (N_14983,N_9109,N_8572);
nor U14984 (N_14984,N_11907,N_11152);
xor U14985 (N_14985,N_9550,N_10561);
or U14986 (N_14986,N_7099,N_10247);
nor U14987 (N_14987,N_10702,N_10512);
nor U14988 (N_14988,N_12352,N_7461);
nand U14989 (N_14989,N_9599,N_8913);
nand U14990 (N_14990,N_10406,N_6854);
and U14991 (N_14991,N_10074,N_8390);
and U14992 (N_14992,N_10625,N_10002);
or U14993 (N_14993,N_9868,N_8609);
or U14994 (N_14994,N_6861,N_10079);
nor U14995 (N_14995,N_7109,N_8229);
and U14996 (N_14996,N_8765,N_10350);
or U14997 (N_14997,N_11182,N_7627);
and U14998 (N_14998,N_8762,N_9814);
xor U14999 (N_14999,N_12019,N_8097);
nand U15000 (N_15000,N_8556,N_11440);
or U15001 (N_15001,N_12020,N_11902);
nor U15002 (N_15002,N_10214,N_9457);
and U15003 (N_15003,N_11850,N_9462);
or U15004 (N_15004,N_10249,N_10133);
nand U15005 (N_15005,N_11632,N_12333);
nor U15006 (N_15006,N_11570,N_11393);
or U15007 (N_15007,N_10721,N_9177);
and U15008 (N_15008,N_10091,N_6443);
or U15009 (N_15009,N_9636,N_6658);
and U15010 (N_15010,N_9981,N_8384);
nand U15011 (N_15011,N_9581,N_6806);
nand U15012 (N_15012,N_11321,N_9335);
xor U15013 (N_15013,N_8804,N_7522);
and U15014 (N_15014,N_9725,N_12440);
nor U15015 (N_15015,N_11031,N_10557);
and U15016 (N_15016,N_8312,N_7097);
nor U15017 (N_15017,N_8710,N_8055);
nor U15018 (N_15018,N_12372,N_9898);
nor U15019 (N_15019,N_10460,N_8917);
nor U15020 (N_15020,N_10379,N_9742);
and U15021 (N_15021,N_12218,N_7352);
nor U15022 (N_15022,N_11412,N_10810);
or U15023 (N_15023,N_11118,N_11861);
xor U15024 (N_15024,N_12078,N_7290);
nand U15025 (N_15025,N_9974,N_6873);
and U15026 (N_15026,N_9654,N_11852);
or U15027 (N_15027,N_9451,N_6614);
or U15028 (N_15028,N_6729,N_6816);
nor U15029 (N_15029,N_6903,N_8522);
and U15030 (N_15030,N_11442,N_8107);
nor U15031 (N_15031,N_7278,N_11914);
nor U15032 (N_15032,N_7214,N_12233);
and U15033 (N_15033,N_10086,N_10056);
nand U15034 (N_15034,N_12191,N_11746);
or U15035 (N_15035,N_8954,N_9677);
nor U15036 (N_15036,N_6948,N_6904);
or U15037 (N_15037,N_11906,N_11895);
nand U15038 (N_15038,N_6256,N_9334);
xnor U15039 (N_15039,N_11957,N_6613);
nand U15040 (N_15040,N_10868,N_7345);
or U15041 (N_15041,N_6317,N_10419);
or U15042 (N_15042,N_7885,N_11499);
xor U15043 (N_15043,N_7074,N_8213);
nor U15044 (N_15044,N_8133,N_8297);
nor U15045 (N_15045,N_6609,N_8040);
xnor U15046 (N_15046,N_10289,N_6285);
xor U15047 (N_15047,N_11408,N_11876);
or U15048 (N_15048,N_8347,N_12355);
nor U15049 (N_15049,N_11034,N_10688);
nand U15050 (N_15050,N_6715,N_11261);
nor U15051 (N_15051,N_11519,N_7242);
nand U15052 (N_15052,N_10157,N_6410);
nand U15053 (N_15053,N_8843,N_6986);
or U15054 (N_15054,N_9873,N_9739);
and U15055 (N_15055,N_6373,N_9658);
nor U15056 (N_15056,N_8247,N_7169);
nand U15057 (N_15057,N_11611,N_9461);
and U15058 (N_15058,N_9943,N_7395);
xor U15059 (N_15059,N_9967,N_10769);
and U15060 (N_15060,N_10300,N_7381);
xor U15061 (N_15061,N_9611,N_10457);
and U15062 (N_15062,N_10844,N_7475);
and U15063 (N_15063,N_9647,N_6312);
xnor U15064 (N_15064,N_7121,N_12141);
xor U15065 (N_15065,N_10995,N_10125);
and U15066 (N_15066,N_7127,N_9609);
xnor U15067 (N_15067,N_6897,N_11190);
nand U15068 (N_15068,N_11263,N_8504);
nand U15069 (N_15069,N_8929,N_10273);
nor U15070 (N_15070,N_11430,N_10898);
nand U15071 (N_15071,N_12499,N_6751);
and U15072 (N_15072,N_9380,N_8957);
nand U15073 (N_15073,N_9585,N_8175);
and U15074 (N_15074,N_8371,N_10693);
nand U15075 (N_15075,N_11456,N_10272);
xnor U15076 (N_15076,N_10595,N_6895);
nand U15077 (N_15077,N_10008,N_6433);
or U15078 (N_15078,N_10036,N_8236);
nor U15079 (N_15079,N_11530,N_9985);
nor U15080 (N_15080,N_8648,N_10967);
nor U15081 (N_15081,N_9377,N_7156);
and U15082 (N_15082,N_8910,N_6769);
nand U15083 (N_15083,N_7334,N_7634);
or U15084 (N_15084,N_6781,N_6950);
nand U15085 (N_15085,N_7061,N_6510);
xnor U15086 (N_15086,N_8501,N_11684);
and U15087 (N_15087,N_7355,N_9118);
and U15088 (N_15088,N_10742,N_7440);
or U15089 (N_15089,N_9754,N_6569);
or U15090 (N_15090,N_8121,N_7502);
and U15091 (N_15091,N_12055,N_11446);
xnor U15092 (N_15092,N_9389,N_9892);
or U15093 (N_15093,N_8858,N_10476);
xnor U15094 (N_15094,N_7260,N_9020);
nand U15095 (N_15095,N_11662,N_11509);
nor U15096 (N_15096,N_8295,N_6752);
xor U15097 (N_15097,N_9813,N_12003);
nand U15098 (N_15098,N_12454,N_11457);
and U15099 (N_15099,N_11574,N_12118);
or U15100 (N_15100,N_11745,N_10635);
or U15101 (N_15101,N_11188,N_7360);
and U15102 (N_15102,N_11936,N_8605);
nor U15103 (N_15103,N_9202,N_6659);
xor U15104 (N_15104,N_9255,N_8178);
nor U15105 (N_15105,N_9699,N_11308);
nand U15106 (N_15106,N_6354,N_9190);
xnor U15107 (N_15107,N_12011,N_9984);
nand U15108 (N_15108,N_11293,N_10761);
xnor U15109 (N_15109,N_9919,N_11816);
nor U15110 (N_15110,N_9166,N_9697);
or U15111 (N_15111,N_9371,N_10554);
and U15112 (N_15112,N_8444,N_11025);
or U15113 (N_15113,N_6625,N_7684);
or U15114 (N_15114,N_11812,N_9953);
nand U15115 (N_15115,N_10384,N_8105);
nand U15116 (N_15116,N_10840,N_6822);
xor U15117 (N_15117,N_8732,N_10896);
nor U15118 (N_15118,N_12015,N_9787);
nand U15119 (N_15119,N_7628,N_8833);
and U15120 (N_15120,N_11385,N_7200);
or U15121 (N_15121,N_12298,N_8281);
nor U15122 (N_15122,N_8008,N_6660);
xnor U15123 (N_15123,N_7307,N_11236);
and U15124 (N_15124,N_9563,N_6699);
xor U15125 (N_15125,N_7726,N_10046);
nor U15126 (N_15126,N_10432,N_8885);
and U15127 (N_15127,N_10357,N_9060);
and U15128 (N_15128,N_9771,N_12321);
xnor U15129 (N_15129,N_9113,N_8543);
or U15130 (N_15130,N_9852,N_12310);
and U15131 (N_15131,N_7499,N_8237);
nor U15132 (N_15132,N_10624,N_11819);
or U15133 (N_15133,N_7586,N_9914);
and U15134 (N_15134,N_12295,N_11158);
and U15135 (N_15135,N_11550,N_7114);
and U15136 (N_15136,N_10359,N_10950);
xor U15137 (N_15137,N_10686,N_12028);
xnor U15138 (N_15138,N_8337,N_7309);
nor U15139 (N_15139,N_12131,N_11094);
nand U15140 (N_15140,N_8027,N_12334);
nor U15141 (N_15141,N_9032,N_10873);
or U15142 (N_15142,N_6496,N_11625);
xor U15143 (N_15143,N_7429,N_12248);
nand U15144 (N_15144,N_12368,N_8471);
xor U15145 (N_15145,N_8488,N_7264);
or U15146 (N_15146,N_11689,N_11204);
nand U15147 (N_15147,N_12360,N_6721);
nor U15148 (N_15148,N_10746,N_11433);
or U15149 (N_15149,N_11073,N_9838);
or U15150 (N_15150,N_10874,N_11599);
or U15151 (N_15151,N_11690,N_8134);
xor U15152 (N_15152,N_7289,N_8979);
nand U15153 (N_15153,N_8754,N_11775);
or U15154 (N_15154,N_10023,N_10398);
nand U15155 (N_15155,N_9672,N_10294);
or U15156 (N_15156,N_8321,N_12446);
and U15157 (N_15157,N_6637,N_10071);
and U15158 (N_15158,N_11119,N_9292);
nor U15159 (N_15159,N_9071,N_7947);
or U15160 (N_15160,N_7299,N_8277);
nor U15161 (N_15161,N_6318,N_6703);
nor U15162 (N_15162,N_7902,N_10570);
nand U15163 (N_15163,N_7733,N_8062);
nor U15164 (N_15164,N_7814,N_11382);
or U15165 (N_15165,N_7526,N_10783);
nand U15166 (N_15166,N_7591,N_12092);
or U15167 (N_15167,N_7433,N_8651);
or U15168 (N_15168,N_12292,N_11125);
nand U15169 (N_15169,N_8812,N_8037);
xor U15170 (N_15170,N_7964,N_12250);
or U15171 (N_15171,N_6839,N_12302);
and U15172 (N_15172,N_6661,N_10369);
nand U15173 (N_15173,N_9853,N_8135);
or U15174 (N_15174,N_6302,N_9273);
or U15175 (N_15175,N_9247,N_11390);
xor U15176 (N_15176,N_8386,N_7955);
nand U15177 (N_15177,N_11127,N_9516);
and U15178 (N_15178,N_9776,N_11713);
nor U15179 (N_15179,N_9842,N_10768);
or U15180 (N_15180,N_6455,N_7581);
nand U15181 (N_15181,N_10179,N_6491);
xnor U15182 (N_15182,N_9504,N_6286);
xor U15183 (N_15183,N_9040,N_12176);
nor U15184 (N_15184,N_10760,N_9798);
or U15185 (N_15185,N_11556,N_9414);
xor U15186 (N_15186,N_9533,N_8798);
xnor U15187 (N_15187,N_9911,N_9079);
nand U15188 (N_15188,N_7075,N_9008);
or U15189 (N_15189,N_11388,N_10408);
nor U15190 (N_15190,N_10616,N_9263);
and U15191 (N_15191,N_7195,N_7488);
and U15192 (N_15192,N_11279,N_6501);
nor U15193 (N_15193,N_7421,N_11155);
or U15194 (N_15194,N_7192,N_8814);
and U15195 (N_15195,N_6530,N_8047);
and U15196 (N_15196,N_6334,N_7357);
and U15197 (N_15197,N_8868,N_10569);
nand U15198 (N_15198,N_10035,N_9534);
or U15199 (N_15199,N_7034,N_8677);
nand U15200 (N_15200,N_12424,N_11323);
and U15201 (N_15201,N_7758,N_7359);
nor U15202 (N_15202,N_8751,N_10517);
nor U15203 (N_15203,N_6595,N_9696);
and U15204 (N_15204,N_6436,N_8778);
xor U15205 (N_15205,N_9524,N_10718);
nand U15206 (N_15206,N_9022,N_12396);
or U15207 (N_15207,N_7678,N_7731);
and U15208 (N_15208,N_9635,N_6967);
and U15209 (N_15209,N_10895,N_12077);
or U15210 (N_15210,N_10882,N_8274);
and U15211 (N_15211,N_11941,N_8839);
and U15212 (N_15212,N_6404,N_10548);
and U15213 (N_15213,N_11444,N_7666);
nand U15214 (N_15214,N_8596,N_9719);
or U15215 (N_15215,N_6584,N_10314);
nor U15216 (N_15216,N_11862,N_11823);
or U15217 (N_15217,N_8085,N_11167);
nor U15218 (N_15218,N_8463,N_11186);
xor U15219 (N_15219,N_8057,N_10842);
nand U15220 (N_15220,N_6336,N_11919);
xnor U15221 (N_15221,N_8408,N_7946);
xnor U15222 (N_15222,N_9816,N_7058);
and U15223 (N_15223,N_11163,N_6402);
xor U15224 (N_15224,N_10197,N_10687);
nand U15225 (N_15225,N_7401,N_7376);
nor U15226 (N_15226,N_12382,N_6764);
or U15227 (N_15227,N_7606,N_8202);
or U15228 (N_15228,N_6937,N_11868);
or U15229 (N_15229,N_10363,N_10533);
or U15230 (N_15230,N_9486,N_12348);
xor U15231 (N_15231,N_9497,N_9913);
or U15232 (N_15232,N_8545,N_8398);
nand U15233 (N_15233,N_11601,N_7325);
xor U15234 (N_15234,N_8553,N_6303);
nor U15235 (N_15235,N_11682,N_12366);
nand U15236 (N_15236,N_11240,N_7585);
nand U15237 (N_15237,N_10637,N_8696);
nor U15238 (N_15238,N_8479,N_9156);
xor U15239 (N_15239,N_7222,N_10891);
xnor U15240 (N_15240,N_7629,N_7677);
nand U15241 (N_15241,N_6378,N_11356);
and U15242 (N_15242,N_9781,N_10069);
nor U15243 (N_15243,N_7989,N_12111);
nand U15244 (N_15244,N_7112,N_9211);
nand U15245 (N_15245,N_6896,N_12167);
or U15246 (N_15246,N_7665,N_9896);
xnor U15247 (N_15247,N_6701,N_10942);
or U15248 (N_15248,N_9571,N_7806);
nand U15249 (N_15249,N_9979,N_12378);
xor U15250 (N_15250,N_10423,N_6405);
xnor U15251 (N_15251,N_10902,N_7837);
nand U15252 (N_15252,N_6490,N_8480);
nand U15253 (N_15253,N_11241,N_7735);
nor U15254 (N_15254,N_8698,N_7654);
xor U15255 (N_15255,N_7111,N_7244);
or U15256 (N_15256,N_10146,N_8425);
nand U15257 (N_15257,N_6810,N_8736);
nand U15258 (N_15258,N_7418,N_6847);
and U15259 (N_15259,N_9894,N_11586);
nand U15260 (N_15260,N_9890,N_9522);
xor U15261 (N_15261,N_10970,N_6988);
or U15262 (N_15262,N_10804,N_8124);
or U15263 (N_15263,N_10251,N_7455);
and U15264 (N_15264,N_12434,N_7259);
nand U15265 (N_15265,N_10378,N_12192);
xnor U15266 (N_15266,N_9900,N_7177);
nor U15267 (N_15267,N_7068,N_8423);
nand U15268 (N_15268,N_6407,N_9319);
nor U15269 (N_15269,N_7011,N_8170);
nor U15270 (N_15270,N_11882,N_7089);
and U15271 (N_15271,N_12479,N_10353);
nor U15272 (N_15272,N_11641,N_9455);
xnor U15273 (N_15273,N_10626,N_10431);
nand U15274 (N_15274,N_7979,N_11973);
nor U15275 (N_15275,N_10161,N_10058);
xnor U15276 (N_15276,N_10105,N_7531);
nand U15277 (N_15277,N_6641,N_8763);
nand U15278 (N_15278,N_11719,N_8616);
and U15279 (N_15279,N_9362,N_10425);
or U15280 (N_15280,N_7981,N_12207);
or U15281 (N_15281,N_10306,N_9664);
nand U15282 (N_15282,N_12135,N_11875);
xor U15283 (N_15283,N_7539,N_7908);
nand U15284 (N_15284,N_6463,N_10986);
and U15285 (N_15285,N_11074,N_9721);
nand U15286 (N_15286,N_11460,N_9127);
nand U15287 (N_15287,N_8618,N_10776);
nor U15288 (N_15288,N_11529,N_7319);
and U15289 (N_15289,N_8820,N_7937);
and U15290 (N_15290,N_9354,N_7505);
nand U15291 (N_15291,N_10407,N_9228);
and U15292 (N_15292,N_11776,N_12258);
and U15293 (N_15293,N_11881,N_10791);
nand U15294 (N_15294,N_10166,N_12270);
xnor U15295 (N_15295,N_7295,N_11173);
nand U15296 (N_15296,N_8823,N_9134);
nor U15297 (N_15297,N_7509,N_9033);
nor U15298 (N_15298,N_11991,N_8665);
nor U15299 (N_15299,N_7203,N_9464);
nand U15300 (N_15300,N_10510,N_9947);
xor U15301 (N_15301,N_11149,N_8892);
xor U15302 (N_15302,N_8169,N_12428);
nand U15303 (N_15303,N_12344,N_7891);
and U15304 (N_15304,N_7310,N_10628);
nor U15305 (N_15305,N_7636,N_11544);
nand U15306 (N_15306,N_7270,N_7459);
nor U15307 (N_15307,N_8491,N_11201);
and U15308 (N_15308,N_11389,N_10150);
or U15309 (N_15309,N_6558,N_9169);
or U15310 (N_15310,N_6352,N_8758);
nor U15311 (N_15311,N_10805,N_10101);
xor U15312 (N_15312,N_7281,N_10480);
xnor U15313 (N_15313,N_7799,N_10167);
and U15314 (N_15314,N_6359,N_9915);
xor U15315 (N_15315,N_6758,N_10826);
xnor U15316 (N_15316,N_12316,N_6498);
and U15317 (N_15317,N_6777,N_9337);
or U15318 (N_15318,N_10674,N_11786);
and U15319 (N_15319,N_7751,N_8587);
nand U15320 (N_15320,N_6601,N_11931);
and U15321 (N_15321,N_8354,N_10541);
nor U15322 (N_15322,N_10929,N_11168);
xnor U15323 (N_15323,N_10513,N_6957);
or U15324 (N_15324,N_12252,N_10061);
and U15325 (N_15325,N_11452,N_9400);
nor U15326 (N_15326,N_9763,N_12087);
nand U15327 (N_15327,N_7104,N_10707);
xnor U15328 (N_15328,N_11959,N_10102);
or U15329 (N_15329,N_8968,N_6344);
nand U15330 (N_15330,N_10190,N_11009);
or U15331 (N_15331,N_11212,N_8527);
xnor U15332 (N_15332,N_10932,N_9126);
nor U15333 (N_15333,N_10936,N_10250);
xor U15334 (N_15334,N_11049,N_7724);
and U15335 (N_15335,N_10943,N_7221);
and U15336 (N_15336,N_8334,N_11353);
nand U15337 (N_15337,N_9718,N_7181);
and U15338 (N_15338,N_9749,N_7851);
and U15339 (N_15339,N_6665,N_11803);
xnor U15340 (N_15340,N_6649,N_10277);
nand U15341 (N_15341,N_7914,N_9093);
or U15342 (N_15342,N_6297,N_8457);
nand U15343 (N_15343,N_12347,N_11116);
xor U15344 (N_15344,N_10184,N_10385);
xnor U15345 (N_15345,N_8259,N_7150);
nand U15346 (N_15346,N_8141,N_10041);
nor U15347 (N_15347,N_7456,N_11836);
or U15348 (N_15348,N_10211,N_9175);
nor U15349 (N_15349,N_11185,N_11988);
nand U15350 (N_15350,N_6428,N_7009);
xnor U15351 (N_15351,N_7463,N_6332);
and U15352 (N_15352,N_10401,N_7582);
nand U15353 (N_15353,N_9653,N_12159);
or U15354 (N_15354,N_12257,N_10737);
or U15355 (N_15355,N_12213,N_11192);
or U15356 (N_15356,N_6438,N_10299);
or U15357 (N_15357,N_12110,N_6619);
or U15358 (N_15358,N_6983,N_8792);
nand U15359 (N_15359,N_6419,N_11292);
and U15360 (N_15360,N_6372,N_7145);
and U15361 (N_15361,N_11056,N_6622);
nand U15362 (N_15362,N_8110,N_8144);
or U15363 (N_15363,N_11272,N_9884);
xnor U15364 (N_15364,N_6567,N_9262);
and U15365 (N_15365,N_6893,N_9729);
and U15366 (N_15366,N_12126,N_7719);
and U15367 (N_15367,N_8682,N_10709);
xor U15368 (N_15368,N_6851,N_9944);
xor U15369 (N_15369,N_11732,N_10683);
or U15370 (N_15370,N_11100,N_10730);
nor U15371 (N_15371,N_9050,N_8207);
and U15372 (N_15372,N_11229,N_8136);
or U15373 (N_15373,N_9909,N_8233);
xnor U15374 (N_15374,N_10691,N_11900);
xor U15375 (N_15375,N_10171,N_9100);
and U15376 (N_15376,N_12460,N_9847);
nand U15377 (N_15377,N_7518,N_10952);
or U15378 (N_15378,N_10195,N_9805);
nand U15379 (N_15379,N_7300,N_11813);
or U15380 (N_15380,N_9307,N_7438);
nor U15381 (N_15381,N_10108,N_8638);
xnor U15382 (N_15382,N_10447,N_10542);
nor U15383 (N_15383,N_9765,N_9288);
nor U15384 (N_15384,N_12143,N_11443);
and U15385 (N_15385,N_12469,N_10656);
or U15386 (N_15386,N_11517,N_6488);
xor U15387 (N_15387,N_6831,N_6998);
xnor U15388 (N_15388,N_9142,N_10612);
nand U15389 (N_15389,N_8939,N_7059);
nand U15390 (N_15390,N_8080,N_8373);
xor U15391 (N_15391,N_7415,N_6672);
nand U15392 (N_15392,N_9075,N_10402);
or U15393 (N_15393,N_9179,N_10634);
or U15394 (N_15394,N_7013,N_9698);
nand U15395 (N_15395,N_12023,N_9931);
nand U15396 (N_15396,N_9988,N_8338);
xor U15397 (N_15397,N_10365,N_6726);
and U15398 (N_15398,N_9519,N_7764);
or U15399 (N_15399,N_7520,N_11166);
nor U15400 (N_15400,N_8857,N_8683);
or U15401 (N_15401,N_10198,N_6461);
nand U15402 (N_15402,N_11762,N_10321);
xnor U15403 (N_15403,N_11749,N_7507);
or U15404 (N_15404,N_9111,N_11359);
xor U15405 (N_15405,N_7215,N_10494);
xor U15406 (N_15406,N_9874,N_10727);
nand U15407 (N_15407,N_11992,N_12012);
nand U15408 (N_15408,N_6598,N_12498);
and U15409 (N_15409,N_12303,N_10713);
nand U15410 (N_15410,N_11218,N_10698);
or U15411 (N_15411,N_6494,N_10640);
or U15412 (N_15412,N_8713,N_9087);
or U15413 (N_15413,N_6688,N_9823);
xor U15414 (N_15414,N_8341,N_9405);
and U15415 (N_15415,N_9492,N_9049);
and U15416 (N_15416,N_7675,N_6295);
xnor U15417 (N_15417,N_8401,N_11298);
or U15418 (N_15418,N_8515,N_7328);
xnor U15419 (N_15419,N_11563,N_10441);
nand U15420 (N_15420,N_9200,N_9361);
nand U15421 (N_15421,N_10525,N_6921);
nor U15422 (N_15422,N_11879,N_7318);
nand U15423 (N_15423,N_8090,N_6580);
nand U15424 (N_15424,N_8712,N_8666);
nor U15425 (N_15425,N_10014,N_9885);
nor U15426 (N_15426,N_7924,N_7028);
or U15427 (N_15427,N_11735,N_8879);
or U15428 (N_15428,N_12301,N_11482);
xor U15429 (N_15429,N_6476,N_8981);
xnor U15430 (N_15430,N_8454,N_11724);
or U15431 (N_15431,N_8396,N_11324);
or U15432 (N_15432,N_8478,N_12374);
or U15433 (N_15433,N_6965,N_10317);
nand U15434 (N_15434,N_6638,N_11417);
xnor U15435 (N_15435,N_6395,N_10953);
xnor U15436 (N_15436,N_8449,N_7794);
xor U15437 (N_15437,N_6273,N_8190);
nand U15438 (N_15438,N_10808,N_6837);
xor U15439 (N_15439,N_8078,N_7250);
or U15440 (N_15440,N_8872,N_12005);
or U15441 (N_15441,N_10522,N_7544);
xnor U15442 (N_15442,N_10140,N_12337);
or U15443 (N_15443,N_8145,N_10417);
or U15444 (N_15444,N_6493,N_9015);
nor U15445 (N_15445,N_9757,N_9249);
nor U15446 (N_15446,N_6949,N_9258);
or U15447 (N_15447,N_7412,N_12098);
nor U15448 (N_15448,N_9507,N_9744);
xnor U15449 (N_15449,N_10831,N_9395);
or U15450 (N_15450,N_10796,N_8126);
nor U15451 (N_15451,N_6449,N_10503);
nor U15452 (N_15452,N_9737,N_7103);
and U15453 (N_15453,N_9831,N_8533);
xnor U15454 (N_15454,N_7584,N_6877);
nand U15455 (N_15455,N_8317,N_9593);
or U15456 (N_15456,N_9570,N_12096);
nor U15457 (N_15457,N_9552,N_11458);
nor U15458 (N_15458,N_12035,N_12280);
or U15459 (N_15459,N_6899,N_9671);
and U15460 (N_15460,N_12245,N_12027);
nor U15461 (N_15461,N_11940,N_10389);
and U15462 (N_15462,N_9628,N_9871);
nor U15463 (N_15463,N_11216,N_6522);
or U15464 (N_15464,N_9619,N_9481);
nand U15465 (N_15465,N_9065,N_9107);
and U15466 (N_15466,N_12201,N_8837);
xor U15467 (N_15467,N_6645,N_10444);
nand U15468 (N_15468,N_10837,N_7559);
nor U15469 (N_15469,N_9728,N_7725);
or U15470 (N_15470,N_11065,N_6710);
or U15471 (N_15471,N_10887,N_8368);
nor U15472 (N_15472,N_7432,N_7839);
nor U15473 (N_15473,N_10820,N_10499);
nor U15474 (N_15474,N_7082,N_10619);
and U15475 (N_15475,N_6675,N_10296);
nand U15476 (N_15476,N_7792,N_11832);
or U15477 (N_15477,N_11915,N_10302);
xnor U15478 (N_15478,N_12282,N_7362);
xnor U15479 (N_15479,N_7261,N_12112);
or U15480 (N_15480,N_11891,N_9991);
nand U15481 (N_15481,N_12066,N_10129);
nand U15482 (N_15482,N_9880,N_11231);
and U15483 (N_15483,N_8842,N_12346);
nand U15484 (N_15484,N_10931,N_6535);
or U15485 (N_15485,N_11738,N_12097);
nor U15486 (N_15486,N_9549,N_11630);
nand U15487 (N_15487,N_10371,N_10427);
xor U15488 (N_15488,N_8882,N_7225);
or U15489 (N_15489,N_8348,N_10839);
xnor U15490 (N_15490,N_8997,N_7283);
or U15491 (N_15491,N_8877,N_6583);
xnor U15492 (N_15492,N_9216,N_12057);
xnor U15493 (N_15493,N_9952,N_10538);
and U15494 (N_15494,N_8331,N_11980);
or U15495 (N_15495,N_10135,N_11785);
or U15496 (N_15496,N_6321,N_12210);
nand U15497 (N_15497,N_8967,N_9882);
xnor U15498 (N_15498,N_6534,N_11824);
or U15499 (N_15499,N_11257,N_9259);
nand U15500 (N_15500,N_6592,N_8140);
or U15501 (N_15501,N_11342,N_8138);
or U15502 (N_15502,N_9790,N_11387);
nand U15503 (N_15503,N_11805,N_6678);
nand U15504 (N_15504,N_8089,N_9797);
xnor U15505 (N_15505,N_9006,N_6919);
and U15506 (N_15506,N_11337,N_10324);
and U15507 (N_15507,N_11479,N_11521);
nor U15508 (N_15508,N_8901,N_7033);
or U15509 (N_15509,N_7115,N_9553);
or U15510 (N_15510,N_11258,N_8171);
and U15511 (N_15511,N_9509,N_8294);
and U15512 (N_15512,N_7000,N_12263);
nor U15513 (N_15513,N_7276,N_8004);
or U15514 (N_15514,N_8518,N_8084);
nand U15515 (N_15515,N_9186,N_9942);
nand U15516 (N_15516,N_6942,N_9956);
and U15517 (N_15517,N_9226,N_9440);
and U15518 (N_15518,N_6707,N_8163);
or U15519 (N_15519,N_10370,N_10555);
nand U15520 (N_15520,N_6947,N_9260);
and U15521 (N_15521,N_7757,N_11334);
and U15522 (N_15522,N_11454,N_9607);
nor U15523 (N_15523,N_7392,N_6953);
nand U15524 (N_15524,N_9605,N_12332);
xnor U15525 (N_15525,N_12288,N_9316);
nand U15526 (N_15526,N_11120,N_11792);
nor U15527 (N_15527,N_9164,N_9406);
xnor U15528 (N_15528,N_9679,N_8448);
or U15529 (N_15529,N_10109,N_9912);
nand U15530 (N_15530,N_10218,N_10516);
nor U15531 (N_15531,N_9573,N_7134);
nor U15532 (N_15532,N_9531,N_9935);
or U15533 (N_15533,N_7886,N_10352);
nor U15534 (N_15534,N_12155,N_7881);
nor U15535 (N_15535,N_6889,N_6862);
or U15536 (N_15536,N_8690,N_12025);
nor U15537 (N_15537,N_7770,N_10667);
nand U15538 (N_15538,N_7460,N_8300);
and U15539 (N_15539,N_9148,N_7165);
and U15540 (N_15540,N_7084,N_10473);
or U15541 (N_15541,N_9401,N_10793);
or U15542 (N_15542,N_12095,N_7468);
or U15543 (N_15543,N_6943,N_7622);
nand U15544 (N_15544,N_10919,N_11351);
nor U15545 (N_15545,N_7696,N_6627);
nand U15546 (N_15546,N_9746,N_9074);
xor U15547 (N_15547,N_12287,N_9133);
or U15548 (N_15548,N_10410,N_7823);
or U15549 (N_15549,N_7971,N_6576);
nor U15550 (N_15550,N_11831,N_9484);
xor U15551 (N_15551,N_10867,N_8571);
and U15552 (N_15552,N_9824,N_6834);
xnor U15553 (N_15553,N_9521,N_11642);
nand U15554 (N_15554,N_9806,N_6817);
xnor U15555 (N_15555,N_8724,N_8046);
nand U15556 (N_15556,N_8660,N_9320);
and U15557 (N_15557,N_11309,N_8965);
nand U15558 (N_15558,N_9829,N_12053);
and U15559 (N_15559,N_9630,N_12497);
nor U15560 (N_15560,N_11797,N_10748);
nor U15561 (N_15561,N_8200,N_11748);
and U15562 (N_15562,N_6444,N_10945);
nor U15563 (N_15563,N_12150,N_10712);
nand U15564 (N_15564,N_9332,N_6666);
xor U15565 (N_15565,N_8509,N_7425);
nand U15566 (N_15566,N_12341,N_7721);
xor U15567 (N_15567,N_9809,N_7607);
nand U15568 (N_15568,N_8285,N_10733);
xnor U15569 (N_15569,N_10981,N_8344);
xor U15570 (N_15570,N_11123,N_9673);
nand U15571 (N_15571,N_9080,N_7689);
xor U15572 (N_15572,N_9128,N_9196);
nor U15573 (N_15573,N_7693,N_12183);
or U15574 (N_15574,N_11952,N_8942);
nor U15575 (N_15575,N_9968,N_12040);
or U15576 (N_15576,N_12099,N_11789);
or U15577 (N_15577,N_7999,N_11378);
nand U15578 (N_15578,N_9875,N_10335);
and U15579 (N_15579,N_7938,N_9314);
nand U15580 (N_15580,N_8249,N_11767);
xor U15581 (N_15581,N_11143,N_9595);
xnor U15582 (N_15582,N_6618,N_6720);
nand U15583 (N_15583,N_6290,N_10740);
nor U15584 (N_15584,N_8436,N_11605);
nor U15585 (N_15585,N_8419,N_11739);
and U15586 (N_15586,N_12076,N_12214);
or U15587 (N_15587,N_7269,N_6848);
and U15588 (N_15588,N_6590,N_10817);
and U15589 (N_15589,N_11392,N_11079);
nor U15590 (N_15590,N_11701,N_10608);
nor U15591 (N_15591,N_12084,N_8284);
nor U15592 (N_15592,N_10292,N_11755);
nand U15593 (N_15593,N_9817,N_10671);
or U15594 (N_15594,N_12452,N_9670);
or U15595 (N_15595,N_9379,N_6801);
nand U15596 (N_15596,N_8566,N_6730);
nor U15597 (N_15597,N_9897,N_11930);
nand U15598 (N_15598,N_11613,N_12388);
or U15599 (N_15599,N_10297,N_9908);
nand U15600 (N_15600,N_7912,N_9001);
xnor U15601 (N_15601,N_11700,N_7390);
xor U15602 (N_15602,N_6426,N_7338);
nor U15603 (N_15603,N_8768,N_7464);
and U15604 (N_15604,N_6475,N_11753);
and U15605 (N_15605,N_6299,N_11644);
nor U15606 (N_15606,N_7640,N_8752);
nor U15607 (N_15607,N_9419,N_8359);
nand U15608 (N_15608,N_6994,N_9483);
xor U15609 (N_15609,N_9237,N_7267);
nor U15610 (N_15610,N_8224,N_6642);
and U15611 (N_15611,N_10054,N_10579);
and U15612 (N_15612,N_8429,N_11555);
and U15613 (N_15613,N_8043,N_12322);
or U15614 (N_15614,N_7056,N_7898);
or U15615 (N_15615,N_11335,N_7577);
and U15616 (N_15616,N_6536,N_10462);
and U15617 (N_15617,N_8550,N_6971);
nor U15618 (N_15618,N_9840,N_8860);
or U15619 (N_15619,N_6482,N_8032);
or U15620 (N_15620,N_7273,N_12177);
or U15621 (N_15621,N_6866,N_12441);
and U15622 (N_15622,N_7621,N_8658);
xnor U15623 (N_15623,N_7110,N_12109);
and U15624 (N_15624,N_8544,N_8561);
nor U15625 (N_15625,N_11616,N_6474);
and U15626 (N_15626,N_8309,N_8754);
nor U15627 (N_15627,N_10245,N_11528);
nor U15628 (N_15628,N_7997,N_10204);
or U15629 (N_15629,N_9013,N_10493);
nand U15630 (N_15630,N_6371,N_8353);
and U15631 (N_15631,N_6424,N_8159);
nand U15632 (N_15632,N_8275,N_6827);
nand U15633 (N_15633,N_7402,N_9397);
nor U15634 (N_15634,N_6975,N_10975);
nor U15635 (N_15635,N_10406,N_6774);
or U15636 (N_15636,N_11601,N_9414);
or U15637 (N_15637,N_8242,N_9740);
xor U15638 (N_15638,N_7392,N_7815);
nand U15639 (N_15639,N_9677,N_6311);
and U15640 (N_15640,N_10653,N_7956);
nand U15641 (N_15641,N_6597,N_9795);
nand U15642 (N_15642,N_11050,N_6508);
or U15643 (N_15643,N_11911,N_7783);
nor U15644 (N_15644,N_6548,N_10067);
nand U15645 (N_15645,N_8499,N_12037);
nand U15646 (N_15646,N_7744,N_9174);
or U15647 (N_15647,N_10368,N_11572);
or U15648 (N_15648,N_12124,N_12141);
or U15649 (N_15649,N_8489,N_6730);
xor U15650 (N_15650,N_6811,N_7999);
xnor U15651 (N_15651,N_6715,N_9474);
and U15652 (N_15652,N_10734,N_11833);
xnor U15653 (N_15653,N_11814,N_12443);
xor U15654 (N_15654,N_8654,N_12003);
or U15655 (N_15655,N_8974,N_9817);
xnor U15656 (N_15656,N_12287,N_7394);
nand U15657 (N_15657,N_6750,N_11155);
or U15658 (N_15658,N_9583,N_10261);
nand U15659 (N_15659,N_7962,N_7734);
nor U15660 (N_15660,N_9428,N_6953);
or U15661 (N_15661,N_7098,N_8072);
nor U15662 (N_15662,N_10688,N_10491);
or U15663 (N_15663,N_8687,N_8004);
or U15664 (N_15664,N_10378,N_9174);
nor U15665 (N_15665,N_7248,N_9653);
nand U15666 (N_15666,N_9969,N_6889);
nor U15667 (N_15667,N_7112,N_12028);
nor U15668 (N_15668,N_8383,N_12217);
xnor U15669 (N_15669,N_10863,N_11270);
and U15670 (N_15670,N_9986,N_7068);
nand U15671 (N_15671,N_7706,N_10630);
and U15672 (N_15672,N_8439,N_8314);
xnor U15673 (N_15673,N_10407,N_6646);
and U15674 (N_15674,N_7747,N_11209);
nor U15675 (N_15675,N_10263,N_9669);
or U15676 (N_15676,N_12070,N_9645);
nand U15677 (N_15677,N_8098,N_12216);
xor U15678 (N_15678,N_8170,N_10005);
or U15679 (N_15679,N_9352,N_7726);
nor U15680 (N_15680,N_6788,N_12485);
nor U15681 (N_15681,N_9315,N_7640);
and U15682 (N_15682,N_11039,N_9453);
xor U15683 (N_15683,N_6494,N_7756);
xnor U15684 (N_15684,N_10751,N_7741);
and U15685 (N_15685,N_9387,N_11970);
xnor U15686 (N_15686,N_9017,N_10446);
nor U15687 (N_15687,N_6848,N_9772);
nor U15688 (N_15688,N_8746,N_7260);
or U15689 (N_15689,N_9641,N_10656);
or U15690 (N_15690,N_11613,N_9262);
nor U15691 (N_15691,N_8121,N_8260);
nor U15692 (N_15692,N_10322,N_12036);
xor U15693 (N_15693,N_9285,N_8019);
nor U15694 (N_15694,N_8914,N_11426);
nand U15695 (N_15695,N_9980,N_7755);
nor U15696 (N_15696,N_9187,N_8619);
or U15697 (N_15697,N_8609,N_9858);
and U15698 (N_15698,N_12470,N_12474);
and U15699 (N_15699,N_9325,N_8450);
and U15700 (N_15700,N_10683,N_8662);
nor U15701 (N_15701,N_9729,N_10892);
or U15702 (N_15702,N_8376,N_7671);
nand U15703 (N_15703,N_8442,N_9374);
nand U15704 (N_15704,N_9291,N_7030);
nor U15705 (N_15705,N_10035,N_10421);
nand U15706 (N_15706,N_6573,N_10786);
and U15707 (N_15707,N_8535,N_7205);
or U15708 (N_15708,N_6504,N_8248);
nand U15709 (N_15709,N_9924,N_7373);
or U15710 (N_15710,N_10951,N_11968);
and U15711 (N_15711,N_11422,N_8496);
or U15712 (N_15712,N_8675,N_9556);
nor U15713 (N_15713,N_9807,N_11559);
xnor U15714 (N_15714,N_7240,N_9573);
and U15715 (N_15715,N_7218,N_9668);
and U15716 (N_15716,N_7052,N_8199);
or U15717 (N_15717,N_7712,N_10258);
or U15718 (N_15718,N_10300,N_9772);
xor U15719 (N_15719,N_7020,N_8703);
or U15720 (N_15720,N_11285,N_11249);
and U15721 (N_15721,N_11499,N_7076);
or U15722 (N_15722,N_6535,N_9523);
xor U15723 (N_15723,N_8905,N_10411);
and U15724 (N_15724,N_9849,N_11219);
nor U15725 (N_15725,N_6317,N_10744);
nor U15726 (N_15726,N_6438,N_11239);
xnor U15727 (N_15727,N_6989,N_10571);
nand U15728 (N_15728,N_6753,N_11629);
and U15729 (N_15729,N_9564,N_10677);
nand U15730 (N_15730,N_10845,N_12294);
nor U15731 (N_15731,N_7049,N_10885);
nand U15732 (N_15732,N_10183,N_6334);
nor U15733 (N_15733,N_8572,N_10379);
or U15734 (N_15734,N_9762,N_11442);
and U15735 (N_15735,N_8326,N_9694);
and U15736 (N_15736,N_9363,N_7380);
nor U15737 (N_15737,N_8645,N_8520);
and U15738 (N_15738,N_9583,N_6927);
or U15739 (N_15739,N_10583,N_10424);
and U15740 (N_15740,N_8342,N_11749);
or U15741 (N_15741,N_7370,N_10801);
or U15742 (N_15742,N_9272,N_9235);
and U15743 (N_15743,N_9425,N_7956);
and U15744 (N_15744,N_12389,N_6411);
or U15745 (N_15745,N_7559,N_12407);
or U15746 (N_15746,N_11534,N_9943);
nand U15747 (N_15747,N_8570,N_9882);
or U15748 (N_15748,N_8460,N_7612);
xor U15749 (N_15749,N_11584,N_8833);
nor U15750 (N_15750,N_12173,N_8810);
nor U15751 (N_15751,N_9228,N_10380);
xnor U15752 (N_15752,N_11326,N_11707);
or U15753 (N_15753,N_12494,N_11282);
or U15754 (N_15754,N_10768,N_12141);
or U15755 (N_15755,N_9507,N_8371);
or U15756 (N_15756,N_11037,N_6306);
nor U15757 (N_15757,N_9725,N_9394);
nand U15758 (N_15758,N_11351,N_11821);
xor U15759 (N_15759,N_6288,N_6657);
nor U15760 (N_15760,N_10301,N_6600);
nor U15761 (N_15761,N_6868,N_10556);
or U15762 (N_15762,N_10417,N_11448);
nand U15763 (N_15763,N_12043,N_9095);
xor U15764 (N_15764,N_7513,N_10100);
and U15765 (N_15765,N_12035,N_9952);
xor U15766 (N_15766,N_11281,N_7380);
or U15767 (N_15767,N_7735,N_10152);
nand U15768 (N_15768,N_9782,N_12441);
or U15769 (N_15769,N_7743,N_8176);
and U15770 (N_15770,N_10521,N_12423);
xor U15771 (N_15771,N_8543,N_6912);
nand U15772 (N_15772,N_10555,N_8789);
or U15773 (N_15773,N_6250,N_8279);
nand U15774 (N_15774,N_8474,N_8646);
xor U15775 (N_15775,N_7993,N_10649);
nor U15776 (N_15776,N_6586,N_8573);
or U15777 (N_15777,N_12499,N_6765);
or U15778 (N_15778,N_9434,N_12144);
nor U15779 (N_15779,N_12494,N_12429);
nor U15780 (N_15780,N_9922,N_9160);
nand U15781 (N_15781,N_8365,N_9916);
nor U15782 (N_15782,N_8406,N_10834);
nand U15783 (N_15783,N_11575,N_10328);
nand U15784 (N_15784,N_10735,N_10164);
or U15785 (N_15785,N_7297,N_7773);
and U15786 (N_15786,N_9285,N_9952);
xor U15787 (N_15787,N_6686,N_7409);
nand U15788 (N_15788,N_8959,N_9357);
nand U15789 (N_15789,N_10996,N_10187);
xnor U15790 (N_15790,N_6347,N_10061);
and U15791 (N_15791,N_10683,N_11059);
nand U15792 (N_15792,N_9439,N_8454);
nor U15793 (N_15793,N_9923,N_10236);
nor U15794 (N_15794,N_9622,N_10914);
nand U15795 (N_15795,N_10884,N_7655);
xnor U15796 (N_15796,N_8459,N_10479);
or U15797 (N_15797,N_6764,N_10591);
xnor U15798 (N_15798,N_10976,N_10500);
xor U15799 (N_15799,N_9264,N_7905);
nor U15800 (N_15800,N_9955,N_6331);
and U15801 (N_15801,N_8737,N_12180);
and U15802 (N_15802,N_10108,N_9020);
or U15803 (N_15803,N_6826,N_9101);
nand U15804 (N_15804,N_10024,N_11885);
or U15805 (N_15805,N_8499,N_7386);
or U15806 (N_15806,N_10438,N_10079);
nand U15807 (N_15807,N_12066,N_6424);
and U15808 (N_15808,N_8861,N_8484);
nand U15809 (N_15809,N_8663,N_7365);
nand U15810 (N_15810,N_11930,N_9008);
xnor U15811 (N_15811,N_7473,N_11063);
xor U15812 (N_15812,N_10314,N_8045);
or U15813 (N_15813,N_10054,N_6611);
and U15814 (N_15814,N_9488,N_7630);
nand U15815 (N_15815,N_6746,N_9960);
nor U15816 (N_15816,N_11349,N_9782);
nand U15817 (N_15817,N_12107,N_11769);
nand U15818 (N_15818,N_7959,N_7699);
xor U15819 (N_15819,N_7933,N_11359);
nand U15820 (N_15820,N_12355,N_9320);
and U15821 (N_15821,N_9941,N_10676);
nor U15822 (N_15822,N_8922,N_7863);
nand U15823 (N_15823,N_7647,N_11428);
xnor U15824 (N_15824,N_11767,N_8021);
nor U15825 (N_15825,N_7397,N_8478);
and U15826 (N_15826,N_8724,N_7686);
xnor U15827 (N_15827,N_7319,N_12032);
xor U15828 (N_15828,N_7916,N_7955);
and U15829 (N_15829,N_10722,N_10494);
xnor U15830 (N_15830,N_6582,N_9304);
xnor U15831 (N_15831,N_9518,N_8421);
and U15832 (N_15832,N_7466,N_10421);
and U15833 (N_15833,N_7920,N_11634);
xnor U15834 (N_15834,N_10403,N_11566);
nand U15835 (N_15835,N_12228,N_11835);
nor U15836 (N_15836,N_11910,N_9425);
nor U15837 (N_15837,N_6257,N_8142);
and U15838 (N_15838,N_7123,N_6664);
and U15839 (N_15839,N_12181,N_10289);
and U15840 (N_15840,N_8240,N_7860);
or U15841 (N_15841,N_10371,N_8788);
nand U15842 (N_15842,N_7541,N_12016);
and U15843 (N_15843,N_7913,N_6980);
and U15844 (N_15844,N_6318,N_12193);
or U15845 (N_15845,N_11978,N_9688);
xnor U15846 (N_15846,N_10359,N_7299);
nor U15847 (N_15847,N_11440,N_10636);
nor U15848 (N_15848,N_11473,N_10739);
xor U15849 (N_15849,N_9961,N_10834);
and U15850 (N_15850,N_11238,N_9486);
nand U15851 (N_15851,N_7252,N_12355);
xnor U15852 (N_15852,N_12026,N_10031);
and U15853 (N_15853,N_10213,N_11206);
nand U15854 (N_15854,N_6870,N_8227);
nor U15855 (N_15855,N_8491,N_8710);
xor U15856 (N_15856,N_9951,N_7518);
or U15857 (N_15857,N_11849,N_10421);
xor U15858 (N_15858,N_6822,N_11224);
and U15859 (N_15859,N_11424,N_7449);
or U15860 (N_15860,N_6734,N_7451);
xnor U15861 (N_15861,N_9361,N_7837);
nor U15862 (N_15862,N_6552,N_10775);
or U15863 (N_15863,N_8102,N_9025);
nand U15864 (N_15864,N_8054,N_8779);
nand U15865 (N_15865,N_12029,N_9538);
or U15866 (N_15866,N_12169,N_7916);
or U15867 (N_15867,N_10881,N_6321);
nor U15868 (N_15868,N_10239,N_9610);
and U15869 (N_15869,N_11717,N_6960);
nor U15870 (N_15870,N_11628,N_8693);
nand U15871 (N_15871,N_12229,N_6331);
nor U15872 (N_15872,N_8571,N_8515);
or U15873 (N_15873,N_8272,N_11149);
nand U15874 (N_15874,N_6792,N_6562);
or U15875 (N_15875,N_10453,N_8638);
and U15876 (N_15876,N_7057,N_10727);
nand U15877 (N_15877,N_7095,N_11987);
nand U15878 (N_15878,N_11096,N_10642);
xor U15879 (N_15879,N_9168,N_9493);
nand U15880 (N_15880,N_7406,N_7889);
xor U15881 (N_15881,N_6675,N_6947);
and U15882 (N_15882,N_7694,N_11433);
nand U15883 (N_15883,N_7888,N_10144);
xor U15884 (N_15884,N_9327,N_7446);
or U15885 (N_15885,N_9139,N_8527);
and U15886 (N_15886,N_8225,N_6941);
nor U15887 (N_15887,N_9920,N_8591);
nor U15888 (N_15888,N_7893,N_8395);
and U15889 (N_15889,N_7781,N_7982);
nand U15890 (N_15890,N_9737,N_7746);
nand U15891 (N_15891,N_11622,N_7508);
nand U15892 (N_15892,N_9245,N_7773);
nand U15893 (N_15893,N_7675,N_7589);
nor U15894 (N_15894,N_11962,N_7471);
and U15895 (N_15895,N_7269,N_10663);
nor U15896 (N_15896,N_9318,N_8546);
and U15897 (N_15897,N_10674,N_10997);
nand U15898 (N_15898,N_9107,N_9177);
xnor U15899 (N_15899,N_6480,N_9921);
or U15900 (N_15900,N_9440,N_11501);
and U15901 (N_15901,N_10991,N_11599);
nand U15902 (N_15902,N_8604,N_7033);
nor U15903 (N_15903,N_10233,N_8719);
nand U15904 (N_15904,N_6706,N_8603);
xor U15905 (N_15905,N_10797,N_6546);
or U15906 (N_15906,N_7678,N_8023);
and U15907 (N_15907,N_7245,N_9261);
xor U15908 (N_15908,N_9536,N_11291);
nor U15909 (N_15909,N_11928,N_7717);
nor U15910 (N_15910,N_12162,N_11897);
xor U15911 (N_15911,N_12482,N_10618);
xor U15912 (N_15912,N_8799,N_8374);
nor U15913 (N_15913,N_11785,N_8517);
and U15914 (N_15914,N_10480,N_9272);
nand U15915 (N_15915,N_8819,N_6544);
xnor U15916 (N_15916,N_7558,N_7825);
nor U15917 (N_15917,N_9132,N_9470);
nor U15918 (N_15918,N_9988,N_11428);
xor U15919 (N_15919,N_6359,N_9978);
or U15920 (N_15920,N_11083,N_10328);
or U15921 (N_15921,N_7179,N_9207);
xnor U15922 (N_15922,N_7434,N_8467);
and U15923 (N_15923,N_8655,N_9198);
and U15924 (N_15924,N_11560,N_8981);
nand U15925 (N_15925,N_9045,N_7962);
nand U15926 (N_15926,N_7691,N_8495);
nor U15927 (N_15927,N_7398,N_9992);
or U15928 (N_15928,N_10653,N_6782);
nand U15929 (N_15929,N_6415,N_6868);
nand U15930 (N_15930,N_8043,N_9198);
and U15931 (N_15931,N_11867,N_10903);
or U15932 (N_15932,N_9204,N_6623);
xor U15933 (N_15933,N_8056,N_6382);
nor U15934 (N_15934,N_7105,N_10821);
and U15935 (N_15935,N_12066,N_8630);
xnor U15936 (N_15936,N_8968,N_9744);
or U15937 (N_15937,N_11437,N_7895);
and U15938 (N_15938,N_8605,N_11070);
xnor U15939 (N_15939,N_8208,N_11370);
xor U15940 (N_15940,N_7331,N_10628);
nand U15941 (N_15941,N_11738,N_8002);
nor U15942 (N_15942,N_9664,N_6786);
or U15943 (N_15943,N_6403,N_10568);
or U15944 (N_15944,N_8747,N_11585);
nand U15945 (N_15945,N_7932,N_10610);
or U15946 (N_15946,N_12198,N_6934);
and U15947 (N_15947,N_8687,N_9062);
and U15948 (N_15948,N_11402,N_10574);
xnor U15949 (N_15949,N_6447,N_7077);
xnor U15950 (N_15950,N_7560,N_9316);
and U15951 (N_15951,N_12190,N_6325);
xnor U15952 (N_15952,N_9892,N_10553);
or U15953 (N_15953,N_12030,N_10857);
and U15954 (N_15954,N_9856,N_9072);
nor U15955 (N_15955,N_10614,N_10482);
nand U15956 (N_15956,N_10221,N_8215);
nand U15957 (N_15957,N_9534,N_11126);
xor U15958 (N_15958,N_7357,N_10923);
xnor U15959 (N_15959,N_12262,N_6393);
nor U15960 (N_15960,N_7861,N_6617);
nor U15961 (N_15961,N_6336,N_6356);
nand U15962 (N_15962,N_9356,N_11865);
xor U15963 (N_15963,N_6921,N_11295);
xnor U15964 (N_15964,N_10899,N_7648);
nand U15965 (N_15965,N_12354,N_10386);
and U15966 (N_15966,N_7840,N_6434);
xnor U15967 (N_15967,N_7254,N_8541);
and U15968 (N_15968,N_10687,N_11642);
or U15969 (N_15969,N_8609,N_6745);
nand U15970 (N_15970,N_12392,N_10528);
nor U15971 (N_15971,N_7869,N_9117);
nand U15972 (N_15972,N_8071,N_10433);
nand U15973 (N_15973,N_8489,N_10394);
xnor U15974 (N_15974,N_11223,N_7409);
nor U15975 (N_15975,N_7384,N_11033);
xnor U15976 (N_15976,N_9512,N_7739);
or U15977 (N_15977,N_8193,N_10888);
nand U15978 (N_15978,N_7906,N_10940);
or U15979 (N_15979,N_9219,N_8224);
nor U15980 (N_15980,N_11572,N_6864);
nor U15981 (N_15981,N_7977,N_12346);
nand U15982 (N_15982,N_11042,N_12054);
xor U15983 (N_15983,N_9472,N_8477);
xnor U15984 (N_15984,N_7263,N_12398);
and U15985 (N_15985,N_11527,N_12135);
xnor U15986 (N_15986,N_7036,N_7105);
or U15987 (N_15987,N_8738,N_11127);
nand U15988 (N_15988,N_11128,N_6451);
or U15989 (N_15989,N_10899,N_8917);
and U15990 (N_15990,N_6447,N_9229);
xor U15991 (N_15991,N_9097,N_11315);
nor U15992 (N_15992,N_9662,N_7696);
and U15993 (N_15993,N_6453,N_11706);
xnor U15994 (N_15994,N_6735,N_11669);
xnor U15995 (N_15995,N_11539,N_10475);
xnor U15996 (N_15996,N_7214,N_12004);
xor U15997 (N_15997,N_9064,N_10623);
and U15998 (N_15998,N_10628,N_8039);
xnor U15999 (N_15999,N_7663,N_9382);
or U16000 (N_16000,N_9832,N_12294);
nor U16001 (N_16001,N_12353,N_10522);
nand U16002 (N_16002,N_8276,N_11044);
and U16003 (N_16003,N_12017,N_9911);
xor U16004 (N_16004,N_11005,N_10773);
nor U16005 (N_16005,N_6537,N_10340);
xnor U16006 (N_16006,N_9099,N_11645);
xnor U16007 (N_16007,N_8926,N_8602);
xnor U16008 (N_16008,N_8007,N_9409);
and U16009 (N_16009,N_9103,N_11314);
nor U16010 (N_16010,N_9982,N_6603);
nor U16011 (N_16011,N_10388,N_11479);
xnor U16012 (N_16012,N_11526,N_9091);
xor U16013 (N_16013,N_11710,N_7527);
or U16014 (N_16014,N_6966,N_10357);
nor U16015 (N_16015,N_10782,N_11885);
xor U16016 (N_16016,N_7251,N_10402);
nand U16017 (N_16017,N_11450,N_12233);
or U16018 (N_16018,N_6622,N_10489);
nor U16019 (N_16019,N_12032,N_12201);
and U16020 (N_16020,N_7774,N_8989);
and U16021 (N_16021,N_9271,N_6250);
or U16022 (N_16022,N_10589,N_8722);
nor U16023 (N_16023,N_9282,N_7315);
and U16024 (N_16024,N_10592,N_7282);
nand U16025 (N_16025,N_11239,N_10684);
and U16026 (N_16026,N_9851,N_6649);
nor U16027 (N_16027,N_7928,N_10734);
or U16028 (N_16028,N_11506,N_6905);
nand U16029 (N_16029,N_11822,N_7459);
and U16030 (N_16030,N_6367,N_10377);
nand U16031 (N_16031,N_7705,N_7063);
nor U16032 (N_16032,N_10299,N_10991);
xor U16033 (N_16033,N_9930,N_10853);
nand U16034 (N_16034,N_12204,N_11442);
nand U16035 (N_16035,N_11150,N_8616);
and U16036 (N_16036,N_8726,N_11442);
and U16037 (N_16037,N_9689,N_7198);
nor U16038 (N_16038,N_11615,N_7452);
and U16039 (N_16039,N_6359,N_8345);
nor U16040 (N_16040,N_10841,N_8417);
nand U16041 (N_16041,N_12325,N_6393);
and U16042 (N_16042,N_8557,N_6289);
or U16043 (N_16043,N_10446,N_7531);
or U16044 (N_16044,N_8942,N_8393);
or U16045 (N_16045,N_10447,N_6438);
and U16046 (N_16046,N_6492,N_10269);
xor U16047 (N_16047,N_11782,N_6322);
nand U16048 (N_16048,N_6547,N_10723);
nand U16049 (N_16049,N_12338,N_9794);
or U16050 (N_16050,N_10254,N_11928);
nand U16051 (N_16051,N_8411,N_8346);
nor U16052 (N_16052,N_8177,N_8628);
and U16053 (N_16053,N_10209,N_10036);
nand U16054 (N_16054,N_10980,N_9354);
or U16055 (N_16055,N_10906,N_7496);
xor U16056 (N_16056,N_9088,N_7386);
and U16057 (N_16057,N_8548,N_11141);
nor U16058 (N_16058,N_10208,N_7796);
or U16059 (N_16059,N_9994,N_11638);
nor U16060 (N_16060,N_9400,N_8482);
or U16061 (N_16061,N_12109,N_9005);
nor U16062 (N_16062,N_12191,N_12249);
and U16063 (N_16063,N_11006,N_8147);
and U16064 (N_16064,N_8476,N_8016);
xor U16065 (N_16065,N_10932,N_9433);
and U16066 (N_16066,N_6813,N_9169);
nor U16067 (N_16067,N_6384,N_10490);
or U16068 (N_16068,N_11996,N_6563);
nand U16069 (N_16069,N_8824,N_12368);
xor U16070 (N_16070,N_9099,N_7902);
xnor U16071 (N_16071,N_9299,N_9613);
nor U16072 (N_16072,N_11037,N_7175);
xor U16073 (N_16073,N_11544,N_10037);
or U16074 (N_16074,N_10147,N_10507);
and U16075 (N_16075,N_7735,N_10240);
xnor U16076 (N_16076,N_12139,N_7671);
or U16077 (N_16077,N_11416,N_7427);
nor U16078 (N_16078,N_8701,N_12287);
or U16079 (N_16079,N_6607,N_9898);
or U16080 (N_16080,N_9611,N_8741);
nand U16081 (N_16081,N_8104,N_7013);
nand U16082 (N_16082,N_8622,N_11189);
and U16083 (N_16083,N_11019,N_10776);
xor U16084 (N_16084,N_9519,N_11253);
and U16085 (N_16085,N_11748,N_8639);
nand U16086 (N_16086,N_7057,N_8636);
and U16087 (N_16087,N_8629,N_8740);
or U16088 (N_16088,N_11721,N_7084);
or U16089 (N_16089,N_9425,N_9104);
and U16090 (N_16090,N_10685,N_8248);
nor U16091 (N_16091,N_9800,N_8712);
and U16092 (N_16092,N_7759,N_7571);
nand U16093 (N_16093,N_8348,N_10643);
and U16094 (N_16094,N_11968,N_7748);
nand U16095 (N_16095,N_8179,N_8127);
nor U16096 (N_16096,N_6671,N_8474);
nor U16097 (N_16097,N_8302,N_8386);
and U16098 (N_16098,N_7996,N_6571);
nor U16099 (N_16099,N_8000,N_6573);
nand U16100 (N_16100,N_9147,N_8082);
nor U16101 (N_16101,N_9622,N_12316);
nor U16102 (N_16102,N_7230,N_7045);
nand U16103 (N_16103,N_8979,N_6869);
or U16104 (N_16104,N_10766,N_12108);
and U16105 (N_16105,N_11613,N_8388);
or U16106 (N_16106,N_6911,N_9947);
and U16107 (N_16107,N_10251,N_12099);
nand U16108 (N_16108,N_10710,N_6989);
and U16109 (N_16109,N_11897,N_7917);
nand U16110 (N_16110,N_7872,N_9596);
and U16111 (N_16111,N_12072,N_11173);
and U16112 (N_16112,N_9760,N_7307);
xor U16113 (N_16113,N_10181,N_6888);
or U16114 (N_16114,N_11189,N_6453);
nor U16115 (N_16115,N_11820,N_10074);
xnor U16116 (N_16116,N_12000,N_7528);
xor U16117 (N_16117,N_9491,N_7691);
nand U16118 (N_16118,N_7803,N_6412);
nor U16119 (N_16119,N_11427,N_12134);
or U16120 (N_16120,N_7918,N_8847);
and U16121 (N_16121,N_10171,N_6472);
or U16122 (N_16122,N_8718,N_10760);
or U16123 (N_16123,N_7382,N_7579);
nor U16124 (N_16124,N_6948,N_9293);
nor U16125 (N_16125,N_9457,N_7739);
and U16126 (N_16126,N_11045,N_11988);
nand U16127 (N_16127,N_8074,N_6984);
xor U16128 (N_16128,N_7564,N_11433);
and U16129 (N_16129,N_7974,N_11549);
nor U16130 (N_16130,N_8792,N_9701);
xor U16131 (N_16131,N_7902,N_12170);
nand U16132 (N_16132,N_7688,N_9497);
nand U16133 (N_16133,N_11207,N_8107);
or U16134 (N_16134,N_10278,N_7132);
xor U16135 (N_16135,N_11426,N_11623);
or U16136 (N_16136,N_7341,N_6974);
or U16137 (N_16137,N_7385,N_10319);
or U16138 (N_16138,N_12140,N_9555);
nor U16139 (N_16139,N_7875,N_6633);
nor U16140 (N_16140,N_12368,N_7592);
xor U16141 (N_16141,N_9850,N_11569);
xnor U16142 (N_16142,N_9844,N_7161);
xnor U16143 (N_16143,N_10821,N_7167);
nand U16144 (N_16144,N_9868,N_12415);
or U16145 (N_16145,N_8491,N_11115);
or U16146 (N_16146,N_12372,N_9282);
and U16147 (N_16147,N_9067,N_7724);
or U16148 (N_16148,N_8627,N_12253);
and U16149 (N_16149,N_12044,N_10511);
nand U16150 (N_16150,N_6544,N_11897);
xnor U16151 (N_16151,N_11434,N_9311);
or U16152 (N_16152,N_10978,N_7378);
or U16153 (N_16153,N_11177,N_6909);
xnor U16154 (N_16154,N_11380,N_9521);
or U16155 (N_16155,N_6750,N_11930);
and U16156 (N_16156,N_6748,N_6499);
and U16157 (N_16157,N_6601,N_11952);
nand U16158 (N_16158,N_9288,N_11037);
nand U16159 (N_16159,N_6347,N_10773);
nor U16160 (N_16160,N_11881,N_9886);
nor U16161 (N_16161,N_10509,N_12271);
nand U16162 (N_16162,N_10409,N_6883);
xor U16163 (N_16163,N_9133,N_8091);
xnor U16164 (N_16164,N_11158,N_9206);
and U16165 (N_16165,N_11143,N_9607);
xnor U16166 (N_16166,N_11786,N_9636);
and U16167 (N_16167,N_12372,N_9788);
and U16168 (N_16168,N_6529,N_10604);
nor U16169 (N_16169,N_10185,N_7669);
xor U16170 (N_16170,N_9548,N_6311);
nor U16171 (N_16171,N_12351,N_6789);
xor U16172 (N_16172,N_10650,N_6910);
nor U16173 (N_16173,N_11980,N_8633);
nand U16174 (N_16174,N_10817,N_7181);
xnor U16175 (N_16175,N_9707,N_12396);
nand U16176 (N_16176,N_11967,N_10257);
and U16177 (N_16177,N_9168,N_7780);
nand U16178 (N_16178,N_7127,N_11490);
nand U16179 (N_16179,N_8550,N_12373);
nand U16180 (N_16180,N_9819,N_7811);
nand U16181 (N_16181,N_11951,N_9696);
or U16182 (N_16182,N_11495,N_9357);
xnor U16183 (N_16183,N_11853,N_7742);
nor U16184 (N_16184,N_12250,N_6383);
and U16185 (N_16185,N_11122,N_9874);
nand U16186 (N_16186,N_8439,N_8687);
or U16187 (N_16187,N_6855,N_8422);
and U16188 (N_16188,N_10400,N_10791);
xnor U16189 (N_16189,N_8349,N_11283);
and U16190 (N_16190,N_7830,N_12468);
nand U16191 (N_16191,N_8342,N_6610);
nor U16192 (N_16192,N_10490,N_11471);
and U16193 (N_16193,N_10694,N_10096);
nor U16194 (N_16194,N_7883,N_9034);
and U16195 (N_16195,N_11161,N_6884);
nand U16196 (N_16196,N_7833,N_9200);
xnor U16197 (N_16197,N_9130,N_10833);
or U16198 (N_16198,N_10916,N_8746);
and U16199 (N_16199,N_6287,N_7724);
or U16200 (N_16200,N_8686,N_11799);
and U16201 (N_16201,N_10899,N_12473);
nor U16202 (N_16202,N_7177,N_8279);
and U16203 (N_16203,N_11645,N_9789);
xor U16204 (N_16204,N_8202,N_10859);
nor U16205 (N_16205,N_6308,N_9816);
and U16206 (N_16206,N_9167,N_10193);
xnor U16207 (N_16207,N_10091,N_10283);
xor U16208 (N_16208,N_9614,N_10411);
and U16209 (N_16209,N_9059,N_10564);
and U16210 (N_16210,N_9136,N_10976);
xor U16211 (N_16211,N_10581,N_12319);
nand U16212 (N_16212,N_9661,N_8347);
nand U16213 (N_16213,N_7542,N_7707);
nor U16214 (N_16214,N_10207,N_8021);
xor U16215 (N_16215,N_12482,N_12472);
nand U16216 (N_16216,N_10085,N_11810);
or U16217 (N_16217,N_8973,N_12186);
and U16218 (N_16218,N_8277,N_10614);
and U16219 (N_16219,N_6690,N_6751);
and U16220 (N_16220,N_9309,N_10737);
or U16221 (N_16221,N_8630,N_10756);
nor U16222 (N_16222,N_8080,N_11321);
or U16223 (N_16223,N_12391,N_10214);
nand U16224 (N_16224,N_12024,N_9782);
nor U16225 (N_16225,N_12353,N_11841);
nand U16226 (N_16226,N_6958,N_12082);
or U16227 (N_16227,N_12094,N_6808);
nor U16228 (N_16228,N_7990,N_8681);
nand U16229 (N_16229,N_9877,N_10952);
or U16230 (N_16230,N_9287,N_11239);
and U16231 (N_16231,N_9453,N_8318);
or U16232 (N_16232,N_8069,N_6797);
nand U16233 (N_16233,N_6835,N_12286);
or U16234 (N_16234,N_11870,N_7872);
nand U16235 (N_16235,N_10741,N_8281);
and U16236 (N_16236,N_11442,N_9119);
and U16237 (N_16237,N_12079,N_12118);
nor U16238 (N_16238,N_10401,N_8714);
xor U16239 (N_16239,N_6273,N_10842);
nor U16240 (N_16240,N_11836,N_6809);
nand U16241 (N_16241,N_11663,N_11316);
nor U16242 (N_16242,N_9047,N_6434);
nand U16243 (N_16243,N_9104,N_8455);
or U16244 (N_16244,N_12114,N_11307);
nor U16245 (N_16245,N_6987,N_11366);
xor U16246 (N_16246,N_6314,N_8922);
or U16247 (N_16247,N_8201,N_11681);
or U16248 (N_16248,N_8947,N_11896);
xor U16249 (N_16249,N_6633,N_11038);
nor U16250 (N_16250,N_11787,N_12236);
or U16251 (N_16251,N_9753,N_10958);
nor U16252 (N_16252,N_10767,N_9919);
xnor U16253 (N_16253,N_12038,N_7456);
nor U16254 (N_16254,N_8798,N_10064);
nand U16255 (N_16255,N_8300,N_8159);
or U16256 (N_16256,N_9941,N_6965);
and U16257 (N_16257,N_11475,N_7769);
nor U16258 (N_16258,N_10477,N_6871);
nor U16259 (N_16259,N_12212,N_10013);
or U16260 (N_16260,N_11676,N_10051);
and U16261 (N_16261,N_11883,N_9939);
xor U16262 (N_16262,N_9386,N_6873);
nand U16263 (N_16263,N_8221,N_8098);
nand U16264 (N_16264,N_10860,N_8789);
or U16265 (N_16265,N_12119,N_9322);
nor U16266 (N_16266,N_11098,N_8969);
nor U16267 (N_16267,N_7541,N_8813);
xor U16268 (N_16268,N_10227,N_9469);
nor U16269 (N_16269,N_8863,N_6506);
nand U16270 (N_16270,N_9808,N_9227);
or U16271 (N_16271,N_7040,N_7840);
xor U16272 (N_16272,N_10459,N_10974);
nor U16273 (N_16273,N_11670,N_9453);
and U16274 (N_16274,N_10491,N_8122);
or U16275 (N_16275,N_12477,N_9294);
nand U16276 (N_16276,N_10654,N_8743);
nand U16277 (N_16277,N_11666,N_10632);
and U16278 (N_16278,N_8156,N_6773);
and U16279 (N_16279,N_8260,N_12203);
or U16280 (N_16280,N_10872,N_7735);
nor U16281 (N_16281,N_8104,N_6967);
and U16282 (N_16282,N_12332,N_7239);
or U16283 (N_16283,N_7850,N_7675);
and U16284 (N_16284,N_8812,N_7227);
or U16285 (N_16285,N_7719,N_9638);
xnor U16286 (N_16286,N_6401,N_8608);
xnor U16287 (N_16287,N_11780,N_12035);
nor U16288 (N_16288,N_9837,N_10508);
and U16289 (N_16289,N_10372,N_10175);
xnor U16290 (N_16290,N_7108,N_9611);
nand U16291 (N_16291,N_8296,N_6501);
nand U16292 (N_16292,N_8997,N_6896);
xnor U16293 (N_16293,N_10246,N_7564);
or U16294 (N_16294,N_9315,N_7207);
nor U16295 (N_16295,N_8551,N_12066);
nand U16296 (N_16296,N_6400,N_6520);
nor U16297 (N_16297,N_9615,N_8139);
xnor U16298 (N_16298,N_6834,N_6818);
or U16299 (N_16299,N_8324,N_9334);
nor U16300 (N_16300,N_7882,N_8261);
and U16301 (N_16301,N_10837,N_7883);
nand U16302 (N_16302,N_10672,N_6261);
xor U16303 (N_16303,N_10755,N_8157);
nand U16304 (N_16304,N_10361,N_12260);
and U16305 (N_16305,N_10170,N_11811);
or U16306 (N_16306,N_10951,N_9564);
nor U16307 (N_16307,N_10104,N_11021);
xnor U16308 (N_16308,N_7226,N_12192);
or U16309 (N_16309,N_10157,N_6351);
xnor U16310 (N_16310,N_8943,N_11420);
nand U16311 (N_16311,N_9058,N_11119);
nor U16312 (N_16312,N_7422,N_11755);
nor U16313 (N_16313,N_9359,N_8977);
nand U16314 (N_16314,N_7217,N_7958);
xor U16315 (N_16315,N_7373,N_12179);
xor U16316 (N_16316,N_8814,N_11157);
nand U16317 (N_16317,N_10943,N_11172);
nor U16318 (N_16318,N_11470,N_8394);
xor U16319 (N_16319,N_7405,N_7172);
nor U16320 (N_16320,N_10319,N_8103);
or U16321 (N_16321,N_10170,N_7013);
nand U16322 (N_16322,N_6993,N_10075);
or U16323 (N_16323,N_11769,N_10394);
or U16324 (N_16324,N_8089,N_7141);
or U16325 (N_16325,N_11028,N_10726);
or U16326 (N_16326,N_7011,N_8260);
and U16327 (N_16327,N_10595,N_10263);
nor U16328 (N_16328,N_9269,N_7019);
xnor U16329 (N_16329,N_8289,N_7384);
xor U16330 (N_16330,N_6956,N_7225);
nor U16331 (N_16331,N_8592,N_8605);
or U16332 (N_16332,N_7052,N_7236);
or U16333 (N_16333,N_12483,N_7420);
xor U16334 (N_16334,N_11402,N_9800);
and U16335 (N_16335,N_11083,N_12359);
and U16336 (N_16336,N_9283,N_9634);
xor U16337 (N_16337,N_9671,N_9672);
nand U16338 (N_16338,N_6839,N_9121);
and U16339 (N_16339,N_8998,N_10516);
or U16340 (N_16340,N_9342,N_9958);
nand U16341 (N_16341,N_7956,N_8794);
nor U16342 (N_16342,N_10655,N_11590);
or U16343 (N_16343,N_6957,N_10799);
xor U16344 (N_16344,N_11090,N_8976);
and U16345 (N_16345,N_12393,N_9390);
or U16346 (N_16346,N_6923,N_8518);
nand U16347 (N_16347,N_10822,N_9718);
or U16348 (N_16348,N_7549,N_6980);
nor U16349 (N_16349,N_8519,N_10288);
xnor U16350 (N_16350,N_8023,N_9360);
and U16351 (N_16351,N_8078,N_11017);
and U16352 (N_16352,N_6581,N_9362);
and U16353 (N_16353,N_9047,N_7049);
nand U16354 (N_16354,N_9531,N_10398);
nand U16355 (N_16355,N_8196,N_12368);
nor U16356 (N_16356,N_9751,N_7534);
nand U16357 (N_16357,N_6366,N_7708);
or U16358 (N_16358,N_9724,N_10334);
and U16359 (N_16359,N_8881,N_12227);
nand U16360 (N_16360,N_9656,N_11011);
and U16361 (N_16361,N_9094,N_11108);
nor U16362 (N_16362,N_7561,N_11177);
nor U16363 (N_16363,N_10344,N_12442);
nor U16364 (N_16364,N_12316,N_7119);
or U16365 (N_16365,N_8503,N_9954);
nor U16366 (N_16366,N_9148,N_9367);
nor U16367 (N_16367,N_9229,N_10778);
nor U16368 (N_16368,N_9921,N_7523);
xor U16369 (N_16369,N_7713,N_7837);
or U16370 (N_16370,N_11228,N_8361);
and U16371 (N_16371,N_10866,N_9704);
xor U16372 (N_16372,N_8407,N_6724);
nor U16373 (N_16373,N_7111,N_7129);
and U16374 (N_16374,N_10464,N_9651);
xnor U16375 (N_16375,N_10777,N_8868);
nand U16376 (N_16376,N_11164,N_11568);
nand U16377 (N_16377,N_6502,N_8009);
or U16378 (N_16378,N_10254,N_8720);
nand U16379 (N_16379,N_6271,N_11595);
nor U16380 (N_16380,N_10062,N_8235);
nor U16381 (N_16381,N_7591,N_11089);
xor U16382 (N_16382,N_11116,N_10642);
nand U16383 (N_16383,N_11364,N_7773);
nand U16384 (N_16384,N_6930,N_12435);
nor U16385 (N_16385,N_12250,N_6928);
or U16386 (N_16386,N_10610,N_12043);
and U16387 (N_16387,N_11493,N_7550);
and U16388 (N_16388,N_7276,N_7267);
xnor U16389 (N_16389,N_9988,N_6516);
nor U16390 (N_16390,N_6568,N_12068);
and U16391 (N_16391,N_9558,N_8879);
and U16392 (N_16392,N_10071,N_9132);
or U16393 (N_16393,N_12474,N_6264);
nand U16394 (N_16394,N_10771,N_9762);
nor U16395 (N_16395,N_9882,N_8990);
or U16396 (N_16396,N_8936,N_7496);
xor U16397 (N_16397,N_12138,N_11544);
xor U16398 (N_16398,N_10490,N_11636);
and U16399 (N_16399,N_11549,N_11656);
xor U16400 (N_16400,N_7917,N_9221);
nor U16401 (N_16401,N_7624,N_7434);
nand U16402 (N_16402,N_9940,N_11715);
or U16403 (N_16403,N_7017,N_7866);
xnor U16404 (N_16404,N_11060,N_11612);
nand U16405 (N_16405,N_10410,N_10062);
xnor U16406 (N_16406,N_12428,N_7976);
and U16407 (N_16407,N_11550,N_9170);
and U16408 (N_16408,N_8300,N_7639);
nand U16409 (N_16409,N_7428,N_12225);
nor U16410 (N_16410,N_8988,N_10276);
or U16411 (N_16411,N_8779,N_8590);
nor U16412 (N_16412,N_11828,N_11709);
nand U16413 (N_16413,N_8669,N_7999);
and U16414 (N_16414,N_6834,N_9082);
and U16415 (N_16415,N_10651,N_8432);
or U16416 (N_16416,N_9631,N_6752);
nor U16417 (N_16417,N_11923,N_9060);
nand U16418 (N_16418,N_11551,N_9203);
xnor U16419 (N_16419,N_12236,N_6308);
and U16420 (N_16420,N_9408,N_7408);
xor U16421 (N_16421,N_9078,N_6573);
xor U16422 (N_16422,N_6253,N_12142);
xnor U16423 (N_16423,N_11438,N_9332);
and U16424 (N_16424,N_7294,N_9057);
xor U16425 (N_16425,N_10532,N_8495);
nand U16426 (N_16426,N_9472,N_10348);
nand U16427 (N_16427,N_7121,N_8372);
xor U16428 (N_16428,N_9756,N_10616);
or U16429 (N_16429,N_11505,N_9593);
and U16430 (N_16430,N_12012,N_8673);
nand U16431 (N_16431,N_9608,N_10037);
nand U16432 (N_16432,N_8497,N_11021);
nand U16433 (N_16433,N_9240,N_6771);
nand U16434 (N_16434,N_10918,N_8692);
nor U16435 (N_16435,N_8540,N_9518);
or U16436 (N_16436,N_11498,N_6652);
nand U16437 (N_16437,N_6481,N_7763);
xor U16438 (N_16438,N_11486,N_10954);
nor U16439 (N_16439,N_7705,N_8804);
nand U16440 (N_16440,N_7539,N_9414);
nand U16441 (N_16441,N_8577,N_9125);
xnor U16442 (N_16442,N_10560,N_9280);
or U16443 (N_16443,N_9253,N_10965);
and U16444 (N_16444,N_6458,N_9363);
nand U16445 (N_16445,N_7601,N_8073);
xor U16446 (N_16446,N_10377,N_6472);
xnor U16447 (N_16447,N_6631,N_11520);
or U16448 (N_16448,N_9212,N_11875);
and U16449 (N_16449,N_10983,N_8907);
nand U16450 (N_16450,N_10256,N_10883);
or U16451 (N_16451,N_9961,N_9762);
xnor U16452 (N_16452,N_8752,N_11738);
nor U16453 (N_16453,N_10188,N_11818);
and U16454 (N_16454,N_8463,N_10723);
nand U16455 (N_16455,N_6715,N_9666);
or U16456 (N_16456,N_10674,N_10139);
nand U16457 (N_16457,N_6824,N_8076);
nor U16458 (N_16458,N_8916,N_10427);
nor U16459 (N_16459,N_11599,N_7494);
and U16460 (N_16460,N_10543,N_12057);
xnor U16461 (N_16461,N_9570,N_11897);
nor U16462 (N_16462,N_10688,N_11401);
xor U16463 (N_16463,N_9453,N_10916);
nand U16464 (N_16464,N_10146,N_10601);
or U16465 (N_16465,N_6736,N_7737);
or U16466 (N_16466,N_8812,N_11957);
and U16467 (N_16467,N_8861,N_7480);
or U16468 (N_16468,N_8805,N_10675);
nor U16469 (N_16469,N_8920,N_11699);
nor U16470 (N_16470,N_11213,N_10873);
nor U16471 (N_16471,N_11208,N_6516);
and U16472 (N_16472,N_8608,N_7132);
nor U16473 (N_16473,N_9578,N_11662);
xnor U16474 (N_16474,N_11905,N_10498);
xor U16475 (N_16475,N_10114,N_11642);
nand U16476 (N_16476,N_7876,N_7903);
nor U16477 (N_16477,N_10367,N_8727);
xor U16478 (N_16478,N_9385,N_6588);
xnor U16479 (N_16479,N_9520,N_11859);
nand U16480 (N_16480,N_8528,N_10057);
or U16481 (N_16481,N_10180,N_7031);
nor U16482 (N_16482,N_8798,N_11265);
xor U16483 (N_16483,N_7371,N_6262);
nor U16484 (N_16484,N_6712,N_11452);
or U16485 (N_16485,N_9340,N_10232);
xnor U16486 (N_16486,N_11510,N_8132);
nand U16487 (N_16487,N_10053,N_9971);
nor U16488 (N_16488,N_6585,N_12420);
or U16489 (N_16489,N_8587,N_7963);
or U16490 (N_16490,N_7344,N_9590);
or U16491 (N_16491,N_6607,N_9368);
or U16492 (N_16492,N_9088,N_11678);
nand U16493 (N_16493,N_7990,N_9554);
nand U16494 (N_16494,N_7888,N_9038);
or U16495 (N_16495,N_10163,N_12452);
nor U16496 (N_16496,N_7029,N_7073);
xor U16497 (N_16497,N_7230,N_10295);
xor U16498 (N_16498,N_12488,N_10312);
nand U16499 (N_16499,N_9471,N_8895);
and U16500 (N_16500,N_6823,N_6975);
xor U16501 (N_16501,N_7702,N_7416);
or U16502 (N_16502,N_9096,N_7795);
nor U16503 (N_16503,N_10050,N_11893);
and U16504 (N_16504,N_9558,N_11382);
nor U16505 (N_16505,N_11934,N_11348);
xnor U16506 (N_16506,N_9848,N_7639);
and U16507 (N_16507,N_10101,N_7296);
or U16508 (N_16508,N_8563,N_6347);
xor U16509 (N_16509,N_10379,N_9110);
or U16510 (N_16510,N_9728,N_8240);
nand U16511 (N_16511,N_9214,N_9881);
nor U16512 (N_16512,N_8068,N_11831);
or U16513 (N_16513,N_10995,N_8530);
or U16514 (N_16514,N_11947,N_8250);
and U16515 (N_16515,N_10343,N_8889);
xor U16516 (N_16516,N_10885,N_8711);
nor U16517 (N_16517,N_8493,N_11018);
or U16518 (N_16518,N_7314,N_12431);
xnor U16519 (N_16519,N_7041,N_7684);
or U16520 (N_16520,N_11921,N_7977);
xor U16521 (N_16521,N_12062,N_6372);
xor U16522 (N_16522,N_6623,N_11243);
nand U16523 (N_16523,N_10129,N_6494);
or U16524 (N_16524,N_7941,N_12334);
or U16525 (N_16525,N_11595,N_11453);
and U16526 (N_16526,N_7273,N_11592);
and U16527 (N_16527,N_11203,N_11195);
or U16528 (N_16528,N_9459,N_8714);
nand U16529 (N_16529,N_9722,N_9582);
xnor U16530 (N_16530,N_7412,N_9222);
or U16531 (N_16531,N_9428,N_9515);
nor U16532 (N_16532,N_11930,N_6487);
and U16533 (N_16533,N_9214,N_9552);
nor U16534 (N_16534,N_12116,N_6394);
or U16535 (N_16535,N_11135,N_6810);
and U16536 (N_16536,N_7392,N_7699);
and U16537 (N_16537,N_7988,N_12394);
or U16538 (N_16538,N_7126,N_9371);
xnor U16539 (N_16539,N_8861,N_11003);
xnor U16540 (N_16540,N_9191,N_8676);
and U16541 (N_16541,N_9451,N_10102);
or U16542 (N_16542,N_8438,N_11129);
nand U16543 (N_16543,N_9431,N_9277);
nor U16544 (N_16544,N_9266,N_7130);
xor U16545 (N_16545,N_7489,N_9763);
nand U16546 (N_16546,N_9308,N_8527);
and U16547 (N_16547,N_6869,N_12226);
xor U16548 (N_16548,N_9187,N_9724);
and U16549 (N_16549,N_7860,N_10306);
or U16550 (N_16550,N_11187,N_7571);
nor U16551 (N_16551,N_12297,N_11717);
xor U16552 (N_16552,N_11258,N_7829);
and U16553 (N_16553,N_9390,N_11202);
and U16554 (N_16554,N_7491,N_12225);
nand U16555 (N_16555,N_9605,N_10566);
xor U16556 (N_16556,N_9463,N_9935);
or U16557 (N_16557,N_11890,N_6725);
xor U16558 (N_16558,N_7043,N_12333);
xnor U16559 (N_16559,N_8508,N_6685);
nand U16560 (N_16560,N_7445,N_9036);
and U16561 (N_16561,N_11585,N_8576);
and U16562 (N_16562,N_6559,N_7708);
xor U16563 (N_16563,N_9913,N_8810);
nand U16564 (N_16564,N_12076,N_8686);
nor U16565 (N_16565,N_9120,N_8306);
xor U16566 (N_16566,N_12255,N_10954);
nand U16567 (N_16567,N_8176,N_11511);
and U16568 (N_16568,N_8939,N_8355);
nor U16569 (N_16569,N_9795,N_8903);
nor U16570 (N_16570,N_9752,N_7878);
and U16571 (N_16571,N_9250,N_10890);
or U16572 (N_16572,N_11610,N_9740);
xnor U16573 (N_16573,N_11397,N_10362);
nor U16574 (N_16574,N_10645,N_6789);
and U16575 (N_16575,N_7703,N_12009);
nor U16576 (N_16576,N_6583,N_10500);
nand U16577 (N_16577,N_9504,N_8498);
xnor U16578 (N_16578,N_8968,N_7133);
xnor U16579 (N_16579,N_12138,N_12339);
xor U16580 (N_16580,N_7045,N_9729);
nor U16581 (N_16581,N_9031,N_10925);
nand U16582 (N_16582,N_8657,N_12149);
or U16583 (N_16583,N_7089,N_9000);
xnor U16584 (N_16584,N_7992,N_8900);
xnor U16585 (N_16585,N_9960,N_12290);
and U16586 (N_16586,N_7301,N_7173);
xor U16587 (N_16587,N_10821,N_8801);
or U16588 (N_16588,N_6351,N_9383);
or U16589 (N_16589,N_8189,N_7146);
and U16590 (N_16590,N_10247,N_6610);
and U16591 (N_16591,N_10448,N_6253);
xnor U16592 (N_16592,N_9097,N_9533);
and U16593 (N_16593,N_11700,N_6595);
xor U16594 (N_16594,N_6713,N_7081);
or U16595 (N_16595,N_7294,N_12024);
nor U16596 (N_16596,N_10597,N_7540);
nor U16597 (N_16597,N_6447,N_11774);
nor U16598 (N_16598,N_7849,N_10967);
xnor U16599 (N_16599,N_8680,N_8281);
nor U16600 (N_16600,N_11914,N_8347);
xnor U16601 (N_16601,N_7236,N_9686);
or U16602 (N_16602,N_7872,N_9545);
and U16603 (N_16603,N_9537,N_11558);
or U16604 (N_16604,N_10060,N_9457);
and U16605 (N_16605,N_8248,N_10884);
nor U16606 (N_16606,N_11821,N_8024);
nor U16607 (N_16607,N_12425,N_9946);
xor U16608 (N_16608,N_7260,N_10369);
or U16609 (N_16609,N_12408,N_9728);
or U16610 (N_16610,N_8288,N_12095);
nor U16611 (N_16611,N_7539,N_10061);
or U16612 (N_16612,N_8037,N_7925);
nand U16613 (N_16613,N_11274,N_12247);
nand U16614 (N_16614,N_10574,N_7541);
nor U16615 (N_16615,N_12230,N_6385);
and U16616 (N_16616,N_8410,N_7455);
or U16617 (N_16617,N_7627,N_9713);
nor U16618 (N_16618,N_9404,N_8609);
nand U16619 (N_16619,N_9244,N_10229);
or U16620 (N_16620,N_9494,N_11381);
and U16621 (N_16621,N_12441,N_8797);
and U16622 (N_16622,N_12381,N_11216);
xnor U16623 (N_16623,N_9799,N_7365);
or U16624 (N_16624,N_9493,N_7979);
or U16625 (N_16625,N_12102,N_8285);
and U16626 (N_16626,N_11107,N_12080);
nor U16627 (N_16627,N_7569,N_9017);
nand U16628 (N_16628,N_8599,N_8764);
xnor U16629 (N_16629,N_9738,N_9526);
xnor U16630 (N_16630,N_6771,N_6521);
xor U16631 (N_16631,N_9882,N_7992);
and U16632 (N_16632,N_11230,N_8192);
xnor U16633 (N_16633,N_7210,N_7765);
or U16634 (N_16634,N_9931,N_6764);
or U16635 (N_16635,N_8332,N_11917);
or U16636 (N_16636,N_9821,N_10335);
nor U16637 (N_16637,N_10631,N_9525);
and U16638 (N_16638,N_11051,N_8668);
or U16639 (N_16639,N_6653,N_6649);
xor U16640 (N_16640,N_10394,N_10237);
or U16641 (N_16641,N_8558,N_9232);
nand U16642 (N_16642,N_8016,N_10387);
xnor U16643 (N_16643,N_6943,N_6835);
nor U16644 (N_16644,N_7793,N_9055);
nor U16645 (N_16645,N_12027,N_7352);
nor U16646 (N_16646,N_6566,N_8679);
xor U16647 (N_16647,N_8456,N_10468);
or U16648 (N_16648,N_8134,N_11705);
nand U16649 (N_16649,N_7815,N_11440);
and U16650 (N_16650,N_6833,N_9376);
xnor U16651 (N_16651,N_6915,N_9477);
or U16652 (N_16652,N_11820,N_11765);
nor U16653 (N_16653,N_7217,N_9505);
or U16654 (N_16654,N_10885,N_10710);
xnor U16655 (N_16655,N_8301,N_10064);
and U16656 (N_16656,N_8095,N_6583);
nor U16657 (N_16657,N_7933,N_9224);
and U16658 (N_16658,N_8907,N_8671);
or U16659 (N_16659,N_9065,N_7256);
nor U16660 (N_16660,N_6910,N_6913);
nor U16661 (N_16661,N_9081,N_7626);
or U16662 (N_16662,N_9549,N_9905);
nand U16663 (N_16663,N_6296,N_11427);
xor U16664 (N_16664,N_8219,N_10133);
or U16665 (N_16665,N_8708,N_12332);
or U16666 (N_16666,N_9137,N_6517);
nand U16667 (N_16667,N_9283,N_11616);
or U16668 (N_16668,N_10279,N_10930);
xor U16669 (N_16669,N_9956,N_7269);
nand U16670 (N_16670,N_7096,N_9583);
and U16671 (N_16671,N_6948,N_10830);
and U16672 (N_16672,N_7918,N_8398);
and U16673 (N_16673,N_11104,N_8366);
or U16674 (N_16674,N_9067,N_10389);
or U16675 (N_16675,N_9703,N_7123);
nand U16676 (N_16676,N_11796,N_9546);
nor U16677 (N_16677,N_8132,N_9092);
and U16678 (N_16678,N_8549,N_6509);
nand U16679 (N_16679,N_10986,N_11313);
and U16680 (N_16680,N_6342,N_11296);
nand U16681 (N_16681,N_9560,N_6664);
and U16682 (N_16682,N_10978,N_11648);
nand U16683 (N_16683,N_9808,N_7753);
xor U16684 (N_16684,N_7985,N_7999);
nand U16685 (N_16685,N_7826,N_8565);
xor U16686 (N_16686,N_8726,N_9149);
and U16687 (N_16687,N_10908,N_8455);
and U16688 (N_16688,N_6365,N_8451);
nor U16689 (N_16689,N_6298,N_8059);
nor U16690 (N_16690,N_11923,N_12254);
and U16691 (N_16691,N_8180,N_9391);
or U16692 (N_16692,N_7316,N_12302);
or U16693 (N_16693,N_9280,N_7872);
and U16694 (N_16694,N_10381,N_7947);
xor U16695 (N_16695,N_7662,N_8785);
and U16696 (N_16696,N_8734,N_11708);
and U16697 (N_16697,N_6554,N_9423);
nand U16698 (N_16698,N_8564,N_7134);
xor U16699 (N_16699,N_7627,N_6489);
nor U16700 (N_16700,N_6293,N_9905);
nor U16701 (N_16701,N_8205,N_6284);
nor U16702 (N_16702,N_10473,N_6817);
xor U16703 (N_16703,N_8967,N_9428);
and U16704 (N_16704,N_7892,N_11660);
or U16705 (N_16705,N_7053,N_10226);
and U16706 (N_16706,N_11139,N_9646);
and U16707 (N_16707,N_6381,N_7065);
or U16708 (N_16708,N_12416,N_10556);
nor U16709 (N_16709,N_7500,N_6444);
nand U16710 (N_16710,N_6512,N_12367);
or U16711 (N_16711,N_6624,N_10611);
nor U16712 (N_16712,N_11451,N_6649);
nand U16713 (N_16713,N_7611,N_8369);
xor U16714 (N_16714,N_9928,N_8014);
xnor U16715 (N_16715,N_11599,N_6944);
or U16716 (N_16716,N_9411,N_12111);
nor U16717 (N_16717,N_9475,N_10643);
or U16718 (N_16718,N_10838,N_10862);
and U16719 (N_16719,N_9938,N_9742);
or U16720 (N_16720,N_10367,N_9954);
nand U16721 (N_16721,N_9819,N_10488);
xor U16722 (N_16722,N_11639,N_10254);
xor U16723 (N_16723,N_9506,N_6774);
nand U16724 (N_16724,N_8520,N_7633);
or U16725 (N_16725,N_9283,N_9614);
or U16726 (N_16726,N_12327,N_12082);
nor U16727 (N_16727,N_8756,N_6833);
or U16728 (N_16728,N_10426,N_6622);
and U16729 (N_16729,N_7307,N_7542);
nand U16730 (N_16730,N_6694,N_10315);
or U16731 (N_16731,N_12210,N_7467);
and U16732 (N_16732,N_12018,N_9402);
nand U16733 (N_16733,N_12341,N_7360);
or U16734 (N_16734,N_8686,N_8219);
nor U16735 (N_16735,N_8316,N_10081);
nand U16736 (N_16736,N_10961,N_8672);
and U16737 (N_16737,N_12008,N_8881);
or U16738 (N_16738,N_6901,N_9392);
nor U16739 (N_16739,N_11599,N_6512);
nand U16740 (N_16740,N_9217,N_6994);
or U16741 (N_16741,N_10145,N_8001);
nand U16742 (N_16742,N_9001,N_12496);
nand U16743 (N_16743,N_7509,N_7470);
xnor U16744 (N_16744,N_8247,N_8170);
and U16745 (N_16745,N_10148,N_7787);
nand U16746 (N_16746,N_9415,N_8314);
nand U16747 (N_16747,N_7553,N_12292);
nand U16748 (N_16748,N_10538,N_12052);
and U16749 (N_16749,N_6929,N_12041);
or U16750 (N_16750,N_11349,N_10842);
nand U16751 (N_16751,N_9588,N_9013);
xnor U16752 (N_16752,N_8539,N_12143);
xnor U16753 (N_16753,N_11680,N_6258);
nor U16754 (N_16754,N_6859,N_10185);
nand U16755 (N_16755,N_10416,N_11941);
xor U16756 (N_16756,N_8608,N_10998);
xnor U16757 (N_16757,N_7010,N_10339);
or U16758 (N_16758,N_6254,N_10973);
and U16759 (N_16759,N_11523,N_11395);
nand U16760 (N_16760,N_12065,N_8465);
nor U16761 (N_16761,N_12118,N_11710);
or U16762 (N_16762,N_12151,N_10243);
and U16763 (N_16763,N_11504,N_12267);
xnor U16764 (N_16764,N_10789,N_9502);
and U16765 (N_16765,N_6834,N_10869);
nand U16766 (N_16766,N_7821,N_8449);
nand U16767 (N_16767,N_7543,N_7230);
xor U16768 (N_16768,N_8585,N_9082);
xnor U16769 (N_16769,N_7210,N_11325);
xor U16770 (N_16770,N_7262,N_8054);
nand U16771 (N_16771,N_7330,N_10484);
xnor U16772 (N_16772,N_7520,N_6927);
or U16773 (N_16773,N_10539,N_6966);
nand U16774 (N_16774,N_12488,N_8778);
nand U16775 (N_16775,N_8925,N_11926);
and U16776 (N_16776,N_11277,N_7947);
and U16777 (N_16777,N_8370,N_10787);
xnor U16778 (N_16778,N_6715,N_6975);
nand U16779 (N_16779,N_11274,N_11286);
nand U16780 (N_16780,N_6268,N_10212);
nor U16781 (N_16781,N_10821,N_7262);
xor U16782 (N_16782,N_6719,N_11688);
nand U16783 (N_16783,N_10902,N_7457);
nor U16784 (N_16784,N_11694,N_10589);
or U16785 (N_16785,N_8833,N_6939);
nor U16786 (N_16786,N_6698,N_6343);
nand U16787 (N_16787,N_11995,N_11017);
nor U16788 (N_16788,N_8910,N_9744);
and U16789 (N_16789,N_10350,N_11709);
and U16790 (N_16790,N_9833,N_9368);
nand U16791 (N_16791,N_8194,N_9144);
and U16792 (N_16792,N_7098,N_9583);
nand U16793 (N_16793,N_11257,N_10840);
nand U16794 (N_16794,N_8289,N_11571);
nand U16795 (N_16795,N_7435,N_12430);
nand U16796 (N_16796,N_10184,N_6547);
xor U16797 (N_16797,N_8197,N_8784);
or U16798 (N_16798,N_6805,N_6365);
nand U16799 (N_16799,N_10181,N_6480);
nor U16800 (N_16800,N_8694,N_8389);
xor U16801 (N_16801,N_11431,N_11783);
nor U16802 (N_16802,N_10675,N_7642);
and U16803 (N_16803,N_11369,N_12204);
nand U16804 (N_16804,N_9131,N_9839);
nor U16805 (N_16805,N_9396,N_7894);
nand U16806 (N_16806,N_12458,N_10858);
and U16807 (N_16807,N_8956,N_8568);
xnor U16808 (N_16808,N_11907,N_6857);
xnor U16809 (N_16809,N_7409,N_7220);
xnor U16810 (N_16810,N_10888,N_8900);
nor U16811 (N_16811,N_9615,N_12341);
xor U16812 (N_16812,N_9225,N_7308);
nand U16813 (N_16813,N_9630,N_10725);
nand U16814 (N_16814,N_8431,N_10985);
xor U16815 (N_16815,N_7019,N_10977);
or U16816 (N_16816,N_11550,N_9613);
nor U16817 (N_16817,N_9726,N_9561);
xor U16818 (N_16818,N_12217,N_9171);
nand U16819 (N_16819,N_7976,N_8770);
nor U16820 (N_16820,N_8560,N_11507);
nor U16821 (N_16821,N_11043,N_8168);
and U16822 (N_16822,N_8104,N_6308);
nand U16823 (N_16823,N_10957,N_11148);
xor U16824 (N_16824,N_8595,N_11849);
and U16825 (N_16825,N_7790,N_8376);
or U16826 (N_16826,N_7776,N_9649);
nand U16827 (N_16827,N_6726,N_11695);
or U16828 (N_16828,N_7030,N_10312);
nor U16829 (N_16829,N_11378,N_6571);
or U16830 (N_16830,N_10930,N_9818);
nor U16831 (N_16831,N_7867,N_6399);
xor U16832 (N_16832,N_6543,N_12450);
and U16833 (N_16833,N_6261,N_9293);
xor U16834 (N_16834,N_9727,N_11241);
xnor U16835 (N_16835,N_12347,N_11288);
nand U16836 (N_16836,N_7503,N_8149);
xor U16837 (N_16837,N_7795,N_8543);
nor U16838 (N_16838,N_9398,N_7091);
nor U16839 (N_16839,N_12302,N_12163);
and U16840 (N_16840,N_10308,N_11224);
nor U16841 (N_16841,N_9719,N_10792);
xor U16842 (N_16842,N_6319,N_9626);
nand U16843 (N_16843,N_8879,N_9981);
nor U16844 (N_16844,N_12025,N_8963);
and U16845 (N_16845,N_11361,N_6833);
xnor U16846 (N_16846,N_7530,N_8966);
xnor U16847 (N_16847,N_7456,N_6554);
or U16848 (N_16848,N_7609,N_10982);
nor U16849 (N_16849,N_11742,N_6987);
and U16850 (N_16850,N_11225,N_6324);
or U16851 (N_16851,N_11712,N_7183);
and U16852 (N_16852,N_8270,N_11594);
xor U16853 (N_16853,N_10066,N_7922);
and U16854 (N_16854,N_7435,N_8542);
nand U16855 (N_16855,N_9692,N_9840);
nor U16856 (N_16856,N_9029,N_9582);
nand U16857 (N_16857,N_12181,N_7182);
nor U16858 (N_16858,N_10714,N_12185);
nor U16859 (N_16859,N_6842,N_8432);
or U16860 (N_16860,N_7115,N_8031);
xor U16861 (N_16861,N_7408,N_7171);
and U16862 (N_16862,N_10202,N_8998);
xnor U16863 (N_16863,N_9987,N_10964);
nor U16864 (N_16864,N_7753,N_9919);
xnor U16865 (N_16865,N_8746,N_8294);
xnor U16866 (N_16866,N_6341,N_6380);
nand U16867 (N_16867,N_9300,N_12350);
nand U16868 (N_16868,N_7785,N_12274);
xor U16869 (N_16869,N_7787,N_9310);
nand U16870 (N_16870,N_10041,N_10060);
or U16871 (N_16871,N_11352,N_10743);
or U16872 (N_16872,N_11700,N_11173);
or U16873 (N_16873,N_8532,N_7271);
xor U16874 (N_16874,N_10687,N_9845);
nor U16875 (N_16875,N_11233,N_10672);
xor U16876 (N_16876,N_12152,N_10730);
nor U16877 (N_16877,N_10738,N_12318);
nor U16878 (N_16878,N_7586,N_6787);
xnor U16879 (N_16879,N_12071,N_6433);
nor U16880 (N_16880,N_10051,N_8669);
and U16881 (N_16881,N_10933,N_10598);
or U16882 (N_16882,N_10212,N_9167);
nand U16883 (N_16883,N_9872,N_9553);
and U16884 (N_16884,N_7296,N_6632);
or U16885 (N_16885,N_7027,N_11357);
xnor U16886 (N_16886,N_11016,N_11253);
and U16887 (N_16887,N_9167,N_6298);
nor U16888 (N_16888,N_12189,N_6527);
nor U16889 (N_16889,N_11395,N_6358);
nor U16890 (N_16890,N_6458,N_12140);
or U16891 (N_16891,N_6967,N_7255);
or U16892 (N_16892,N_9298,N_7624);
nand U16893 (N_16893,N_9174,N_9788);
nor U16894 (N_16894,N_8195,N_7809);
or U16895 (N_16895,N_8892,N_6940);
nand U16896 (N_16896,N_11871,N_7338);
nand U16897 (N_16897,N_10178,N_7388);
xnor U16898 (N_16898,N_9417,N_8388);
or U16899 (N_16899,N_8408,N_8477);
and U16900 (N_16900,N_9960,N_8387);
or U16901 (N_16901,N_11010,N_8145);
nor U16902 (N_16902,N_6700,N_12238);
and U16903 (N_16903,N_11458,N_11590);
nor U16904 (N_16904,N_12316,N_8960);
or U16905 (N_16905,N_8798,N_6442);
and U16906 (N_16906,N_9518,N_10873);
nand U16907 (N_16907,N_10546,N_7454);
nor U16908 (N_16908,N_11175,N_8450);
and U16909 (N_16909,N_6591,N_9750);
and U16910 (N_16910,N_7122,N_8710);
xnor U16911 (N_16911,N_6319,N_8296);
nor U16912 (N_16912,N_9072,N_12117);
and U16913 (N_16913,N_10488,N_9463);
or U16914 (N_16914,N_12381,N_6511);
or U16915 (N_16915,N_10817,N_11253);
nand U16916 (N_16916,N_11022,N_8072);
xnor U16917 (N_16917,N_9724,N_10314);
and U16918 (N_16918,N_6957,N_11851);
nor U16919 (N_16919,N_11549,N_10187);
xnor U16920 (N_16920,N_8948,N_11504);
nor U16921 (N_16921,N_10574,N_6432);
nor U16922 (N_16922,N_10091,N_9275);
xnor U16923 (N_16923,N_11435,N_7453);
xor U16924 (N_16924,N_8326,N_8858);
and U16925 (N_16925,N_8773,N_12256);
and U16926 (N_16926,N_11246,N_11936);
nor U16927 (N_16927,N_9579,N_6899);
nor U16928 (N_16928,N_9855,N_7590);
nor U16929 (N_16929,N_9458,N_10312);
nand U16930 (N_16930,N_8304,N_6409);
or U16931 (N_16931,N_6623,N_6970);
nor U16932 (N_16932,N_7831,N_7707);
and U16933 (N_16933,N_9094,N_7177);
nand U16934 (N_16934,N_9868,N_10852);
or U16935 (N_16935,N_7017,N_11749);
nand U16936 (N_16936,N_8461,N_10233);
nor U16937 (N_16937,N_9607,N_7881);
nand U16938 (N_16938,N_9429,N_6574);
nor U16939 (N_16939,N_9540,N_10309);
and U16940 (N_16940,N_8362,N_10774);
nand U16941 (N_16941,N_6561,N_11017);
or U16942 (N_16942,N_10064,N_7098);
and U16943 (N_16943,N_7269,N_8848);
nand U16944 (N_16944,N_11315,N_7580);
or U16945 (N_16945,N_6748,N_6855);
nand U16946 (N_16946,N_6354,N_7466);
or U16947 (N_16947,N_8864,N_7147);
xnor U16948 (N_16948,N_10346,N_10237);
xor U16949 (N_16949,N_10237,N_8736);
xnor U16950 (N_16950,N_6455,N_7858);
xor U16951 (N_16951,N_9931,N_6988);
xor U16952 (N_16952,N_8156,N_12401);
and U16953 (N_16953,N_9701,N_10473);
nor U16954 (N_16954,N_11489,N_7853);
xnor U16955 (N_16955,N_7955,N_7190);
or U16956 (N_16956,N_10311,N_6601);
or U16957 (N_16957,N_8129,N_8600);
nand U16958 (N_16958,N_9375,N_8485);
nor U16959 (N_16959,N_10519,N_9350);
and U16960 (N_16960,N_7376,N_6323);
or U16961 (N_16961,N_12219,N_9895);
or U16962 (N_16962,N_10403,N_8999);
nor U16963 (N_16963,N_6712,N_10895);
or U16964 (N_16964,N_10997,N_12186);
xor U16965 (N_16965,N_6767,N_6326);
xor U16966 (N_16966,N_10600,N_7055);
nand U16967 (N_16967,N_7309,N_10525);
xor U16968 (N_16968,N_7712,N_6755);
nor U16969 (N_16969,N_11957,N_12081);
xor U16970 (N_16970,N_7182,N_7375);
nor U16971 (N_16971,N_9089,N_8167);
or U16972 (N_16972,N_11707,N_10676);
nand U16973 (N_16973,N_8677,N_6540);
and U16974 (N_16974,N_11666,N_6455);
nand U16975 (N_16975,N_10928,N_8738);
or U16976 (N_16976,N_10296,N_9210);
nand U16977 (N_16977,N_6859,N_8969);
xor U16978 (N_16978,N_12329,N_10911);
nor U16979 (N_16979,N_11607,N_10069);
and U16980 (N_16980,N_7428,N_11718);
and U16981 (N_16981,N_12009,N_6440);
xor U16982 (N_16982,N_11636,N_7471);
xor U16983 (N_16983,N_8527,N_11316);
nand U16984 (N_16984,N_7832,N_8927);
nand U16985 (N_16985,N_11234,N_7094);
and U16986 (N_16986,N_8083,N_6854);
or U16987 (N_16987,N_8318,N_6846);
nor U16988 (N_16988,N_7246,N_7053);
nor U16989 (N_16989,N_7042,N_11829);
nor U16990 (N_16990,N_9796,N_6359);
xor U16991 (N_16991,N_9270,N_10877);
or U16992 (N_16992,N_9116,N_9212);
xnor U16993 (N_16993,N_8479,N_8428);
xnor U16994 (N_16994,N_9208,N_6305);
or U16995 (N_16995,N_10359,N_8559);
or U16996 (N_16996,N_11263,N_7981);
or U16997 (N_16997,N_7849,N_8286);
nor U16998 (N_16998,N_9701,N_9625);
xnor U16999 (N_16999,N_9529,N_12066);
and U17000 (N_17000,N_11138,N_6722);
and U17001 (N_17001,N_10902,N_10295);
and U17002 (N_17002,N_10274,N_6803);
xnor U17003 (N_17003,N_10567,N_8701);
nor U17004 (N_17004,N_11529,N_12137);
nand U17005 (N_17005,N_11210,N_11285);
or U17006 (N_17006,N_9741,N_6392);
xor U17007 (N_17007,N_6411,N_8977);
or U17008 (N_17008,N_8643,N_8266);
and U17009 (N_17009,N_6645,N_10574);
xnor U17010 (N_17010,N_11117,N_11506);
and U17011 (N_17011,N_9611,N_8407);
nor U17012 (N_17012,N_7216,N_6501);
and U17013 (N_17013,N_9882,N_7813);
nand U17014 (N_17014,N_9110,N_12343);
nand U17015 (N_17015,N_8358,N_8681);
and U17016 (N_17016,N_9562,N_8627);
or U17017 (N_17017,N_7105,N_8831);
nor U17018 (N_17018,N_9638,N_11651);
xor U17019 (N_17019,N_10351,N_11059);
nor U17020 (N_17020,N_7203,N_9172);
and U17021 (N_17021,N_7261,N_10949);
and U17022 (N_17022,N_10100,N_10369);
nand U17023 (N_17023,N_12227,N_7702);
xor U17024 (N_17024,N_10763,N_7008);
or U17025 (N_17025,N_9708,N_8742);
or U17026 (N_17026,N_8118,N_8129);
xnor U17027 (N_17027,N_8223,N_6777);
and U17028 (N_17028,N_9973,N_11569);
or U17029 (N_17029,N_10540,N_8219);
nor U17030 (N_17030,N_7615,N_10581);
and U17031 (N_17031,N_7125,N_9358);
xor U17032 (N_17032,N_7833,N_9087);
or U17033 (N_17033,N_10302,N_7441);
or U17034 (N_17034,N_8344,N_10826);
or U17035 (N_17035,N_11533,N_12380);
and U17036 (N_17036,N_8869,N_9136);
or U17037 (N_17037,N_10054,N_7435);
xnor U17038 (N_17038,N_10828,N_9985);
nor U17039 (N_17039,N_10122,N_10917);
and U17040 (N_17040,N_9595,N_7664);
nor U17041 (N_17041,N_8257,N_9319);
and U17042 (N_17042,N_7451,N_10407);
nand U17043 (N_17043,N_9622,N_12003);
or U17044 (N_17044,N_9639,N_12198);
or U17045 (N_17045,N_10308,N_9695);
nand U17046 (N_17046,N_7046,N_9057);
and U17047 (N_17047,N_7483,N_10789);
and U17048 (N_17048,N_9497,N_7250);
or U17049 (N_17049,N_9847,N_11682);
and U17050 (N_17050,N_7496,N_7010);
or U17051 (N_17051,N_10867,N_6796);
nor U17052 (N_17052,N_8127,N_6830);
and U17053 (N_17053,N_7864,N_11157);
or U17054 (N_17054,N_9423,N_12153);
nor U17055 (N_17055,N_7079,N_9055);
nor U17056 (N_17056,N_6470,N_10031);
and U17057 (N_17057,N_10867,N_7868);
nor U17058 (N_17058,N_10735,N_9825);
xor U17059 (N_17059,N_9993,N_9175);
and U17060 (N_17060,N_11719,N_10399);
nor U17061 (N_17061,N_8335,N_12062);
and U17062 (N_17062,N_9700,N_7958);
and U17063 (N_17063,N_11123,N_7460);
nand U17064 (N_17064,N_12221,N_7934);
and U17065 (N_17065,N_7725,N_9700);
and U17066 (N_17066,N_10301,N_10240);
and U17067 (N_17067,N_6660,N_10633);
nor U17068 (N_17068,N_7689,N_11951);
and U17069 (N_17069,N_9299,N_9872);
xor U17070 (N_17070,N_7266,N_7921);
nor U17071 (N_17071,N_6672,N_6482);
xor U17072 (N_17072,N_9560,N_7423);
xor U17073 (N_17073,N_6451,N_11694);
or U17074 (N_17074,N_7836,N_10971);
and U17075 (N_17075,N_12334,N_7221);
or U17076 (N_17076,N_6629,N_8688);
or U17077 (N_17077,N_11905,N_12320);
xnor U17078 (N_17078,N_7117,N_11232);
nand U17079 (N_17079,N_7688,N_9370);
xnor U17080 (N_17080,N_8578,N_7916);
or U17081 (N_17081,N_6693,N_7040);
nor U17082 (N_17082,N_10992,N_12452);
xor U17083 (N_17083,N_10179,N_12025);
or U17084 (N_17084,N_11368,N_10571);
xor U17085 (N_17085,N_7949,N_7449);
nand U17086 (N_17086,N_12356,N_9148);
nand U17087 (N_17087,N_8141,N_10929);
and U17088 (N_17088,N_9272,N_9680);
and U17089 (N_17089,N_8834,N_9269);
and U17090 (N_17090,N_8817,N_8183);
nor U17091 (N_17091,N_8733,N_11510);
xor U17092 (N_17092,N_10352,N_12215);
and U17093 (N_17093,N_11736,N_6880);
xor U17094 (N_17094,N_9039,N_7480);
nand U17095 (N_17095,N_11037,N_10657);
and U17096 (N_17096,N_11524,N_6772);
and U17097 (N_17097,N_7994,N_11727);
and U17098 (N_17098,N_11692,N_6902);
xor U17099 (N_17099,N_9560,N_9180);
xnor U17100 (N_17100,N_11058,N_11192);
nor U17101 (N_17101,N_8966,N_9799);
nor U17102 (N_17102,N_12094,N_6359);
and U17103 (N_17103,N_9219,N_10191);
and U17104 (N_17104,N_11837,N_6926);
nand U17105 (N_17105,N_10980,N_7053);
nand U17106 (N_17106,N_11359,N_7887);
xnor U17107 (N_17107,N_8267,N_11175);
xor U17108 (N_17108,N_8827,N_6797);
and U17109 (N_17109,N_6506,N_10747);
xor U17110 (N_17110,N_8839,N_10874);
xor U17111 (N_17111,N_9242,N_10979);
or U17112 (N_17112,N_12369,N_7709);
nor U17113 (N_17113,N_11152,N_11351);
nor U17114 (N_17114,N_9328,N_8739);
nor U17115 (N_17115,N_9724,N_7526);
nor U17116 (N_17116,N_12090,N_7645);
or U17117 (N_17117,N_6784,N_7819);
nand U17118 (N_17118,N_9640,N_10305);
or U17119 (N_17119,N_7973,N_8010);
or U17120 (N_17120,N_10243,N_11647);
and U17121 (N_17121,N_11176,N_10564);
nand U17122 (N_17122,N_8834,N_12277);
and U17123 (N_17123,N_7355,N_10716);
and U17124 (N_17124,N_10771,N_8373);
xor U17125 (N_17125,N_8729,N_8111);
or U17126 (N_17126,N_10905,N_10429);
xnor U17127 (N_17127,N_12205,N_9104);
and U17128 (N_17128,N_9310,N_11859);
or U17129 (N_17129,N_10144,N_8128);
or U17130 (N_17130,N_9683,N_9900);
xor U17131 (N_17131,N_10392,N_11939);
nor U17132 (N_17132,N_6579,N_8748);
or U17133 (N_17133,N_8200,N_10718);
or U17134 (N_17134,N_6746,N_7235);
nor U17135 (N_17135,N_9631,N_11883);
and U17136 (N_17136,N_12378,N_7104);
nand U17137 (N_17137,N_12061,N_6350);
nor U17138 (N_17138,N_9946,N_12357);
and U17139 (N_17139,N_7568,N_7697);
nand U17140 (N_17140,N_9220,N_9883);
nand U17141 (N_17141,N_7890,N_12202);
nand U17142 (N_17142,N_8598,N_9873);
xnor U17143 (N_17143,N_11017,N_11764);
or U17144 (N_17144,N_10772,N_12086);
xor U17145 (N_17145,N_8319,N_9335);
or U17146 (N_17146,N_9985,N_11370);
or U17147 (N_17147,N_8760,N_11155);
nand U17148 (N_17148,N_7092,N_11356);
nand U17149 (N_17149,N_10878,N_6431);
nand U17150 (N_17150,N_11347,N_8518);
or U17151 (N_17151,N_9873,N_7127);
and U17152 (N_17152,N_7060,N_11614);
xnor U17153 (N_17153,N_9915,N_6497);
nor U17154 (N_17154,N_7441,N_10653);
nand U17155 (N_17155,N_9107,N_9427);
nor U17156 (N_17156,N_9086,N_8333);
nor U17157 (N_17157,N_8466,N_8918);
nand U17158 (N_17158,N_10586,N_6504);
xor U17159 (N_17159,N_8105,N_9880);
or U17160 (N_17160,N_10257,N_11292);
xnor U17161 (N_17161,N_11603,N_12365);
nand U17162 (N_17162,N_7819,N_10016);
and U17163 (N_17163,N_6679,N_9599);
and U17164 (N_17164,N_6814,N_10129);
nand U17165 (N_17165,N_10057,N_8215);
nand U17166 (N_17166,N_7783,N_8089);
xnor U17167 (N_17167,N_6989,N_6299);
and U17168 (N_17168,N_11399,N_8416);
xor U17169 (N_17169,N_10363,N_8455);
nand U17170 (N_17170,N_6357,N_6537);
xnor U17171 (N_17171,N_11063,N_11590);
nor U17172 (N_17172,N_6730,N_10409);
xor U17173 (N_17173,N_7365,N_10914);
xor U17174 (N_17174,N_6494,N_9778);
and U17175 (N_17175,N_9500,N_7653);
and U17176 (N_17176,N_12400,N_6485);
or U17177 (N_17177,N_7507,N_6976);
or U17178 (N_17178,N_11481,N_12144);
and U17179 (N_17179,N_10004,N_11335);
xor U17180 (N_17180,N_6735,N_7876);
nor U17181 (N_17181,N_6265,N_12389);
nand U17182 (N_17182,N_7019,N_7826);
or U17183 (N_17183,N_8293,N_11259);
xnor U17184 (N_17184,N_8212,N_7710);
nand U17185 (N_17185,N_6590,N_12373);
nand U17186 (N_17186,N_10303,N_7037);
and U17187 (N_17187,N_11146,N_12029);
or U17188 (N_17188,N_11817,N_10688);
or U17189 (N_17189,N_7140,N_9451);
or U17190 (N_17190,N_8189,N_9360);
and U17191 (N_17191,N_11176,N_9627);
nor U17192 (N_17192,N_8285,N_7776);
nand U17193 (N_17193,N_10483,N_7242);
and U17194 (N_17194,N_6528,N_10990);
nand U17195 (N_17195,N_6611,N_6866);
nand U17196 (N_17196,N_9415,N_9338);
and U17197 (N_17197,N_6394,N_11862);
nand U17198 (N_17198,N_7795,N_10765);
or U17199 (N_17199,N_12353,N_9959);
or U17200 (N_17200,N_11093,N_7717);
nand U17201 (N_17201,N_6893,N_9751);
and U17202 (N_17202,N_7816,N_10341);
nand U17203 (N_17203,N_6768,N_10290);
xnor U17204 (N_17204,N_11688,N_6956);
nand U17205 (N_17205,N_10871,N_9010);
nor U17206 (N_17206,N_12496,N_6517);
nand U17207 (N_17207,N_12081,N_7630);
xor U17208 (N_17208,N_7005,N_10787);
nor U17209 (N_17209,N_10332,N_9380);
nand U17210 (N_17210,N_8547,N_11969);
or U17211 (N_17211,N_9038,N_8475);
xnor U17212 (N_17212,N_12472,N_10656);
nand U17213 (N_17213,N_8911,N_8942);
nor U17214 (N_17214,N_6973,N_11185);
or U17215 (N_17215,N_6274,N_8940);
or U17216 (N_17216,N_11030,N_10199);
and U17217 (N_17217,N_9093,N_12497);
nor U17218 (N_17218,N_7976,N_11651);
nand U17219 (N_17219,N_11030,N_8071);
and U17220 (N_17220,N_8999,N_9757);
nor U17221 (N_17221,N_7440,N_8887);
and U17222 (N_17222,N_12240,N_8604);
and U17223 (N_17223,N_6969,N_6270);
or U17224 (N_17224,N_10990,N_7243);
xor U17225 (N_17225,N_9511,N_7178);
or U17226 (N_17226,N_9825,N_8367);
nand U17227 (N_17227,N_7939,N_11069);
and U17228 (N_17228,N_8269,N_11407);
nor U17229 (N_17229,N_6801,N_11180);
and U17230 (N_17230,N_10257,N_7532);
and U17231 (N_17231,N_8509,N_7351);
xor U17232 (N_17232,N_12005,N_11248);
nor U17233 (N_17233,N_12401,N_10945);
and U17234 (N_17234,N_7499,N_8601);
nand U17235 (N_17235,N_8013,N_8562);
and U17236 (N_17236,N_6406,N_8755);
nor U17237 (N_17237,N_10828,N_6874);
or U17238 (N_17238,N_10750,N_7136);
nor U17239 (N_17239,N_11105,N_7000);
nand U17240 (N_17240,N_8169,N_8622);
xnor U17241 (N_17241,N_9889,N_6388);
nand U17242 (N_17242,N_11393,N_10044);
nor U17243 (N_17243,N_9689,N_10816);
nand U17244 (N_17244,N_11627,N_10556);
or U17245 (N_17245,N_7968,N_9114);
and U17246 (N_17246,N_12041,N_11458);
and U17247 (N_17247,N_12243,N_9001);
xor U17248 (N_17248,N_6609,N_7451);
or U17249 (N_17249,N_6652,N_6584);
xnor U17250 (N_17250,N_6708,N_11752);
or U17251 (N_17251,N_11677,N_12109);
or U17252 (N_17252,N_9993,N_8939);
nor U17253 (N_17253,N_9517,N_9856);
nor U17254 (N_17254,N_7637,N_9367);
nand U17255 (N_17255,N_6537,N_11723);
xor U17256 (N_17256,N_10201,N_10473);
and U17257 (N_17257,N_9337,N_10412);
xnor U17258 (N_17258,N_10815,N_8469);
xnor U17259 (N_17259,N_8193,N_12047);
or U17260 (N_17260,N_6482,N_11638);
nand U17261 (N_17261,N_11908,N_8113);
and U17262 (N_17262,N_9688,N_8058);
xnor U17263 (N_17263,N_6757,N_6489);
nand U17264 (N_17264,N_6627,N_12062);
or U17265 (N_17265,N_7125,N_9504);
and U17266 (N_17266,N_8779,N_8417);
or U17267 (N_17267,N_7603,N_11646);
xnor U17268 (N_17268,N_6431,N_12379);
or U17269 (N_17269,N_7881,N_6969);
nand U17270 (N_17270,N_8117,N_10716);
xor U17271 (N_17271,N_7203,N_10587);
xnor U17272 (N_17272,N_11955,N_6290);
xor U17273 (N_17273,N_10338,N_8990);
or U17274 (N_17274,N_6759,N_9573);
and U17275 (N_17275,N_7752,N_10772);
and U17276 (N_17276,N_11241,N_8290);
nor U17277 (N_17277,N_12296,N_6517);
nor U17278 (N_17278,N_7695,N_11219);
xor U17279 (N_17279,N_7158,N_7491);
and U17280 (N_17280,N_7986,N_11371);
nor U17281 (N_17281,N_9620,N_12172);
nand U17282 (N_17282,N_9329,N_11598);
nand U17283 (N_17283,N_7995,N_9528);
nand U17284 (N_17284,N_11884,N_7616);
nand U17285 (N_17285,N_10149,N_9695);
xor U17286 (N_17286,N_7292,N_7413);
nand U17287 (N_17287,N_11720,N_7811);
nor U17288 (N_17288,N_9380,N_6333);
and U17289 (N_17289,N_11562,N_10411);
xor U17290 (N_17290,N_11731,N_11972);
nor U17291 (N_17291,N_7540,N_9788);
and U17292 (N_17292,N_10080,N_7221);
xnor U17293 (N_17293,N_6433,N_6324);
xor U17294 (N_17294,N_7651,N_10555);
xnor U17295 (N_17295,N_11553,N_10779);
nor U17296 (N_17296,N_12422,N_9207);
nor U17297 (N_17297,N_7193,N_6380);
and U17298 (N_17298,N_9231,N_10227);
xor U17299 (N_17299,N_8741,N_7727);
xnor U17300 (N_17300,N_11313,N_6418);
or U17301 (N_17301,N_8766,N_7266);
xor U17302 (N_17302,N_6623,N_9312);
and U17303 (N_17303,N_6879,N_10264);
nand U17304 (N_17304,N_10075,N_6526);
or U17305 (N_17305,N_10781,N_8126);
xnor U17306 (N_17306,N_7146,N_7931);
and U17307 (N_17307,N_10120,N_7490);
nand U17308 (N_17308,N_7385,N_10378);
nand U17309 (N_17309,N_10965,N_8089);
nor U17310 (N_17310,N_7948,N_10378);
xnor U17311 (N_17311,N_7009,N_12104);
or U17312 (N_17312,N_8089,N_8742);
xor U17313 (N_17313,N_12191,N_11417);
nor U17314 (N_17314,N_6409,N_7415);
xnor U17315 (N_17315,N_11094,N_9153);
xnor U17316 (N_17316,N_10875,N_10381);
nor U17317 (N_17317,N_7913,N_8451);
and U17318 (N_17318,N_6736,N_7966);
nand U17319 (N_17319,N_8984,N_12335);
or U17320 (N_17320,N_6929,N_8431);
nor U17321 (N_17321,N_7689,N_6857);
xor U17322 (N_17322,N_11269,N_9139);
xnor U17323 (N_17323,N_8360,N_10490);
or U17324 (N_17324,N_11370,N_10142);
xnor U17325 (N_17325,N_12000,N_10216);
nor U17326 (N_17326,N_8983,N_8721);
and U17327 (N_17327,N_8430,N_12073);
or U17328 (N_17328,N_6431,N_9693);
and U17329 (N_17329,N_9283,N_6824);
and U17330 (N_17330,N_7920,N_9267);
and U17331 (N_17331,N_11888,N_11839);
nand U17332 (N_17332,N_10008,N_8372);
or U17333 (N_17333,N_11105,N_8209);
and U17334 (N_17334,N_8674,N_9484);
and U17335 (N_17335,N_6696,N_7523);
or U17336 (N_17336,N_6312,N_9909);
nand U17337 (N_17337,N_10875,N_9667);
and U17338 (N_17338,N_12294,N_7875);
nor U17339 (N_17339,N_7707,N_8570);
or U17340 (N_17340,N_9789,N_9079);
xor U17341 (N_17341,N_12152,N_6843);
and U17342 (N_17342,N_12172,N_9988);
xnor U17343 (N_17343,N_6384,N_11675);
or U17344 (N_17344,N_11747,N_12093);
or U17345 (N_17345,N_10828,N_11042);
nand U17346 (N_17346,N_10749,N_9294);
nand U17347 (N_17347,N_9361,N_8653);
nor U17348 (N_17348,N_10079,N_10136);
nand U17349 (N_17349,N_8241,N_9026);
xor U17350 (N_17350,N_9116,N_8884);
nor U17351 (N_17351,N_8905,N_7747);
nor U17352 (N_17352,N_8300,N_12400);
xor U17353 (N_17353,N_10009,N_6797);
and U17354 (N_17354,N_8796,N_8781);
and U17355 (N_17355,N_10594,N_7088);
nand U17356 (N_17356,N_6923,N_10639);
and U17357 (N_17357,N_9729,N_10405);
xor U17358 (N_17358,N_10313,N_9960);
xor U17359 (N_17359,N_11238,N_7371);
or U17360 (N_17360,N_9906,N_10865);
or U17361 (N_17361,N_10658,N_10670);
xnor U17362 (N_17362,N_9791,N_11874);
nand U17363 (N_17363,N_8589,N_8477);
xor U17364 (N_17364,N_9573,N_12474);
nand U17365 (N_17365,N_10560,N_9373);
xor U17366 (N_17366,N_12490,N_7907);
xnor U17367 (N_17367,N_9476,N_9912);
xor U17368 (N_17368,N_11023,N_10654);
and U17369 (N_17369,N_11790,N_10657);
nand U17370 (N_17370,N_9045,N_9185);
or U17371 (N_17371,N_11775,N_10597);
xor U17372 (N_17372,N_10148,N_8390);
xnor U17373 (N_17373,N_7039,N_7131);
nor U17374 (N_17374,N_9128,N_7006);
nor U17375 (N_17375,N_8801,N_11164);
xnor U17376 (N_17376,N_10220,N_8115);
or U17377 (N_17377,N_9288,N_6679);
xor U17378 (N_17378,N_6349,N_11713);
nor U17379 (N_17379,N_7031,N_12421);
or U17380 (N_17380,N_8609,N_9994);
xnor U17381 (N_17381,N_6750,N_11915);
nor U17382 (N_17382,N_11626,N_11096);
nand U17383 (N_17383,N_12202,N_8463);
nor U17384 (N_17384,N_9763,N_11271);
and U17385 (N_17385,N_11887,N_12238);
or U17386 (N_17386,N_10921,N_8815);
and U17387 (N_17387,N_9498,N_11625);
xnor U17388 (N_17388,N_7058,N_8359);
nand U17389 (N_17389,N_10785,N_8770);
xnor U17390 (N_17390,N_11131,N_12018);
nand U17391 (N_17391,N_7515,N_9442);
nand U17392 (N_17392,N_10689,N_11249);
or U17393 (N_17393,N_8538,N_10012);
nor U17394 (N_17394,N_12458,N_9958);
and U17395 (N_17395,N_7803,N_9454);
nand U17396 (N_17396,N_10821,N_9537);
xnor U17397 (N_17397,N_10182,N_8742);
and U17398 (N_17398,N_11309,N_8183);
nand U17399 (N_17399,N_8446,N_8590);
nor U17400 (N_17400,N_8038,N_6783);
or U17401 (N_17401,N_7721,N_8492);
xnor U17402 (N_17402,N_9137,N_11539);
and U17403 (N_17403,N_6447,N_10335);
or U17404 (N_17404,N_10190,N_7971);
nor U17405 (N_17405,N_9392,N_8762);
or U17406 (N_17406,N_6449,N_11015);
or U17407 (N_17407,N_11268,N_10368);
nand U17408 (N_17408,N_7736,N_9694);
xnor U17409 (N_17409,N_7819,N_11478);
nand U17410 (N_17410,N_11933,N_7514);
and U17411 (N_17411,N_9412,N_6326);
xnor U17412 (N_17412,N_9200,N_10710);
xor U17413 (N_17413,N_7847,N_10884);
xor U17414 (N_17414,N_8362,N_8830);
xnor U17415 (N_17415,N_10606,N_7206);
or U17416 (N_17416,N_9958,N_11440);
xor U17417 (N_17417,N_11099,N_7387);
or U17418 (N_17418,N_8813,N_8501);
or U17419 (N_17419,N_9161,N_7625);
or U17420 (N_17420,N_7030,N_12176);
and U17421 (N_17421,N_7138,N_11996);
or U17422 (N_17422,N_10000,N_7814);
xnor U17423 (N_17423,N_9070,N_11709);
or U17424 (N_17424,N_10942,N_6962);
nand U17425 (N_17425,N_8466,N_7952);
or U17426 (N_17426,N_10284,N_6476);
xnor U17427 (N_17427,N_6485,N_7579);
nor U17428 (N_17428,N_11290,N_11044);
and U17429 (N_17429,N_8756,N_7099);
or U17430 (N_17430,N_12264,N_7420);
nor U17431 (N_17431,N_10161,N_10477);
or U17432 (N_17432,N_9446,N_9306);
and U17433 (N_17433,N_12310,N_10147);
nand U17434 (N_17434,N_12298,N_8902);
or U17435 (N_17435,N_6696,N_8192);
nand U17436 (N_17436,N_10165,N_7892);
and U17437 (N_17437,N_12406,N_9606);
and U17438 (N_17438,N_8923,N_6364);
and U17439 (N_17439,N_10484,N_9859);
and U17440 (N_17440,N_9846,N_7326);
or U17441 (N_17441,N_9164,N_9612);
xnor U17442 (N_17442,N_12049,N_8371);
and U17443 (N_17443,N_7272,N_10212);
nand U17444 (N_17444,N_10238,N_11319);
nor U17445 (N_17445,N_9295,N_11018);
nor U17446 (N_17446,N_8604,N_7310);
nor U17447 (N_17447,N_6311,N_11158);
or U17448 (N_17448,N_9648,N_8998);
nor U17449 (N_17449,N_12401,N_11679);
xnor U17450 (N_17450,N_11818,N_11113);
nand U17451 (N_17451,N_7261,N_8380);
nor U17452 (N_17452,N_7994,N_9098);
or U17453 (N_17453,N_10581,N_9436);
and U17454 (N_17454,N_9015,N_8862);
xor U17455 (N_17455,N_10465,N_6856);
nor U17456 (N_17456,N_6413,N_12364);
or U17457 (N_17457,N_7325,N_8381);
and U17458 (N_17458,N_7701,N_7092);
or U17459 (N_17459,N_9789,N_8804);
xnor U17460 (N_17460,N_10725,N_6747);
and U17461 (N_17461,N_9910,N_6796);
nor U17462 (N_17462,N_8783,N_6359);
nand U17463 (N_17463,N_11426,N_6335);
and U17464 (N_17464,N_8758,N_12243);
or U17465 (N_17465,N_11138,N_10505);
or U17466 (N_17466,N_11508,N_12176);
xnor U17467 (N_17467,N_7535,N_11033);
nand U17468 (N_17468,N_7204,N_10354);
nor U17469 (N_17469,N_10775,N_6937);
xnor U17470 (N_17470,N_11718,N_7391);
nand U17471 (N_17471,N_12090,N_7011);
or U17472 (N_17472,N_9569,N_11654);
and U17473 (N_17473,N_11963,N_6964);
or U17474 (N_17474,N_8481,N_9105);
or U17475 (N_17475,N_8154,N_12443);
nor U17476 (N_17476,N_10563,N_6267);
xor U17477 (N_17477,N_9143,N_11435);
xnor U17478 (N_17478,N_6309,N_7931);
xor U17479 (N_17479,N_7423,N_7661);
or U17480 (N_17480,N_11571,N_9311);
and U17481 (N_17481,N_9118,N_11629);
or U17482 (N_17482,N_12322,N_10365);
nand U17483 (N_17483,N_8682,N_10737);
nor U17484 (N_17484,N_9632,N_7452);
xor U17485 (N_17485,N_6726,N_11138);
xor U17486 (N_17486,N_8022,N_8185);
or U17487 (N_17487,N_9734,N_12372);
nand U17488 (N_17488,N_6840,N_7437);
and U17489 (N_17489,N_11951,N_6554);
and U17490 (N_17490,N_11620,N_9900);
and U17491 (N_17491,N_11539,N_9147);
nor U17492 (N_17492,N_6649,N_10703);
nor U17493 (N_17493,N_11725,N_9692);
xnor U17494 (N_17494,N_8924,N_11845);
or U17495 (N_17495,N_12011,N_7784);
or U17496 (N_17496,N_6554,N_12429);
and U17497 (N_17497,N_6620,N_9667);
xor U17498 (N_17498,N_11649,N_11934);
nand U17499 (N_17499,N_11874,N_7503);
xor U17500 (N_17500,N_7365,N_11533);
and U17501 (N_17501,N_9076,N_8262);
and U17502 (N_17502,N_10523,N_7573);
nand U17503 (N_17503,N_6825,N_12015);
nand U17504 (N_17504,N_8519,N_7847);
nor U17505 (N_17505,N_9896,N_10077);
xnor U17506 (N_17506,N_8427,N_6499);
and U17507 (N_17507,N_12456,N_9066);
and U17508 (N_17508,N_9262,N_7559);
nand U17509 (N_17509,N_10574,N_8082);
nand U17510 (N_17510,N_12000,N_7658);
and U17511 (N_17511,N_7503,N_12041);
nand U17512 (N_17512,N_7309,N_9863);
xor U17513 (N_17513,N_9276,N_6828);
xor U17514 (N_17514,N_10519,N_8711);
xor U17515 (N_17515,N_8021,N_8224);
or U17516 (N_17516,N_7252,N_6322);
and U17517 (N_17517,N_10094,N_6509);
xor U17518 (N_17518,N_6468,N_6833);
nand U17519 (N_17519,N_7703,N_7585);
xnor U17520 (N_17520,N_9362,N_9092);
or U17521 (N_17521,N_7279,N_8887);
nor U17522 (N_17522,N_9580,N_11900);
nand U17523 (N_17523,N_7800,N_11057);
nor U17524 (N_17524,N_9808,N_9514);
nand U17525 (N_17525,N_11886,N_9782);
and U17526 (N_17526,N_6300,N_10218);
nor U17527 (N_17527,N_9126,N_10531);
nand U17528 (N_17528,N_9447,N_7597);
and U17529 (N_17529,N_10250,N_10454);
or U17530 (N_17530,N_11166,N_10636);
or U17531 (N_17531,N_11765,N_6471);
xor U17532 (N_17532,N_11242,N_12224);
nand U17533 (N_17533,N_12233,N_8023);
and U17534 (N_17534,N_9510,N_6431);
nand U17535 (N_17535,N_12021,N_7376);
nand U17536 (N_17536,N_10799,N_6468);
and U17537 (N_17537,N_11274,N_10425);
nor U17538 (N_17538,N_9289,N_12151);
xnor U17539 (N_17539,N_10007,N_8735);
xor U17540 (N_17540,N_11264,N_8684);
nand U17541 (N_17541,N_9585,N_9858);
xor U17542 (N_17542,N_11662,N_6453);
xor U17543 (N_17543,N_7106,N_9359);
nand U17544 (N_17544,N_6363,N_7459);
nand U17545 (N_17545,N_7340,N_9144);
xnor U17546 (N_17546,N_8124,N_7664);
nor U17547 (N_17547,N_8703,N_12415);
and U17548 (N_17548,N_11623,N_6980);
nand U17549 (N_17549,N_12139,N_10638);
nor U17550 (N_17550,N_9238,N_11283);
nor U17551 (N_17551,N_8534,N_9231);
and U17552 (N_17552,N_10797,N_7459);
or U17553 (N_17553,N_12270,N_7945);
xor U17554 (N_17554,N_11574,N_12042);
xor U17555 (N_17555,N_6614,N_10815);
xor U17556 (N_17556,N_10004,N_7435);
or U17557 (N_17557,N_12008,N_7644);
nor U17558 (N_17558,N_8484,N_9534);
nand U17559 (N_17559,N_6376,N_9284);
and U17560 (N_17560,N_7522,N_12465);
or U17561 (N_17561,N_9941,N_9846);
nor U17562 (N_17562,N_7834,N_11921);
nand U17563 (N_17563,N_7199,N_9560);
and U17564 (N_17564,N_6250,N_9989);
and U17565 (N_17565,N_11889,N_6823);
nand U17566 (N_17566,N_11516,N_9264);
nand U17567 (N_17567,N_8226,N_9429);
xnor U17568 (N_17568,N_7905,N_11332);
and U17569 (N_17569,N_7121,N_11140);
nor U17570 (N_17570,N_8257,N_8382);
or U17571 (N_17571,N_6714,N_7418);
nand U17572 (N_17572,N_7326,N_10116);
xnor U17573 (N_17573,N_7526,N_8600);
and U17574 (N_17574,N_9290,N_10605);
nand U17575 (N_17575,N_6686,N_11844);
or U17576 (N_17576,N_6308,N_7401);
nor U17577 (N_17577,N_10170,N_9236);
and U17578 (N_17578,N_10852,N_7364);
xnor U17579 (N_17579,N_7986,N_6822);
nor U17580 (N_17580,N_9812,N_10859);
or U17581 (N_17581,N_6300,N_9681);
nor U17582 (N_17582,N_7815,N_6967);
nand U17583 (N_17583,N_10169,N_12037);
nor U17584 (N_17584,N_9208,N_11886);
xnor U17585 (N_17585,N_8124,N_12409);
xor U17586 (N_17586,N_12109,N_12283);
nor U17587 (N_17587,N_12169,N_7861);
and U17588 (N_17588,N_9668,N_9704);
xor U17589 (N_17589,N_7795,N_7392);
xor U17590 (N_17590,N_7150,N_9695);
nor U17591 (N_17591,N_6804,N_7945);
and U17592 (N_17592,N_10995,N_9564);
xor U17593 (N_17593,N_7782,N_9320);
nand U17594 (N_17594,N_10471,N_10617);
nand U17595 (N_17595,N_10839,N_9109);
and U17596 (N_17596,N_8267,N_11774);
nor U17597 (N_17597,N_10766,N_6785);
nand U17598 (N_17598,N_7094,N_9029);
xnor U17599 (N_17599,N_8626,N_11908);
nand U17600 (N_17600,N_9938,N_10953);
or U17601 (N_17601,N_10091,N_7885);
xnor U17602 (N_17602,N_7669,N_6914);
xnor U17603 (N_17603,N_6966,N_11534);
xnor U17604 (N_17604,N_7294,N_7482);
and U17605 (N_17605,N_10743,N_7711);
nor U17606 (N_17606,N_10141,N_12456);
nor U17607 (N_17607,N_8121,N_9185);
nand U17608 (N_17608,N_10581,N_8322);
xor U17609 (N_17609,N_8600,N_9807);
nor U17610 (N_17610,N_9332,N_11253);
xnor U17611 (N_17611,N_6805,N_8693);
xor U17612 (N_17612,N_9347,N_10633);
nand U17613 (N_17613,N_8256,N_12178);
or U17614 (N_17614,N_9790,N_8218);
nand U17615 (N_17615,N_12390,N_11567);
nand U17616 (N_17616,N_7312,N_9661);
nand U17617 (N_17617,N_10171,N_6851);
and U17618 (N_17618,N_10811,N_6347);
nand U17619 (N_17619,N_8415,N_11995);
or U17620 (N_17620,N_7543,N_8796);
xor U17621 (N_17621,N_6307,N_11270);
xor U17622 (N_17622,N_11164,N_10560);
and U17623 (N_17623,N_9348,N_8888);
or U17624 (N_17624,N_7745,N_9018);
nor U17625 (N_17625,N_8025,N_8588);
nor U17626 (N_17626,N_7079,N_6644);
and U17627 (N_17627,N_8341,N_12374);
xor U17628 (N_17628,N_12441,N_9108);
or U17629 (N_17629,N_9322,N_6804);
nand U17630 (N_17630,N_11932,N_6839);
nand U17631 (N_17631,N_12301,N_8667);
nand U17632 (N_17632,N_8664,N_10118);
nand U17633 (N_17633,N_12024,N_8863);
nor U17634 (N_17634,N_7924,N_6895);
nor U17635 (N_17635,N_6484,N_7833);
xnor U17636 (N_17636,N_12326,N_7931);
nand U17637 (N_17637,N_8681,N_11323);
xor U17638 (N_17638,N_10664,N_9392);
or U17639 (N_17639,N_6555,N_7712);
nand U17640 (N_17640,N_7039,N_7759);
nand U17641 (N_17641,N_9866,N_11643);
nand U17642 (N_17642,N_11060,N_9055);
and U17643 (N_17643,N_8182,N_12390);
xnor U17644 (N_17644,N_8932,N_12370);
nor U17645 (N_17645,N_11091,N_9408);
or U17646 (N_17646,N_8665,N_9469);
nor U17647 (N_17647,N_8381,N_11586);
or U17648 (N_17648,N_11692,N_11703);
xor U17649 (N_17649,N_9804,N_8973);
xor U17650 (N_17650,N_11490,N_8492);
nor U17651 (N_17651,N_8032,N_11907);
or U17652 (N_17652,N_8450,N_7802);
nor U17653 (N_17653,N_8597,N_9596);
nor U17654 (N_17654,N_8804,N_9991);
nor U17655 (N_17655,N_6353,N_11532);
and U17656 (N_17656,N_12397,N_8849);
or U17657 (N_17657,N_11949,N_10395);
nand U17658 (N_17658,N_8063,N_7681);
nand U17659 (N_17659,N_9011,N_8829);
xor U17660 (N_17660,N_7181,N_8576);
nand U17661 (N_17661,N_6456,N_6634);
or U17662 (N_17662,N_6987,N_6481);
xnor U17663 (N_17663,N_10400,N_11892);
and U17664 (N_17664,N_7966,N_7311);
xor U17665 (N_17665,N_11820,N_11731);
and U17666 (N_17666,N_11476,N_11338);
xnor U17667 (N_17667,N_10053,N_11356);
and U17668 (N_17668,N_8618,N_10132);
and U17669 (N_17669,N_6579,N_10349);
and U17670 (N_17670,N_6701,N_9551);
xor U17671 (N_17671,N_8876,N_7424);
or U17672 (N_17672,N_11907,N_11911);
and U17673 (N_17673,N_8597,N_6758);
nor U17674 (N_17674,N_11364,N_10776);
nand U17675 (N_17675,N_6369,N_6378);
nor U17676 (N_17676,N_7678,N_8548);
and U17677 (N_17677,N_8909,N_9635);
and U17678 (N_17678,N_11800,N_8601);
or U17679 (N_17679,N_9246,N_8172);
nor U17680 (N_17680,N_6642,N_12204);
and U17681 (N_17681,N_9507,N_9657);
or U17682 (N_17682,N_12009,N_10451);
nand U17683 (N_17683,N_10910,N_10201);
or U17684 (N_17684,N_6665,N_9186);
nand U17685 (N_17685,N_7537,N_7143);
xnor U17686 (N_17686,N_11026,N_11930);
xor U17687 (N_17687,N_8985,N_12328);
nand U17688 (N_17688,N_7886,N_9668);
and U17689 (N_17689,N_6726,N_11481);
nor U17690 (N_17690,N_8296,N_8328);
xnor U17691 (N_17691,N_10474,N_7414);
or U17692 (N_17692,N_7354,N_12225);
nand U17693 (N_17693,N_9923,N_11801);
xor U17694 (N_17694,N_11786,N_8918);
nand U17695 (N_17695,N_10637,N_7499);
xnor U17696 (N_17696,N_8546,N_6642);
or U17697 (N_17697,N_11226,N_6918);
nor U17698 (N_17698,N_6999,N_12166);
and U17699 (N_17699,N_8201,N_8727);
and U17700 (N_17700,N_10057,N_9479);
nor U17701 (N_17701,N_11172,N_12391);
xor U17702 (N_17702,N_7973,N_8461);
nand U17703 (N_17703,N_6452,N_7656);
or U17704 (N_17704,N_6320,N_9514);
nand U17705 (N_17705,N_11810,N_7266);
xnor U17706 (N_17706,N_9282,N_11871);
nor U17707 (N_17707,N_7227,N_11555);
or U17708 (N_17708,N_11460,N_8989);
xnor U17709 (N_17709,N_8953,N_11459);
nor U17710 (N_17710,N_9863,N_11644);
and U17711 (N_17711,N_8919,N_10595);
or U17712 (N_17712,N_10535,N_6625);
xnor U17713 (N_17713,N_6904,N_11500);
xor U17714 (N_17714,N_11014,N_10353);
nor U17715 (N_17715,N_11880,N_10006);
or U17716 (N_17716,N_9103,N_11955);
nor U17717 (N_17717,N_9416,N_7007);
or U17718 (N_17718,N_11787,N_7242);
nand U17719 (N_17719,N_12172,N_11337);
or U17720 (N_17720,N_7053,N_7294);
and U17721 (N_17721,N_7768,N_9851);
xor U17722 (N_17722,N_9557,N_6856);
nor U17723 (N_17723,N_11764,N_6883);
nand U17724 (N_17724,N_12440,N_9487);
nor U17725 (N_17725,N_9814,N_6675);
nor U17726 (N_17726,N_9702,N_9717);
and U17727 (N_17727,N_12389,N_9376);
or U17728 (N_17728,N_8922,N_10394);
nor U17729 (N_17729,N_9578,N_8924);
nand U17730 (N_17730,N_6659,N_9015);
and U17731 (N_17731,N_8722,N_9252);
nand U17732 (N_17732,N_9405,N_11206);
or U17733 (N_17733,N_10917,N_10141);
or U17734 (N_17734,N_8716,N_7476);
and U17735 (N_17735,N_10150,N_8944);
nand U17736 (N_17736,N_10571,N_8188);
nand U17737 (N_17737,N_8006,N_10878);
nor U17738 (N_17738,N_9165,N_7647);
nor U17739 (N_17739,N_8369,N_6441);
nand U17740 (N_17740,N_6729,N_8729);
nand U17741 (N_17741,N_12096,N_10077);
xnor U17742 (N_17742,N_11571,N_11503);
xnor U17743 (N_17743,N_10721,N_8112);
nand U17744 (N_17744,N_6935,N_8920);
or U17745 (N_17745,N_9661,N_9142);
nor U17746 (N_17746,N_12333,N_8398);
or U17747 (N_17747,N_12130,N_7072);
xor U17748 (N_17748,N_11927,N_8004);
xnor U17749 (N_17749,N_9339,N_8553);
and U17750 (N_17750,N_10564,N_10369);
xor U17751 (N_17751,N_6535,N_12133);
and U17752 (N_17752,N_12119,N_9820);
or U17753 (N_17753,N_10913,N_10251);
and U17754 (N_17754,N_8743,N_9123);
nor U17755 (N_17755,N_7271,N_10735);
nor U17756 (N_17756,N_6829,N_8037);
or U17757 (N_17757,N_6646,N_8175);
nand U17758 (N_17758,N_11425,N_6437);
xnor U17759 (N_17759,N_8134,N_8457);
xnor U17760 (N_17760,N_7203,N_6774);
nand U17761 (N_17761,N_10254,N_6755);
nand U17762 (N_17762,N_10008,N_6400);
xor U17763 (N_17763,N_8072,N_8710);
xnor U17764 (N_17764,N_12242,N_11819);
nand U17765 (N_17765,N_7776,N_6973);
or U17766 (N_17766,N_8782,N_11700);
xnor U17767 (N_17767,N_6778,N_10954);
nor U17768 (N_17768,N_10590,N_6341);
and U17769 (N_17769,N_7977,N_6308);
nor U17770 (N_17770,N_11615,N_7562);
nand U17771 (N_17771,N_12074,N_12313);
nor U17772 (N_17772,N_7517,N_7042);
or U17773 (N_17773,N_11089,N_11685);
and U17774 (N_17774,N_11686,N_7572);
or U17775 (N_17775,N_10037,N_11621);
xnor U17776 (N_17776,N_11129,N_7524);
and U17777 (N_17777,N_11134,N_9134);
nor U17778 (N_17778,N_10037,N_8432);
xnor U17779 (N_17779,N_7086,N_12019);
nor U17780 (N_17780,N_10364,N_6548);
and U17781 (N_17781,N_6847,N_8453);
or U17782 (N_17782,N_9937,N_9235);
and U17783 (N_17783,N_10356,N_8378);
nor U17784 (N_17784,N_11836,N_11177);
and U17785 (N_17785,N_7419,N_8706);
and U17786 (N_17786,N_11991,N_6634);
or U17787 (N_17787,N_10400,N_9615);
and U17788 (N_17788,N_7389,N_6643);
nor U17789 (N_17789,N_8403,N_8810);
and U17790 (N_17790,N_10800,N_7699);
xnor U17791 (N_17791,N_7638,N_6304);
or U17792 (N_17792,N_12213,N_7023);
nand U17793 (N_17793,N_11474,N_11317);
or U17794 (N_17794,N_10050,N_7057);
nor U17795 (N_17795,N_11486,N_9911);
nor U17796 (N_17796,N_8090,N_9042);
and U17797 (N_17797,N_11009,N_10922);
or U17798 (N_17798,N_7797,N_8989);
nand U17799 (N_17799,N_6726,N_10700);
nor U17800 (N_17800,N_12050,N_8438);
or U17801 (N_17801,N_10181,N_11693);
nor U17802 (N_17802,N_11376,N_11580);
or U17803 (N_17803,N_11560,N_11628);
or U17804 (N_17804,N_11120,N_7574);
xor U17805 (N_17805,N_9295,N_12044);
xnor U17806 (N_17806,N_8398,N_8955);
nor U17807 (N_17807,N_10370,N_10264);
and U17808 (N_17808,N_11956,N_7710);
nor U17809 (N_17809,N_11262,N_8336);
nand U17810 (N_17810,N_9292,N_12203);
nand U17811 (N_17811,N_12243,N_10132);
or U17812 (N_17812,N_10732,N_9063);
nor U17813 (N_17813,N_8545,N_7666);
nand U17814 (N_17814,N_9380,N_11992);
xor U17815 (N_17815,N_8606,N_7401);
nand U17816 (N_17816,N_6784,N_6664);
nand U17817 (N_17817,N_9588,N_6605);
xnor U17818 (N_17818,N_12132,N_6749);
nor U17819 (N_17819,N_9910,N_11182);
and U17820 (N_17820,N_9330,N_9140);
xor U17821 (N_17821,N_9510,N_9801);
and U17822 (N_17822,N_10002,N_11585);
nand U17823 (N_17823,N_10617,N_7936);
xnor U17824 (N_17824,N_8418,N_6256);
nor U17825 (N_17825,N_6840,N_11090);
nor U17826 (N_17826,N_10520,N_8437);
xor U17827 (N_17827,N_6312,N_11834);
or U17828 (N_17828,N_12310,N_8406);
nor U17829 (N_17829,N_7778,N_9958);
nor U17830 (N_17830,N_11765,N_11918);
nand U17831 (N_17831,N_11276,N_10560);
xor U17832 (N_17832,N_10184,N_9310);
nor U17833 (N_17833,N_7307,N_10833);
xnor U17834 (N_17834,N_12108,N_9214);
nand U17835 (N_17835,N_10105,N_7451);
nor U17836 (N_17836,N_7363,N_11275);
and U17837 (N_17837,N_9504,N_6711);
nand U17838 (N_17838,N_11974,N_8665);
nor U17839 (N_17839,N_10479,N_10401);
nor U17840 (N_17840,N_8138,N_10838);
and U17841 (N_17841,N_9081,N_6968);
nand U17842 (N_17842,N_9900,N_6300);
nor U17843 (N_17843,N_7916,N_9185);
nor U17844 (N_17844,N_11666,N_7907);
xnor U17845 (N_17845,N_10377,N_8906);
or U17846 (N_17846,N_9126,N_6324);
xnor U17847 (N_17847,N_11217,N_7848);
nand U17848 (N_17848,N_7008,N_9290);
nand U17849 (N_17849,N_12164,N_11730);
and U17850 (N_17850,N_7405,N_8308);
and U17851 (N_17851,N_12329,N_12385);
or U17852 (N_17852,N_8862,N_10566);
nor U17853 (N_17853,N_8220,N_9719);
xnor U17854 (N_17854,N_11152,N_10888);
xnor U17855 (N_17855,N_6659,N_11795);
and U17856 (N_17856,N_9451,N_9093);
or U17857 (N_17857,N_9624,N_6275);
xnor U17858 (N_17858,N_11138,N_10280);
and U17859 (N_17859,N_9135,N_12372);
or U17860 (N_17860,N_12166,N_11940);
or U17861 (N_17861,N_7973,N_6966);
nand U17862 (N_17862,N_10720,N_10007);
nor U17863 (N_17863,N_11358,N_9403);
and U17864 (N_17864,N_10145,N_8569);
and U17865 (N_17865,N_7246,N_6855);
and U17866 (N_17866,N_12129,N_8433);
nor U17867 (N_17867,N_8349,N_7077);
nand U17868 (N_17868,N_11489,N_10519);
xor U17869 (N_17869,N_6996,N_11696);
and U17870 (N_17870,N_10149,N_9665);
nor U17871 (N_17871,N_6881,N_7024);
xor U17872 (N_17872,N_10052,N_8986);
nand U17873 (N_17873,N_10320,N_8253);
nor U17874 (N_17874,N_12410,N_8463);
or U17875 (N_17875,N_12179,N_11619);
and U17876 (N_17876,N_11793,N_10263);
nor U17877 (N_17877,N_6363,N_7420);
or U17878 (N_17878,N_7373,N_8453);
xor U17879 (N_17879,N_11706,N_10274);
nor U17880 (N_17880,N_11000,N_6497);
nand U17881 (N_17881,N_6924,N_9135);
and U17882 (N_17882,N_10139,N_11096);
nor U17883 (N_17883,N_7022,N_12365);
and U17884 (N_17884,N_7865,N_12124);
and U17885 (N_17885,N_10752,N_9875);
or U17886 (N_17886,N_11020,N_11322);
and U17887 (N_17887,N_9630,N_7219);
and U17888 (N_17888,N_10145,N_6578);
or U17889 (N_17889,N_9461,N_10632);
xor U17890 (N_17890,N_10417,N_9009);
xor U17891 (N_17891,N_10721,N_9840);
nand U17892 (N_17892,N_7107,N_9387);
or U17893 (N_17893,N_8332,N_12199);
or U17894 (N_17894,N_7012,N_7032);
and U17895 (N_17895,N_10843,N_7782);
and U17896 (N_17896,N_8497,N_7221);
xnor U17897 (N_17897,N_6736,N_8988);
nor U17898 (N_17898,N_10216,N_11544);
xnor U17899 (N_17899,N_8687,N_10240);
and U17900 (N_17900,N_11919,N_6903);
nand U17901 (N_17901,N_7182,N_6655);
nand U17902 (N_17902,N_9637,N_8365);
nor U17903 (N_17903,N_6254,N_12019);
nand U17904 (N_17904,N_10218,N_11283);
nor U17905 (N_17905,N_6890,N_11278);
nor U17906 (N_17906,N_7560,N_6806);
or U17907 (N_17907,N_9920,N_8663);
nor U17908 (N_17908,N_8310,N_10412);
and U17909 (N_17909,N_10576,N_9437);
or U17910 (N_17910,N_11747,N_8434);
xor U17911 (N_17911,N_10854,N_8029);
and U17912 (N_17912,N_7690,N_7199);
nand U17913 (N_17913,N_7632,N_10570);
nand U17914 (N_17914,N_12139,N_12159);
and U17915 (N_17915,N_12241,N_6551);
nand U17916 (N_17916,N_11972,N_7569);
or U17917 (N_17917,N_7055,N_11179);
or U17918 (N_17918,N_12176,N_11995);
nor U17919 (N_17919,N_11259,N_10479);
and U17920 (N_17920,N_11608,N_7975);
xor U17921 (N_17921,N_6641,N_10407);
xor U17922 (N_17922,N_7113,N_11770);
xnor U17923 (N_17923,N_10064,N_9911);
nor U17924 (N_17924,N_8486,N_9718);
and U17925 (N_17925,N_9784,N_7543);
and U17926 (N_17926,N_7986,N_7350);
nor U17927 (N_17927,N_11148,N_11378);
nor U17928 (N_17928,N_11135,N_10867);
or U17929 (N_17929,N_11987,N_8533);
or U17930 (N_17930,N_9911,N_11936);
xor U17931 (N_17931,N_10479,N_8707);
xor U17932 (N_17932,N_11356,N_11922);
xnor U17933 (N_17933,N_10754,N_8030);
nand U17934 (N_17934,N_10510,N_7267);
or U17935 (N_17935,N_10155,N_12488);
nor U17936 (N_17936,N_9614,N_8729);
and U17937 (N_17937,N_10307,N_11814);
nor U17938 (N_17938,N_10573,N_12091);
nand U17939 (N_17939,N_10347,N_6477);
or U17940 (N_17940,N_11818,N_12354);
and U17941 (N_17941,N_9665,N_12240);
nand U17942 (N_17942,N_9197,N_10693);
nand U17943 (N_17943,N_11561,N_11597);
nand U17944 (N_17944,N_7353,N_9223);
nand U17945 (N_17945,N_12417,N_9621);
xnor U17946 (N_17946,N_10136,N_8823);
nand U17947 (N_17947,N_10903,N_12399);
or U17948 (N_17948,N_11588,N_9143);
nor U17949 (N_17949,N_8755,N_11917);
and U17950 (N_17950,N_10466,N_11642);
nand U17951 (N_17951,N_9902,N_6691);
nor U17952 (N_17952,N_7837,N_6470);
or U17953 (N_17953,N_7276,N_10848);
nor U17954 (N_17954,N_9461,N_10416);
nor U17955 (N_17955,N_6986,N_10161);
nor U17956 (N_17956,N_7834,N_10617);
nand U17957 (N_17957,N_9374,N_11421);
or U17958 (N_17958,N_7739,N_10599);
or U17959 (N_17959,N_9930,N_7049);
nor U17960 (N_17960,N_9876,N_7005);
nor U17961 (N_17961,N_6886,N_8108);
and U17962 (N_17962,N_7213,N_7015);
or U17963 (N_17963,N_12099,N_7941);
or U17964 (N_17964,N_10815,N_6969);
xnor U17965 (N_17965,N_9552,N_10107);
xnor U17966 (N_17966,N_8862,N_10600);
xor U17967 (N_17967,N_9972,N_10650);
xor U17968 (N_17968,N_11660,N_8198);
xnor U17969 (N_17969,N_8218,N_6265);
nor U17970 (N_17970,N_11220,N_9034);
nand U17971 (N_17971,N_8943,N_10520);
and U17972 (N_17972,N_6820,N_10537);
and U17973 (N_17973,N_7694,N_9441);
or U17974 (N_17974,N_10415,N_9565);
xnor U17975 (N_17975,N_9557,N_10807);
or U17976 (N_17976,N_7350,N_6784);
nor U17977 (N_17977,N_9469,N_11570);
xnor U17978 (N_17978,N_11703,N_9686);
and U17979 (N_17979,N_8786,N_9049);
xor U17980 (N_17980,N_9347,N_6675);
xor U17981 (N_17981,N_10914,N_10478);
nand U17982 (N_17982,N_7573,N_10311);
and U17983 (N_17983,N_10705,N_7245);
nand U17984 (N_17984,N_10936,N_6780);
xnor U17985 (N_17985,N_7950,N_9065);
or U17986 (N_17986,N_11208,N_10791);
and U17987 (N_17987,N_8149,N_6365);
or U17988 (N_17988,N_11462,N_11796);
xnor U17989 (N_17989,N_8572,N_6737);
and U17990 (N_17990,N_8743,N_11140);
or U17991 (N_17991,N_11749,N_8103);
and U17992 (N_17992,N_6775,N_9573);
nand U17993 (N_17993,N_10943,N_8868);
nor U17994 (N_17994,N_7907,N_6841);
nor U17995 (N_17995,N_11361,N_9440);
nor U17996 (N_17996,N_12169,N_11450);
nor U17997 (N_17997,N_10631,N_11544);
and U17998 (N_17998,N_8519,N_7249);
nand U17999 (N_17999,N_11347,N_10060);
or U18000 (N_18000,N_6485,N_6569);
nor U18001 (N_18001,N_7045,N_8139);
or U18002 (N_18002,N_9537,N_12405);
nand U18003 (N_18003,N_8388,N_8155);
xor U18004 (N_18004,N_11440,N_12395);
and U18005 (N_18005,N_11654,N_8284);
nor U18006 (N_18006,N_7610,N_6910);
xor U18007 (N_18007,N_10528,N_11562);
or U18008 (N_18008,N_10770,N_8327);
and U18009 (N_18009,N_11627,N_8307);
and U18010 (N_18010,N_6276,N_6469);
or U18011 (N_18011,N_11148,N_7751);
xor U18012 (N_18012,N_7244,N_9702);
nand U18013 (N_18013,N_11118,N_10076);
xor U18014 (N_18014,N_10459,N_8487);
or U18015 (N_18015,N_12336,N_9514);
nor U18016 (N_18016,N_9270,N_8991);
and U18017 (N_18017,N_7446,N_12362);
nand U18018 (N_18018,N_9861,N_7054);
nand U18019 (N_18019,N_8898,N_11978);
nor U18020 (N_18020,N_11494,N_11344);
and U18021 (N_18021,N_10548,N_7345);
and U18022 (N_18022,N_8440,N_7550);
nand U18023 (N_18023,N_7881,N_12196);
xor U18024 (N_18024,N_8607,N_6858);
xnor U18025 (N_18025,N_9199,N_7864);
or U18026 (N_18026,N_11870,N_9092);
or U18027 (N_18027,N_10179,N_8132);
and U18028 (N_18028,N_8469,N_8531);
nand U18029 (N_18029,N_8190,N_10923);
and U18030 (N_18030,N_9502,N_11262);
or U18031 (N_18031,N_10656,N_6536);
or U18032 (N_18032,N_7232,N_8410);
nand U18033 (N_18033,N_7101,N_7062);
xor U18034 (N_18034,N_6847,N_8014);
and U18035 (N_18035,N_11683,N_12447);
xor U18036 (N_18036,N_12195,N_8052);
xor U18037 (N_18037,N_6590,N_7720);
or U18038 (N_18038,N_7158,N_6588);
xor U18039 (N_18039,N_10871,N_11707);
and U18040 (N_18040,N_12088,N_12228);
or U18041 (N_18041,N_9011,N_6413);
xor U18042 (N_18042,N_7468,N_9063);
and U18043 (N_18043,N_10744,N_7161);
xor U18044 (N_18044,N_10918,N_7195);
nand U18045 (N_18045,N_11114,N_9797);
nor U18046 (N_18046,N_8155,N_9939);
and U18047 (N_18047,N_8589,N_7412);
nand U18048 (N_18048,N_6822,N_7656);
nand U18049 (N_18049,N_11887,N_9729);
and U18050 (N_18050,N_12351,N_9974);
nor U18051 (N_18051,N_10523,N_7842);
nand U18052 (N_18052,N_11363,N_9104);
nor U18053 (N_18053,N_11589,N_7955);
and U18054 (N_18054,N_8336,N_10938);
nor U18055 (N_18055,N_8555,N_11890);
nand U18056 (N_18056,N_10730,N_9387);
nand U18057 (N_18057,N_6969,N_11464);
and U18058 (N_18058,N_10791,N_10147);
xor U18059 (N_18059,N_9211,N_6304);
nand U18060 (N_18060,N_7887,N_11273);
nor U18061 (N_18061,N_12339,N_7123);
nor U18062 (N_18062,N_9698,N_10298);
nand U18063 (N_18063,N_6474,N_10046);
nand U18064 (N_18064,N_11422,N_11734);
nand U18065 (N_18065,N_11161,N_10858);
xnor U18066 (N_18066,N_8913,N_10518);
xnor U18067 (N_18067,N_10077,N_9137);
or U18068 (N_18068,N_10114,N_8499);
xor U18069 (N_18069,N_10883,N_11364);
or U18070 (N_18070,N_10806,N_8407);
or U18071 (N_18071,N_9954,N_6495);
and U18072 (N_18072,N_6569,N_9849);
nand U18073 (N_18073,N_11546,N_11816);
nand U18074 (N_18074,N_9470,N_8261);
or U18075 (N_18075,N_6552,N_9516);
and U18076 (N_18076,N_8785,N_10314);
nand U18077 (N_18077,N_6883,N_9338);
and U18078 (N_18078,N_10766,N_8255);
nor U18079 (N_18079,N_6695,N_8933);
xor U18080 (N_18080,N_10779,N_7221);
or U18081 (N_18081,N_7250,N_7892);
nor U18082 (N_18082,N_8465,N_8038);
and U18083 (N_18083,N_8869,N_12252);
nand U18084 (N_18084,N_11275,N_9939);
nand U18085 (N_18085,N_10474,N_7482);
xnor U18086 (N_18086,N_9060,N_10844);
or U18087 (N_18087,N_9883,N_9785);
or U18088 (N_18088,N_9665,N_10391);
or U18089 (N_18089,N_7792,N_8984);
xnor U18090 (N_18090,N_9153,N_12450);
nor U18091 (N_18091,N_11768,N_10968);
or U18092 (N_18092,N_10316,N_9642);
xnor U18093 (N_18093,N_12468,N_7940);
and U18094 (N_18094,N_7790,N_12002);
or U18095 (N_18095,N_7366,N_8061);
nor U18096 (N_18096,N_9661,N_10624);
nand U18097 (N_18097,N_9316,N_8642);
nor U18098 (N_18098,N_7863,N_8576);
and U18099 (N_18099,N_6870,N_7715);
xor U18100 (N_18100,N_8903,N_11208);
or U18101 (N_18101,N_7351,N_8950);
nand U18102 (N_18102,N_11824,N_8417);
xnor U18103 (N_18103,N_11754,N_11990);
xor U18104 (N_18104,N_10595,N_11555);
nor U18105 (N_18105,N_10434,N_9739);
nor U18106 (N_18106,N_7838,N_7189);
xor U18107 (N_18107,N_9424,N_10203);
xor U18108 (N_18108,N_6419,N_7645);
xor U18109 (N_18109,N_9545,N_10188);
and U18110 (N_18110,N_10465,N_8038);
xnor U18111 (N_18111,N_7054,N_8767);
nor U18112 (N_18112,N_8452,N_9592);
xor U18113 (N_18113,N_6409,N_9960);
nor U18114 (N_18114,N_12191,N_10749);
and U18115 (N_18115,N_7139,N_11290);
xor U18116 (N_18116,N_10750,N_6578);
nor U18117 (N_18117,N_8569,N_10386);
or U18118 (N_18118,N_7797,N_9401);
or U18119 (N_18119,N_7399,N_8030);
nand U18120 (N_18120,N_9085,N_11796);
nand U18121 (N_18121,N_12182,N_6532);
nand U18122 (N_18122,N_12223,N_12395);
nand U18123 (N_18123,N_9876,N_7105);
nand U18124 (N_18124,N_7909,N_8557);
nor U18125 (N_18125,N_10563,N_9673);
and U18126 (N_18126,N_11048,N_10511);
or U18127 (N_18127,N_9956,N_11539);
nor U18128 (N_18128,N_7137,N_9129);
or U18129 (N_18129,N_8823,N_10084);
nor U18130 (N_18130,N_12226,N_10399);
nand U18131 (N_18131,N_7849,N_7807);
or U18132 (N_18132,N_10012,N_8780);
and U18133 (N_18133,N_11408,N_11497);
nor U18134 (N_18134,N_11672,N_7280);
xor U18135 (N_18135,N_8425,N_9015);
or U18136 (N_18136,N_12466,N_8933);
nor U18137 (N_18137,N_11523,N_9345);
or U18138 (N_18138,N_7566,N_9634);
nor U18139 (N_18139,N_10003,N_7154);
nand U18140 (N_18140,N_11796,N_7732);
or U18141 (N_18141,N_7871,N_8110);
or U18142 (N_18142,N_10907,N_10546);
or U18143 (N_18143,N_8245,N_7771);
or U18144 (N_18144,N_11048,N_6845);
nand U18145 (N_18145,N_6989,N_7435);
nor U18146 (N_18146,N_12432,N_9721);
and U18147 (N_18147,N_7082,N_11901);
or U18148 (N_18148,N_12230,N_10603);
and U18149 (N_18149,N_9981,N_12160);
nor U18150 (N_18150,N_10104,N_10389);
nand U18151 (N_18151,N_12255,N_7088);
nand U18152 (N_18152,N_11305,N_9987);
or U18153 (N_18153,N_10886,N_10074);
nand U18154 (N_18154,N_7316,N_8613);
nand U18155 (N_18155,N_8367,N_11916);
nor U18156 (N_18156,N_11338,N_9677);
and U18157 (N_18157,N_11109,N_8223);
and U18158 (N_18158,N_6813,N_8064);
or U18159 (N_18159,N_11031,N_12311);
xor U18160 (N_18160,N_9565,N_11265);
nor U18161 (N_18161,N_8623,N_6542);
nor U18162 (N_18162,N_11269,N_10601);
or U18163 (N_18163,N_6690,N_10048);
nand U18164 (N_18164,N_12174,N_6982);
or U18165 (N_18165,N_10558,N_7268);
nor U18166 (N_18166,N_7894,N_7025);
or U18167 (N_18167,N_9443,N_11569);
nor U18168 (N_18168,N_9139,N_8639);
and U18169 (N_18169,N_7581,N_11553);
nand U18170 (N_18170,N_8246,N_11366);
nor U18171 (N_18171,N_6566,N_12410);
xor U18172 (N_18172,N_9130,N_9023);
nand U18173 (N_18173,N_11745,N_7250);
or U18174 (N_18174,N_11645,N_8763);
or U18175 (N_18175,N_8018,N_6473);
and U18176 (N_18176,N_7826,N_12381);
nor U18177 (N_18177,N_7085,N_9944);
and U18178 (N_18178,N_7534,N_11518);
and U18179 (N_18179,N_12435,N_12056);
nand U18180 (N_18180,N_11521,N_9656);
xnor U18181 (N_18181,N_11497,N_9138);
and U18182 (N_18182,N_11027,N_11857);
or U18183 (N_18183,N_9778,N_10099);
xnor U18184 (N_18184,N_9180,N_6716);
and U18185 (N_18185,N_8222,N_12356);
xnor U18186 (N_18186,N_7313,N_8125);
or U18187 (N_18187,N_7258,N_9692);
and U18188 (N_18188,N_8303,N_10004);
and U18189 (N_18189,N_7958,N_7874);
xor U18190 (N_18190,N_10564,N_12461);
and U18191 (N_18191,N_9597,N_6369);
xor U18192 (N_18192,N_10378,N_6923);
nand U18193 (N_18193,N_7829,N_10195);
or U18194 (N_18194,N_9888,N_10021);
nand U18195 (N_18195,N_6857,N_7267);
xnor U18196 (N_18196,N_7303,N_6418);
nand U18197 (N_18197,N_12013,N_12054);
and U18198 (N_18198,N_10541,N_8955);
or U18199 (N_18199,N_9412,N_7494);
and U18200 (N_18200,N_7207,N_10910);
xnor U18201 (N_18201,N_12176,N_8455);
xor U18202 (N_18202,N_8664,N_11219);
xor U18203 (N_18203,N_11081,N_9399);
xor U18204 (N_18204,N_6472,N_9337);
and U18205 (N_18205,N_9608,N_9375);
or U18206 (N_18206,N_8389,N_11175);
or U18207 (N_18207,N_7490,N_6877);
and U18208 (N_18208,N_6440,N_8741);
nor U18209 (N_18209,N_9923,N_7098);
nand U18210 (N_18210,N_11723,N_11286);
nand U18211 (N_18211,N_8350,N_7360);
xor U18212 (N_18212,N_10923,N_11565);
nor U18213 (N_18213,N_7064,N_6497);
xor U18214 (N_18214,N_11946,N_10663);
xnor U18215 (N_18215,N_11355,N_9821);
xor U18216 (N_18216,N_8376,N_6918);
nand U18217 (N_18217,N_8806,N_8364);
nor U18218 (N_18218,N_7297,N_7391);
and U18219 (N_18219,N_7580,N_9775);
nand U18220 (N_18220,N_6309,N_8859);
nor U18221 (N_18221,N_6517,N_11924);
and U18222 (N_18222,N_8128,N_11127);
nor U18223 (N_18223,N_10193,N_9549);
nand U18224 (N_18224,N_7421,N_7553);
nand U18225 (N_18225,N_10762,N_7210);
or U18226 (N_18226,N_11296,N_7482);
nor U18227 (N_18227,N_12221,N_10056);
nor U18228 (N_18228,N_10356,N_9649);
xnor U18229 (N_18229,N_11639,N_6832);
nor U18230 (N_18230,N_7982,N_6883);
or U18231 (N_18231,N_7365,N_7331);
xnor U18232 (N_18232,N_9970,N_9618);
xor U18233 (N_18233,N_9945,N_8214);
nand U18234 (N_18234,N_7090,N_6268);
and U18235 (N_18235,N_6818,N_10990);
nand U18236 (N_18236,N_6360,N_9894);
xnor U18237 (N_18237,N_7028,N_12036);
nand U18238 (N_18238,N_10897,N_8928);
nand U18239 (N_18239,N_10909,N_12468);
xor U18240 (N_18240,N_10476,N_6571);
xor U18241 (N_18241,N_10690,N_11246);
and U18242 (N_18242,N_12438,N_9756);
or U18243 (N_18243,N_11605,N_11508);
nand U18244 (N_18244,N_9019,N_11889);
nor U18245 (N_18245,N_6879,N_10059);
nand U18246 (N_18246,N_11788,N_12074);
xor U18247 (N_18247,N_9772,N_9393);
or U18248 (N_18248,N_6910,N_8761);
or U18249 (N_18249,N_6322,N_6971);
or U18250 (N_18250,N_9430,N_9933);
nand U18251 (N_18251,N_10198,N_8645);
nor U18252 (N_18252,N_7277,N_10513);
xnor U18253 (N_18253,N_9360,N_8482);
nand U18254 (N_18254,N_10438,N_8046);
nor U18255 (N_18255,N_11239,N_12005);
or U18256 (N_18256,N_6628,N_8597);
xnor U18257 (N_18257,N_7228,N_7335);
and U18258 (N_18258,N_8360,N_10118);
xnor U18259 (N_18259,N_12431,N_11694);
or U18260 (N_18260,N_6547,N_6594);
xor U18261 (N_18261,N_7071,N_8867);
nor U18262 (N_18262,N_11179,N_9888);
and U18263 (N_18263,N_6730,N_11440);
and U18264 (N_18264,N_6942,N_6465);
and U18265 (N_18265,N_9805,N_10305);
or U18266 (N_18266,N_7142,N_9035);
nand U18267 (N_18267,N_8310,N_10246);
and U18268 (N_18268,N_10315,N_9388);
and U18269 (N_18269,N_7784,N_7783);
and U18270 (N_18270,N_8797,N_11453);
nand U18271 (N_18271,N_8619,N_9148);
nand U18272 (N_18272,N_12223,N_8551);
xor U18273 (N_18273,N_8050,N_7407);
xnor U18274 (N_18274,N_11680,N_9251);
nand U18275 (N_18275,N_12195,N_9560);
nor U18276 (N_18276,N_8935,N_8083);
or U18277 (N_18277,N_9933,N_6836);
and U18278 (N_18278,N_9028,N_10935);
or U18279 (N_18279,N_7246,N_9312);
or U18280 (N_18280,N_6738,N_11106);
nor U18281 (N_18281,N_9053,N_11606);
and U18282 (N_18282,N_6668,N_8121);
or U18283 (N_18283,N_10117,N_6805);
nand U18284 (N_18284,N_8540,N_11467);
and U18285 (N_18285,N_10475,N_6659);
nor U18286 (N_18286,N_11277,N_6275);
or U18287 (N_18287,N_7887,N_7686);
nand U18288 (N_18288,N_12112,N_6619);
nand U18289 (N_18289,N_6986,N_7001);
or U18290 (N_18290,N_10010,N_7114);
and U18291 (N_18291,N_12002,N_7806);
and U18292 (N_18292,N_8268,N_6264);
or U18293 (N_18293,N_11166,N_7667);
nand U18294 (N_18294,N_6877,N_11714);
xnor U18295 (N_18295,N_10667,N_11293);
nor U18296 (N_18296,N_9059,N_9113);
nor U18297 (N_18297,N_9692,N_9898);
nor U18298 (N_18298,N_10069,N_8740);
and U18299 (N_18299,N_9462,N_6770);
and U18300 (N_18300,N_9997,N_8430);
xor U18301 (N_18301,N_12046,N_9436);
and U18302 (N_18302,N_11433,N_9440);
nor U18303 (N_18303,N_7022,N_8690);
or U18304 (N_18304,N_9467,N_8403);
or U18305 (N_18305,N_7555,N_9716);
and U18306 (N_18306,N_12480,N_11529);
and U18307 (N_18307,N_9204,N_7725);
xor U18308 (N_18308,N_8907,N_8732);
nor U18309 (N_18309,N_11925,N_10062);
or U18310 (N_18310,N_6623,N_11085);
or U18311 (N_18311,N_10420,N_6706);
xnor U18312 (N_18312,N_8229,N_10203);
nand U18313 (N_18313,N_9675,N_8100);
and U18314 (N_18314,N_9182,N_8453);
and U18315 (N_18315,N_10733,N_11584);
nor U18316 (N_18316,N_7775,N_10946);
or U18317 (N_18317,N_10232,N_9220);
and U18318 (N_18318,N_10724,N_6481);
nor U18319 (N_18319,N_6649,N_10113);
nor U18320 (N_18320,N_7245,N_8298);
or U18321 (N_18321,N_8780,N_8945);
nor U18322 (N_18322,N_9537,N_12270);
nand U18323 (N_18323,N_6393,N_7697);
or U18324 (N_18324,N_7906,N_6363);
or U18325 (N_18325,N_12121,N_9337);
and U18326 (N_18326,N_11903,N_11074);
xnor U18327 (N_18327,N_9471,N_7091);
and U18328 (N_18328,N_10815,N_7996);
nand U18329 (N_18329,N_10853,N_8871);
xnor U18330 (N_18330,N_9642,N_7558);
nor U18331 (N_18331,N_7949,N_9468);
nand U18332 (N_18332,N_7272,N_8461);
and U18333 (N_18333,N_6820,N_6865);
nor U18334 (N_18334,N_11832,N_9993);
nor U18335 (N_18335,N_7902,N_6763);
or U18336 (N_18336,N_10869,N_8191);
or U18337 (N_18337,N_6634,N_8496);
or U18338 (N_18338,N_10573,N_8558);
nor U18339 (N_18339,N_10673,N_9735);
nand U18340 (N_18340,N_6556,N_7851);
xnor U18341 (N_18341,N_11925,N_9955);
xor U18342 (N_18342,N_6631,N_9896);
and U18343 (N_18343,N_11258,N_6358);
xnor U18344 (N_18344,N_11862,N_9835);
or U18345 (N_18345,N_8509,N_6834);
or U18346 (N_18346,N_9839,N_7773);
or U18347 (N_18347,N_11441,N_11931);
nor U18348 (N_18348,N_7495,N_8565);
nor U18349 (N_18349,N_8515,N_8687);
or U18350 (N_18350,N_8550,N_10527);
nor U18351 (N_18351,N_9813,N_8127);
and U18352 (N_18352,N_10558,N_9768);
nand U18353 (N_18353,N_11796,N_10307);
nand U18354 (N_18354,N_7279,N_7259);
xor U18355 (N_18355,N_11714,N_9383);
nor U18356 (N_18356,N_9825,N_11505);
nor U18357 (N_18357,N_11045,N_6585);
and U18358 (N_18358,N_8929,N_11987);
and U18359 (N_18359,N_11202,N_6555);
nand U18360 (N_18360,N_10880,N_9602);
nand U18361 (N_18361,N_10439,N_11666);
xnor U18362 (N_18362,N_11080,N_9173);
nand U18363 (N_18363,N_11436,N_12286);
and U18364 (N_18364,N_12469,N_7830);
or U18365 (N_18365,N_7743,N_8268);
or U18366 (N_18366,N_9921,N_10167);
nand U18367 (N_18367,N_10280,N_7382);
or U18368 (N_18368,N_11735,N_9412);
or U18369 (N_18369,N_11117,N_6668);
and U18370 (N_18370,N_7258,N_11575);
or U18371 (N_18371,N_6677,N_7979);
xor U18372 (N_18372,N_10324,N_9424);
and U18373 (N_18373,N_8215,N_9449);
or U18374 (N_18374,N_6646,N_11272);
nor U18375 (N_18375,N_6487,N_11074);
or U18376 (N_18376,N_11456,N_11280);
nand U18377 (N_18377,N_10685,N_11530);
nor U18378 (N_18378,N_10461,N_8698);
nand U18379 (N_18379,N_7084,N_10437);
xor U18380 (N_18380,N_11492,N_11018);
or U18381 (N_18381,N_11458,N_6909);
xnor U18382 (N_18382,N_8285,N_10072);
xnor U18383 (N_18383,N_9324,N_6440);
xor U18384 (N_18384,N_11638,N_12065);
xnor U18385 (N_18385,N_6575,N_8480);
xnor U18386 (N_18386,N_6310,N_8500);
xnor U18387 (N_18387,N_8167,N_9624);
xnor U18388 (N_18388,N_9136,N_6948);
and U18389 (N_18389,N_12072,N_8920);
and U18390 (N_18390,N_6735,N_8451);
nand U18391 (N_18391,N_8261,N_7869);
and U18392 (N_18392,N_12210,N_8616);
nand U18393 (N_18393,N_7152,N_6944);
nand U18394 (N_18394,N_8864,N_12356);
nand U18395 (N_18395,N_11127,N_9054);
or U18396 (N_18396,N_8542,N_8471);
nor U18397 (N_18397,N_8348,N_11276);
and U18398 (N_18398,N_10058,N_8016);
xnor U18399 (N_18399,N_6550,N_11246);
nand U18400 (N_18400,N_7757,N_8619);
and U18401 (N_18401,N_11655,N_8159);
xor U18402 (N_18402,N_10910,N_11641);
and U18403 (N_18403,N_11648,N_11828);
or U18404 (N_18404,N_7683,N_6389);
xnor U18405 (N_18405,N_6417,N_9941);
xnor U18406 (N_18406,N_9424,N_8338);
nor U18407 (N_18407,N_11811,N_9833);
and U18408 (N_18408,N_10599,N_8054);
xor U18409 (N_18409,N_7570,N_6398);
or U18410 (N_18410,N_7590,N_9714);
or U18411 (N_18411,N_6379,N_7328);
nor U18412 (N_18412,N_9949,N_7553);
nand U18413 (N_18413,N_6646,N_9430);
or U18414 (N_18414,N_10752,N_6409);
xor U18415 (N_18415,N_8327,N_6480);
nor U18416 (N_18416,N_11324,N_9299);
nand U18417 (N_18417,N_12350,N_6521);
or U18418 (N_18418,N_9051,N_12185);
or U18419 (N_18419,N_12497,N_7496);
xor U18420 (N_18420,N_11876,N_11923);
xnor U18421 (N_18421,N_9627,N_10902);
nand U18422 (N_18422,N_11493,N_9404);
xnor U18423 (N_18423,N_11790,N_8524);
or U18424 (N_18424,N_11784,N_10072);
xor U18425 (N_18425,N_11981,N_6609);
or U18426 (N_18426,N_9669,N_8583);
nand U18427 (N_18427,N_6365,N_6331);
or U18428 (N_18428,N_10209,N_11344);
nand U18429 (N_18429,N_8239,N_10473);
and U18430 (N_18430,N_9790,N_7714);
xnor U18431 (N_18431,N_7152,N_11640);
or U18432 (N_18432,N_7743,N_7860);
or U18433 (N_18433,N_11105,N_7418);
and U18434 (N_18434,N_10926,N_7259);
and U18435 (N_18435,N_8210,N_10608);
nand U18436 (N_18436,N_7815,N_11595);
nand U18437 (N_18437,N_12393,N_10110);
and U18438 (N_18438,N_9935,N_9769);
nor U18439 (N_18439,N_6333,N_6638);
xor U18440 (N_18440,N_10728,N_9673);
xor U18441 (N_18441,N_11307,N_12286);
and U18442 (N_18442,N_7397,N_8932);
nor U18443 (N_18443,N_10472,N_6481);
nand U18444 (N_18444,N_12447,N_10332);
or U18445 (N_18445,N_7270,N_12489);
nand U18446 (N_18446,N_9287,N_8414);
nor U18447 (N_18447,N_12018,N_6826);
or U18448 (N_18448,N_6734,N_6501);
and U18449 (N_18449,N_11167,N_6301);
and U18450 (N_18450,N_6737,N_11502);
nand U18451 (N_18451,N_11761,N_12429);
xor U18452 (N_18452,N_7796,N_7322);
xnor U18453 (N_18453,N_9775,N_7135);
nor U18454 (N_18454,N_11323,N_10112);
nor U18455 (N_18455,N_7494,N_12332);
and U18456 (N_18456,N_8817,N_8053);
and U18457 (N_18457,N_12393,N_11197);
nor U18458 (N_18458,N_9814,N_6626);
xnor U18459 (N_18459,N_11472,N_9332);
or U18460 (N_18460,N_9833,N_10282);
nor U18461 (N_18461,N_8426,N_11297);
or U18462 (N_18462,N_6686,N_8206);
nand U18463 (N_18463,N_11738,N_8310);
nand U18464 (N_18464,N_6451,N_8776);
nand U18465 (N_18465,N_6673,N_8710);
xnor U18466 (N_18466,N_11018,N_11137);
xnor U18467 (N_18467,N_7819,N_9004);
nand U18468 (N_18468,N_11468,N_10211);
xor U18469 (N_18469,N_8989,N_9222);
xor U18470 (N_18470,N_6424,N_6468);
xor U18471 (N_18471,N_9033,N_10632);
xor U18472 (N_18472,N_11691,N_8976);
and U18473 (N_18473,N_8221,N_10398);
nand U18474 (N_18474,N_11644,N_11614);
or U18475 (N_18475,N_6424,N_6554);
nor U18476 (N_18476,N_9527,N_9218);
xor U18477 (N_18477,N_9977,N_9118);
nand U18478 (N_18478,N_10232,N_12387);
nor U18479 (N_18479,N_6529,N_8923);
nor U18480 (N_18480,N_12493,N_8005);
xor U18481 (N_18481,N_11367,N_11306);
nor U18482 (N_18482,N_7744,N_8697);
nor U18483 (N_18483,N_6836,N_8253);
xor U18484 (N_18484,N_11565,N_7595);
nand U18485 (N_18485,N_7935,N_7293);
xor U18486 (N_18486,N_7592,N_9778);
nand U18487 (N_18487,N_6380,N_10532);
and U18488 (N_18488,N_8775,N_7845);
nor U18489 (N_18489,N_8776,N_10230);
nand U18490 (N_18490,N_11218,N_7679);
nor U18491 (N_18491,N_11581,N_11191);
and U18492 (N_18492,N_8141,N_11997);
nor U18493 (N_18493,N_9371,N_9535);
xnor U18494 (N_18494,N_9233,N_7497);
and U18495 (N_18495,N_9847,N_8242);
or U18496 (N_18496,N_11674,N_9237);
nand U18497 (N_18497,N_11101,N_10964);
or U18498 (N_18498,N_10787,N_7617);
and U18499 (N_18499,N_12377,N_9244);
and U18500 (N_18500,N_8820,N_11301);
nand U18501 (N_18501,N_11934,N_10224);
xor U18502 (N_18502,N_8333,N_10429);
xor U18503 (N_18503,N_7417,N_10538);
or U18504 (N_18504,N_9275,N_11442);
nor U18505 (N_18505,N_10730,N_6390);
or U18506 (N_18506,N_7877,N_6507);
nor U18507 (N_18507,N_10392,N_7986);
or U18508 (N_18508,N_8190,N_11221);
and U18509 (N_18509,N_9372,N_8543);
or U18510 (N_18510,N_9219,N_7745);
and U18511 (N_18511,N_9797,N_6673);
nor U18512 (N_18512,N_12009,N_7639);
nand U18513 (N_18513,N_8979,N_8915);
nand U18514 (N_18514,N_11958,N_11043);
or U18515 (N_18515,N_10687,N_11900);
or U18516 (N_18516,N_7383,N_9776);
and U18517 (N_18517,N_6523,N_7943);
nand U18518 (N_18518,N_11495,N_10496);
or U18519 (N_18519,N_8157,N_9210);
or U18520 (N_18520,N_6587,N_6554);
and U18521 (N_18521,N_6743,N_10865);
xor U18522 (N_18522,N_6995,N_6648);
and U18523 (N_18523,N_10512,N_12486);
or U18524 (N_18524,N_8660,N_9486);
xnor U18525 (N_18525,N_10326,N_11536);
and U18526 (N_18526,N_7924,N_10106);
nand U18527 (N_18527,N_10169,N_10524);
nor U18528 (N_18528,N_7130,N_11296);
or U18529 (N_18529,N_7203,N_6986);
nand U18530 (N_18530,N_8384,N_10841);
nor U18531 (N_18531,N_9460,N_9097);
or U18532 (N_18532,N_10128,N_10508);
xnor U18533 (N_18533,N_7260,N_6897);
xor U18534 (N_18534,N_9744,N_8201);
and U18535 (N_18535,N_10855,N_10914);
or U18536 (N_18536,N_6474,N_8161);
or U18537 (N_18537,N_9596,N_7614);
and U18538 (N_18538,N_12461,N_10133);
and U18539 (N_18539,N_6985,N_6635);
nand U18540 (N_18540,N_7728,N_7603);
and U18541 (N_18541,N_6910,N_11555);
nor U18542 (N_18542,N_12310,N_7157);
nor U18543 (N_18543,N_10872,N_8338);
nor U18544 (N_18544,N_9375,N_12181);
xnor U18545 (N_18545,N_7085,N_10128);
and U18546 (N_18546,N_6528,N_9049);
nand U18547 (N_18547,N_7274,N_10443);
and U18548 (N_18548,N_7805,N_11944);
xor U18549 (N_18549,N_8635,N_9940);
and U18550 (N_18550,N_11310,N_11656);
or U18551 (N_18551,N_7483,N_9740);
and U18552 (N_18552,N_10960,N_10226);
or U18553 (N_18553,N_11181,N_9280);
nor U18554 (N_18554,N_6427,N_10447);
xor U18555 (N_18555,N_8867,N_11521);
nor U18556 (N_18556,N_6454,N_10011);
or U18557 (N_18557,N_11955,N_10428);
xnor U18558 (N_18558,N_11968,N_8601);
nand U18559 (N_18559,N_8632,N_7713);
nand U18560 (N_18560,N_6306,N_11836);
nand U18561 (N_18561,N_9637,N_10934);
nand U18562 (N_18562,N_11065,N_9310);
xor U18563 (N_18563,N_8486,N_9558);
nor U18564 (N_18564,N_11939,N_10400);
and U18565 (N_18565,N_12422,N_9062);
nand U18566 (N_18566,N_11713,N_11734);
or U18567 (N_18567,N_9471,N_7557);
and U18568 (N_18568,N_8949,N_9236);
nor U18569 (N_18569,N_9087,N_8555);
and U18570 (N_18570,N_11240,N_8335);
nor U18571 (N_18571,N_10237,N_8785);
xor U18572 (N_18572,N_11952,N_7604);
xnor U18573 (N_18573,N_11263,N_9596);
and U18574 (N_18574,N_7741,N_7298);
nand U18575 (N_18575,N_7417,N_9705);
or U18576 (N_18576,N_10061,N_11432);
and U18577 (N_18577,N_10431,N_9222);
nor U18578 (N_18578,N_6482,N_7958);
nand U18579 (N_18579,N_10862,N_7401);
nand U18580 (N_18580,N_9315,N_10056);
nor U18581 (N_18581,N_11374,N_11025);
and U18582 (N_18582,N_7105,N_9176);
xor U18583 (N_18583,N_8504,N_8303);
and U18584 (N_18584,N_8341,N_7544);
and U18585 (N_18585,N_8831,N_7330);
nand U18586 (N_18586,N_9848,N_8218);
nor U18587 (N_18587,N_12030,N_7810);
nor U18588 (N_18588,N_9028,N_7528);
nor U18589 (N_18589,N_9161,N_9219);
xor U18590 (N_18590,N_11307,N_6718);
nor U18591 (N_18591,N_11272,N_9105);
nand U18592 (N_18592,N_11077,N_9051);
xor U18593 (N_18593,N_10673,N_11614);
or U18594 (N_18594,N_12213,N_11762);
xnor U18595 (N_18595,N_9116,N_12389);
nand U18596 (N_18596,N_6600,N_11688);
nand U18597 (N_18597,N_11053,N_8655);
or U18598 (N_18598,N_11436,N_9975);
and U18599 (N_18599,N_6301,N_6627);
nand U18600 (N_18600,N_11070,N_6340);
xnor U18601 (N_18601,N_8948,N_7098);
nor U18602 (N_18602,N_11568,N_8383);
or U18603 (N_18603,N_10871,N_9619);
nand U18604 (N_18604,N_7570,N_11816);
xor U18605 (N_18605,N_8144,N_11168);
xor U18606 (N_18606,N_7897,N_7109);
or U18607 (N_18607,N_9998,N_12321);
or U18608 (N_18608,N_9074,N_11098);
xor U18609 (N_18609,N_11173,N_11306);
nor U18610 (N_18610,N_10620,N_7036);
xor U18611 (N_18611,N_10945,N_8105);
and U18612 (N_18612,N_8902,N_10835);
or U18613 (N_18613,N_6839,N_10222);
and U18614 (N_18614,N_7042,N_9765);
xnor U18615 (N_18615,N_7088,N_9844);
nor U18616 (N_18616,N_10663,N_12442);
xnor U18617 (N_18617,N_10782,N_11113);
and U18618 (N_18618,N_6901,N_6479);
xor U18619 (N_18619,N_11636,N_6704);
and U18620 (N_18620,N_8756,N_8710);
xor U18621 (N_18621,N_11442,N_8674);
nand U18622 (N_18622,N_7189,N_10467);
and U18623 (N_18623,N_7883,N_6777);
or U18624 (N_18624,N_11902,N_8049);
nand U18625 (N_18625,N_6306,N_7435);
nor U18626 (N_18626,N_11987,N_10269);
and U18627 (N_18627,N_6377,N_11467);
xnor U18628 (N_18628,N_11757,N_10013);
nand U18629 (N_18629,N_8319,N_11384);
nor U18630 (N_18630,N_11200,N_6618);
or U18631 (N_18631,N_10220,N_11448);
xnor U18632 (N_18632,N_12071,N_10206);
and U18633 (N_18633,N_8942,N_8078);
or U18634 (N_18634,N_9979,N_11132);
nand U18635 (N_18635,N_12171,N_11545);
xor U18636 (N_18636,N_10144,N_9741);
nor U18637 (N_18637,N_8031,N_11063);
and U18638 (N_18638,N_10615,N_11676);
and U18639 (N_18639,N_12059,N_10708);
or U18640 (N_18640,N_6684,N_11149);
and U18641 (N_18641,N_11927,N_10750);
and U18642 (N_18642,N_6836,N_7393);
xor U18643 (N_18643,N_7603,N_6919);
xnor U18644 (N_18644,N_9261,N_8196);
nand U18645 (N_18645,N_9807,N_12342);
xnor U18646 (N_18646,N_12148,N_9917);
xor U18647 (N_18647,N_9792,N_7652);
xnor U18648 (N_18648,N_7100,N_9954);
nand U18649 (N_18649,N_6365,N_12473);
or U18650 (N_18650,N_10760,N_6816);
nand U18651 (N_18651,N_11851,N_11004);
nand U18652 (N_18652,N_8517,N_9780);
nand U18653 (N_18653,N_10053,N_9621);
nand U18654 (N_18654,N_10732,N_10154);
nand U18655 (N_18655,N_11264,N_12314);
nor U18656 (N_18656,N_12370,N_10930);
or U18657 (N_18657,N_7699,N_10163);
and U18658 (N_18658,N_9678,N_7818);
nor U18659 (N_18659,N_9887,N_7828);
nor U18660 (N_18660,N_10115,N_11561);
or U18661 (N_18661,N_7741,N_11641);
or U18662 (N_18662,N_9453,N_6695);
or U18663 (N_18663,N_12130,N_8378);
xnor U18664 (N_18664,N_11786,N_6995);
nand U18665 (N_18665,N_10283,N_12445);
or U18666 (N_18666,N_11940,N_6574);
xor U18667 (N_18667,N_9172,N_10359);
or U18668 (N_18668,N_9121,N_10790);
or U18669 (N_18669,N_11029,N_6420);
xor U18670 (N_18670,N_9967,N_9617);
xor U18671 (N_18671,N_7818,N_9738);
nand U18672 (N_18672,N_9595,N_6345);
nand U18673 (N_18673,N_7410,N_10596);
nor U18674 (N_18674,N_11714,N_8957);
or U18675 (N_18675,N_10596,N_10061);
nand U18676 (N_18676,N_6624,N_9632);
nor U18677 (N_18677,N_8152,N_11234);
nor U18678 (N_18678,N_6824,N_11706);
and U18679 (N_18679,N_8526,N_11599);
and U18680 (N_18680,N_10226,N_11730);
or U18681 (N_18681,N_10548,N_12419);
or U18682 (N_18682,N_12341,N_8683);
and U18683 (N_18683,N_11419,N_9952);
xnor U18684 (N_18684,N_11985,N_10972);
and U18685 (N_18685,N_6794,N_7598);
or U18686 (N_18686,N_11767,N_8004);
nor U18687 (N_18687,N_10242,N_10812);
xnor U18688 (N_18688,N_7073,N_12436);
nor U18689 (N_18689,N_9560,N_10108);
xnor U18690 (N_18690,N_9163,N_7523);
or U18691 (N_18691,N_7344,N_7252);
xnor U18692 (N_18692,N_9953,N_7706);
nor U18693 (N_18693,N_6867,N_10038);
xor U18694 (N_18694,N_11812,N_12033);
and U18695 (N_18695,N_6932,N_11229);
or U18696 (N_18696,N_8167,N_9597);
or U18697 (N_18697,N_10714,N_8581);
nand U18698 (N_18698,N_9694,N_10553);
nand U18699 (N_18699,N_10259,N_10555);
or U18700 (N_18700,N_6708,N_8117);
or U18701 (N_18701,N_6982,N_10795);
and U18702 (N_18702,N_9888,N_10736);
nand U18703 (N_18703,N_8875,N_7387);
and U18704 (N_18704,N_11621,N_12115);
xnor U18705 (N_18705,N_11119,N_6403);
nand U18706 (N_18706,N_7834,N_9619);
nor U18707 (N_18707,N_9023,N_8513);
or U18708 (N_18708,N_11366,N_12158);
nand U18709 (N_18709,N_11294,N_10696);
nand U18710 (N_18710,N_10094,N_10150);
and U18711 (N_18711,N_8160,N_8255);
and U18712 (N_18712,N_7500,N_8117);
xor U18713 (N_18713,N_9024,N_6864);
nor U18714 (N_18714,N_11216,N_7773);
nand U18715 (N_18715,N_11177,N_7768);
or U18716 (N_18716,N_8879,N_9262);
nand U18717 (N_18717,N_6787,N_12336);
or U18718 (N_18718,N_11404,N_8942);
xnor U18719 (N_18719,N_11677,N_12262);
or U18720 (N_18720,N_7478,N_9676);
or U18721 (N_18721,N_12185,N_11445);
xor U18722 (N_18722,N_7910,N_10656);
xnor U18723 (N_18723,N_8590,N_10739);
nor U18724 (N_18724,N_7159,N_9112);
nor U18725 (N_18725,N_11538,N_9387);
and U18726 (N_18726,N_6770,N_9438);
nor U18727 (N_18727,N_10296,N_10749);
xnor U18728 (N_18728,N_8511,N_11928);
or U18729 (N_18729,N_8844,N_7406);
xor U18730 (N_18730,N_9710,N_7646);
nor U18731 (N_18731,N_9143,N_6573);
nor U18732 (N_18732,N_9782,N_6974);
and U18733 (N_18733,N_11084,N_8689);
xor U18734 (N_18734,N_8218,N_8187);
nor U18735 (N_18735,N_10992,N_9772);
and U18736 (N_18736,N_7237,N_12111);
or U18737 (N_18737,N_8582,N_8713);
and U18738 (N_18738,N_9630,N_12184);
nand U18739 (N_18739,N_11564,N_6342);
and U18740 (N_18740,N_8903,N_9392);
nand U18741 (N_18741,N_8778,N_8769);
nor U18742 (N_18742,N_7596,N_11616);
or U18743 (N_18743,N_12478,N_11001);
nand U18744 (N_18744,N_7877,N_7723);
and U18745 (N_18745,N_10031,N_7621);
and U18746 (N_18746,N_12317,N_11627);
nand U18747 (N_18747,N_10839,N_10210);
nor U18748 (N_18748,N_11976,N_11575);
nor U18749 (N_18749,N_12313,N_7140);
nor U18750 (N_18750,N_17558,N_14226);
and U18751 (N_18751,N_16306,N_12987);
or U18752 (N_18752,N_18068,N_16827);
and U18753 (N_18753,N_12975,N_18200);
nand U18754 (N_18754,N_14658,N_16889);
nor U18755 (N_18755,N_13590,N_12566);
nor U18756 (N_18756,N_16986,N_13428);
or U18757 (N_18757,N_12595,N_14865);
or U18758 (N_18758,N_17231,N_15175);
and U18759 (N_18759,N_16681,N_15490);
nand U18760 (N_18760,N_17130,N_18640);
and U18761 (N_18761,N_17957,N_13154);
and U18762 (N_18762,N_15792,N_17490);
nand U18763 (N_18763,N_16143,N_17912);
nor U18764 (N_18764,N_15363,N_15550);
nor U18765 (N_18765,N_15627,N_12531);
nor U18766 (N_18766,N_17870,N_15110);
and U18767 (N_18767,N_13491,N_18426);
nand U18768 (N_18768,N_12839,N_17062);
or U18769 (N_18769,N_16828,N_17250);
nand U18770 (N_18770,N_17152,N_15973);
nand U18771 (N_18771,N_13955,N_13555);
and U18772 (N_18772,N_13144,N_16377);
nor U18773 (N_18773,N_16231,N_17642);
xor U18774 (N_18774,N_17183,N_13357);
or U18775 (N_18775,N_14590,N_16529);
xor U18776 (N_18776,N_15016,N_17486);
and U18777 (N_18777,N_16560,N_13438);
xor U18778 (N_18778,N_13224,N_15401);
and U18779 (N_18779,N_13306,N_13320);
nand U18780 (N_18780,N_17001,N_12548);
xor U18781 (N_18781,N_18501,N_17655);
or U18782 (N_18782,N_14855,N_13009);
nand U18783 (N_18783,N_18514,N_17314);
nand U18784 (N_18784,N_17125,N_13313);
and U18785 (N_18785,N_14260,N_18669);
nor U18786 (N_18786,N_17953,N_16267);
nand U18787 (N_18787,N_13189,N_13010);
nand U18788 (N_18788,N_14376,N_15036);
xor U18789 (N_18789,N_13708,N_17790);
xor U18790 (N_18790,N_13921,N_18741);
xor U18791 (N_18791,N_18295,N_13731);
and U18792 (N_18792,N_18745,N_15287);
and U18793 (N_18793,N_12673,N_14467);
and U18794 (N_18794,N_14718,N_14979);
and U18795 (N_18795,N_12596,N_15727);
xnor U18796 (N_18796,N_16477,N_17452);
and U18797 (N_18797,N_14712,N_17975);
and U18798 (N_18798,N_18471,N_15601);
nand U18799 (N_18799,N_12961,N_16795);
nand U18800 (N_18800,N_14672,N_13474);
nand U18801 (N_18801,N_16951,N_12901);
nor U18802 (N_18802,N_13255,N_17536);
or U18803 (N_18803,N_15289,N_13656);
and U18804 (N_18804,N_14724,N_16884);
and U18805 (N_18805,N_16848,N_12789);
or U18806 (N_18806,N_15201,N_13429);
and U18807 (N_18807,N_14551,N_16208);
xor U18808 (N_18808,N_12685,N_18266);
or U18809 (N_18809,N_18289,N_15311);
nand U18810 (N_18810,N_17833,N_16935);
nand U18811 (N_18811,N_13246,N_15904);
nor U18812 (N_18812,N_17078,N_14659);
nor U18813 (N_18813,N_17432,N_18198);
and U18814 (N_18814,N_15648,N_17520);
or U18815 (N_18815,N_18711,N_18575);
and U18816 (N_18816,N_16695,N_15246);
nand U18817 (N_18817,N_14219,N_16983);
or U18818 (N_18818,N_12679,N_15147);
xor U18819 (N_18819,N_18151,N_16329);
nand U18820 (N_18820,N_16045,N_13751);
xnor U18821 (N_18821,N_13460,N_15894);
nand U18822 (N_18822,N_14611,N_16134);
or U18823 (N_18823,N_17441,N_14612);
nor U18824 (N_18824,N_18152,N_16342);
nand U18825 (N_18825,N_17017,N_16437);
nand U18826 (N_18826,N_17259,N_16422);
or U18827 (N_18827,N_17748,N_15074);
and U18828 (N_18828,N_15661,N_18002);
nor U18829 (N_18829,N_16398,N_17681);
xnor U18830 (N_18830,N_18272,N_18732);
nor U18831 (N_18831,N_12842,N_15086);
and U18832 (N_18832,N_16977,N_14577);
nand U18833 (N_18833,N_16486,N_12833);
nand U18834 (N_18834,N_15134,N_12787);
nand U18835 (N_18835,N_15681,N_13942);
nand U18836 (N_18836,N_18400,N_13545);
and U18837 (N_18837,N_13185,N_17906);
or U18838 (N_18838,N_13220,N_15475);
xor U18839 (N_18839,N_17493,N_15859);
and U18840 (N_18840,N_12616,N_14939);
and U18841 (N_18841,N_18603,N_13549);
and U18842 (N_18842,N_15438,N_13200);
and U18843 (N_18843,N_18605,N_13177);
nor U18844 (N_18844,N_16663,N_18218);
and U18845 (N_18845,N_17847,N_14727);
and U18846 (N_18846,N_16467,N_14579);
xnor U18847 (N_18847,N_13591,N_17856);
or U18848 (N_18848,N_15983,N_13886);
nand U18849 (N_18849,N_16016,N_13569);
or U18850 (N_18850,N_16771,N_18608);
nor U18851 (N_18851,N_16315,N_15162);
nand U18852 (N_18852,N_17397,N_16172);
xnor U18853 (N_18853,N_17469,N_18389);
xor U18854 (N_18854,N_17508,N_18247);
and U18855 (N_18855,N_14852,N_13210);
nand U18856 (N_18856,N_14300,N_14937);
nor U18857 (N_18857,N_18609,N_18549);
or U18858 (N_18858,N_13365,N_13114);
nand U18859 (N_18859,N_14386,N_14571);
xnor U18860 (N_18860,N_18148,N_18197);
nand U18861 (N_18861,N_14860,N_16714);
and U18862 (N_18862,N_15804,N_14918);
nor U18863 (N_18863,N_15950,N_15053);
xnor U18864 (N_18864,N_17290,N_15213);
and U18865 (N_18865,N_15451,N_16968);
xnor U18866 (N_18866,N_17304,N_17589);
or U18867 (N_18867,N_16969,N_17818);
nor U18868 (N_18868,N_15666,N_13923);
and U18869 (N_18869,N_15420,N_16772);
or U18870 (N_18870,N_14794,N_15834);
and U18871 (N_18871,N_18487,N_12910);
nor U18872 (N_18872,N_17881,N_12504);
or U18873 (N_18873,N_15729,N_16945);
and U18874 (N_18874,N_12551,N_13831);
and U18875 (N_18875,N_15798,N_15486);
or U18876 (N_18876,N_18070,N_14771);
nand U18877 (N_18877,N_17134,N_12998);
xnor U18878 (N_18878,N_17208,N_15252);
nor U18879 (N_18879,N_14265,N_12657);
nor U18880 (N_18880,N_17179,N_13269);
and U18881 (N_18881,N_18593,N_14209);
xnor U18882 (N_18882,N_16193,N_17745);
nor U18883 (N_18883,N_15535,N_18730);
and U18884 (N_18884,N_15527,N_13499);
and U18885 (N_18885,N_16929,N_18582);
or U18886 (N_18886,N_14597,N_18693);
nor U18887 (N_18887,N_17170,N_13825);
or U18888 (N_18888,N_13485,N_16523);
nor U18889 (N_18889,N_14801,N_17994);
nand U18890 (N_18890,N_14299,N_15421);
nand U18891 (N_18891,N_16404,N_18089);
xor U18892 (N_18892,N_14482,N_13716);
or U18893 (N_18893,N_17090,N_14772);
nor U18894 (N_18894,N_15699,N_14240);
nor U18895 (N_18895,N_13363,N_15072);
nand U18896 (N_18896,N_16475,N_17444);
and U18897 (N_18897,N_13713,N_16985);
or U18898 (N_18898,N_16163,N_15967);
nor U18899 (N_18899,N_12852,N_17067);
nor U18900 (N_18900,N_15127,N_14923);
nand U18901 (N_18901,N_17116,N_17186);
xor U18902 (N_18902,N_14746,N_13128);
nor U18903 (N_18903,N_15788,N_16954);
or U18904 (N_18904,N_13015,N_18257);
xor U18905 (N_18905,N_17879,N_13355);
or U18906 (N_18906,N_18393,N_16413);
or U18907 (N_18907,N_14459,N_17162);
nor U18908 (N_18908,N_16156,N_14307);
and U18909 (N_18909,N_15519,N_16494);
or U18910 (N_18910,N_14877,N_15885);
xnor U18911 (N_18911,N_15651,N_18668);
nor U18912 (N_18912,N_17047,N_12986);
xnor U18913 (N_18913,N_18182,N_17239);
xor U18914 (N_18914,N_14804,N_17466);
nor U18915 (N_18915,N_15168,N_17316);
nor U18916 (N_18916,N_13655,N_15516);
or U18917 (N_18917,N_13290,N_14043);
or U18918 (N_18918,N_15653,N_14983);
and U18919 (N_18919,N_17206,N_14706);
nand U18920 (N_18920,N_12742,N_14441);
nor U18921 (N_18921,N_16325,N_16819);
or U18922 (N_18922,N_15657,N_14038);
or U18923 (N_18923,N_16743,N_14595);
or U18924 (N_18924,N_14763,N_15954);
nand U18925 (N_18925,N_13771,N_15910);
and U18926 (N_18926,N_16744,N_17301);
nand U18927 (N_18927,N_18294,N_13403);
nand U18928 (N_18928,N_14092,N_13020);
nand U18929 (N_18929,N_18607,N_18240);
or U18930 (N_18930,N_13594,N_18168);
xor U18931 (N_18931,N_16387,N_15120);
nand U18932 (N_18932,N_15492,N_17942);
and U18933 (N_18933,N_15732,N_17031);
xor U18934 (N_18934,N_15735,N_14780);
nand U18935 (N_18935,N_12555,N_12632);
nor U18936 (N_18936,N_17335,N_15538);
xor U18937 (N_18937,N_13524,N_15595);
or U18938 (N_18938,N_15158,N_18001);
xnor U18939 (N_18939,N_13453,N_15341);
nand U18940 (N_18940,N_13073,N_16755);
xnor U18941 (N_18941,N_14208,N_16470);
and U18942 (N_18942,N_12713,N_12812);
or U18943 (N_18943,N_13121,N_15887);
nand U18944 (N_18944,N_17665,N_13547);
nand U18945 (N_18945,N_17085,N_15019);
or U18946 (N_18946,N_13407,N_17641);
and U18947 (N_18947,N_13568,N_16502);
nand U18948 (N_18948,N_17049,N_16824);
and U18949 (N_18949,N_15044,N_17232);
nor U18950 (N_18950,N_17042,N_13452);
xor U18951 (N_18951,N_17312,N_16854);
nand U18952 (N_18952,N_16294,N_13054);
nand U18953 (N_18953,N_12874,N_14816);
and U18954 (N_18954,N_12774,N_15095);
nor U18955 (N_18955,N_14641,N_16460);
or U18956 (N_18956,N_13959,N_15769);
nor U18957 (N_18957,N_18192,N_13593);
nor U18958 (N_18958,N_14497,N_15922);
xor U18959 (N_18959,N_16682,N_18298);
and U18960 (N_18960,N_15596,N_15011);
nand U18961 (N_18961,N_16576,N_14256);
and U18962 (N_18962,N_17238,N_13141);
nand U18963 (N_18963,N_14848,N_13150);
nand U18964 (N_18964,N_16149,N_13425);
nor U18965 (N_18965,N_17997,N_12667);
xnor U18966 (N_18966,N_17524,N_17340);
and U18967 (N_18967,N_12997,N_15961);
nor U18968 (N_18968,N_15046,N_12953);
and U18969 (N_18969,N_17715,N_18436);
and U18970 (N_18970,N_13149,N_13634);
xnor U18971 (N_18971,N_13245,N_15335);
or U18972 (N_18972,N_14451,N_12898);
nand U18973 (N_18973,N_15917,N_16555);
nor U18974 (N_18974,N_14834,N_14084);
and U18975 (N_18975,N_17960,N_13342);
and U18976 (N_18976,N_14969,N_12593);
xnor U18977 (N_18977,N_15774,N_14129);
nand U18978 (N_18978,N_17652,N_17150);
or U18979 (N_18979,N_14608,N_13080);
or U18980 (N_18980,N_17408,N_16836);
nand U18981 (N_18981,N_14170,N_16433);
xnor U18982 (N_18982,N_15427,N_14536);
xnor U18983 (N_18983,N_13686,N_18321);
nor U18984 (N_18984,N_12829,N_16664);
nor U18985 (N_18985,N_13789,N_15224);
and U18986 (N_18986,N_17288,N_14044);
or U18987 (N_18987,N_14588,N_14316);
or U18988 (N_18988,N_18425,N_15070);
or U18989 (N_18989,N_12920,N_18191);
nand U18990 (N_18990,N_17630,N_17889);
and U18991 (N_18991,N_14963,N_16481);
nor U18992 (N_18992,N_14311,N_16952);
xnor U18993 (N_18993,N_15106,N_14133);
or U18994 (N_18994,N_18021,N_13592);
nor U18995 (N_18995,N_13102,N_12984);
xor U18996 (N_18996,N_17549,N_18111);
or U18997 (N_18997,N_12582,N_14753);
and U18998 (N_18998,N_16288,N_17999);
or U18999 (N_18999,N_16811,N_18147);
xor U19000 (N_19000,N_14700,N_13448);
or U19001 (N_19001,N_15027,N_18153);
and U19002 (N_19002,N_12883,N_18035);
or U19003 (N_19003,N_16943,N_13117);
xnor U19004 (N_19004,N_13755,N_16212);
nor U19005 (N_19005,N_13865,N_16409);
xnor U19006 (N_19006,N_12958,N_16173);
and U19007 (N_19007,N_14964,N_15015);
or U19008 (N_19008,N_18359,N_14840);
and U19009 (N_19009,N_15431,N_14738);
xnor U19010 (N_19010,N_17801,N_17683);
xnor U19011 (N_19011,N_15534,N_14532);
or U19012 (N_19012,N_14762,N_15157);
xnor U19013 (N_19013,N_13626,N_17192);
nor U19014 (N_19014,N_14480,N_18217);
nand U19015 (N_19015,N_13377,N_17352);
and U19016 (N_19016,N_18597,N_13527);
or U19017 (N_19017,N_13884,N_14466);
nand U19018 (N_19018,N_13120,N_15563);
nor U19019 (N_19019,N_17088,N_16967);
and U19020 (N_19020,N_13092,N_18476);
nand U19021 (N_19021,N_18051,N_17199);
and U19022 (N_19022,N_13465,N_12957);
or U19023 (N_19023,N_18233,N_17657);
nand U19024 (N_19024,N_14907,N_13875);
and U19025 (N_19025,N_16721,N_15496);
nand U19026 (N_19026,N_17653,N_15925);
nand U19027 (N_19027,N_14910,N_14268);
and U19028 (N_19028,N_13617,N_17229);
xor U19029 (N_19029,N_17754,N_15066);
nor U19030 (N_19030,N_14392,N_17809);
xnor U19031 (N_19031,N_15059,N_14616);
or U19032 (N_19032,N_12722,N_12635);
xnor U19033 (N_19033,N_17362,N_14057);
or U19034 (N_19034,N_18533,N_16947);
xor U19035 (N_19035,N_18167,N_13833);
and U19036 (N_19036,N_18695,N_18063);
xor U19037 (N_19037,N_15476,N_16674);
and U19038 (N_19038,N_12978,N_12610);
nand U19039 (N_19039,N_15980,N_14107);
and U19040 (N_19040,N_12516,N_16202);
or U19041 (N_19041,N_15819,N_16634);
nand U19042 (N_19042,N_15674,N_13791);
nor U19043 (N_19043,N_16505,N_17048);
or U19044 (N_19044,N_13935,N_17323);
and U19045 (N_19045,N_12581,N_15458);
and U19046 (N_19046,N_13866,N_18709);
nand U19047 (N_19047,N_18241,N_15277);
xor U19048 (N_19048,N_13059,N_13885);
nor U19049 (N_19049,N_18412,N_15814);
and U19050 (N_19050,N_12557,N_16292);
xor U19051 (N_19051,N_14011,N_15189);
nand U19052 (N_19052,N_16590,N_13649);
nor U19053 (N_19053,N_17979,N_14207);
xor U19054 (N_19054,N_17507,N_14808);
nor U19055 (N_19055,N_13086,N_14003);
nor U19056 (N_19056,N_16885,N_15270);
nand U19057 (N_19057,N_15465,N_15726);
or U19058 (N_19058,N_15564,N_13180);
and U19059 (N_19059,N_17566,N_18009);
xor U19060 (N_19060,N_13480,N_15809);
xnor U19061 (N_19061,N_14345,N_14610);
nor U19062 (N_19062,N_12682,N_14061);
nand U19063 (N_19063,N_12553,N_16356);
xor U19064 (N_19064,N_18660,N_12908);
xor U19065 (N_19065,N_18539,N_16620);
and U19066 (N_19066,N_14190,N_13603);
xor U19067 (N_19067,N_15480,N_13648);
nand U19068 (N_19068,N_14193,N_14246);
nand U19069 (N_19069,N_16726,N_16676);
or U19070 (N_19070,N_12932,N_13945);
nand U19071 (N_19071,N_17504,N_12868);
or U19072 (N_19072,N_15028,N_17546);
nand U19073 (N_19073,N_12505,N_17036);
xor U19074 (N_19074,N_16476,N_15235);
and U19075 (N_19075,N_14534,N_14460);
xnor U19076 (N_19076,N_14598,N_16660);
nor U19077 (N_19077,N_16363,N_18285);
xnor U19078 (N_19078,N_16277,N_12625);
nand U19079 (N_19079,N_16264,N_15455);
xnor U19080 (N_19080,N_14785,N_17509);
nor U19081 (N_19081,N_14118,N_13960);
xnor U19082 (N_19082,N_14552,N_14817);
nand U19083 (N_19083,N_13842,N_14350);
or U19084 (N_19084,N_18427,N_14777);
nand U19085 (N_19085,N_13608,N_15688);
nand U19086 (N_19086,N_15787,N_17387);
nand U19087 (N_19087,N_17599,N_15380);
or U19088 (N_19088,N_14956,N_16395);
nand U19089 (N_19089,N_15082,N_12659);
xor U19090 (N_19090,N_14032,N_17988);
nand U19091 (N_19091,N_15881,N_13249);
and U19092 (N_19092,N_14862,N_16993);
nor U19093 (N_19093,N_14132,N_14618);
nor U19094 (N_19094,N_17253,N_13676);
xnor U19095 (N_19095,N_13042,N_13829);
xnor U19096 (N_19096,N_18394,N_16093);
nor U19097 (N_19097,N_14033,N_13427);
nand U19098 (N_19098,N_12799,N_14285);
nor U19099 (N_19099,N_13937,N_16822);
xor U19100 (N_19100,N_15355,N_13466);
nand U19101 (N_19101,N_14085,N_16987);
and U19102 (N_19102,N_12913,N_16251);
nor U19103 (N_19103,N_14624,N_17069);
or U19104 (N_19104,N_18517,N_14934);
nor U19105 (N_19105,N_15903,N_13419);
nand U19106 (N_19106,N_16246,N_15460);
or U19107 (N_19107,N_14416,N_17635);
nor U19108 (N_19108,N_14449,N_15195);
nor U19109 (N_19109,N_13788,N_17396);
nand U19110 (N_19110,N_12822,N_13761);
or U19111 (N_19111,N_17808,N_14131);
nor U19112 (N_19112,N_13878,N_18073);
and U19113 (N_19113,N_14121,N_14112);
nand U19114 (N_19114,N_13490,N_17488);
nor U19115 (N_19115,N_14888,N_14580);
and U19116 (N_19116,N_17629,N_15518);
nand U19117 (N_19117,N_16767,N_16168);
nor U19118 (N_19118,N_17919,N_15071);
nand U19119 (N_19119,N_18408,N_14568);
nor U19120 (N_19120,N_13239,N_16556);
nor U19121 (N_19121,N_13038,N_16488);
nor U19122 (N_19122,N_16571,N_13680);
and U19123 (N_19123,N_14348,N_16863);
nor U19124 (N_19124,N_15414,N_13505);
xnor U19125 (N_19125,N_13288,N_12994);
nand U19126 (N_19126,N_14798,N_14250);
nor U19127 (N_19127,N_12550,N_12993);
nor U19128 (N_19128,N_16281,N_16964);
or U19129 (N_19129,N_18339,N_16650);
nand U19130 (N_19130,N_14912,N_17177);
or U19131 (N_19131,N_17105,N_13197);
xor U19132 (N_19132,N_16920,N_18061);
or U19133 (N_19133,N_13016,N_15907);
xor U19134 (N_19134,N_14468,N_18529);
or U19135 (N_19135,N_13785,N_13230);
nor U19136 (N_19136,N_14339,N_12525);
nor U19137 (N_19137,N_17103,N_13675);
and U19138 (N_19138,N_14055,N_14884);
or U19139 (N_19139,N_16835,N_16763);
or U19140 (N_19140,N_13665,N_17738);
xor U19141 (N_19141,N_15358,N_17060);
and U19142 (N_19142,N_16328,N_15330);
nand U19143 (N_19143,N_16895,N_13175);
nand U19144 (N_19144,N_17435,N_13550);
xor U19145 (N_19145,N_14503,N_14947);
and U19146 (N_19146,N_13219,N_16937);
or U19147 (N_19147,N_18567,N_14864);
nor U19148 (N_19148,N_14555,N_18645);
nor U19149 (N_19149,N_15343,N_13976);
nor U19150 (N_19150,N_16057,N_17694);
nor U19151 (N_19151,N_13947,N_16610);
and U19152 (N_19152,N_17223,N_15411);
and U19153 (N_19153,N_15276,N_14788);
xor U19154 (N_19154,N_15823,N_14470);
nor U19155 (N_19155,N_15462,N_16719);
xnor U19156 (N_19156,N_18520,N_16852);
nand U19157 (N_19157,N_14446,N_16867);
and U19158 (N_19158,N_16207,N_15700);
or U19159 (N_19159,N_14187,N_13027);
and U19160 (N_19160,N_16781,N_18411);
and U19161 (N_19161,N_14009,N_15269);
and U19162 (N_19162,N_16940,N_15280);
nand U19163 (N_19163,N_16754,N_16578);
xnor U19164 (N_19164,N_16091,N_17485);
nor U19165 (N_19165,N_12518,N_17235);
nand U19166 (N_19166,N_16715,N_16785);
xor U19167 (N_19167,N_13880,N_17914);
nor U19168 (N_19168,N_15064,N_14664);
or U19169 (N_19169,N_18523,N_12549);
nor U19170 (N_19170,N_17968,N_16381);
or U19171 (N_19171,N_16160,N_14324);
nor U19172 (N_19172,N_14232,N_16462);
nand U19173 (N_19173,N_18156,N_16542);
xor U19174 (N_19174,N_17632,N_16751);
or U19175 (N_19175,N_13134,N_14485);
nand U19176 (N_19176,N_13874,N_18004);
or U19177 (N_19177,N_18223,N_14745);
nor U19178 (N_19178,N_17849,N_18444);
or U19179 (N_19179,N_13889,N_16549);
nor U19180 (N_19180,N_13164,N_12554);
and U19181 (N_19181,N_15014,N_13234);
or U19182 (N_19182,N_12583,N_18185);
nand U19183 (N_19183,N_14262,N_12598);
xnor U19184 (N_19184,N_12627,N_14797);
or U19185 (N_19185,N_14191,N_18030);
nand U19186 (N_19186,N_15990,N_14053);
and U19187 (N_19187,N_18193,N_16056);
and U19188 (N_19188,N_18022,N_14781);
or U19189 (N_19189,N_18729,N_15763);
xnor U19190 (N_19190,N_18356,N_16118);
or U19191 (N_19191,N_15042,N_12574);
nor U19192 (N_19192,N_16028,N_16565);
xnor U19193 (N_19193,N_17735,N_16197);
nand U19194 (N_19194,N_13922,N_14439);
nand U19195 (N_19195,N_14231,N_13450);
nor U19196 (N_19196,N_14836,N_14136);
or U19197 (N_19197,N_14980,N_17770);
nand U19198 (N_19198,N_15687,N_14389);
nor U19199 (N_19199,N_15102,N_13966);
and U19200 (N_19200,N_14830,N_17249);
nor U19201 (N_19201,N_13050,N_13621);
nor U19202 (N_19202,N_17104,N_16535);
nand U19203 (N_19203,N_13734,N_16581);
xor U19204 (N_19204,N_13849,N_15302);
nand U19205 (N_19205,N_15299,N_15829);
xor U19206 (N_19206,N_15013,N_17024);
nor U19207 (N_19207,N_13746,N_13596);
xnor U19208 (N_19208,N_16067,N_16641);
nor U19209 (N_19209,N_14374,N_14946);
or U19210 (N_19210,N_17859,N_17443);
nor U19211 (N_19211,N_17560,N_18591);
xor U19212 (N_19212,N_16871,N_13254);
and U19213 (N_19213,N_13289,N_15223);
nor U19214 (N_19214,N_16095,N_15507);
nor U19215 (N_19215,N_17730,N_13541);
nor U19216 (N_19216,N_12615,N_17122);
and U19217 (N_19217,N_16766,N_13696);
nand U19218 (N_19218,N_17424,N_14182);
xor U19219 (N_19219,N_16793,N_14525);
nor U19220 (N_19220,N_17187,N_13691);
and U19221 (N_19221,N_17300,N_17938);
nor U19222 (N_19222,N_18428,N_14405);
and U19223 (N_19223,N_13599,N_16047);
nand U19224 (N_19224,N_17718,N_15061);
nor U19225 (N_19225,N_17554,N_15007);
nor U19226 (N_19226,N_18731,N_14362);
or U19227 (N_19227,N_14224,N_14357);
xor U19228 (N_19228,N_14896,N_18460);
nor U19229 (N_19229,N_18599,N_16575);
and U19230 (N_19230,N_16309,N_16319);
or U19231 (N_19231,N_15248,N_13604);
xnor U19232 (N_19232,N_13522,N_12796);
xnor U19233 (N_19233,N_17117,N_18540);
xnor U19234 (N_19234,N_16688,N_16675);
or U19235 (N_19235,N_13238,N_14795);
nand U19236 (N_19236,N_16868,N_14211);
nand U19237 (N_19237,N_17143,N_18250);
nor U19238 (N_19238,N_13406,N_14991);
and U19239 (N_19239,N_16471,N_13887);
and U19240 (N_19240,N_15261,N_12959);
or U19241 (N_19241,N_17065,N_13404);
nand U19242 (N_19242,N_12572,N_13692);
xor U19243 (N_19243,N_14770,N_18509);
or U19244 (N_19244,N_12541,N_14221);
nand U19245 (N_19245,N_15831,N_17713);
nand U19246 (N_19246,N_15911,N_15097);
or U19247 (N_19247,N_12513,N_14626);
nor U19248 (N_19248,N_16907,N_16587);
xnor U19249 (N_19249,N_17716,N_16652);
and U19250 (N_19250,N_16052,N_14444);
and U19251 (N_19251,N_13066,N_14068);
and U19252 (N_19252,N_13623,N_16770);
xnor U19253 (N_19253,N_16419,N_15893);
nor U19254 (N_19254,N_18438,N_14164);
or U19255 (N_19255,N_12732,N_15909);
or U19256 (N_19256,N_18449,N_16996);
and U19257 (N_19257,N_14022,N_14786);
or U19258 (N_19258,N_16392,N_15386);
nor U19259 (N_19259,N_14596,N_17992);
nand U19260 (N_19260,N_13546,N_13468);
or U19261 (N_19261,N_15669,N_16326);
nor U19262 (N_19262,N_13784,N_16321);
nand U19263 (N_19263,N_17415,N_16138);
xnor U19264 (N_19264,N_15430,N_13919);
or U19265 (N_19265,N_12892,N_12857);
and U19266 (N_19266,N_16830,N_15599);
xor U19267 (N_19267,N_13390,N_15432);
nand U19268 (N_19268,N_17580,N_16021);
and U19269 (N_19269,N_12559,N_12628);
xnor U19270 (N_19270,N_16158,N_14683);
or U19271 (N_19271,N_14401,N_13916);
nor U19272 (N_19272,N_18551,N_16802);
or U19273 (N_19273,N_18722,N_17752);
nor U19274 (N_19274,N_12600,N_16960);
xor U19275 (N_19275,N_18406,N_14733);
nor U19276 (N_19276,N_16085,N_14635);
nand U19277 (N_19277,N_18503,N_15410);
nand U19278 (N_19278,N_14719,N_12939);
xor U19279 (N_19279,N_14083,N_18634);
and U19280 (N_19280,N_13852,N_12836);
nor U19281 (N_19281,N_13236,N_14506);
xnor U19282 (N_19282,N_12545,N_17107);
nand U19283 (N_19283,N_14775,N_16457);
nor U19284 (N_19284,N_12500,N_13104);
and U19285 (N_19285,N_15413,N_17261);
and U19286 (N_19286,N_15360,N_18346);
and U19287 (N_19287,N_14399,N_17543);
and U19288 (N_19288,N_12652,N_14515);
or U19289 (N_19289,N_14023,N_17654);
or U19290 (N_19290,N_12784,N_15286);
and U19291 (N_19291,N_12613,N_14120);
nand U19292 (N_19292,N_14422,N_18433);
nand U19293 (N_19293,N_17310,N_16019);
and U19294 (N_19294,N_14500,N_14548);
nor U19295 (N_19295,N_16849,N_16786);
or U19296 (N_19296,N_13732,N_14874);
nand U19297 (N_19297,N_13996,N_17869);
and U19298 (N_19298,N_13241,N_17428);
or U19299 (N_19299,N_17234,N_18364);
xor U19300 (N_19300,N_16094,N_13683);
nor U19301 (N_19301,N_12696,N_15370);
or U19302 (N_19302,N_14294,N_18654);
or U19303 (N_19303,N_16635,N_18513);
xor U19304 (N_19304,N_15495,N_17133);
or U19305 (N_19305,N_13948,N_18666);
or U19306 (N_19306,N_18313,N_16366);
xor U19307 (N_19307,N_18748,N_16606);
and U19308 (N_19308,N_14212,N_13272);
nor U19309 (N_19309,N_14421,N_13684);
nand U19310 (N_19310,N_16098,N_16004);
or U19311 (N_19311,N_15778,N_17557);
or U19312 (N_19312,N_16667,N_18131);
xor U19313 (N_19313,N_15029,N_12644);
nand U19314 (N_19314,N_17567,N_16918);
or U19315 (N_19315,N_14743,N_18450);
and U19316 (N_19316,N_16099,N_14867);
nand U19317 (N_19317,N_16778,N_15205);
nand U19318 (N_19318,N_15452,N_17463);
or U19319 (N_19319,N_18532,N_15434);
xnor U19320 (N_19320,N_17623,N_17297);
and U19321 (N_19321,N_13385,N_12942);
or U19322 (N_19322,N_16374,N_17838);
xor U19323 (N_19323,N_13139,N_18093);
or U19324 (N_19324,N_14866,N_18173);
or U19325 (N_19325,N_17837,N_16685);
nand U19326 (N_19326,N_15618,N_15841);
nor U19327 (N_19327,N_17032,N_17902);
nand U19328 (N_19328,N_13291,N_15931);
xor U19329 (N_19329,N_18323,N_18472);
nor U19330 (N_19330,N_13443,N_14544);
nand U19331 (N_19331,N_16648,N_14842);
nand U19332 (N_19332,N_16307,N_15470);
or U19333 (N_19333,N_14483,N_13244);
xnor U19334 (N_19334,N_14931,N_15031);
and U19335 (N_19335,N_13790,N_18054);
xnor U19336 (N_19336,N_17305,N_15582);
xnor U19337 (N_19337,N_16613,N_16383);
nor U19338 (N_19338,N_16238,N_18362);
and U19339 (N_19339,N_18318,N_12717);
or U19340 (N_19340,N_15136,N_18287);
nand U19341 (N_19341,N_18160,N_14958);
nor U19342 (N_19342,N_13389,N_13388);
or U19343 (N_19343,N_17886,N_17939);
or U19344 (N_19344,N_15544,N_18424);
nor U19345 (N_19345,N_14042,N_13069);
or U19346 (N_19346,N_17658,N_18194);
nor U19347 (N_19347,N_13048,N_13077);
nand U19348 (N_19348,N_15997,N_12743);
and U19349 (N_19349,N_15958,N_14234);
nand U19350 (N_19350,N_17144,N_14223);
xnor U19351 (N_19351,N_15955,N_13259);
xnor U19352 (N_19352,N_18564,N_16566);
nand U19353 (N_19353,N_14437,N_14759);
nor U19354 (N_19354,N_17556,N_14378);
or U19355 (N_19355,N_13216,N_17040);
nor U19356 (N_19356,N_16239,N_15226);
or U19357 (N_19357,N_15691,N_16787);
or U19358 (N_19358,N_17846,N_17076);
and U19359 (N_19359,N_13497,N_13808);
or U19360 (N_19360,N_14204,N_13304);
xor U19361 (N_19361,N_14058,N_13266);
nand U19362 (N_19362,N_16268,N_15324);
nand U19363 (N_19363,N_16077,N_17220);
nand U19364 (N_19364,N_18170,N_15919);
nor U19365 (N_19365,N_16493,N_13830);
xor U19366 (N_19366,N_13125,N_17618);
nor U19367 (N_19367,N_13152,N_13479);
or U19368 (N_19368,N_17110,N_13917);
nor U19369 (N_19369,N_16516,N_15442);
nand U19370 (N_19370,N_12607,N_16064);
xor U19371 (N_19371,N_14589,N_13101);
or U19372 (N_19372,N_15832,N_16563);
and U19373 (N_19373,N_17878,N_16128);
nand U19374 (N_19374,N_14387,N_18349);
nor U19375 (N_19375,N_15636,N_13477);
or U19376 (N_19376,N_18596,N_17501);
and U19377 (N_19377,N_16847,N_15600);
nor U19378 (N_19378,N_17820,N_17733);
or U19379 (N_19379,N_13412,N_14424);
and U19380 (N_19380,N_15838,N_14513);
and U19381 (N_19381,N_17829,N_17781);
nor U19382 (N_19382,N_14197,N_15030);
xnor U19383 (N_19383,N_17273,N_16414);
or U19384 (N_19384,N_18270,N_15836);
xor U19385 (N_19385,N_18494,N_16725);
and U19386 (N_19386,N_14566,N_12899);
and U19387 (N_19387,N_15112,N_14553);
nor U19388 (N_19388,N_14791,N_14900);
nand U19389 (N_19389,N_15171,N_16804);
or U19390 (N_19390,N_18464,N_17964);
nor U19391 (N_19391,N_16009,N_17918);
and U19392 (N_19392,N_18039,N_13828);
and U19393 (N_19393,N_15159,N_13142);
xor U19394 (N_19394,N_15759,N_13381);
and U19395 (N_19395,N_13011,N_18475);
nor U19396 (N_19396,N_18391,N_15474);
or U19397 (N_19397,N_16970,N_16014);
nor U19398 (N_19398,N_12885,N_13183);
nor U19399 (N_19399,N_18327,N_16196);
or U19400 (N_19400,N_18655,N_13169);
xor U19401 (N_19401,N_14139,N_16266);
and U19402 (N_19402,N_12974,N_14457);
xor U19403 (N_19403,N_15234,N_13752);
nand U19404 (N_19404,N_17484,N_14127);
xnor U19405 (N_19405,N_15542,N_17926);
nand U19406 (N_19406,N_15617,N_18211);
xnor U19407 (N_19407,N_17602,N_17570);
nand U19408 (N_19408,N_14008,N_12648);
nand U19409 (N_19409,N_17245,N_14490);
or U19410 (N_19410,N_14545,N_16540);
nor U19411 (N_19411,N_17522,N_14429);
or U19412 (N_19412,N_14585,N_15867);
or U19413 (N_19413,N_13638,N_13287);
nand U19414 (N_19414,N_18442,N_17924);
and U19415 (N_19415,N_14657,N_12968);
nand U19416 (N_19416,N_16602,N_14259);
nor U19417 (N_19417,N_12925,N_14846);
or U19418 (N_19418,N_17499,N_17850);
and U19419 (N_19419,N_17483,N_13278);
nor U19420 (N_19420,N_17679,N_18018);
xnor U19421 (N_19421,N_14819,N_16988);
nor U19422 (N_19422,N_15923,N_13826);
nor U19423 (N_19423,N_13132,N_17639);
and U19424 (N_19424,N_18474,N_17603);
nor U19425 (N_19425,N_13578,N_16547);
or U19426 (N_19426,N_18245,N_17863);
nand U19427 (N_19427,N_15616,N_15154);
nand U19428 (N_19428,N_16761,N_16204);
xnor U19429 (N_19429,N_18341,N_16015);
xnor U19430 (N_19430,N_15847,N_15536);
or U19431 (N_19431,N_17098,N_17815);
and U19432 (N_19432,N_15350,N_16205);
or U19433 (N_19433,N_16005,N_14652);
xnor U19434 (N_19434,N_12864,N_14229);
nor U19435 (N_19435,N_13565,N_18548);
and U19436 (N_19436,N_17277,N_16466);
or U19437 (N_19437,N_17740,N_13756);
and U19438 (N_19438,N_12624,N_12886);
xor U19439 (N_19439,N_18186,N_12825);
nand U19440 (N_19440,N_17895,N_14415);
xnor U19441 (N_19441,N_18521,N_13981);
and U19442 (N_19442,N_12952,N_16459);
nor U19443 (N_19443,N_14688,N_14965);
or U19444 (N_19444,N_13079,N_18251);
nor U19445 (N_19445,N_14572,N_18606);
nor U19446 (N_19446,N_17996,N_13325);
or U19447 (N_19447,N_17000,N_17553);
and U19448 (N_19448,N_17534,N_14440);
nor U19449 (N_19449,N_14060,N_14052);
nand U19450 (N_19450,N_14478,N_18589);
or U19451 (N_19451,N_17315,N_15025);
xnor U19452 (N_19452,N_15231,N_18102);
xor U19453 (N_19453,N_13977,N_14674);
xnor U19454 (N_19454,N_17527,N_14847);
or U19455 (N_19455,N_16931,N_17080);
xor U19456 (N_19456,N_14407,N_17822);
or U19457 (N_19457,N_18468,N_15200);
or U19458 (N_19458,N_13943,N_13644);
xnor U19459 (N_19459,N_12621,N_17225);
nand U19460 (N_19460,N_14504,N_18264);
or U19461 (N_19461,N_13036,N_14064);
nand U19462 (N_19462,N_13435,N_16046);
xnor U19463 (N_19463,N_17695,N_16922);
xnor U19464 (N_19464,N_17542,N_16224);
or U19465 (N_19465,N_15143,N_15970);
or U19466 (N_19466,N_17579,N_17330);
nand U19467 (N_19467,N_17375,N_17064);
and U19468 (N_19468,N_14681,N_17548);
or U19469 (N_19469,N_17771,N_12967);
nand U19470 (N_19470,N_15827,N_12684);
xnor U19471 (N_19471,N_14687,N_15852);
or U19472 (N_19472,N_15630,N_13993);
nand U19473 (N_19473,N_13103,N_16712);
or U19474 (N_19474,N_14729,N_17329);
and U19475 (N_19475,N_17216,N_16886);
nand U19476 (N_19476,N_18271,N_13487);
nand U19477 (N_19477,N_14406,N_17736);
xor U19478 (N_19478,N_13766,N_18696);
xor U19479 (N_19479,N_13498,N_15292);
or U19480 (N_19480,N_14177,N_14741);
or U19481 (N_19481,N_18028,N_17897);
xnor U19482 (N_19482,N_14831,N_17724);
nand U19483 (N_19483,N_16534,N_13515);
xor U19484 (N_19484,N_18623,N_16011);
nor U19485 (N_19485,N_18048,N_17153);
xnor U19486 (N_19486,N_14021,N_18179);
nor U19487 (N_19487,N_17081,N_18635);
or U19488 (N_19488,N_17591,N_16962);
or U19489 (N_19489,N_15433,N_13773);
and U19490 (N_19490,N_14995,N_17697);
nor U19491 (N_19491,N_16088,N_14695);
xnor U19492 (N_19492,N_12938,N_17773);
and U19493 (N_19493,N_18541,N_12956);
xor U19494 (N_19494,N_16144,N_14269);
or U19495 (N_19495,N_14135,N_13076);
nor U19496 (N_19496,N_15121,N_14062);
xor U19497 (N_19497,N_17875,N_16519);
and U19498 (N_19498,N_13774,N_15103);
xnor U19499 (N_19499,N_17782,N_15230);
nor U19500 (N_19500,N_13040,N_14241);
or U19501 (N_19501,N_13736,N_16564);
xnor U19502 (N_19502,N_13606,N_14990);
nor U19503 (N_19503,N_14007,N_18561);
and U19504 (N_19504,N_16062,N_17664);
nor U19505 (N_19505,N_17289,N_15837);
nor U19506 (N_19506,N_16483,N_12654);
nor U19507 (N_19507,N_16798,N_18095);
or U19508 (N_19508,N_15384,N_14283);
and U19509 (N_19509,N_13516,N_13769);
and U19510 (N_19510,N_17243,N_14857);
nor U19511 (N_19511,N_13562,N_13240);
xnor U19512 (N_19512,N_13472,N_18601);
xor U19513 (N_19513,N_17927,N_15946);
nor U19514 (N_19514,N_15683,N_12636);
nor U19515 (N_19515,N_17359,N_14692);
xor U19516 (N_19516,N_12765,N_18662);
xnor U19517 (N_19517,N_17731,N_15253);
or U19518 (N_19518,N_17834,N_17616);
or U19519 (N_19519,N_12777,N_17840);
and U19520 (N_19520,N_16774,N_15367);
nand U19521 (N_19521,N_12676,N_18094);
or U19522 (N_19522,N_15797,N_15356);
nand U19523 (N_19523,N_14200,N_17255);
or U19524 (N_19524,N_16237,N_13494);
xnor U19525 (N_19525,N_16588,N_13386);
xnor U19526 (N_19526,N_14111,N_17188);
xor U19527 (N_19527,N_15587,N_16496);
nand U19528 (N_19528,N_18319,N_12605);
nand U19529 (N_19529,N_18714,N_17126);
and U19530 (N_19530,N_13525,N_18273);
nor U19531 (N_19531,N_15854,N_12837);
nor U19532 (N_19532,N_15746,N_15948);
nor U19533 (N_19533,N_13850,N_15344);
nor U19534 (N_19534,N_14333,N_15730);
and U19535 (N_19535,N_17203,N_18683);
nand U19536 (N_19536,N_13409,N_16706);
nand U19537 (N_19537,N_12589,N_17005);
or U19538 (N_19538,N_18091,N_16910);
or U19539 (N_19539,N_12951,N_12780);
nor U19540 (N_19540,N_14296,N_17739);
or U19541 (N_19541,N_15406,N_13612);
or U19542 (N_19542,N_18062,N_16112);
nand U19543 (N_19543,N_15672,N_12580);
and U19544 (N_19544,N_17796,N_16082);
nand U19545 (N_19545,N_17762,N_12775);
or U19546 (N_19546,N_17129,N_13558);
and U19547 (N_19547,N_17194,N_15679);
nor U19548 (N_19548,N_18719,N_16815);
xnor U19549 (N_19549,N_17202,N_13297);
and U19550 (N_19550,N_18171,N_17828);
xnor U19551 (N_19551,N_17169,N_16936);
or U19552 (N_19552,N_16119,N_17516);
nand U19553 (N_19553,N_13387,N_15076);
xnor U19554 (N_19554,N_14462,N_16882);
or U19555 (N_19555,N_16375,N_18299);
or U19556 (N_19556,N_16557,N_15454);
xnor U19557 (N_19557,N_18144,N_16553);
or U19558 (N_19558,N_16076,N_16407);
and U19559 (N_19559,N_14889,N_13379);
nand U19560 (N_19560,N_18157,N_18451);
nor U19561 (N_19561,N_13455,N_16216);
and U19562 (N_19562,N_14975,N_18263);
nand U19563 (N_19563,N_14036,N_13580);
nor U19564 (N_19564,N_14933,N_16691);
and U19565 (N_19565,N_13859,N_14461);
and U19566 (N_19566,N_17146,N_13999);
nand U19567 (N_19567,N_15924,N_13107);
nand U19568 (N_19568,N_12808,N_14163);
nand U19569 (N_19569,N_13195,N_18692);
and U19570 (N_19570,N_17181,N_14575);
nand U19571 (N_19571,N_12646,N_17720);
xor U19572 (N_19572,N_14172,N_17690);
or U19573 (N_19573,N_14400,N_14481);
nor U19574 (N_19574,N_15240,N_18497);
nand U19575 (N_19575,N_14748,N_14134);
nor U19576 (N_19576,N_15409,N_15212);
and U19577 (N_19577,N_13687,N_13834);
nand U19578 (N_19578,N_18130,N_17744);
or U19579 (N_19579,N_16153,N_12801);
nand U19580 (N_19580,N_13160,N_14465);
nand U19581 (N_19581,N_13292,N_18262);
and U19582 (N_19582,N_18316,N_18116);
nor U19583 (N_19583,N_13314,N_15926);
and U19584 (N_19584,N_13229,N_16203);
nand U19585 (N_19585,N_15187,N_12879);
nand U19586 (N_19586,N_13726,N_12965);
and U19587 (N_19587,N_12608,N_14445);
xor U19588 (N_19588,N_16278,N_13112);
or U19589 (N_19589,N_15712,N_18036);
xor U19590 (N_19590,N_18122,N_16741);
and U19591 (N_19591,N_16963,N_14761);
nand U19592 (N_19592,N_14565,N_12532);
or U19593 (N_19593,N_13349,N_17112);
or U19594 (N_19594,N_15347,N_17409);
nor U19595 (N_19595,N_18677,N_15100);
xor U19596 (N_19596,N_17271,N_17650);
xor U19597 (N_19597,N_16994,N_16360);
nor U19598 (N_19598,N_17788,N_18355);
and U19599 (N_19599,N_13492,N_18081);
or U19600 (N_19600,N_13820,N_13065);
nand U19601 (N_19601,N_13818,N_18379);
or U19602 (N_19602,N_17728,N_15346);
or U19603 (N_19603,N_13082,N_14395);
or U19604 (N_19604,N_16898,N_14144);
and U19605 (N_19605,N_13658,N_18003);
nor U19606 (N_19606,N_14332,N_16037);
xor U19607 (N_19607,N_18616,N_16784);
nand U19608 (N_19608,N_14284,N_15810);
nand U19609 (N_19609,N_16522,N_17418);
or U19610 (N_19610,N_17872,N_17743);
or U19611 (N_19611,N_17535,N_12735);
or U19612 (N_19612,N_14411,N_12662);
or U19613 (N_19613,N_15780,N_14100);
and U19614 (N_19614,N_16299,N_17331);
xor U19615 (N_19615,N_17185,N_15238);
xor U19616 (N_19616,N_17191,N_18701);
and U19617 (N_19617,N_13869,N_17322);
or U19618 (N_19618,N_12631,N_17096);
and U19619 (N_19619,N_16817,N_14199);
and U19620 (N_19620,N_16869,N_16858);
and U19621 (N_19621,N_18132,N_18614);
or U19622 (N_19622,N_18096,N_16717);
nor U19623 (N_19623,N_15142,N_12982);
nor U19624 (N_19624,N_13824,N_14206);
nand U19625 (N_19625,N_15003,N_16508);
and U19626 (N_19626,N_17114,N_13679);
or U19627 (N_19627,N_13360,N_13561);
nor U19628 (N_19628,N_12750,N_17686);
nor U19629 (N_19629,N_16218,N_14488);
nor U19630 (N_19630,N_13136,N_15993);
nor U19631 (N_19631,N_13051,N_13228);
and U19632 (N_19632,N_15428,N_15232);
xnor U19633 (N_19633,N_16035,N_17705);
and U19634 (N_19634,N_14323,N_13988);
nor U19635 (N_19635,N_15285,N_17166);
xor U19636 (N_19636,N_14986,N_14522);
and U19637 (N_19637,N_14020,N_15960);
xor U19638 (N_19638,N_18113,N_15621);
xnor U19639 (N_19639,N_16311,N_15441);
nor U19640 (N_19640,N_16102,N_16242);
nand U19641 (N_19641,N_17257,N_16832);
and U19642 (N_19642,N_18358,N_13252);
xnor U19643 (N_19643,N_17789,N_15489);
xnor U19644 (N_19644,N_13827,N_14870);
or U19645 (N_19645,N_17390,N_17931);
and U19646 (N_19646,N_12564,N_15004);
and U19647 (N_19647,N_17514,N_15043);
or U19648 (N_19648,N_18199,N_16177);
nand U19649 (N_19649,N_18071,N_15779);
xor U19650 (N_19650,N_12633,N_17357);
nor U19651 (N_19651,N_12521,N_16129);
nor U19652 (N_19652,N_14341,N_13968);
xor U19653 (N_19653,N_13029,N_18420);
or U19654 (N_19654,N_14298,N_18309);
nor U19655 (N_19655,N_16870,N_16272);
nand U19656 (N_19656,N_18432,N_14643);
xor U19657 (N_19657,N_14728,N_15193);
nor U19658 (N_19658,N_14477,N_16909);
or U19659 (N_19659,N_14868,N_16044);
or U19660 (N_19660,N_17861,N_17442);
and U19661 (N_19661,N_14601,N_16545);
and U19662 (N_19662,N_12519,N_13031);
nand U19663 (N_19663,N_17656,N_16928);
and U19664 (N_19664,N_12737,N_18502);
nand U19665 (N_19665,N_14410,N_12736);
nor U19666 (N_19666,N_12614,N_17175);
xnor U19667 (N_19667,N_14878,N_14824);
nor U19668 (N_19668,N_18139,N_18288);
nand U19669 (N_19669,N_14880,N_13801);
nor U19670 (N_19670,N_13049,N_12797);
or U19671 (N_19671,N_17356,N_12510);
nand U19672 (N_19672,N_16609,N_15598);
nand U19673 (N_19673,N_17698,N_12767);
nor U19674 (N_19674,N_15090,N_17858);
nand U19675 (N_19675,N_16126,N_17925);
nor U19676 (N_19676,N_15777,N_13815);
nor U19677 (N_19677,N_15244,N_18354);
nor U19678 (N_19678,N_17475,N_16680);
xnor U19679 (N_19679,N_14334,N_17783);
xor U19680 (N_19680,N_12544,N_15040);
or U19681 (N_19681,N_16449,N_17399);
nand U19682 (N_19682,N_18384,N_12517);
and U19683 (N_19683,N_13913,N_13096);
or U19684 (N_19684,N_17075,N_17894);
nor U19685 (N_19685,N_14554,N_15368);
or U19686 (N_19686,N_13434,N_13182);
and U19687 (N_19687,N_15918,N_12683);
nand U19688 (N_19688,N_16117,N_16388);
or U19689 (N_19689,N_14110,N_16255);
xnor U19690 (N_19690,N_12623,N_17969);
nand U19691 (N_19691,N_13991,N_17280);
nand U19692 (N_19692,N_18553,N_18187);
xor U19693 (N_19693,N_16807,N_14556);
and U19694 (N_19694,N_15078,N_14649);
xor U19695 (N_19695,N_13130,N_18680);
and U19696 (N_19696,N_14145,N_13378);
nor U19697 (N_19697,N_16551,N_18176);
nand U19698 (N_19698,N_13034,N_16391);
xor U19699 (N_19699,N_14301,N_18166);
nor U19700 (N_19700,N_15400,N_16365);
xnor U19701 (N_19701,N_16274,N_17097);
nor U19702 (N_19702,N_13441,N_18342);
or U19703 (N_19703,N_15447,N_15088);
nor U19704 (N_19704,N_13964,N_17317);
xnor U19705 (N_19705,N_16921,N_16078);
nor U19706 (N_19706,N_16484,N_14394);
xnor U19707 (N_19707,N_12511,N_13095);
xnor U19708 (N_19708,N_16689,N_14631);
xor U19709 (N_19709,N_12805,N_14275);
nor U19710 (N_19710,N_13643,N_18739);
xor U19711 (N_19711,N_15975,N_15466);
and U19712 (N_19712,N_17093,N_18703);
nand U19713 (N_19713,N_18628,N_13368);
nor U19714 (N_19714,N_13375,N_14264);
or U19715 (N_19715,N_16103,N_12828);
nor U19716 (N_19716,N_13167,N_18164);
or U19717 (N_19717,N_15625,N_13436);
or U19718 (N_19718,N_12941,N_15992);
xor U19719 (N_19719,N_14079,N_15008);
xor U19720 (N_19720,N_16265,N_18467);
nor U19721 (N_19721,N_12604,N_18254);
or U19722 (N_19722,N_18707,N_15999);
and U19723 (N_19723,N_16023,N_13307);
and U19724 (N_19724,N_18632,N_17767);
nand U19725 (N_19725,N_16759,N_16364);
nand U19726 (N_19726,N_15108,N_14822);
and U19727 (N_19727,N_13930,N_16683);
and U19728 (N_19728,N_15845,N_13295);
and U19729 (N_19729,N_14351,N_17381);
xor U19730 (N_19730,N_16703,N_13879);
and U19731 (N_19731,N_16220,N_17030);
nor U19732 (N_19732,N_16949,N_12816);
and U19733 (N_19733,N_15619,N_14489);
xnor U19734 (N_19734,N_15880,N_13576);
nor U19735 (N_19735,N_15731,N_16861);
and U19736 (N_19736,N_15654,N_12862);
and U19737 (N_19737,N_14915,N_16166);
xnor U19738 (N_19738,N_16199,N_15956);
and U19739 (N_19739,N_18737,N_17467);
or U19740 (N_19740,N_14730,N_18246);
or U19741 (N_19741,N_15868,N_14331);
xnor U19742 (N_19742,N_17587,N_15192);
nor U19743 (N_19743,N_14130,N_13315);
or U19744 (N_19744,N_14217,N_17174);
and U19745 (N_19745,N_15225,N_14603);
xor U19746 (N_19746,N_13170,N_17227);
or U19747 (N_19747,N_14382,N_13137);
nor U19748 (N_19748,N_15807,N_16027);
or U19749 (N_19749,N_13748,N_16644);
or U19750 (N_19750,N_14744,N_14518);
and U19751 (N_19751,N_12588,N_15791);
or U19752 (N_19752,N_16698,N_17779);
xnor U19753 (N_19753,N_13093,N_17446);
nor U19754 (N_19754,N_15606,N_12786);
xor U19755 (N_19755,N_13893,N_15038);
xnor U19756 (N_19756,N_17719,N_16337);
nand U19757 (N_19757,N_14274,N_13060);
xor U19758 (N_19758,N_13710,N_18508);
xnor U19759 (N_19759,N_13654,N_17171);
and U19760 (N_19760,N_17687,N_12740);
nand U19761 (N_19761,N_17101,N_14844);
nand U19762 (N_19762,N_13888,N_18092);
xor U19763 (N_19763,N_14502,N_13446);
and U19764 (N_19764,N_18337,N_16312);
nor U19765 (N_19765,N_13963,N_16443);
xor U19766 (N_19766,N_13361,N_15995);
and U19767 (N_19767,N_14528,N_16105);
nor U19768 (N_19768,N_13892,N_16773);
nor U19769 (N_19769,N_15650,N_15895);
nor U19770 (N_19770,N_15624,N_17476);
nor U19771 (N_19771,N_17286,N_18259);
or U19772 (N_19772,N_17775,N_12991);
and U19773 (N_19773,N_15815,N_13003);
or U19774 (N_19774,N_18516,N_15259);
nand U19775 (N_19775,N_18243,N_13542);
nor U19776 (N_19776,N_14653,N_14581);
nand U19777 (N_19777,N_15208,N_18495);
xnor U19778 (N_19778,N_14327,N_15826);
xnor U19779 (N_19779,N_15890,N_15340);
or U19780 (N_19780,N_14479,N_12587);
nor U19781 (N_19781,N_16750,N_18455);
nor U19782 (N_19782,N_14675,N_18500);
nor U19783 (N_19783,N_17693,N_14869);
xor U19784 (N_19784,N_16378,N_14125);
xnor U19785 (N_19785,N_15098,N_16317);
and U19786 (N_19786,N_13796,N_18103);
and U19787 (N_19787,N_13056,N_14124);
xnor U19788 (N_19788,N_14902,N_15884);
nor U19789 (N_19789,N_15713,N_17296);
and U19790 (N_19790,N_15715,N_16332);
nor U19791 (N_19791,N_17998,N_12856);
nor U19792 (N_19792,N_12893,N_17473);
nand U19793 (N_19793,N_15387,N_13274);
and U19794 (N_19794,N_18631,N_15858);
nand U19795 (N_19795,N_17050,N_13473);
nand U19796 (N_19796,N_17436,N_15614);
nor U19797 (N_19797,N_14994,N_16497);
nand U19798 (N_19798,N_12575,N_13566);
xnor U19799 (N_19799,N_15936,N_17597);
nand U19800 (N_19800,N_15914,N_13367);
nand U19801 (N_19801,N_12653,N_15793);
and U19802 (N_19802,N_16958,N_18137);
xnor U19803 (N_19803,N_14974,N_15677);
and U19804 (N_19804,N_13537,N_12776);
nor U19805 (N_19805,N_14147,N_14828);
xnor U19806 (N_19806,N_14742,N_17427);
nand U19807 (N_19807,N_14920,N_12763);
xnor U19808 (N_19808,N_17363,N_16915);
and U19809 (N_19809,N_13722,N_12573);
xnor U19810 (N_19810,N_18244,N_15723);
nand U19811 (N_19811,N_15457,N_16900);
or U19812 (N_19812,N_14035,N_17029);
xnor U19813 (N_19813,N_17393,N_18180);
nand U19814 (N_19814,N_15129,N_17157);
nor U19815 (N_19815,N_14546,N_13765);
nand U19816 (N_19816,N_13868,N_12954);
and U19817 (N_19817,N_15114,N_18562);
and U19818 (N_19818,N_15118,N_18610);
nor U19819 (N_19819,N_15423,N_14099);
or U19820 (N_19820,N_16405,N_18489);
xor U19821 (N_19821,N_14606,N_13690);
or U19822 (N_19822,N_16941,N_15722);
or U19823 (N_19823,N_16379,N_13353);
and U19824 (N_19824,N_14845,N_18734);
nor U19825 (N_19825,N_12851,N_15509);
nor U19826 (N_19826,N_15939,N_12522);
and U19827 (N_19827,N_14651,N_16247);
xnor U19828 (N_19828,N_18208,N_13701);
and U19829 (N_19829,N_14691,N_17423);
and U19830 (N_19830,N_15620,N_15796);
xor U19831 (N_19831,N_14087,N_17318);
nand U19832 (N_19832,N_18518,N_13398);
or U19833 (N_19833,N_16448,N_16180);
and U19834 (N_19834,N_15196,N_17015);
nand U19835 (N_19835,N_15105,N_12768);
and U19836 (N_19836,N_14018,N_17482);
nand U19837 (N_19837,N_13041,N_13166);
and U19838 (N_19838,N_16679,N_16686);
xnor U19839 (N_19839,N_15942,N_16972);
and U19840 (N_19840,N_15179,N_13618);
nand U19841 (N_19841,N_16738,N_15631);
nand U19842 (N_19842,N_17711,N_12558);
or U19843 (N_19843,N_12618,N_18690);
nor U19844 (N_19844,N_16580,N_18134);
or U19845 (N_19845,N_13163,N_15844);
and U19846 (N_19846,N_18446,N_16577);
or U19847 (N_19847,N_13579,N_16932);
or U19848 (N_19848,N_18329,N_12866);
nor U19849 (N_19849,N_15637,N_16894);
and U19850 (N_19850,N_16926,N_12811);
nor U19851 (N_19851,N_16072,N_18704);
nor U19852 (N_19852,N_16999,N_15635);
nand U19853 (N_19853,N_12928,N_15545);
nand U19854 (N_19854,N_16594,N_16346);
nand U19855 (N_19855,N_15049,N_13595);
or U19856 (N_19856,N_18363,N_15591);
xor U19857 (N_19857,N_17962,N_17577);
nor U19858 (N_19858,N_17817,N_16673);
nor U19859 (N_19859,N_13819,N_17865);
and U19860 (N_19860,N_14094,N_16527);
nand U19861 (N_19861,N_16060,N_17372);
or U19862 (N_19862,N_16668,N_13268);
nor U19863 (N_19863,N_15479,N_15293);
nor U19864 (N_19864,N_17823,N_18465);
nand U19865 (N_19865,N_16039,N_12803);
and U19866 (N_19866,N_18429,N_17923);
and U19867 (N_19867,N_18531,N_18260);
xnor U19868 (N_19868,N_14146,N_12909);
nand U19869 (N_19869,N_15952,N_17278);
nor U19870 (N_19870,N_12844,N_13470);
xor U19871 (N_19871,N_15181,N_17518);
or U19872 (N_19872,N_13109,N_16195);
nand U19873 (N_19873,N_13426,N_14458);
xnor U19874 (N_19874,N_13573,N_17394);
or U19875 (N_19875,N_13018,N_14929);
nand U19876 (N_19876,N_18661,N_15644);
nand U19877 (N_19877,N_18419,N_13214);
nand U19878 (N_19878,N_17763,N_18473);
or U19879 (N_19879,N_15866,N_17385);
and U19880 (N_19880,N_16521,N_12649);
and U19881 (N_19881,N_17008,N_13763);
and U19882 (N_19882,N_15382,N_13871);
xor U19883 (N_19883,N_17173,N_18202);
xor U19884 (N_19884,N_13347,N_14976);
xor U19885 (N_19885,N_13622,N_16385);
or U19886 (N_19886,N_16879,N_14368);
xor U19887 (N_19887,N_12912,N_15245);
or U19888 (N_19888,N_14168,N_16705);
or U19889 (N_19889,N_17013,N_17092);
and U19890 (N_19890,N_14682,N_16041);
or U19891 (N_19891,N_18212,N_14438);
and U19892 (N_19892,N_13282,N_17274);
xor U19893 (N_19893,N_13273,N_12918);
and U19894 (N_19894,N_14962,N_13127);
xnor U19895 (N_19895,N_15957,N_15565);
xor U19896 (N_19896,N_13025,N_17247);
xnor U19897 (N_19897,N_14358,N_15334);
or U19898 (N_19898,N_16718,N_16896);
or U19899 (N_19899,N_18457,N_14188);
nand U19900 (N_19900,N_14196,N_12727);
or U19901 (N_19901,N_16517,N_17260);
nor U19902 (N_19902,N_17971,N_12539);
nor U19903 (N_19903,N_16690,N_13793);
and U19904 (N_19904,N_17966,N_16732);
nor U19905 (N_19905,N_13705,N_16603);
xnor U19906 (N_19906,N_12745,N_17649);
or U19907 (N_19907,N_17525,N_17195);
nand U19908 (N_19908,N_13517,N_16473);
or U19909 (N_19909,N_17209,N_18538);
or U19910 (N_19910,N_12508,N_18535);
xnor U19911 (N_19911,N_15329,N_15912);
and U19912 (N_19912,N_18466,N_15077);
or U19913 (N_19913,N_12933,N_15472);
nor U19914 (N_19914,N_17913,N_17908);
or U19915 (N_19915,N_14815,N_15972);
xor U19916 (N_19916,N_12744,N_18519);
xnor U19917 (N_19917,N_17420,N_17197);
or U19918 (N_19918,N_18338,N_15145);
nand U19919 (N_19919,N_16808,N_15022);
and U19920 (N_19920,N_13148,N_14849);
and U19921 (N_19921,N_18374,N_16720);
xor U19922 (N_19922,N_14642,N_13283);
xor U19923 (N_19923,N_14640,N_17035);
xor U19924 (N_19924,N_16748,N_14093);
nand U19925 (N_19925,N_17455,N_16089);
nand U19926 (N_19926,N_12711,N_18024);
or U19927 (N_19927,N_12947,N_17951);
nor U19928 (N_19928,N_18463,N_15148);
nand U19929 (N_19929,N_12520,N_13535);
or U19930 (N_19930,N_15348,N_18204);
and U19931 (N_19931,N_14086,N_12626);
nor U19932 (N_19932,N_18522,N_14220);
and U19933 (N_19933,N_18563,N_13222);
and U19934 (N_19934,N_15081,N_13877);
xor U19935 (N_19935,N_13078,N_15642);
xor U19936 (N_19936,N_18050,N_15191);
xor U19937 (N_19937,N_15740,N_15247);
nand U19938 (N_19938,N_15321,N_14203);
nand U19939 (N_19939,N_13697,N_17670);
or U19940 (N_19940,N_14476,N_17037);
xnor U19941 (N_19941,N_18012,N_16981);
and U19942 (N_19942,N_18629,N_13070);
nor U19943 (N_19943,N_16873,N_16890);
and U19944 (N_19944,N_13564,N_16393);
or U19945 (N_19945,N_17226,N_13053);
or U19946 (N_19946,N_16503,N_13615);
xor U19947 (N_19947,N_18586,N_18396);
or U19948 (N_19948,N_16504,N_15744);
nand U19949 (N_19949,N_15592,N_14533);
or U19950 (N_19950,N_12761,N_13106);
and U19951 (N_19951,N_17364,N_17377);
nand U19952 (N_19952,N_14216,N_14945);
xnor U19953 (N_19953,N_17071,N_15773);
xnor U19954 (N_19954,N_17388,N_13970);
nor U19955 (N_19955,N_18437,N_16728);
and U19956 (N_19956,N_16131,N_14473);
and U19957 (N_19957,N_14721,N_12612);
or U19958 (N_19958,N_14004,N_18005);
or U19959 (N_19959,N_15638,N_14379);
or U19960 (N_19960,N_12906,N_15485);
xnor U19961 (N_19961,N_15900,N_13235);
nor U19962 (N_19962,N_18658,N_15304);
xnor U19963 (N_19963,N_13544,N_18469);
nor U19964 (N_19964,N_15524,N_15174);
and U19965 (N_19965,N_13215,N_18641);
nor U19966 (N_19966,N_17155,N_17373);
xor U19967 (N_19967,N_13925,N_18480);
nor U19968 (N_19968,N_17453,N_18674);
xnor U19969 (N_19969,N_13895,N_16618);
nor U19970 (N_19970,N_13715,N_13971);
xor U19971 (N_19971,N_14752,N_14677);
and U19972 (N_19972,N_18159,N_12976);
nand U19973 (N_19973,N_15281,N_13896);
xnor U19974 (N_19974,N_17774,N_17468);
xnor U19975 (N_19975,N_16190,N_15585);
nor U19976 (N_19976,N_12770,N_17342);
xnor U19977 (N_19977,N_17921,N_13218);
or U19978 (N_19978,N_12845,N_17764);
or U19979 (N_19979,N_17011,N_15236);
nor U19980 (N_19980,N_16357,N_16270);
nor U19981 (N_19981,N_13607,N_12706);
xnor U19982 (N_19982,N_17140,N_13354);
or U19983 (N_19983,N_15928,N_15932);
nor U19984 (N_19984,N_14663,N_18277);
or U19985 (N_19985,N_15006,N_12751);
and U19986 (N_19986,N_17685,N_13411);
and U19987 (N_19987,N_14427,N_15647);
nand U19988 (N_19988,N_17523,N_17079);
nor U19989 (N_19989,N_17671,N_12645);
nor U19990 (N_19990,N_15376,N_15589);
nand U19991 (N_19991,N_18074,N_13262);
nand U19992 (N_19992,N_15278,N_17127);
and U19993 (N_19993,N_16127,N_16136);
or U19994 (N_19994,N_12747,N_18007);
xor U19995 (N_19995,N_17989,N_13173);
nand U19996 (N_19996,N_13758,N_14989);
xnor U19997 (N_19997,N_15211,N_15113);
nand U19998 (N_19998,N_14486,N_15794);
and U19999 (N_19999,N_13151,N_17562);
nor U20000 (N_20000,N_14342,N_16826);
nor U20001 (N_20001,N_17344,N_12641);
nand U20002 (N_20002,N_15684,N_15228);
nand U20003 (N_20003,N_12617,N_15254);
or U20004 (N_20004,N_16825,N_12937);
or U20005 (N_20005,N_18558,N_12769);
nor U20006 (N_20006,N_15767,N_15725);
or U20007 (N_20007,N_18084,N_14156);
xnor U20008 (N_20008,N_18196,N_16211);
nand U20009 (N_20009,N_15056,N_13619);
and U20010 (N_20010,N_16887,N_13854);
and U20011 (N_20011,N_15981,N_12668);
xor U20012 (N_20012,N_13035,N_17070);
and U20013 (N_20013,N_14319,N_18454);
nor U20014 (N_20014,N_14594,N_13779);
xnor U20015 (N_20015,N_17360,N_16939);
and U20016 (N_20016,N_17366,N_13213);
xnor U20017 (N_20017,N_16111,N_18443);
and U20018 (N_20018,N_14725,N_13211);
nand U20019 (N_20019,N_17980,N_14623);
or U20020 (N_20020,N_18430,N_15902);
nand U20021 (N_20021,N_14271,N_17659);
or U20022 (N_20022,N_16631,N_15588);
or U20023 (N_20023,N_17440,N_15668);
nand U20024 (N_20024,N_14760,N_14843);
nand U20025 (N_20025,N_17439,N_16853);
xor U20026 (N_20026,N_17108,N_14280);
nand U20027 (N_20027,N_16995,N_14563);
nor U20028 (N_20028,N_16338,N_12739);
or U20029 (N_20029,N_13495,N_16498);
nand U20030 (N_20030,N_14091,N_13669);
nand U20031 (N_20031,N_16284,N_14027);
and U20032 (N_20032,N_14070,N_14805);
and U20033 (N_20033,N_16411,N_15075);
and U20034 (N_20034,N_15425,N_16692);
or U20035 (N_20035,N_17413,N_13703);
nor U20036 (N_20036,N_18117,N_15905);
nand U20037 (N_20037,N_16074,N_16614);
and U20038 (N_20038,N_18112,N_18146);
and U20039 (N_20039,N_13129,N_18281);
xnor U20040 (N_20040,N_15921,N_17876);
or U20041 (N_20041,N_16905,N_16823);
or U20042 (N_20042,N_18336,N_17617);
nand U20043 (N_20043,N_18238,N_17757);
xor U20044 (N_20044,N_14895,N_18069);
and U20045 (N_20045,N_15747,N_14602);
and U20046 (N_20046,N_13764,N_15692);
or U20047 (N_20047,N_16908,N_16038);
xnor U20048 (N_20048,N_14821,N_15573);
nor U20049 (N_20049,N_15214,N_15094);
nand U20050 (N_20050,N_13202,N_18431);
nor U20051 (N_20051,N_13585,N_15000);
or U20052 (N_20052,N_18619,N_15801);
nand U20053 (N_20053,N_16140,N_14981);
nand U20054 (N_20054,N_15394,N_13780);
xnor U20055 (N_20055,N_18686,N_13023);
and U20056 (N_20056,N_16839,N_16253);
xnor U20057 (N_20057,N_13417,N_16539);
or U20058 (N_20058,N_15851,N_12691);
xnor U20059 (N_20059,N_16532,N_15037);
nor U20060 (N_20060,N_12565,N_16106);
and U20061 (N_20061,N_13664,N_15660);
or U20062 (N_20062,N_18253,N_17382);
nor U20063 (N_20063,N_14065,N_15396);
nand U20064 (N_20064,N_14968,N_16627);
xor U20065 (N_20065,N_13090,N_18622);
and U20066 (N_20066,N_17645,N_13798);
nand U20067 (N_20067,N_13633,N_13969);
xnor U20068 (N_20068,N_17692,N_16821);
and U20069 (N_20069,N_13281,N_16633);
or U20070 (N_20070,N_14922,N_13371);
and U20071 (N_20071,N_18195,N_13915);
xor U20072 (N_20072,N_15312,N_14778);
and U20073 (N_20073,N_15020,N_17487);
nor U20074 (N_20074,N_14173,N_13954);
and U20075 (N_20075,N_13511,N_15935);
xor U20076 (N_20076,N_12850,N_18080);
xor U20077 (N_20077,N_14122,N_16124);
xor U20078 (N_20078,N_13028,N_16426);
or U20079 (N_20079,N_15886,N_17089);
and U20080 (N_20080,N_15745,N_15711);
and U20081 (N_20081,N_13351,N_14326);
nand U20082 (N_20082,N_16147,N_17512);
or U20083 (N_20083,N_14680,N_17292);
xor U20084 (N_20084,N_13091,N_16007);
or U20085 (N_20085,N_13442,N_13588);
nor U20086 (N_20086,N_18178,N_15696);
and U20087 (N_20087,N_17198,N_18105);
and U20088 (N_20088,N_15054,N_16298);
nor U20089 (N_20089,N_14448,N_17252);
or U20090 (N_20090,N_15920,N_16888);
and U20091 (N_20091,N_16148,N_18366);
or U20092 (N_20092,N_13227,N_15695);
xnor U20093 (N_20093,N_14138,N_16441);
xor U20094 (N_20094,N_13231,N_14693);
nand U20095 (N_20095,N_18588,N_18568);
nor U20096 (N_20096,N_18530,N_14984);
xnor U20097 (N_20097,N_15153,N_15079);
and U20098 (N_20098,N_17237,N_13504);
nor U20099 (N_20099,N_15559,N_13521);
xor U20100 (N_20100,N_14012,N_17009);
and U20101 (N_20101,N_13782,N_15488);
and U20102 (N_20102,N_15824,N_16244);
nand U20103 (N_20103,N_18511,N_14810);
or U20104 (N_20104,N_13768,N_13720);
or U20105 (N_20105,N_18715,N_13695);
and U20106 (N_20106,N_12757,N_17811);
and U20107 (N_20107,N_14430,N_14318);
or U20108 (N_20108,N_12884,N_18720);
or U20109 (N_20109,N_14678,N_15172);
nor U20110 (N_20110,N_14291,N_13639);
or U20111 (N_20111,N_16183,N_14517);
nor U20112 (N_20112,N_13335,N_14491);
xor U20113 (N_20113,N_17978,N_12680);
and U20114 (N_20114,N_17634,N_16245);
nor U20115 (N_20115,N_13704,N_18647);
nand U20116 (N_20116,N_18373,N_16651);
nand U20117 (N_20117,N_14450,N_12710);
or U20118 (N_20118,N_12537,N_14615);
xnor U20119 (N_20119,N_13248,N_15772);
nor U20120 (N_20120,N_18570,N_16293);
and U20121 (N_20121,N_17149,N_15906);
nor U20122 (N_20122,N_14669,N_18727);
xor U20123 (N_20123,N_14310,N_14175);
nor U20124 (N_20124,N_15566,N_16980);
or U20125 (N_20125,N_15005,N_17920);
nand U20126 (N_20126,N_13706,N_15720);
xnor U20127 (N_20127,N_15111,N_17426);
or U20128 (N_20128,N_16260,N_12936);
or U20129 (N_20129,N_17995,N_16803);
nor U20130 (N_20130,N_16054,N_18064);
and U20131 (N_20131,N_14827,N_14435);
or U20132 (N_20132,N_15045,N_15342);
and U20133 (N_20133,N_15327,N_17498);
or U20134 (N_20134,N_12914,N_12814);
or U20135 (N_20135,N_12843,N_13043);
and U20136 (N_20136,N_15494,N_15359);
and U20137 (N_20137,N_14709,N_16188);
nand U20138 (N_20138,N_12716,N_15561);
nor U20139 (N_20139,N_17343,N_18214);
xor U20140 (N_20140,N_14793,N_18461);
nor U20141 (N_20141,N_13198,N_14524);
or U20142 (N_20142,N_18716,N_12677);
and U20143 (N_20143,N_14006,N_18554);
xnor U20144 (N_20144,N_15099,N_14178);
xnor U20145 (N_20145,N_18351,N_14509);
and U20146 (N_20146,N_16012,N_14806);
nor U20147 (N_20147,N_17831,N_15822);
and U20148 (N_20148,N_17708,N_14025);
xnor U20149 (N_20149,N_16913,N_13528);
nor U20150 (N_20150,N_16630,N_15697);
xnor U20151 (N_20151,N_13844,N_16380);
nor U20152 (N_20152,N_16092,N_12859);
xnor U20153 (N_20153,N_13279,N_15491);
nand U20154 (N_20154,N_18667,N_15352);
xnor U20155 (N_20155,N_14397,N_15255);
nor U20156 (N_20156,N_13776,N_13369);
or U20157 (N_20157,N_14447,N_12718);
xnor U20158 (N_20158,N_13933,N_13519);
nor U20159 (N_20159,N_18300,N_13444);
nand U20160 (N_20160,N_15165,N_13712);
and U20161 (N_20161,N_16499,N_13217);
or U20162 (N_20162,N_13374,N_17417);
nor U20163 (N_20163,N_15623,N_15477);
nand U20164 (N_20164,N_15197,N_17772);
xor U20165 (N_20165,N_16657,N_13237);
and U20166 (N_20166,N_18347,N_13072);
nor U20167 (N_20167,N_17503,N_15083);
and U20168 (N_20168,N_14105,N_13711);
nand U20169 (N_20169,N_13261,N_12647);
xor U20170 (N_20170,N_13311,N_18330);
and U20171 (N_20171,N_17056,N_14646);
xor U20172 (N_20172,N_14375,N_17821);
nand U20173 (N_20173,N_13767,N_17977);
xor U20174 (N_20174,N_15916,N_17880);
nor U20175 (N_20175,N_13496,N_14266);
nand U20176 (N_20176,N_13157,N_13629);
and U20177 (N_20177,N_13986,N_13620);
and U20178 (N_20178,N_16071,N_15742);
nor U20179 (N_20179,N_17590,N_13642);
nand U20180 (N_20180,N_13994,N_13610);
nand U20181 (N_20181,N_17240,N_17884);
and U20182 (N_20182,N_17633,N_15511);
xnor U20183 (N_20183,N_15429,N_12916);
or U20184 (N_20184,N_14493,N_18286);
nor U20185 (N_20185,N_14668,N_14573);
or U20186 (N_20186,N_16150,N_16125);
nor U20187 (N_20187,N_16450,N_15087);
and U20188 (N_20188,N_15104,N_13876);
or U20189 (N_20189,N_14535,N_16447);
nand U20190 (N_20190,N_16788,N_14255);
and U20191 (N_20191,N_13927,N_13902);
nor U20192 (N_20192,N_16322,N_17961);
and U20193 (N_20193,N_13476,N_14614);
and U20194 (N_20194,N_15424,N_18651);
and U20195 (N_20195,N_15017,N_14607);
or U20196 (N_20196,N_17233,N_17095);
and U20197 (N_20197,N_14697,N_18422);
nor U20198 (N_20198,N_14487,N_18670);
nor U20199 (N_20199,N_15622,N_15602);
nand U20200 (N_20200,N_13190,N_13205);
nand U20201 (N_20201,N_15018,N_17898);
nand U20202 (N_20202,N_18315,N_16961);
nand U20203 (N_20203,N_14340,N_13837);
and U20204 (N_20204,N_13373,N_16389);
xor U20205 (N_20205,N_16455,N_17839);
and U20206 (N_20206,N_16872,N_18107);
nor U20207 (N_20207,N_15693,N_14841);
xor U20208 (N_20208,N_16359,N_13039);
nand U20209 (N_20209,N_12876,N_14904);
and U20210 (N_20210,N_14629,N_14560);
xnor U20211 (N_20211,N_14897,N_17349);
nor U20212 (N_20212,N_18310,N_14670);
nor U20213 (N_20213,N_17248,N_14423);
nand U20214 (N_20214,N_13250,N_13395);
or U20215 (N_20215,N_16182,N_16418);
xnor U20216 (N_20216,N_17714,N_18056);
nand U20217 (N_20217,N_16034,N_15149);
xor U20218 (N_20218,N_12950,N_12530);
nand U20219 (N_20219,N_16169,N_17200);
and U20220 (N_20220,N_13640,N_17615);
nand U20221 (N_20221,N_13098,N_14160);
nor U20222 (N_20222,N_17531,N_17844);
xnor U20223 (N_20223,N_13253,N_15555);
and U20224 (N_20224,N_16585,N_17967);
nand U20225 (N_20225,N_18507,N_16925);
nor U20226 (N_20226,N_18694,N_16607);
xnor U20227 (N_20227,N_17365,N_16579);
and U20228 (N_20228,N_16942,N_14305);
or U20229 (N_20229,N_14754,N_13437);
or U20230 (N_20230,N_13482,N_17674);
or U20231 (N_20231,N_18090,N_17709);
and U20232 (N_20232,N_15362,N_16438);
nand U20233 (N_20233,N_18348,N_17180);
and U20234 (N_20234,N_16876,N_17769);
xor U20235 (N_20235,N_17578,N_16561);
nand U20236 (N_20236,N_18435,N_16068);
and U20237 (N_20237,N_18221,N_13299);
or U20238 (N_20238,N_12800,N_15282);
or U20239 (N_20239,N_14708,N_18546);
xor U20240 (N_20240,N_14344,N_14909);
and U20241 (N_20241,N_12778,N_14800);
and U20242 (N_20242,N_17910,N_14523);
and U20243 (N_20243,N_15663,N_13757);
and U20244 (N_20244,N_16275,N_13179);
nand U20245 (N_20245,N_13483,N_13836);
nand U20246 (N_20246,N_13440,N_17094);
nand U20247 (N_20247,N_15849,N_17899);
and U20248 (N_20248,N_14967,N_14047);
and U20249 (N_20249,N_17555,N_16314);
xnor U20250 (N_20250,N_16083,N_12512);
or U20251 (N_20251,N_16982,N_18276);
and U20252 (N_20252,N_14839,N_15320);
xor U20253 (N_20253,N_18158,N_14161);
or U20254 (N_20254,N_16184,N_17976);
nand U20255 (N_20255,N_15233,N_15461);
nor U20256 (N_20256,N_18335,N_17643);
and U20257 (N_20257,N_17973,N_13770);
nor U20258 (N_20258,N_16334,N_17137);
and U20259 (N_20259,N_17256,N_14703);
xnor U20260 (N_20260,N_13433,N_17059);
xnor U20261 (N_20261,N_16305,N_13670);
nor U20262 (N_20262,N_14932,N_13475);
or U20263 (N_20263,N_17332,N_12748);
xnor U20264 (N_20264,N_17276,N_18296);
and U20265 (N_20265,N_14355,N_16101);
nand U20266 (N_20266,N_13225,N_16115);
xnor U20267 (N_20267,N_16079,N_16176);
or U20268 (N_20268,N_14903,N_14414);
nor U20269 (N_20269,N_15850,N_14769);
nand U20270 (N_20270,N_12979,N_16979);
or U20271 (N_20271,N_18033,N_13328);
nor U20272 (N_20272,N_16893,N_16370);
or U20273 (N_20273,N_17113,N_14249);
or U20274 (N_20274,N_12666,N_13145);
xnor U20275 (N_20275,N_15404,N_14978);
nor U20276 (N_20276,N_13045,N_13085);
nand U20277 (N_20277,N_16159,N_14218);
xnor U20278 (N_20278,N_18700,N_12538);
nor U20279 (N_20279,N_13992,N_12639);
and U20280 (N_20280,N_15876,N_14393);
nand U20281 (N_20281,N_16186,N_14561);
xor U20282 (N_20282,N_17379,N_17106);
nor U20283 (N_20283,N_15256,N_16797);
nor U20284 (N_20284,N_14787,N_13531);
nor U20285 (N_20285,N_14505,N_17647);
nand U20286 (N_20286,N_17798,N_17328);
or U20287 (N_20287,N_16877,N_16572);
nand U20288 (N_20288,N_13459,N_16891);
nand U20289 (N_20289,N_12858,N_17528);
xor U20290 (N_20290,N_16769,N_18718);
nor U20291 (N_20291,N_17915,N_15803);
nor U20292 (N_20292,N_12507,N_12637);
and U20293 (N_20293,N_15708,N_17722);
and U20294 (N_20294,N_14059,N_18038);
nand U20295 (N_20295,N_13600,N_14113);
or U20296 (N_20296,N_17339,N_15833);
or U20297 (N_20297,N_18267,N_13667);
nand U20298 (N_20298,N_18581,N_16625);
nor U20299 (N_20299,N_18368,N_14702);
or U20300 (N_20300,N_17660,N_17182);
nand U20301 (N_20301,N_17529,N_15216);
nor U20302 (N_20302,N_17172,N_17825);
xnor U20303 (N_20303,N_14184,N_18542);
nor U20304 (N_20304,N_16524,N_18685);
or U20305 (N_20305,N_13714,N_15323);
nand U20306 (N_20306,N_16428,N_14954);
xor U20307 (N_20307,N_14349,N_15673);
and U20308 (N_20308,N_13536,N_15656);
xor U20309 (N_20309,N_18456,N_18165);
and U20310 (N_20310,N_17147,N_17254);
xor U20311 (N_20311,N_18041,N_15273);
and U20312 (N_20312,N_13484,N_15150);
and U20313 (N_20313,N_12534,N_16665);
and U20314 (N_20314,N_14936,N_12815);
or U20315 (N_20315,N_15266,N_15539);
xor U20316 (N_20316,N_18082,N_13493);
and U20317 (N_20317,N_16917,N_18646);
nor U20318 (N_20318,N_13206,N_14270);
nand U20319 (N_20319,N_15556,N_13735);
or U20320 (N_20320,N_18203,N_12971);
or U20321 (N_20321,N_12665,N_16010);
nor U20322 (N_20322,N_14015,N_16881);
or U20323 (N_20323,N_14853,N_14484);
or U20324 (N_20324,N_17319,N_12702);
xor U20325 (N_20325,N_17810,N_14192);
xor U20326 (N_20326,N_18526,N_18106);
nand U20327 (N_20327,N_13358,N_16454);
and U20328 (N_20328,N_12785,N_13559);
and U20329 (N_20329,N_13193,N_16367);
and U20330 (N_20330,N_14711,N_13777);
nor U20331 (N_20331,N_13118,N_13613);
nand U20332 (N_20332,N_16729,N_15332);
nor U20333 (N_20333,N_18602,N_16782);
xor U20334 (N_20334,N_15445,N_12891);
nor U20335 (N_20335,N_12528,N_14764);
or U20336 (N_20336,N_16509,N_16269);
xnor U20337 (N_20337,N_14564,N_15493);
or U20338 (N_20338,N_17950,N_18404);
and U20339 (N_20339,N_17052,N_17928);
nor U20340 (N_20340,N_13380,N_13464);
nand U20341 (N_20341,N_14050,N_16541);
or U20342 (N_20342,N_14328,N_14353);
xor U20343 (N_20343,N_16022,N_13628);
nor U20344 (N_20344,N_15298,N_16582);
xor U20345 (N_20345,N_18045,N_16347);
and U20346 (N_20346,N_16087,N_15641);
nor U20347 (N_20347,N_13660,N_16711);
nand U20348 (N_20348,N_16416,N_12562);
and U20349 (N_20349,N_14570,N_15522);
nand U20350 (N_20350,N_18006,N_17974);
nand U20351 (N_20351,N_18598,N_12847);
or U20352 (N_20352,N_12895,N_16934);
nand U20353 (N_20353,N_13203,N_17947);
or U20354 (N_20354,N_15487,N_14183);
or U20355 (N_20355,N_17018,N_13026);
nor U20356 (N_20356,N_13753,N_16290);
nand U20357 (N_20357,N_15878,N_16514);
or U20358 (N_20358,N_12560,N_15237);
or U20359 (N_20359,N_14128,N_14116);
or U20360 (N_20360,N_15463,N_16050);
xor U20361 (N_20361,N_14010,N_17600);
nor U20362 (N_20362,N_16735,N_17479);
and U20363 (N_20363,N_14655,N_14499);
nor U20364 (N_20364,N_18060,N_16070);
and U20365 (N_20365,N_13191,N_12719);
or U20366 (N_20366,N_14245,N_12728);
nand U20367 (N_20367,N_18626,N_18499);
nor U20368 (N_20368,N_16765,N_12806);
nand U20369 (N_20369,N_15194,N_17389);
and U20370 (N_20370,N_14041,N_16386);
xor U20371 (N_20371,N_12881,N_15319);
and U20372 (N_20372,N_15934,N_13105);
or U20373 (N_20373,N_15578,N_12855);
and U20374 (N_20374,N_18201,N_17970);
nand U20375 (N_20375,N_17306,N_18543);
and U20376 (N_20376,N_13171,N_18292);
and U20377 (N_20377,N_17123,N_15575);
xor U20378 (N_20378,N_16104,N_15389);
and U20379 (N_20379,N_14749,N_13838);
nor U20380 (N_20380,N_18405,N_13081);
or U20381 (N_20381,N_16206,N_15395);
nor U20382 (N_20382,N_16569,N_12760);
nor U20383 (N_20383,N_17450,N_16175);
xnor U20384 (N_20384,N_12651,N_13804);
and U20385 (N_20385,N_14736,N_17026);
nor U20386 (N_20386,N_18659,N_12999);
nand U20387 (N_20387,N_17303,N_13759);
nor U20388 (N_20388,N_14302,N_13570);
xnor U20389 (N_20389,N_13394,N_17299);
nor U20390 (N_20390,N_14811,N_15166);
xnor U20391 (N_20391,N_17515,N_13931);
nor U20392 (N_20392,N_17474,N_12540);
nand U20393 (N_20393,N_15689,N_16860);
or U20394 (N_20394,N_15326,N_14796);
nor U20395 (N_20395,N_14297,N_14512);
nand U20396 (N_20396,N_18689,N_18587);
xor U20397 (N_20397,N_14069,N_15840);
or U20398 (N_20398,N_17412,N_12983);
xor U20399 (N_20399,N_17778,N_16646);
nor U20400 (N_20400,N_13754,N_14315);
nor U20401 (N_20401,N_16946,N_14281);
and U20402 (N_20402,N_17291,N_14550);
or U20403 (N_20403,N_13794,N_15128);
or U20404 (N_20404,N_16130,N_14707);
or U20405 (N_20405,N_14977,N_16899);
xnor U20406 (N_20406,N_15399,N_13668);
nand U20407 (N_20407,N_14661,N_15949);
xor U20408 (N_20408,N_16991,N_13806);
nor U20409 (N_20409,N_14498,N_15659);
nand U20410 (N_20410,N_13135,N_13414);
nand U20411 (N_20411,N_16300,N_13165);
xnor U20412 (N_20412,N_14768,N_15567);
or U20413 (N_20413,N_13007,N_15422);
nand U20414 (N_20414,N_15675,N_15354);
and U20415 (N_20415,N_14166,N_18537);
xnor U20416 (N_20416,N_16026,N_17091);
and U20417 (N_20417,N_16591,N_14883);
nand U20418 (N_20418,N_17124,N_13920);
nand U20419 (N_20419,N_14710,N_13232);
or U20420 (N_20420,N_17640,N_17732);
xor U20421 (N_20421,N_17749,N_17053);
and U20422 (N_20422,N_13730,N_18306);
xor U20423 (N_20423,N_16862,N_14576);
nand U20424 (N_20424,N_14391,N_17707);
or U20425 (N_20425,N_13467,N_18372);
xor U20426 (N_20426,N_15204,N_12687);
xnor U20427 (N_20427,N_16452,N_12922);
nand U20428 (N_20428,N_14149,N_14049);
and U20429 (N_20429,N_13337,N_15530);
or U20430 (N_20430,N_14999,N_18140);
nand U20431 (N_20431,N_17401,N_16018);
nand U20432 (N_20432,N_14243,N_18031);
nand U20433 (N_20433,N_18423,N_16468);
and U20434 (N_20434,N_18077,N_17935);
xor U20435 (N_20435,N_15707,N_16733);
nor U20436 (N_20436,N_15453,N_17932);
or U20437 (N_20437,N_15966,N_13742);
nor U20438 (N_20438,N_18044,N_15378);
nor U20439 (N_20439,N_12989,N_16974);
or U20440 (N_20440,N_13393,N_12730);
and U20441 (N_20441,N_13345,N_13956);
xor U20442 (N_20442,N_17346,N_18417);
and U20443 (N_20443,N_13540,N_18109);
nand U20444 (N_20444,N_15188,N_15915);
nor U20445 (N_20445,N_14464,N_18402);
nand U20446 (N_20446,N_12820,N_17706);
xnor U20447 (N_20447,N_17454,N_15508);
or U20448 (N_20448,N_15580,N_17012);
nand U20449 (N_20449,N_13958,N_14222);
nand U20450 (N_20450,N_17696,N_17043);
nor U20451 (N_20451,N_15757,N_18594);
and U20452 (N_20452,N_14766,N_14157);
nand U20453 (N_20453,N_13781,N_15124);
and U20454 (N_20454,N_17211,N_12835);
xnor U20455 (N_20455,N_13449,N_14858);
xor U20456 (N_20456,N_15055,N_14632);
nand U20457 (N_20457,N_18544,N_15316);
xor U20458 (N_20458,N_15375,N_12547);
xnor U20459 (N_20459,N_15898,N_18079);
or U20460 (N_20460,N_16084,N_12703);
nand U20461 (N_20461,N_16813,N_17269);
or U20462 (N_20462,N_18136,N_15543);
and U20463 (N_20463,N_14757,N_12609);
or U20464 (N_20464,N_18579,N_14126);
nand U20465 (N_20465,N_12655,N_14599);
nor U20466 (N_20466,N_15440,N_16210);
xor U20467 (N_20467,N_18101,N_12670);
and U20468 (N_20468,N_13396,N_18304);
or U20469 (N_20469,N_14527,N_16444);
nor U20470 (N_20470,N_15888,N_16155);
and U20471 (N_20471,N_17295,N_15716);
xor U20472 (N_20472,N_15686,N_13745);
or U20473 (N_20473,N_14381,N_16593);
xor U20474 (N_20474,N_13589,N_16469);
xnor U20475 (N_20475,N_15843,N_18332);
nand U20476 (N_20476,N_12597,N_13597);
nand U20477 (N_20477,N_15057,N_15190);
nor U20478 (N_20478,N_17055,N_14143);
xnor U20479 (N_20479,N_15080,N_15800);
nor U20480 (N_20480,N_18498,N_17178);
nand U20481 (N_20481,N_18625,N_17689);
or U20482 (N_20482,N_17258,N_18496);
nand U20483 (N_20483,N_14953,N_14809);
or U20484 (N_20484,N_14630,N_14366);
nor U20485 (N_20485,N_15755,N_16997);
xnor U20486 (N_20486,N_18100,N_16864);
xor U20487 (N_20487,N_14665,N_18133);
and U20488 (N_20488,N_14247,N_12686);
and U20489 (N_20489,N_15050,N_17320);
or U20490 (N_20490,N_18057,N_13153);
and U20491 (N_20491,N_13718,N_17700);
xnor U20492 (N_20492,N_17460,N_18630);
nor U20493 (N_20493,N_16485,N_16063);
or U20494 (N_20494,N_13783,N_17729);
nand U20495 (N_20495,N_12723,N_13953);
nand U20496 (N_20496,N_16624,N_15307);
xnor U20497 (N_20497,N_17370,N_15897);
or U20498 (N_20498,N_16201,N_18236);
or U20499 (N_20499,N_17721,N_12734);
or U20500 (N_20500,N_13822,N_14263);
nand U20501 (N_20501,N_18470,N_18512);
or U20502 (N_20502,N_17057,N_16384);
nor U20503 (N_20503,N_18642,N_13631);
or U20504 (N_20504,N_15146,N_12896);
xor U20505 (N_20505,N_17845,N_13721);
or U20506 (N_20506,N_18413,N_14820);
and U20507 (N_20507,N_17353,N_14704);
and U20508 (N_20508,N_17606,N_18378);
or U20509 (N_20509,N_15178,N_15435);
and U20510 (N_20510,N_16530,N_17627);
and U20511 (N_20511,N_17434,N_13439);
and U20512 (N_20512,N_12810,N_18085);
and U20513 (N_20513,N_17517,N_15219);
and U20514 (N_20514,N_13431,N_13560);
nand U20515 (N_20515,N_16339,N_16024);
or U20516 (N_20516,N_17930,N_12819);
xnor U20517 (N_20517,N_14540,N_17341);
xor U20518 (N_20518,N_17022,N_15505);
and U20519 (N_20519,N_16756,N_16369);
or U20520 (N_20520,N_14359,N_14198);
nand U20521 (N_20521,N_13017,N_16959);
xnor U20522 (N_20522,N_16417,N_15010);
or U20523 (N_20523,N_15393,N_13872);
or U20524 (N_20524,N_15583,N_18382);
nor U20525 (N_20525,N_16258,N_16794);
or U20526 (N_20526,N_15085,N_14650);
xnor U20527 (N_20527,N_16865,N_16742);
and U20528 (N_20528,N_18550,N_12563);
and U20529 (N_20529,N_17521,N_17841);
nand U20530 (N_20530,N_15753,N_13506);
and U20531 (N_20531,N_13574,N_12840);
nand U20532 (N_20532,N_13940,N_17904);
and U20533 (N_20533,N_18395,N_13908);
and U20534 (N_20534,N_18269,N_17688);
or U20535 (N_20535,N_14031,N_15215);
and U20536 (N_20536,N_13581,N_16109);
nand U20537 (N_20537,N_13338,N_17701);
xnor U20538 (N_20538,N_18370,N_17572);
xnor U20539 (N_20539,N_15875,N_18013);
nor U20540 (N_20540,N_15869,N_18633);
nand U20541 (N_20541,N_16531,N_17526);
or U20542 (N_20542,N_16796,N_18371);
and U20543 (N_20543,N_17462,N_17449);
xnor U20544 (N_20544,N_14562,N_13456);
nand U20545 (N_20545,N_14740,N_15976);
xor U20546 (N_20546,N_17827,N_17425);
and U20547 (N_20547,N_16343,N_17678);
xnor U20548 (N_20548,N_16313,N_16382);
and U20549 (N_20549,N_13341,N_14295);
nand U20550 (N_20550,N_15182,N_12630);
xor U20551 (N_20551,N_14656,N_15590);
or U20552 (N_20552,N_13209,N_16507);
and U20553 (N_20553,N_14279,N_17661);
nor U20554 (N_20554,N_16029,N_17852);
or U20555 (N_20555,N_17972,N_13138);
xor U20556 (N_20556,N_16837,N_18086);
xor U20557 (N_20557,N_18392,N_13309);
and U20558 (N_20558,N_12813,N_18040);
xnor U20559 (N_20559,N_18478,N_15497);
or U20560 (N_20560,N_13063,N_17221);
nand U20561 (N_20561,N_12779,N_14838);
nor U20562 (N_20562,N_14213,N_13853);
and U20563 (N_20563,N_17326,N_14673);
xnor U20564 (N_20564,N_16789,N_15523);
or U20565 (N_20565,N_12788,N_13924);
and U20566 (N_20566,N_18665,N_14325);
nand U20567 (N_20567,N_12824,N_14309);
nand U20568 (N_20568,N_16318,N_13832);
xnor U20569 (N_20569,N_15163,N_13864);
nor U20570 (N_20570,N_17836,N_15469);
or U20571 (N_20571,N_14654,N_16235);
xor U20572 (N_20572,N_14747,N_16859);
or U20573 (N_20573,N_18687,N_17607);
nor U20574 (N_20574,N_17016,N_14030);
nand U20575 (N_20575,N_16254,N_13415);
xnor U20576 (N_20576,N_12963,N_15818);
nand U20577 (N_20577,N_15609,N_14317);
nand U20578 (N_20578,N_16906,N_15448);
or U20579 (N_20579,N_15260,N_15605);
or U20580 (N_20580,N_17753,N_16295);
xor U20581 (N_20581,N_13906,N_14790);
nor U20582 (N_20582,N_18052,N_14095);
or U20583 (N_20583,N_14115,N_15351);
nand U20584 (N_20584,N_13803,N_17218);
nand U20585 (N_20585,N_14148,N_17128);
xor U20586 (N_20586,N_15264,N_16075);
nor U20587 (N_20587,N_14037,N_16841);
nor U20588 (N_20588,N_14993,N_16487);
and U20589 (N_20589,N_15940,N_16659);
xnor U20590 (N_20590,N_13952,N_16709);
nand U20591 (N_20591,N_15558,N_14501);
nand U20592 (N_20592,N_18740,N_15864);
or U20593 (N_20593,N_15680,N_12980);
nor U20594 (N_20594,N_13400,N_16303);
nor U20595 (N_20595,N_17492,N_14593);
nor U20596 (N_20596,N_15865,N_17746);
and U20597 (N_20597,N_17569,N_15611);
and U20598 (N_20598,N_18326,N_15283);
or U20599 (N_20599,N_13862,N_13296);
nand U20600 (N_20600,N_15639,N_16394);
nand U20601 (N_20601,N_12695,N_16492);
and U20602 (N_20602,N_16107,N_14835);
nor U20603 (N_20603,N_18617,N_14179);
or U20604 (N_20604,N_18303,N_12873);
or U20605 (N_20605,N_15579,N_13666);
nor U20606 (N_20606,N_17552,N_15862);
or U20607 (N_20607,N_15927,N_15156);
or U20608 (N_20608,N_12578,N_13951);
nor U20609 (N_20609,N_15979,N_13058);
and U20610 (N_20610,N_13270,N_15023);
and U20611 (N_20611,N_17438,N_15987);
or U20612 (N_20612,N_17883,N_12571);
or U20613 (N_20613,N_16232,N_15517);
nor U20614 (N_20614,N_18127,N_16145);
nor U20615 (N_20615,N_16349,N_12611);
nand U20616 (N_20616,N_18087,N_16435);
nor U20617 (N_20617,N_13551,N_15372);
xnor U20618 (N_20618,N_18059,N_18224);
and U20619 (N_20619,N_18458,N_15514);
or U20620 (N_20620,N_12766,N_14321);
and U20621 (N_20621,N_17668,N_18150);
or U20622 (N_20622,N_16308,N_13199);
or U20623 (N_20623,N_16080,N_15033);
and U20624 (N_20624,N_17002,N_13911);
xor U20625 (N_20625,N_15361,N_12902);
and U20626 (N_20626,N_15547,N_16133);
xor U20627 (N_20627,N_17954,N_15795);
or U20628 (N_20628,N_16031,N_14715);
xor U20629 (N_20629,N_15528,N_18401);
or U20630 (N_20630,N_15379,N_12514);
or U20631 (N_20631,N_14005,N_18115);
nand U20632 (N_20632,N_16178,N_18155);
xnor U20633 (N_20633,N_15743,N_13032);
or U20634 (N_20634,N_14236,N_15322);
nor U20635 (N_20635,N_14080,N_13727);
xor U20636 (N_20636,N_15217,N_13980);
xnor U20637 (N_20637,N_16955,N_12985);
or U20638 (N_20638,N_17756,N_17471);
and U20639 (N_20639,N_12960,N_16213);
and U20640 (N_20640,N_17184,N_13530);
xnor U20641 (N_20641,N_17495,N_17539);
or U20642 (N_20642,N_15135,N_17929);
and U20643 (N_20643,N_13340,N_16137);
nand U20644 (N_20644,N_13894,N_15155);
or U20645 (N_20645,N_16727,N_15041);
xnor U20646 (N_20646,N_13305,N_13548);
and U20647 (N_20647,N_13973,N_12832);
or U20648 (N_20648,N_16479,N_12697);
or U20649 (N_20649,N_14046,N_18008);
nor U20650 (N_20650,N_13707,N_17384);
and U20651 (N_20651,N_13523,N_12669);
and U20652 (N_20652,N_14238,N_14526);
or U20653 (N_20653,N_17727,N_17345);
xor U20654 (N_20654,N_15209,N_17985);
xor U20655 (N_20655,N_15183,N_16053);
or U20656 (N_20656,N_12798,N_12935);
nand U20657 (N_20657,N_13747,N_18675);
xnor U20658 (N_20658,N_17270,N_18453);
and U20659 (N_20659,N_15964,N_13327);
or U20660 (N_20660,N_12576,N_15784);
nand U20661 (N_20661,N_14453,N_18129);
and U20662 (N_20662,N_15930,N_13162);
and U20663 (N_20663,N_18682,N_12794);
nor U20664 (N_20664,N_13899,N_16241);
nand U20665 (N_20665,N_13778,N_17156);
nor U20666 (N_20666,N_18672,N_16713);
xnor U20667 (N_20667,N_18227,N_15577);
xnor U20668 (N_20668,N_17422,N_14261);
xor U20669 (N_20669,N_17946,N_16653);
nand U20670 (N_20670,N_17584,N_18017);
nor U20671 (N_20671,N_13294,N_14142);
nor U20672 (N_20672,N_17864,N_15369);
xor U20673 (N_20673,N_13413,N_14633);
xnor U20674 (N_20674,N_13882,N_16989);
or U20675 (N_20675,N_13507,N_13317);
xnor U20676 (N_20676,N_15024,N_15220);
nand U20677 (N_20677,N_15771,N_12731);
or U20678 (N_20678,N_14051,N_16978);
nor U20679 (N_20679,N_15811,N_12945);
nor U20680 (N_20680,N_12931,N_13904);
or U20681 (N_20681,N_14195,N_18163);
or U20682 (N_20682,N_14737,N_16604);
nor U20683 (N_20683,N_12753,N_14322);
nor U20684 (N_20684,N_16086,N_13319);
and U20685 (N_20685,N_18657,N_16701);
nand U20686 (N_20686,N_12729,N_15109);
nor U20687 (N_20687,N_18697,N_15581);
nand U20688 (N_20688,N_17083,N_16301);
and U20689 (N_20689,N_17551,N_14257);
and U20690 (N_20690,N_13855,N_16403);
or U20691 (N_20691,N_18383,N_12861);
nor U20692 (N_20692,N_17530,N_14419);
or U20693 (N_20693,N_18376,N_17750);
and U20694 (N_20694,N_16240,N_16114);
xnor U20695 (N_20695,N_18462,N_12791);
xor U20696 (N_20696,N_13055,N_17598);
nand U20697 (N_20697,N_16595,N_17262);
nor U20698 (N_20698,N_16217,N_17909);
or U20699 (N_20699,N_13961,N_15937);
and U20700 (N_20700,N_13563,N_17311);
nor U20701 (N_20701,N_15913,N_12877);
nor U20702 (N_20702,N_15249,N_12620);
xnor U20703 (N_20703,N_14081,N_17787);
and U20704 (N_20704,N_13840,N_12543);
nor U20705 (N_20705,N_15710,N_18302);
nand U20706 (N_20706,N_18110,N_17862);
nand U20707 (N_20707,N_13575,N_17922);
nand U20708 (N_20708,N_15786,N_13949);
nor U20709 (N_20709,N_16764,N_16948);
or U20710 (N_20710,N_16990,N_14096);
xnor U20711 (N_20711,N_12917,N_16171);
nand U20712 (N_20712,N_17333,N_18569);
xor U20713 (N_20713,N_15736,N_18713);
nor U20714 (N_20714,N_14851,N_15703);
and U20715 (N_20715,N_15317,N_16809);
or U20716 (N_20716,N_15830,N_13057);
and U20717 (N_20717,N_16757,N_17073);
or U20718 (N_20718,N_13630,N_15945);
nor U20719 (N_20719,N_16831,N_16666);
nand U20720 (N_20720,N_16702,N_16810);
xnor U20721 (N_20721,N_17848,N_18620);
and U20722 (N_20722,N_16397,N_14017);
xor U20723 (N_20723,N_16626,N_14346);
nand U20724 (N_20724,N_14519,N_12992);
nand U20725 (N_20725,N_16662,N_12973);
and U20726 (N_20726,N_18679,N_13362);
nor U20727 (N_20727,N_15705,N_17433);
nor U20728 (N_20728,N_15065,N_14871);
nor U20729 (N_20729,N_16373,N_17758);
nor U20730 (N_20730,N_12940,N_15473);
nor U20731 (N_20731,N_16878,N_17903);
nor U20732 (N_20732,N_16372,N_14894);
nor U20733 (N_20733,N_18367,N_13624);
nand U20734 (N_20734,N_13301,N_16800);
or U20735 (N_20735,N_17900,N_17901);
xor U20736 (N_20736,N_14082,N_17506);
nor U20737 (N_20737,N_15161,N_15537);
nor U20738 (N_20738,N_13099,N_18049);
xor U20739 (N_20739,N_17891,N_12714);
and U20740 (N_20740,N_16724,N_17819);
xnor U20741 (N_20741,N_16643,N_18556);
or U20742 (N_20742,N_14751,N_16048);
nand U20743 (N_20743,N_18231,N_18104);
nand U20744 (N_20744,N_13702,N_17236);
nand U20745 (N_20745,N_15572,N_14940);
xor U20746 (N_20746,N_13502,N_15719);
nor U20747 (N_20747,N_15310,N_16857);
xor U20748 (N_20748,N_18252,N_14765);
nand U20749 (N_20749,N_16570,N_17135);
nand U20750 (N_20750,N_13967,N_12536);
nand U20751 (N_20751,N_13422,N_16157);
xor U20752 (N_20752,N_13392,N_15613);
xor U20753 (N_20753,N_16649,N_15418);
nand U20754 (N_20754,N_15782,N_14906);
xnor U20755 (N_20755,N_14537,N_16194);
or U20756 (N_20756,N_17851,N_13410);
xor U20757 (N_20757,N_18083,N_15863);
xnor U20758 (N_20758,N_13635,N_13817);
xor U20759 (N_20759,N_16511,N_12542);
nand U20760 (N_20760,N_14066,N_13738);
nor U20761 (N_20761,N_13489,N_12860);
nand U20762 (N_20762,N_14235,N_16654);
xor U20763 (N_20763,N_16167,N_15694);
and U20764 (N_20764,N_12619,N_15515);
or U20765 (N_20765,N_17807,N_18369);
nand U20766 (N_20766,N_14985,N_18066);
nor U20767 (N_20767,N_14338,N_17952);
or U20768 (N_20768,N_13663,N_14273);
xnor U20769 (N_20769,N_17421,N_15652);
nand U20770 (N_20770,N_13586,N_17785);
nor U20771 (N_20771,N_14684,N_15879);
xnor U20772 (N_20772,N_16834,N_18572);
or U20773 (N_20773,N_17936,N_13799);
nand U20774 (N_20774,N_13936,N_13376);
and U20775 (N_20775,N_17755,N_13399);
xnor U20776 (N_20776,N_12990,N_15883);
xnor U20777 (N_20777,N_15775,N_15764);
nor U20778 (N_20778,N_12688,N_13944);
nand U20779 (N_20779,N_15506,N_13221);
or U20780 (N_20780,N_17826,N_13860);
or U20781 (N_20781,N_12919,N_15846);
nor U20782 (N_20782,N_13518,N_14685);
nor U20783 (N_20783,N_12929,N_12793);
nand U20784 (N_20784,N_18078,N_15604);
nor U20785 (N_20785,N_18352,N_15301);
nand U20786 (N_20786,N_14090,N_13926);
xnor U20787 (N_20787,N_17768,N_13334);
nor U20788 (N_20788,N_15336,N_18439);
nor U20789 (N_20789,N_16687,N_17832);
nor U20790 (N_20790,N_17307,N_12704);
nor U20791 (N_20791,N_13348,N_14365);
nor U20792 (N_20792,N_17651,N_16775);
nand U20793 (N_20793,N_15374,N_14420);
nor U20794 (N_20794,N_12944,N_14620);
and U20795 (N_20795,N_14807,N_13002);
xnor U20796 (N_20796,N_18142,N_18305);
nand U20797 (N_20797,N_12533,N_13807);
and U20798 (N_20798,N_14312,N_17759);
xor U20799 (N_20799,N_13883,N_15817);
nand U20800 (N_20800,N_18149,N_12592);
nand U20801 (N_20801,N_14882,N_16592);
and U20802 (N_20802,N_13391,N_18621);
and U20803 (N_20803,N_17532,N_15766);
or U20804 (N_20804,N_13408,N_13264);
nor U20805 (N_20805,N_12762,N_15670);
xor U20806 (N_20806,N_16324,N_17547);
xor U20807 (N_20807,N_16957,N_12924);
nand U20808 (N_20808,N_16637,N_14253);
xor U20809 (N_20809,N_16777,N_13553);
and U20810 (N_20810,N_14716,N_16434);
and U20811 (N_20811,N_14832,N_14604);
xnor U20812 (N_20812,N_13900,N_13424);
nor U20813 (N_20813,N_14567,N_12561);
xor U20814 (N_20814,N_13932,N_13133);
or U20815 (N_20815,N_18576,N_14644);
nor U20816 (N_20816,N_14609,N_14970);
or U20817 (N_20817,N_12915,N_17410);
nor U20818 (N_20818,N_18552,N_13802);
nand U20819 (N_20819,N_14412,N_13212);
nor U20820 (N_20820,N_15734,N_17793);
nor U20821 (N_20821,N_14171,N_16008);
and U20822 (N_20822,N_16327,N_15685);
and U20823 (N_20823,N_12904,N_16984);
nand U20824 (N_20824,N_17611,N_15366);
nor U20825 (N_20825,N_18020,N_16515);
and U20826 (N_20826,N_15965,N_18415);
nand U20827 (N_20827,N_12708,N_17624);
nor U20828 (N_20828,N_18324,N_16506);
nor U20829 (N_20829,N_16543,N_15690);
xnor U20830 (N_20830,N_15540,N_13775);
nand U20831 (N_20831,N_17151,N_13725);
and U20832 (N_20832,N_17077,N_14181);
nor U20833 (N_20833,N_16162,N_13698);
or U20834 (N_20834,N_18220,N_13998);
xor U20835 (N_20835,N_18229,N_16333);
xor U20836 (N_20836,N_14469,N_13532);
nand U20837 (N_20837,N_17161,N_18525);
nor U20838 (N_20838,N_13168,N_14384);
xnor U20839 (N_20839,N_15210,N_13420);
or U20840 (N_20840,N_16933,N_14303);
and U20841 (N_20841,N_12894,N_18248);
nand U20842 (N_20842,N_17351,N_17321);
xor U20843 (N_20843,N_13863,N_18205);
xnor U20844 (N_20844,N_17893,N_15313);
nand U20845 (N_20845,N_13694,N_17594);
and U20846 (N_20846,N_18239,N_16696);
or U20847 (N_20847,N_16191,N_13662);
xor U20848 (N_20848,N_16002,N_14549);
nand U20849 (N_20849,N_18128,N_12870);
nand U20850 (N_20850,N_15403,N_17984);
nor U20851 (N_20851,N_15610,N_16096);
nand U20852 (N_20852,N_17917,N_15459);
xor U20853 (N_20853,N_16538,N_15871);
nor U20854 (N_20854,N_14919,N_18702);
nand U20855 (N_20855,N_13192,N_16883);
or U20856 (N_20856,N_17601,N_12854);
and U20857 (N_20857,N_18723,N_14072);
xnor U20858 (N_20858,N_16707,N_18445);
or U20859 (N_20859,N_15959,N_16297);
nor U20860 (N_20860,N_14356,N_14039);
xnor U20861 (N_20861,N_15357,N_13204);
nor U20862 (N_20862,N_17361,N_17268);
and U20863 (N_20863,N_13813,N_17888);
or U20864 (N_20864,N_18615,N_17885);
xnor U20865 (N_20865,N_17045,N_18459);
nand U20866 (N_20866,N_12523,N_18585);
and U20867 (N_20867,N_13277,N_13336);
nand U20868 (N_20868,N_18671,N_13693);
xnor U20869 (N_20869,N_17214,N_16622);
nand U20870 (N_20870,N_17281,N_18414);
xnor U20871 (N_20871,N_14167,N_16930);
or U20872 (N_20872,N_18088,N_14329);
or U20873 (N_20873,N_17472,N_12664);
nor U20874 (N_20874,N_16436,N_15002);
or U20875 (N_20875,N_17367,N_18708);
and U20876 (N_20876,N_16658,N_15943);
xnor U20877 (N_20877,N_16513,N_13979);
nor U20878 (N_20878,N_17074,N_14330);
or U20879 (N_20879,N_15607,N_16001);
nand U20880 (N_20880,N_15737,N_12733);
nand U20881 (N_20881,N_17559,N_13554);
and U20882 (N_20882,N_15820,N_14048);
xnor U20883 (N_20883,N_14557,N_18484);
nor U20884 (N_20884,N_15101,N_16446);
nand U20885 (N_20885,N_15398,N_16812);
nor U20886 (N_20886,N_16108,N_17786);
nor U20887 (N_20887,N_14701,N_13350);
nand U20888 (N_20888,N_16851,N_14921);
nand U20889 (N_20889,N_18691,N_16567);
and U20890 (N_20890,N_14924,N_16495);
nand U20891 (N_20891,N_14583,N_14531);
and U20892 (N_20892,N_15701,N_17699);
xnor U20893 (N_20893,N_13950,N_15698);
or U20894 (N_20894,N_16916,N_15717);
nor U20895 (N_20895,N_15646,N_13601);
xor U20896 (N_20896,N_17193,N_14194);
nand U20897 (N_20897,N_15047,N_13251);
nand U20898 (N_20898,N_14119,N_17293);
or U20899 (N_20899,N_15671,N_16249);
nand U20900 (N_20900,N_16601,N_15416);
and U20901 (N_20901,N_16671,N_14950);
and U20902 (N_20902,N_17605,N_17480);
or U20903 (N_20903,N_16621,N_17537);
xnor U20904 (N_20904,N_13512,N_17063);
nor U20905 (N_20905,N_15034,N_17857);
or U20906 (N_20906,N_15521,N_14180);
xnor U20907 (N_20907,N_17145,N_12656);
nor U20908 (N_20908,N_13823,N_17934);
nand U20909 (N_20909,N_13022,N_15603);
nor U20910 (N_20910,N_14074,N_18624);
and U20911 (N_20911,N_13719,N_16749);
and U20912 (N_20912,N_14720,N_15947);
and U20913 (N_20913,N_12502,N_18710);
nand U20914 (N_20914,N_13131,N_16806);
or U20915 (N_20915,N_12888,N_16752);
xor U20916 (N_20916,N_17044,N_16161);
or U20917 (N_20917,N_18175,N_17027);
xnor U20918 (N_20918,N_16066,N_12878);
nor U20919 (N_20919,N_12501,N_13298);
or U20920 (N_20920,N_14605,N_14731);
or U20921 (N_20921,N_14282,N_15891);
xnor U20922 (N_20922,N_12943,N_14098);
nor U20923 (N_20923,N_15586,N_13652);
and U20924 (N_20924,N_15167,N_18398);
nor U20925 (N_20925,N_18145,N_13372);
xor U20926 (N_20926,N_15439,N_16747);
xor U20927 (N_20927,N_18584,N_14876);
and U20928 (N_20928,N_18452,N_13897);
nor U20929 (N_20929,N_12962,N_13321);
nand U20930 (N_20930,N_13870,N_15901);
nor U20931 (N_20931,N_18639,N_12712);
or U20932 (N_20932,N_16605,N_18357);
nand U20933 (N_20933,N_15397,N_13178);
nor U20934 (N_20934,N_16289,N_17667);
nor U20935 (N_20935,N_13678,N_17025);
xnor U20936 (N_20936,N_14875,N_13384);
xor U20937 (N_20937,N_17666,N_15513);
and U20938 (N_20938,N_16596,N_16192);
xnor U20939 (N_20939,N_14417,N_15144);
xor U20940 (N_20940,N_14948,N_15816);
nand U20941 (N_20941,N_16716,N_17550);
nand U20942 (N_20942,N_12709,N_17777);
nand U20943 (N_20943,N_15265,N_18399);
xor U20944 (N_20944,N_15655,N_12602);
nor U20945 (N_20945,N_14137,N_12905);
nor U20946 (N_20946,N_16279,N_16302);
nand U20947 (N_20947,N_16225,N_16855);
nor U20948 (N_20948,N_17702,N_13577);
nor U20949 (N_20949,N_18547,N_13310);
or U20950 (N_20950,N_17581,N_17201);
nor U20951 (N_20951,N_16228,N_16866);
xor U20952 (N_20952,N_16838,N_18574);
nand U20953 (N_20953,N_13851,N_15364);
xor U20954 (N_20954,N_17544,N_17347);
xnor U20955 (N_20955,N_16790,N_16376);
nor U20956 (N_20956,N_15267,N_14992);
or U20957 (N_20957,N_16221,N_14001);
or U20958 (N_20958,N_13614,N_16110);
and U20959 (N_20959,N_18282,N_13809);
xnor U20960 (N_20960,N_12882,N_12689);
and U20961 (N_20961,N_13071,N_16762);
nor U20962 (N_20962,N_13653,N_18174);
and U20963 (N_20963,N_18481,N_13188);
xor U20964 (N_20964,N_12603,N_14750);
or U20965 (N_20965,N_16760,N_13682);
or U20966 (N_20966,N_16677,N_14916);
nand U20967 (N_20967,N_16170,N_15177);
xnor U20968 (N_20968,N_16259,N_14613);
or U20969 (N_20969,N_15986,N_12698);
nand U20970 (N_20970,N_18663,N_15962);
nand U20971 (N_20971,N_12970,N_17154);
nand U20972 (N_20972,N_13421,N_12701);
nand U20973 (N_20973,N_16971,N_17136);
nor U20974 (N_20974,N_14162,N_14516);
and U20975 (N_20975,N_16033,N_17737);
and U20976 (N_20976,N_16820,N_18583);
nand U20977 (N_20977,N_12756,N_13326);
nor U20978 (N_20978,N_16608,N_14833);
xnor U20979 (N_20979,N_18717,N_14383);
nand U20980 (N_20980,N_12552,N_17937);
and U20981 (N_20981,N_14109,N_14117);
and U20982 (N_20982,N_13324,N_13280);
nor U20983 (N_20983,N_15032,N_12773);
nor U20984 (N_20984,N_17158,N_15173);
nor U20985 (N_20985,N_13331,N_15325);
or U20986 (N_20986,N_16151,N_16758);
or U20987 (N_20987,N_17784,N_17402);
nor U20988 (N_20988,N_17896,N_17447);
nand U20989 (N_20989,N_18643,N_16412);
or U20990 (N_20990,N_17406,N_13989);
or U20991 (N_20991,N_18613,N_13233);
nand U20992 (N_20992,N_16472,N_16746);
and U20993 (N_20993,N_15126,N_17497);
xnor U20994 (N_20994,N_14705,N_15718);
and U20995 (N_20995,N_13208,N_18749);
or U20996 (N_20996,N_12823,N_18291);
xnor U20997 (N_20997,N_17336,N_12758);
and U20998 (N_20998,N_15241,N_18648);
and U20999 (N_20999,N_17160,N_13737);
xnor U21000 (N_21000,N_12790,N_17283);
nand U21001 (N_21001,N_14913,N_17298);
and U21002 (N_21002,N_14367,N_18265);
nor U21003 (N_21003,N_17887,N_18043);
nand U21004 (N_21004,N_17669,N_18482);
nand U21005 (N_21005,N_15785,N_18328);
xnor U21006 (N_21006,N_12783,N_16856);
xnor U21007 (N_21007,N_13001,N_17470);
xnor U21008 (N_21008,N_17626,N_15353);
nand U21009 (N_21009,N_15186,N_16722);
nor U21010 (N_21010,N_16730,N_16753);
and U21011 (N_21011,N_17168,N_17327);
nor U21012 (N_21012,N_13583,N_15021);
xnor U21013 (N_21013,N_15721,N_12643);
nor U21014 (N_21014,N_16768,N_17119);
or U21015 (N_21015,N_18125,N_14776);
nand U21016 (N_21016,N_17494,N_18653);
or U21017 (N_21017,N_13843,N_15608);
and U21018 (N_21018,N_18014,N_17215);
nand U21019 (N_21019,N_13087,N_15337);
xnor U21020 (N_21020,N_14242,N_17369);
nand U21021 (N_21021,N_13673,N_17804);
xor U21022 (N_21022,N_15984,N_12869);
nor U21023 (N_21023,N_15482,N_14911);
nand U21024 (N_21024,N_16003,N_17061);
xor U21025 (N_21025,N_13526,N_15770);
or U21026 (N_21026,N_14617,N_15227);
nand U21027 (N_21027,N_16611,N_14951);
and U21028 (N_21028,N_16684,N_12969);
and U21029 (N_21029,N_16669,N_18578);
nor U21030 (N_21030,N_14343,N_18510);
xor U21031 (N_21031,N_13529,N_17457);
and U21032 (N_21032,N_13339,N_16042);
xor U21033 (N_21033,N_13126,N_18184);
nand U21034 (N_21034,N_18534,N_17943);
nor U21035 (N_21035,N_17282,N_14648);
nand U21036 (N_21036,N_15570,N_17742);
xor U21037 (N_21037,N_18638,N_16142);
nand U21038 (N_21038,N_18678,N_15929);
and U21039 (N_21039,N_17682,N_17241);
or U21040 (N_21040,N_17628,N_17676);
nand U21041 (N_21041,N_18580,N_14854);
nor U21042 (N_21042,N_16655,N_18076);
or U21043 (N_21043,N_15089,N_15009);
nor U21044 (N_21044,N_18652,N_17448);
nor U21045 (N_21045,N_16699,N_14930);
nor U21046 (N_21046,N_17068,N_17854);
nand U21047 (N_21047,N_17324,N_18138);
and U21048 (N_21048,N_13709,N_17251);
xnor U21049 (N_21049,N_18448,N_17205);
nand U21050 (N_21050,N_17374,N_12946);
xnor U21051 (N_21051,N_12772,N_15553);
nand U21052 (N_21052,N_14881,N_16482);
or U21053 (N_21053,N_13352,N_13645);
nor U21054 (N_21054,N_16463,N_18029);
or U21055 (N_21055,N_17806,N_15749);
nor U21056 (N_21056,N_16304,N_17585);
nor U21057 (N_21057,N_12930,N_13641);
xor U21058 (N_21058,N_15768,N_18037);
and U21059 (N_21059,N_13263,N_16154);
nand U21060 (N_21060,N_17780,N_18256);
xor U21061 (N_21061,N_13567,N_15345);
nand U21062 (N_21062,N_14040,N_15856);
xor U21063 (N_21063,N_13510,N_15125);
and U21064 (N_21064,N_14971,N_18377);
nor U21065 (N_21065,N_14873,N_12872);
nor U21066 (N_21066,N_14150,N_18237);
xnor U21067 (N_21067,N_15107,N_17637);
nand U21068 (N_21068,N_13116,N_17350);
nand U21069 (N_21069,N_15848,N_18046);
xor U21070 (N_21070,N_16842,N_15279);
nand U21071 (N_21071,N_14818,N_18565);
nand U21072 (N_21072,N_13461,N_16355);
nand U21073 (N_21073,N_13401,N_15733);
or U21074 (N_21074,N_14957,N_15842);
or U21075 (N_21075,N_13454,N_18350);
xor U21076 (N_21076,N_13861,N_17956);
or U21077 (N_21077,N_17163,N_17228);
or U21078 (N_21078,N_12675,N_13792);
or U21079 (N_21079,N_18216,N_18114);
or U21080 (N_21080,N_15184,N_17795);
nor U21081 (N_21081,N_16950,N_18015);
nor U21082 (N_21082,N_16400,N_17141);
nor U21083 (N_21083,N_18441,N_14103);
nand U21084 (N_21084,N_18274,N_14287);
and U21085 (N_21085,N_18278,N_16636);
nand U21086 (N_21086,N_15284,N_14850);
nor U21087 (N_21087,N_17717,N_16973);
nor U21088 (N_21088,N_13909,N_16723);
and U21089 (N_21089,N_14941,N_18637);
nor U21090 (N_21090,N_14019,N_18258);
or U21091 (N_21091,N_13478,N_13539);
nand U21092 (N_21092,N_17824,N_18011);
xnor U21093 (N_21093,N_15944,N_12699);
nor U21094 (N_21094,N_16799,N_17620);
nor U21095 (N_21095,N_17582,N_15291);
and U21096 (N_21096,N_14959,N_16780);
nor U21097 (N_21097,N_15806,N_17054);
xnor U21098 (N_21098,N_12995,N_16040);
nand U21099 (N_21099,N_18097,N_12577);
nor U21100 (N_21100,N_17033,N_13397);
nor U21101 (N_21101,N_15333,N_13119);
xnor U21102 (N_21102,N_12955,N_15309);
nor U21103 (N_21103,N_18725,N_17058);
nor U21104 (N_21104,N_12746,N_14803);
nor U21105 (N_21105,N_18261,N_17596);
nor U21106 (N_21106,N_15805,N_17867);
nor U21107 (N_21107,N_17445,N_14592);
nor U21108 (N_21108,N_18524,N_13223);
nor U21109 (N_21109,N_13047,N_15199);
or U21110 (N_21110,N_16396,N_15789);
nand U21111 (N_21111,N_14667,N_17100);
and U21112 (N_21112,N_18490,N_17965);
xnor U21113 (N_21113,N_16697,N_16537);
xnor U21114 (N_21114,N_15426,N_16464);
and U21115 (N_21115,N_16362,N_17916);
nor U21116 (N_21116,N_16049,N_14071);
nand U21117 (N_21117,N_17892,N_18283);
and U21118 (N_21118,N_17398,N_18736);
nand U21119 (N_21119,N_13800,N_16840);
nand U21120 (N_21120,N_13848,N_13037);
nor U21121 (N_21121,N_13689,N_15629);
nor U21122 (N_21122,N_18249,N_17391);
nor U21123 (N_21123,N_13845,N_18228);
nand U21124 (N_21124,N_17510,N_15835);
or U21125 (N_21125,N_15408,N_15257);
nand U21126 (N_21126,N_14689,N_13303);
or U21127 (N_21127,N_13602,N_12880);
and U21128 (N_21128,N_18536,N_15392);
xor U21129 (N_21129,N_12830,N_13962);
nand U21130 (N_21130,N_13929,N_13247);
nor U21131 (N_21131,N_15667,N_17378);
nand U21132 (N_21132,N_12503,N_17308);
and U21133 (N_21133,N_12927,N_14634);
xor U21134 (N_21134,N_12663,N_13094);
nand U21135 (N_21135,N_14542,N_15169);
nor U21136 (N_21136,N_13115,N_13062);
and U21137 (N_21137,N_17765,N_14926);
xnor U21138 (N_21138,N_17102,N_13242);
and U21139 (N_21139,N_15117,N_16801);
nand U21140 (N_21140,N_13671,N_17691);
or U21141 (N_21141,N_14024,N_18397);
or U21142 (N_21142,N_16456,N_13488);
xnor U21143 (N_21143,N_14289,N_14288);
xnor U21144 (N_21144,N_18676,N_18235);
xnor U21145 (N_21145,N_13743,N_18515);
or U21146 (N_21146,N_15576,N_17456);
or U21147 (N_21147,N_16598,N_13430);
nand U21148 (N_21148,N_14267,N_16629);
nor U21149 (N_21149,N_13760,N_13370);
xor U21150 (N_21150,N_16976,N_15185);
nand U21151 (N_21151,N_16390,N_16335);
or U21152 (N_21152,N_18334,N_14893);
or U21153 (N_21153,N_13513,N_16938);
nor U21154 (N_21154,N_18023,N_18387);
xor U21155 (N_21155,N_15295,N_15825);
nand U21156 (N_21156,N_16323,N_13975);
nor U21157 (N_21157,N_15218,N_13795);
or U21158 (N_21158,N_17573,N_16296);
xor U21159 (N_21159,N_15554,N_18219);
nor U21160 (N_21160,N_13293,N_17383);
nor U21161 (N_21161,N_17776,N_15678);
nor U21162 (N_21162,N_14402,N_18344);
nand U21163 (N_21163,N_16287,N_13835);
xor U21164 (N_21164,N_12693,N_13176);
and U21165 (N_21165,N_14089,N_17963);
nor U21166 (N_21166,N_14756,N_15464);
or U21167 (N_21167,N_15951,N_16520);
nand U21168 (N_21168,N_15138,N_14073);
xnor U21169 (N_21169,N_13616,N_13685);
nor U21170 (N_21170,N_13108,N_15741);
nor U21171 (N_21171,N_16548,N_13520);
or U21172 (N_21172,N_13741,N_14000);
and U21173 (N_21173,N_16661,N_13322);
and U21174 (N_21174,N_14666,N_15206);
and U21175 (N_21175,N_14628,N_16731);
or U21176 (N_21176,N_16139,N_17358);
nor U21177 (N_21177,N_16992,N_12569);
and U21178 (N_21178,N_16845,N_14890);
nor U21179 (N_21179,N_16924,N_15908);
xnor U21180 (N_21180,N_18172,N_12792);
nand U21181 (N_21181,N_18311,N_15860);
xor U21182 (N_21182,N_14313,N_17196);
or U21183 (N_21183,N_12721,N_15481);
or U21184 (N_21184,N_16573,N_16361);
nor U21185 (N_21185,N_12586,N_15058);
xor U21186 (N_21186,N_13258,N_15052);
nor U21187 (N_21187,N_15390,N_12724);
xnor U21188 (N_21188,N_15828,N_17519);
nand U21189 (N_21189,N_14404,N_13856);
and U21190 (N_21190,N_13572,N_12515);
nand U21191 (N_21191,N_13672,N_13587);
and U21192 (N_21192,N_14063,N_14293);
nand U21193 (N_21193,N_16431,N_15813);
xnor U21194 (N_21194,N_13285,N_17066);
and U21195 (N_21195,N_15202,N_15436);
nor U21196 (N_21196,N_17955,N_15417);
nor U21197 (N_21197,N_16214,N_18290);
xor U21198 (N_21198,N_12782,N_14337);
xor U21199 (N_21199,N_14812,N_16233);
or U21200 (N_21200,N_17302,N_13302);
xor U21201 (N_21201,N_15303,N_14758);
and U21202 (N_21202,N_13749,N_16597);
nand U21203 (N_21203,N_15574,N_14861);
and U21204 (N_21204,N_16647,N_14141);
nor U21205 (N_21205,N_14428,N_15243);
xnor U21206 (N_21206,N_13984,N_17164);
xor U21207 (N_21207,N_14225,N_13046);
nand U21208 (N_21208,N_13858,N_16875);
or U21209 (N_21209,N_16558,N_13300);
nand U21210 (N_21210,N_14248,N_14114);
or U21211 (N_21211,N_13286,N_17545);
or U21212 (N_21212,N_16461,N_15119);
or U21213 (N_21213,N_16536,N_15349);
xor U21214 (N_21214,N_16615,N_14558);
xor U21215 (N_21215,N_18255,N_16745);
nor U21216 (N_21216,N_13928,N_13147);
nor U21217 (N_21217,N_15405,N_14408);
and U21218 (N_21218,N_15665,N_13124);
or U21219 (N_21219,N_12926,N_17007);
nand U21220 (N_21220,N_16737,N_15739);
nand U21221 (N_21221,N_14856,N_17843);
xor U21222 (N_21222,N_16638,N_12900);
nand U21223 (N_21223,N_14227,N_15664);
nand U21224 (N_21224,N_17933,N_13811);
and U21225 (N_21225,N_16283,N_18226);
or U21226 (N_21226,N_14879,N_18242);
or U21227 (N_21227,N_15989,N_13343);
nand U21228 (N_21228,N_18612,N_13797);
nor U21229 (N_21229,N_13194,N_17407);
or U21230 (N_21230,N_16406,N_14372);
xor U21231 (N_21231,N_14928,N_17500);
and U21232 (N_21232,N_16181,N_16552);
nor U21233 (N_21233,N_13905,N_15557);
or U21234 (N_21234,N_15758,N_14185);
and U21235 (N_21235,N_17574,N_14396);
or U21236 (N_21236,N_17741,N_12817);
or U21237 (N_21237,N_15531,N_16371);
nor U21238 (N_21238,N_15449,N_14863);
xnor U21239 (N_21239,N_16965,N_17451);
or U21240 (N_21240,N_12725,N_14292);
nand U21241 (N_21241,N_17800,N_14336);
xnor U21242 (N_21242,N_13557,N_12996);
and U21243 (N_21243,N_14938,N_18604);
or U21244 (N_21244,N_17176,N_14942);
nor U21245 (N_21245,N_14076,N_14028);
and U21246 (N_21246,N_17496,N_16546);
and U21247 (N_21247,N_15221,N_18410);
or U21248 (N_21248,N_18026,N_16006);
nand U21249 (N_21249,N_13155,N_16252);
nand U21250 (N_21250,N_15998,N_17949);
or U21251 (N_21251,N_15963,N_18390);
nand U21252 (N_21252,N_15388,N_13097);
nor U21253 (N_21253,N_12720,N_16583);
xnor U21254 (N_21254,N_14314,N_18307);
nand U21255 (N_21255,N_14802,N_16429);
nand U21256 (N_21256,N_14521,N_14966);
nand U21257 (N_21257,N_14755,N_17712);
xor U21258 (N_21258,N_16704,N_17429);
nand U21259 (N_21259,N_14176,N_16120);
nor U21260 (N_21260,N_17207,N_15412);
nor U21261 (N_21261,N_15985,N_12804);
xor U21262 (N_21262,N_18403,N_15502);
or U21263 (N_21263,N_13997,N_13810);
xnor U21264 (N_21264,N_14539,N_16271);
nand U21265 (N_21265,N_13052,N_18483);
nand U21266 (N_21266,N_15092,N_15640);
xor U21267 (N_21267,N_14773,N_16234);
nand U21268 (N_21268,N_16368,N_15318);
or U21269 (N_21269,N_16345,N_17038);
nand U21270 (N_21270,N_16025,N_18733);
nand U21271 (N_21271,N_18738,N_18380);
nor U21272 (N_21272,N_12849,N_18590);
xor U21273 (N_21273,N_16904,N_12529);
or U21274 (N_21274,N_13284,N_12650);
nand U21275 (N_21275,N_17568,N_13005);
nor U21276 (N_21276,N_18025,N_18317);
or U21277 (N_21277,N_18225,N_17595);
and U21278 (N_21278,N_13486,N_15314);
nor U21279 (N_21279,N_17403,N_18280);
or U21280 (N_21280,N_16892,N_15899);
or U21281 (N_21281,N_13903,N_13659);
and U21282 (N_21282,N_14277,N_16280);
xor U21283 (N_21283,N_17491,N_14547);
and U21284 (N_21284,N_18325,N_13605);
nor U21285 (N_21285,N_14433,N_17313);
nand U21286 (N_21286,N_18034,N_15137);
nand U21287 (N_21287,N_17541,N_14290);
nand U21288 (N_21288,N_16445,N_13717);
nor U21289 (N_21289,N_13019,N_14186);
nor U21290 (N_21290,N_12700,N_13733);
and U21291 (N_21291,N_13323,N_12781);
or U21292 (N_21292,N_13814,N_12671);
nor U21293 (N_21293,N_17586,N_12755);
or U21294 (N_21294,N_15632,N_14472);
nand U21295 (N_21295,N_13584,N_13471);
nand U21296 (N_21296,N_13839,N_18222);
and U21297 (N_21297,N_17677,N_17612);
and U21298 (N_21298,N_12678,N_15662);
nor U21299 (N_21299,N_14813,N_16927);
and U21300 (N_21300,N_13275,N_18418);
nand U21301 (N_21301,N_16164,N_17625);
and U21302 (N_21302,N_17416,N_15091);
xor U21303 (N_21303,N_13184,N_15738);
and U21304 (N_21304,N_18555,N_12795);
and U21305 (N_21305,N_18124,N_15251);
nor U21306 (N_21306,N_13901,N_12826);
xor U21307 (N_21307,N_14494,N_14306);
xor U21308 (N_21308,N_16358,N_12715);
nand U21309 (N_21309,N_12584,N_18492);
xnor U21310 (N_21310,N_18047,N_17131);
or U21311 (N_21311,N_12661,N_16586);
or U21312 (N_21312,N_15450,N_17511);
xnor U21313 (N_21313,N_16097,N_16399);
nor U21314 (N_21314,N_15084,N_15628);
nor U21315 (N_21315,N_12660,N_14639);
or U21316 (N_21316,N_14779,N_18099);
or U21317 (N_21317,N_15338,N_12568);
and U21318 (N_21318,N_13786,N_13637);
and U21319 (N_21319,N_12707,N_15889);
nand U21320 (N_21320,N_14662,N_15709);
nand U21321 (N_21321,N_14783,N_15714);
nand U21322 (N_21322,N_18673,N_15063);
and U21323 (N_21323,N_17028,N_15296);
xor U21324 (N_21324,N_18742,N_17086);
or U21325 (N_21325,N_13805,N_17354);
nand U21326 (N_21326,N_15377,N_17868);
nand U21327 (N_21327,N_18314,N_17242);
xor U21328 (N_21328,N_14972,N_17489);
xnor U21329 (N_21329,N_16874,N_16073);
nor U21330 (N_21330,N_14686,N_13729);
xor U21331 (N_21331,N_13632,N_15026);
or U21332 (N_21332,N_14507,N_17609);
nor U21333 (N_21333,N_13012,N_16670);
and U21334 (N_21334,N_16589,N_13111);
nand U21335 (N_21335,N_17614,N_15857);
or U21336 (N_21336,N_18688,N_14914);
or U21337 (N_21337,N_13965,N_13907);
nand U21338 (N_21338,N_14898,N_12818);
or U21339 (N_21339,N_15839,N_18016);
nand U21340 (N_21340,N_16710,N_16351);
xor U21341 (N_21341,N_13308,N_13890);
xnor U21342 (N_21342,N_18019,N_17023);
xnor U21343 (N_21343,N_14885,N_16465);
nor U21344 (N_21344,N_15568,N_17672);
nor U21345 (N_21345,N_18353,N_13681);
and U21346 (N_21346,N_15262,N_15207);
and U21347 (N_21347,N_12579,N_13013);
xnor U21348 (N_21348,N_17805,N_18545);
or U21349 (N_21349,N_16656,N_16628);
and U21350 (N_21350,N_17561,N_17189);
xnor U21351 (N_21351,N_13014,N_17430);
or U21352 (N_21352,N_18135,N_16911);
nand U21353 (N_21353,N_17039,N_17477);
and U21354 (N_21354,N_13912,N_16846);
nand U21355 (N_21355,N_17575,N_12934);
or U21356 (N_21356,N_18322,N_15164);
and U21357 (N_21357,N_15096,N_13772);
or U21358 (N_21358,N_16844,N_14056);
or U21359 (N_21359,N_17563,N_16510);
nor U21360 (N_21360,N_17604,N_16276);
nor U21361 (N_21361,N_14077,N_16501);
or U21362 (N_21362,N_15533,N_17797);
nor U21363 (N_21363,N_18595,N_12622);
or U21364 (N_21364,N_13075,N_16902);
and U21365 (N_21365,N_15991,N_18618);
nand U21366 (N_21366,N_15974,N_17761);
or U21367 (N_21367,N_13402,N_16000);
and U21368 (N_21368,N_14627,N_16250);
nand U21369 (N_21369,N_14514,N_17983);
or U21370 (N_21370,N_17540,N_13469);
or U21371 (N_21371,N_15977,N_15873);
nand U21372 (N_21372,N_15140,N_18447);
xor U21373 (N_21373,N_15468,N_15467);
nand U21374 (N_21374,N_17680,N_14886);
nor U21375 (N_21375,N_14714,N_17010);
nand U21376 (N_21376,N_18118,N_16432);
or U21377 (N_21377,N_14823,N_13974);
nand U21378 (N_21378,N_17263,N_18684);
nand U21379 (N_21379,N_14454,N_17405);
and U21380 (N_21380,N_13083,N_16525);
or U21381 (N_21381,N_16816,N_17437);
nor U21382 (N_21382,N_14825,N_18032);
nor U21383 (N_21383,N_12506,N_14541);
xor U21384 (N_21384,N_13571,N_16500);
nor U21385 (N_21385,N_15529,N_18275);
nand U21386 (N_21386,N_13276,N_14215);
nand U21387 (N_21387,N_15645,N_16316);
or U21388 (N_21388,N_18360,N_15706);
nand U21389 (N_21389,N_18656,N_16229);
nor U21390 (N_21390,N_18207,N_18181);
and U21391 (N_21391,N_16833,N_12606);
xnor U21392 (N_21392,N_17814,N_18177);
or U21393 (N_21393,N_16439,N_18230);
xor U21394 (N_21394,N_13688,N_16286);
nor U21395 (N_21395,N_14152,N_15994);
or U21396 (N_21396,N_13156,N_15437);
nor U21397 (N_21397,N_14511,N_12853);
xnor U21398 (N_21398,N_13533,N_18189);
xnor U21399 (N_21399,N_12834,N_13344);
xor U21400 (N_21400,N_16632,N_13739);
or U21401 (N_21401,N_15308,N_18143);
nor U21402 (N_21402,N_17940,N_17087);
or U21403 (N_21403,N_16533,N_17148);
or U21404 (N_21404,N_17538,N_13226);
and U21405 (N_21405,N_16619,N_14456);
xor U21406 (N_21406,N_13257,N_18053);
nor U21407 (N_21407,N_12629,N_13265);
nor U21408 (N_21408,N_15160,N_18644);
and U21409 (N_21409,N_15724,N_17619);
nor U21410 (N_21410,N_14360,N_16783);
or U21411 (N_21411,N_16672,N_13100);
nand U21412 (N_21412,N_17505,N_18611);
and U21413 (N_21413,N_17006,N_14621);
and U21414 (N_21414,N_14625,N_15203);
nand U21415 (N_21415,N_14988,N_15969);
xnor U21416 (N_21416,N_13113,N_15560);
or U21417 (N_21417,N_18206,N_15407);
nand U21418 (N_21418,N_12988,N_18154);
xor U21419 (N_21419,N_15271,N_15402);
nor U21420 (N_21420,N_17760,N_16017);
and U21421 (N_21421,N_17217,N_16043);
and U21422 (N_21422,N_16230,N_14584);
nand U21423 (N_21423,N_12949,N_13534);
and U21424 (N_21424,N_15478,N_15941);
xor U21425 (N_21425,N_18301,N_17109);
nor U21426 (N_21426,N_17812,N_18559);
and U21427 (N_21427,N_17622,N_13918);
nand U21428 (N_21428,N_18488,N_17663);
and U21429 (N_21429,N_14097,N_16420);
or U21430 (N_21430,N_15501,N_13978);
or U21431 (N_21431,N_17646,N_18527);
xor U21432 (N_21432,N_16215,N_14371);
nand U21433 (N_21433,N_14637,N_16491);
nand U21434 (N_21434,N_12964,N_16736);
and U21435 (N_21435,N_13146,N_12875);
or U21436 (N_21436,N_15170,N_16341);
nand U21437 (N_21437,N_14997,N_16061);
xnor U21438 (N_21438,N_14530,N_17941);
or U21439 (N_21439,N_12599,N_14887);
or U21440 (N_21440,N_14432,N_17593);
and U21441 (N_21441,N_18735,N_17583);
nor U21442 (N_21442,N_17419,N_17608);
nand U21443 (N_21443,N_18075,N_16427);
nor U21444 (N_21444,N_14799,N_16402);
nor U21445 (N_21445,N_16152,N_16791);
nand U21446 (N_21446,N_12846,N_14636);
nand U21447 (N_21447,N_16776,N_18067);
or U21448 (N_21448,N_17592,N_16880);
nand U21449 (N_21449,N_14578,N_15781);
nor U21450 (N_21450,N_16453,N_13008);
and U21451 (N_21451,N_14398,N_14679);
nor U21452 (N_21452,N_13481,N_15615);
or U21453 (N_21453,N_15060,N_16518);
and U21454 (N_21454,N_17464,N_17386);
and U21455 (N_21455,N_18409,N_15968);
or U21456 (N_21456,N_15704,N_13088);
xor U21457 (N_21457,N_15446,N_12887);
xor U21458 (N_21458,N_13006,N_16897);
and U21459 (N_21459,N_14153,N_15520);
and U21460 (N_21460,N_14455,N_16425);
or U21461 (N_21461,N_15799,N_16141);
nor U21462 (N_21462,N_16792,N_15268);
and U21463 (N_21463,N_18706,N_13089);
and U21464 (N_21464,N_16458,N_17334);
nand U21465 (N_21465,N_13187,N_17003);
and U21466 (N_21466,N_12966,N_17987);
nor U21467 (N_21467,N_14373,N_15306);
or U21468 (N_21468,N_17284,N_17710);
nor U21469 (N_21469,N_15503,N_18577);
or U21470 (N_21470,N_15139,N_16998);
or U21471 (N_21471,N_16291,N_14723);
and U21472 (N_21472,N_17725,N_14258);
nand U21473 (N_21473,N_18636,N_16451);
nor U21474 (N_21474,N_17905,N_13995);
nor U21475 (N_21475,N_13366,N_13611);
and U21476 (N_21476,N_15419,N_15512);
xor U21477 (N_21477,N_17644,N_14201);
nand U21478 (N_21478,N_16694,N_15853);
xor U21479 (N_21479,N_15571,N_15373);
or U21480 (N_21480,N_15498,N_13677);
or U21481 (N_21481,N_18571,N_12841);
or U21482 (N_21482,N_13359,N_16440);
xor U21483 (N_21483,N_14899,N_14619);
nor U21484 (N_21484,N_18705,N_17638);
nand U21485 (N_21485,N_16734,N_15597);
and U21486 (N_21486,N_16340,N_15551);
nand U21487 (N_21487,N_17675,N_14676);
and U21488 (N_21488,N_17882,N_13462);
nand U21489 (N_21489,N_17958,N_17478);
nor U21490 (N_21490,N_12634,N_17986);
nand U21491 (N_21491,N_13432,N_17287);
or U21492 (N_21492,N_17275,N_15385);
and U21493 (N_21493,N_18479,N_16544);
or U21494 (N_21494,N_13021,N_18010);
nor U21495 (N_21495,N_14925,N_14426);
xnor U21496 (N_21496,N_18234,N_18268);
nand U21497 (N_21497,N_16401,N_16081);
xor U21498 (N_21498,N_14104,N_17813);
and U21499 (N_21499,N_16923,N_18746);
nand U21500 (N_21500,N_16639,N_14155);
xnor U21501 (N_21501,N_13987,N_17803);
and U21502 (N_21502,N_15067,N_15250);
or U21503 (N_21503,N_15180,N_16219);
xor U21504 (N_21504,N_14029,N_18340);
and U21505 (N_21505,N_17684,N_17791);
and U21506 (N_21506,N_13445,N_18042);
nor U21507 (N_21507,N_16065,N_16528);
xnor U21508 (N_21508,N_13033,N_16236);
nor U21509 (N_21509,N_17244,N_14574);
or U21510 (N_21510,N_15152,N_12726);
nor U21511 (N_21511,N_17371,N_15444);
and U21512 (N_21512,N_14088,N_14403);
xor U21513 (N_21513,N_14347,N_17662);
xor U21514 (N_21514,N_13382,N_12921);
xor U21515 (N_21515,N_13064,N_12601);
or U21516 (N_21516,N_14442,N_15988);
nand U21517 (N_21517,N_16165,N_12638);
nand U21518 (N_21518,N_14872,N_16209);
nor U21519 (N_21519,N_18120,N_18381);
nor U21520 (N_21520,N_14586,N_15750);
xnor U21521 (N_21521,N_16600,N_14690);
nor U21522 (N_21522,N_15982,N_17465);
xnor U21523 (N_21523,N_12827,N_16353);
nor U21524 (N_21524,N_14917,N_13207);
or U21525 (N_21525,N_15861,N_17959);
nor U21526 (N_21526,N_12903,N_17459);
and U21527 (N_21527,N_13318,N_16248);
nor U21528 (N_21528,N_14944,N_15933);
and U21529 (N_21529,N_13181,N_13657);
nor U21530 (N_21530,N_17945,N_15776);
nand U21531 (N_21531,N_17210,N_14837);
nor U21532 (N_21532,N_15039,N_16693);
nor U21533 (N_21533,N_17230,N_17565);
nand U21534 (N_21534,N_16421,N_17704);
xor U21535 (N_21535,N_18183,N_13423);
xor U21536 (N_21536,N_15754,N_13463);
nor U21537 (N_21537,N_14174,N_13312);
xor U21538 (N_21538,N_15874,N_13938);
or U21539 (N_21539,N_18477,N_14698);
xnor U21540 (N_21540,N_12705,N_16256);
nor U21541 (N_21541,N_17513,N_12749);
or U21542 (N_21542,N_13159,N_12865);
xor U21543 (N_21543,N_16285,N_17613);
nor U21544 (N_21544,N_14508,N_17392);
nor U21545 (N_21545,N_13172,N_16263);
and U21546 (N_21546,N_13501,N_15297);
nor U21547 (N_21547,N_18434,N_16843);
and U21548 (N_21548,N_14363,N_13914);
and U21549 (N_21549,N_17380,N_16850);
xor U21550 (N_21550,N_12594,N_13538);
or U21551 (N_21551,N_16975,N_14202);
nand U21552 (N_21552,N_14377,N_18440);
or U21553 (N_21553,N_15971,N_16032);
nor U21554 (N_21554,N_16901,N_16550);
nor U21555 (N_21555,N_16116,N_13196);
or U21556 (N_21556,N_14320,N_13067);
nor U21557 (N_21557,N_17747,N_14354);
or U21558 (N_21558,N_14996,N_17246);
xnor U21559 (N_21559,N_17873,N_16423);
xnor U21560 (N_21560,N_14638,N_16562);
or U21561 (N_21561,N_14520,N_13972);
nor U21562 (N_21562,N_17871,N_15239);
or U21563 (N_21563,N_18421,N_17014);
xor U21564 (N_21564,N_16914,N_17842);
and U21565 (N_21565,N_14463,N_14026);
xor U21566 (N_21566,N_13110,N_17703);
xnor U21567 (N_21567,N_15676,N_16912);
xor U21568 (N_21568,N_18699,N_15702);
nand U21569 (N_21569,N_18126,N_13661);
xor U21570 (N_21570,N_17404,N_18712);
nor U21571 (N_21571,N_15300,N_15484);
xor U21572 (N_21572,N_15131,N_16956);
or U21573 (N_21573,N_14905,N_14569);
or U21574 (N_21574,N_17431,N_18293);
and U21575 (N_21575,N_13316,N_13609);
nor U21576 (N_21576,N_15068,N_14364);
nor U21577 (N_21577,N_17142,N_15093);
xor U21578 (N_21578,N_13744,N_15812);
and U21579 (N_21579,N_14496,N_14151);
and U21580 (N_21580,N_15728,N_12863);
nor U21581 (N_21581,N_13556,N_14169);
and U21582 (N_21582,N_14529,N_16100);
xor U21583 (N_21583,N_14436,N_14385);
or U21584 (N_21584,N_17799,N_14782);
or U21585 (N_21585,N_16966,N_12911);
nor U21586 (N_21586,N_12570,N_17111);
nand U21587 (N_21587,N_14002,N_14390);
nand U21588 (N_21588,N_13724,N_17866);
or U21589 (N_21589,N_17138,N_17673);
or U21590 (N_21590,N_13543,N_14434);
nand U21591 (N_21591,N_17860,N_18600);
and U21592 (N_21592,N_12642,N_14123);
or U21593 (N_21593,N_17120,N_17348);
xnor U21594 (N_21594,N_18724,N_13030);
xnor U21595 (N_21595,N_14722,N_12897);
xnor U21596 (N_21596,N_14582,N_17816);
nor U21597 (N_21597,N_15141,N_16135);
or U21598 (N_21598,N_18331,N_17279);
and U21599 (N_21599,N_15821,N_14543);
xor U21600 (N_21600,N_14495,N_16410);
and U21601 (N_21601,N_15808,N_12674);
and U21602 (N_21602,N_15305,N_15682);
and U21603 (N_21603,N_17051,N_17877);
and U21604 (N_21604,N_16036,N_14108);
or U21605 (N_21605,N_17481,N_16344);
and U21606 (N_21606,N_15549,N_15073);
xnor U21607 (N_21607,N_12509,N_16430);
xnor U21608 (N_21608,N_16616,N_12759);
nor U21609 (N_21609,N_18493,N_14647);
xnor U21610 (N_21610,N_13000,N_15123);
and U21611 (N_21611,N_13750,N_17400);
nor U21612 (N_21612,N_12658,N_15315);
nand U21613 (N_21613,N_16352,N_14826);
nand U21614 (N_21614,N_13787,N_14784);
or U21615 (N_21615,N_18098,N_14908);
xor U21616 (N_21616,N_14154,N_15783);
xor U21617 (N_21617,N_16623,N_13514);
and U21618 (N_21618,N_15328,N_13552);
or U21619 (N_21619,N_17265,N_14101);
and U21620 (N_21620,N_14067,N_15762);
nand U21621 (N_21621,N_16330,N_16818);
nand U21622 (N_21622,N_12754,N_13447);
nand U21623 (N_21623,N_17723,N_14431);
nor U21624 (N_21624,N_14474,N_17021);
or U21625 (N_21625,N_14960,N_14254);
nor U21626 (N_21626,N_17911,N_18627);
nor U21627 (N_21627,N_17115,N_14789);
or U21628 (N_21628,N_13762,N_14694);
and U21629 (N_21629,N_14418,N_13946);
nor U21630 (N_21630,N_12681,N_14492);
nor U21631 (N_21631,N_12890,N_17084);
nand U21632 (N_21632,N_13451,N_13329);
xor U21633 (N_21633,N_18361,N_13812);
nand U21634 (N_21634,N_16678,N_16489);
nor U21635 (N_21635,N_15062,N_14559);
xnor U21636 (N_21636,N_17726,N_16708);
or U21637 (N_21637,N_15288,N_15525);
and U21638 (N_21638,N_14214,N_14054);
or U21639 (N_21639,N_14443,N_18491);
nor U21640 (N_21640,N_18065,N_15365);
xnor U21641 (N_21641,N_16174,N_15765);
and U21642 (N_21642,N_16480,N_16055);
or U21643 (N_21643,N_12672,N_15371);
nand U21644 (N_21644,N_14369,N_15381);
nand U21645 (N_21645,N_16645,N_14361);
and U21646 (N_21646,N_14034,N_17204);
nor U21647 (N_21647,N_13846,N_18215);
and U21648 (N_21648,N_13647,N_13260);
or U21649 (N_21649,N_14538,N_13457);
nor U21650 (N_21650,N_12524,N_12527);
xor U21651 (N_21651,N_18386,N_14370);
or U21652 (N_21652,N_16408,N_16442);
xor U21653 (N_21653,N_17835,N_13841);
and U21654 (N_21654,N_12809,N_16310);
nand U21655 (N_21655,N_14252,N_14413);
xnor U21656 (N_21656,N_12981,N_16779);
xnor U21657 (N_21657,N_14380,N_17368);
and U21658 (N_21658,N_13416,N_17564);
nor U21659 (N_21659,N_16739,N_12907);
nand U21660 (N_21660,N_18121,N_12690);
xnor U21661 (N_21661,N_14717,N_15275);
and U21662 (N_21662,N_16226,N_18000);
xor U21663 (N_21663,N_18506,N_12871);
nor U21664 (N_21664,N_13857,N_13418);
or U21665 (N_21665,N_18169,N_13625);
nand U21666 (N_21666,N_14587,N_17139);
nand U21667 (N_21667,N_17734,N_17267);
nor U21668 (N_21668,N_16090,N_18072);
xnor U21669 (N_21669,N_16953,N_18119);
and U21670 (N_21670,N_18027,N_15756);
nor U21671 (N_21671,N_18343,N_14732);
and U21672 (N_21672,N_18485,N_12923);
and U21673 (N_21673,N_13186,N_15133);
nand U21674 (N_21674,N_14140,N_18681);
and U21675 (N_21675,N_15751,N_13201);
nor U21676 (N_21676,N_18232,N_13267);
nor U21677 (N_21677,N_14078,N_17118);
and U21678 (N_21678,N_17041,N_13509);
nor U21679 (N_21679,N_15760,N_17948);
or U21680 (N_21680,N_15122,N_17285);
nand U21681 (N_21681,N_15532,N_13364);
nor U21682 (N_21682,N_14165,N_17355);
xnor U21683 (N_21683,N_15272,N_18058);
or U21684 (N_21684,N_18649,N_16122);
and U21685 (N_21685,N_16058,N_15130);
nor U21686 (N_21686,N_14210,N_17046);
and U21687 (N_21687,N_15504,N_17213);
and U21688 (N_21688,N_14935,N_17309);
nand U21689 (N_21689,N_18108,N_12831);
nand U21690 (N_21690,N_18744,N_17072);
or U21691 (N_21691,N_15198,N_14045);
or U21692 (N_21692,N_17907,N_13990);
nand U21693 (N_21693,N_17571,N_15996);
nand U21694 (N_21694,N_15649,N_15048);
nand U21695 (N_21695,N_18213,N_14600);
xnor U21696 (N_21696,N_14973,N_13503);
or U21697 (N_21697,N_16331,N_18560);
and U21698 (N_21698,N_17212,N_14102);
nor U21699 (N_21699,N_13330,N_15612);
xor U21700 (N_21700,N_14671,N_14734);
and U21701 (N_21701,N_14961,N_17648);
nand U21702 (N_21702,N_18188,N_17165);
nand U21703 (N_21703,N_13074,N_18528);
xnor U21704 (N_21704,N_17588,N_15500);
or U21705 (N_21705,N_17533,N_16320);
and U21706 (N_21706,N_16574,N_15115);
nor U21707 (N_21707,N_13356,N_18650);
nand U21708 (N_21708,N_15870,N_16121);
xor U21709 (N_21709,N_17636,N_17376);
xor U21710 (N_21710,N_16350,N_16261);
and U21711 (N_21711,N_14949,N_15658);
xnor U21712 (N_21712,N_15443,N_17830);
xnor U21713 (N_21713,N_12867,N_15748);
nand U21714 (N_21714,N_13024,N_17874);
and U21715 (N_21715,N_16474,N_13061);
or U21716 (N_21716,N_17266,N_13636);
or U21717 (N_21717,N_14987,N_13158);
and U21718 (N_21718,N_16490,N_16059);
or U21719 (N_21719,N_14276,N_16526);
and U21720 (N_21720,N_17019,N_17853);
nand U21721 (N_21721,N_16189,N_13004);
nand U21722 (N_21722,N_13084,N_15584);
xor U21723 (N_21723,N_17004,N_14352);
nor U21724 (N_21724,N_12771,N_16568);
xnor U21725 (N_21725,N_15802,N_14814);
nor U21726 (N_21726,N_16123,N_13816);
or U21727 (N_21727,N_18698,N_17222);
nand U21728 (N_21728,N_14237,N_15391);
or U21729 (N_21729,N_16262,N_13985);
or U21730 (N_21730,N_12848,N_15552);
or U21731 (N_21731,N_17792,N_15978);
xor U21732 (N_21732,N_14471,N_14622);
xnor U21733 (N_21733,N_13174,N_18161);
xor U21734 (N_21734,N_13650,N_18365);
nand U21735 (N_21735,N_15499,N_15242);
nor U21736 (N_21736,N_18592,N_14452);
nand U21737 (N_21737,N_13068,N_15562);
or U21738 (N_21738,N_16829,N_14645);
or U21739 (N_21739,N_16559,N_16013);
nand U21740 (N_21740,N_13674,N_15896);
nand U21741 (N_21741,N_14982,N_13123);
nor U21742 (N_21742,N_18505,N_14510);
xnor U21743 (N_21743,N_13383,N_16243);
nand U21744 (N_21744,N_14425,N_15483);
xor U21745 (N_21745,N_15938,N_16617);
nor U21746 (N_21746,N_17132,N_13957);
or U21747 (N_21747,N_16222,N_15953);
nor U21748 (N_21748,N_15274,N_18504);
nor U21749 (N_21749,N_18747,N_18388);
nor U21750 (N_21750,N_15526,N_14859);
xnor U21751 (N_21751,N_18308,N_18284);
nand U21752 (N_21752,N_16700,N_16273);
nor U21753 (N_21753,N_17082,N_17461);
xor U21754 (N_21754,N_13821,N_17264);
or U21755 (N_21755,N_18209,N_15294);
and U21756 (N_21756,N_15290,N_14735);
nor U21757 (N_21757,N_17325,N_17190);
and U21758 (N_21758,N_17099,N_17802);
nor U21759 (N_21759,N_15877,N_14016);
or U21760 (N_21760,N_13982,N_13910);
and U21761 (N_21761,N_17167,N_14228);
xnor U21762 (N_21762,N_14205,N_14014);
nand U21763 (N_21763,N_12556,N_16612);
nand U21764 (N_21764,N_17981,N_14943);
or U21765 (N_21765,N_13044,N_12821);
nor U21766 (N_21766,N_18055,N_13891);
or U21767 (N_21767,N_18297,N_13508);
and U21768 (N_21768,N_18726,N_14726);
xnor U21769 (N_21769,N_15035,N_16227);
nor U21770 (N_21770,N_16354,N_17621);
and U21771 (N_21771,N_14286,N_14106);
nand U21772 (N_21772,N_14774,N_17458);
or U21773 (N_21773,N_15229,N_16336);
xnor U21774 (N_21774,N_15594,N_12738);
nor U21775 (N_21775,N_14475,N_13122);
xnor U21776 (N_21776,N_13271,N_16424);
and U21777 (N_21777,N_13939,N_15132);
and U21778 (N_21778,N_14013,N_12535);
nor U21779 (N_21779,N_14901,N_18721);
and U21780 (N_21780,N_16069,N_18345);
or U21781 (N_21781,N_14591,N_13699);
nand U21782 (N_21782,N_17610,N_16051);
or U21783 (N_21783,N_14159,N_16257);
nand U21784 (N_21784,N_16740,N_13847);
nand U21785 (N_21785,N_16805,N_18210);
nor U21786 (N_21786,N_15012,N_15456);
nand U21787 (N_21787,N_16415,N_14767);
or U21788 (N_21788,N_14075,N_18486);
nand U21789 (N_21789,N_14792,N_12972);
and U21790 (N_21790,N_18407,N_15752);
and U21791 (N_21791,N_18123,N_16919);
nand U21792 (N_21792,N_14998,N_15872);
xor U21793 (N_21793,N_17411,N_16512);
and U21794 (N_21794,N_15051,N_14696);
nand U21795 (N_21795,N_12977,N_13983);
or U21796 (N_21796,N_15643,N_17751);
and U21797 (N_21797,N_13898,N_14713);
or U21798 (N_21798,N_17414,N_15415);
nor U21799 (N_21799,N_14244,N_12567);
or U21800 (N_21800,N_15761,N_14891);
xor U21801 (N_21801,N_17121,N_17982);
and U21802 (N_21802,N_15116,N_17294);
xor U21803 (N_21803,N_15510,N_14829);
and U21804 (N_21804,N_12752,N_12585);
nand U21805 (N_21805,N_17159,N_12741);
nand U21806 (N_21806,N_13728,N_16179);
xor U21807 (N_21807,N_18416,N_12692);
and U21808 (N_21808,N_15258,N_17219);
and U21809 (N_21809,N_14335,N_15790);
or U21810 (N_21810,N_18312,N_17991);
xnor U21811 (N_21811,N_16944,N_16030);
nand U21812 (N_21812,N_15855,N_16640);
xnor U21813 (N_21813,N_18566,N_15339);
xor U21814 (N_21814,N_17502,N_13700);
or U21815 (N_21815,N_14230,N_13458);
or U21816 (N_21816,N_13651,N_13405);
xor U21817 (N_21817,N_17766,N_12838);
or U21818 (N_21818,N_13646,N_14892);
xor U21819 (N_21819,N_18141,N_14272);
and U21820 (N_21820,N_12694,N_18162);
or U21821 (N_21821,N_14239,N_13161);
xor U21822 (N_21822,N_17395,N_12802);
nand U21823 (N_21823,N_17890,N_12546);
nor U21824 (N_21824,N_14739,N_17631);
or U21825 (N_21825,N_16282,N_16348);
or U21826 (N_21826,N_18728,N_15548);
nand U21827 (N_21827,N_16478,N_17034);
or U21828 (N_21828,N_15331,N_13256);
nand U21829 (N_21829,N_14955,N_15383);
or U21830 (N_21830,N_18190,N_14660);
nand U21831 (N_21831,N_13333,N_15001);
and U21832 (N_21832,N_17855,N_15546);
nand U21833 (N_21833,N_12526,N_12764);
nor U21834 (N_21834,N_13598,N_16642);
nor U21835 (N_21835,N_12590,N_16132);
nand U21836 (N_21836,N_17990,N_13740);
xor U21837 (N_21837,N_14233,N_17944);
and U21838 (N_21838,N_13723,N_13140);
and U21839 (N_21839,N_18333,N_14699);
xor U21840 (N_21840,N_13500,N_16198);
xnor U21841 (N_21841,N_15069,N_18557);
or U21842 (N_21842,N_15633,N_15569);
nand U21843 (N_21843,N_16187,N_17020);
nor U21844 (N_21844,N_13934,N_16200);
and U21845 (N_21845,N_17337,N_13873);
nand U21846 (N_21846,N_14308,N_16903);
nand U21847 (N_21847,N_18573,N_13941);
and U21848 (N_21848,N_17576,N_16814);
xnor U21849 (N_21849,N_12948,N_14251);
and U21850 (N_21850,N_15593,N_16223);
or U21851 (N_21851,N_13627,N_15634);
and U21852 (N_21852,N_12591,N_13332);
nand U21853 (N_21853,N_12640,N_15626);
xnor U21854 (N_21854,N_15263,N_16146);
xor U21855 (N_21855,N_16113,N_17338);
or U21856 (N_21856,N_13582,N_15541);
nor U21857 (N_21857,N_16599,N_18385);
or U21858 (N_21858,N_17794,N_18664);
and U21859 (N_21859,N_15222,N_12807);
and U21860 (N_21860,N_17224,N_18279);
and U21861 (N_21861,N_14927,N_15471);
or U21862 (N_21862,N_17272,N_13143);
or U21863 (N_21863,N_13243,N_18320);
or U21864 (N_21864,N_13867,N_15892);
nand U21865 (N_21865,N_14952,N_14388);
nor U21866 (N_21866,N_15151,N_12889);
and U21867 (N_21867,N_13346,N_15882);
or U21868 (N_21868,N_14189,N_16554);
nor U21869 (N_21869,N_14158,N_16584);
nor U21870 (N_21870,N_13881,N_14304);
and U21871 (N_21871,N_16185,N_17993);
nand U21872 (N_21872,N_18743,N_18375);
xnor U21873 (N_21873,N_16020,N_14409);
or U21874 (N_21874,N_14278,N_15176);
or U21875 (N_21875,N_18438,N_16452);
nor U21876 (N_21876,N_12529,N_18007);
nand U21877 (N_21877,N_14083,N_14485);
nor U21878 (N_21878,N_12747,N_13868);
and U21879 (N_21879,N_13996,N_14379);
nand U21880 (N_21880,N_12714,N_17714);
or U21881 (N_21881,N_18717,N_12607);
nand U21882 (N_21882,N_17417,N_14500);
xor U21883 (N_21883,N_16969,N_16171);
nand U21884 (N_21884,N_17328,N_12652);
xor U21885 (N_21885,N_14660,N_17186);
nand U21886 (N_21886,N_14323,N_15006);
xor U21887 (N_21887,N_15156,N_16392);
nor U21888 (N_21888,N_18544,N_18324);
xnor U21889 (N_21889,N_17686,N_16959);
nand U21890 (N_21890,N_18206,N_17759);
nand U21891 (N_21891,N_18255,N_15502);
xnor U21892 (N_21892,N_17268,N_14710);
xnor U21893 (N_21893,N_15048,N_17893);
nand U21894 (N_21894,N_13886,N_18713);
xor U21895 (N_21895,N_13922,N_18186);
nand U21896 (N_21896,N_18410,N_18497);
xnor U21897 (N_21897,N_17961,N_16803);
nor U21898 (N_21898,N_13680,N_14616);
xnor U21899 (N_21899,N_18497,N_14840);
or U21900 (N_21900,N_16562,N_18287);
or U21901 (N_21901,N_14970,N_14758);
nand U21902 (N_21902,N_13101,N_17865);
xor U21903 (N_21903,N_16794,N_17291);
nor U21904 (N_21904,N_17481,N_18622);
nor U21905 (N_21905,N_17851,N_17992);
or U21906 (N_21906,N_18698,N_15516);
xor U21907 (N_21907,N_13853,N_14925);
and U21908 (N_21908,N_15621,N_17689);
nand U21909 (N_21909,N_18353,N_16887);
and U21910 (N_21910,N_18467,N_14315);
xnor U21911 (N_21911,N_17207,N_12632);
nor U21912 (N_21912,N_13792,N_15072);
or U21913 (N_21913,N_13650,N_14961);
or U21914 (N_21914,N_15027,N_14362);
nand U21915 (N_21915,N_14720,N_14007);
nor U21916 (N_21916,N_17477,N_15937);
and U21917 (N_21917,N_15397,N_15024);
nor U21918 (N_21918,N_16662,N_15458);
nor U21919 (N_21919,N_15018,N_13626);
nor U21920 (N_21920,N_13898,N_15269);
xor U21921 (N_21921,N_13858,N_16027);
or U21922 (N_21922,N_16985,N_15826);
and U21923 (N_21923,N_15789,N_16573);
and U21924 (N_21924,N_16694,N_12642);
or U21925 (N_21925,N_12689,N_14702);
xor U21926 (N_21926,N_17878,N_17010);
and U21927 (N_21927,N_18159,N_18620);
xor U21928 (N_21928,N_17357,N_15066);
nor U21929 (N_21929,N_13583,N_16248);
or U21930 (N_21930,N_12697,N_13390);
xor U21931 (N_21931,N_16072,N_13960);
nand U21932 (N_21932,N_13519,N_16091);
nand U21933 (N_21933,N_16539,N_17129);
and U21934 (N_21934,N_13508,N_14005);
and U21935 (N_21935,N_18152,N_17927);
nor U21936 (N_21936,N_12684,N_17161);
xor U21937 (N_21937,N_12632,N_16719);
nor U21938 (N_21938,N_14351,N_15984);
nand U21939 (N_21939,N_13970,N_17610);
nor U21940 (N_21940,N_14461,N_14653);
nand U21941 (N_21941,N_16514,N_13005);
nor U21942 (N_21942,N_17070,N_15707);
nor U21943 (N_21943,N_12659,N_15524);
nand U21944 (N_21944,N_15533,N_18337);
nor U21945 (N_21945,N_17879,N_16740);
nor U21946 (N_21946,N_16156,N_14812);
and U21947 (N_21947,N_18595,N_16014);
nor U21948 (N_21948,N_12742,N_16161);
nand U21949 (N_21949,N_15661,N_17761);
nand U21950 (N_21950,N_16930,N_12779);
nand U21951 (N_21951,N_14221,N_13750);
nand U21952 (N_21952,N_17610,N_16379);
nand U21953 (N_21953,N_14846,N_15497);
or U21954 (N_21954,N_15430,N_15038);
xor U21955 (N_21955,N_13854,N_17067);
nor U21956 (N_21956,N_17546,N_15994);
or U21957 (N_21957,N_17959,N_14394);
nand U21958 (N_21958,N_15095,N_15817);
and U21959 (N_21959,N_18019,N_14806);
and U21960 (N_21960,N_16126,N_13834);
and U21961 (N_21961,N_15051,N_18663);
or U21962 (N_21962,N_14186,N_16351);
and U21963 (N_21963,N_15211,N_18034);
and U21964 (N_21964,N_15182,N_12999);
xnor U21965 (N_21965,N_16635,N_13950);
and U21966 (N_21966,N_14651,N_17731);
nand U21967 (N_21967,N_16723,N_12930);
nor U21968 (N_21968,N_15466,N_18693);
nand U21969 (N_21969,N_18241,N_12630);
and U21970 (N_21970,N_16492,N_13495);
or U21971 (N_21971,N_16270,N_15334);
xor U21972 (N_21972,N_15641,N_16421);
nand U21973 (N_21973,N_13559,N_12711);
xnor U21974 (N_21974,N_13498,N_16348);
nand U21975 (N_21975,N_17058,N_17105);
and U21976 (N_21976,N_17110,N_13750);
or U21977 (N_21977,N_15647,N_15190);
or U21978 (N_21978,N_12855,N_18211);
nor U21979 (N_21979,N_15192,N_16799);
or U21980 (N_21980,N_17988,N_15232);
xor U21981 (N_21981,N_14262,N_18212);
nand U21982 (N_21982,N_16166,N_13995);
nand U21983 (N_21983,N_18184,N_16440);
nand U21984 (N_21984,N_17199,N_14713);
and U21985 (N_21985,N_14583,N_18123);
nor U21986 (N_21986,N_13424,N_17405);
or U21987 (N_21987,N_17788,N_12897);
nand U21988 (N_21988,N_16735,N_13929);
and U21989 (N_21989,N_13777,N_12800);
or U21990 (N_21990,N_18519,N_16689);
xnor U21991 (N_21991,N_15803,N_17454);
nand U21992 (N_21992,N_17539,N_16144);
and U21993 (N_21993,N_13510,N_14176);
and U21994 (N_21994,N_14007,N_18020);
xor U21995 (N_21995,N_13403,N_15890);
or U21996 (N_21996,N_18341,N_13877);
xor U21997 (N_21997,N_14618,N_17878);
xor U21998 (N_21998,N_14806,N_14981);
xnor U21999 (N_21999,N_14846,N_15151);
and U22000 (N_22000,N_12964,N_16992);
or U22001 (N_22001,N_17533,N_15736);
nand U22002 (N_22002,N_14071,N_12725);
and U22003 (N_22003,N_13942,N_16533);
and U22004 (N_22004,N_15772,N_16916);
nor U22005 (N_22005,N_17858,N_15031);
nand U22006 (N_22006,N_14946,N_14188);
and U22007 (N_22007,N_16204,N_16767);
nor U22008 (N_22008,N_15381,N_16922);
xnor U22009 (N_22009,N_13345,N_17738);
nor U22010 (N_22010,N_14313,N_18305);
or U22011 (N_22011,N_15856,N_16034);
xnor U22012 (N_22012,N_12626,N_14739);
and U22013 (N_22013,N_16816,N_15425);
and U22014 (N_22014,N_16274,N_13888);
xnor U22015 (N_22015,N_18505,N_16459);
or U22016 (N_22016,N_18599,N_12811);
or U22017 (N_22017,N_17086,N_17938);
nand U22018 (N_22018,N_17546,N_15810);
nand U22019 (N_22019,N_16101,N_16325);
xor U22020 (N_22020,N_13906,N_12583);
nor U22021 (N_22021,N_16653,N_13241);
nor U22022 (N_22022,N_15973,N_14867);
nand U22023 (N_22023,N_16645,N_15230);
xnor U22024 (N_22024,N_14746,N_12863);
xor U22025 (N_22025,N_17168,N_17370);
and U22026 (N_22026,N_14829,N_18428);
and U22027 (N_22027,N_18271,N_14733);
and U22028 (N_22028,N_15949,N_14023);
xnor U22029 (N_22029,N_13242,N_14945);
nand U22030 (N_22030,N_14628,N_17800);
or U22031 (N_22031,N_12741,N_13924);
nor U22032 (N_22032,N_15437,N_17571);
and U22033 (N_22033,N_15285,N_16924);
and U22034 (N_22034,N_16187,N_17634);
and U22035 (N_22035,N_17869,N_14077);
nor U22036 (N_22036,N_13031,N_12602);
or U22037 (N_22037,N_16672,N_17404);
or U22038 (N_22038,N_17183,N_13889);
nor U22039 (N_22039,N_14580,N_13819);
and U22040 (N_22040,N_14412,N_17760);
nand U22041 (N_22041,N_12552,N_13227);
or U22042 (N_22042,N_15349,N_14117);
nand U22043 (N_22043,N_15740,N_18212);
nand U22044 (N_22044,N_17802,N_14776);
xor U22045 (N_22045,N_14828,N_12544);
nand U22046 (N_22046,N_17357,N_15193);
nand U22047 (N_22047,N_15168,N_16510);
and U22048 (N_22048,N_16397,N_18576);
nand U22049 (N_22049,N_16588,N_13412);
and U22050 (N_22050,N_17413,N_18458);
and U22051 (N_22051,N_13666,N_14349);
nor U22052 (N_22052,N_16781,N_12576);
nand U22053 (N_22053,N_16966,N_14309);
and U22054 (N_22054,N_12603,N_13690);
nor U22055 (N_22055,N_15130,N_14036);
and U22056 (N_22056,N_17840,N_13135);
nor U22057 (N_22057,N_13489,N_14976);
xnor U22058 (N_22058,N_12782,N_13499);
and U22059 (N_22059,N_15992,N_13495);
nand U22060 (N_22060,N_16865,N_13934);
xor U22061 (N_22061,N_14222,N_12919);
and U22062 (N_22062,N_12652,N_18303);
xor U22063 (N_22063,N_18743,N_17842);
or U22064 (N_22064,N_14304,N_18466);
nor U22065 (N_22065,N_13190,N_17465);
or U22066 (N_22066,N_15486,N_13599);
and U22067 (N_22067,N_16119,N_17937);
xor U22068 (N_22068,N_13897,N_15883);
nand U22069 (N_22069,N_18699,N_13398);
xor U22070 (N_22070,N_13563,N_18569);
or U22071 (N_22071,N_15986,N_13296);
and U22072 (N_22072,N_17273,N_13977);
nor U22073 (N_22073,N_13329,N_13569);
xor U22074 (N_22074,N_15279,N_13477);
and U22075 (N_22075,N_16685,N_12893);
nand U22076 (N_22076,N_14755,N_14205);
xnor U22077 (N_22077,N_15039,N_14320);
and U22078 (N_22078,N_16160,N_16601);
nand U22079 (N_22079,N_17859,N_17701);
and U22080 (N_22080,N_18630,N_14025);
xor U22081 (N_22081,N_12649,N_13129);
xor U22082 (N_22082,N_12684,N_16698);
and U22083 (N_22083,N_13418,N_13798);
and U22084 (N_22084,N_16693,N_14796);
nor U22085 (N_22085,N_16865,N_14173);
xnor U22086 (N_22086,N_17506,N_15434);
xor U22087 (N_22087,N_15556,N_13585);
nor U22088 (N_22088,N_14668,N_15280);
nand U22089 (N_22089,N_18190,N_15397);
nand U22090 (N_22090,N_17098,N_12849);
nand U22091 (N_22091,N_16730,N_16144);
nand U22092 (N_22092,N_14079,N_17024);
nor U22093 (N_22093,N_17962,N_15328);
xor U22094 (N_22094,N_14866,N_16162);
xnor U22095 (N_22095,N_14788,N_16348);
nor U22096 (N_22096,N_17787,N_15093);
xnor U22097 (N_22097,N_14418,N_14902);
and U22098 (N_22098,N_17342,N_13778);
and U22099 (N_22099,N_17903,N_13863);
nor U22100 (N_22100,N_16390,N_17529);
nand U22101 (N_22101,N_14368,N_14661);
or U22102 (N_22102,N_12900,N_13255);
nand U22103 (N_22103,N_17698,N_18539);
and U22104 (N_22104,N_12705,N_16548);
or U22105 (N_22105,N_17492,N_18556);
nand U22106 (N_22106,N_15109,N_12839);
nor U22107 (N_22107,N_17285,N_14918);
and U22108 (N_22108,N_13318,N_15563);
and U22109 (N_22109,N_17904,N_15200);
and U22110 (N_22110,N_16691,N_17066);
or U22111 (N_22111,N_15834,N_14690);
xor U22112 (N_22112,N_12710,N_14129);
xor U22113 (N_22113,N_12510,N_15046);
and U22114 (N_22114,N_13577,N_17470);
or U22115 (N_22115,N_14686,N_18247);
or U22116 (N_22116,N_16210,N_13913);
and U22117 (N_22117,N_15736,N_14345);
and U22118 (N_22118,N_14549,N_17602);
nor U22119 (N_22119,N_14831,N_16792);
xnor U22120 (N_22120,N_15654,N_17104);
nor U22121 (N_22121,N_15723,N_16851);
nor U22122 (N_22122,N_15448,N_15686);
or U22123 (N_22123,N_15026,N_17206);
xor U22124 (N_22124,N_18495,N_16984);
or U22125 (N_22125,N_16893,N_12819);
xor U22126 (N_22126,N_17360,N_12976);
xor U22127 (N_22127,N_18435,N_18710);
nor U22128 (N_22128,N_16838,N_14880);
and U22129 (N_22129,N_13746,N_15218);
xnor U22130 (N_22130,N_17549,N_12585);
or U22131 (N_22131,N_14348,N_17104);
nor U22132 (N_22132,N_12996,N_17757);
nor U22133 (N_22133,N_14554,N_17764);
or U22134 (N_22134,N_13034,N_16996);
nand U22135 (N_22135,N_14786,N_17471);
or U22136 (N_22136,N_18522,N_18245);
and U22137 (N_22137,N_18460,N_15384);
nand U22138 (N_22138,N_14635,N_14433);
xor U22139 (N_22139,N_15603,N_18367);
or U22140 (N_22140,N_15319,N_14672);
nand U22141 (N_22141,N_18105,N_18085);
and U22142 (N_22142,N_14057,N_17580);
or U22143 (N_22143,N_13596,N_13120);
nor U22144 (N_22144,N_12904,N_18087);
or U22145 (N_22145,N_16920,N_13874);
nor U22146 (N_22146,N_14155,N_14938);
and U22147 (N_22147,N_13882,N_14994);
nand U22148 (N_22148,N_17601,N_16113);
xor U22149 (N_22149,N_15487,N_17152);
and U22150 (N_22150,N_14990,N_16649);
xor U22151 (N_22151,N_18441,N_16277);
nand U22152 (N_22152,N_18306,N_18319);
nand U22153 (N_22153,N_12864,N_16039);
xor U22154 (N_22154,N_17644,N_15559);
xor U22155 (N_22155,N_14251,N_17508);
xnor U22156 (N_22156,N_16087,N_12699);
and U22157 (N_22157,N_17361,N_15337);
or U22158 (N_22158,N_13924,N_14603);
nand U22159 (N_22159,N_18674,N_17770);
nand U22160 (N_22160,N_13740,N_13138);
and U22161 (N_22161,N_14957,N_17369);
or U22162 (N_22162,N_16703,N_18401);
nor U22163 (N_22163,N_15378,N_17228);
xor U22164 (N_22164,N_13578,N_16616);
and U22165 (N_22165,N_14221,N_15966);
or U22166 (N_22166,N_13571,N_13268);
or U22167 (N_22167,N_16348,N_15427);
and U22168 (N_22168,N_17788,N_16758);
nand U22169 (N_22169,N_14893,N_14422);
or U22170 (N_22170,N_18559,N_14406);
nor U22171 (N_22171,N_14683,N_12924);
xor U22172 (N_22172,N_17087,N_13183);
or U22173 (N_22173,N_16913,N_12613);
nor U22174 (N_22174,N_14136,N_12576);
nand U22175 (N_22175,N_17789,N_15628);
and U22176 (N_22176,N_14051,N_13348);
nor U22177 (N_22177,N_14208,N_18575);
nand U22178 (N_22178,N_16795,N_13030);
and U22179 (N_22179,N_16659,N_17081);
nand U22180 (N_22180,N_18739,N_13408);
or U22181 (N_22181,N_16308,N_14492);
nor U22182 (N_22182,N_14718,N_15634);
or U22183 (N_22183,N_17915,N_18177);
or U22184 (N_22184,N_17087,N_17762);
nor U22185 (N_22185,N_14052,N_16660);
xnor U22186 (N_22186,N_12852,N_15872);
nand U22187 (N_22187,N_16480,N_16337);
and U22188 (N_22188,N_13907,N_16861);
and U22189 (N_22189,N_14467,N_16321);
xor U22190 (N_22190,N_18132,N_18272);
nand U22191 (N_22191,N_14801,N_14911);
nor U22192 (N_22192,N_14393,N_13354);
xor U22193 (N_22193,N_14452,N_14660);
or U22194 (N_22194,N_17043,N_18641);
nor U22195 (N_22195,N_16463,N_18626);
xnor U22196 (N_22196,N_13236,N_12858);
or U22197 (N_22197,N_18704,N_14059);
or U22198 (N_22198,N_17993,N_14658);
xor U22199 (N_22199,N_18272,N_16527);
xnor U22200 (N_22200,N_15980,N_16318);
and U22201 (N_22201,N_16015,N_17622);
and U22202 (N_22202,N_12594,N_14637);
or U22203 (N_22203,N_14646,N_16149);
or U22204 (N_22204,N_15778,N_18345);
or U22205 (N_22205,N_15216,N_15829);
nand U22206 (N_22206,N_15113,N_15136);
or U22207 (N_22207,N_18393,N_13088);
nor U22208 (N_22208,N_14510,N_14532);
nor U22209 (N_22209,N_15303,N_15496);
and U22210 (N_22210,N_13318,N_13401);
nor U22211 (N_22211,N_13126,N_14188);
nor U22212 (N_22212,N_13391,N_13619);
xnor U22213 (N_22213,N_13904,N_17399);
xnor U22214 (N_22214,N_18313,N_13598);
nand U22215 (N_22215,N_17710,N_16770);
and U22216 (N_22216,N_16668,N_17032);
and U22217 (N_22217,N_18490,N_18113);
and U22218 (N_22218,N_15405,N_14574);
xnor U22219 (N_22219,N_15503,N_17218);
xnor U22220 (N_22220,N_17459,N_13354);
xor U22221 (N_22221,N_16241,N_16758);
and U22222 (N_22222,N_18531,N_18504);
nor U22223 (N_22223,N_12913,N_14726);
xnor U22224 (N_22224,N_14966,N_13560);
nand U22225 (N_22225,N_14417,N_18123);
or U22226 (N_22226,N_14414,N_13625);
and U22227 (N_22227,N_15478,N_14571);
and U22228 (N_22228,N_16783,N_17183);
nand U22229 (N_22229,N_15635,N_13794);
nand U22230 (N_22230,N_15834,N_15943);
xnor U22231 (N_22231,N_14944,N_15684);
and U22232 (N_22232,N_13200,N_13707);
nand U22233 (N_22233,N_17843,N_15649);
and U22234 (N_22234,N_16031,N_16492);
nand U22235 (N_22235,N_15154,N_17279);
xnor U22236 (N_22236,N_17077,N_17865);
nor U22237 (N_22237,N_16532,N_16973);
nand U22238 (N_22238,N_14311,N_18078);
and U22239 (N_22239,N_15481,N_13968);
or U22240 (N_22240,N_14045,N_12592);
and U22241 (N_22241,N_17477,N_14722);
or U22242 (N_22242,N_13505,N_12893);
and U22243 (N_22243,N_18361,N_14943);
xor U22244 (N_22244,N_13378,N_13148);
nor U22245 (N_22245,N_17493,N_16848);
nand U22246 (N_22246,N_15954,N_15588);
nand U22247 (N_22247,N_15021,N_13340);
nand U22248 (N_22248,N_15760,N_13857);
and U22249 (N_22249,N_17015,N_13141);
xnor U22250 (N_22250,N_16997,N_14254);
or U22251 (N_22251,N_15184,N_14986);
nor U22252 (N_22252,N_17022,N_16960);
or U22253 (N_22253,N_15690,N_14886);
or U22254 (N_22254,N_17159,N_16560);
nor U22255 (N_22255,N_13980,N_17857);
or U22256 (N_22256,N_15446,N_16748);
nand U22257 (N_22257,N_18525,N_15460);
xor U22258 (N_22258,N_17947,N_13593);
and U22259 (N_22259,N_16880,N_13527);
nor U22260 (N_22260,N_18468,N_17158);
and U22261 (N_22261,N_16010,N_13234);
nor U22262 (N_22262,N_15090,N_13456);
xor U22263 (N_22263,N_13857,N_16285);
and U22264 (N_22264,N_13041,N_12955);
or U22265 (N_22265,N_14316,N_16870);
nor U22266 (N_22266,N_18598,N_18660);
and U22267 (N_22267,N_16177,N_16058);
and U22268 (N_22268,N_17350,N_17853);
nand U22269 (N_22269,N_12971,N_13507);
and U22270 (N_22270,N_13854,N_16150);
nor U22271 (N_22271,N_14395,N_18445);
and U22272 (N_22272,N_15351,N_13049);
nand U22273 (N_22273,N_13828,N_15748);
xor U22274 (N_22274,N_13654,N_16288);
and U22275 (N_22275,N_12810,N_15190);
nand U22276 (N_22276,N_18734,N_14079);
nor U22277 (N_22277,N_13260,N_13423);
xnor U22278 (N_22278,N_13896,N_18290);
xor U22279 (N_22279,N_18037,N_17197);
nand U22280 (N_22280,N_15097,N_16667);
nand U22281 (N_22281,N_17303,N_16299);
nand U22282 (N_22282,N_14033,N_17325);
nand U22283 (N_22283,N_17172,N_17882);
or U22284 (N_22284,N_15079,N_13640);
nor U22285 (N_22285,N_17602,N_14997);
or U22286 (N_22286,N_16399,N_17002);
nand U22287 (N_22287,N_12734,N_13457);
xnor U22288 (N_22288,N_18704,N_13793);
and U22289 (N_22289,N_13507,N_14186);
and U22290 (N_22290,N_14665,N_16111);
or U22291 (N_22291,N_14334,N_13335);
or U22292 (N_22292,N_14275,N_17322);
nand U22293 (N_22293,N_18737,N_15215);
or U22294 (N_22294,N_18258,N_13671);
nor U22295 (N_22295,N_15024,N_15089);
and U22296 (N_22296,N_15021,N_13104);
xor U22297 (N_22297,N_13052,N_13990);
xor U22298 (N_22298,N_17670,N_14234);
nand U22299 (N_22299,N_12550,N_13000);
or U22300 (N_22300,N_14663,N_14264);
or U22301 (N_22301,N_16372,N_16132);
xor U22302 (N_22302,N_16093,N_17051);
nor U22303 (N_22303,N_15121,N_17738);
and U22304 (N_22304,N_16478,N_18485);
nor U22305 (N_22305,N_14224,N_14591);
and U22306 (N_22306,N_17213,N_15691);
nand U22307 (N_22307,N_13910,N_15273);
nor U22308 (N_22308,N_17665,N_14527);
nor U22309 (N_22309,N_12574,N_18348);
or U22310 (N_22310,N_15442,N_15324);
nand U22311 (N_22311,N_14491,N_14836);
nand U22312 (N_22312,N_15593,N_15131);
xor U22313 (N_22313,N_18644,N_12570);
nor U22314 (N_22314,N_18293,N_15197);
and U22315 (N_22315,N_12698,N_14013);
nand U22316 (N_22316,N_13108,N_13746);
xor U22317 (N_22317,N_14578,N_18262);
nand U22318 (N_22318,N_16491,N_15976);
and U22319 (N_22319,N_18569,N_13018);
nand U22320 (N_22320,N_18398,N_17641);
nor U22321 (N_22321,N_15535,N_14697);
xnor U22322 (N_22322,N_18158,N_14607);
and U22323 (N_22323,N_16481,N_13491);
and U22324 (N_22324,N_17780,N_15771);
and U22325 (N_22325,N_16170,N_15730);
xor U22326 (N_22326,N_15085,N_18509);
or U22327 (N_22327,N_17594,N_12745);
nand U22328 (N_22328,N_16611,N_14288);
and U22329 (N_22329,N_17387,N_15391);
or U22330 (N_22330,N_13289,N_13307);
or U22331 (N_22331,N_14951,N_16279);
xnor U22332 (N_22332,N_16745,N_13957);
and U22333 (N_22333,N_13100,N_14353);
nand U22334 (N_22334,N_18442,N_14337);
and U22335 (N_22335,N_13809,N_15372);
nand U22336 (N_22336,N_14850,N_14653);
or U22337 (N_22337,N_15012,N_15120);
xnor U22338 (N_22338,N_18159,N_13285);
nand U22339 (N_22339,N_14653,N_17360);
and U22340 (N_22340,N_13153,N_15593);
nand U22341 (N_22341,N_16583,N_16449);
xnor U22342 (N_22342,N_12551,N_15323);
nor U22343 (N_22343,N_14755,N_13532);
or U22344 (N_22344,N_13036,N_17738);
nor U22345 (N_22345,N_14941,N_15304);
or U22346 (N_22346,N_13156,N_12521);
nor U22347 (N_22347,N_13914,N_18369);
xor U22348 (N_22348,N_17591,N_17450);
nor U22349 (N_22349,N_12622,N_16585);
nor U22350 (N_22350,N_16169,N_17349);
and U22351 (N_22351,N_17946,N_16248);
and U22352 (N_22352,N_17565,N_17938);
or U22353 (N_22353,N_15798,N_15544);
or U22354 (N_22354,N_15218,N_14641);
nor U22355 (N_22355,N_17338,N_14516);
nand U22356 (N_22356,N_16057,N_18600);
and U22357 (N_22357,N_14898,N_13813);
nor U22358 (N_22358,N_15941,N_14612);
or U22359 (N_22359,N_15491,N_12728);
nand U22360 (N_22360,N_12582,N_15279);
xor U22361 (N_22361,N_17477,N_14075);
and U22362 (N_22362,N_13882,N_13472);
nor U22363 (N_22363,N_12615,N_18376);
nand U22364 (N_22364,N_15138,N_17072);
nand U22365 (N_22365,N_13371,N_13918);
or U22366 (N_22366,N_18590,N_17197);
nand U22367 (N_22367,N_13617,N_16613);
nand U22368 (N_22368,N_18130,N_16316);
xor U22369 (N_22369,N_17303,N_14028);
nand U22370 (N_22370,N_14567,N_18543);
and U22371 (N_22371,N_18244,N_12684);
and U22372 (N_22372,N_14291,N_18647);
nand U22373 (N_22373,N_13931,N_14716);
nand U22374 (N_22374,N_17856,N_14082);
and U22375 (N_22375,N_13694,N_18691);
or U22376 (N_22376,N_13669,N_14738);
xor U22377 (N_22377,N_15574,N_12523);
or U22378 (N_22378,N_17005,N_17182);
nand U22379 (N_22379,N_12914,N_12678);
and U22380 (N_22380,N_13628,N_14565);
or U22381 (N_22381,N_17104,N_14074);
nor U22382 (N_22382,N_12577,N_16367);
nor U22383 (N_22383,N_18319,N_16588);
or U22384 (N_22384,N_17783,N_17146);
or U22385 (N_22385,N_16773,N_18118);
nand U22386 (N_22386,N_13076,N_16389);
xor U22387 (N_22387,N_17863,N_15236);
nand U22388 (N_22388,N_17544,N_15697);
and U22389 (N_22389,N_15416,N_13270);
xor U22390 (N_22390,N_12980,N_18364);
xnor U22391 (N_22391,N_12517,N_14026);
nor U22392 (N_22392,N_15020,N_13594);
xnor U22393 (N_22393,N_14718,N_18020);
and U22394 (N_22394,N_17570,N_13669);
nand U22395 (N_22395,N_16032,N_16752);
or U22396 (N_22396,N_18437,N_18064);
xor U22397 (N_22397,N_13622,N_15186);
and U22398 (N_22398,N_12984,N_14820);
xnor U22399 (N_22399,N_12896,N_15865);
or U22400 (N_22400,N_15037,N_14478);
and U22401 (N_22401,N_15142,N_13607);
nand U22402 (N_22402,N_18499,N_14333);
nor U22403 (N_22403,N_14077,N_12803);
and U22404 (N_22404,N_13698,N_15321);
xnor U22405 (N_22405,N_14999,N_14599);
or U22406 (N_22406,N_13481,N_18033);
nor U22407 (N_22407,N_14483,N_17203);
or U22408 (N_22408,N_13871,N_15235);
and U22409 (N_22409,N_18513,N_14560);
nor U22410 (N_22410,N_14514,N_17407);
or U22411 (N_22411,N_13894,N_18109);
xor U22412 (N_22412,N_15723,N_17096);
xnor U22413 (N_22413,N_18225,N_18085);
and U22414 (N_22414,N_13305,N_12726);
xnor U22415 (N_22415,N_13920,N_17065);
nor U22416 (N_22416,N_16501,N_16978);
and U22417 (N_22417,N_17070,N_16864);
nor U22418 (N_22418,N_13274,N_15490);
nand U22419 (N_22419,N_16343,N_14134);
nor U22420 (N_22420,N_12589,N_15322);
nor U22421 (N_22421,N_12604,N_13361);
nor U22422 (N_22422,N_14843,N_16774);
nand U22423 (N_22423,N_14912,N_14110);
xnor U22424 (N_22424,N_17282,N_15048);
nand U22425 (N_22425,N_15851,N_16549);
xnor U22426 (N_22426,N_18237,N_15464);
and U22427 (N_22427,N_18107,N_18034);
or U22428 (N_22428,N_14703,N_17814);
nor U22429 (N_22429,N_16724,N_13829);
nor U22430 (N_22430,N_13957,N_17719);
nand U22431 (N_22431,N_17285,N_13100);
or U22432 (N_22432,N_14277,N_13078);
xor U22433 (N_22433,N_17970,N_16092);
or U22434 (N_22434,N_17554,N_17235);
nand U22435 (N_22435,N_12575,N_18092);
or U22436 (N_22436,N_15375,N_17889);
nand U22437 (N_22437,N_18712,N_12935);
xor U22438 (N_22438,N_13134,N_13873);
nor U22439 (N_22439,N_13904,N_17489);
nand U22440 (N_22440,N_18075,N_13897);
nor U22441 (N_22441,N_15486,N_14211);
or U22442 (N_22442,N_16296,N_12639);
nand U22443 (N_22443,N_13513,N_15846);
xnor U22444 (N_22444,N_18016,N_18381);
nand U22445 (N_22445,N_17099,N_16346);
nor U22446 (N_22446,N_14344,N_17165);
xnor U22447 (N_22447,N_14447,N_14836);
nor U22448 (N_22448,N_16168,N_12860);
xnor U22449 (N_22449,N_12584,N_16031);
and U22450 (N_22450,N_17107,N_14098);
or U22451 (N_22451,N_14796,N_13441);
nor U22452 (N_22452,N_15181,N_17270);
xnor U22453 (N_22453,N_17891,N_18037);
nor U22454 (N_22454,N_15247,N_14149);
and U22455 (N_22455,N_17445,N_17003);
nor U22456 (N_22456,N_16951,N_15344);
or U22457 (N_22457,N_12951,N_16727);
or U22458 (N_22458,N_13714,N_15521);
xor U22459 (N_22459,N_18490,N_17929);
nor U22460 (N_22460,N_12657,N_14841);
and U22461 (N_22461,N_15016,N_15512);
or U22462 (N_22462,N_16801,N_18089);
xnor U22463 (N_22463,N_14768,N_13393);
and U22464 (N_22464,N_16975,N_14360);
xor U22465 (N_22465,N_14411,N_13512);
xnor U22466 (N_22466,N_12915,N_14722);
and U22467 (N_22467,N_17709,N_18149);
nor U22468 (N_22468,N_18582,N_14563);
nand U22469 (N_22469,N_15283,N_16061);
xnor U22470 (N_22470,N_14365,N_17610);
nand U22471 (N_22471,N_17929,N_15482);
and U22472 (N_22472,N_15250,N_16922);
nand U22473 (N_22473,N_18475,N_13663);
or U22474 (N_22474,N_17950,N_14772);
and U22475 (N_22475,N_16422,N_15537);
or U22476 (N_22476,N_15102,N_15749);
nand U22477 (N_22477,N_17460,N_15818);
nand U22478 (N_22478,N_13568,N_14343);
xor U22479 (N_22479,N_12660,N_15120);
or U22480 (N_22480,N_17880,N_13521);
nand U22481 (N_22481,N_12789,N_15686);
xnor U22482 (N_22482,N_15023,N_15104);
xor U22483 (N_22483,N_12828,N_14723);
or U22484 (N_22484,N_16867,N_13201);
nand U22485 (N_22485,N_14716,N_15972);
nor U22486 (N_22486,N_17983,N_12528);
xnor U22487 (N_22487,N_12559,N_13229);
nor U22488 (N_22488,N_16143,N_15783);
xnor U22489 (N_22489,N_13273,N_15748);
nor U22490 (N_22490,N_17745,N_13022);
and U22491 (N_22491,N_14121,N_16144);
nor U22492 (N_22492,N_16073,N_13553);
xor U22493 (N_22493,N_16079,N_13746);
xor U22494 (N_22494,N_17920,N_16830);
and U22495 (N_22495,N_18300,N_17689);
xnor U22496 (N_22496,N_14913,N_18589);
and U22497 (N_22497,N_14037,N_13205);
and U22498 (N_22498,N_17958,N_15729);
or U22499 (N_22499,N_14751,N_16410);
and U22500 (N_22500,N_13694,N_14097);
nand U22501 (N_22501,N_17686,N_15966);
nand U22502 (N_22502,N_15160,N_18005);
and U22503 (N_22503,N_14803,N_14231);
nand U22504 (N_22504,N_18144,N_13980);
nor U22505 (N_22505,N_18576,N_16321);
nor U22506 (N_22506,N_14835,N_13880);
and U22507 (N_22507,N_16913,N_12972);
xnor U22508 (N_22508,N_13304,N_15667);
xnor U22509 (N_22509,N_18069,N_13778);
nand U22510 (N_22510,N_17270,N_14459);
nor U22511 (N_22511,N_12661,N_16702);
and U22512 (N_22512,N_15610,N_16266);
xor U22513 (N_22513,N_17196,N_14068);
xor U22514 (N_22514,N_17433,N_16526);
or U22515 (N_22515,N_13571,N_18725);
and U22516 (N_22516,N_14029,N_13587);
nand U22517 (N_22517,N_15717,N_15069);
xor U22518 (N_22518,N_15719,N_14282);
and U22519 (N_22519,N_14584,N_16208);
xor U22520 (N_22520,N_14685,N_16721);
xor U22521 (N_22521,N_13359,N_13615);
or U22522 (N_22522,N_13018,N_18590);
or U22523 (N_22523,N_15266,N_13283);
or U22524 (N_22524,N_18125,N_12910);
nor U22525 (N_22525,N_18169,N_14938);
nand U22526 (N_22526,N_13179,N_17828);
and U22527 (N_22527,N_15866,N_15855);
or U22528 (N_22528,N_14013,N_13939);
xor U22529 (N_22529,N_16865,N_14586);
or U22530 (N_22530,N_15533,N_15870);
nor U22531 (N_22531,N_16089,N_18322);
nor U22532 (N_22532,N_16766,N_13728);
nand U22533 (N_22533,N_15629,N_16198);
nand U22534 (N_22534,N_14521,N_12731);
xor U22535 (N_22535,N_18034,N_17393);
and U22536 (N_22536,N_14879,N_14199);
and U22537 (N_22537,N_13630,N_14185);
xor U22538 (N_22538,N_12500,N_18342);
nor U22539 (N_22539,N_18005,N_14021);
and U22540 (N_22540,N_17803,N_14407);
or U22541 (N_22541,N_17840,N_15741);
and U22542 (N_22542,N_14007,N_16470);
nor U22543 (N_22543,N_18170,N_12528);
xor U22544 (N_22544,N_13211,N_18045);
nor U22545 (N_22545,N_12785,N_15163);
nor U22546 (N_22546,N_15605,N_12822);
or U22547 (N_22547,N_16262,N_18303);
xnor U22548 (N_22548,N_13747,N_16728);
and U22549 (N_22549,N_17358,N_14897);
nand U22550 (N_22550,N_16040,N_17744);
nand U22551 (N_22551,N_15074,N_15067);
or U22552 (N_22552,N_16062,N_15869);
nand U22553 (N_22553,N_13875,N_17025);
xor U22554 (N_22554,N_15663,N_18227);
nor U22555 (N_22555,N_16243,N_15345);
nand U22556 (N_22556,N_12778,N_17398);
nand U22557 (N_22557,N_14079,N_15921);
and U22558 (N_22558,N_15128,N_17888);
and U22559 (N_22559,N_18122,N_18520);
xnor U22560 (N_22560,N_15001,N_17410);
or U22561 (N_22561,N_14343,N_16741);
xnor U22562 (N_22562,N_18344,N_15966);
xor U22563 (N_22563,N_13806,N_15994);
xnor U22564 (N_22564,N_14600,N_15884);
nand U22565 (N_22565,N_16655,N_13841);
or U22566 (N_22566,N_17883,N_12820);
and U22567 (N_22567,N_18122,N_15392);
and U22568 (N_22568,N_16277,N_17423);
nand U22569 (N_22569,N_12542,N_14265);
or U22570 (N_22570,N_17272,N_18585);
xnor U22571 (N_22571,N_17390,N_15643);
and U22572 (N_22572,N_14015,N_12957);
or U22573 (N_22573,N_18486,N_15602);
and U22574 (N_22574,N_12939,N_12995);
or U22575 (N_22575,N_12896,N_16093);
or U22576 (N_22576,N_18157,N_17829);
and U22577 (N_22577,N_12982,N_15874);
nor U22578 (N_22578,N_14531,N_16400);
and U22579 (N_22579,N_18086,N_14712);
nor U22580 (N_22580,N_16902,N_14917);
nor U22581 (N_22581,N_13420,N_17123);
xor U22582 (N_22582,N_12512,N_18313);
and U22583 (N_22583,N_13039,N_16347);
xor U22584 (N_22584,N_13083,N_15609);
and U22585 (N_22585,N_18335,N_13940);
and U22586 (N_22586,N_18575,N_14112);
nor U22587 (N_22587,N_13976,N_13005);
xnor U22588 (N_22588,N_14188,N_17298);
or U22589 (N_22589,N_17516,N_13060);
nor U22590 (N_22590,N_15440,N_12504);
xnor U22591 (N_22591,N_17694,N_14772);
nand U22592 (N_22592,N_14827,N_18413);
or U22593 (N_22593,N_15002,N_13499);
or U22594 (N_22594,N_12718,N_15553);
nand U22595 (N_22595,N_13323,N_15854);
nor U22596 (N_22596,N_17212,N_16431);
xnor U22597 (N_22597,N_12598,N_17138);
nand U22598 (N_22598,N_17348,N_17724);
or U22599 (N_22599,N_15931,N_13456);
xor U22600 (N_22600,N_13920,N_18466);
nand U22601 (N_22601,N_13240,N_13196);
or U22602 (N_22602,N_12890,N_17614);
nor U22603 (N_22603,N_13931,N_15055);
and U22604 (N_22604,N_14034,N_12645);
or U22605 (N_22605,N_15197,N_13134);
nand U22606 (N_22606,N_17419,N_13066);
nand U22607 (N_22607,N_16521,N_17608);
nand U22608 (N_22608,N_17158,N_18749);
xor U22609 (N_22609,N_16015,N_17077);
or U22610 (N_22610,N_13917,N_13409);
nand U22611 (N_22611,N_14550,N_15194);
xnor U22612 (N_22612,N_14899,N_13186);
nand U22613 (N_22613,N_18255,N_12813);
xor U22614 (N_22614,N_14430,N_18497);
nor U22615 (N_22615,N_16839,N_16339);
xor U22616 (N_22616,N_16308,N_16186);
and U22617 (N_22617,N_17676,N_13819);
nor U22618 (N_22618,N_14341,N_18109);
nand U22619 (N_22619,N_13613,N_16736);
nand U22620 (N_22620,N_17247,N_16609);
or U22621 (N_22621,N_14712,N_13343);
nor U22622 (N_22622,N_14484,N_14507);
nand U22623 (N_22623,N_16838,N_14713);
or U22624 (N_22624,N_17455,N_16355);
nor U22625 (N_22625,N_14644,N_14642);
nand U22626 (N_22626,N_13976,N_15250);
xor U22627 (N_22627,N_16670,N_13431);
nand U22628 (N_22628,N_15291,N_15165);
xnor U22629 (N_22629,N_12906,N_17582);
xnor U22630 (N_22630,N_16983,N_15809);
nand U22631 (N_22631,N_13452,N_12563);
and U22632 (N_22632,N_13147,N_13287);
nand U22633 (N_22633,N_15190,N_16165);
or U22634 (N_22634,N_16636,N_15711);
xnor U22635 (N_22635,N_13594,N_17248);
and U22636 (N_22636,N_14000,N_15680);
nand U22637 (N_22637,N_15438,N_14229);
or U22638 (N_22638,N_15301,N_14640);
or U22639 (N_22639,N_14065,N_14041);
and U22640 (N_22640,N_17595,N_17254);
xor U22641 (N_22641,N_15079,N_16445);
xor U22642 (N_22642,N_17887,N_15933);
and U22643 (N_22643,N_13772,N_18479);
nand U22644 (N_22644,N_13437,N_15868);
xnor U22645 (N_22645,N_13194,N_13555);
nor U22646 (N_22646,N_15836,N_16969);
xnor U22647 (N_22647,N_15108,N_17287);
and U22648 (N_22648,N_14407,N_18262);
nand U22649 (N_22649,N_16701,N_14646);
xor U22650 (N_22650,N_17120,N_15571);
or U22651 (N_22651,N_13609,N_16868);
and U22652 (N_22652,N_13975,N_14556);
nand U22653 (N_22653,N_16543,N_17155);
nand U22654 (N_22654,N_16480,N_17969);
nand U22655 (N_22655,N_15894,N_15209);
or U22656 (N_22656,N_16156,N_12677);
nor U22657 (N_22657,N_17620,N_14586);
xor U22658 (N_22658,N_17564,N_17995);
xor U22659 (N_22659,N_18185,N_12567);
xnor U22660 (N_22660,N_18657,N_17818);
xor U22661 (N_22661,N_16998,N_17017);
or U22662 (N_22662,N_12895,N_13949);
and U22663 (N_22663,N_15608,N_15245);
xnor U22664 (N_22664,N_15236,N_15696);
nor U22665 (N_22665,N_13996,N_15782);
nand U22666 (N_22666,N_17814,N_12980);
and U22667 (N_22667,N_16316,N_16896);
xnor U22668 (N_22668,N_17411,N_14722);
nand U22669 (N_22669,N_14202,N_15174);
and U22670 (N_22670,N_18348,N_18533);
xnor U22671 (N_22671,N_13129,N_15571);
and U22672 (N_22672,N_16663,N_13373);
nor U22673 (N_22673,N_18708,N_17679);
nand U22674 (N_22674,N_15376,N_17536);
nand U22675 (N_22675,N_14824,N_13281);
or U22676 (N_22676,N_14552,N_17365);
or U22677 (N_22677,N_13924,N_13901);
nand U22678 (N_22678,N_16494,N_17877);
nor U22679 (N_22679,N_15890,N_12925);
nand U22680 (N_22680,N_14664,N_16755);
and U22681 (N_22681,N_18352,N_14836);
nor U22682 (N_22682,N_14030,N_15811);
and U22683 (N_22683,N_16115,N_14413);
and U22684 (N_22684,N_14293,N_14404);
and U22685 (N_22685,N_13691,N_15338);
and U22686 (N_22686,N_17574,N_16572);
nand U22687 (N_22687,N_13226,N_17989);
nand U22688 (N_22688,N_16016,N_16556);
nor U22689 (N_22689,N_18718,N_13013);
or U22690 (N_22690,N_14615,N_13540);
nor U22691 (N_22691,N_15796,N_15686);
nand U22692 (N_22692,N_15457,N_17232);
xnor U22693 (N_22693,N_16574,N_13366);
and U22694 (N_22694,N_12767,N_15293);
xnor U22695 (N_22695,N_16173,N_15814);
xor U22696 (N_22696,N_14325,N_17071);
nor U22697 (N_22697,N_16200,N_12785);
or U22698 (N_22698,N_14155,N_17299);
xnor U22699 (N_22699,N_18475,N_17122);
nor U22700 (N_22700,N_16664,N_15367);
or U22701 (N_22701,N_16451,N_17077);
and U22702 (N_22702,N_14042,N_17605);
xnor U22703 (N_22703,N_12897,N_14738);
and U22704 (N_22704,N_18482,N_16807);
xnor U22705 (N_22705,N_17681,N_18224);
nand U22706 (N_22706,N_15844,N_12768);
or U22707 (N_22707,N_16383,N_16361);
and U22708 (N_22708,N_12595,N_15343);
and U22709 (N_22709,N_14975,N_18032);
nand U22710 (N_22710,N_14102,N_12558);
nor U22711 (N_22711,N_12681,N_17573);
xor U22712 (N_22712,N_16773,N_15435);
xnor U22713 (N_22713,N_17629,N_16641);
nand U22714 (N_22714,N_17274,N_14321);
xor U22715 (N_22715,N_15906,N_15530);
and U22716 (N_22716,N_14443,N_16613);
and U22717 (N_22717,N_13708,N_13011);
xnor U22718 (N_22718,N_15453,N_17474);
or U22719 (N_22719,N_13236,N_14910);
and U22720 (N_22720,N_15852,N_15729);
nand U22721 (N_22721,N_14625,N_18461);
nand U22722 (N_22722,N_14496,N_14610);
and U22723 (N_22723,N_16723,N_12808);
nor U22724 (N_22724,N_15983,N_12875);
nand U22725 (N_22725,N_16463,N_15910);
xnor U22726 (N_22726,N_15684,N_17220);
and U22727 (N_22727,N_15888,N_15513);
and U22728 (N_22728,N_12875,N_18466);
nor U22729 (N_22729,N_12509,N_17049);
nor U22730 (N_22730,N_16312,N_15581);
and U22731 (N_22731,N_12890,N_17193);
and U22732 (N_22732,N_18011,N_12792);
or U22733 (N_22733,N_13037,N_16183);
nor U22734 (N_22734,N_15909,N_15518);
nand U22735 (N_22735,N_17614,N_17787);
nor U22736 (N_22736,N_15054,N_15379);
or U22737 (N_22737,N_12946,N_18167);
and U22738 (N_22738,N_13603,N_16689);
nor U22739 (N_22739,N_17099,N_14487);
and U22740 (N_22740,N_18627,N_18639);
or U22741 (N_22741,N_15149,N_13149);
or U22742 (N_22742,N_14581,N_13961);
xor U22743 (N_22743,N_17236,N_18251);
nand U22744 (N_22744,N_13814,N_16542);
nand U22745 (N_22745,N_13639,N_13230);
nor U22746 (N_22746,N_13403,N_13834);
or U22747 (N_22747,N_12709,N_18697);
and U22748 (N_22748,N_18482,N_12951);
nand U22749 (N_22749,N_15460,N_13563);
and U22750 (N_22750,N_15943,N_13192);
and U22751 (N_22751,N_17963,N_18272);
nand U22752 (N_22752,N_15260,N_15596);
xor U22753 (N_22753,N_18135,N_14011);
and U22754 (N_22754,N_16789,N_13291);
and U22755 (N_22755,N_17460,N_15855);
or U22756 (N_22756,N_14000,N_13843);
nand U22757 (N_22757,N_16741,N_16240);
nor U22758 (N_22758,N_15510,N_14145);
xor U22759 (N_22759,N_15608,N_17253);
nand U22760 (N_22760,N_14464,N_16160);
or U22761 (N_22761,N_12833,N_16130);
nand U22762 (N_22762,N_16891,N_18731);
nand U22763 (N_22763,N_13381,N_14949);
nor U22764 (N_22764,N_17637,N_16003);
xnor U22765 (N_22765,N_13326,N_16625);
nand U22766 (N_22766,N_13003,N_17053);
and U22767 (N_22767,N_14876,N_17611);
or U22768 (N_22768,N_15198,N_17822);
nor U22769 (N_22769,N_17149,N_14032);
or U22770 (N_22770,N_17367,N_16759);
xor U22771 (N_22771,N_15362,N_18386);
and U22772 (N_22772,N_17226,N_17421);
nor U22773 (N_22773,N_18326,N_13227);
and U22774 (N_22774,N_16284,N_15497);
nand U22775 (N_22775,N_15083,N_18511);
xor U22776 (N_22776,N_13777,N_17606);
and U22777 (N_22777,N_17070,N_15582);
nand U22778 (N_22778,N_13727,N_13613);
nand U22779 (N_22779,N_14129,N_13215);
nand U22780 (N_22780,N_16867,N_13811);
and U22781 (N_22781,N_15788,N_13402);
xor U22782 (N_22782,N_15288,N_18126);
xnor U22783 (N_22783,N_18143,N_15444);
or U22784 (N_22784,N_16356,N_14281);
xnor U22785 (N_22785,N_14006,N_14611);
nand U22786 (N_22786,N_16080,N_18145);
or U22787 (N_22787,N_17950,N_13967);
and U22788 (N_22788,N_14226,N_17403);
nand U22789 (N_22789,N_14569,N_14149);
and U22790 (N_22790,N_18009,N_16464);
xor U22791 (N_22791,N_16834,N_16154);
and U22792 (N_22792,N_14357,N_15078);
or U22793 (N_22793,N_15459,N_17236);
or U22794 (N_22794,N_16209,N_15658);
nor U22795 (N_22795,N_15735,N_13829);
or U22796 (N_22796,N_13176,N_15718);
xnor U22797 (N_22797,N_18177,N_12799);
nor U22798 (N_22798,N_18477,N_16342);
nor U22799 (N_22799,N_17418,N_13383);
or U22800 (N_22800,N_15115,N_14480);
xnor U22801 (N_22801,N_16058,N_17319);
nand U22802 (N_22802,N_18241,N_18736);
xnor U22803 (N_22803,N_16980,N_16413);
or U22804 (N_22804,N_16373,N_18749);
xnor U22805 (N_22805,N_17584,N_13644);
nor U22806 (N_22806,N_12820,N_13362);
or U22807 (N_22807,N_17399,N_14655);
nand U22808 (N_22808,N_18075,N_18122);
nand U22809 (N_22809,N_17006,N_17753);
xnor U22810 (N_22810,N_13188,N_14662);
xor U22811 (N_22811,N_17850,N_14774);
and U22812 (N_22812,N_16136,N_13305);
or U22813 (N_22813,N_15501,N_14159);
xnor U22814 (N_22814,N_16443,N_14586);
or U22815 (N_22815,N_13500,N_13573);
and U22816 (N_22816,N_18272,N_12578);
and U22817 (N_22817,N_14620,N_16408);
xor U22818 (N_22818,N_18520,N_16886);
nor U22819 (N_22819,N_14836,N_13286);
nor U22820 (N_22820,N_16062,N_15855);
xor U22821 (N_22821,N_15590,N_12619);
and U22822 (N_22822,N_14998,N_14373);
nor U22823 (N_22823,N_18247,N_18711);
xor U22824 (N_22824,N_17519,N_13022);
nor U22825 (N_22825,N_16028,N_17988);
nor U22826 (N_22826,N_16678,N_17764);
nor U22827 (N_22827,N_12968,N_16373);
xor U22828 (N_22828,N_13075,N_13605);
nor U22829 (N_22829,N_13664,N_16756);
nand U22830 (N_22830,N_12567,N_15515);
nor U22831 (N_22831,N_17865,N_14742);
nand U22832 (N_22832,N_13549,N_17916);
xor U22833 (N_22833,N_17471,N_16816);
nor U22834 (N_22834,N_18462,N_17014);
nand U22835 (N_22835,N_14519,N_14925);
nand U22836 (N_22836,N_14808,N_13851);
xor U22837 (N_22837,N_15843,N_17843);
nor U22838 (N_22838,N_14318,N_15216);
nor U22839 (N_22839,N_16995,N_13796);
xnor U22840 (N_22840,N_14205,N_17531);
nand U22841 (N_22841,N_14756,N_18656);
or U22842 (N_22842,N_17260,N_13869);
and U22843 (N_22843,N_17610,N_15868);
xor U22844 (N_22844,N_14933,N_14603);
xor U22845 (N_22845,N_16791,N_17072);
xnor U22846 (N_22846,N_15031,N_15379);
nor U22847 (N_22847,N_18707,N_12878);
xnor U22848 (N_22848,N_18673,N_15223);
or U22849 (N_22849,N_14108,N_18206);
nor U22850 (N_22850,N_14957,N_15023);
xor U22851 (N_22851,N_15440,N_18571);
or U22852 (N_22852,N_17268,N_13014);
or U22853 (N_22853,N_18678,N_14866);
nor U22854 (N_22854,N_15269,N_17052);
or U22855 (N_22855,N_18690,N_17609);
xor U22856 (N_22856,N_12572,N_16907);
nor U22857 (N_22857,N_15506,N_14136);
nand U22858 (N_22858,N_16666,N_17741);
xor U22859 (N_22859,N_17206,N_15167);
xnor U22860 (N_22860,N_16575,N_13106);
and U22861 (N_22861,N_15979,N_14100);
nor U22862 (N_22862,N_13217,N_17236);
xnor U22863 (N_22863,N_16866,N_17902);
or U22864 (N_22864,N_18340,N_18299);
or U22865 (N_22865,N_14220,N_13117);
nor U22866 (N_22866,N_13969,N_13067);
xor U22867 (N_22867,N_15246,N_16342);
or U22868 (N_22868,N_18109,N_15515);
and U22869 (N_22869,N_15701,N_12729);
or U22870 (N_22870,N_18594,N_16914);
nor U22871 (N_22871,N_13150,N_15714);
xor U22872 (N_22872,N_13327,N_17938);
and U22873 (N_22873,N_14982,N_15421);
xor U22874 (N_22874,N_14148,N_14028);
or U22875 (N_22875,N_15991,N_14773);
nand U22876 (N_22876,N_13189,N_15156);
and U22877 (N_22877,N_14311,N_14075);
or U22878 (N_22878,N_17457,N_15828);
nor U22879 (N_22879,N_16266,N_18534);
and U22880 (N_22880,N_13910,N_14032);
or U22881 (N_22881,N_17741,N_12787);
or U22882 (N_22882,N_12970,N_12557);
nor U22883 (N_22883,N_16484,N_18730);
nand U22884 (N_22884,N_16267,N_14259);
nor U22885 (N_22885,N_16122,N_13778);
and U22886 (N_22886,N_17307,N_13883);
nor U22887 (N_22887,N_16888,N_13007);
xnor U22888 (N_22888,N_13165,N_17787);
and U22889 (N_22889,N_17195,N_14545);
nor U22890 (N_22890,N_14683,N_18389);
nand U22891 (N_22891,N_16972,N_14398);
or U22892 (N_22892,N_17580,N_16236);
and U22893 (N_22893,N_16604,N_13368);
xnor U22894 (N_22894,N_17064,N_16185);
nor U22895 (N_22895,N_13580,N_17666);
xor U22896 (N_22896,N_18251,N_12892);
nand U22897 (N_22897,N_14686,N_14509);
xnor U22898 (N_22898,N_15024,N_18044);
xor U22899 (N_22899,N_13365,N_12810);
and U22900 (N_22900,N_15443,N_14010);
and U22901 (N_22901,N_14735,N_18381);
and U22902 (N_22902,N_17643,N_16821);
or U22903 (N_22903,N_13336,N_18415);
nor U22904 (N_22904,N_18001,N_16072);
and U22905 (N_22905,N_16858,N_13200);
nor U22906 (N_22906,N_13390,N_13045);
nor U22907 (N_22907,N_12874,N_17244);
nand U22908 (N_22908,N_18141,N_18203);
nand U22909 (N_22909,N_18331,N_18519);
or U22910 (N_22910,N_18145,N_17535);
nor U22911 (N_22911,N_14414,N_16014);
nor U22912 (N_22912,N_18361,N_12611);
xnor U22913 (N_22913,N_14078,N_13785);
or U22914 (N_22914,N_13171,N_16664);
nand U22915 (N_22915,N_14257,N_15038);
or U22916 (N_22916,N_14269,N_16088);
and U22917 (N_22917,N_15676,N_15488);
or U22918 (N_22918,N_12640,N_15383);
or U22919 (N_22919,N_16136,N_18145);
and U22920 (N_22920,N_14636,N_13972);
nand U22921 (N_22921,N_17652,N_17740);
xor U22922 (N_22922,N_13789,N_13954);
and U22923 (N_22923,N_13050,N_14691);
nand U22924 (N_22924,N_17608,N_14040);
nand U22925 (N_22925,N_17763,N_15405);
nand U22926 (N_22926,N_18404,N_14080);
and U22927 (N_22927,N_14064,N_17376);
nand U22928 (N_22928,N_16284,N_17106);
and U22929 (N_22929,N_15879,N_12812);
nand U22930 (N_22930,N_14809,N_15811);
xor U22931 (N_22931,N_13281,N_18145);
nor U22932 (N_22932,N_13805,N_15959);
nor U22933 (N_22933,N_15056,N_15256);
nand U22934 (N_22934,N_16419,N_17671);
or U22935 (N_22935,N_13930,N_16236);
nand U22936 (N_22936,N_16489,N_15004);
nand U22937 (N_22937,N_14965,N_14007);
nand U22938 (N_22938,N_16167,N_16415);
or U22939 (N_22939,N_12800,N_15169);
or U22940 (N_22940,N_17308,N_16664);
nand U22941 (N_22941,N_16257,N_17055);
nor U22942 (N_22942,N_14759,N_15134);
or U22943 (N_22943,N_18343,N_13705);
and U22944 (N_22944,N_14950,N_12536);
nand U22945 (N_22945,N_15895,N_15379);
xor U22946 (N_22946,N_12632,N_13024);
nand U22947 (N_22947,N_16855,N_15434);
nand U22948 (N_22948,N_16400,N_18094);
nor U22949 (N_22949,N_18597,N_12543);
or U22950 (N_22950,N_15519,N_13170);
or U22951 (N_22951,N_13162,N_18470);
nand U22952 (N_22952,N_16136,N_16058);
xor U22953 (N_22953,N_15347,N_12943);
and U22954 (N_22954,N_18472,N_18291);
and U22955 (N_22955,N_17481,N_14744);
xnor U22956 (N_22956,N_18663,N_17953);
nand U22957 (N_22957,N_18348,N_13660);
xor U22958 (N_22958,N_15294,N_17255);
and U22959 (N_22959,N_17182,N_18406);
nor U22960 (N_22960,N_15259,N_16815);
and U22961 (N_22961,N_15738,N_12958);
or U22962 (N_22962,N_18067,N_18026);
xnor U22963 (N_22963,N_17671,N_16799);
or U22964 (N_22964,N_18395,N_15700);
xnor U22965 (N_22965,N_15658,N_14064);
nand U22966 (N_22966,N_18660,N_13884);
or U22967 (N_22967,N_14102,N_15017);
nand U22968 (N_22968,N_15557,N_16971);
nor U22969 (N_22969,N_14318,N_14417);
xnor U22970 (N_22970,N_12618,N_12949);
or U22971 (N_22971,N_12524,N_16089);
nor U22972 (N_22972,N_18419,N_17929);
and U22973 (N_22973,N_18009,N_16146);
and U22974 (N_22974,N_17039,N_14693);
and U22975 (N_22975,N_17202,N_15982);
nand U22976 (N_22976,N_16584,N_13088);
or U22977 (N_22977,N_14629,N_15802);
nand U22978 (N_22978,N_13234,N_13338);
nand U22979 (N_22979,N_13672,N_15088);
and U22980 (N_22980,N_15422,N_17294);
and U22981 (N_22981,N_16455,N_15976);
and U22982 (N_22982,N_14028,N_18051);
and U22983 (N_22983,N_14933,N_15325);
and U22984 (N_22984,N_16380,N_14290);
nand U22985 (N_22985,N_14996,N_16007);
nor U22986 (N_22986,N_13875,N_15923);
xnor U22987 (N_22987,N_15194,N_15332);
or U22988 (N_22988,N_17292,N_12504);
or U22989 (N_22989,N_14278,N_16905);
xor U22990 (N_22990,N_16793,N_16578);
or U22991 (N_22991,N_15572,N_15808);
xor U22992 (N_22992,N_15260,N_12894);
nor U22993 (N_22993,N_18355,N_14047);
or U22994 (N_22994,N_12605,N_14811);
nand U22995 (N_22995,N_14132,N_12709);
or U22996 (N_22996,N_13728,N_15614);
or U22997 (N_22997,N_15220,N_16753);
nand U22998 (N_22998,N_15476,N_15413);
and U22999 (N_22999,N_12792,N_16892);
or U23000 (N_23000,N_16649,N_16965);
xnor U23001 (N_23001,N_14881,N_16605);
and U23002 (N_23002,N_16227,N_18589);
xnor U23003 (N_23003,N_14689,N_15728);
or U23004 (N_23004,N_15777,N_17997);
or U23005 (N_23005,N_15102,N_14455);
nand U23006 (N_23006,N_16777,N_12520);
nand U23007 (N_23007,N_15193,N_18147);
xor U23008 (N_23008,N_13243,N_15180);
nand U23009 (N_23009,N_16152,N_17448);
nor U23010 (N_23010,N_17402,N_14850);
or U23011 (N_23011,N_16710,N_15651);
or U23012 (N_23012,N_13619,N_16156);
xnor U23013 (N_23013,N_13417,N_13984);
and U23014 (N_23014,N_15315,N_17125);
nor U23015 (N_23015,N_15757,N_15128);
nand U23016 (N_23016,N_15173,N_16144);
or U23017 (N_23017,N_13477,N_15395);
and U23018 (N_23018,N_18616,N_14043);
nor U23019 (N_23019,N_16166,N_17988);
xor U23020 (N_23020,N_12583,N_14919);
or U23021 (N_23021,N_12512,N_15389);
nand U23022 (N_23022,N_15629,N_13646);
xor U23023 (N_23023,N_17306,N_17292);
nand U23024 (N_23024,N_13612,N_15348);
xnor U23025 (N_23025,N_17646,N_13211);
or U23026 (N_23026,N_16117,N_18682);
or U23027 (N_23027,N_16799,N_15704);
and U23028 (N_23028,N_17160,N_17612);
nor U23029 (N_23029,N_15436,N_17287);
nor U23030 (N_23030,N_13632,N_12921);
xnor U23031 (N_23031,N_12758,N_17006);
or U23032 (N_23032,N_17752,N_17429);
xor U23033 (N_23033,N_13945,N_15941);
and U23034 (N_23034,N_17184,N_14202);
or U23035 (N_23035,N_15785,N_12675);
nand U23036 (N_23036,N_13875,N_14774);
xor U23037 (N_23037,N_13935,N_13754);
xor U23038 (N_23038,N_18279,N_18299);
or U23039 (N_23039,N_18369,N_18099);
nand U23040 (N_23040,N_17387,N_13111);
xor U23041 (N_23041,N_18591,N_12960);
and U23042 (N_23042,N_18020,N_18093);
or U23043 (N_23043,N_17754,N_18545);
xnor U23044 (N_23044,N_18676,N_16871);
nor U23045 (N_23045,N_13551,N_17339);
and U23046 (N_23046,N_17381,N_16440);
or U23047 (N_23047,N_15803,N_18699);
and U23048 (N_23048,N_17771,N_14554);
or U23049 (N_23049,N_17537,N_18674);
xnor U23050 (N_23050,N_16341,N_17625);
and U23051 (N_23051,N_16018,N_13687);
nor U23052 (N_23052,N_15227,N_15721);
and U23053 (N_23053,N_16834,N_12882);
xor U23054 (N_23054,N_13700,N_17214);
nand U23055 (N_23055,N_12541,N_14760);
nor U23056 (N_23056,N_15375,N_14110);
xor U23057 (N_23057,N_17843,N_13514);
or U23058 (N_23058,N_16163,N_15578);
nor U23059 (N_23059,N_13191,N_16976);
nor U23060 (N_23060,N_15995,N_15739);
nand U23061 (N_23061,N_17769,N_12773);
xnor U23062 (N_23062,N_16229,N_16588);
nand U23063 (N_23063,N_18635,N_18128);
and U23064 (N_23064,N_18608,N_18087);
or U23065 (N_23065,N_16697,N_17356);
and U23066 (N_23066,N_13818,N_14653);
and U23067 (N_23067,N_14185,N_14301);
and U23068 (N_23068,N_12821,N_15384);
or U23069 (N_23069,N_15806,N_14113);
nor U23070 (N_23070,N_15776,N_17620);
xor U23071 (N_23071,N_16528,N_14777);
or U23072 (N_23072,N_16187,N_15752);
or U23073 (N_23073,N_13519,N_16267);
and U23074 (N_23074,N_16013,N_15232);
xor U23075 (N_23075,N_18696,N_14303);
nand U23076 (N_23076,N_13861,N_17340);
xor U23077 (N_23077,N_14280,N_14835);
and U23078 (N_23078,N_13395,N_16287);
or U23079 (N_23079,N_16586,N_13445);
and U23080 (N_23080,N_13525,N_14855);
nand U23081 (N_23081,N_17898,N_12861);
nor U23082 (N_23082,N_13011,N_13123);
xnor U23083 (N_23083,N_13206,N_14722);
nand U23084 (N_23084,N_12634,N_14964);
nor U23085 (N_23085,N_16645,N_14672);
nand U23086 (N_23086,N_16732,N_18078);
xnor U23087 (N_23087,N_16015,N_18236);
xnor U23088 (N_23088,N_12662,N_14840);
or U23089 (N_23089,N_14189,N_12716);
xor U23090 (N_23090,N_15225,N_18646);
and U23091 (N_23091,N_17749,N_18489);
or U23092 (N_23092,N_12689,N_17793);
or U23093 (N_23093,N_14920,N_17637);
or U23094 (N_23094,N_13865,N_15361);
nor U23095 (N_23095,N_17307,N_15005);
nand U23096 (N_23096,N_17579,N_17841);
nor U23097 (N_23097,N_15432,N_17967);
or U23098 (N_23098,N_16128,N_13349);
and U23099 (N_23099,N_14490,N_12672);
or U23100 (N_23100,N_13262,N_13823);
or U23101 (N_23101,N_17255,N_15358);
nand U23102 (N_23102,N_17284,N_16620);
xor U23103 (N_23103,N_14858,N_16989);
nor U23104 (N_23104,N_12574,N_14986);
and U23105 (N_23105,N_15502,N_13975);
nand U23106 (N_23106,N_15117,N_13957);
nor U23107 (N_23107,N_13611,N_16620);
and U23108 (N_23108,N_13759,N_16221);
nand U23109 (N_23109,N_14043,N_13452);
xor U23110 (N_23110,N_13745,N_13660);
nor U23111 (N_23111,N_18280,N_14069);
or U23112 (N_23112,N_17814,N_17961);
and U23113 (N_23113,N_15714,N_14423);
nand U23114 (N_23114,N_17201,N_15222);
or U23115 (N_23115,N_18024,N_15092);
and U23116 (N_23116,N_14502,N_16268);
nor U23117 (N_23117,N_18321,N_17173);
xor U23118 (N_23118,N_17816,N_15573);
nor U23119 (N_23119,N_16211,N_14383);
and U23120 (N_23120,N_17196,N_17254);
nor U23121 (N_23121,N_15984,N_15356);
and U23122 (N_23122,N_17834,N_15541);
and U23123 (N_23123,N_17506,N_14768);
and U23124 (N_23124,N_18250,N_12984);
nand U23125 (N_23125,N_16966,N_12953);
xor U23126 (N_23126,N_12952,N_17374);
and U23127 (N_23127,N_15447,N_13573);
xnor U23128 (N_23128,N_14312,N_17547);
or U23129 (N_23129,N_15634,N_18639);
or U23130 (N_23130,N_16992,N_14273);
xor U23131 (N_23131,N_13678,N_15351);
and U23132 (N_23132,N_12949,N_12981);
nand U23133 (N_23133,N_18080,N_16167);
xnor U23134 (N_23134,N_17404,N_16630);
or U23135 (N_23135,N_16640,N_15817);
nor U23136 (N_23136,N_18737,N_18045);
or U23137 (N_23137,N_17763,N_13414);
nand U23138 (N_23138,N_15235,N_14620);
nand U23139 (N_23139,N_13096,N_17537);
nor U23140 (N_23140,N_16254,N_18418);
xor U23141 (N_23141,N_18149,N_13024);
nor U23142 (N_23142,N_16639,N_16641);
or U23143 (N_23143,N_13488,N_16151);
and U23144 (N_23144,N_13751,N_13346);
nand U23145 (N_23145,N_16877,N_16595);
nand U23146 (N_23146,N_15581,N_15846);
nor U23147 (N_23147,N_13993,N_12996);
and U23148 (N_23148,N_18293,N_13101);
xor U23149 (N_23149,N_13178,N_16177);
and U23150 (N_23150,N_17993,N_15193);
xnor U23151 (N_23151,N_17872,N_16504);
nand U23152 (N_23152,N_18338,N_16803);
nor U23153 (N_23153,N_17752,N_14130);
nand U23154 (N_23154,N_16146,N_13259);
or U23155 (N_23155,N_15345,N_16540);
or U23156 (N_23156,N_17037,N_15647);
or U23157 (N_23157,N_16624,N_13526);
or U23158 (N_23158,N_14005,N_16910);
nor U23159 (N_23159,N_15143,N_16386);
nand U23160 (N_23160,N_16026,N_12623);
and U23161 (N_23161,N_14452,N_16785);
xor U23162 (N_23162,N_16294,N_13441);
or U23163 (N_23163,N_14297,N_13268);
or U23164 (N_23164,N_17128,N_14088);
xnor U23165 (N_23165,N_17438,N_13775);
xor U23166 (N_23166,N_12528,N_17123);
and U23167 (N_23167,N_18690,N_15390);
nand U23168 (N_23168,N_18672,N_13745);
nand U23169 (N_23169,N_12843,N_18661);
nor U23170 (N_23170,N_17420,N_17377);
or U23171 (N_23171,N_14087,N_17062);
nand U23172 (N_23172,N_14215,N_13318);
nand U23173 (N_23173,N_13472,N_12684);
and U23174 (N_23174,N_13919,N_12770);
nor U23175 (N_23175,N_15786,N_17517);
nor U23176 (N_23176,N_14424,N_13944);
nor U23177 (N_23177,N_13833,N_14422);
and U23178 (N_23178,N_12917,N_15662);
nor U23179 (N_23179,N_13887,N_13984);
and U23180 (N_23180,N_13289,N_16110);
nand U23181 (N_23181,N_14329,N_17864);
xor U23182 (N_23182,N_16991,N_18635);
nand U23183 (N_23183,N_17551,N_14290);
or U23184 (N_23184,N_15329,N_16019);
nand U23185 (N_23185,N_18618,N_16711);
nand U23186 (N_23186,N_14269,N_16695);
or U23187 (N_23187,N_17762,N_14759);
or U23188 (N_23188,N_15144,N_18367);
nor U23189 (N_23189,N_17168,N_15549);
and U23190 (N_23190,N_13930,N_18152);
nand U23191 (N_23191,N_15169,N_18732);
and U23192 (N_23192,N_17173,N_17938);
nor U23193 (N_23193,N_16897,N_14508);
nand U23194 (N_23194,N_18483,N_12833);
nand U23195 (N_23195,N_18619,N_17293);
xnor U23196 (N_23196,N_18668,N_16859);
or U23197 (N_23197,N_14772,N_13727);
and U23198 (N_23198,N_13363,N_15001);
and U23199 (N_23199,N_12920,N_14776);
and U23200 (N_23200,N_12925,N_15511);
and U23201 (N_23201,N_15634,N_12616);
nand U23202 (N_23202,N_14605,N_15922);
nor U23203 (N_23203,N_16715,N_14368);
xor U23204 (N_23204,N_17687,N_17166);
nand U23205 (N_23205,N_18221,N_16745);
or U23206 (N_23206,N_17009,N_18474);
and U23207 (N_23207,N_14266,N_13954);
and U23208 (N_23208,N_14047,N_14108);
xnor U23209 (N_23209,N_14837,N_16457);
and U23210 (N_23210,N_14459,N_13718);
nand U23211 (N_23211,N_17709,N_12706);
nor U23212 (N_23212,N_15146,N_15631);
nor U23213 (N_23213,N_17871,N_13723);
nor U23214 (N_23214,N_18125,N_17446);
or U23215 (N_23215,N_12765,N_15695);
xnor U23216 (N_23216,N_17093,N_14363);
xor U23217 (N_23217,N_18324,N_17740);
and U23218 (N_23218,N_18287,N_17307);
nand U23219 (N_23219,N_15598,N_13045);
nor U23220 (N_23220,N_13350,N_13785);
and U23221 (N_23221,N_17384,N_13781);
and U23222 (N_23222,N_17025,N_13969);
or U23223 (N_23223,N_13281,N_14426);
nand U23224 (N_23224,N_15988,N_13801);
nand U23225 (N_23225,N_17373,N_16991);
nand U23226 (N_23226,N_16454,N_16216);
nand U23227 (N_23227,N_15880,N_12812);
nand U23228 (N_23228,N_14039,N_13816);
nor U23229 (N_23229,N_16449,N_16434);
and U23230 (N_23230,N_15915,N_14407);
nand U23231 (N_23231,N_13758,N_17580);
nand U23232 (N_23232,N_14190,N_15616);
nor U23233 (N_23233,N_17268,N_14619);
nand U23234 (N_23234,N_13050,N_14906);
or U23235 (N_23235,N_16810,N_16441);
and U23236 (N_23236,N_13551,N_18089);
nor U23237 (N_23237,N_13077,N_15277);
or U23238 (N_23238,N_15833,N_13553);
or U23239 (N_23239,N_17136,N_17707);
or U23240 (N_23240,N_17908,N_17088);
nor U23241 (N_23241,N_16093,N_16640);
nor U23242 (N_23242,N_18252,N_14417);
xor U23243 (N_23243,N_17533,N_13558);
nor U23244 (N_23244,N_18296,N_15016);
xor U23245 (N_23245,N_12653,N_14168);
xor U23246 (N_23246,N_16427,N_15496);
nor U23247 (N_23247,N_12938,N_18552);
xor U23248 (N_23248,N_17146,N_18290);
xor U23249 (N_23249,N_15595,N_15738);
nor U23250 (N_23250,N_17835,N_13639);
and U23251 (N_23251,N_14656,N_15333);
xor U23252 (N_23252,N_16584,N_16355);
or U23253 (N_23253,N_15616,N_17364);
or U23254 (N_23254,N_15115,N_16287);
xnor U23255 (N_23255,N_15166,N_18009);
nand U23256 (N_23256,N_18176,N_18150);
nand U23257 (N_23257,N_15501,N_15554);
and U23258 (N_23258,N_12580,N_12749);
and U23259 (N_23259,N_14246,N_13737);
nor U23260 (N_23260,N_16986,N_16165);
xnor U23261 (N_23261,N_13390,N_18253);
and U23262 (N_23262,N_16544,N_15174);
nand U23263 (N_23263,N_17108,N_17556);
or U23264 (N_23264,N_16052,N_17774);
or U23265 (N_23265,N_15478,N_13349);
xnor U23266 (N_23266,N_14531,N_18245);
nand U23267 (N_23267,N_17640,N_13360);
and U23268 (N_23268,N_15392,N_14818);
nand U23269 (N_23269,N_13531,N_16369);
nand U23270 (N_23270,N_17030,N_12756);
and U23271 (N_23271,N_17952,N_18724);
and U23272 (N_23272,N_16076,N_14356);
and U23273 (N_23273,N_15581,N_17516);
xnor U23274 (N_23274,N_18530,N_17119);
nand U23275 (N_23275,N_16825,N_15705);
or U23276 (N_23276,N_13387,N_15243);
or U23277 (N_23277,N_12745,N_16850);
nor U23278 (N_23278,N_13092,N_13043);
nor U23279 (N_23279,N_16025,N_16409);
nor U23280 (N_23280,N_17177,N_18298);
xnor U23281 (N_23281,N_14336,N_16362);
nand U23282 (N_23282,N_14596,N_18309);
or U23283 (N_23283,N_15373,N_17390);
and U23284 (N_23284,N_17599,N_17472);
nand U23285 (N_23285,N_15655,N_15740);
nand U23286 (N_23286,N_17338,N_15728);
or U23287 (N_23287,N_12527,N_14062);
nor U23288 (N_23288,N_14309,N_15758);
xor U23289 (N_23289,N_13417,N_18575);
nand U23290 (N_23290,N_14751,N_16869);
nor U23291 (N_23291,N_17647,N_17937);
or U23292 (N_23292,N_15353,N_15313);
or U23293 (N_23293,N_16369,N_15954);
nand U23294 (N_23294,N_16999,N_14024);
nor U23295 (N_23295,N_17330,N_17372);
nor U23296 (N_23296,N_13124,N_14284);
nand U23297 (N_23297,N_13221,N_14332);
nand U23298 (N_23298,N_16768,N_17671);
or U23299 (N_23299,N_17699,N_16581);
xnor U23300 (N_23300,N_14872,N_18160);
and U23301 (N_23301,N_18506,N_15742);
xnor U23302 (N_23302,N_18445,N_16094);
nand U23303 (N_23303,N_15489,N_12791);
nand U23304 (N_23304,N_16871,N_17102);
nor U23305 (N_23305,N_18700,N_15309);
nand U23306 (N_23306,N_13931,N_15153);
nand U23307 (N_23307,N_16012,N_13678);
nand U23308 (N_23308,N_16413,N_15411);
xnor U23309 (N_23309,N_13043,N_16171);
and U23310 (N_23310,N_16529,N_18501);
nand U23311 (N_23311,N_16269,N_14095);
nor U23312 (N_23312,N_17335,N_16780);
or U23313 (N_23313,N_17799,N_17254);
xnor U23314 (N_23314,N_18211,N_15840);
xnor U23315 (N_23315,N_15511,N_15189);
nand U23316 (N_23316,N_14732,N_17665);
nand U23317 (N_23317,N_15629,N_18481);
and U23318 (N_23318,N_12904,N_17474);
xnor U23319 (N_23319,N_13569,N_17355);
or U23320 (N_23320,N_14154,N_17834);
nor U23321 (N_23321,N_16504,N_14265);
and U23322 (N_23322,N_18332,N_15407);
or U23323 (N_23323,N_18111,N_16472);
or U23324 (N_23324,N_12792,N_17472);
and U23325 (N_23325,N_13110,N_15574);
nand U23326 (N_23326,N_16457,N_16149);
nand U23327 (N_23327,N_14080,N_12523);
and U23328 (N_23328,N_13119,N_16027);
nor U23329 (N_23329,N_16561,N_13812);
nor U23330 (N_23330,N_17751,N_14372);
and U23331 (N_23331,N_16933,N_16032);
or U23332 (N_23332,N_13448,N_13532);
nor U23333 (N_23333,N_13052,N_15079);
or U23334 (N_23334,N_17971,N_14521);
or U23335 (N_23335,N_13763,N_18388);
and U23336 (N_23336,N_15294,N_17574);
and U23337 (N_23337,N_17764,N_16827);
nor U23338 (N_23338,N_18190,N_16928);
and U23339 (N_23339,N_13923,N_16095);
xor U23340 (N_23340,N_12798,N_13217);
nor U23341 (N_23341,N_15559,N_14277);
nand U23342 (N_23342,N_18260,N_16963);
nor U23343 (N_23343,N_17269,N_17605);
nand U23344 (N_23344,N_16891,N_14247);
nand U23345 (N_23345,N_12827,N_17347);
or U23346 (N_23346,N_13867,N_16662);
nor U23347 (N_23347,N_13139,N_18459);
xor U23348 (N_23348,N_14691,N_14047);
or U23349 (N_23349,N_18024,N_14353);
and U23350 (N_23350,N_16173,N_18182);
xnor U23351 (N_23351,N_13469,N_15958);
or U23352 (N_23352,N_15039,N_15151);
nor U23353 (N_23353,N_12510,N_16667);
nand U23354 (N_23354,N_17145,N_16011);
xor U23355 (N_23355,N_17407,N_13330);
and U23356 (N_23356,N_18531,N_14182);
and U23357 (N_23357,N_13791,N_13411);
xnor U23358 (N_23358,N_18122,N_17380);
xor U23359 (N_23359,N_17858,N_13621);
nor U23360 (N_23360,N_13578,N_17295);
xor U23361 (N_23361,N_18597,N_15486);
nor U23362 (N_23362,N_13735,N_16982);
and U23363 (N_23363,N_15083,N_12946);
nand U23364 (N_23364,N_17366,N_17495);
xnor U23365 (N_23365,N_15019,N_12879);
nor U23366 (N_23366,N_15669,N_17951);
xor U23367 (N_23367,N_15076,N_18366);
or U23368 (N_23368,N_14764,N_13835);
or U23369 (N_23369,N_13799,N_17066);
nor U23370 (N_23370,N_13440,N_16201);
nand U23371 (N_23371,N_15219,N_12859);
xor U23372 (N_23372,N_17746,N_15945);
nor U23373 (N_23373,N_16599,N_13409);
nor U23374 (N_23374,N_13135,N_15154);
and U23375 (N_23375,N_16633,N_14020);
xor U23376 (N_23376,N_15012,N_15139);
nand U23377 (N_23377,N_17406,N_18154);
nand U23378 (N_23378,N_16123,N_14982);
nor U23379 (N_23379,N_14477,N_17804);
and U23380 (N_23380,N_15016,N_13395);
nand U23381 (N_23381,N_16429,N_15254);
nor U23382 (N_23382,N_17990,N_13822);
xor U23383 (N_23383,N_18076,N_13237);
or U23384 (N_23384,N_16082,N_17366);
nor U23385 (N_23385,N_18270,N_13347);
and U23386 (N_23386,N_14926,N_17850);
nor U23387 (N_23387,N_15507,N_15269);
nand U23388 (N_23388,N_15299,N_15825);
and U23389 (N_23389,N_18171,N_18246);
nor U23390 (N_23390,N_13171,N_15773);
nand U23391 (N_23391,N_15498,N_15696);
xnor U23392 (N_23392,N_16116,N_13819);
nor U23393 (N_23393,N_18195,N_18169);
and U23394 (N_23394,N_18241,N_18639);
nand U23395 (N_23395,N_17234,N_16502);
nand U23396 (N_23396,N_14864,N_16837);
nand U23397 (N_23397,N_16232,N_15845);
nand U23398 (N_23398,N_17117,N_14896);
and U23399 (N_23399,N_14329,N_15230);
nand U23400 (N_23400,N_15736,N_16927);
nor U23401 (N_23401,N_15723,N_14035);
nand U23402 (N_23402,N_13757,N_16294);
or U23403 (N_23403,N_13660,N_17925);
xnor U23404 (N_23404,N_15537,N_16259);
nand U23405 (N_23405,N_14126,N_18174);
or U23406 (N_23406,N_14702,N_16562);
xor U23407 (N_23407,N_12603,N_14371);
or U23408 (N_23408,N_13939,N_17300);
xnor U23409 (N_23409,N_16693,N_14210);
or U23410 (N_23410,N_16075,N_17313);
or U23411 (N_23411,N_18016,N_12946);
or U23412 (N_23412,N_15980,N_18638);
xor U23413 (N_23413,N_18658,N_13637);
xor U23414 (N_23414,N_14684,N_16912);
xnor U23415 (N_23415,N_14047,N_16261);
nand U23416 (N_23416,N_17144,N_17546);
nor U23417 (N_23417,N_17753,N_13002);
nor U23418 (N_23418,N_17734,N_13531);
and U23419 (N_23419,N_14637,N_14451);
or U23420 (N_23420,N_17945,N_16078);
nor U23421 (N_23421,N_14331,N_15070);
nand U23422 (N_23422,N_17705,N_14667);
nand U23423 (N_23423,N_17997,N_13719);
nand U23424 (N_23424,N_13302,N_15118);
xor U23425 (N_23425,N_13814,N_17562);
or U23426 (N_23426,N_13326,N_15538);
xor U23427 (N_23427,N_13204,N_14761);
nand U23428 (N_23428,N_17698,N_18716);
or U23429 (N_23429,N_16701,N_18472);
nand U23430 (N_23430,N_16478,N_13892);
and U23431 (N_23431,N_18528,N_17238);
xor U23432 (N_23432,N_17838,N_16184);
and U23433 (N_23433,N_18201,N_18191);
nor U23434 (N_23434,N_17038,N_14027);
nand U23435 (N_23435,N_16072,N_14252);
nor U23436 (N_23436,N_15658,N_13665);
xnor U23437 (N_23437,N_15736,N_13577);
nand U23438 (N_23438,N_13040,N_16825);
or U23439 (N_23439,N_15528,N_16294);
nor U23440 (N_23440,N_13781,N_17890);
and U23441 (N_23441,N_15602,N_16883);
or U23442 (N_23442,N_17636,N_13991);
and U23443 (N_23443,N_14598,N_17242);
xor U23444 (N_23444,N_13515,N_18088);
xor U23445 (N_23445,N_15482,N_17669);
or U23446 (N_23446,N_16504,N_16563);
nand U23447 (N_23447,N_18550,N_16380);
or U23448 (N_23448,N_14279,N_13878);
nand U23449 (N_23449,N_16363,N_17784);
nor U23450 (N_23450,N_13579,N_15246);
xor U23451 (N_23451,N_17189,N_16086);
xor U23452 (N_23452,N_13686,N_18672);
or U23453 (N_23453,N_18571,N_13507);
and U23454 (N_23454,N_13865,N_13389);
or U23455 (N_23455,N_17340,N_13424);
and U23456 (N_23456,N_17232,N_17171);
or U23457 (N_23457,N_17202,N_18604);
xnor U23458 (N_23458,N_15869,N_17347);
xor U23459 (N_23459,N_18482,N_15394);
nor U23460 (N_23460,N_13003,N_16391);
nand U23461 (N_23461,N_14177,N_14253);
xnor U23462 (N_23462,N_14033,N_12890);
xor U23463 (N_23463,N_18155,N_16464);
nand U23464 (N_23464,N_13678,N_18594);
xor U23465 (N_23465,N_15807,N_16454);
nor U23466 (N_23466,N_17962,N_18465);
nor U23467 (N_23467,N_16727,N_13026);
or U23468 (N_23468,N_18006,N_15574);
nand U23469 (N_23469,N_12795,N_14168);
nand U23470 (N_23470,N_13101,N_14416);
nand U23471 (N_23471,N_15217,N_13410);
xnor U23472 (N_23472,N_14269,N_17839);
or U23473 (N_23473,N_17246,N_14376);
and U23474 (N_23474,N_16735,N_15821);
nor U23475 (N_23475,N_15138,N_16701);
nand U23476 (N_23476,N_16731,N_16958);
nor U23477 (N_23477,N_12581,N_15226);
and U23478 (N_23478,N_15068,N_16464);
and U23479 (N_23479,N_12604,N_16532);
nand U23480 (N_23480,N_13788,N_16527);
nor U23481 (N_23481,N_13132,N_15576);
or U23482 (N_23482,N_15056,N_13493);
nor U23483 (N_23483,N_15181,N_13327);
nor U23484 (N_23484,N_13936,N_18294);
nand U23485 (N_23485,N_13446,N_18450);
nand U23486 (N_23486,N_16244,N_17208);
or U23487 (N_23487,N_13429,N_13526);
or U23488 (N_23488,N_14067,N_12651);
xnor U23489 (N_23489,N_15761,N_18519);
and U23490 (N_23490,N_14351,N_18492);
nand U23491 (N_23491,N_17879,N_15883);
xor U23492 (N_23492,N_14063,N_16662);
nor U23493 (N_23493,N_17245,N_14262);
xnor U23494 (N_23494,N_14971,N_17311);
nor U23495 (N_23495,N_12763,N_15252);
xnor U23496 (N_23496,N_17958,N_18274);
or U23497 (N_23497,N_17179,N_15500);
and U23498 (N_23498,N_13268,N_16440);
xor U23499 (N_23499,N_14156,N_17280);
and U23500 (N_23500,N_18085,N_16300);
nor U23501 (N_23501,N_14227,N_12953);
or U23502 (N_23502,N_13877,N_13099);
nand U23503 (N_23503,N_17287,N_12781);
or U23504 (N_23504,N_14697,N_15107);
nor U23505 (N_23505,N_15850,N_18640);
xor U23506 (N_23506,N_16572,N_18427);
nand U23507 (N_23507,N_14010,N_15650);
nand U23508 (N_23508,N_15159,N_15547);
nand U23509 (N_23509,N_13378,N_16480);
and U23510 (N_23510,N_13513,N_18008);
nand U23511 (N_23511,N_14273,N_17113);
xor U23512 (N_23512,N_16281,N_16413);
or U23513 (N_23513,N_18533,N_16238);
and U23514 (N_23514,N_17393,N_13866);
and U23515 (N_23515,N_14332,N_13710);
nor U23516 (N_23516,N_16879,N_18209);
nand U23517 (N_23517,N_14698,N_12871);
or U23518 (N_23518,N_12805,N_13684);
or U23519 (N_23519,N_13262,N_14174);
nand U23520 (N_23520,N_17882,N_18380);
or U23521 (N_23521,N_14910,N_16319);
and U23522 (N_23522,N_17929,N_18573);
or U23523 (N_23523,N_17291,N_15695);
nor U23524 (N_23524,N_13841,N_15571);
nor U23525 (N_23525,N_17741,N_14331);
nand U23526 (N_23526,N_14876,N_15392);
xnor U23527 (N_23527,N_13013,N_13540);
nor U23528 (N_23528,N_14017,N_15290);
nand U23529 (N_23529,N_17522,N_17979);
and U23530 (N_23530,N_17116,N_16518);
xor U23531 (N_23531,N_15807,N_16081);
and U23532 (N_23532,N_18421,N_13542);
xor U23533 (N_23533,N_16394,N_16744);
nor U23534 (N_23534,N_13876,N_13820);
or U23535 (N_23535,N_13963,N_14035);
or U23536 (N_23536,N_18588,N_18494);
nor U23537 (N_23537,N_18633,N_18588);
xnor U23538 (N_23538,N_16112,N_13601);
nor U23539 (N_23539,N_18200,N_16068);
xnor U23540 (N_23540,N_17687,N_16979);
nor U23541 (N_23541,N_13933,N_13918);
nor U23542 (N_23542,N_13984,N_14315);
nor U23543 (N_23543,N_17788,N_16036);
or U23544 (N_23544,N_17574,N_12707);
and U23545 (N_23545,N_14543,N_15171);
xor U23546 (N_23546,N_14186,N_17410);
or U23547 (N_23547,N_12701,N_14243);
nor U23548 (N_23548,N_13133,N_15722);
xor U23549 (N_23549,N_15688,N_17886);
xor U23550 (N_23550,N_17361,N_17367);
xor U23551 (N_23551,N_14656,N_18413);
nor U23552 (N_23552,N_13666,N_12860);
or U23553 (N_23553,N_14878,N_17406);
or U23554 (N_23554,N_16051,N_16758);
xnor U23555 (N_23555,N_16060,N_16144);
nand U23556 (N_23556,N_16836,N_16548);
or U23557 (N_23557,N_14267,N_13580);
and U23558 (N_23558,N_15962,N_13356);
xor U23559 (N_23559,N_16074,N_16659);
nand U23560 (N_23560,N_15024,N_18372);
nor U23561 (N_23561,N_13434,N_14074);
nor U23562 (N_23562,N_18467,N_12828);
nor U23563 (N_23563,N_15869,N_12514);
nor U23564 (N_23564,N_16189,N_17189);
xor U23565 (N_23565,N_18651,N_16583);
nor U23566 (N_23566,N_16192,N_15694);
nand U23567 (N_23567,N_12650,N_15141);
xnor U23568 (N_23568,N_18416,N_14740);
nand U23569 (N_23569,N_16943,N_13662);
and U23570 (N_23570,N_14030,N_18030);
nor U23571 (N_23571,N_16774,N_15133);
xnor U23572 (N_23572,N_18024,N_14665);
nand U23573 (N_23573,N_17506,N_18418);
nand U23574 (N_23574,N_14512,N_14487);
and U23575 (N_23575,N_15019,N_18611);
nor U23576 (N_23576,N_18328,N_15661);
or U23577 (N_23577,N_17748,N_12518);
xnor U23578 (N_23578,N_15015,N_12618);
nand U23579 (N_23579,N_15009,N_15290);
nand U23580 (N_23580,N_14211,N_18393);
or U23581 (N_23581,N_16461,N_16900);
xnor U23582 (N_23582,N_17685,N_17113);
nor U23583 (N_23583,N_14472,N_14300);
and U23584 (N_23584,N_17170,N_16631);
and U23585 (N_23585,N_17092,N_17266);
nand U23586 (N_23586,N_18597,N_13971);
or U23587 (N_23587,N_13280,N_15949);
nor U23588 (N_23588,N_15474,N_14502);
or U23589 (N_23589,N_16984,N_17689);
or U23590 (N_23590,N_14002,N_17426);
or U23591 (N_23591,N_15360,N_17945);
xor U23592 (N_23592,N_15409,N_16997);
or U23593 (N_23593,N_12912,N_17464);
xor U23594 (N_23594,N_17979,N_14730);
xor U23595 (N_23595,N_16918,N_13449);
nor U23596 (N_23596,N_18683,N_15620);
xor U23597 (N_23597,N_13237,N_13007);
nand U23598 (N_23598,N_16113,N_15877);
nand U23599 (N_23599,N_17424,N_18006);
xor U23600 (N_23600,N_13487,N_13850);
or U23601 (N_23601,N_14828,N_15873);
or U23602 (N_23602,N_18300,N_14753);
nor U23603 (N_23603,N_15151,N_13093);
nor U23604 (N_23604,N_15493,N_15787);
and U23605 (N_23605,N_16944,N_18459);
and U23606 (N_23606,N_16142,N_14334);
nor U23607 (N_23607,N_14951,N_13677);
or U23608 (N_23608,N_16269,N_12875);
nor U23609 (N_23609,N_17363,N_12523);
nor U23610 (N_23610,N_17764,N_15648);
xor U23611 (N_23611,N_13637,N_18661);
nand U23612 (N_23612,N_13123,N_12643);
and U23613 (N_23613,N_13824,N_16469);
and U23614 (N_23614,N_16100,N_16827);
nor U23615 (N_23615,N_13608,N_18624);
nor U23616 (N_23616,N_13849,N_16701);
nand U23617 (N_23617,N_18724,N_16864);
nor U23618 (N_23618,N_14219,N_16034);
nand U23619 (N_23619,N_15659,N_14501);
xor U23620 (N_23620,N_14273,N_13825);
nor U23621 (N_23621,N_16501,N_18252);
and U23622 (N_23622,N_12550,N_14032);
nand U23623 (N_23623,N_13990,N_17622);
nor U23624 (N_23624,N_15038,N_14236);
nand U23625 (N_23625,N_18246,N_13425);
and U23626 (N_23626,N_16833,N_18544);
nand U23627 (N_23627,N_18206,N_14940);
xor U23628 (N_23628,N_15276,N_15428);
nand U23629 (N_23629,N_16139,N_12690);
and U23630 (N_23630,N_18260,N_16905);
or U23631 (N_23631,N_16777,N_18574);
and U23632 (N_23632,N_14802,N_15558);
nor U23633 (N_23633,N_12931,N_13436);
nand U23634 (N_23634,N_15787,N_13587);
or U23635 (N_23635,N_16979,N_12818);
xnor U23636 (N_23636,N_16685,N_15996);
and U23637 (N_23637,N_15343,N_12560);
and U23638 (N_23638,N_14221,N_14598);
xor U23639 (N_23639,N_14608,N_17239);
xnor U23640 (N_23640,N_18069,N_18052);
or U23641 (N_23641,N_18245,N_13347);
and U23642 (N_23642,N_14694,N_14471);
and U23643 (N_23643,N_12654,N_16745);
and U23644 (N_23644,N_14840,N_17523);
xor U23645 (N_23645,N_16819,N_13886);
and U23646 (N_23646,N_14055,N_15825);
nand U23647 (N_23647,N_16220,N_15127);
and U23648 (N_23648,N_16263,N_12535);
xnor U23649 (N_23649,N_17805,N_12729);
xnor U23650 (N_23650,N_16122,N_15116);
or U23651 (N_23651,N_15204,N_12529);
xor U23652 (N_23652,N_17551,N_17933);
nand U23653 (N_23653,N_17480,N_16504);
nand U23654 (N_23654,N_17258,N_14294);
nor U23655 (N_23655,N_15919,N_14123);
xnor U23656 (N_23656,N_14773,N_14127);
or U23657 (N_23657,N_13313,N_13192);
nor U23658 (N_23658,N_12694,N_13036);
nor U23659 (N_23659,N_18199,N_18179);
nand U23660 (N_23660,N_18634,N_12601);
nand U23661 (N_23661,N_15563,N_16204);
and U23662 (N_23662,N_13010,N_13055);
xor U23663 (N_23663,N_14792,N_16022);
nand U23664 (N_23664,N_14192,N_18464);
nor U23665 (N_23665,N_16967,N_15317);
nor U23666 (N_23666,N_16627,N_17428);
nor U23667 (N_23667,N_15882,N_16225);
xor U23668 (N_23668,N_18328,N_13531);
xor U23669 (N_23669,N_16069,N_16237);
and U23670 (N_23670,N_13713,N_15967);
nor U23671 (N_23671,N_17722,N_13382);
xnor U23672 (N_23672,N_18090,N_14758);
xor U23673 (N_23673,N_16090,N_13326);
xnor U23674 (N_23674,N_15448,N_14016);
nor U23675 (N_23675,N_13990,N_16162);
nand U23676 (N_23676,N_17233,N_14951);
nand U23677 (N_23677,N_13009,N_17184);
nor U23678 (N_23678,N_16262,N_15942);
nor U23679 (N_23679,N_13350,N_17600);
and U23680 (N_23680,N_15632,N_13850);
nor U23681 (N_23681,N_15661,N_15560);
xor U23682 (N_23682,N_18741,N_16537);
xor U23683 (N_23683,N_17102,N_14627);
nor U23684 (N_23684,N_16434,N_18563);
or U23685 (N_23685,N_13371,N_15606);
xor U23686 (N_23686,N_16517,N_15886);
or U23687 (N_23687,N_18026,N_12809);
and U23688 (N_23688,N_16502,N_14337);
xor U23689 (N_23689,N_15519,N_13043);
xor U23690 (N_23690,N_15332,N_12600);
and U23691 (N_23691,N_17097,N_14931);
and U23692 (N_23692,N_13322,N_13029);
and U23693 (N_23693,N_13312,N_15256);
nand U23694 (N_23694,N_16769,N_13276);
nand U23695 (N_23695,N_16805,N_12665);
and U23696 (N_23696,N_12807,N_17189);
and U23697 (N_23697,N_16795,N_18291);
nand U23698 (N_23698,N_13993,N_16512);
nor U23699 (N_23699,N_15717,N_15130);
and U23700 (N_23700,N_14143,N_14247);
and U23701 (N_23701,N_12628,N_15169);
nor U23702 (N_23702,N_17755,N_18563);
nor U23703 (N_23703,N_17638,N_12532);
nand U23704 (N_23704,N_14693,N_15921);
and U23705 (N_23705,N_18020,N_17232);
or U23706 (N_23706,N_17155,N_14997);
nor U23707 (N_23707,N_16912,N_17229);
nor U23708 (N_23708,N_16563,N_18744);
nand U23709 (N_23709,N_13837,N_13259);
and U23710 (N_23710,N_17511,N_13176);
nand U23711 (N_23711,N_13796,N_18467);
xor U23712 (N_23712,N_15264,N_13855);
or U23713 (N_23713,N_17039,N_16766);
and U23714 (N_23714,N_12872,N_18668);
nand U23715 (N_23715,N_13217,N_17497);
or U23716 (N_23716,N_18010,N_13455);
nor U23717 (N_23717,N_15637,N_13921);
nand U23718 (N_23718,N_12620,N_15911);
or U23719 (N_23719,N_15922,N_12640);
xnor U23720 (N_23720,N_16217,N_13559);
or U23721 (N_23721,N_13221,N_17893);
or U23722 (N_23722,N_16600,N_12671);
or U23723 (N_23723,N_14619,N_12948);
xnor U23724 (N_23724,N_15544,N_15334);
nand U23725 (N_23725,N_16647,N_12763);
and U23726 (N_23726,N_17789,N_18122);
and U23727 (N_23727,N_13809,N_15542);
xor U23728 (N_23728,N_14840,N_16024);
xor U23729 (N_23729,N_17291,N_15920);
and U23730 (N_23730,N_14993,N_17365);
nand U23731 (N_23731,N_16578,N_16237);
and U23732 (N_23732,N_15713,N_12709);
or U23733 (N_23733,N_18472,N_15555);
and U23734 (N_23734,N_18441,N_14764);
nand U23735 (N_23735,N_17358,N_15139);
and U23736 (N_23736,N_17219,N_14580);
or U23737 (N_23737,N_14134,N_15139);
or U23738 (N_23738,N_14012,N_13622);
xor U23739 (N_23739,N_13438,N_15205);
xnor U23740 (N_23740,N_15390,N_18237);
xor U23741 (N_23741,N_17873,N_17591);
nand U23742 (N_23742,N_13379,N_12506);
nand U23743 (N_23743,N_18279,N_15458);
nand U23744 (N_23744,N_13164,N_16324);
nand U23745 (N_23745,N_17654,N_16457);
xor U23746 (N_23746,N_15450,N_16047);
and U23747 (N_23747,N_16979,N_17506);
or U23748 (N_23748,N_16056,N_16696);
nand U23749 (N_23749,N_13515,N_17783);
nor U23750 (N_23750,N_15122,N_13887);
and U23751 (N_23751,N_14962,N_16476);
nor U23752 (N_23752,N_15773,N_18531);
nand U23753 (N_23753,N_14830,N_12542);
xor U23754 (N_23754,N_17016,N_12619);
and U23755 (N_23755,N_13689,N_16096);
nand U23756 (N_23756,N_16096,N_12869);
xnor U23757 (N_23757,N_14764,N_18437);
xnor U23758 (N_23758,N_18070,N_17629);
and U23759 (N_23759,N_16536,N_18333);
and U23760 (N_23760,N_13378,N_18580);
and U23761 (N_23761,N_16894,N_12894);
and U23762 (N_23762,N_16187,N_12693);
or U23763 (N_23763,N_16644,N_18522);
xnor U23764 (N_23764,N_13026,N_17697);
and U23765 (N_23765,N_14708,N_15996);
nor U23766 (N_23766,N_14315,N_18593);
or U23767 (N_23767,N_13086,N_14452);
xor U23768 (N_23768,N_13925,N_17571);
and U23769 (N_23769,N_14780,N_17431);
and U23770 (N_23770,N_15141,N_14785);
or U23771 (N_23771,N_14871,N_15389);
or U23772 (N_23772,N_13756,N_15695);
nor U23773 (N_23773,N_15149,N_15572);
or U23774 (N_23774,N_13798,N_14316);
xnor U23775 (N_23775,N_13191,N_18472);
nor U23776 (N_23776,N_12766,N_14903);
nor U23777 (N_23777,N_18469,N_15436);
and U23778 (N_23778,N_15397,N_13030);
nand U23779 (N_23779,N_14262,N_18375);
nand U23780 (N_23780,N_16589,N_17923);
nor U23781 (N_23781,N_17088,N_16507);
and U23782 (N_23782,N_14427,N_17712);
nand U23783 (N_23783,N_12959,N_15998);
or U23784 (N_23784,N_17579,N_17418);
xor U23785 (N_23785,N_13858,N_18232);
nand U23786 (N_23786,N_13546,N_15902);
nand U23787 (N_23787,N_18049,N_17000);
and U23788 (N_23788,N_14056,N_13817);
nor U23789 (N_23789,N_18712,N_13771);
and U23790 (N_23790,N_17439,N_16856);
xor U23791 (N_23791,N_18229,N_15767);
nand U23792 (N_23792,N_18343,N_12582);
and U23793 (N_23793,N_16285,N_16782);
nand U23794 (N_23794,N_15053,N_13774);
or U23795 (N_23795,N_16952,N_14530);
nor U23796 (N_23796,N_16153,N_14069);
nor U23797 (N_23797,N_15214,N_13053);
and U23798 (N_23798,N_13568,N_16074);
or U23799 (N_23799,N_13657,N_16953);
nor U23800 (N_23800,N_14227,N_14819);
nand U23801 (N_23801,N_17297,N_15585);
xnor U23802 (N_23802,N_14123,N_17075);
and U23803 (N_23803,N_13243,N_17362);
nand U23804 (N_23804,N_12965,N_12759);
and U23805 (N_23805,N_13301,N_18504);
nand U23806 (N_23806,N_16817,N_15247);
xor U23807 (N_23807,N_14395,N_14622);
nand U23808 (N_23808,N_12762,N_15397);
nor U23809 (N_23809,N_17111,N_14409);
and U23810 (N_23810,N_13064,N_15384);
and U23811 (N_23811,N_15606,N_16427);
and U23812 (N_23812,N_16564,N_13671);
nand U23813 (N_23813,N_16571,N_14784);
and U23814 (N_23814,N_13057,N_14093);
or U23815 (N_23815,N_17228,N_17700);
or U23816 (N_23816,N_17338,N_15651);
and U23817 (N_23817,N_16012,N_15031);
xnor U23818 (N_23818,N_13220,N_14983);
xor U23819 (N_23819,N_17048,N_17972);
nand U23820 (N_23820,N_13889,N_13567);
nand U23821 (N_23821,N_15205,N_15037);
or U23822 (N_23822,N_18666,N_14127);
xnor U23823 (N_23823,N_14325,N_14393);
or U23824 (N_23824,N_16264,N_12855);
nand U23825 (N_23825,N_14636,N_13534);
nor U23826 (N_23826,N_16742,N_17451);
xor U23827 (N_23827,N_14561,N_15222);
xor U23828 (N_23828,N_16424,N_16091);
or U23829 (N_23829,N_17801,N_15245);
or U23830 (N_23830,N_12889,N_12771);
xnor U23831 (N_23831,N_18571,N_13387);
nand U23832 (N_23832,N_14592,N_16323);
and U23833 (N_23833,N_13891,N_17369);
and U23834 (N_23834,N_18104,N_18264);
xor U23835 (N_23835,N_17493,N_12994);
nor U23836 (N_23836,N_17195,N_15657);
nand U23837 (N_23837,N_12642,N_14196);
and U23838 (N_23838,N_16840,N_14518);
nor U23839 (N_23839,N_18145,N_16381);
xor U23840 (N_23840,N_17991,N_13242);
or U23841 (N_23841,N_18342,N_17001);
and U23842 (N_23842,N_15898,N_15815);
or U23843 (N_23843,N_12992,N_12828);
or U23844 (N_23844,N_17523,N_18100);
or U23845 (N_23845,N_17014,N_16639);
xor U23846 (N_23846,N_14912,N_16300);
nand U23847 (N_23847,N_17907,N_17974);
xor U23848 (N_23848,N_15659,N_13619);
nand U23849 (N_23849,N_13587,N_12937);
nor U23850 (N_23850,N_17276,N_16225);
and U23851 (N_23851,N_16246,N_16828);
or U23852 (N_23852,N_14180,N_17641);
or U23853 (N_23853,N_14622,N_13826);
nand U23854 (N_23854,N_13692,N_13879);
nor U23855 (N_23855,N_18396,N_16205);
xor U23856 (N_23856,N_15978,N_16825);
and U23857 (N_23857,N_17257,N_18584);
and U23858 (N_23858,N_15189,N_17471);
or U23859 (N_23859,N_15851,N_13927);
nand U23860 (N_23860,N_12596,N_17154);
xnor U23861 (N_23861,N_16889,N_12715);
xnor U23862 (N_23862,N_13857,N_13632);
or U23863 (N_23863,N_17267,N_15305);
or U23864 (N_23864,N_18073,N_16707);
xor U23865 (N_23865,N_13345,N_13903);
xor U23866 (N_23866,N_12820,N_15974);
or U23867 (N_23867,N_12945,N_15222);
or U23868 (N_23868,N_14501,N_17817);
and U23869 (N_23869,N_16052,N_13080);
nor U23870 (N_23870,N_15232,N_13694);
or U23871 (N_23871,N_14773,N_14312);
or U23872 (N_23872,N_16849,N_15247);
and U23873 (N_23873,N_17425,N_13079);
xnor U23874 (N_23874,N_15948,N_13740);
and U23875 (N_23875,N_16117,N_13034);
nor U23876 (N_23876,N_14211,N_17071);
and U23877 (N_23877,N_16344,N_13110);
and U23878 (N_23878,N_12658,N_18622);
nor U23879 (N_23879,N_16025,N_14112);
and U23880 (N_23880,N_15530,N_18510);
nand U23881 (N_23881,N_12913,N_17261);
and U23882 (N_23882,N_14724,N_17271);
xor U23883 (N_23883,N_14603,N_16470);
and U23884 (N_23884,N_16793,N_13026);
nand U23885 (N_23885,N_16498,N_14224);
nor U23886 (N_23886,N_14158,N_15312);
or U23887 (N_23887,N_13377,N_16842);
and U23888 (N_23888,N_15832,N_16581);
xor U23889 (N_23889,N_16327,N_12690);
or U23890 (N_23890,N_12918,N_17551);
nand U23891 (N_23891,N_14191,N_15411);
nand U23892 (N_23892,N_13608,N_13332);
or U23893 (N_23893,N_12816,N_14069);
nor U23894 (N_23894,N_17371,N_13217);
nor U23895 (N_23895,N_17287,N_17301);
xor U23896 (N_23896,N_17971,N_17442);
xnor U23897 (N_23897,N_17967,N_12758);
and U23898 (N_23898,N_15803,N_15539);
xor U23899 (N_23899,N_14082,N_13505);
or U23900 (N_23900,N_12628,N_16348);
nand U23901 (N_23901,N_16802,N_14146);
and U23902 (N_23902,N_18263,N_16514);
or U23903 (N_23903,N_18688,N_16154);
nand U23904 (N_23904,N_13617,N_17729);
nand U23905 (N_23905,N_13639,N_17194);
and U23906 (N_23906,N_17088,N_14444);
xor U23907 (N_23907,N_14499,N_16549);
nor U23908 (N_23908,N_18534,N_12602);
nand U23909 (N_23909,N_13736,N_15013);
or U23910 (N_23910,N_17817,N_16701);
nand U23911 (N_23911,N_18078,N_14903);
nor U23912 (N_23912,N_16369,N_15048);
nand U23913 (N_23913,N_18680,N_17299);
xor U23914 (N_23914,N_17623,N_12800);
and U23915 (N_23915,N_14897,N_18108);
and U23916 (N_23916,N_17445,N_15090);
or U23917 (N_23917,N_13164,N_13152);
and U23918 (N_23918,N_17116,N_18016);
nor U23919 (N_23919,N_15148,N_13369);
or U23920 (N_23920,N_13759,N_15868);
or U23921 (N_23921,N_16246,N_17636);
or U23922 (N_23922,N_16115,N_16096);
nor U23923 (N_23923,N_13545,N_15718);
or U23924 (N_23924,N_15935,N_15952);
nand U23925 (N_23925,N_13414,N_17429);
nor U23926 (N_23926,N_18435,N_18233);
nand U23927 (N_23927,N_16118,N_17075);
nor U23928 (N_23928,N_13772,N_16607);
nor U23929 (N_23929,N_13535,N_17645);
nand U23930 (N_23930,N_13396,N_16894);
or U23931 (N_23931,N_14794,N_14051);
xor U23932 (N_23932,N_16391,N_15383);
xor U23933 (N_23933,N_16586,N_16718);
and U23934 (N_23934,N_16055,N_13073);
nor U23935 (N_23935,N_16132,N_14911);
and U23936 (N_23936,N_17570,N_13870);
nand U23937 (N_23937,N_17357,N_12529);
xor U23938 (N_23938,N_18476,N_12674);
or U23939 (N_23939,N_16172,N_15244);
and U23940 (N_23940,N_14073,N_12757);
and U23941 (N_23941,N_14696,N_13167);
or U23942 (N_23942,N_18464,N_13381);
or U23943 (N_23943,N_12851,N_16895);
nor U23944 (N_23944,N_12693,N_16908);
or U23945 (N_23945,N_15057,N_12888);
and U23946 (N_23946,N_13863,N_13399);
nor U23947 (N_23947,N_15580,N_14394);
nand U23948 (N_23948,N_17765,N_16186);
and U23949 (N_23949,N_16201,N_15170);
and U23950 (N_23950,N_14414,N_16672);
xnor U23951 (N_23951,N_15014,N_15830);
or U23952 (N_23952,N_13796,N_13719);
nor U23953 (N_23953,N_18201,N_17856);
or U23954 (N_23954,N_18206,N_14757);
nand U23955 (N_23955,N_17775,N_16676);
nand U23956 (N_23956,N_13172,N_14333);
nor U23957 (N_23957,N_17455,N_15155);
nor U23958 (N_23958,N_17527,N_14380);
xnor U23959 (N_23959,N_13006,N_14277);
nand U23960 (N_23960,N_14229,N_13905);
xnor U23961 (N_23961,N_12660,N_15624);
and U23962 (N_23962,N_15806,N_14049);
xor U23963 (N_23963,N_17397,N_14090);
xnor U23964 (N_23964,N_18638,N_12926);
and U23965 (N_23965,N_15943,N_15383);
or U23966 (N_23966,N_14414,N_16078);
and U23967 (N_23967,N_13924,N_13683);
xor U23968 (N_23968,N_18451,N_16280);
nand U23969 (N_23969,N_18190,N_15018);
nor U23970 (N_23970,N_13236,N_18518);
and U23971 (N_23971,N_16768,N_15275);
xor U23972 (N_23972,N_15814,N_14602);
nor U23973 (N_23973,N_16430,N_13978);
nand U23974 (N_23974,N_16674,N_12892);
nor U23975 (N_23975,N_13680,N_14277);
xor U23976 (N_23976,N_16192,N_15689);
and U23977 (N_23977,N_12755,N_12728);
nand U23978 (N_23978,N_13292,N_15141);
or U23979 (N_23979,N_13725,N_13081);
or U23980 (N_23980,N_18591,N_17013);
or U23981 (N_23981,N_15312,N_12827);
and U23982 (N_23982,N_14254,N_14766);
xnor U23983 (N_23983,N_12511,N_14477);
and U23984 (N_23984,N_14058,N_14857);
nand U23985 (N_23985,N_15039,N_16588);
nor U23986 (N_23986,N_18506,N_16975);
or U23987 (N_23987,N_12671,N_13779);
or U23988 (N_23988,N_16352,N_13914);
xnor U23989 (N_23989,N_17852,N_15962);
nand U23990 (N_23990,N_17285,N_16265);
and U23991 (N_23991,N_17360,N_17773);
xor U23992 (N_23992,N_18214,N_16724);
nand U23993 (N_23993,N_14314,N_16265);
nand U23994 (N_23994,N_13640,N_14694);
nand U23995 (N_23995,N_16045,N_17554);
or U23996 (N_23996,N_18333,N_15627);
or U23997 (N_23997,N_15132,N_16808);
xor U23998 (N_23998,N_16696,N_15318);
and U23999 (N_23999,N_17365,N_15644);
and U24000 (N_24000,N_16352,N_14233);
nand U24001 (N_24001,N_18494,N_13670);
or U24002 (N_24002,N_16378,N_16335);
xnor U24003 (N_24003,N_15502,N_15411);
nor U24004 (N_24004,N_16495,N_15600);
or U24005 (N_24005,N_14577,N_16139);
xnor U24006 (N_24006,N_18262,N_17307);
or U24007 (N_24007,N_14388,N_17623);
and U24008 (N_24008,N_14994,N_12933);
nand U24009 (N_24009,N_17154,N_15709);
xnor U24010 (N_24010,N_15660,N_13624);
nor U24011 (N_24011,N_17174,N_14927);
and U24012 (N_24012,N_12950,N_16229);
xor U24013 (N_24013,N_14037,N_15535);
xnor U24014 (N_24014,N_14574,N_17773);
and U24015 (N_24015,N_15248,N_17325);
nor U24016 (N_24016,N_16931,N_16930);
xnor U24017 (N_24017,N_16291,N_15478);
and U24018 (N_24018,N_14747,N_13646);
and U24019 (N_24019,N_13611,N_12520);
nand U24020 (N_24020,N_17527,N_15699);
or U24021 (N_24021,N_17281,N_14950);
xnor U24022 (N_24022,N_15100,N_15722);
nand U24023 (N_24023,N_13192,N_17555);
and U24024 (N_24024,N_16318,N_14903);
nor U24025 (N_24025,N_13537,N_13121);
nor U24026 (N_24026,N_17272,N_15975);
xnor U24027 (N_24027,N_16612,N_13079);
nor U24028 (N_24028,N_12890,N_14741);
or U24029 (N_24029,N_18198,N_13916);
or U24030 (N_24030,N_15640,N_12797);
nor U24031 (N_24031,N_13304,N_15000);
and U24032 (N_24032,N_16963,N_13304);
or U24033 (N_24033,N_12991,N_17217);
nor U24034 (N_24034,N_15925,N_14177);
or U24035 (N_24035,N_18096,N_13482);
nor U24036 (N_24036,N_18002,N_15295);
nand U24037 (N_24037,N_17806,N_15685);
and U24038 (N_24038,N_13065,N_18186);
nor U24039 (N_24039,N_18163,N_12929);
xor U24040 (N_24040,N_15132,N_17988);
or U24041 (N_24041,N_17678,N_14557);
nor U24042 (N_24042,N_14214,N_13589);
nor U24043 (N_24043,N_18185,N_16553);
or U24044 (N_24044,N_13197,N_13880);
nor U24045 (N_24045,N_15649,N_17527);
and U24046 (N_24046,N_17925,N_15385);
xor U24047 (N_24047,N_17020,N_18315);
nor U24048 (N_24048,N_17140,N_13975);
or U24049 (N_24049,N_14617,N_16152);
or U24050 (N_24050,N_18523,N_13077);
or U24051 (N_24051,N_17327,N_16995);
or U24052 (N_24052,N_16943,N_13768);
or U24053 (N_24053,N_14465,N_14551);
xnor U24054 (N_24054,N_16080,N_15717);
xnor U24055 (N_24055,N_15612,N_17615);
and U24056 (N_24056,N_14452,N_18734);
xnor U24057 (N_24057,N_15822,N_15610);
and U24058 (N_24058,N_15231,N_15115);
and U24059 (N_24059,N_15868,N_15167);
nor U24060 (N_24060,N_18107,N_17443);
nor U24061 (N_24061,N_16315,N_14235);
nor U24062 (N_24062,N_18166,N_12975);
nand U24063 (N_24063,N_13128,N_18080);
xor U24064 (N_24064,N_16122,N_17636);
xnor U24065 (N_24065,N_13008,N_17938);
nor U24066 (N_24066,N_16899,N_16921);
nand U24067 (N_24067,N_17856,N_14037);
xor U24068 (N_24068,N_17980,N_16176);
or U24069 (N_24069,N_16569,N_15184);
xnor U24070 (N_24070,N_17278,N_16029);
nand U24071 (N_24071,N_17494,N_16004);
or U24072 (N_24072,N_16724,N_14059);
nor U24073 (N_24073,N_16578,N_16568);
and U24074 (N_24074,N_16755,N_13399);
and U24075 (N_24075,N_18633,N_17928);
or U24076 (N_24076,N_14600,N_13653);
and U24077 (N_24077,N_12572,N_16554);
and U24078 (N_24078,N_15500,N_16902);
nor U24079 (N_24079,N_15675,N_17908);
or U24080 (N_24080,N_15312,N_15573);
and U24081 (N_24081,N_13151,N_13947);
xnor U24082 (N_24082,N_15048,N_14525);
nor U24083 (N_24083,N_16901,N_12677);
nor U24084 (N_24084,N_17233,N_17219);
nor U24085 (N_24085,N_14462,N_16656);
nand U24086 (N_24086,N_13112,N_17272);
xor U24087 (N_24087,N_17964,N_12768);
nor U24088 (N_24088,N_18396,N_18484);
and U24089 (N_24089,N_16242,N_14186);
xnor U24090 (N_24090,N_12924,N_18465);
and U24091 (N_24091,N_17473,N_12589);
nand U24092 (N_24092,N_14904,N_17008);
nand U24093 (N_24093,N_16090,N_13498);
nor U24094 (N_24094,N_15647,N_14086);
nand U24095 (N_24095,N_14901,N_15628);
nand U24096 (N_24096,N_16853,N_13318);
or U24097 (N_24097,N_15637,N_13020);
nor U24098 (N_24098,N_17492,N_12789);
xor U24099 (N_24099,N_16606,N_17647);
nand U24100 (N_24100,N_15193,N_17949);
nor U24101 (N_24101,N_14428,N_13484);
nor U24102 (N_24102,N_13198,N_14178);
nor U24103 (N_24103,N_15321,N_15560);
nand U24104 (N_24104,N_18725,N_13149);
or U24105 (N_24105,N_18608,N_14285);
xnor U24106 (N_24106,N_13257,N_13317);
nand U24107 (N_24107,N_15156,N_18475);
or U24108 (N_24108,N_15741,N_17870);
or U24109 (N_24109,N_12544,N_15522);
or U24110 (N_24110,N_15301,N_12747);
or U24111 (N_24111,N_12911,N_16970);
or U24112 (N_24112,N_16849,N_14567);
and U24113 (N_24113,N_16130,N_13633);
and U24114 (N_24114,N_16342,N_18524);
xor U24115 (N_24115,N_17949,N_15084);
and U24116 (N_24116,N_18314,N_15029);
xnor U24117 (N_24117,N_17206,N_18221);
nand U24118 (N_24118,N_13208,N_12812);
xnor U24119 (N_24119,N_16930,N_15997);
and U24120 (N_24120,N_13819,N_14815);
and U24121 (N_24121,N_13419,N_13772);
nor U24122 (N_24122,N_14128,N_17822);
and U24123 (N_24123,N_14427,N_16974);
and U24124 (N_24124,N_15534,N_15954);
nor U24125 (N_24125,N_14566,N_15548);
nor U24126 (N_24126,N_13048,N_17265);
or U24127 (N_24127,N_13803,N_14017);
nand U24128 (N_24128,N_16825,N_15004);
and U24129 (N_24129,N_13336,N_16330);
xnor U24130 (N_24130,N_16571,N_14603);
nand U24131 (N_24131,N_13436,N_16797);
and U24132 (N_24132,N_17976,N_14659);
nand U24133 (N_24133,N_16820,N_15748);
nand U24134 (N_24134,N_16665,N_18631);
nand U24135 (N_24135,N_17033,N_12866);
nor U24136 (N_24136,N_18027,N_17260);
nor U24137 (N_24137,N_13668,N_14964);
nor U24138 (N_24138,N_14582,N_16360);
and U24139 (N_24139,N_16095,N_15279);
or U24140 (N_24140,N_17598,N_18540);
or U24141 (N_24141,N_12573,N_16250);
nand U24142 (N_24142,N_16119,N_16003);
xnor U24143 (N_24143,N_15395,N_16306);
and U24144 (N_24144,N_16205,N_16658);
nand U24145 (N_24145,N_14022,N_14311);
or U24146 (N_24146,N_16073,N_14150);
or U24147 (N_24147,N_18096,N_18015);
nand U24148 (N_24148,N_14749,N_12521);
xnor U24149 (N_24149,N_15280,N_17896);
xnor U24150 (N_24150,N_18512,N_14236);
nand U24151 (N_24151,N_13153,N_12966);
xor U24152 (N_24152,N_18079,N_16845);
nand U24153 (N_24153,N_15073,N_18724);
and U24154 (N_24154,N_15036,N_13369);
nor U24155 (N_24155,N_15430,N_17316);
and U24156 (N_24156,N_17171,N_14590);
xor U24157 (N_24157,N_16470,N_14100);
nand U24158 (N_24158,N_14121,N_13358);
nor U24159 (N_24159,N_18091,N_14838);
nand U24160 (N_24160,N_18723,N_16334);
or U24161 (N_24161,N_14862,N_14590);
nand U24162 (N_24162,N_15234,N_18480);
nand U24163 (N_24163,N_16439,N_16900);
nand U24164 (N_24164,N_15964,N_15097);
nor U24165 (N_24165,N_16130,N_12975);
nand U24166 (N_24166,N_18720,N_14606);
and U24167 (N_24167,N_16943,N_13087);
and U24168 (N_24168,N_14876,N_16207);
and U24169 (N_24169,N_17824,N_12680);
xnor U24170 (N_24170,N_18416,N_14616);
or U24171 (N_24171,N_15083,N_13942);
nor U24172 (N_24172,N_13987,N_17478);
or U24173 (N_24173,N_14891,N_15604);
or U24174 (N_24174,N_15400,N_13757);
xnor U24175 (N_24175,N_18381,N_13214);
nor U24176 (N_24176,N_13673,N_17092);
nor U24177 (N_24177,N_15146,N_14916);
and U24178 (N_24178,N_17977,N_14150);
or U24179 (N_24179,N_15347,N_17828);
and U24180 (N_24180,N_18570,N_16781);
and U24181 (N_24181,N_18523,N_15413);
nor U24182 (N_24182,N_14237,N_14568);
and U24183 (N_24183,N_17406,N_16907);
xor U24184 (N_24184,N_14063,N_17439);
and U24185 (N_24185,N_14436,N_16082);
or U24186 (N_24186,N_12558,N_15339);
xnor U24187 (N_24187,N_17270,N_18740);
or U24188 (N_24188,N_15275,N_12994);
nand U24189 (N_24189,N_18676,N_16482);
xor U24190 (N_24190,N_15203,N_15770);
nor U24191 (N_24191,N_17130,N_16135);
nor U24192 (N_24192,N_16382,N_16401);
nor U24193 (N_24193,N_16223,N_16220);
nor U24194 (N_24194,N_17929,N_16100);
xor U24195 (N_24195,N_13404,N_13081);
xor U24196 (N_24196,N_18111,N_14879);
xnor U24197 (N_24197,N_13034,N_16666);
nand U24198 (N_24198,N_13786,N_15140);
nor U24199 (N_24199,N_17917,N_18654);
nor U24200 (N_24200,N_14164,N_13224);
and U24201 (N_24201,N_18320,N_17603);
nand U24202 (N_24202,N_12770,N_14577);
or U24203 (N_24203,N_18660,N_16648);
or U24204 (N_24204,N_14603,N_14625);
nand U24205 (N_24205,N_13674,N_13147);
nand U24206 (N_24206,N_12587,N_12867);
nand U24207 (N_24207,N_15770,N_17769);
xor U24208 (N_24208,N_15807,N_17773);
xnor U24209 (N_24209,N_13809,N_16900);
nor U24210 (N_24210,N_14153,N_16522);
nand U24211 (N_24211,N_15846,N_13161);
xor U24212 (N_24212,N_17270,N_18001);
nand U24213 (N_24213,N_16604,N_16214);
and U24214 (N_24214,N_16349,N_18624);
xnor U24215 (N_24215,N_14690,N_14647);
and U24216 (N_24216,N_18714,N_16484);
nor U24217 (N_24217,N_14547,N_15502);
xor U24218 (N_24218,N_14337,N_14702);
nand U24219 (N_24219,N_13297,N_17585);
xnor U24220 (N_24220,N_14596,N_17632);
nand U24221 (N_24221,N_15800,N_14425);
nor U24222 (N_24222,N_17007,N_12588);
nand U24223 (N_24223,N_17286,N_13343);
and U24224 (N_24224,N_15630,N_17479);
xor U24225 (N_24225,N_17352,N_13198);
nor U24226 (N_24226,N_17375,N_17568);
nor U24227 (N_24227,N_15499,N_14712);
nand U24228 (N_24228,N_16745,N_14967);
nand U24229 (N_24229,N_15614,N_17037);
or U24230 (N_24230,N_14836,N_12772);
xor U24231 (N_24231,N_15824,N_17334);
nand U24232 (N_24232,N_16888,N_13269);
nor U24233 (N_24233,N_13515,N_14206);
or U24234 (N_24234,N_17918,N_18398);
nand U24235 (N_24235,N_14931,N_16294);
nor U24236 (N_24236,N_18138,N_14082);
and U24237 (N_24237,N_13727,N_14625);
and U24238 (N_24238,N_15952,N_17364);
or U24239 (N_24239,N_14515,N_15048);
or U24240 (N_24240,N_18046,N_15885);
or U24241 (N_24241,N_16610,N_15554);
nand U24242 (N_24242,N_17694,N_18582);
or U24243 (N_24243,N_15255,N_18534);
nor U24244 (N_24244,N_14577,N_16034);
nor U24245 (N_24245,N_12811,N_15688);
or U24246 (N_24246,N_12681,N_15223);
xor U24247 (N_24247,N_14236,N_15283);
nor U24248 (N_24248,N_15923,N_16782);
xor U24249 (N_24249,N_13750,N_14786);
nor U24250 (N_24250,N_13683,N_18421);
nand U24251 (N_24251,N_16977,N_16771);
or U24252 (N_24252,N_15860,N_16610);
nor U24253 (N_24253,N_15601,N_15396);
or U24254 (N_24254,N_13145,N_18289);
or U24255 (N_24255,N_15922,N_15018);
nor U24256 (N_24256,N_17982,N_17972);
and U24257 (N_24257,N_12654,N_12787);
or U24258 (N_24258,N_14099,N_17165);
xor U24259 (N_24259,N_18283,N_14377);
and U24260 (N_24260,N_13861,N_12879);
xnor U24261 (N_24261,N_15533,N_18474);
or U24262 (N_24262,N_15310,N_16714);
or U24263 (N_24263,N_16703,N_16042);
nor U24264 (N_24264,N_18562,N_15928);
and U24265 (N_24265,N_15346,N_12991);
xor U24266 (N_24266,N_18364,N_15586);
nand U24267 (N_24267,N_12736,N_13428);
or U24268 (N_24268,N_18087,N_18219);
nor U24269 (N_24269,N_13150,N_12752);
or U24270 (N_24270,N_18588,N_12555);
nand U24271 (N_24271,N_15601,N_13933);
and U24272 (N_24272,N_16729,N_14342);
xnor U24273 (N_24273,N_18660,N_14026);
and U24274 (N_24274,N_15852,N_17781);
or U24275 (N_24275,N_12650,N_18213);
or U24276 (N_24276,N_18621,N_15945);
nor U24277 (N_24277,N_16637,N_14553);
or U24278 (N_24278,N_12739,N_14699);
nor U24279 (N_24279,N_17052,N_16607);
nand U24280 (N_24280,N_15425,N_18454);
or U24281 (N_24281,N_18129,N_16891);
xor U24282 (N_24282,N_12617,N_16718);
nor U24283 (N_24283,N_18059,N_15940);
or U24284 (N_24284,N_12829,N_18474);
or U24285 (N_24285,N_15595,N_17097);
nand U24286 (N_24286,N_13346,N_14173);
nand U24287 (N_24287,N_16027,N_15458);
and U24288 (N_24288,N_14990,N_17186);
nor U24289 (N_24289,N_15045,N_13893);
or U24290 (N_24290,N_16063,N_17903);
and U24291 (N_24291,N_13644,N_18352);
xor U24292 (N_24292,N_14619,N_18464);
and U24293 (N_24293,N_15124,N_14910);
and U24294 (N_24294,N_14700,N_13702);
or U24295 (N_24295,N_15595,N_17754);
and U24296 (N_24296,N_16095,N_14838);
or U24297 (N_24297,N_14466,N_16669);
nand U24298 (N_24298,N_16299,N_18102);
nor U24299 (N_24299,N_15850,N_17788);
or U24300 (N_24300,N_14879,N_15446);
xor U24301 (N_24301,N_13477,N_17749);
or U24302 (N_24302,N_13681,N_16258);
nor U24303 (N_24303,N_15562,N_14341);
xnor U24304 (N_24304,N_15818,N_13768);
nand U24305 (N_24305,N_17267,N_15412);
xnor U24306 (N_24306,N_18019,N_13452);
nand U24307 (N_24307,N_15007,N_14256);
and U24308 (N_24308,N_15940,N_17312);
and U24309 (N_24309,N_13264,N_18045);
nor U24310 (N_24310,N_16592,N_16701);
and U24311 (N_24311,N_18333,N_13576);
xnor U24312 (N_24312,N_17269,N_17770);
nor U24313 (N_24313,N_14095,N_16446);
nand U24314 (N_24314,N_12681,N_13374);
nand U24315 (N_24315,N_14262,N_14026);
nor U24316 (N_24316,N_13790,N_17313);
nor U24317 (N_24317,N_17659,N_16657);
nand U24318 (N_24318,N_15780,N_18515);
nand U24319 (N_24319,N_17289,N_17181);
and U24320 (N_24320,N_13457,N_16390);
and U24321 (N_24321,N_12983,N_14504);
nand U24322 (N_24322,N_13452,N_15155);
or U24323 (N_24323,N_18121,N_14537);
and U24324 (N_24324,N_17094,N_15816);
and U24325 (N_24325,N_16651,N_15450);
or U24326 (N_24326,N_18255,N_18614);
and U24327 (N_24327,N_18034,N_17846);
xnor U24328 (N_24328,N_14931,N_18153);
or U24329 (N_24329,N_18362,N_12597);
or U24330 (N_24330,N_17385,N_14253);
xor U24331 (N_24331,N_13821,N_17215);
and U24332 (N_24332,N_17568,N_17962);
or U24333 (N_24333,N_18004,N_12668);
nand U24334 (N_24334,N_18377,N_15042);
nor U24335 (N_24335,N_15387,N_12682);
or U24336 (N_24336,N_15034,N_16639);
xor U24337 (N_24337,N_18617,N_13854);
nand U24338 (N_24338,N_12919,N_17061);
nor U24339 (N_24339,N_14936,N_14914);
or U24340 (N_24340,N_13930,N_14646);
nor U24341 (N_24341,N_13069,N_17404);
xor U24342 (N_24342,N_17137,N_14506);
nor U24343 (N_24343,N_15258,N_17792);
or U24344 (N_24344,N_15963,N_17690);
nand U24345 (N_24345,N_17195,N_15945);
nor U24346 (N_24346,N_17899,N_14697);
xnor U24347 (N_24347,N_16281,N_13611);
or U24348 (N_24348,N_17781,N_14759);
and U24349 (N_24349,N_15315,N_17149);
and U24350 (N_24350,N_12891,N_18524);
xnor U24351 (N_24351,N_14381,N_13712);
nor U24352 (N_24352,N_14855,N_17646);
or U24353 (N_24353,N_14047,N_14526);
nor U24354 (N_24354,N_13979,N_18445);
nor U24355 (N_24355,N_13574,N_18593);
xnor U24356 (N_24356,N_17415,N_14337);
nor U24357 (N_24357,N_13905,N_15279);
nand U24358 (N_24358,N_14955,N_15166);
and U24359 (N_24359,N_15775,N_17025);
and U24360 (N_24360,N_12768,N_18624);
nor U24361 (N_24361,N_16380,N_16041);
nor U24362 (N_24362,N_17436,N_15173);
xor U24363 (N_24363,N_18426,N_16630);
xnor U24364 (N_24364,N_14816,N_14360);
and U24365 (N_24365,N_15438,N_15833);
and U24366 (N_24366,N_12693,N_17276);
or U24367 (N_24367,N_13672,N_18234);
or U24368 (N_24368,N_17104,N_18442);
and U24369 (N_24369,N_13380,N_13279);
and U24370 (N_24370,N_14408,N_14429);
and U24371 (N_24371,N_16019,N_17009);
and U24372 (N_24372,N_14878,N_18017);
nor U24373 (N_24373,N_17751,N_16274);
nand U24374 (N_24374,N_17280,N_18198);
nor U24375 (N_24375,N_14517,N_14637);
xnor U24376 (N_24376,N_18490,N_18274);
xor U24377 (N_24377,N_12945,N_15706);
or U24378 (N_24378,N_13990,N_13747);
or U24379 (N_24379,N_15307,N_14739);
xnor U24380 (N_24380,N_17890,N_13447);
or U24381 (N_24381,N_15820,N_18333);
nand U24382 (N_24382,N_18589,N_16948);
xnor U24383 (N_24383,N_16461,N_18418);
nand U24384 (N_24384,N_15380,N_16787);
xor U24385 (N_24385,N_13525,N_14874);
nand U24386 (N_24386,N_18695,N_17090);
or U24387 (N_24387,N_13651,N_14372);
nor U24388 (N_24388,N_14195,N_17042);
nand U24389 (N_24389,N_14544,N_16837);
and U24390 (N_24390,N_16593,N_12816);
and U24391 (N_24391,N_17014,N_17617);
xor U24392 (N_24392,N_14367,N_13789);
xnor U24393 (N_24393,N_14648,N_17738);
nand U24394 (N_24394,N_15513,N_15221);
nand U24395 (N_24395,N_14540,N_17049);
xor U24396 (N_24396,N_17114,N_18471);
and U24397 (N_24397,N_16781,N_17137);
nand U24398 (N_24398,N_13707,N_14208);
nor U24399 (N_24399,N_17597,N_17043);
nand U24400 (N_24400,N_12830,N_16933);
nor U24401 (N_24401,N_17552,N_16947);
nand U24402 (N_24402,N_18514,N_17157);
xor U24403 (N_24403,N_13695,N_13026);
nor U24404 (N_24404,N_12855,N_13838);
xnor U24405 (N_24405,N_15161,N_17045);
xnor U24406 (N_24406,N_18622,N_17031);
nand U24407 (N_24407,N_18262,N_16220);
nor U24408 (N_24408,N_16804,N_15145);
nand U24409 (N_24409,N_14377,N_17925);
nand U24410 (N_24410,N_18001,N_16282);
nand U24411 (N_24411,N_13247,N_15090);
nand U24412 (N_24412,N_16140,N_16206);
nor U24413 (N_24413,N_16358,N_13473);
xnor U24414 (N_24414,N_17617,N_14512);
nor U24415 (N_24415,N_14820,N_17367);
or U24416 (N_24416,N_15553,N_15239);
xnor U24417 (N_24417,N_13709,N_13723);
or U24418 (N_24418,N_17925,N_16421);
xnor U24419 (N_24419,N_18141,N_16366);
nor U24420 (N_24420,N_13399,N_17575);
nor U24421 (N_24421,N_14428,N_18652);
and U24422 (N_24422,N_13203,N_12817);
or U24423 (N_24423,N_14110,N_12969);
nor U24424 (N_24424,N_13299,N_15385);
nor U24425 (N_24425,N_13035,N_16496);
or U24426 (N_24426,N_13871,N_17189);
and U24427 (N_24427,N_16045,N_17464);
and U24428 (N_24428,N_15507,N_14307);
xnor U24429 (N_24429,N_12868,N_13312);
or U24430 (N_24430,N_12706,N_18137);
and U24431 (N_24431,N_12818,N_15626);
nand U24432 (N_24432,N_18719,N_13797);
or U24433 (N_24433,N_15706,N_12600);
or U24434 (N_24434,N_16494,N_17674);
or U24435 (N_24435,N_13772,N_15894);
nand U24436 (N_24436,N_12986,N_13305);
nand U24437 (N_24437,N_17691,N_17225);
or U24438 (N_24438,N_14208,N_14123);
and U24439 (N_24439,N_12742,N_17849);
or U24440 (N_24440,N_13920,N_18365);
or U24441 (N_24441,N_16756,N_18215);
and U24442 (N_24442,N_15096,N_15446);
nor U24443 (N_24443,N_12528,N_15097);
or U24444 (N_24444,N_18335,N_13620);
and U24445 (N_24445,N_12991,N_13725);
xnor U24446 (N_24446,N_13701,N_17758);
nand U24447 (N_24447,N_13274,N_13064);
or U24448 (N_24448,N_16262,N_14264);
or U24449 (N_24449,N_17752,N_17262);
or U24450 (N_24450,N_13063,N_18476);
nand U24451 (N_24451,N_15237,N_16102);
or U24452 (N_24452,N_15548,N_15184);
or U24453 (N_24453,N_18562,N_18263);
nor U24454 (N_24454,N_17127,N_18128);
or U24455 (N_24455,N_15445,N_13667);
nand U24456 (N_24456,N_13222,N_14834);
and U24457 (N_24457,N_17936,N_15048);
xnor U24458 (N_24458,N_15832,N_16017);
nor U24459 (N_24459,N_16471,N_13187);
or U24460 (N_24460,N_17848,N_16292);
and U24461 (N_24461,N_18441,N_12917);
xor U24462 (N_24462,N_13412,N_13348);
xnor U24463 (N_24463,N_18112,N_15819);
or U24464 (N_24464,N_13822,N_14677);
xnor U24465 (N_24465,N_15095,N_16612);
or U24466 (N_24466,N_17463,N_16235);
and U24467 (N_24467,N_16934,N_18263);
or U24468 (N_24468,N_14321,N_14393);
and U24469 (N_24469,N_13413,N_14265);
or U24470 (N_24470,N_13990,N_17684);
and U24471 (N_24471,N_13027,N_13487);
nand U24472 (N_24472,N_16701,N_18523);
xnor U24473 (N_24473,N_16124,N_16282);
xnor U24474 (N_24474,N_14641,N_16185);
or U24475 (N_24475,N_15132,N_13408);
and U24476 (N_24476,N_13017,N_17155);
xor U24477 (N_24477,N_16437,N_12973);
nand U24478 (N_24478,N_13139,N_15854);
nor U24479 (N_24479,N_12605,N_18455);
nand U24480 (N_24480,N_13612,N_17143);
and U24481 (N_24481,N_16767,N_14071);
or U24482 (N_24482,N_13342,N_16908);
nor U24483 (N_24483,N_18208,N_12614);
and U24484 (N_24484,N_15830,N_15057);
or U24485 (N_24485,N_15827,N_13168);
and U24486 (N_24486,N_16105,N_18655);
xor U24487 (N_24487,N_18349,N_17767);
or U24488 (N_24488,N_16459,N_17047);
nand U24489 (N_24489,N_17677,N_18155);
nor U24490 (N_24490,N_14329,N_12564);
xor U24491 (N_24491,N_14983,N_12964);
or U24492 (N_24492,N_17897,N_16297);
or U24493 (N_24493,N_12629,N_13381);
xor U24494 (N_24494,N_15347,N_18677);
nor U24495 (N_24495,N_14155,N_13817);
nand U24496 (N_24496,N_12783,N_14471);
and U24497 (N_24497,N_15275,N_15881);
xnor U24498 (N_24498,N_14922,N_13701);
and U24499 (N_24499,N_12935,N_15157);
nor U24500 (N_24500,N_13269,N_15569);
nand U24501 (N_24501,N_14792,N_16858);
xnor U24502 (N_24502,N_17543,N_15312);
or U24503 (N_24503,N_16535,N_14378);
nand U24504 (N_24504,N_16637,N_14423);
nand U24505 (N_24505,N_14794,N_14223);
or U24506 (N_24506,N_18218,N_14615);
nand U24507 (N_24507,N_15546,N_16364);
and U24508 (N_24508,N_16926,N_15712);
xor U24509 (N_24509,N_17308,N_13815);
and U24510 (N_24510,N_15423,N_18061);
or U24511 (N_24511,N_12941,N_18098);
nand U24512 (N_24512,N_13847,N_14870);
nand U24513 (N_24513,N_16293,N_15297);
nor U24514 (N_24514,N_15315,N_13250);
xor U24515 (N_24515,N_16755,N_16115);
nand U24516 (N_24516,N_18570,N_13004);
and U24517 (N_24517,N_14148,N_14694);
xor U24518 (N_24518,N_16966,N_17502);
or U24519 (N_24519,N_17940,N_13229);
and U24520 (N_24520,N_15432,N_14591);
nor U24521 (N_24521,N_17546,N_13450);
and U24522 (N_24522,N_15732,N_14537);
nand U24523 (N_24523,N_12758,N_16060);
and U24524 (N_24524,N_16754,N_16111);
nand U24525 (N_24525,N_16390,N_16851);
or U24526 (N_24526,N_16591,N_15119);
nor U24527 (N_24527,N_15472,N_13084);
or U24528 (N_24528,N_17477,N_14743);
nand U24529 (N_24529,N_18153,N_17710);
or U24530 (N_24530,N_15478,N_18132);
and U24531 (N_24531,N_17125,N_17737);
or U24532 (N_24532,N_17557,N_16809);
and U24533 (N_24533,N_12932,N_14714);
nor U24534 (N_24534,N_13045,N_16266);
xor U24535 (N_24535,N_14420,N_16863);
nor U24536 (N_24536,N_13755,N_14689);
nand U24537 (N_24537,N_12541,N_14357);
nor U24538 (N_24538,N_14323,N_15458);
and U24539 (N_24539,N_14335,N_18513);
nor U24540 (N_24540,N_14908,N_15483);
and U24541 (N_24541,N_15537,N_16567);
xnor U24542 (N_24542,N_16969,N_17648);
and U24543 (N_24543,N_13546,N_12563);
or U24544 (N_24544,N_12567,N_15017);
and U24545 (N_24545,N_18683,N_15611);
or U24546 (N_24546,N_13015,N_13183);
nand U24547 (N_24547,N_17386,N_16340);
nand U24548 (N_24548,N_15573,N_14839);
and U24549 (N_24549,N_16842,N_14196);
nor U24550 (N_24550,N_14518,N_16395);
xor U24551 (N_24551,N_13835,N_13262);
nor U24552 (N_24552,N_15133,N_14191);
or U24553 (N_24553,N_14329,N_13438);
nor U24554 (N_24554,N_16282,N_16927);
xnor U24555 (N_24555,N_16832,N_18497);
nor U24556 (N_24556,N_14177,N_14173);
xnor U24557 (N_24557,N_15657,N_18019);
nand U24558 (N_24558,N_14684,N_18267);
and U24559 (N_24559,N_12989,N_17527);
or U24560 (N_24560,N_14101,N_13320);
and U24561 (N_24561,N_18033,N_17807);
and U24562 (N_24562,N_13308,N_15863);
or U24563 (N_24563,N_13210,N_16454);
nor U24564 (N_24564,N_14749,N_16143);
nor U24565 (N_24565,N_14071,N_16063);
nor U24566 (N_24566,N_15525,N_13843);
xnor U24567 (N_24567,N_16921,N_13624);
or U24568 (N_24568,N_17625,N_14759);
and U24569 (N_24569,N_13806,N_12840);
nor U24570 (N_24570,N_14973,N_18534);
xor U24571 (N_24571,N_15431,N_16749);
and U24572 (N_24572,N_17545,N_16554);
xor U24573 (N_24573,N_14526,N_17984);
xor U24574 (N_24574,N_16149,N_14757);
or U24575 (N_24575,N_15992,N_12918);
or U24576 (N_24576,N_13335,N_18013);
nor U24577 (N_24577,N_14486,N_13922);
nand U24578 (N_24578,N_15778,N_15425);
xor U24579 (N_24579,N_12763,N_18409);
nand U24580 (N_24580,N_16651,N_13371);
and U24581 (N_24581,N_13538,N_15198);
or U24582 (N_24582,N_17544,N_16918);
nand U24583 (N_24583,N_14219,N_16771);
nor U24584 (N_24584,N_18617,N_18522);
xnor U24585 (N_24585,N_16533,N_13894);
xor U24586 (N_24586,N_18684,N_15254);
or U24587 (N_24587,N_15941,N_16619);
or U24588 (N_24588,N_16665,N_18003);
or U24589 (N_24589,N_15428,N_14379);
xnor U24590 (N_24590,N_17067,N_14373);
or U24591 (N_24591,N_13864,N_13663);
xnor U24592 (N_24592,N_18655,N_18150);
xor U24593 (N_24593,N_13837,N_15330);
xnor U24594 (N_24594,N_16560,N_13819);
nor U24595 (N_24595,N_12726,N_14075);
xor U24596 (N_24596,N_13063,N_16478);
nor U24597 (N_24597,N_16546,N_15634);
and U24598 (N_24598,N_15052,N_12879);
nand U24599 (N_24599,N_16882,N_13048);
or U24600 (N_24600,N_18338,N_13448);
or U24601 (N_24601,N_14377,N_16520);
and U24602 (N_24602,N_17669,N_13359);
or U24603 (N_24603,N_13489,N_15739);
nor U24604 (N_24604,N_15864,N_15871);
or U24605 (N_24605,N_14113,N_16865);
and U24606 (N_24606,N_17625,N_14775);
xor U24607 (N_24607,N_13723,N_14203);
xnor U24608 (N_24608,N_17493,N_12764);
xnor U24609 (N_24609,N_14157,N_17523);
or U24610 (N_24610,N_13630,N_16349);
xnor U24611 (N_24611,N_13842,N_18177);
xnor U24612 (N_24612,N_13015,N_13068);
xnor U24613 (N_24613,N_17952,N_16147);
nor U24614 (N_24614,N_14254,N_13330);
and U24615 (N_24615,N_18230,N_18687);
xnor U24616 (N_24616,N_14515,N_16378);
nand U24617 (N_24617,N_13578,N_13624);
or U24618 (N_24618,N_15898,N_17953);
nand U24619 (N_24619,N_16912,N_15394);
xor U24620 (N_24620,N_18294,N_15119);
and U24621 (N_24621,N_14452,N_13600);
nand U24622 (N_24622,N_16249,N_13370);
nand U24623 (N_24623,N_18656,N_13064);
and U24624 (N_24624,N_15790,N_14673);
or U24625 (N_24625,N_13094,N_16733);
or U24626 (N_24626,N_14905,N_17446);
xor U24627 (N_24627,N_13459,N_17805);
or U24628 (N_24628,N_14915,N_14648);
and U24629 (N_24629,N_16950,N_17463);
nand U24630 (N_24630,N_13626,N_17083);
and U24631 (N_24631,N_17567,N_12936);
nand U24632 (N_24632,N_13572,N_16165);
xor U24633 (N_24633,N_15488,N_15258);
xor U24634 (N_24634,N_12566,N_13460);
nand U24635 (N_24635,N_13386,N_13793);
nor U24636 (N_24636,N_14782,N_15409);
or U24637 (N_24637,N_17049,N_16583);
xor U24638 (N_24638,N_14866,N_17239);
xor U24639 (N_24639,N_12553,N_16525);
nor U24640 (N_24640,N_17928,N_14779);
and U24641 (N_24641,N_15897,N_16589);
nor U24642 (N_24642,N_12608,N_14854);
xor U24643 (N_24643,N_17919,N_12926);
and U24644 (N_24644,N_15192,N_13055);
or U24645 (N_24645,N_16062,N_12749);
or U24646 (N_24646,N_13615,N_12512);
xnor U24647 (N_24647,N_15499,N_14539);
or U24648 (N_24648,N_17186,N_16489);
nand U24649 (N_24649,N_15625,N_16466);
or U24650 (N_24650,N_14333,N_18202);
nor U24651 (N_24651,N_12669,N_15741);
nand U24652 (N_24652,N_17608,N_17233);
or U24653 (N_24653,N_18697,N_14928);
nor U24654 (N_24654,N_12510,N_16628);
and U24655 (N_24655,N_12511,N_14106);
nor U24656 (N_24656,N_14738,N_17867);
nand U24657 (N_24657,N_13766,N_16083);
and U24658 (N_24658,N_13225,N_18302);
nand U24659 (N_24659,N_13592,N_14021);
nor U24660 (N_24660,N_14939,N_17697);
nor U24661 (N_24661,N_17540,N_13674);
xor U24662 (N_24662,N_16493,N_15079);
xnor U24663 (N_24663,N_17716,N_14347);
or U24664 (N_24664,N_15941,N_16301);
nor U24665 (N_24665,N_13062,N_16936);
xor U24666 (N_24666,N_15246,N_16244);
and U24667 (N_24667,N_18740,N_18377);
or U24668 (N_24668,N_13528,N_17340);
and U24669 (N_24669,N_15276,N_16053);
nor U24670 (N_24670,N_15940,N_14349);
and U24671 (N_24671,N_14434,N_12716);
nand U24672 (N_24672,N_12860,N_18560);
nor U24673 (N_24673,N_13999,N_13108);
or U24674 (N_24674,N_13206,N_17087);
nor U24675 (N_24675,N_15330,N_17606);
or U24676 (N_24676,N_17493,N_13429);
or U24677 (N_24677,N_15136,N_14722);
nand U24678 (N_24678,N_16421,N_14306);
nor U24679 (N_24679,N_15293,N_16369);
and U24680 (N_24680,N_16085,N_13712);
and U24681 (N_24681,N_15238,N_18050);
nor U24682 (N_24682,N_15494,N_18399);
and U24683 (N_24683,N_13408,N_14730);
nand U24684 (N_24684,N_17844,N_12715);
nand U24685 (N_24685,N_16777,N_12698);
xor U24686 (N_24686,N_17555,N_17340);
and U24687 (N_24687,N_18566,N_14764);
or U24688 (N_24688,N_18095,N_15933);
xnor U24689 (N_24689,N_17243,N_13757);
or U24690 (N_24690,N_17521,N_15468);
nor U24691 (N_24691,N_18235,N_12887);
nor U24692 (N_24692,N_14453,N_13414);
nand U24693 (N_24693,N_14368,N_16702);
nand U24694 (N_24694,N_13841,N_13923);
or U24695 (N_24695,N_12844,N_16900);
nand U24696 (N_24696,N_17937,N_17679);
nor U24697 (N_24697,N_18029,N_12952);
and U24698 (N_24698,N_17431,N_16913);
xnor U24699 (N_24699,N_14275,N_17300);
xnor U24700 (N_24700,N_13754,N_13287);
and U24701 (N_24701,N_13680,N_15532);
xnor U24702 (N_24702,N_14617,N_18568);
or U24703 (N_24703,N_14859,N_18322);
or U24704 (N_24704,N_15793,N_14571);
nor U24705 (N_24705,N_18425,N_17399);
nand U24706 (N_24706,N_14229,N_12909);
and U24707 (N_24707,N_16103,N_15348);
xnor U24708 (N_24708,N_15143,N_13441);
and U24709 (N_24709,N_16160,N_16595);
xnor U24710 (N_24710,N_13821,N_13677);
or U24711 (N_24711,N_13224,N_17435);
nor U24712 (N_24712,N_14787,N_16142);
and U24713 (N_24713,N_16752,N_17787);
or U24714 (N_24714,N_18315,N_12595);
and U24715 (N_24715,N_13481,N_15823);
or U24716 (N_24716,N_15680,N_16262);
or U24717 (N_24717,N_15009,N_15344);
nand U24718 (N_24718,N_18522,N_17101);
nand U24719 (N_24719,N_13333,N_14623);
nor U24720 (N_24720,N_15339,N_13648);
xnor U24721 (N_24721,N_16032,N_17209);
or U24722 (N_24722,N_13473,N_14247);
and U24723 (N_24723,N_16416,N_12754);
and U24724 (N_24724,N_18682,N_17518);
and U24725 (N_24725,N_15770,N_13595);
and U24726 (N_24726,N_14385,N_12666);
nor U24727 (N_24727,N_15369,N_16024);
nand U24728 (N_24728,N_16542,N_12630);
xor U24729 (N_24729,N_17398,N_15311);
nor U24730 (N_24730,N_13392,N_17240);
xor U24731 (N_24731,N_18720,N_15236);
and U24732 (N_24732,N_16096,N_14962);
nor U24733 (N_24733,N_14838,N_13496);
xor U24734 (N_24734,N_13254,N_17958);
xnor U24735 (N_24735,N_14881,N_16702);
nor U24736 (N_24736,N_18154,N_15706);
nand U24737 (N_24737,N_15110,N_14095);
nand U24738 (N_24738,N_17423,N_16310);
or U24739 (N_24739,N_16448,N_17211);
xor U24740 (N_24740,N_14612,N_18687);
or U24741 (N_24741,N_13189,N_17962);
and U24742 (N_24742,N_16603,N_17530);
and U24743 (N_24743,N_15710,N_17882);
or U24744 (N_24744,N_13653,N_16244);
and U24745 (N_24745,N_14181,N_17489);
nand U24746 (N_24746,N_13025,N_13571);
or U24747 (N_24747,N_15699,N_16020);
or U24748 (N_24748,N_14160,N_16777);
nor U24749 (N_24749,N_15213,N_15142);
or U24750 (N_24750,N_17375,N_15981);
xor U24751 (N_24751,N_16320,N_18030);
nand U24752 (N_24752,N_18618,N_14618);
xnor U24753 (N_24753,N_15669,N_16404);
or U24754 (N_24754,N_14567,N_13926);
xor U24755 (N_24755,N_18421,N_13988);
xnor U24756 (N_24756,N_14227,N_17243);
and U24757 (N_24757,N_18297,N_12922);
nor U24758 (N_24758,N_18280,N_16628);
nand U24759 (N_24759,N_13367,N_17421);
and U24760 (N_24760,N_15665,N_13619);
nor U24761 (N_24761,N_17811,N_13518);
nand U24762 (N_24762,N_16986,N_12698);
xnor U24763 (N_24763,N_18302,N_18207);
xor U24764 (N_24764,N_12701,N_15009);
xor U24765 (N_24765,N_15118,N_16743);
and U24766 (N_24766,N_16616,N_14497);
nor U24767 (N_24767,N_18000,N_14394);
or U24768 (N_24768,N_18670,N_13427);
or U24769 (N_24769,N_15499,N_13471);
and U24770 (N_24770,N_13303,N_18011);
or U24771 (N_24771,N_13494,N_14856);
nand U24772 (N_24772,N_17604,N_18006);
nand U24773 (N_24773,N_17166,N_13934);
and U24774 (N_24774,N_15779,N_13463);
nor U24775 (N_24775,N_16548,N_17481);
nor U24776 (N_24776,N_15225,N_16312);
and U24777 (N_24777,N_16852,N_17454);
and U24778 (N_24778,N_16019,N_16048);
and U24779 (N_24779,N_16994,N_16170);
nor U24780 (N_24780,N_12579,N_15694);
xnor U24781 (N_24781,N_14531,N_13573);
or U24782 (N_24782,N_18496,N_15682);
nor U24783 (N_24783,N_13673,N_14494);
or U24784 (N_24784,N_16366,N_15608);
nand U24785 (N_24785,N_15904,N_15719);
nor U24786 (N_24786,N_16586,N_18140);
nand U24787 (N_24787,N_16793,N_12715);
and U24788 (N_24788,N_18106,N_18440);
and U24789 (N_24789,N_18411,N_18144);
nor U24790 (N_24790,N_18347,N_18558);
xor U24791 (N_24791,N_16949,N_13280);
nand U24792 (N_24792,N_14404,N_17813);
or U24793 (N_24793,N_16834,N_16034);
or U24794 (N_24794,N_16302,N_15134);
xnor U24795 (N_24795,N_13813,N_17862);
and U24796 (N_24796,N_13685,N_15285);
nor U24797 (N_24797,N_17631,N_17638);
nand U24798 (N_24798,N_18126,N_17909);
xnor U24799 (N_24799,N_17953,N_17326);
nor U24800 (N_24800,N_14350,N_16786);
nor U24801 (N_24801,N_17408,N_17592);
xor U24802 (N_24802,N_17201,N_16469);
or U24803 (N_24803,N_15931,N_14742);
nor U24804 (N_24804,N_17102,N_18449);
xnor U24805 (N_24805,N_17481,N_15964);
or U24806 (N_24806,N_13564,N_13469);
nand U24807 (N_24807,N_15771,N_16009);
nand U24808 (N_24808,N_16347,N_13082);
nor U24809 (N_24809,N_15742,N_18098);
or U24810 (N_24810,N_14537,N_15906);
nor U24811 (N_24811,N_15301,N_17300);
xor U24812 (N_24812,N_15940,N_17833);
nand U24813 (N_24813,N_16716,N_14433);
or U24814 (N_24814,N_15583,N_13418);
nor U24815 (N_24815,N_15447,N_18602);
or U24816 (N_24816,N_14240,N_13487);
and U24817 (N_24817,N_15886,N_12772);
nor U24818 (N_24818,N_12701,N_17064);
or U24819 (N_24819,N_13114,N_14256);
nand U24820 (N_24820,N_14227,N_14988);
nand U24821 (N_24821,N_17672,N_16055);
and U24822 (N_24822,N_13123,N_17505);
nand U24823 (N_24823,N_16648,N_14351);
xnor U24824 (N_24824,N_18081,N_18066);
xnor U24825 (N_24825,N_14052,N_14841);
or U24826 (N_24826,N_14865,N_13857);
nand U24827 (N_24827,N_13662,N_13980);
nand U24828 (N_24828,N_16372,N_17416);
nand U24829 (N_24829,N_14673,N_16385);
xnor U24830 (N_24830,N_14610,N_12576);
or U24831 (N_24831,N_18499,N_15396);
nor U24832 (N_24832,N_14412,N_16232);
or U24833 (N_24833,N_12874,N_18483);
nor U24834 (N_24834,N_14934,N_15332);
or U24835 (N_24835,N_15938,N_12784);
nand U24836 (N_24836,N_15335,N_18190);
nor U24837 (N_24837,N_18015,N_13171);
xor U24838 (N_24838,N_15099,N_14665);
nor U24839 (N_24839,N_14747,N_16095);
xor U24840 (N_24840,N_16519,N_18489);
and U24841 (N_24841,N_17172,N_13908);
and U24842 (N_24842,N_15226,N_17622);
nor U24843 (N_24843,N_15714,N_16394);
nor U24844 (N_24844,N_16058,N_15008);
xor U24845 (N_24845,N_17889,N_15183);
or U24846 (N_24846,N_15561,N_16712);
and U24847 (N_24847,N_18511,N_16914);
or U24848 (N_24848,N_13558,N_16462);
or U24849 (N_24849,N_14571,N_14543);
or U24850 (N_24850,N_15904,N_17154);
and U24851 (N_24851,N_18199,N_18399);
nor U24852 (N_24852,N_16845,N_14446);
xnor U24853 (N_24853,N_15272,N_15531);
and U24854 (N_24854,N_13697,N_14981);
xnor U24855 (N_24855,N_16682,N_15930);
nand U24856 (N_24856,N_15890,N_15560);
or U24857 (N_24857,N_15439,N_12817);
xnor U24858 (N_24858,N_13849,N_16132);
or U24859 (N_24859,N_14875,N_13583);
xnor U24860 (N_24860,N_14022,N_14222);
nand U24861 (N_24861,N_16200,N_16768);
xor U24862 (N_24862,N_16578,N_15256);
xnor U24863 (N_24863,N_15170,N_15332);
nor U24864 (N_24864,N_17104,N_17285);
nor U24865 (N_24865,N_16908,N_15009);
nor U24866 (N_24866,N_16760,N_13986);
and U24867 (N_24867,N_14684,N_15013);
xnor U24868 (N_24868,N_15008,N_12971);
nor U24869 (N_24869,N_16746,N_14747);
nor U24870 (N_24870,N_13473,N_15326);
nor U24871 (N_24871,N_13945,N_14883);
xor U24872 (N_24872,N_16444,N_18180);
nand U24873 (N_24873,N_13118,N_18280);
nor U24874 (N_24874,N_12886,N_14151);
or U24875 (N_24875,N_16244,N_15410);
nor U24876 (N_24876,N_17386,N_14162);
or U24877 (N_24877,N_14131,N_13515);
or U24878 (N_24878,N_15561,N_17274);
xor U24879 (N_24879,N_18360,N_13250);
xor U24880 (N_24880,N_17309,N_13305);
or U24881 (N_24881,N_17159,N_16973);
or U24882 (N_24882,N_14745,N_18123);
and U24883 (N_24883,N_16191,N_13443);
nor U24884 (N_24884,N_14239,N_12973);
nor U24885 (N_24885,N_18173,N_17151);
and U24886 (N_24886,N_16956,N_18443);
or U24887 (N_24887,N_17665,N_12591);
nand U24888 (N_24888,N_15626,N_18214);
and U24889 (N_24889,N_18679,N_12606);
and U24890 (N_24890,N_12644,N_17588);
or U24891 (N_24891,N_18324,N_18150);
nand U24892 (N_24892,N_15756,N_12581);
xor U24893 (N_24893,N_12771,N_17574);
nor U24894 (N_24894,N_16865,N_13793);
and U24895 (N_24895,N_14506,N_15639);
nor U24896 (N_24896,N_14263,N_16219);
and U24897 (N_24897,N_17599,N_17850);
nor U24898 (N_24898,N_15232,N_13740);
or U24899 (N_24899,N_17131,N_18689);
or U24900 (N_24900,N_14304,N_16687);
and U24901 (N_24901,N_13881,N_17753);
xnor U24902 (N_24902,N_14613,N_14444);
nand U24903 (N_24903,N_13506,N_17280);
or U24904 (N_24904,N_13703,N_18606);
or U24905 (N_24905,N_18708,N_17265);
and U24906 (N_24906,N_16504,N_13670);
xor U24907 (N_24907,N_13555,N_16482);
xor U24908 (N_24908,N_13927,N_13797);
xnor U24909 (N_24909,N_14620,N_15053);
nand U24910 (N_24910,N_14117,N_13720);
nor U24911 (N_24911,N_15549,N_13250);
xor U24912 (N_24912,N_16076,N_15380);
nor U24913 (N_24913,N_15390,N_13489);
or U24914 (N_24914,N_12796,N_14063);
nand U24915 (N_24915,N_18320,N_17453);
and U24916 (N_24916,N_18080,N_15123);
xnor U24917 (N_24917,N_16987,N_16590);
nand U24918 (N_24918,N_18268,N_16202);
nand U24919 (N_24919,N_17376,N_15907);
nand U24920 (N_24920,N_18463,N_14557);
and U24921 (N_24921,N_16132,N_13192);
and U24922 (N_24922,N_17785,N_13731);
and U24923 (N_24923,N_16816,N_15118);
nand U24924 (N_24924,N_16542,N_16830);
and U24925 (N_24925,N_13987,N_15549);
xnor U24926 (N_24926,N_14270,N_18271);
xnor U24927 (N_24927,N_14286,N_17245);
nand U24928 (N_24928,N_13305,N_16064);
nor U24929 (N_24929,N_14616,N_13200);
xnor U24930 (N_24930,N_16283,N_13287);
nor U24931 (N_24931,N_13121,N_16437);
and U24932 (N_24932,N_15007,N_17493);
and U24933 (N_24933,N_14816,N_18079);
nand U24934 (N_24934,N_18586,N_16622);
or U24935 (N_24935,N_17933,N_15903);
xnor U24936 (N_24936,N_14841,N_13529);
nand U24937 (N_24937,N_18567,N_17271);
or U24938 (N_24938,N_15918,N_17078);
nand U24939 (N_24939,N_17760,N_16445);
xnor U24940 (N_24940,N_15869,N_17520);
nand U24941 (N_24941,N_12772,N_13958);
nor U24942 (N_24942,N_18407,N_14922);
nor U24943 (N_24943,N_12539,N_13005);
xnor U24944 (N_24944,N_13219,N_17382);
or U24945 (N_24945,N_17628,N_17587);
nor U24946 (N_24946,N_15339,N_13163);
nor U24947 (N_24947,N_13709,N_18121);
and U24948 (N_24948,N_13450,N_14925);
nor U24949 (N_24949,N_18565,N_15792);
xor U24950 (N_24950,N_13360,N_14741);
xnor U24951 (N_24951,N_14281,N_15853);
xnor U24952 (N_24952,N_18679,N_15417);
xnor U24953 (N_24953,N_14340,N_17558);
nand U24954 (N_24954,N_13346,N_17583);
and U24955 (N_24955,N_18252,N_15512);
nand U24956 (N_24956,N_12974,N_14643);
or U24957 (N_24957,N_14064,N_12613);
or U24958 (N_24958,N_14083,N_13828);
xnor U24959 (N_24959,N_12691,N_15133);
nor U24960 (N_24960,N_13609,N_13532);
nor U24961 (N_24961,N_18446,N_15447);
xnor U24962 (N_24962,N_17622,N_15057);
nand U24963 (N_24963,N_15734,N_12734);
and U24964 (N_24964,N_18133,N_13857);
nor U24965 (N_24965,N_14027,N_17840);
and U24966 (N_24966,N_17690,N_16222);
or U24967 (N_24967,N_13055,N_18660);
and U24968 (N_24968,N_13339,N_16614);
or U24969 (N_24969,N_18455,N_15645);
or U24970 (N_24970,N_12567,N_13383);
and U24971 (N_24971,N_14251,N_14343);
xnor U24972 (N_24972,N_14748,N_18118);
xor U24973 (N_24973,N_14581,N_15513);
xnor U24974 (N_24974,N_14886,N_17684);
and U24975 (N_24975,N_16395,N_18512);
xor U24976 (N_24976,N_16205,N_14777);
or U24977 (N_24977,N_13501,N_14153);
and U24978 (N_24978,N_13585,N_12989);
nand U24979 (N_24979,N_15022,N_16544);
nand U24980 (N_24980,N_17752,N_14023);
nor U24981 (N_24981,N_15040,N_16382);
and U24982 (N_24982,N_17879,N_14712);
xnor U24983 (N_24983,N_12866,N_13415);
nor U24984 (N_24984,N_18398,N_13531);
nor U24985 (N_24985,N_15278,N_16287);
xor U24986 (N_24986,N_15376,N_17432);
xnor U24987 (N_24987,N_14567,N_17234);
and U24988 (N_24988,N_16829,N_16116);
or U24989 (N_24989,N_12947,N_17943);
xnor U24990 (N_24990,N_13307,N_15802);
nor U24991 (N_24991,N_17916,N_13596);
nand U24992 (N_24992,N_15046,N_17401);
nor U24993 (N_24993,N_16142,N_17937);
or U24994 (N_24994,N_18149,N_18292);
xnor U24995 (N_24995,N_14103,N_15420);
nor U24996 (N_24996,N_17329,N_12646);
nor U24997 (N_24997,N_14061,N_14068);
or U24998 (N_24998,N_18709,N_17207);
and U24999 (N_24999,N_16263,N_14277);
nand UO_0 (O_0,N_22925,N_21369);
xor UO_1 (O_1,N_20701,N_24384);
nor UO_2 (O_2,N_24664,N_22521);
xnor UO_3 (O_3,N_19215,N_19408);
nand UO_4 (O_4,N_19418,N_19632);
nand UO_5 (O_5,N_21333,N_21043);
and UO_6 (O_6,N_18876,N_19011);
and UO_7 (O_7,N_20006,N_21719);
and UO_8 (O_8,N_21404,N_21950);
xor UO_9 (O_9,N_18998,N_19535);
and UO_10 (O_10,N_20676,N_22571);
xnor UO_11 (O_11,N_23289,N_24980);
nand UO_12 (O_12,N_21812,N_20881);
or UO_13 (O_13,N_22203,N_21936);
xnor UO_14 (O_14,N_20506,N_21656);
xnor UO_15 (O_15,N_19096,N_24360);
or UO_16 (O_16,N_22313,N_19920);
nor UO_17 (O_17,N_24894,N_23616);
nand UO_18 (O_18,N_24608,N_22901);
or UO_19 (O_19,N_22886,N_23480);
nor UO_20 (O_20,N_22380,N_22813);
and UO_21 (O_21,N_22047,N_18960);
nand UO_22 (O_22,N_18976,N_20234);
or UO_23 (O_23,N_19177,N_24299);
nand UO_24 (O_24,N_20409,N_20995);
nand UO_25 (O_25,N_19650,N_24146);
nand UO_26 (O_26,N_21984,N_21946);
or UO_27 (O_27,N_22093,N_23935);
or UO_28 (O_28,N_23320,N_22974);
and UO_29 (O_29,N_21356,N_21045);
nor UO_30 (O_30,N_20978,N_20094);
xor UO_31 (O_31,N_23813,N_20810);
xor UO_32 (O_32,N_24305,N_20025);
or UO_33 (O_33,N_21086,N_21491);
xnor UO_34 (O_34,N_24656,N_21835);
nor UO_35 (O_35,N_21989,N_19162);
xnor UO_36 (O_36,N_19298,N_23632);
nor UO_37 (O_37,N_20690,N_23629);
or UO_38 (O_38,N_19022,N_24239);
nor UO_39 (O_39,N_20937,N_21374);
or UO_40 (O_40,N_24307,N_20572);
xor UO_41 (O_41,N_23266,N_20704);
and UO_42 (O_42,N_24069,N_21585);
nor UO_43 (O_43,N_20003,N_23386);
nor UO_44 (O_44,N_22956,N_19017);
or UO_45 (O_45,N_20430,N_21629);
or UO_46 (O_46,N_22645,N_19361);
nor UO_47 (O_47,N_22557,N_21772);
or UO_48 (O_48,N_21108,N_21484);
and UO_49 (O_49,N_24851,N_21923);
and UO_50 (O_50,N_24815,N_19123);
and UO_51 (O_51,N_23137,N_23850);
or UO_52 (O_52,N_24210,N_20962);
nand UO_53 (O_53,N_22719,N_18944);
xor UO_54 (O_54,N_20418,N_22844);
nor UO_55 (O_55,N_19611,N_21994);
nor UO_56 (O_56,N_21534,N_22800);
nor UO_57 (O_57,N_19240,N_19502);
or UO_58 (O_58,N_18811,N_22845);
and UO_59 (O_59,N_21031,N_21283);
xor UO_60 (O_60,N_24694,N_22466);
or UO_61 (O_61,N_18886,N_19191);
or UO_62 (O_62,N_24992,N_20903);
or UO_63 (O_63,N_24927,N_21582);
xnor UO_64 (O_64,N_20406,N_23930);
or UO_65 (O_65,N_24734,N_24657);
xnor UO_66 (O_66,N_20100,N_21420);
and UO_67 (O_67,N_23640,N_20186);
nor UO_68 (O_68,N_20687,N_24497);
nand UO_69 (O_69,N_21345,N_24603);
nor UO_70 (O_70,N_24433,N_23102);
nand UO_71 (O_71,N_21864,N_23905);
nand UO_72 (O_72,N_22105,N_21865);
nand UO_73 (O_73,N_20432,N_23955);
nand UO_74 (O_74,N_23599,N_19027);
nand UO_75 (O_75,N_18987,N_21872);
nor UO_76 (O_76,N_23942,N_23365);
xor UO_77 (O_77,N_20885,N_21640);
xor UO_78 (O_78,N_24775,N_19972);
or UO_79 (O_79,N_22605,N_23756);
nor UO_80 (O_80,N_19385,N_24364);
and UO_81 (O_81,N_20139,N_19855);
and UO_82 (O_82,N_22708,N_20161);
nor UO_83 (O_83,N_24692,N_19796);
or UO_84 (O_84,N_19763,N_19308);
xor UO_85 (O_85,N_23626,N_22268);
nor UO_86 (O_86,N_24139,N_24501);
and UO_87 (O_87,N_24285,N_20815);
and UO_88 (O_88,N_23001,N_22164);
nand UO_89 (O_89,N_20012,N_23400);
or UO_90 (O_90,N_23807,N_20498);
and UO_91 (O_91,N_19599,N_24401);
xnor UO_92 (O_92,N_24665,N_20279);
and UO_93 (O_93,N_19380,N_20171);
xor UO_94 (O_94,N_22447,N_23095);
or UO_95 (O_95,N_22256,N_19866);
xor UO_96 (O_96,N_22285,N_24088);
and UO_97 (O_97,N_19830,N_19672);
nand UO_98 (O_98,N_24674,N_18908);
and UO_99 (O_99,N_23451,N_24796);
and UO_100 (O_100,N_21882,N_22084);
xnor UO_101 (O_101,N_20589,N_19346);
nand UO_102 (O_102,N_22910,N_22151);
and UO_103 (O_103,N_23624,N_19420);
xnor UO_104 (O_104,N_20327,N_20452);
nand UO_105 (O_105,N_24746,N_20342);
nand UO_106 (O_106,N_24250,N_22420);
or UO_107 (O_107,N_23529,N_24414);
nand UO_108 (O_108,N_22930,N_19433);
nor UO_109 (O_109,N_24207,N_21120);
or UO_110 (O_110,N_24846,N_22599);
or UO_111 (O_111,N_19384,N_22860);
or UO_112 (O_112,N_20276,N_21712);
nor UO_113 (O_113,N_21925,N_23628);
nor UO_114 (O_114,N_21189,N_18843);
or UO_115 (O_115,N_23117,N_24074);
or UO_116 (O_116,N_19442,N_20608);
and UO_117 (O_117,N_22622,N_24131);
and UO_118 (O_118,N_24975,N_23646);
nand UO_119 (O_119,N_22887,N_19147);
xnor UO_120 (O_120,N_23174,N_21439);
or UO_121 (O_121,N_24693,N_21735);
nor UO_122 (O_122,N_22903,N_24300);
or UO_123 (O_123,N_24647,N_19540);
xnor UO_124 (O_124,N_19768,N_19640);
nand UO_125 (O_125,N_19102,N_21178);
nand UO_126 (O_126,N_23555,N_24278);
and UO_127 (O_127,N_24281,N_23871);
nand UO_128 (O_128,N_21126,N_23333);
nand UO_129 (O_129,N_24643,N_22265);
xnor UO_130 (O_130,N_20669,N_22733);
xor UO_131 (O_131,N_19862,N_18757);
and UO_132 (O_132,N_24486,N_23424);
or UO_133 (O_133,N_24151,N_19293);
nor UO_134 (O_134,N_23188,N_21163);
nand UO_135 (O_135,N_18924,N_24130);
xnor UO_136 (O_136,N_23917,N_24725);
or UO_137 (O_137,N_22003,N_21753);
or UO_138 (O_138,N_19890,N_21760);
xor UO_139 (O_139,N_19974,N_23432);
nand UO_140 (O_140,N_22350,N_21742);
and UO_141 (O_141,N_20880,N_19549);
and UO_142 (O_142,N_19787,N_21687);
and UO_143 (O_143,N_21986,N_19133);
and UO_144 (O_144,N_23833,N_21727);
nand UO_145 (O_145,N_20359,N_19633);
or UO_146 (O_146,N_23715,N_23338);
and UO_147 (O_147,N_22361,N_23517);
nand UO_148 (O_148,N_19000,N_22549);
nand UO_149 (O_149,N_24524,N_19350);
and UO_150 (O_150,N_22102,N_22324);
nor UO_151 (O_151,N_21911,N_19739);
nand UO_152 (O_152,N_18991,N_20874);
and UO_153 (O_153,N_20629,N_20328);
xnor UO_154 (O_154,N_21442,N_20622);
nor UO_155 (O_155,N_18899,N_23429);
and UO_156 (O_156,N_21059,N_23893);
and UO_157 (O_157,N_21039,N_24472);
and UO_158 (O_158,N_21739,N_21583);
xor UO_159 (O_159,N_20079,N_23571);
or UO_160 (O_160,N_21533,N_20996);
or UO_161 (O_161,N_24425,N_24500);
nor UO_162 (O_162,N_22527,N_22160);
nor UO_163 (O_163,N_24771,N_22184);
and UO_164 (O_164,N_23892,N_19223);
or UO_165 (O_165,N_19994,N_21868);
nor UO_166 (O_166,N_23090,N_20239);
xor UO_167 (O_167,N_20592,N_20886);
nor UO_168 (O_168,N_21386,N_20770);
and UO_169 (O_169,N_23855,N_23869);
nor UO_170 (O_170,N_24566,N_18895);
and UO_171 (O_171,N_23899,N_21990);
and UO_172 (O_172,N_20068,N_21317);
nor UO_173 (O_173,N_19959,N_19853);
nand UO_174 (O_174,N_19288,N_23346);
and UO_175 (O_175,N_23963,N_20296);
or UO_176 (O_176,N_22700,N_22567);
nand UO_177 (O_177,N_22713,N_24764);
and UO_178 (O_178,N_24323,N_19557);
nor UO_179 (O_179,N_19092,N_22033);
xnor UO_180 (O_180,N_19124,N_20421);
or UO_181 (O_181,N_24957,N_20210);
nor UO_182 (O_182,N_21274,N_19815);
or UO_183 (O_183,N_21612,N_24451);
nor UO_184 (O_184,N_20797,N_22192);
nor UO_185 (O_185,N_21871,N_23933);
and UO_186 (O_186,N_19860,N_21110);
or UO_187 (O_187,N_20242,N_19750);
nand UO_188 (O_188,N_21441,N_20864);
or UO_189 (O_189,N_19833,N_24881);
or UO_190 (O_190,N_22913,N_21768);
xor UO_191 (O_191,N_22769,N_19643);
and UO_192 (O_192,N_21941,N_19926);
xor UO_193 (O_193,N_21508,N_20520);
nand UO_194 (O_194,N_23351,N_23687);
xnor UO_195 (O_195,N_21607,N_23790);
nand UO_196 (O_196,N_21236,N_20415);
nand UO_197 (O_197,N_21409,N_24464);
xor UO_198 (O_198,N_20146,N_23383);
nand UO_199 (O_199,N_18817,N_21958);
nor UO_200 (O_200,N_24782,N_19211);
or UO_201 (O_201,N_18766,N_22520);
nor UO_202 (O_202,N_21118,N_19314);
nor UO_203 (O_203,N_22660,N_22847);
nand UO_204 (O_204,N_20464,N_21197);
nand UO_205 (O_205,N_21769,N_24411);
or UO_206 (O_206,N_20916,N_20753);
nor UO_207 (O_207,N_24367,N_21650);
xnor UO_208 (O_208,N_23401,N_23142);
xor UO_209 (O_209,N_22635,N_24294);
xor UO_210 (O_210,N_23528,N_23032);
nor UO_211 (O_211,N_21631,N_22185);
nand UO_212 (O_212,N_24595,N_24208);
or UO_213 (O_213,N_23431,N_24644);
and UO_214 (O_214,N_21857,N_24906);
or UO_215 (O_215,N_24826,N_21453);
or UO_216 (O_216,N_24996,N_23055);
nand UO_217 (O_217,N_20732,N_24910);
xnor UO_218 (O_218,N_19539,N_21006);
nand UO_219 (O_219,N_22042,N_18837);
nor UO_220 (O_220,N_23825,N_24466);
xnor UO_221 (O_221,N_21960,N_20783);
nor UO_222 (O_222,N_22048,N_20293);
nor UO_223 (O_223,N_19619,N_24289);
and UO_224 (O_224,N_22743,N_22777);
xnor UO_225 (O_225,N_19915,N_20787);
nor UO_226 (O_226,N_19699,N_20580);
nor UO_227 (O_227,N_20290,N_19425);
xnor UO_228 (O_228,N_19700,N_20788);
or UO_229 (O_229,N_24287,N_21850);
and UO_230 (O_230,N_23921,N_19575);
xnor UO_231 (O_231,N_23826,N_20420);
nand UO_232 (O_232,N_20685,N_24564);
and UO_233 (O_233,N_20212,N_22728);
nand UO_234 (O_234,N_20448,N_24193);
or UO_235 (O_235,N_24850,N_24741);
xnor UO_236 (O_236,N_21047,N_23399);
and UO_237 (O_237,N_20192,N_20260);
or UO_238 (O_238,N_23827,N_20429);
and UO_239 (O_239,N_24126,N_24690);
nand UO_240 (O_240,N_24017,N_21526);
nor UO_241 (O_241,N_24532,N_24276);
nand UO_242 (O_242,N_20084,N_24891);
and UO_243 (O_243,N_24298,N_20411);
xnor UO_244 (O_244,N_19289,N_19881);
and UO_245 (O_245,N_21830,N_24018);
and UO_246 (O_246,N_19591,N_19546);
or UO_247 (O_247,N_19208,N_20808);
xor UO_248 (O_248,N_19332,N_22906);
nand UO_249 (O_249,N_23284,N_21599);
xnor UO_250 (O_250,N_22207,N_21461);
or UO_251 (O_251,N_21483,N_22029);
nand UO_252 (O_252,N_24991,N_24633);
or UO_253 (O_253,N_24217,N_19989);
nor UO_254 (O_254,N_21618,N_22392);
and UO_255 (O_255,N_23758,N_23736);
xor UO_256 (O_256,N_24026,N_22623);
nor UO_257 (O_257,N_20958,N_18874);
nand UO_258 (O_258,N_19170,N_23627);
nor UO_259 (O_259,N_20743,N_23091);
xor UO_260 (O_260,N_19788,N_23291);
xor UO_261 (O_261,N_22628,N_22723);
nor UO_262 (O_262,N_20948,N_22378);
nor UO_263 (O_263,N_20579,N_24301);
nand UO_264 (O_264,N_24256,N_23258);
and UO_265 (O_265,N_24964,N_23221);
nand UO_266 (O_266,N_20835,N_21912);
nor UO_267 (O_267,N_24786,N_22684);
nor UO_268 (O_268,N_23033,N_18931);
and UO_269 (O_269,N_24450,N_24123);
or UO_270 (O_270,N_20221,N_24215);
nand UO_271 (O_271,N_23547,N_20697);
and UO_272 (O_272,N_22952,N_20266);
nand UO_273 (O_273,N_19279,N_22587);
xor UO_274 (O_274,N_23046,N_22811);
xnor UO_275 (O_275,N_21744,N_24283);
and UO_276 (O_276,N_24629,N_22725);
and UO_277 (O_277,N_24393,N_21549);
and UO_278 (O_278,N_21931,N_22095);
xnor UO_279 (O_279,N_21754,N_20173);
nand UO_280 (O_280,N_19685,N_24578);
xnor UO_281 (O_281,N_22341,N_20154);
xor UO_282 (O_282,N_21568,N_23428);
nand UO_283 (O_283,N_23314,N_22123);
xor UO_284 (O_284,N_20258,N_24610);
and UO_285 (O_285,N_24574,N_24843);
nor UO_286 (O_286,N_22022,N_24435);
nand UO_287 (O_287,N_21643,N_19261);
or UO_288 (O_288,N_23743,N_23515);
xor UO_289 (O_289,N_20957,N_21054);
nor UO_290 (O_290,N_24547,N_21259);
nand UO_291 (O_291,N_19448,N_21474);
and UO_292 (O_292,N_18910,N_20241);
nor UO_293 (O_293,N_21904,N_20153);
nor UO_294 (O_294,N_19886,N_19104);
xor UO_295 (O_295,N_22821,N_23106);
and UO_296 (O_296,N_22891,N_20534);
nor UO_297 (O_297,N_20603,N_22376);
xor UO_298 (O_298,N_23471,N_20722);
xor UO_299 (O_299,N_24672,N_19450);
and UO_300 (O_300,N_21562,N_22301);
and UO_301 (O_301,N_23922,N_18810);
or UO_302 (O_302,N_21713,N_21610);
nor UO_303 (O_303,N_18964,N_23250);
nor UO_304 (O_304,N_20116,N_19501);
or UO_305 (O_305,N_24392,N_20953);
and UO_306 (O_306,N_21214,N_23603);
or UO_307 (O_307,N_22976,N_19099);
or UO_308 (O_308,N_21094,N_23569);
xor UO_309 (O_309,N_22546,N_20673);
and UO_310 (O_310,N_20046,N_18751);
xor UO_311 (O_311,N_20301,N_21200);
nand UO_312 (O_312,N_21069,N_22693);
or UO_313 (O_313,N_22331,N_18863);
and UO_314 (O_314,N_21968,N_24068);
and UO_315 (O_315,N_21630,N_19166);
or UO_316 (O_316,N_22210,N_23889);
and UO_317 (O_317,N_20535,N_24302);
nand UO_318 (O_318,N_23862,N_19719);
and UO_319 (O_319,N_21127,N_20219);
nand UO_320 (O_320,N_23031,N_18940);
or UO_321 (O_321,N_24935,N_19230);
xor UO_322 (O_322,N_23296,N_21244);
or UO_323 (O_323,N_19838,N_19766);
or UO_324 (O_324,N_22866,N_20122);
xnor UO_325 (O_325,N_23859,N_23232);
nand UO_326 (O_326,N_20112,N_20405);
or UO_327 (O_327,N_20879,N_23113);
and UO_328 (O_328,N_22602,N_23194);
nor UO_329 (O_329,N_23262,N_22625);
or UO_330 (O_330,N_20220,N_23822);
and UO_331 (O_331,N_24836,N_19963);
nor UO_332 (O_332,N_22058,N_22319);
and UO_333 (O_333,N_23948,N_19832);
xnor UO_334 (O_334,N_24284,N_24196);
and UO_335 (O_335,N_21135,N_24765);
or UO_336 (O_336,N_21873,N_21927);
and UO_337 (O_337,N_21588,N_19082);
nand UO_338 (O_338,N_23466,N_23037);
xor UO_339 (O_339,N_21522,N_24915);
nand UO_340 (O_340,N_21352,N_22037);
or UO_341 (O_341,N_20264,N_23153);
or UO_342 (O_342,N_21264,N_24858);
or UO_343 (O_343,N_22892,N_20939);
and UO_344 (O_344,N_20232,N_18777);
nand UO_345 (O_345,N_20842,N_19837);
xnor UO_346 (O_346,N_21211,N_19392);
nor UO_347 (O_347,N_18770,N_20272);
and UO_348 (O_348,N_22509,N_19688);
or UO_349 (O_349,N_21041,N_22505);
nand UO_350 (O_350,N_19792,N_22055);
nand UO_351 (O_351,N_21034,N_22568);
nor UO_352 (O_352,N_19052,N_23760);
nand UO_353 (O_353,N_22985,N_24295);
nand UO_354 (O_354,N_24899,N_20928);
or UO_355 (O_355,N_22070,N_20726);
xnor UO_356 (O_356,N_22992,N_20960);
nand UO_357 (O_357,N_22773,N_19906);
xor UO_358 (O_358,N_21036,N_20636);
nand UO_359 (O_359,N_23805,N_20019);
and UO_360 (O_360,N_22208,N_19522);
nor UO_361 (O_361,N_22146,N_20964);
nand UO_362 (O_362,N_24127,N_19214);
nand UO_363 (O_363,N_23573,N_24675);
xnor UO_364 (O_364,N_21308,N_24112);
nor UO_365 (O_365,N_23853,N_18975);
or UO_366 (O_366,N_23768,N_22656);
xnor UO_367 (O_367,N_18865,N_20688);
nor UO_368 (O_368,N_24105,N_20354);
xor UO_369 (O_369,N_23092,N_23220);
or UO_370 (O_370,N_22372,N_22008);
nand UO_371 (O_371,N_22683,N_19771);
and UO_372 (O_372,N_23298,N_20717);
and UO_373 (O_373,N_18805,N_24175);
nor UO_374 (O_374,N_24546,N_20609);
xnor UO_375 (O_375,N_20064,N_24738);
xor UO_376 (O_376,N_23638,N_19966);
nor UO_377 (O_377,N_23260,N_20247);
or UO_378 (O_378,N_23941,N_24994);
or UO_379 (O_379,N_19013,N_19379);
xnor UO_380 (O_380,N_20035,N_20522);
xor UO_381 (O_381,N_19859,N_21444);
or UO_382 (O_382,N_20215,N_21296);
nand UO_383 (O_383,N_23196,N_19556);
and UO_384 (O_384,N_21171,N_22444);
xnor UO_385 (O_385,N_23903,N_19794);
nor UO_386 (O_386,N_24878,N_21518);
nand UO_387 (O_387,N_20977,N_21013);
xor UO_388 (O_388,N_23389,N_22260);
and UO_389 (O_389,N_24999,N_24928);
nor UO_390 (O_390,N_23882,N_19905);
nand UO_391 (O_391,N_21875,N_22438);
and UO_392 (O_392,N_23211,N_19362);
and UO_393 (O_393,N_21255,N_19300);
xnor UO_394 (O_394,N_21448,N_19823);
xor UO_395 (O_395,N_23361,N_22619);
and UO_396 (O_396,N_21072,N_23710);
or UO_397 (O_397,N_19574,N_22929);
nand UO_398 (O_398,N_19336,N_22791);
or UO_399 (O_399,N_21416,N_20250);
nor UO_400 (O_400,N_22765,N_21295);
xor UO_401 (O_401,N_18973,N_19212);
nor UO_402 (O_402,N_20013,N_19315);
nor UO_403 (O_403,N_20795,N_21813);
or UO_404 (O_404,N_24249,N_23403);
nand UO_405 (O_405,N_18848,N_24240);
xor UO_406 (O_406,N_20184,N_19868);
nand UO_407 (O_407,N_20807,N_22441);
nor UO_408 (O_408,N_22277,N_24029);
or UO_409 (O_409,N_23230,N_19709);
or UO_410 (O_410,N_19459,N_23663);
and UO_411 (O_411,N_21303,N_22933);
or UO_412 (O_412,N_18896,N_20703);
xnor UO_413 (O_413,N_20399,N_23372);
xnor UO_414 (O_414,N_19554,N_23285);
and UO_415 (O_415,N_21575,N_20867);
and UO_416 (O_416,N_24940,N_19274);
xnor UO_417 (O_417,N_24518,N_23879);
xnor UO_418 (O_418,N_18968,N_20336);
nand UO_419 (O_419,N_20126,N_19564);
xor UO_420 (O_420,N_19998,N_24280);
nor UO_421 (O_421,N_21903,N_22720);
or UO_422 (O_422,N_20281,N_23182);
xnor UO_423 (O_423,N_24039,N_24315);
or UO_424 (O_424,N_22018,N_19059);
nor UO_425 (O_425,N_23550,N_23252);
nand UO_426 (O_426,N_21350,N_21866);
and UO_427 (O_427,N_24970,N_23759);
nor UO_428 (O_428,N_20053,N_20321);
nand UO_429 (O_429,N_20785,N_22173);
xnor UO_430 (O_430,N_24918,N_21210);
or UO_431 (O_431,N_24988,N_23349);
xor UO_432 (O_432,N_21910,N_22220);
xor UO_433 (O_433,N_23047,N_21022);
or UO_434 (O_434,N_19250,N_22071);
nor UO_435 (O_435,N_22815,N_20600);
nand UO_436 (O_436,N_19990,N_19036);
or UO_437 (O_437,N_20459,N_23614);
xor UO_438 (O_438,N_19140,N_23895);
nor UO_439 (O_439,N_23875,N_24013);
and UO_440 (O_440,N_22532,N_21577);
xor UO_441 (O_441,N_19993,N_19169);
and UO_442 (O_442,N_23890,N_23730);
nor UO_443 (O_443,N_21029,N_19087);
xnor UO_444 (O_444,N_21062,N_24947);
and UO_445 (O_445,N_24154,N_22292);
or UO_446 (O_446,N_19533,N_20532);
xor UO_447 (O_447,N_20476,N_18860);
nor UO_448 (O_448,N_23313,N_24260);
nand UO_449 (O_449,N_23511,N_20142);
nand UO_450 (O_450,N_24598,N_19666);
or UO_451 (O_451,N_24145,N_19493);
or UO_452 (O_452,N_19049,N_21645);
and UO_453 (O_453,N_19296,N_24321);
and UO_454 (O_454,N_19186,N_23487);
and UO_455 (O_455,N_19563,N_24370);
and UO_456 (O_456,N_23133,N_21090);
nor UO_457 (O_457,N_22415,N_21675);
xnor UO_458 (O_458,N_20822,N_19146);
and UO_459 (O_459,N_19470,N_22281);
nand UO_460 (O_460,N_22456,N_24452);
nand UO_461 (O_461,N_24758,N_22867);
or UO_462 (O_462,N_22135,N_18984);
nand UO_463 (O_463,N_19641,N_23253);
and UO_464 (O_464,N_23322,N_22965);
or UO_465 (O_465,N_21359,N_20955);
nand UO_466 (O_466,N_21435,N_23427);
nor UO_467 (O_467,N_22746,N_23385);
or UO_468 (O_468,N_19515,N_21563);
and UO_469 (O_469,N_22167,N_23910);
and UO_470 (O_470,N_21726,N_24865);
nand UO_471 (O_471,N_19851,N_19410);
nor UO_472 (O_472,N_19468,N_24049);
or UO_473 (O_473,N_24785,N_24562);
and UO_474 (O_474,N_22764,N_20905);
nor UO_475 (O_475,N_19421,N_23447);
nor UO_476 (O_476,N_24969,N_23559);
xor UO_477 (O_477,N_19577,N_19318);
and UO_478 (O_478,N_22465,N_22830);
or UO_479 (O_479,N_20714,N_19680);
nor UO_480 (O_480,N_20208,N_21798);
nor UO_481 (O_481,N_24953,N_24591);
xnor UO_482 (O_482,N_20437,N_22573);
and UO_483 (O_483,N_23327,N_21185);
nand UO_484 (O_484,N_21113,N_24925);
nand UO_485 (O_485,N_23208,N_23473);
nand UO_486 (O_486,N_24063,N_23123);
nand UO_487 (O_487,N_20101,N_24254);
or UO_488 (O_488,N_18997,N_19108);
or UO_489 (O_489,N_18844,N_19582);
or UO_490 (O_490,N_18824,N_22468);
nor UO_491 (O_491,N_23004,N_23460);
xnor UO_492 (O_492,N_20729,N_19106);
or UO_493 (O_493,N_22857,N_20853);
nand UO_494 (O_494,N_20512,N_23064);
or UO_495 (O_495,N_22542,N_24535);
nor UO_496 (O_496,N_19085,N_22594);
nor UO_497 (O_497,N_19128,N_20470);
xnor UO_498 (O_498,N_21180,N_22963);
xnor UO_499 (O_499,N_22025,N_23934);
and UO_500 (O_500,N_19578,N_21218);
nand UO_501 (O_501,N_20027,N_23006);
xor UO_502 (O_502,N_24646,N_22560);
nand UO_503 (O_503,N_21566,N_20992);
xnor UO_504 (O_504,N_20474,N_24902);
or UO_505 (O_505,N_24628,N_20625);
nor UO_506 (O_506,N_19716,N_20615);
nand UO_507 (O_507,N_21157,N_21933);
or UO_508 (O_508,N_24877,N_24199);
and UO_509 (O_509,N_23504,N_24893);
nand UO_510 (O_510,N_20151,N_21479);
nand UO_511 (O_511,N_23158,N_20896);
xnor UO_512 (O_512,N_21692,N_23352);
nor UO_513 (O_513,N_21433,N_24757);
and UO_514 (O_514,N_22971,N_19940);
or UO_515 (O_515,N_23908,N_22407);
and UO_516 (O_516,N_24654,N_20741);
nand UO_517 (O_517,N_24430,N_23947);
xor UO_518 (O_518,N_23848,N_23765);
and UO_519 (O_519,N_22592,N_23397);
or UO_520 (O_520,N_23304,N_24181);
or UO_521 (O_521,N_22237,N_20680);
nand UO_522 (O_522,N_24660,N_21025);
nand UO_523 (O_523,N_24386,N_23588);
xor UO_524 (O_524,N_21421,N_20398);
xnor UO_525 (O_525,N_21601,N_22885);
nor UO_526 (O_526,N_19805,N_24417);
nand UO_527 (O_527,N_24638,N_19934);
and UO_528 (O_528,N_19387,N_19413);
nand UO_529 (O_529,N_20376,N_23493);
nand UO_530 (O_530,N_22564,N_18866);
or UO_531 (O_531,N_24005,N_22702);
xnor UO_532 (O_532,N_18905,N_20963);
or UO_533 (O_533,N_21111,N_21506);
or UO_534 (O_534,N_19791,N_18945);
xor UO_535 (O_535,N_19356,N_19046);
nor UO_536 (O_536,N_21260,N_24985);
nor UO_537 (O_537,N_24194,N_23734);
nor UO_538 (O_538,N_21053,N_22340);
xnor UO_539 (O_539,N_22601,N_20134);
nor UO_540 (O_540,N_22670,N_21394);
and UO_541 (O_541,N_23809,N_22132);
or UO_542 (O_542,N_20251,N_22804);
nand UO_543 (O_543,N_22240,N_18930);
xnor UO_544 (O_544,N_23733,N_23448);
or UO_545 (O_545,N_20725,N_24818);
xnor UO_546 (O_546,N_22789,N_23433);
nor UO_547 (O_547,N_22259,N_18826);
or UO_548 (O_548,N_18812,N_24368);
and UO_549 (O_549,N_23104,N_23755);
or UO_550 (O_550,N_24369,N_21824);
xnor UO_551 (O_551,N_20983,N_23754);
nand UO_552 (O_552,N_20255,N_23317);
xnor UO_553 (O_553,N_23017,N_19724);
nor UO_554 (O_554,N_24548,N_20631);
nand UO_555 (O_555,N_20630,N_24042);
nand UO_556 (O_556,N_22597,N_20924);
or UO_557 (O_557,N_19977,N_19759);
nand UO_558 (O_558,N_22828,N_22349);
nor UO_559 (O_559,N_24230,N_24073);
nand UO_560 (O_560,N_22106,N_23245);
xor UO_561 (O_561,N_22390,N_21862);
nand UO_562 (O_562,N_22442,N_20728);
or UO_563 (O_563,N_23362,N_24875);
nand UO_564 (O_564,N_21331,N_24787);
nor UO_565 (O_565,N_19485,N_20227);
nor UO_566 (O_566,N_22943,N_24982);
and UO_567 (O_567,N_23829,N_21551);
and UO_568 (O_568,N_21455,N_23919);
or UO_569 (O_569,N_21251,N_23029);
nand UO_570 (O_570,N_23508,N_22862);
xor UO_571 (O_571,N_24752,N_19799);
xnor UO_572 (O_572,N_19403,N_19116);
and UO_573 (O_573,N_19151,N_23568);
or UO_574 (O_574,N_24615,N_24036);
or UO_575 (O_575,N_21932,N_19592);
or UO_576 (O_576,N_21098,N_19071);
nor UO_577 (O_577,N_21361,N_20902);
nand UO_578 (O_578,N_19237,N_20740);
xor UO_579 (O_579,N_23516,N_24636);
nand UO_580 (O_580,N_20036,N_23580);
nor UO_581 (O_581,N_18806,N_19946);
xnor UO_582 (O_582,N_23572,N_19216);
nand UO_583 (O_583,N_20730,N_19431);
xnor UO_584 (O_584,N_22329,N_23608);
xnor UO_585 (O_585,N_19360,N_19035);
and UO_586 (O_586,N_23381,N_20206);
nand UO_587 (O_587,N_20480,N_24890);
nand UO_588 (O_588,N_23617,N_20674);
xor UO_589 (O_589,N_24530,N_24550);
nand UO_590 (O_590,N_22216,N_21653);
nand UO_591 (O_591,N_23651,N_22890);
and UO_592 (O_592,N_22082,N_23688);
or UO_593 (O_593,N_21079,N_21801);
or UO_594 (O_594,N_19246,N_21124);
nor UO_595 (O_595,N_23154,N_24035);
and UO_596 (O_596,N_22816,N_21139);
nand UO_597 (O_597,N_22550,N_24745);
and UO_598 (O_598,N_21665,N_21774);
xor UO_599 (O_599,N_19093,N_24604);
nand UO_600 (O_600,N_24388,N_24076);
or UO_601 (O_601,N_24596,N_22271);
and UO_602 (O_602,N_21281,N_22807);
or UO_603 (O_603,N_21540,N_24889);
and UO_604 (O_604,N_19321,N_24027);
and UO_605 (O_605,N_21363,N_19630);
nor UO_606 (O_606,N_23356,N_20510);
xor UO_607 (O_607,N_21081,N_19232);
or UO_608 (O_608,N_18969,N_21907);
xnor UO_609 (O_609,N_20384,N_22473);
xor UO_610 (O_610,N_20552,N_23127);
nand UO_611 (O_611,N_20789,N_22267);
nor UO_612 (O_612,N_19658,N_19199);
and UO_613 (O_613,N_24271,N_20032);
xor UO_614 (O_614,N_23575,N_23810);
nand UO_615 (O_615,N_24541,N_23357);
and UO_616 (O_616,N_18934,N_21194);
nor UO_617 (O_617,N_23436,N_24116);
nand UO_618 (O_618,N_18881,N_24346);
and UO_619 (O_619,N_23967,N_21714);
and UO_620 (O_620,N_22545,N_20771);
or UO_621 (O_621,N_23950,N_21136);
nand UO_622 (O_622,N_23554,N_21908);
nor UO_623 (O_623,N_20229,N_21112);
or UO_624 (O_624,N_20809,N_23691);
nand UO_625 (O_625,N_19445,N_22264);
and UO_626 (O_626,N_23881,N_24586);
and UO_627 (O_627,N_21524,N_21626);
nor UO_628 (O_628,N_19876,N_21354);
or UO_629 (O_629,N_20403,N_21877);
xnor UO_630 (O_630,N_19987,N_22286);
xor UO_631 (O_631,N_19769,N_19550);
and UO_632 (O_632,N_21838,N_22876);
or UO_633 (O_633,N_20854,N_18758);
xnor UO_634 (O_634,N_19953,N_22351);
nor UO_635 (O_635,N_21007,N_21815);
xor UO_636 (O_636,N_20889,N_18761);
and UO_637 (O_637,N_20851,N_18902);
and UO_638 (O_638,N_20311,N_22704);
nor UO_639 (O_639,N_24492,N_21215);
nor UO_640 (O_640,N_24328,N_20419);
or UO_641 (O_641,N_20371,N_20875);
xnor UO_642 (O_642,N_23574,N_19932);
nor UO_643 (O_643,N_21065,N_23169);
and UO_644 (O_644,N_21240,N_24565);
nand UO_645 (O_645,N_21179,N_24898);
xnor UO_646 (O_646,N_19033,N_19505);
nand UO_647 (O_647,N_19648,N_20706);
and UO_648 (O_648,N_22366,N_19921);
xnor UO_649 (O_649,N_19477,N_22767);
or UO_650 (O_650,N_24955,N_18979);
nor UO_651 (O_651,N_18774,N_23486);
xnor UO_652 (O_652,N_19708,N_21743);
or UO_653 (O_653,N_22787,N_20616);
nand UO_654 (O_654,N_20776,N_23778);
xor UO_655 (O_655,N_20517,N_21005);
or UO_656 (O_656,N_22007,N_19901);
and UO_657 (O_657,N_24440,N_20014);
nand UO_658 (O_658,N_22266,N_24959);
and UO_659 (O_659,N_19499,N_21107);
nand UO_660 (O_660,N_22051,N_24101);
or UO_661 (O_661,N_24405,N_20361);
nor UO_662 (O_662,N_24859,N_21087);
xor UO_663 (O_663,N_20516,N_23593);
nand UO_664 (O_664,N_19095,N_21998);
xnor UO_665 (O_665,N_20548,N_23844);
xor UO_666 (O_666,N_19002,N_24247);
nand UO_667 (O_667,N_22308,N_24834);
or UO_668 (O_668,N_23268,N_20107);
nor UO_669 (O_669,N_23079,N_22873);
xnor UO_670 (O_670,N_19810,N_21988);
nand UO_671 (O_671,N_19441,N_20216);
nor UO_672 (O_672,N_19626,N_20009);
and UO_673 (O_673,N_21611,N_22458);
or UO_674 (O_674,N_20038,N_24688);
and UO_675 (O_675,N_22419,N_24410);
nand UO_676 (O_676,N_24735,N_21940);
nand UO_677 (O_677,N_24186,N_19583);
nor UO_678 (O_678,N_22273,N_22405);
or UO_679 (O_679,N_19939,N_23631);
xnor UO_680 (O_680,N_24028,N_19964);
or UO_681 (O_681,N_23125,N_20066);
xnor UO_682 (O_682,N_20727,N_19891);
nor UO_683 (O_683,N_19319,N_22606);
or UO_684 (O_684,N_23699,N_23610);
nor UO_685 (O_685,N_19679,N_24047);
xor UO_686 (O_686,N_23728,N_24882);
nor UO_687 (O_687,N_20489,N_22779);
or UO_688 (O_688,N_20098,N_23929);
or UO_689 (O_689,N_19561,N_24759);
or UO_690 (O_690,N_21570,N_19462);
nand UO_691 (O_691,N_19790,N_19465);
and UO_692 (O_692,N_22138,N_23774);
nand UO_693 (O_693,N_20643,N_21372);
or UO_694 (O_694,N_24762,N_20110);
or UO_695 (O_695,N_21033,N_19607);
or UO_696 (O_696,N_21595,N_21710);
nand UO_697 (O_697,N_20130,N_23785);
xnor UO_698 (O_698,N_22035,N_20458);
xnor UO_699 (O_699,N_22482,N_22792);
and UO_700 (O_700,N_22293,N_24493);
nor UO_701 (O_701,N_23019,N_19677);
or UO_702 (O_702,N_22707,N_19887);
and UO_703 (O_703,N_24442,N_19342);
nand UO_704 (O_704,N_19194,N_20526);
or UO_705 (O_705,N_19969,N_22417);
xnor UO_706 (O_706,N_18996,N_21561);
nand UO_707 (O_707,N_22650,N_23187);
and UO_708 (O_708,N_20467,N_23179);
xor UO_709 (O_709,N_21145,N_21542);
nor UO_710 (O_710,N_21917,N_24936);
or UO_711 (O_711,N_23462,N_24352);
nor UO_712 (O_712,N_21431,N_21963);
nor UO_713 (O_713,N_24823,N_20541);
or UO_714 (O_714,N_23985,N_24077);
or UO_715 (O_715,N_23426,N_22411);
or UO_716 (O_716,N_21503,N_22307);
or UO_717 (O_717,N_19836,N_24099);
xnor UO_718 (O_718,N_19266,N_18833);
nand UO_719 (O_719,N_20573,N_23557);
or UO_720 (O_720,N_19174,N_24463);
nand UO_721 (O_721,N_22006,N_23742);
xnor UO_722 (O_722,N_24161,N_23505);
and UO_723 (O_723,N_20640,N_23111);
nand UO_724 (O_724,N_19304,N_23552);
nor UO_725 (O_725,N_22671,N_24236);
nand UO_726 (O_726,N_19711,N_22227);
or UO_727 (O_727,N_20554,N_18907);
or UO_728 (O_728,N_24623,N_20340);
nand UO_729 (O_729,N_20650,N_18900);
nor UO_730 (O_730,N_23666,N_21831);
nor UO_731 (O_731,N_20075,N_23797);
xor UO_732 (O_732,N_23078,N_23097);
nand UO_733 (O_733,N_20745,N_24849);
nor UO_734 (O_734,N_20176,N_23420);
xnor UO_735 (O_735,N_20447,N_19786);
xnor UO_736 (O_736,N_19062,N_19909);
xnor UO_737 (O_737,N_21225,N_24783);
nor UO_738 (O_738,N_18807,N_20042);
nand UO_739 (O_739,N_19532,N_21557);
nand UO_740 (O_740,N_23139,N_24291);
nor UO_741 (O_741,N_24066,N_21429);
nor UO_742 (O_742,N_24286,N_23788);
or UO_743 (O_743,N_23576,N_20908);
xor UO_744 (O_744,N_19222,N_21026);
or UO_745 (O_745,N_19593,N_23987);
nor UO_746 (O_746,N_22849,N_21327);
and UO_747 (O_747,N_20656,N_23094);
xnor UO_748 (O_748,N_20550,N_24052);
and UO_749 (O_749,N_20664,N_22059);
nand UO_750 (O_750,N_19024,N_19278);
xnor UO_751 (O_751,N_21096,N_18923);
or UO_752 (O_752,N_20076,N_21024);
xnor UO_753 (O_753,N_19614,N_22621);
or UO_754 (O_754,N_21979,N_22839);
or UO_755 (O_755,N_22663,N_19741);
nand UO_756 (O_756,N_19590,N_23622);
xor UO_757 (O_757,N_22757,N_21076);
and UO_758 (O_758,N_24560,N_24325);
or UO_759 (O_759,N_21187,N_19736);
nor UO_760 (O_760,N_20030,N_19506);
or UO_761 (O_761,N_20883,N_20649);
nand UO_762 (O_762,N_19600,N_22881);
or UO_763 (O_763,N_21449,N_24444);
or UO_764 (O_764,N_20540,N_22763);
or UO_765 (O_765,N_23749,N_19925);
and UO_766 (O_766,N_19047,N_21749);
nor UO_767 (O_767,N_24912,N_22072);
and UO_768 (O_768,N_22806,N_23946);
nor UO_769 (O_769,N_23525,N_23521);
nand UO_770 (O_770,N_24805,N_22190);
nand UO_771 (O_771,N_22245,N_23157);
nand UO_772 (O_772,N_23446,N_19311);
nand UO_773 (O_773,N_22242,N_21014);
nor UO_774 (O_774,N_24446,N_21492);
nor UO_775 (O_775,N_24172,N_24223);
nand UO_776 (O_776,N_23149,N_19954);
nor UO_777 (O_777,N_19262,N_19547);
or UO_778 (O_778,N_24736,N_20318);
nand UO_779 (O_779,N_23911,N_21537);
xnor UO_780 (O_780,N_24259,N_23277);
nor UO_781 (O_781,N_21012,N_22348);
nand UO_782 (O_782,N_21430,N_21913);
nand UO_783 (O_783,N_23767,N_24170);
nor UO_784 (O_784,N_19331,N_22032);
xnor UO_785 (O_785,N_19776,N_22403);
and UO_786 (O_786,N_21893,N_24051);
nand UO_787 (O_787,N_20335,N_23015);
nand UO_788 (O_788,N_22309,N_23130);
xnor UO_789 (O_789,N_24945,N_20275);
and UO_790 (O_790,N_19055,N_19587);
or UO_791 (O_791,N_21440,N_24205);
and UO_792 (O_792,N_20422,N_20179);
nor UO_793 (O_793,N_22443,N_24704);
nand UO_794 (O_794,N_19455,N_19486);
nand UO_795 (O_795,N_19843,N_24443);
and UO_796 (O_796,N_19762,N_18846);
nor UO_797 (O_797,N_19748,N_20026);
nor UO_798 (O_798,N_20792,N_20751);
or UO_799 (O_799,N_23162,N_21114);
nor UO_800 (O_800,N_21867,N_23163);
or UO_801 (O_801,N_22884,N_24707);
and UO_802 (O_802,N_20016,N_21015);
xnor UO_803 (O_803,N_21246,N_22360);
or UO_804 (O_804,N_19025,N_19615);
nor UO_805 (O_805,N_22480,N_22452);
nor UO_806 (O_806,N_20423,N_22904);
xnor UO_807 (O_807,N_20966,N_22882);
or UO_808 (O_808,N_24117,N_24220);
nor UO_809 (O_809,N_19467,N_19238);
and UO_810 (O_810,N_23753,N_24998);
nor UO_811 (O_811,N_18791,N_19241);
nor UO_812 (O_812,N_21962,N_18936);
or UO_813 (O_813,N_24983,N_18955);
nor UO_814 (O_814,N_20531,N_24371);
and UO_815 (O_815,N_23982,N_21238);
nand UO_816 (O_816,N_22843,N_22522);
or UO_817 (O_817,N_21740,N_24700);
nor UO_818 (O_818,N_20979,N_24508);
nand UO_819 (O_819,N_21293,N_21624);
or UO_820 (O_820,N_20605,N_23566);
nor UO_821 (O_821,N_21450,N_23184);
and UO_822 (O_822,N_20954,N_22250);
nand UO_823 (O_823,N_21089,N_19348);
xnor UO_824 (O_824,N_23497,N_21312);
nor UO_825 (O_825,N_18767,N_22437);
and UO_826 (O_826,N_24432,N_20157);
or UO_827 (O_827,N_24706,N_20779);
nand UO_828 (O_828,N_22610,N_22261);
nor UO_829 (O_829,N_18962,N_22368);
or UO_830 (O_830,N_21184,N_22988);
and UO_831 (O_831,N_24685,N_22636);
or UO_832 (O_832,N_20710,N_21016);
xnor UO_833 (O_833,N_23458,N_20353);
nor UO_834 (O_834,N_20428,N_23541);
and UO_835 (O_835,N_22896,N_23145);
xor UO_836 (O_836,N_23852,N_23368);
nand UO_837 (O_837,N_21291,N_19073);
and UO_838 (O_838,N_22507,N_22894);
nand UO_839 (O_839,N_19941,N_24337);
and UO_840 (O_840,N_20007,N_24447);
or UO_841 (O_841,N_23714,N_22877);
nor UO_842 (O_842,N_22932,N_23254);
xnor UO_843 (O_843,N_21558,N_20226);
nand UO_844 (O_844,N_20170,N_24791);
xor UO_845 (O_845,N_24743,N_23997);
or UO_846 (O_846,N_21482,N_22129);
nand UO_847 (O_847,N_20425,N_21275);
or UO_848 (O_848,N_24978,N_19312);
nor UO_849 (O_849,N_21955,N_22049);
xor UO_850 (O_850,N_20444,N_22603);
and UO_851 (O_851,N_20599,N_23553);
or UO_852 (O_852,N_22658,N_21972);
nand UO_853 (O_853,N_22320,N_21038);
nor UO_854 (O_854,N_22688,N_20465);
and UO_855 (O_855,N_23858,N_23434);
and UO_856 (O_856,N_19610,N_22381);
and UO_857 (O_857,N_20951,N_20925);
nand UO_858 (O_858,N_24222,N_19432);
xor UO_859 (O_859,N_19405,N_21949);
nor UO_860 (O_860,N_21552,N_21035);
nand UO_861 (O_861,N_21131,N_20218);
and UO_862 (O_862,N_24822,N_19565);
xor UO_863 (O_863,N_22436,N_24922);
nand UO_864 (O_864,N_21426,N_24363);
nor UO_865 (O_865,N_22296,N_21729);
xnor UO_866 (O_866,N_24290,N_19487);
xnor UO_867 (O_867,N_22820,N_24382);
or UO_868 (O_868,N_24645,N_21802);
or UO_869 (O_869,N_19043,N_22096);
and UO_870 (O_870,N_23831,N_23526);
xor UO_871 (O_871,N_22026,N_21401);
nand UO_872 (O_872,N_19031,N_19411);
and UO_873 (O_873,N_23010,N_24226);
or UO_874 (O_874,N_20196,N_24357);
xor UO_875 (O_875,N_19783,N_22944);
and UO_876 (O_876,N_22327,N_22170);
nor UO_877 (O_877,N_24016,N_19021);
nand UO_878 (O_878,N_22194,N_20862);
nand UO_879 (O_879,N_23747,N_21258);
or UO_880 (O_880,N_23049,N_20388);
or UO_881 (O_881,N_24514,N_20087);
or UO_882 (O_882,N_23007,N_21276);
and UO_883 (O_883,N_22162,N_21888);
and UO_884 (O_884,N_21341,N_22870);
or UO_885 (O_885,N_21326,N_23944);
and UO_886 (O_886,N_21103,N_24793);
nor UO_887 (O_887,N_21186,N_22841);
nand UO_888 (O_888,N_22255,N_23792);
and UO_889 (O_889,N_24424,N_23932);
and UO_890 (O_890,N_19682,N_21423);
and UO_891 (O_891,N_22345,N_23703);
and UO_892 (O_892,N_21371,N_23332);
xnor UO_893 (O_893,N_23949,N_18885);
xor UO_894 (O_894,N_19531,N_24056);
xor UO_895 (O_895,N_22682,N_19306);
and UO_896 (O_896,N_18912,N_24094);
or UO_897 (O_897,N_19686,N_21858);
and UO_898 (O_898,N_22928,N_24350);
nor UO_899 (O_899,N_19968,N_24523);
or UO_900 (O_900,N_23025,N_23148);
and UO_901 (O_901,N_20922,N_20621);
and UO_902 (O_902,N_18783,N_22247);
nor UO_903 (O_903,N_23281,N_24776);
xor UO_904 (O_904,N_21381,N_23301);
xor UO_905 (O_905,N_23720,N_21939);
and UO_906 (O_906,N_23457,N_24534);
or UO_907 (O_907,N_19944,N_24195);
or UO_908 (O_908,N_23093,N_19008);
xor UO_909 (O_909,N_19176,N_20627);
nor UO_910 (O_910,N_21502,N_24520);
nand UO_911 (O_911,N_19882,N_19798);
xor UO_912 (O_912,N_22449,N_19156);
nor UO_913 (O_913,N_21693,N_24933);
xor UO_914 (O_914,N_21948,N_23067);
or UO_915 (O_915,N_21344,N_24800);
or UO_916 (O_916,N_24045,N_19086);
xor UO_917 (O_917,N_21397,N_20846);
nor UO_918 (O_918,N_21088,N_23272);
or UO_919 (O_919,N_21728,N_22861);
xnor UO_920 (O_920,N_23325,N_20099);
nor UO_921 (O_921,N_23701,N_23558);
or UO_922 (O_922,N_22611,N_23718);
xnor UO_923 (O_923,N_20794,N_23763);
or UO_924 (O_924,N_23321,N_23925);
xor UO_925 (O_925,N_23983,N_23570);
nor UO_926 (O_926,N_24821,N_20364);
nor UO_927 (O_927,N_21918,N_18911);
or UO_928 (O_928,N_23854,N_20989);
nand UO_929 (O_929,N_22687,N_20986);
nand UO_930 (O_930,N_20800,N_24602);
nand UO_931 (O_931,N_23068,N_19884);
or UO_932 (O_932,N_22012,N_19136);
or UO_933 (O_933,N_23725,N_24914);
nand UO_934 (O_934,N_19772,N_21733);
or UO_935 (O_935,N_19635,N_19273);
or UO_936 (O_936,N_23804,N_20500);
nor UO_937 (O_937,N_20659,N_22961);
xnor UO_938 (O_938,N_22824,N_19777);
or UO_939 (O_939,N_19057,N_21414);
and UO_940 (O_940,N_24798,N_20556);
nand UO_941 (O_941,N_19299,N_23936);
or UO_942 (O_942,N_23864,N_24904);
and UO_943 (O_943,N_20141,N_19795);
and UO_944 (O_944,N_24561,N_22879);
and UO_945 (O_945,N_21619,N_22955);
and UO_946 (O_946,N_24742,N_18878);
nor UO_947 (O_947,N_22142,N_23069);
nor UO_948 (O_948,N_21646,N_20976);
or UO_949 (O_949,N_22524,N_22315);
and UO_950 (O_950,N_22498,N_19406);
and UO_951 (O_951,N_20124,N_23203);
nand UO_952 (O_952,N_23847,N_21898);
or UO_953 (O_953,N_19858,N_24573);
or UO_954 (O_954,N_24129,N_23178);
nand UO_955 (O_955,N_20781,N_22501);
nand UO_956 (O_956,N_19358,N_20372);
xor UO_957 (O_957,N_19704,N_21790);
nor UO_958 (O_958,N_22580,N_23878);
xor UO_959 (O_959,N_19461,N_23680);
and UO_960 (O_960,N_21230,N_21494);
or UO_961 (O_961,N_20906,N_23565);
or UO_962 (O_962,N_24020,N_23814);
nor UO_963 (O_963,N_21883,N_20760);
nor UO_964 (O_964,N_22262,N_23897);
and UO_965 (O_965,N_19524,N_20460);
nand UO_966 (O_966,N_22064,N_21309);
nor UO_967 (O_967,N_24833,N_18756);
nand UO_968 (O_968,N_23449,N_21762);
nor UO_969 (O_969,N_24810,N_21261);
nand UO_970 (O_970,N_20628,N_19537);
nand UO_971 (O_971,N_23464,N_20365);
nand UO_972 (O_972,N_23951,N_24870);
nor UO_973 (O_973,N_20439,N_19519);
nand UO_974 (O_974,N_21436,N_23437);
or UO_975 (O_975,N_20029,N_19126);
and UO_976 (O_976,N_21935,N_22783);
or UO_977 (O_977,N_22041,N_22629);
nand UO_978 (O_978,N_19452,N_24924);
or UO_979 (O_979,N_24642,N_23970);
or UO_980 (O_980,N_20648,N_19430);
nand UO_981 (O_981,N_22433,N_19138);
xnor UO_982 (O_982,N_24917,N_24083);
xnor UO_983 (O_983,N_24583,N_24163);
xor UO_984 (O_984,N_23278,N_22742);
or UO_985 (O_985,N_21365,N_23350);
xnor UO_986 (O_986,N_20546,N_20197);
nand UO_987 (O_987,N_21447,N_19365);
nand UO_988 (O_988,N_22187,N_23315);
nor UO_989 (O_989,N_20494,N_24937);
nor UO_990 (O_990,N_21349,N_24314);
nand UO_991 (O_991,N_18901,N_23344);
or UO_992 (O_992,N_20923,N_22298);
nor UO_993 (O_993,N_20270,N_20533);
nor UO_994 (O_994,N_20926,N_19758);
xor UO_995 (O_995,N_23794,N_19390);
nand UO_996 (O_996,N_19153,N_21699);
or UO_997 (O_997,N_20268,N_19895);
or UO_998 (O_998,N_19345,N_19809);
or UO_999 (O_999,N_19847,N_23308);
or UO_1000 (O_1000,N_24232,N_22141);
xor UO_1001 (O_1001,N_20265,N_24778);
nand UO_1002 (O_1002,N_22276,N_23363);
nor UO_1003 (O_1003,N_23562,N_19144);
xnor UO_1004 (O_1004,N_19302,N_22131);
nand UO_1005 (O_1005,N_21651,N_22196);
nand UO_1006 (O_1006,N_22949,N_24829);
and UO_1007 (O_1007,N_20045,N_20826);
nand UO_1008 (O_1008,N_23695,N_19856);
nor UO_1009 (O_1009,N_22859,N_23379);
and UO_1010 (O_1010,N_23952,N_24923);
xor UO_1011 (O_1011,N_20559,N_21392);
nand UO_1012 (O_1012,N_24768,N_19101);
nor UO_1013 (O_1013,N_19344,N_19456);
and UO_1014 (O_1014,N_20876,N_20897);
nand UO_1015 (O_1015,N_19623,N_22101);
nor UO_1016 (O_1016,N_23976,N_22463);
and UO_1017 (O_1017,N_23347,N_22993);
nand UO_1018 (O_1018,N_20655,N_20699);
nand UO_1019 (O_1019,N_21282,N_23808);
nand UO_1020 (O_1020,N_19638,N_18851);
xor UO_1021 (O_1021,N_19628,N_24122);
nand UO_1022 (O_1022,N_24863,N_21254);
nand UO_1023 (O_1023,N_21091,N_21080);
or UO_1024 (O_1024,N_20553,N_24059);
xor UO_1025 (O_1025,N_22069,N_22364);
nand UO_1026 (O_1026,N_22299,N_21639);
and UO_1027 (O_1027,N_24570,N_23928);
or UO_1028 (O_1028,N_24587,N_24739);
and UO_1029 (O_1029,N_20525,N_19620);
xor UO_1030 (O_1030,N_23081,N_24468);
nand UO_1031 (O_1031,N_24317,N_19316);
nor UO_1032 (O_1032,N_21143,N_23439);
nor UO_1033 (O_1033,N_24931,N_23524);
or UO_1034 (O_1034,N_20040,N_20750);
xnor UO_1035 (O_1035,N_21860,N_20331);
or UO_1036 (O_1036,N_19007,N_23679);
or UO_1037 (O_1037,N_19005,N_21358);
and UO_1038 (O_1038,N_23336,N_18971);
xnor UO_1039 (O_1039,N_19094,N_24506);
and UO_1040 (O_1040,N_24718,N_23035);
nor UO_1041 (O_1041,N_18861,N_22040);
xnor UO_1042 (O_1042,N_23454,N_21245);
or UO_1043 (O_1043,N_24984,N_21212);
xnor UO_1044 (O_1044,N_24942,N_20152);
or UO_1045 (O_1045,N_24231,N_24809);
xor UO_1046 (O_1046,N_20067,N_23945);
and UO_1047 (O_1047,N_21722,N_23787);
nand UO_1048 (O_1048,N_20502,N_21270);
or UO_1049 (O_1049,N_20074,N_23650);
nor UO_1050 (O_1050,N_18919,N_24089);
and UO_1051 (O_1051,N_23072,N_24797);
nor UO_1052 (O_1052,N_23226,N_24869);
xor UO_1053 (O_1053,N_21298,N_19965);
and UO_1054 (O_1054,N_23239,N_24431);
xnor UO_1055 (O_1055,N_19584,N_22143);
xnor UO_1056 (O_1056,N_24211,N_20082);
nor UO_1057 (O_1057,N_21307,N_24394);
nor UO_1058 (O_1058,N_18943,N_22038);
or UO_1059 (O_1059,N_21773,N_18830);
and UO_1060 (O_1060,N_18950,N_24082);
nand UO_1061 (O_1061,N_18906,N_22469);
xor UO_1062 (O_1062,N_18875,N_22079);
nand UO_1063 (O_1063,N_23107,N_22584);
and UO_1064 (O_1064,N_23939,N_21523);
nor UO_1065 (O_1065,N_20877,N_24986);
and UO_1066 (O_1066,N_23609,N_20274);
and UO_1067 (O_1067,N_21207,N_24505);
xor UO_1068 (O_1068,N_22530,N_22057);
nand UO_1069 (O_1069,N_20128,N_21828);
nand UO_1070 (O_1070,N_22631,N_23456);
or UO_1071 (O_1071,N_20780,N_20764);
nor UO_1072 (O_1072,N_22477,N_22609);
and UO_1073 (O_1073,N_19040,N_23777);
xor UO_1074 (O_1074,N_24580,N_21242);
and UO_1075 (O_1075,N_20117,N_19054);
or UO_1076 (O_1076,N_20718,N_19848);
nor UO_1077 (O_1077,N_21199,N_23533);
or UO_1078 (O_1078,N_20899,N_24389);
or UO_1079 (O_1079,N_20191,N_21707);
and UO_1080 (O_1080,N_24668,N_21471);
nand UO_1081 (O_1081,N_20455,N_24777);
and UO_1082 (O_1082,N_19454,N_21055);
or UO_1083 (O_1083,N_19164,N_18929);
and UO_1084 (O_1084,N_23920,N_20791);
nor UO_1085 (O_1085,N_21785,N_19598);
and UO_1086 (O_1086,N_23175,N_22659);
xor UO_1087 (O_1087,N_21140,N_19399);
nor UO_1088 (O_1088,N_23977,N_21547);
xor UO_1089 (O_1089,N_23668,N_19644);
nor UO_1090 (O_1090,N_22782,N_20187);
nor UO_1091 (O_1091,N_22183,N_20684);
nor UO_1092 (O_1092,N_23185,N_21205);
nand UO_1093 (O_1093,N_23883,N_22013);
nand UO_1094 (O_1094,N_22681,N_19091);
and UO_1095 (O_1095,N_22569,N_19518);
nand UO_1096 (O_1096,N_24001,N_22499);
nor UO_1097 (O_1097,N_24219,N_23819);
xor UO_1098 (O_1098,N_23131,N_21525);
and UO_1099 (O_1099,N_22595,N_18889);
nor UO_1100 (O_1100,N_20366,N_24731);
nand UO_1101 (O_1101,N_23112,N_21408);
xnor UO_1102 (O_1102,N_19081,N_24961);
xnor UO_1103 (O_1103,N_19072,N_22278);
nor UO_1104 (O_1104,N_24140,N_19409);
or UO_1105 (O_1105,N_21586,N_22063);
nand UO_1106 (O_1106,N_19429,N_24490);
or UO_1107 (O_1107,N_21761,N_24963);
nand UO_1108 (O_1108,N_24847,N_22251);
nand UO_1109 (O_1109,N_23531,N_19080);
nand UO_1110 (O_1110,N_20985,N_22163);
xor UO_1111 (O_1111,N_20298,N_19355);
or UO_1112 (O_1112,N_24008,N_20782);
nand UO_1113 (O_1113,N_19875,N_20731);
xor UO_1114 (O_1114,N_23633,N_24844);
and UO_1115 (O_1115,N_19481,N_23816);
and UO_1116 (O_1116,N_22516,N_19605);
nor UO_1117 (O_1117,N_20374,N_19270);
nor UO_1118 (O_1118,N_22525,N_24190);
nand UO_1119 (O_1119,N_20635,N_24118);
nand UO_1120 (O_1120,N_24407,N_19165);
xnor UO_1121 (O_1121,N_23190,N_23353);
nor UO_1122 (O_1122,N_20921,N_18993);
nor UO_1123 (O_1123,N_22289,N_24968);
nand UO_1124 (O_1124,N_21425,N_24277);
or UO_1125 (O_1125,N_21669,N_23996);
and UO_1126 (O_1126,N_22150,N_24737);
or UO_1127 (O_1127,N_22137,N_20386);
nor UO_1128 (O_1128,N_24641,N_23249);
xor UO_1129 (O_1129,N_22454,N_20873);
nor UO_1130 (O_1130,N_21162,N_20334);
or UO_1131 (O_1131,N_20160,N_21578);
nor UO_1132 (O_1132,N_20988,N_23662);
nor UO_1133 (O_1133,N_21781,N_19291);
nor UO_1134 (O_1134,N_21550,N_19236);
or UO_1135 (O_1135,N_20839,N_22919);
and UO_1136 (O_1136,N_21237,N_19912);
and UO_1137 (O_1137,N_24475,N_21977);
nor UO_1138 (O_1138,N_21700,N_20481);
xnor UO_1139 (O_1139,N_22978,N_19137);
nor UO_1140 (O_1140,N_24862,N_22751);
nor UO_1141 (O_1141,N_20528,N_24434);
xnor UO_1142 (O_1142,N_23089,N_23675);
or UO_1143 (O_1143,N_24781,N_20189);
and UO_1144 (O_1144,N_21576,N_24114);
or UO_1145 (O_1145,N_19732,N_20590);
nand UO_1146 (O_1146,N_21616,N_22115);
and UO_1147 (O_1147,N_22646,N_20195);
nor UO_1148 (O_1148,N_20720,N_23637);
and UO_1149 (O_1149,N_22416,N_20938);
and UO_1150 (O_1150,N_20172,N_19588);
xor UO_1151 (O_1151,N_23468,N_24098);
or UO_1152 (O_1152,N_24972,N_20857);
or UO_1153 (O_1153,N_24202,N_21776);
or UO_1154 (O_1154,N_20982,N_20934);
nor UO_1155 (O_1155,N_23041,N_22840);
nor UO_1156 (O_1156,N_19551,N_24183);
xor UO_1157 (O_1157,N_24744,N_22097);
and UO_1158 (O_1158,N_22627,N_20763);
and UO_1159 (O_1159,N_18760,N_19111);
and UO_1160 (O_1160,N_20209,N_24311);
nor UO_1161 (O_1161,N_24631,N_23863);
nand UO_1162 (O_1162,N_22342,N_19867);
nor UO_1163 (O_1163,N_22691,N_21334);
nor UO_1164 (O_1164,N_23371,N_20940);
xor UO_1165 (O_1165,N_24799,N_23238);
nor UO_1166 (O_1166,N_23776,N_21377);
and UO_1167 (O_1167,N_22999,N_20893);
nor UO_1168 (O_1168,N_21342,N_20959);
or UO_1169 (O_1169,N_21339,N_22418);
and UO_1170 (O_1170,N_21256,N_22786);
xor UO_1171 (O_1171,N_19984,N_20705);
nand UO_1172 (O_1172,N_24419,N_19829);
or UO_1173 (O_1173,N_20020,N_21324);
xnor UO_1174 (O_1174,N_23926,N_19943);
and UO_1175 (O_1175,N_23764,N_23748);
or UO_1176 (O_1176,N_19579,N_23212);
nand UO_1177 (O_1177,N_21391,N_20243);
xnor UO_1178 (O_1178,N_22028,N_21485);
nor UO_1179 (O_1179,N_20083,N_23136);
or UO_1180 (O_1180,N_20675,N_22576);
nor UO_1181 (O_1181,N_24330,N_24253);
nand UO_1182 (O_1182,N_19782,N_21501);
xnor UO_1183 (O_1183,N_23189,N_20319);
and UO_1184 (O_1184,N_19813,N_19646);
or UO_1185 (O_1185,N_20295,N_23986);
xnor UO_1186 (O_1186,N_21042,N_21418);
xor UO_1187 (O_1187,N_20441,N_20894);
xor UO_1188 (O_1188,N_20380,N_20587);
xnor UO_1189 (O_1189,N_23737,N_20224);
or UO_1190 (O_1190,N_19414,N_20496);
xor UO_1191 (O_1191,N_24655,N_19509);
or UO_1192 (O_1192,N_20471,N_19353);
or UO_1193 (O_1193,N_23053,N_22159);
xnor UO_1194 (O_1194,N_21702,N_18953);
xnor UO_1195 (O_1195,N_19438,N_23311);
and UO_1196 (O_1196,N_24513,N_19395);
and UO_1197 (O_1197,N_24507,N_24903);
nand UO_1198 (O_1198,N_24568,N_19423);
xnor UO_1199 (O_1199,N_21846,N_22238);
or UO_1200 (O_1200,N_23587,N_24110);
nand UO_1201 (O_1201,N_23199,N_23696);
xnor UO_1202 (O_1202,N_21947,N_22397);
nand UO_1203 (O_1203,N_22665,N_23909);
xor UO_1204 (O_1204,N_18948,N_24966);
xnor UO_1205 (O_1205,N_20761,N_24477);
nor UO_1206 (O_1206,N_21589,N_20499);
xnor UO_1207 (O_1207,N_20758,N_23495);
nor UO_1208 (O_1208,N_22206,N_20424);
nand UO_1209 (O_1209,N_19200,N_24584);
or UO_1210 (O_1210,N_18967,N_21839);
or UO_1211 (O_1211,N_20970,N_19220);
and UO_1212 (O_1212,N_23509,N_21560);
xnor UO_1213 (O_1213,N_22440,N_19168);
or UO_1214 (O_1214,N_23507,N_24397);
or UO_1215 (O_1215,N_19877,N_23305);
nor UO_1216 (O_1216,N_21900,N_24569);
and UO_1217 (O_1217,N_19606,N_20947);
nor UO_1218 (O_1218,N_23307,N_24415);
xnor UO_1219 (O_1219,N_20798,N_18789);
nand UO_1220 (O_1220,N_21532,N_19067);
or UO_1221 (O_1221,N_18882,N_20694);
and UO_1222 (O_1222,N_23008,N_23160);
nor UO_1223 (O_1223,N_20446,N_22994);
nand UO_1224 (O_1224,N_23116,N_22470);
nor UO_1225 (O_1225,N_20133,N_18928);
xnor UO_1226 (O_1226,N_24747,N_22230);
nand UO_1227 (O_1227,N_21415,N_22200);
nor UO_1228 (O_1228,N_22756,N_20869);
xor UO_1229 (O_1229,N_21660,N_21288);
and UO_1230 (O_1230,N_21373,N_20156);
xor UO_1231 (O_1231,N_20747,N_18832);
nand UO_1232 (O_1232,N_19451,N_20382);
nand UO_1233 (O_1233,N_21796,N_20070);
and UO_1234 (O_1234,N_21082,N_20485);
xnor UO_1235 (O_1235,N_23978,N_20950);
nor UO_1236 (O_1236,N_22445,N_24263);
and UO_1237 (O_1237,N_22092,N_21137);
nand UO_1238 (O_1238,N_23530,N_24921);
xor UO_1239 (O_1239,N_22798,N_23283);
and UO_1240 (O_1240,N_22827,N_22563);
or UO_1241 (O_1241,N_23605,N_23677);
nand UO_1242 (O_1242,N_20912,N_21679);
or UO_1243 (O_1243,N_23973,N_22673);
nor UO_1244 (O_1244,N_22204,N_18954);
or UO_1245 (O_1245,N_19260,N_21870);
nand UO_1246 (O_1246,N_22496,N_20245);
and UO_1247 (O_1247,N_19694,N_23988);
nand UO_1248 (O_1248,N_20041,N_22004);
or UO_1249 (O_1249,N_22078,N_23334);
and UO_1250 (O_1250,N_21971,N_24150);
nor UO_1251 (O_1251,N_20681,N_24527);
nor UO_1252 (O_1252,N_24091,N_20246);
xor UO_1253 (O_1253,N_20238,N_22157);
nor UO_1254 (O_1254,N_24132,N_23421);
or UO_1255 (O_1255,N_22429,N_22788);
nor UO_1256 (O_1256,N_19317,N_22703);
nor UO_1257 (O_1257,N_21539,N_24174);
xor UO_1258 (O_1258,N_22977,N_24306);
nor UO_1259 (O_1259,N_19801,N_19604);
or UO_1260 (O_1260,N_20400,N_20249);
and UO_1261 (O_1261,N_19203,N_19436);
xnor UO_1262 (O_1262,N_20623,N_21765);
nand UO_1263 (O_1263,N_20769,N_20352);
or UO_1264 (O_1264,N_19979,N_19616);
xnor UO_1265 (O_1265,N_24911,N_24916);
nor UO_1266 (O_1266,N_19160,N_24188);
or UO_1267 (O_1267,N_20713,N_21721);
or UO_1268 (O_1268,N_19713,N_24380);
nor UO_1269 (O_1269,N_19861,N_22676);
nor UO_1270 (O_1270,N_22715,N_18784);
and UO_1271 (O_1271,N_23360,N_22148);
nand UO_1272 (O_1272,N_20575,N_23009);
and UO_1273 (O_1273,N_21648,N_19570);
or UO_1274 (O_1274,N_21412,N_24885);
and UO_1275 (O_1275,N_22893,N_24695);
xnor UO_1276 (O_1276,N_24592,N_24137);
xor UO_1277 (O_1277,N_24255,N_20585);
nand UO_1278 (O_1278,N_19807,N_20283);
and UO_1279 (O_1279,N_20658,N_23012);
nor UO_1280 (O_1280,N_22596,N_23045);
nor UO_1281 (O_1281,N_20332,N_20315);
nor UO_1282 (O_1282,N_23492,N_22067);
nor UO_1283 (O_1283,N_19352,N_21470);
nand UO_1284 (O_1284,N_20393,N_19576);
and UO_1285 (O_1285,N_20292,N_22982);
or UO_1286 (O_1286,N_24134,N_24679);
nand UO_1287 (O_1287,N_20878,N_21789);
xnor UO_1288 (O_1288,N_19427,N_20855);
xor UO_1289 (O_1289,N_21879,N_18999);
nand UO_1290 (O_1290,N_23886,N_21973);
and UO_1291 (O_1291,N_19585,N_19703);
and UO_1292 (O_1292,N_24488,N_21101);
and UO_1293 (O_1293,N_19363,N_20935);
or UO_1294 (O_1294,N_18978,N_22335);
xnor UO_1295 (O_1295,N_24377,N_23267);
nor UO_1296 (O_1296,N_24320,N_21198);
nor UO_1297 (O_1297,N_23011,N_19676);
xnor UO_1298 (O_1298,N_21398,N_22109);
nor UO_1299 (O_1299,N_21848,N_21498);
and UO_1300 (O_1300,N_19464,N_22471);
and UO_1301 (O_1301,N_18856,N_23016);
xnor UO_1302 (O_1302,N_24125,N_23475);
nand UO_1303 (O_1303,N_19328,N_19573);
and UO_1304 (O_1304,N_21438,N_24080);
nor UO_1305 (O_1305,N_20309,N_23181);
nor UO_1306 (O_1306,N_24334,N_21268);
nand UO_1307 (O_1307,N_23323,N_21176);
nand UO_1308 (O_1308,N_24812,N_19500);
nand UO_1309 (O_1309,N_19970,N_24620);
nor UO_1310 (O_1310,N_24454,N_20860);
nor UO_1311 (O_1311,N_22710,N_22107);
or UO_1312 (O_1312,N_20001,N_24245);
nand UO_1313 (O_1313,N_24238,N_19283);
xnor UO_1314 (O_1314,N_20257,N_18869);
nor UO_1315 (O_1315,N_20530,N_22983);
nand UO_1316 (O_1316,N_23299,N_24168);
xor UO_1317 (O_1317,N_22486,N_23088);
xor UO_1318 (O_1318,N_19045,N_23180);
and UO_1319 (O_1319,N_22410,N_21511);
and UO_1320 (O_1320,N_20391,N_21289);
nor UO_1321 (O_1321,N_23202,N_23770);
nand UO_1322 (O_1322,N_23721,N_19910);
and UO_1323 (O_1323,N_21099,N_23402);
xnor UO_1324 (O_1324,N_23704,N_23479);
nand UO_1325 (O_1325,N_23341,N_18941);
nand UO_1326 (O_1326,N_21316,N_24216);
nor UO_1327 (O_1327,N_19529,N_19187);
or UO_1328 (O_1328,N_24609,N_19391);
nor UO_1329 (O_1329,N_20121,N_24483);
or UO_1330 (O_1330,N_22912,N_20436);
or UO_1331 (O_1331,N_22692,N_21916);
and UO_1332 (O_1332,N_24981,N_21228);
nor UO_1333 (O_1333,N_22145,N_24766);
xor UO_1334 (O_1334,N_23172,N_21168);
nand UO_1335 (O_1335,N_21849,N_24455);
or UO_1336 (O_1336,N_22518,N_19396);
nand UO_1337 (O_1337,N_24616,N_24662);
or UO_1338 (O_1338,N_20861,N_20390);
and UO_1339 (O_1339,N_18801,N_21516);
or UO_1340 (O_1340,N_23745,N_21141);
nand UO_1341 (O_1341,N_20555,N_21966);
nor UO_1342 (O_1342,N_19567,N_22014);
xnor UO_1343 (O_1343,N_20194,N_19935);
and UO_1344 (O_1344,N_24974,N_23722);
nand UO_1345 (O_1345,N_19484,N_22797);
or UO_1346 (O_1346,N_19219,N_22356);
xor UO_1347 (O_1347,N_19852,N_22989);
nand UO_1348 (O_1348,N_19817,N_21008);
xor UO_1349 (O_1349,N_19077,N_21691);
or UO_1350 (O_1350,N_19981,N_20305);
xnor UO_1351 (O_1351,N_24855,N_21641);
or UO_1352 (O_1352,N_21682,N_22186);
nor UO_1353 (O_1353,N_21064,N_23022);
or UO_1354 (O_1354,N_20050,N_19878);
and UO_1355 (O_1355,N_23129,N_23582);
xor UO_1356 (O_1356,N_23705,N_23649);
and UO_1357 (O_1357,N_19050,N_23670);
nor UO_1358 (O_1358,N_24689,N_21169);
and UO_1359 (O_1359,N_19897,N_20356);
and UO_1360 (O_1360,N_24267,N_23802);
nor UO_1361 (O_1361,N_20063,N_19645);
xor UO_1362 (O_1362,N_22446,N_23483);
nand UO_1363 (O_1363,N_24730,N_21360);
nor UO_1364 (O_1364,N_21219,N_24009);
or UO_1365 (O_1365,N_20558,N_21952);
and UO_1366 (O_1366,N_20859,N_20339);
nor UO_1367 (O_1367,N_20051,N_22358);
nand UO_1368 (O_1368,N_21703,N_19388);
or UO_1369 (O_1369,N_24155,N_22152);
xnor UO_1370 (O_1370,N_20344,N_19827);
nand UO_1371 (O_1371,N_21427,N_20524);
nor UO_1372 (O_1372,N_23465,N_18803);
nor UO_1373 (O_1373,N_21970,N_22819);
and UO_1374 (O_1374,N_22675,N_19367);
nor UO_1375 (O_1375,N_23876,N_23636);
nand UO_1376 (O_1376,N_24038,N_21078);
or UO_1377 (O_1377,N_18904,N_23527);
or UO_1378 (O_1378,N_20849,N_22212);
nor UO_1379 (O_1379,N_24659,N_23583);
xor UO_1380 (O_1380,N_22114,N_24767);
nor UO_1381 (O_1381,N_21267,N_23821);
or UO_1382 (O_1382,N_22174,N_19003);
or UO_1383 (O_1383,N_21819,N_19653);
nand UO_1384 (O_1384,N_22727,N_22853);
nor UO_1385 (O_1385,N_24839,N_23689);
and UO_1386 (O_1386,N_22231,N_19415);
nand UO_1387 (O_1387,N_19014,N_23664);
nor UO_1388 (O_1388,N_24244,N_21884);
nand UO_1389 (O_1389,N_20752,N_23110);
or UO_1390 (O_1390,N_22937,N_19609);
nand UO_1391 (O_1391,N_19366,N_23059);
nand UO_1392 (O_1392,N_23120,N_24880);
xor UO_1393 (O_1393,N_21188,N_19831);
or UO_1394 (O_1394,N_22528,N_19712);
and UO_1395 (O_1395,N_23256,N_23065);
nor UO_1396 (O_1396,N_23472,N_18775);
nor UO_1397 (O_1397,N_22863,N_20200);
and UO_1398 (O_1398,N_23500,N_19275);
xnor UO_1399 (O_1399,N_18917,N_24390);
xor UO_1400 (O_1400,N_19446,N_20092);
and UO_1401 (O_1401,N_24579,N_24445);
nand UO_1402 (O_1402,N_19542,N_21591);
nand UO_1403 (O_1403,N_21943,N_19552);
nor UO_1404 (O_1404,N_19401,N_23660);
and UO_1405 (O_1405,N_21320,N_23207);
and UO_1406 (O_1406,N_19555,N_22579);
xor UO_1407 (O_1407,N_20198,N_20145);
or UO_1408 (O_1408,N_22716,N_23164);
or UO_1409 (O_1409,N_19754,N_19132);
or UO_1410 (O_1410,N_21277,N_19651);
or UO_1411 (O_1411,N_23270,N_19204);
and UO_1412 (O_1412,N_22270,N_22431);
xor UO_1413 (O_1413,N_21732,N_22717);
or UO_1414 (O_1414,N_22888,N_20445);
nor UO_1415 (O_1415,N_23326,N_18958);
nor UO_1416 (O_1416,N_23998,N_22297);
nand UO_1417 (O_1417,N_21476,N_19254);
and UO_1418 (O_1418,N_20518,N_24779);
and UO_1419 (O_1419,N_22379,N_20123);
and UO_1420 (O_1420,N_24896,N_18918);
and UO_1421 (O_1421,N_20262,N_19654);
or UO_1422 (O_1422,N_23560,N_23023);
and UO_1423 (O_1423,N_19320,N_20320);
nand UO_1424 (O_1424,N_23729,N_19437);
nor UO_1425 (O_1425,N_23419,N_22802);
or UO_1426 (O_1426,N_24147,N_20987);
nor UO_1427 (O_1427,N_19976,N_20814);
nand UO_1428 (O_1428,N_19541,N_23667);
xor UO_1429 (O_1429,N_24516,N_20672);
xor UO_1430 (O_1430,N_23048,N_19372);
xor UO_1431 (O_1431,N_18893,N_21343);
nor UO_1432 (O_1432,N_22334,N_23880);
or UO_1433 (O_1433,N_24081,N_24436);
xor UO_1434 (O_1434,N_19339,N_24667);
nand UO_1435 (O_1435,N_23060,N_21969);
nor UO_1436 (O_1436,N_23405,N_23843);
nor UO_1437 (O_1437,N_19264,N_24228);
nand UO_1438 (O_1438,N_24938,N_22317);
nand UO_1439 (O_1439,N_22784,N_24934);
xnor UO_1440 (O_1440,N_22630,N_22171);
nand UO_1441 (O_1441,N_22754,N_22274);
xor UO_1442 (O_1442,N_20163,N_21854);
and UO_1443 (O_1443,N_19928,N_22352);
and UO_1444 (O_1444,N_20168,N_20801);
nand UO_1445 (O_1445,N_22491,N_23108);
or UO_1446 (O_1446,N_21928,N_23659);
and UO_1447 (O_1447,N_21655,N_22781);
and UO_1448 (O_1448,N_21637,N_20866);
xnor UO_1449 (O_1449,N_21902,N_19330);
nor UO_1450 (O_1450,N_23489,N_24095);
nor UO_1451 (O_1451,N_19738,N_19060);
or UO_1452 (O_1452,N_24167,N_23954);
or UO_1453 (O_1453,N_23594,N_21368);
and UO_1454 (O_1454,N_20389,N_24157);
nand UO_1455 (O_1455,N_19340,N_19765);
nor UO_1456 (O_1456,N_23026,N_24422);
nor UO_1457 (O_1457,N_23735,N_21997);
nor UO_1458 (O_1458,N_23682,N_23958);
nor UO_1459 (O_1459,N_19068,N_20028);
xnor UO_1460 (O_1460,N_23751,N_21698);
nor UO_1461 (O_1461,N_23518,N_20071);
xnor UO_1462 (O_1462,N_23975,N_24037);
nand UO_1463 (O_1463,N_22771,N_23906);
nand UO_1464 (O_1464,N_20942,N_21154);
xnor UO_1465 (O_1465,N_24600,N_19955);
nand UO_1466 (O_1466,N_22428,N_19382);
nor UO_1467 (O_1467,N_19566,N_21805);
xnor UO_1468 (O_1468,N_23837,N_19394);
and UO_1469 (O_1469,N_20162,N_19824);
nor UO_1470 (O_1470,N_21353,N_22165);
nand UO_1471 (O_1471,N_19995,N_20683);
nor UO_1472 (O_1472,N_24770,N_19997);
and UO_1473 (O_1473,N_19806,N_22483);
nand UO_1474 (O_1474,N_22404,N_19916);
and UO_1475 (O_1475,N_22399,N_24067);
xor UO_1476 (O_1476,N_20975,N_19351);
nor UO_1477 (O_1477,N_23414,N_20438);
nand UO_1478 (O_1478,N_22661,N_24381);
and UO_1479 (O_1479,N_20858,N_22314);
and UO_1480 (O_1480,N_21306,N_22258);
nand UO_1481 (O_1481,N_19207,N_19569);
or UO_1482 (O_1482,N_23545,N_22139);
or UO_1483 (O_1483,N_20577,N_24832);
xor UO_1484 (O_1484,N_21376,N_19865);
xor UO_1485 (O_1485,N_18884,N_22236);
nor UO_1486 (O_1486,N_21121,N_23343);
or UO_1487 (O_1487,N_24261,N_20288);
nand UO_1488 (O_1488,N_23798,N_20547);
nand UO_1489 (O_1489,N_18966,N_22931);
nor UO_1490 (O_1490,N_21191,N_22591);
xor UO_1491 (O_1491,N_18823,N_19902);
and UO_1492 (O_1492,N_19109,N_23586);
nand UO_1493 (O_1493,N_20790,N_20566);
nand UO_1494 (O_1494,N_20927,N_20824);
xor UO_1495 (O_1495,N_24159,N_21202);
nor UO_1496 (O_1496,N_21690,N_20564);
and UO_1497 (O_1497,N_18871,N_20777);
and UO_1498 (O_1498,N_19740,N_22620);
xor UO_1499 (O_1499,N_22808,N_22248);
nor UO_1500 (O_1500,N_19192,N_19755);
nand UO_1501 (O_1501,N_24710,N_19814);
xor UO_1502 (O_1502,N_19324,N_22426);
or UO_1503 (O_1503,N_21527,N_21659);
or UO_1504 (O_1504,N_24987,N_22504);
nand UO_1505 (O_1505,N_20733,N_24801);
nor UO_1506 (O_1506,N_18903,N_22668);
and UO_1507 (O_1507,N_21348,N_24652);
or UO_1508 (O_1508,N_22188,N_22814);
or UO_1509 (O_1509,N_20475,N_19665);
nor UO_1510 (O_1510,N_18894,N_19323);
xor UO_1511 (O_1511,N_19898,N_19907);
xor UO_1512 (O_1512,N_24421,N_23604);
nand UO_1513 (O_1513,N_23697,N_19184);
and UO_1514 (O_1514,N_22618,N_21400);
or UO_1515 (O_1515,N_23820,N_23634);
nor UO_1516 (O_1516,N_19595,N_23210);
nor UO_1517 (O_1517,N_20000,N_23918);
and UO_1518 (O_1518,N_21956,N_24055);
or UO_1519 (O_1519,N_23872,N_18887);
or UO_1520 (O_1520,N_22272,N_22432);
or UO_1521 (O_1521,N_19511,N_23684);
or UO_1522 (O_1522,N_24774,N_19098);
or UO_1523 (O_1523,N_22617,N_18822);
xnor UO_1524 (O_1524,N_20416,N_20058);
or UO_1525 (O_1525,N_24634,N_23597);
and UO_1526 (O_1526,N_19061,N_20254);
xor UO_1527 (O_1527,N_24556,N_22060);
or UO_1528 (O_1528,N_22154,N_24504);
xnor UO_1529 (O_1529,N_23724,N_22481);
and UO_1530 (O_1530,N_22339,N_22453);
and UO_1531 (O_1531,N_21147,N_19951);
and UO_1532 (O_1532,N_23044,N_23470);
nand UO_1533 (O_1533,N_23643,N_19018);
and UO_1534 (O_1534,N_20638,N_19113);
or UO_1535 (O_1535,N_20759,N_19930);
and UO_1536 (O_1536,N_19701,N_20767);
and UO_1537 (O_1537,N_19234,N_18750);
and UO_1538 (O_1538,N_20972,N_19937);
or UO_1539 (O_1539,N_24729,N_19371);
nor UO_1540 (O_1540,N_21297,N_24119);
xor UO_1541 (O_1541,N_23964,N_20562);
or UO_1542 (O_1542,N_21419,N_21663);
xor UO_1543 (O_1543,N_24750,N_22263);
or UO_1544 (O_1544,N_21203,N_23542);
nor UO_1545 (O_1545,N_22249,N_22149);
and UO_1546 (O_1546,N_24104,N_23443);
or UO_1547 (O_1547,N_19718,N_24078);
or UO_1548 (O_1548,N_24340,N_19996);
nand UO_1549 (O_1549,N_20594,N_23857);
and UO_1550 (O_1550,N_22555,N_22283);
nor UO_1551 (O_1551,N_19272,N_20278);
and UO_1552 (O_1552,N_20828,N_20077);
nand UO_1553 (O_1553,N_20306,N_23367);
xor UO_1554 (O_1554,N_23913,N_20716);
xor UO_1555 (O_1555,N_21302,N_23904);
xnor UO_1556 (O_1556,N_19864,N_23707);
and UO_1557 (O_1557,N_22554,N_24413);
and UO_1558 (O_1558,N_23138,N_23602);
and UO_1559 (O_1559,N_23192,N_22088);
nand UO_1560 (O_1560,N_20299,N_21737);
nand UO_1561 (O_1561,N_20302,N_24251);
nand UO_1562 (O_1562,N_20653,N_24649);
xor UO_1563 (O_1563,N_20601,N_24160);
or UO_1564 (O_1564,N_19089,N_24336);
nor UO_1565 (O_1565,N_24427,N_23459);
xor UO_1566 (O_1566,N_22547,N_23723);
nand UO_1567 (O_1567,N_23786,N_22193);
nand UO_1568 (O_1568,N_19329,N_20078);
nor UO_1569 (O_1569,N_20852,N_20164);
nand UO_1570 (O_1570,N_19338,N_22305);
nor UO_1571 (O_1571,N_22218,N_23375);
nand UO_1572 (O_1572,N_19290,N_21222);
nand UO_1573 (O_1573,N_18957,N_23713);
nand UO_1574 (O_1574,N_23376,N_21010);
and UO_1575 (O_1575,N_20529,N_21486);
nor UO_1576 (O_1576,N_21451,N_20887);
nand UO_1577 (O_1577,N_23084,N_19779);
or UO_1578 (O_1578,N_20557,N_21894);
or UO_1579 (O_1579,N_23727,N_21891);
xor UO_1580 (O_1580,N_24682,N_19373);
xor UO_1581 (O_1581,N_21122,N_22517);
or UO_1582 (O_1582,N_22031,N_24715);
nor UO_1583 (O_1583,N_22083,N_19190);
nand UO_1584 (O_1584,N_24481,N_22975);
and UO_1585 (O_1585,N_24087,N_18981);
nor UO_1586 (O_1586,N_22257,N_23563);
nand UO_1587 (O_1587,N_20396,N_24399);
nor UO_1588 (O_1588,N_23075,N_20999);
nand UO_1589 (O_1589,N_24845,N_20837);
xnor UO_1590 (O_1590,N_20719,N_20468);
nand UO_1591 (O_1591,N_22909,N_21325);
xor UO_1592 (O_1592,N_23694,N_24558);
nor UO_1593 (O_1593,N_23404,N_24909);
or UO_1594 (O_1594,N_20634,N_20884);
or UO_1595 (O_1595,N_19281,N_24439);
or UO_1596 (O_1596,N_21800,N_21565);
nand UO_1597 (O_1597,N_19039,N_24577);
or UO_1598 (O_1598,N_20091,N_20433);
or UO_1599 (O_1599,N_19224,N_21174);
nand UO_1600 (O_1600,N_24549,N_20586);
nand UO_1601 (O_1601,N_22221,N_21155);
nand UO_1602 (O_1602,N_22074,N_18879);
nor UO_1603 (O_1603,N_21546,N_24288);
or UO_1604 (O_1604,N_23261,N_24156);
or UO_1605 (O_1605,N_20841,N_22640);
nand UO_1606 (O_1606,N_20803,N_20932);
and UO_1607 (O_1607,N_23773,N_20610);
nor UO_1608 (O_1608,N_21688,N_20872);
and UO_1609 (O_1609,N_20061,N_24926);
and UO_1610 (O_1610,N_21976,N_19286);
or UO_1611 (O_1611,N_24470,N_23124);
or UO_1612 (O_1612,N_22243,N_24941);
xnor UO_1613 (O_1613,N_22895,N_22321);
and UO_1614 (O_1614,N_24557,N_22613);
nor UO_1615 (O_1615,N_22878,N_18891);
and UO_1616 (O_1616,N_20108,N_19751);
nand UO_1617 (O_1617,N_20736,N_23215);
or UO_1618 (O_1618,N_19142,N_22908);
or UO_1619 (O_1619,N_22642,N_21424);
and UO_1620 (O_1620,N_23295,N_23815);
nand UO_1621 (O_1621,N_24333,N_20178);
xor UO_1622 (O_1622,N_21843,N_21759);
or UO_1623 (O_1623,N_24031,N_21017);
nor UO_1624 (O_1624,N_24218,N_22034);
and UO_1625 (O_1625,N_23924,N_23849);
nand UO_1626 (O_1626,N_24176,N_22749);
nor UO_1627 (O_1627,N_19343,N_21677);
xor UO_1628 (O_1628,N_22981,N_20351);
xor UO_1629 (O_1629,N_22940,N_24003);
nand UO_1630 (O_1630,N_21074,N_23514);
nor UO_1631 (O_1631,N_22363,N_21142);
nand UO_1632 (O_1632,N_20362,N_22288);
nand UO_1633 (O_1633,N_22081,N_19435);
and UO_1634 (O_1634,N_21347,N_19114);
and UO_1635 (O_1635,N_23791,N_19152);
or UO_1636 (O_1636,N_22616,N_21623);
nand UO_1637 (O_1637,N_21763,N_19571);
nor UO_1638 (O_1638,N_21937,N_19479);
nor UO_1639 (O_1639,N_20015,N_22809);
or UO_1640 (O_1640,N_22729,N_18781);
nand UO_1641 (O_1641,N_18916,N_19702);
nor UO_1642 (O_1642,N_20214,N_24993);
xor UO_1643 (O_1643,N_21285,N_24597);
nor UO_1644 (O_1644,N_19209,N_24883);
and UO_1645 (O_1645,N_24133,N_23700);
or UO_1646 (O_1646,N_24990,N_18799);
or UO_1647 (O_1647,N_19625,N_20316);
xor UO_1648 (O_1648,N_23851,N_19637);
xnor UO_1649 (O_1649,N_22946,N_19282);
nand UO_1650 (O_1650,N_23167,N_21664);
or UO_1651 (O_1651,N_23417,N_21378);
and UO_1652 (O_1652,N_22678,N_20484);
or UO_1653 (O_1653,N_20267,N_21901);
and UO_1654 (O_1654,N_19800,N_21313);
nand UO_1655 (O_1655,N_22973,N_23259);
xnor UO_1656 (O_1656,N_22829,N_22395);
and UO_1657 (O_1657,N_20089,N_22412);
nor UO_1658 (O_1658,N_24048,N_24857);
or UO_1659 (O_1659,N_19397,N_24726);
nor UO_1660 (O_1660,N_22328,N_23042);
nor UO_1661 (O_1661,N_22785,N_22695);
nor UO_1662 (O_1662,N_21383,N_23265);
and UO_1663 (O_1663,N_24469,N_22633);
xnor UO_1664 (O_1664,N_22168,N_21905);
and UO_1665 (O_1665,N_21644,N_22838);
nor UO_1666 (O_1666,N_18780,N_19982);
or UO_1667 (O_1667,N_22552,N_24461);
and UO_1668 (O_1668,N_22169,N_20816);
nor UO_1669 (O_1669,N_21336,N_22558);
or UO_1670 (O_1670,N_21437,N_22652);
nand UO_1671 (O_1671,N_20980,N_23761);
nand UO_1672 (O_1672,N_21403,N_20657);
nor UO_1673 (O_1673,N_23532,N_23834);
nor UO_1674 (O_1674,N_23364,N_19931);
and UO_1675 (O_1675,N_22195,N_20289);
xnor UO_1676 (O_1676,N_21636,N_18850);
or UO_1677 (O_1677,N_23039,N_22434);
nand UO_1678 (O_1678,N_19961,N_24551);
xnor UO_1679 (O_1679,N_23887,N_22667);
or UO_1680 (O_1680,N_20147,N_23510);
xnor UO_1681 (O_1681,N_22686,N_21489);
and UO_1682 (O_1682,N_20431,N_24438);
nor UO_1683 (O_1683,N_21109,N_21657);
and UO_1684 (O_1684,N_22036,N_21070);
or UO_1685 (O_1685,N_23625,N_22053);
xnor UO_1686 (O_1686,N_19924,N_21217);
and UO_1687 (O_1687,N_21788,N_20341);
nor UO_1688 (O_1688,N_23806,N_19695);
and UO_1689 (O_1689,N_23824,N_18965);
nor UO_1690 (O_1690,N_18854,N_21417);
nand UO_1691 (O_1691,N_22502,N_23151);
or UO_1692 (O_1692,N_18920,N_24920);
and UO_1693 (O_1693,N_23070,N_22825);
nor UO_1694 (O_1694,N_23832,N_23146);
nand UO_1695 (O_1695,N_23801,N_22375);
nor UO_1696 (O_1696,N_24416,N_22118);
xor UO_1697 (O_1697,N_23166,N_21959);
nor UO_1698 (O_1698,N_21764,N_22353);
nand UO_1699 (O_1699,N_21967,N_23132);
nor UO_1700 (O_1700,N_22935,N_23028);
or UO_1701 (O_1701,N_19596,N_20345);
nor UO_1702 (O_1702,N_19874,N_24100);
nand UO_1703 (O_1703,N_21684,N_22831);
xnor UO_1704 (O_1704,N_20211,N_20702);
nor UO_1705 (O_1705,N_20892,N_22531);
nor UO_1706 (O_1706,N_19917,N_19673);
and UO_1707 (O_1707,N_21123,N_24819);
and UO_1708 (O_1708,N_22054,N_24773);
xnor UO_1709 (O_1709,N_22541,N_22122);
or UO_1710 (O_1710,N_23741,N_19722);
nor UO_1711 (O_1711,N_19121,N_19548);
xor UO_1712 (O_1712,N_21869,N_22110);
nand UO_1713 (O_1713,N_23498,N_21367);
nand UO_1714 (O_1714,N_23712,N_21263);
xor UO_1715 (O_1715,N_19636,N_19357);
nor UO_1716 (O_1716,N_20991,N_23057);
or UO_1717 (O_1717,N_19603,N_23264);
nor UO_1718 (O_1718,N_22864,N_23177);
nand UO_1719 (O_1719,N_20363,N_22514);
and UO_1720 (O_1720,N_23387,N_22304);
nor UO_1721 (O_1721,N_22347,N_19842);
nand UO_1722 (O_1722,N_20611,N_19873);
nand UO_1723 (O_1723,N_19999,N_19428);
or UO_1724 (O_1724,N_23463,N_22607);
xor UO_1725 (O_1725,N_21980,N_19737);
and UO_1726 (O_1726,N_19967,N_19154);
nand UO_1727 (O_1727,N_20734,N_23902);
nor UO_1728 (O_1728,N_19649,N_19301);
nor UO_1729 (O_1729,N_20307,N_21102);
or UO_1730 (O_1730,N_24351,N_23306);
nor UO_1731 (O_1731,N_20833,N_20343);
nand UO_1732 (O_1732,N_24375,N_20169);
nor UO_1733 (O_1733,N_24058,N_23216);
nand UO_1734 (O_1734,N_19945,N_21674);
or UO_1735 (O_1735,N_20190,N_24958);
nor UO_1736 (O_1736,N_20137,N_21856);
nand UO_1737 (O_1737,N_20708,N_23841);
nor UO_1738 (O_1738,N_23237,N_20282);
nand UO_1739 (O_1739,N_21248,N_21146);
nor UO_1740 (O_1740,N_18794,N_20968);
xor UO_1741 (O_1741,N_22987,N_20410);
nand UO_1742 (O_1742,N_20900,N_18897);
nand UO_1743 (O_1743,N_21750,N_19227);
nor UO_1744 (O_1744,N_24939,N_20450);
and UO_1745 (O_1745,N_19652,N_21792);
xnor UO_1746 (O_1746,N_19692,N_23144);
and UO_1747 (O_1747,N_24272,N_22178);
xnor UO_1748 (O_1748,N_22582,N_20297);
xor UO_1749 (O_1749,N_23369,N_19006);
nor UO_1750 (O_1750,N_21859,N_21335);
nand UO_1751 (O_1751,N_24624,N_23063);
and UO_1752 (O_1752,N_24448,N_22637);
xnor UO_1753 (O_1753,N_20330,N_21472);
nand UO_1754 (O_1754,N_20140,N_20756);
nor UO_1755 (O_1755,N_22388,N_24895);
nand UO_1756 (O_1756,N_21208,N_24197);
nand UO_1757 (O_1757,N_24429,N_23885);
and UO_1758 (O_1758,N_22689,N_23407);
and UO_1759 (O_1759,N_20104,N_23957);
xor UO_1760 (O_1760,N_19157,N_19255);
nor UO_1761 (O_1761,N_19188,N_22736);
nor UO_1762 (O_1762,N_22677,N_19297);
or UO_1763 (O_1763,N_19687,N_22112);
or UO_1764 (O_1764,N_22941,N_21945);
nand UO_1765 (O_1765,N_19753,N_23330);
and UO_1766 (O_1766,N_23739,N_21784);
nand UO_1767 (O_1767,N_22089,N_19307);
and UO_1768 (O_1768,N_24732,N_19205);
or UO_1769 (O_1769,N_21921,N_20057);
or UO_1770 (O_1770,N_19942,N_23096);
or UO_1771 (O_1771,N_22990,N_24070);
xor UO_1772 (O_1772,N_20017,N_21782);
nand UO_1773 (O_1773,N_24467,N_19919);
xnor UO_1774 (O_1774,N_20588,N_24203);
nand UO_1775 (O_1775,N_22672,N_22984);
or UO_1776 (O_1776,N_23653,N_24835);
xor UO_1777 (O_1777,N_21253,N_24687);
nand UO_1778 (O_1778,N_22180,N_20501);
and UO_1779 (O_1779,N_20910,N_24772);
xnor UO_1780 (O_1780,N_22874,N_23901);
nor UO_1781 (O_1781,N_19044,N_23303);
or UO_1782 (O_1782,N_22748,N_24173);
or UO_1783 (O_1783,N_21841,N_22581);
nand UO_1784 (O_1784,N_23971,N_19904);
or UO_1785 (O_1785,N_20149,N_24041);
or UO_1786 (O_1786,N_22755,N_21314);
or UO_1787 (O_1787,N_23972,N_22942);
xor UO_1788 (O_1788,N_21132,N_19259);
and UO_1789 (O_1789,N_22588,N_21787);
or UO_1790 (O_1790,N_21544,N_20073);
xor UO_1791 (O_1791,N_23642,N_23923);
xnor UO_1792 (O_1792,N_24023,N_24589);
or UO_1793 (O_1793,N_22577,N_18754);
nand UO_1794 (O_1794,N_22116,N_23915);
or UO_1795 (O_1795,N_24784,N_21681);
nand UO_1796 (O_1796,N_24108,N_24004);
and UO_1797 (O_1797,N_19911,N_19475);
nand UO_1798 (O_1798,N_22311,N_19457);
or UO_1799 (O_1799,N_19295,N_19770);
nor UO_1800 (O_1800,N_24838,N_20284);
or UO_1801 (O_1801,N_19820,N_22472);
and UO_1802 (O_1802,N_20310,N_23109);
and UO_1803 (O_1803,N_21294,N_21837);
or UO_1804 (O_1804,N_20700,N_24012);
and UO_1805 (O_1805,N_24143,N_22235);
xor UO_1806 (O_1806,N_22181,N_20820);
nor UO_1807 (O_1807,N_20370,N_24697);
and UO_1808 (O_1808,N_22880,N_19030);
or UO_1809 (O_1809,N_21152,N_24816);
nand UO_1810 (O_1810,N_21104,N_19534);
nor UO_1811 (O_1811,N_19143,N_22002);
nand UO_1812 (O_1812,N_19019,N_20565);
and UO_1813 (O_1813,N_20472,N_19818);
nand UO_1814 (O_1814,N_18842,N_21840);
nor UO_1815 (O_1815,N_24820,N_21375);
nor UO_1816 (O_1816,N_23601,N_21571);
xor UO_1817 (O_1817,N_20394,N_24473);
and UO_1818 (O_1818,N_22176,N_19678);
and UO_1819 (O_1819,N_22600,N_23018);
xnor UO_1820 (O_1820,N_19458,N_20479);
xor UO_1821 (O_1821,N_19841,N_18792);
and UO_1822 (O_1822,N_23244,N_21567);
xnor UO_1823 (O_1823,N_22553,N_23539);
nand UO_1824 (O_1824,N_20909,N_20244);
and UO_1825 (O_1825,N_22834,N_19163);
or UO_1826 (O_1826,N_22529,N_23781);
or UO_1827 (O_1827,N_21592,N_18825);
nor UO_1828 (O_1828,N_22953,N_20413);
or UO_1829 (O_1829,N_23991,N_23503);
xnor UO_1830 (O_1830,N_23121,N_21885);
nor UO_1831 (O_1831,N_22653,N_20090);
nand UO_1832 (O_1832,N_21689,N_21330);
and UO_1833 (O_1833,N_21514,N_20291);
nor UO_1834 (O_1834,N_24673,N_20263);
nor UO_1835 (O_1835,N_23690,N_22027);
and UO_1836 (O_1836,N_21748,N_23128);
xnor UO_1837 (O_1837,N_24022,N_20738);
and UO_1838 (O_1838,N_22920,N_21027);
xnor UO_1839 (O_1839,N_19206,N_18769);
nand UO_1840 (O_1840,N_23907,N_24404);
and UO_1841 (O_1841,N_24234,N_19839);
nand UO_1842 (O_1842,N_19069,N_22513);
nand UO_1843 (O_1843,N_18864,N_19923);
nor UO_1844 (O_1844,N_20604,N_24663);
nor UO_1845 (O_1845,N_21667,N_21148);
nand UO_1846 (O_1846,N_20973,N_22384);
nand UO_1847 (O_1847,N_18753,N_23784);
and UO_1848 (O_1848,N_19347,N_22969);
or UO_1849 (O_1849,N_21604,N_20004);
xor UO_1850 (O_1850,N_23251,N_18961);
nor UO_1851 (O_1851,N_19715,N_24756);
nand UO_1852 (O_1852,N_22735,N_23898);
nand UO_1853 (O_1853,N_23891,N_18952);
or UO_1854 (O_1854,N_18840,N_22252);
and UO_1855 (O_1855,N_24751,N_19053);
and UO_1856 (O_1856,N_22699,N_22338);
or UO_1857 (O_1857,N_18772,N_21816);
xor UO_1858 (O_1858,N_24722,N_19517);
or UO_1859 (O_1859,N_23378,N_20845);
xor UO_1860 (O_1860,N_20412,N_24184);
or UO_1861 (O_1861,N_24025,N_22312);
or UO_1862 (O_1862,N_20167,N_22537);
nor UO_1863 (O_1863,N_23213,N_24072);
xnor UO_1864 (O_1864,N_21044,N_19078);
xor UO_1865 (O_1865,N_24032,N_24007);
and UO_1866 (O_1866,N_19325,N_22883);
nand UO_1867 (O_1867,N_19835,N_20620);
nand UO_1868 (O_1868,N_21758,N_22233);
and UO_1869 (O_1869,N_23927,N_24886);
nor UO_1870 (O_1870,N_24378,N_24423);
and UO_1871 (O_1871,N_21661,N_19404);
and UO_1872 (O_1872,N_23540,N_24960);
nand UO_1873 (O_1873,N_21243,N_19327);
and UO_1874 (O_1874,N_22774,N_23953);
nor UO_1875 (O_1875,N_20159,N_21478);
xnor UO_1876 (O_1876,N_24814,N_20271);
nand UO_1877 (O_1877,N_22768,N_19494);
xnor UO_1878 (O_1878,N_21481,N_22077);
nor UO_1879 (O_1879,N_22972,N_21346);
xnor UO_1880 (O_1880,N_22980,N_20049);
and UO_1881 (O_1881,N_24178,N_20549);
nand UO_1882 (O_1882,N_23005,N_20969);
nor UO_1883 (O_1883,N_23960,N_20786);
and UO_1884 (O_1884,N_19764,N_23681);
and UO_1885 (O_1885,N_21250,N_21564);
or UO_1886 (O_1886,N_21957,N_23441);
xnor UO_1887 (O_1887,N_19516,N_18972);
and UO_1888 (O_1888,N_20177,N_24971);
or UO_1889 (O_1889,N_24304,N_23596);
or UO_1890 (O_1890,N_24711,N_22479);
nor UO_1891 (O_1891,N_20904,N_20633);
or UO_1892 (O_1892,N_19378,N_18814);
and UO_1893 (O_1893,N_21160,N_22614);
xnor UO_1894 (O_1894,N_19134,N_19370);
nand UO_1895 (O_1895,N_24748,N_22355);
or UO_1896 (O_1896,N_23223,N_22117);
and UO_1897 (O_1897,N_19079,N_20383);
or UO_1898 (O_1898,N_21456,N_24269);
or UO_1899 (O_1899,N_23746,N_21389);
or UO_1900 (O_1900,N_19158,N_20784);
nor UO_1901 (O_1901,N_23288,N_24420);
nor UO_1902 (O_1902,N_20888,N_22370);
or UO_1903 (O_1903,N_23543,N_21825);
nor UO_1904 (O_1904,N_23585,N_24769);
nor UO_1905 (O_1905,N_20217,N_24618);
nor UO_1906 (O_1906,N_20661,N_19507);
nor UO_1907 (O_1907,N_18752,N_22222);
and UO_1908 (O_1908,N_24494,N_19526);
or UO_1909 (O_1909,N_22711,N_19508);
nand UO_1910 (O_1910,N_22229,N_18994);
and UO_1911 (O_1911,N_24102,N_21097);
and UO_1912 (O_1912,N_23318,N_24491);
nand UO_1913 (O_1913,N_19443,N_23348);
nor UO_1914 (O_1914,N_19217,N_21370);
or UO_1915 (O_1915,N_22590,N_22023);
or UO_1916 (O_1916,N_22950,N_22211);
xnor UO_1917 (O_1917,N_21206,N_20054);
or UO_1918 (O_1918,N_23840,N_20085);
nand UO_1919 (O_1919,N_21826,N_19287);
xnor UO_1920 (O_1920,N_24142,N_20806);
nor UO_1921 (O_1921,N_21783,N_20919);
nand UO_1922 (O_1922,N_21020,N_19819);
and UO_1923 (O_1923,N_21092,N_19460);
xor UO_1924 (O_1924,N_20961,N_18818);
or UO_1925 (O_1925,N_23141,N_22572);
nand UO_1926 (O_1926,N_23171,N_22697);
and UO_1927 (O_1927,N_20607,N_22374);
nor UO_1928 (O_1928,N_20913,N_20358);
or UO_1929 (O_1929,N_21642,N_20031);
nor UO_1930 (O_1930,N_19150,N_19426);
or UO_1931 (O_1931,N_18980,N_22911);
and UO_1932 (O_1932,N_19757,N_20602);
or UO_1933 (O_1933,N_20870,N_18834);
and UO_1934 (O_1934,N_22794,N_18937);
or UO_1935 (O_1935,N_20567,N_19453);
and UO_1936 (O_1936,N_19226,N_24522);
and UO_1937 (O_1937,N_18831,N_24837);
and UO_1938 (O_1938,N_22039,N_23740);
nor UO_1939 (O_1939,N_19560,N_20047);
nand UO_1940 (O_1940,N_23257,N_19333);
xnor UO_1941 (O_1941,N_24808,N_24266);
xnor UO_1942 (O_1942,N_24353,N_18802);
xor UO_1943 (O_1943,N_24313,N_19051);
nor UO_1944 (O_1944,N_22253,N_19243);
and UO_1945 (O_1945,N_20560,N_23393);
xor UO_1946 (O_1946,N_22810,N_23083);
or UO_1947 (O_1947,N_19210,N_24198);
nor UO_1948 (O_1948,N_22215,N_21975);
and UO_1949 (O_1949,N_20836,N_18809);
nand UO_1950 (O_1950,N_24827,N_22837);
nand UO_1951 (O_1951,N_24456,N_21605);
or UO_1952 (O_1952,N_20813,N_21896);
or UO_1953 (O_1953,N_24900,N_22359);
nor UO_1954 (O_1954,N_23440,N_22075);
nand UO_1955 (O_1955,N_18759,N_21529);
nand UO_1956 (O_1956,N_24379,N_19572);
and UO_1957 (O_1957,N_22009,N_24678);
or UO_1958 (O_1958,N_20679,N_22968);
or UO_1959 (O_1959,N_24593,N_24613);
or UO_1960 (O_1960,N_20236,N_23501);
xnor UO_1961 (O_1961,N_23780,N_20735);
xor UO_1962 (O_1962,N_21771,N_23279);
or UO_1963 (O_1963,N_23394,N_23085);
xnor UO_1964 (O_1964,N_20109,N_24115);
and UO_1965 (O_1965,N_19489,N_22565);
nor UO_1966 (O_1966,N_21459,N_21321);
or UO_1967 (O_1967,N_19826,N_19498);
and UO_1968 (O_1968,N_21158,N_18880);
and UO_1969 (O_1969,N_20695,N_19900);
nor UO_1970 (O_1970,N_24418,N_21919);
nand UO_1971 (O_1971,N_24760,N_24293);
or UO_1972 (O_1972,N_21954,N_19689);
nor UO_1973 (O_1973,N_20451,N_19784);
and UO_1974 (O_1974,N_23335,N_20434);
or UO_1975 (O_1975,N_20120,N_20993);
nand UO_1976 (O_1976,N_23795,N_24282);
and UO_1977 (O_1977,N_24179,N_22585);
or UO_1978 (O_1978,N_23423,N_22487);
nand UO_1979 (O_1979,N_22485,N_19066);
and UO_1980 (O_1980,N_23621,N_21151);
xor UO_1981 (O_1981,N_21647,N_19354);
or UO_1982 (O_1982,N_23038,N_20918);
nor UO_1983 (O_1983,N_19023,N_20105);
xor UO_1984 (O_1984,N_21232,N_19948);
nand UO_1985 (O_1985,N_22369,N_21011);
and UO_1986 (O_1986,N_24209,N_19721);
or UO_1987 (O_1987,N_20691,N_21399);
or UO_1988 (O_1988,N_19957,N_22467);
or UO_1989 (O_1989,N_19141,N_19009);
nor UO_1990 (O_1990,N_19631,N_23205);
nor UO_1991 (O_1991,N_24054,N_22795);
and UO_1992 (O_1992,N_19767,N_21701);
nand UO_1993 (O_1993,N_23269,N_23173);
nor UO_1994 (O_1994,N_24496,N_24374);
xnor UO_1995 (O_1995,N_20848,N_19076);
nor UO_1996 (O_1996,N_21554,N_19349);
xnor UO_1997 (O_1997,N_20584,N_19183);
xnor UO_1998 (O_1998,N_22586,N_19480);
and UO_1999 (O_1999,N_24428,N_24103);
xor UO_2000 (O_2000,N_19202,N_20646);
or UO_2001 (O_2001,N_24866,N_20127);
nand UO_2002 (O_2002,N_22290,N_23054);
and UO_2003 (O_2003,N_24341,N_19305);
xnor UO_2004 (O_2004,N_23726,N_22801);
nor UO_2005 (O_2005,N_21493,N_24000);
xnor UO_2006 (O_2006,N_22761,N_21617);
nand UO_2007 (O_2007,N_22898,N_21106);
and UO_2008 (O_2008,N_24225,N_19634);
and UO_2009 (O_2009,N_21379,N_21475);
nand UO_2010 (O_2010,N_24571,N_22001);
and UO_2011 (O_2011,N_22643,N_20175);
and UO_2012 (O_2012,N_19084,N_21249);
or UO_2013 (O_2013,N_20115,N_21395);
xnor UO_2014 (O_2014,N_23678,N_18913);
or UO_2015 (O_2015,N_19728,N_22391);
xnor UO_2016 (O_2016,N_19239,N_24536);
nand UO_2017 (O_2017,N_20165,N_23959);
and UO_2018 (O_2018,N_20965,N_20724);
nor UO_2019 (O_2019,N_23981,N_21897);
or UO_2020 (O_2020,N_23198,N_23150);
and UO_2021 (O_2021,N_22731,N_22239);
or UO_2022 (O_2022,N_22228,N_23100);
or UO_2023 (O_2023,N_23328,N_22179);
and UO_2024 (O_2024,N_22010,N_22280);
nor UO_2025 (O_2025,N_18845,N_23556);
or UO_2026 (O_2026,N_24165,N_19473);
nand UO_2027 (O_2027,N_19707,N_21413);
nor UO_2028 (O_2028,N_23453,N_21115);
and UO_2029 (O_2029,N_18852,N_20303);
nand UO_2030 (O_2030,N_20811,N_24650);
and UO_2031 (O_2031,N_19947,N_20059);
or UO_2032 (O_2032,N_22644,N_22875);
or UO_2033 (O_2033,N_23442,N_21654);
xor UO_2034 (O_2034,N_22738,N_24478);
nor UO_2035 (O_2035,N_21063,N_20150);
or UO_2036 (O_2036,N_19171,N_23884);
xnor UO_2037 (O_2037,N_21133,N_23248);
xor UO_2038 (O_2038,N_24111,N_23937);
or UO_2039 (O_2039,N_22900,N_22664);
and UO_2040 (O_2040,N_24329,N_24632);
nand UO_2041 (O_2041,N_21861,N_23415);
and UO_2042 (O_2042,N_23769,N_19115);
xor UO_2043 (O_2043,N_23744,N_19933);
nor UO_2044 (O_2044,N_22130,N_19145);
nand UO_2045 (O_2045,N_24326,N_22234);
nand UO_2046 (O_2046,N_20285,N_20917);
xnor UO_2047 (O_2047,N_24034,N_20360);
and UO_2048 (O_2048,N_22061,N_21987);
or UO_2049 (O_2049,N_22365,N_21680);
xor UO_2050 (O_2050,N_23276,N_19846);
or UO_2051 (O_2051,N_20454,N_22385);
xnor UO_2052 (O_2052,N_21895,N_22914);
or UO_2053 (O_2053,N_24402,N_23779);
nand UO_2054 (O_2054,N_23600,N_23147);
nor UO_2055 (O_2055,N_19671,N_24913);
and UO_2056 (O_2056,N_24484,N_19326);
and UO_2057 (O_2057,N_24727,N_19870);
or UO_2058 (O_2058,N_18959,N_24908);
and UO_2059 (O_2059,N_21332,N_21716);
or UO_2060 (O_2060,N_20561,N_22515);
and UO_2061 (O_2061,N_20595,N_21579);
nor UO_2062 (O_2062,N_21300,N_23979);
xor UO_2063 (O_2063,N_22897,N_23686);
or UO_2064 (O_2064,N_24525,N_20542);
xnor UO_2065 (O_2065,N_23611,N_23943);
nand UO_2066 (O_2066,N_22770,N_23337);
nor UO_2067 (O_2067,N_21806,N_21718);
xor UO_2068 (O_2068,N_19696,N_20825);
nand UO_2069 (O_2069,N_22371,N_22570);
nand UO_2070 (O_2070,N_18835,N_24533);
and UO_2071 (O_2071,N_23485,N_24064);
or UO_2072 (O_2072,N_22015,N_24802);
and UO_2073 (O_2073,N_23484,N_23865);
xor UO_2074 (O_2074,N_19196,N_24997);
xnor UO_2075 (O_2075,N_19647,N_19918);
nand UO_2076 (O_2076,N_22111,N_21920);
xnor UO_2077 (O_2077,N_23293,N_22459);
and UO_2078 (O_2078,N_24932,N_20709);
nand UO_2079 (O_2079,N_18764,N_24962);
nand UO_2080 (O_2080,N_23655,N_20817);
nor UO_2081 (O_2081,N_19280,N_19908);
xor UO_2082 (O_2082,N_23241,N_24354);
or UO_2083 (O_2083,N_19655,N_20606);
nor UO_2084 (O_2084,N_21004,N_18947);
or UO_2085 (O_2085,N_19127,N_19037);
nand UO_2086 (O_2086,N_23590,N_23358);
xor UO_2087 (O_2087,N_24347,N_21003);
xor UO_2088 (O_2088,N_23021,N_21071);
nor UO_2089 (O_2089,N_24905,N_20392);
or UO_2090 (O_2090,N_24666,N_24907);
or UO_2091 (O_2091,N_21574,N_24790);
xor UO_2092 (O_2092,N_24268,N_19181);
and UO_2093 (O_2093,N_23034,N_21262);
and UO_2094 (O_2094,N_21548,N_24519);
nand UO_2095 (O_2095,N_24989,N_24152);
nand UO_2096 (O_2096,N_24817,N_19245);
and UO_2097 (O_2097,N_23444,N_22153);
and UO_2098 (O_2098,N_18827,N_24487);
nand UO_2099 (O_2099,N_20182,N_20056);
nor UO_2100 (O_2100,N_24864,N_23783);
and UO_2101 (O_2101,N_24356,N_22556);
and UO_2102 (O_2102,N_20491,N_21711);
nor UO_2103 (O_2103,N_19510,N_20478);
or UO_2104 (O_2104,N_20527,N_18828);
and UO_2105 (O_2105,N_24136,N_19528);
or UO_2106 (O_2106,N_21019,N_23345);
or UO_2107 (O_2107,N_24135,N_20692);
nor UO_2108 (O_2108,N_24651,N_22536);
nor UO_2109 (O_2109,N_24096,N_21221);
or UO_2110 (O_2110,N_24868,N_22709);
xor UO_2111 (O_2111,N_19495,N_20544);
nor UO_2112 (O_2112,N_20225,N_21755);
and UO_2113 (O_2113,N_19309,N_19975);
or UO_2114 (O_2114,N_22921,N_22734);
nand UO_2115 (O_2115,N_20772,N_21930);
nand UO_2116 (O_2116,N_18963,N_19962);
nand UO_2117 (O_2117,N_19735,N_19376);
nor UO_2118 (O_2118,N_24614,N_21832);
xnor UO_2119 (O_2119,N_22144,N_18849);
xnor UO_2120 (O_2120,N_20865,N_23618);
xnor UO_2121 (O_2121,N_24243,N_22091);
xor UO_2122 (O_2122,N_23409,N_18836);
and UO_2123 (O_2123,N_20521,N_24621);
or UO_2124 (O_2124,N_24719,N_19172);
xnor UO_2125 (O_2125,N_18983,N_19491);
xnor UO_2126 (O_2126,N_18839,N_20737);
and UO_2127 (O_2127,N_23494,N_23200);
nand UO_2128 (O_2128,N_21770,N_23546);
nor UO_2129 (O_2129,N_18798,N_23416);
or UO_2130 (O_2130,N_21487,N_20155);
nand UO_2131 (O_2131,N_19434,N_23118);
nor UO_2132 (O_2132,N_24162,N_19624);
nor UO_2133 (O_2133,N_22947,N_20619);
and UO_2134 (O_2134,N_24852,N_20654);
or UO_2135 (O_2135,N_19256,N_23467);
nand UO_2136 (O_2136,N_24495,N_19781);
nand UO_2137 (O_2137,N_20974,N_24044);
and UO_2138 (O_2138,N_23410,N_19513);
nor UO_2139 (O_2139,N_20222,N_22156);
nand UO_2140 (O_2140,N_20930,N_23273);
nand UO_2141 (O_2141,N_18796,N_23800);
nor UO_2142 (O_2142,N_23024,N_19889);
xnor UO_2143 (O_2143,N_23297,N_23274);
nand UO_2144 (O_2144,N_24708,N_23966);
nand UO_2145 (O_2145,N_18909,N_24763);
nor UO_2146 (O_2146,N_23374,N_20469);
nand UO_2147 (O_2147,N_22724,N_22450);
and UO_2148 (O_2148,N_24965,N_21580);
and UO_2149 (O_2149,N_20571,N_22021);
or UO_2150 (O_2150,N_23126,N_24348);
nor UO_2151 (O_2151,N_21777,N_19581);
and UO_2152 (O_2152,N_22624,N_24789);
xor UO_2153 (O_2153,N_24676,N_19490);
or UO_2154 (O_2154,N_23615,N_22213);
nor UO_2155 (O_2155,N_23732,N_24831);
nand UO_2156 (O_2156,N_20005,N_22199);
nor UO_2157 (O_2157,N_22120,N_22902);
and UO_2158 (O_2158,N_19986,N_18816);
xor UO_2159 (O_2159,N_19228,N_24338);
and UO_2160 (O_2160,N_19956,N_20818);
nand UO_2161 (O_2161,N_23782,N_24967);
nor UO_2162 (O_2162,N_21292,N_23647);
nor UO_2163 (O_2163,N_23359,N_22705);
xor UO_2164 (O_2164,N_18956,N_22225);
xnor UO_2165 (O_2165,N_19778,N_24274);
or UO_2166 (O_2166,N_20838,N_19697);
or UO_2167 (O_2167,N_20349,N_24498);
or UO_2168 (O_2168,N_24526,N_24062);
and UO_2169 (O_2169,N_18795,N_21676);
or UO_2170 (O_2170,N_22858,N_21452);
and UO_2171 (O_2171,N_24128,N_24554);
and UO_2172 (O_2172,N_23099,N_21229);
nand UO_2173 (O_2173,N_20408,N_19803);
nor UO_2174 (O_2174,N_19896,N_20652);
nand UO_2175 (O_2175,N_18951,N_23989);
or UO_2176 (O_2176,N_23225,N_22872);
nand UO_2177 (O_2177,N_23512,N_21531);
xor UO_2178 (O_2178,N_20235,N_24235);
and UO_2179 (O_2179,N_21490,N_18946);
nor UO_2180 (O_2180,N_23074,N_22494);
or UO_2181 (O_2181,N_22344,N_24755);
and UO_2182 (O_2182,N_23873,N_21183);
nand UO_2183 (O_2183,N_23683,N_22753);
or UO_2184 (O_2184,N_23534,N_24043);
xnor UO_2185 (O_2185,N_22354,N_20941);
nand UO_2186 (O_2186,N_23657,N_23086);
and UO_2187 (O_2187,N_19472,N_22927);
or UO_2188 (O_2188,N_19251,N_20440);
xor UO_2189 (O_2189,N_21974,N_19894);
and UO_2190 (O_2190,N_19893,N_22393);
or UO_2191 (O_2191,N_20778,N_22759);
nand UO_2192 (O_2192,N_18820,N_23654);
nor UO_2193 (O_2193,N_21581,N_23812);
xor UO_2194 (O_2194,N_21996,N_20911);
nand UO_2195 (O_2195,N_20802,N_23719);
or UO_2196 (O_2196,N_20689,N_19785);
or UO_2197 (O_2197,N_24871,N_19271);
xor UO_2198 (O_2198,N_23418,N_24828);
or UO_2199 (O_2199,N_19504,N_24292);
or UO_2200 (O_2200,N_22657,N_20166);
nor UO_2201 (O_2201,N_20185,N_22387);
nand UO_2202 (O_2202,N_21505,N_22330);
xor UO_2203 (O_2203,N_19553,N_19960);
nand UO_2204 (O_2204,N_24876,N_20022);
nand UO_2205 (O_2205,N_19449,N_23549);
or UO_2206 (O_2206,N_21827,N_23623);
nor UO_2207 (O_2207,N_21951,N_23606);
and UO_2208 (O_2208,N_23652,N_21520);
nand UO_2209 (O_2209,N_23676,N_21890);
or UO_2210 (O_2210,N_19482,N_19558);
or UO_2211 (O_2211,N_22016,N_23134);
and UO_2212 (O_2212,N_20095,N_21037);
nor UO_2213 (O_2213,N_24639,N_18797);
xor UO_2214 (O_2214,N_22747,N_24897);
xor UO_2215 (O_2215,N_21266,N_20385);
nand UO_2216 (O_2216,N_21521,N_24539);
nand UO_2217 (O_2217,N_23082,N_20804);
or UO_2218 (O_2218,N_23388,N_21725);
or UO_2219 (O_2219,N_21328,N_21834);
or UO_2220 (O_2220,N_22011,N_21396);
nand UO_2221 (O_2221,N_23052,N_24572);
and UO_2222 (O_2222,N_20775,N_19131);
and UO_2223 (O_2223,N_24319,N_20313);
and UO_2224 (O_2224,N_19949,N_19568);
or UO_2225 (O_2225,N_19476,N_23103);
and UO_2226 (O_2226,N_24318,N_22832);
nand UO_2227 (O_2227,N_19083,N_21786);
nand UO_2228 (O_2228,N_22478,N_21995);
xor UO_2229 (O_2229,N_21134,N_20793);
or UO_2230 (O_2230,N_19914,N_22455);
or UO_2231 (O_2231,N_24331,N_23477);
and UO_2232 (O_2232,N_20427,N_18926);
or UO_2233 (O_2233,N_19233,N_19149);
nand UO_2234 (O_2234,N_23030,N_23435);
or UO_2235 (O_2235,N_21723,N_24241);
xnor UO_2236 (O_2236,N_22306,N_21609);
or UO_2237 (O_2237,N_22495,N_20180);
nand UO_2238 (O_2238,N_22424,N_22332);
and UO_2239 (O_2239,N_20174,N_20671);
or UO_2240 (O_2240,N_24359,N_20739);
or UO_2241 (O_2241,N_19412,N_22907);
nor UO_2242 (O_2242,N_19269,N_20929);
xor UO_2243 (O_2243,N_19562,N_19559);
or UO_2244 (O_2244,N_21290,N_20093);
or UO_2245 (O_2245,N_21638,N_18763);
xnor UO_2246 (O_2246,N_24169,N_21938);
and UO_2247 (O_2247,N_19661,N_21555);
nand UO_2248 (O_2248,N_23499,N_20757);
xor UO_2249 (O_2249,N_21048,N_20668);
or UO_2250 (O_2250,N_21810,N_22918);
nand UO_2251 (O_2251,N_24011,N_20138);
nor UO_2252 (O_2252,N_23589,N_19322);
nand UO_2253 (O_2253,N_24605,N_24361);
xnor UO_2254 (O_2254,N_23066,N_24362);
nor UO_2255 (O_2255,N_22133,N_23823);
or UO_2256 (O_2256,N_21049,N_20840);
xor UO_2257 (O_2257,N_24824,N_20513);
and UO_2258 (O_2258,N_21273,N_24185);
and UO_2259 (O_2259,N_23856,N_24275);
and UO_2260 (O_2260,N_20677,N_23020);
xor UO_2261 (O_2261,N_22406,N_21594);
xnor UO_2262 (O_2262,N_24648,N_21556);
nor UO_2263 (O_2263,N_21337,N_23231);
nand UO_2264 (O_2264,N_24030,N_20463);
xnor UO_2265 (O_2265,N_23217,N_19871);
or UO_2266 (O_2266,N_20647,N_23391);
or UO_2267 (O_2267,N_23229,N_24310);
nand UO_2268 (O_2268,N_22113,N_21668);
xnor UO_2269 (O_2269,N_24398,N_18859);
and UO_2270 (O_2270,N_22778,N_21670);
xnor UO_2271 (O_2271,N_18915,N_19492);
nor UO_2272 (O_2272,N_21058,N_19938);
or UO_2273 (O_2273,N_20832,N_22046);
or UO_2274 (O_2274,N_24949,N_21541);
nor UO_2275 (O_2275,N_21628,N_22856);
or UO_2276 (O_2276,N_19012,N_19161);
and UO_2277 (O_2277,N_24537,N_23775);
nand UO_2278 (O_2278,N_21000,N_22382);
nand UO_2279 (O_2279,N_18921,N_24761);
xor UO_2280 (O_2280,N_22484,N_20256);
or UO_2281 (O_2281,N_23706,N_19743);
and UO_2282 (O_2282,N_22690,N_19936);
or UO_2283 (O_2283,N_22752,N_19720);
xor UO_2284 (O_2284,N_19364,N_22493);
xnor UO_2285 (O_2285,N_20551,N_23672);
xor UO_2286 (O_2286,N_23247,N_24607);
and UO_2287 (O_2287,N_24671,N_19026);
and UO_2288 (O_2288,N_21795,N_22523);
xnor UO_2289 (O_2289,N_24303,N_22080);
and UO_2290 (O_2290,N_24385,N_23613);
xnor UO_2291 (O_2291,N_20693,N_19375);
or UO_2292 (O_2292,N_20956,N_24637);
or UO_2293 (O_2293,N_19747,N_22073);
nand UO_2294 (O_2294,N_22121,N_20443);
or UO_2295 (O_2295,N_20023,N_24409);
and UO_2296 (O_2296,N_23395,N_22497);
xnor UO_2297 (O_2297,N_19586,N_23685);
or UO_2298 (O_2298,N_20682,N_19218);
xor UO_2299 (O_2299,N_24453,N_21807);
xor UO_2300 (O_2300,N_24973,N_22254);
nor UO_2301 (O_2301,N_21953,N_19811);
xor UO_2302 (O_2302,N_23101,N_21021);
xnor UO_2303 (O_2303,N_22161,N_21138);
nor UO_2304 (O_2304,N_20721,N_21204);
or UO_2305 (O_2305,N_19828,N_24171);
nor UO_2306 (O_2306,N_23766,N_22960);
and UO_2307 (O_2307,N_22103,N_19195);
nand UO_2308 (O_2308,N_20473,N_21559);
xnor UO_2309 (O_2309,N_23282,N_22638);
and UO_2310 (O_2310,N_21182,N_22425);
or UO_2311 (O_2311,N_22136,N_21720);
or UO_2312 (O_2312,N_23224,N_20350);
xor UO_2313 (O_2313,N_24258,N_24515);
or UO_2314 (O_2314,N_23838,N_21741);
and UO_2315 (O_2315,N_24002,N_22679);
or UO_2316 (O_2316,N_21469,N_20097);
nor UO_2317 (O_2317,N_23990,N_24977);
and UO_2318 (O_2318,N_22852,N_23938);
nand UO_2319 (O_2319,N_22979,N_23888);
nor UO_2320 (O_2320,N_19885,N_23098);
or UO_2321 (O_2321,N_21028,N_20644);
and UO_2322 (O_2322,N_23143,N_19065);
nand UO_2323 (O_2323,N_21105,N_24408);
nand UO_2324 (O_2324,N_22938,N_22647);
xor UO_2325 (O_2325,N_20578,N_20080);
or UO_2326 (O_2326,N_23673,N_23940);
and UO_2327 (O_2327,N_23339,N_18800);
nand UO_2328 (O_2328,N_21814,N_21465);
xor UO_2329 (O_2329,N_18942,N_21596);
nand UO_2330 (O_2330,N_21734,N_19466);
nand UO_2331 (O_2331,N_18808,N_21434);
nor UO_2332 (O_2332,N_22543,N_20819);
or UO_2333 (O_2333,N_20641,N_23811);
or UO_2334 (O_2334,N_20612,N_20799);
or UO_2335 (O_2335,N_22316,N_19112);
or UO_2336 (O_2336,N_19148,N_24788);
nor UO_2337 (O_2337,N_24670,N_23392);
and UO_2338 (O_2338,N_19872,N_21319);
xor UO_2339 (O_2339,N_19888,N_23544);
nand UO_2340 (O_2340,N_19463,N_23658);
xnor UO_2341 (O_2341,N_19285,N_24714);
and UO_2342 (O_2342,N_24691,N_24033);
or UO_2343 (O_2343,N_20944,N_22632);
xor UO_2344 (O_2344,N_20805,N_22812);
nand UO_2345 (O_2345,N_22310,N_22020);
and UO_2346 (O_2346,N_23255,N_21553);
nand UO_2347 (O_2347,N_22439,N_21272);
nor UO_2348 (O_2348,N_20598,N_19249);
or UO_2349 (O_2349,N_21535,N_22970);
and UO_2350 (O_2350,N_19496,N_22598);
nand UO_2351 (O_2351,N_21793,N_24040);
and UO_2352 (O_2352,N_22457,N_21652);
xor UO_2353 (O_2353,N_20333,N_21863);
nor UO_2354 (O_2354,N_21463,N_19119);
or UO_2355 (O_2355,N_21724,N_22333);
nor UO_2356 (O_2356,N_21095,N_19857);
or UO_2357 (O_2357,N_21201,N_22712);
nor UO_2358 (O_2358,N_18898,N_21166);
xnor UO_2359 (O_2359,N_21694,N_20369);
xnor UO_2360 (O_2360,N_21052,N_24180);
xnor UO_2361 (O_2361,N_21808,N_23382);
and UO_2362 (O_2362,N_23469,N_23455);
and UO_2363 (O_2363,N_21153,N_21794);
and UO_2364 (O_2364,N_24387,N_21318);
nor UO_2365 (O_2365,N_23551,N_23115);
and UO_2366 (O_2366,N_20203,N_20868);
nand UO_2367 (O_2367,N_24867,N_20379);
nor UO_2368 (O_2368,N_20698,N_23581);
xor UO_2369 (O_2369,N_21961,N_22826);
or UO_2370 (O_2370,N_20850,N_23370);
xor UO_2371 (O_2371,N_18838,N_22275);
or UO_2372 (O_2372,N_23329,N_21621);
nor UO_2373 (O_2373,N_19189,N_20228);
nand UO_2374 (O_2374,N_18778,N_19265);
nor UO_2375 (O_2375,N_21060,N_22721);
and UO_2376 (O_2376,N_24109,N_21751);
xor UO_2377 (O_2377,N_22386,N_20453);
nand UO_2378 (O_2378,N_24733,N_21226);
and UO_2379 (O_2379,N_24542,N_20723);
and UO_2380 (O_2380,N_24187,N_22548);
and UO_2381 (O_2381,N_22421,N_23002);
xor UO_2382 (O_2382,N_20280,N_23914);
and UO_2383 (O_2383,N_24061,N_20407);
and UO_2384 (O_2384,N_22269,N_21833);
nand UO_2385 (O_2385,N_23522,N_23861);
nand UO_2386 (O_2386,N_19193,N_19334);
or UO_2387 (O_2387,N_18870,N_19705);
and UO_2388 (O_2388,N_23240,N_18779);
and UO_2389 (O_2389,N_23040,N_19167);
nand UO_2390 (O_2390,N_24403,N_24010);
xnor UO_2391 (O_2391,N_21745,N_19440);
nand UO_2392 (O_2392,N_19657,N_20183);
xnor UO_2393 (O_2393,N_24943,N_23656);
nand UO_2394 (O_2394,N_24854,N_20294);
nor UO_2395 (O_2395,N_24322,N_19662);
and UO_2396 (O_2396,N_22957,N_20048);
xnor UO_2397 (O_2397,N_23302,N_21278);
nand UO_2398 (O_2398,N_24803,N_19118);
xor UO_2399 (O_2399,N_21164,N_21817);
xnor UO_2400 (O_2400,N_24581,N_21299);
or UO_2401 (O_2401,N_20755,N_23793);
nor UO_2402 (O_2402,N_23752,N_20213);
and UO_2403 (O_2403,N_18762,N_24092);
and UO_2404 (O_2404,N_23165,N_22805);
and UO_2405 (O_2405,N_20890,N_22394);
xnor UO_2406 (O_2406,N_24619,N_21513);
nor UO_2407 (O_2407,N_20304,N_19090);
nor UO_2408 (O_2408,N_22739,N_22357);
and UO_2409 (O_2409,N_18872,N_19393);
nand UO_2410 (O_2410,N_22422,N_20286);
xor UO_2411 (O_2411,N_24709,N_19690);
and UO_2412 (O_2412,N_20984,N_21388);
xnor UO_2413 (O_2413,N_20482,N_24270);
and UO_2414 (O_2414,N_19041,N_19849);
nand UO_2415 (O_2415,N_19580,N_22343);
xor UO_2416 (O_2416,N_24555,N_19863);
or UO_2417 (O_2417,N_23438,N_21881);
xnor UO_2418 (O_2418,N_19797,N_19730);
xor UO_2419 (O_2419,N_24640,N_22926);
nand UO_2420 (O_2420,N_20223,N_23980);
nor UO_2421 (O_2421,N_19048,N_19015);
and UO_2422 (O_2422,N_19627,N_18776);
nor UO_2423 (O_2423,N_23050,N_23830);
nand UO_2424 (O_2424,N_19663,N_24856);
nor UO_2425 (O_2425,N_20490,N_21876);
nand UO_2426 (O_2426,N_20461,N_22279);
nand UO_2427 (O_2427,N_22383,N_21766);
xnor UO_2428 (O_2428,N_22214,N_20103);
or UO_2429 (O_2429,N_24723,N_21747);
nand UO_2430 (O_2430,N_22126,N_19369);
nor UO_2431 (O_2431,N_24153,N_19958);
and UO_2432 (O_2432,N_21620,N_22696);
or UO_2433 (O_2433,N_22775,N_20338);
xor UO_2434 (O_2434,N_19074,N_19056);
or UO_2435 (O_2435,N_21172,N_24677);
or UO_2436 (O_2436,N_21614,N_20945);
nand UO_2437 (O_2437,N_20768,N_22198);
xor UO_2438 (O_2438,N_19543,N_20678);
and UO_2439 (O_2439,N_22851,N_21752);
or UO_2440 (O_2440,N_23300,N_23474);
and UO_2441 (O_2441,N_24345,N_23481);
or UO_2442 (O_2442,N_21340,N_23828);
nor UO_2443 (O_2443,N_22835,N_19129);
nand UO_2444 (O_2444,N_19004,N_24441);
or UO_2445 (O_2445,N_24006,N_19693);
nand UO_2446 (O_2446,N_24705,N_22065);
xnor UO_2447 (O_2447,N_23598,N_24625);
nand UO_2448 (O_2448,N_24521,N_20322);
xor UO_2449 (O_2449,N_22669,N_18815);
or UO_2450 (O_2450,N_19107,N_22100);
nand UO_2451 (O_2451,N_21818,N_22954);
nand UO_2452 (O_2452,N_18927,N_22958);
xnor UO_2453 (O_2453,N_22217,N_20503);
or UO_2454 (O_2454,N_20018,N_20457);
nor UO_2455 (O_2455,N_22995,N_24754);
nand UO_2456 (O_2456,N_21985,N_19601);
nand UO_2457 (O_2457,N_24841,N_24480);
nor UO_2458 (O_2458,N_19225,N_22674);
nor UO_2459 (O_2459,N_19386,N_23709);
nor UO_2460 (O_2460,N_24019,N_23422);
nor UO_2461 (O_2461,N_21504,N_21322);
or UO_2462 (O_2462,N_21083,N_20519);
xor UO_2463 (O_2463,N_24366,N_20205);
nand UO_2464 (O_2464,N_20844,N_21775);
and UO_2465 (O_2465,N_21598,N_18939);
and UO_2466 (O_2466,N_24976,N_20596);
and UO_2467 (O_2467,N_21068,N_20901);
xor UO_2468 (O_2468,N_20823,N_21030);
nand UO_2469 (O_2469,N_21446,N_24191);
or UO_2470 (O_2470,N_20515,N_19525);
nand UO_2471 (O_2471,N_24669,N_23711);
or UO_2472 (O_2472,N_24681,N_24684);
or UO_2473 (O_2473,N_23354,N_19268);
or UO_2474 (O_2474,N_22869,N_19793);
nand UO_2475 (O_2475,N_22099,N_24930);
or UO_2476 (O_2476,N_20483,N_21018);
nor UO_2477 (O_2477,N_19775,N_19185);
and UO_2478 (O_2478,N_20639,N_24952);
nor UO_2479 (O_2479,N_24395,N_21512);
xor UO_2480 (O_2480,N_21252,N_19621);
or UO_2481 (O_2481,N_18990,N_22604);
nor UO_2482 (O_2482,N_19122,N_23193);
xnor UO_2483 (O_2483,N_24686,N_24065);
and UO_2484 (O_2484,N_20665,N_19034);
xnor UO_2485 (O_2485,N_20898,N_19263);
or UO_2486 (O_2486,N_24517,N_20008);
nor UO_2487 (O_2487,N_19668,N_20240);
nand UO_2488 (O_2488,N_22796,N_20821);
or UO_2489 (O_2489,N_18787,N_21315);
and UO_2490 (O_2490,N_24312,N_20508);
nor UO_2491 (O_2491,N_22846,N_19729);
nand UO_2492 (O_2492,N_24531,N_20326);
xor UO_2493 (O_2493,N_22098,N_19731);
nor UO_2494 (O_2494,N_22654,N_22964);
nor UO_2495 (O_2495,N_24794,N_18782);
and UO_2496 (O_2496,N_23845,N_24071);
and UO_2497 (O_2497,N_21173,N_22741);
nor UO_2498 (O_2498,N_22959,N_19952);
nor UO_2499 (O_2499,N_20574,N_20417);
xor UO_2500 (O_2500,N_24474,N_21517);
xnor UO_2501 (O_2501,N_24874,N_19257);
nand UO_2502 (O_2502,N_20617,N_24559);
nor UO_2503 (O_2503,N_24701,N_19618);
xnor UO_2504 (O_2504,N_21981,N_19589);
nor UO_2505 (O_2505,N_22068,N_21149);
and UO_2506 (O_2506,N_19016,N_24528);
nand UO_2507 (O_2507,N_23619,N_22030);
and UO_2508 (O_2508,N_19155,N_22362);
nand UO_2509 (O_2509,N_20081,N_19670);
nor UO_2510 (O_2510,N_20387,N_19028);
xnor UO_2511 (O_2511,N_21051,N_20662);
nand UO_2512 (O_2512,N_22318,N_21697);
or UO_2513 (O_2513,N_22780,N_24499);
or UO_2514 (O_2514,N_23645,N_23214);
nand UO_2515 (O_2515,N_19139,N_24476);
and UO_2516 (O_2516,N_20055,N_22533);
nand UO_2517 (O_2517,N_21633,N_18974);
xor UO_2518 (O_2518,N_20404,N_24552);
nand UO_2519 (O_2519,N_23197,N_24273);
and UO_2520 (O_2520,N_20943,N_20269);
xnor UO_2521 (O_2521,N_23698,N_24995);
or UO_2522 (O_2522,N_24324,N_23331);
or UO_2523 (O_2523,N_22056,N_20744);
xnor UO_2524 (O_2524,N_22295,N_19742);
nand UO_2525 (O_2525,N_23877,N_24296);
or UO_2526 (O_2526,N_23984,N_21231);
nor UO_2527 (O_2527,N_18883,N_21224);
xnor UO_2528 (O_2528,N_21649,N_24148);
xor UO_2529 (O_2529,N_24804,N_20487);
nor UO_2530 (O_2530,N_22219,N_23176);
nand UO_2531 (O_2531,N_23316,N_19310);
nor UO_2532 (O_2532,N_23159,N_24724);
or UO_2533 (O_2533,N_21590,N_22766);
nor UO_2534 (O_2534,N_21075,N_21311);
xnor UO_2535 (O_2535,N_22639,N_24696);
or UO_2536 (O_2536,N_20259,N_19821);
xor UO_2537 (O_2537,N_19368,N_21284);
nor UO_2538 (O_2538,N_24948,N_24842);
and UO_2539 (O_2539,N_18977,N_23661);
and UO_2540 (O_2540,N_22730,N_19424);
xor UO_2541 (O_2541,N_22714,N_21301);
nor UO_2542 (O_2542,N_20062,N_21233);
nor UO_2543 (O_2543,N_23445,N_22559);
and UO_2544 (O_2544,N_22732,N_24884);
and UO_2545 (O_2545,N_22086,N_22934);
and UO_2546 (O_2546,N_22172,N_23408);
nand UO_2547 (O_2547,N_22414,N_23564);
and UO_2548 (O_2548,N_22760,N_21170);
or UO_2549 (O_2549,N_20011,N_20660);
xnor UO_2550 (O_2550,N_21922,N_21799);
nand UO_2551 (O_2551,N_23835,N_24699);
or UO_2552 (O_2552,N_24106,N_20119);
and UO_2553 (O_2553,N_21978,N_19760);
xor UO_2554 (O_2554,N_24121,N_21234);
nand UO_2555 (O_2555,N_22104,N_19135);
nor UO_2556 (O_2556,N_22050,N_24229);
or UO_2557 (O_2557,N_23425,N_20102);
or UO_2558 (O_2558,N_22649,N_22325);
or UO_2559 (O_2559,N_21050,N_19612);
or UO_2560 (O_2560,N_18890,N_21889);
and UO_2561 (O_2561,N_21362,N_22574);
nand UO_2562 (O_2562,N_20624,N_24412);
nor UO_2563 (O_2563,N_24053,N_21886);
or UO_2564 (O_2564,N_20666,N_19520);
nand UO_2565 (O_2565,N_21150,N_21432);
nor UO_2566 (O_2566,N_24929,N_19276);
and UO_2567 (O_2567,N_21845,N_23309);
or UO_2568 (O_2568,N_23962,N_18949);
and UO_2569 (O_2569,N_19617,N_22593);
or UO_2570 (O_2570,N_22474,N_23817);
nand UO_2571 (O_2571,N_23665,N_21829);
or UO_2572 (O_2572,N_24811,N_19978);
xor UO_2573 (O_2573,N_24489,N_20181);
nand UO_2574 (O_2574,N_22423,N_21731);
and UO_2575 (O_2575,N_20039,N_22539);
or UO_2576 (O_2576,N_21310,N_24563);
nand UO_2577 (O_2577,N_22655,N_19691);
and UO_2578 (O_2578,N_21497,N_19292);
nor UO_2579 (O_2579,N_22854,N_23287);
or UO_2580 (O_2580,N_24192,N_23478);
or UO_2581 (O_2581,N_23461,N_20711);
nor UO_2582 (O_2582,N_19359,N_24716);
nand UO_2583 (O_2583,N_23561,N_22799);
nand UO_2584 (O_2584,N_22166,N_20088);
nor UO_2585 (O_2585,N_22303,N_21393);
or UO_2586 (O_2586,N_23003,N_20132);
xor UO_2587 (O_2587,N_22087,N_23496);
or UO_2588 (O_2588,N_22535,N_19683);
nor UO_2589 (O_2589,N_21046,N_20435);
nand UO_2590 (O_2590,N_22134,N_23140);
nand UO_2591 (O_2591,N_20990,N_19913);
xor UO_2592 (O_2592,N_24626,N_19503);
xor UO_2593 (O_2593,N_21067,N_20148);
and UO_2594 (O_2594,N_24252,N_21001);
and UO_2595 (O_2595,N_20308,N_19512);
or UO_2596 (O_2596,N_23324,N_24406);
xor UO_2597 (O_2597,N_21887,N_22718);
nand UO_2598 (O_2598,N_24177,N_21384);
or UO_2599 (O_2599,N_21462,N_22991);
or UO_2600 (O_2600,N_21569,N_20347);
nor UO_2601 (O_2601,N_23630,N_22962);
nor UO_2602 (O_2602,N_23135,N_19416);
and UO_2603 (O_2603,N_24449,N_24853);
and UO_2604 (O_2604,N_23271,N_23771);
and UO_2605 (O_2605,N_24545,N_24919);
nand UO_2606 (O_2606,N_24079,N_21603);
nand UO_2607 (O_2607,N_21717,N_22024);
and UO_2608 (O_2608,N_22124,N_19103);
or UO_2609 (O_2609,N_21093,N_19110);
or UO_2610 (O_2610,N_20773,N_24309);
and UO_2611 (O_2611,N_23073,N_20543);
and UO_2612 (O_2612,N_23152,N_24888);
xor UO_2613 (O_2613,N_19681,N_19213);
or UO_2614 (O_2614,N_19822,N_20199);
xnor UO_2615 (O_2615,N_24601,N_21899);
nor UO_2616 (O_2616,N_21608,N_24365);
nor UO_2617 (O_2617,N_24437,N_24221);
or UO_2618 (O_2618,N_18858,N_19070);
xor UO_2619 (O_2619,N_23243,N_21820);
or UO_2620 (O_2620,N_24242,N_24611);
xor UO_2621 (O_2621,N_24075,N_21357);
nand UO_2622 (O_2622,N_19927,N_19389);
nor UO_2623 (O_2623,N_24021,N_22396);
xor UO_2624 (O_2624,N_22492,N_20317);
nor UO_2625 (O_2625,N_19398,N_22401);
or UO_2626 (O_2626,N_20253,N_20368);
nand UO_2627 (O_2627,N_19159,N_23209);
nor UO_2628 (O_2628,N_23513,N_22246);
nor UO_2629 (O_2629,N_19303,N_21736);
xnor UO_2630 (O_2630,N_22490,N_19698);
xnor UO_2631 (O_2631,N_24458,N_21280);
nor UO_2632 (O_2632,N_18765,N_23413);
or UO_2633 (O_2633,N_22191,N_23592);
nand UO_2634 (O_2634,N_23860,N_22836);
and UO_2635 (O_2635,N_23595,N_20754);
nor UO_2636 (O_2636,N_22140,N_20829);
or UO_2637 (O_2637,N_21422,N_24630);
xnor UO_2638 (O_2638,N_22090,N_20696);
nor UO_2639 (O_2639,N_24622,N_18988);
nor UO_2640 (O_2640,N_21181,N_21584);
nand UO_2641 (O_2641,N_19744,N_18985);
and UO_2642 (O_2642,N_19471,N_24097);
nand UO_2643 (O_2643,N_21538,N_23292);
nand UO_2644 (O_2644,N_23077,N_19726);
or UO_2645 (O_2645,N_21480,N_19756);
nor UO_2646 (O_2646,N_23731,N_20847);
or UO_2647 (O_2647,N_22511,N_18938);
or UO_2648 (O_2648,N_21507,N_21791);
or UO_2649 (O_2649,N_21445,N_20593);
and UO_2650 (O_2650,N_21002,N_23280);
xor UO_2651 (O_2651,N_22476,N_20582);
nand UO_2652 (O_2652,N_19469,N_24308);
and UO_2653 (O_2653,N_23155,N_19313);
and UO_2654 (O_2654,N_23620,N_24227);
or UO_2655 (O_2655,N_21809,N_21991);
or UO_2656 (O_2656,N_22346,N_19075);
or UO_2657 (O_2657,N_20106,N_20952);
and UO_2658 (O_2658,N_22966,N_20114);
nand UO_2659 (O_2659,N_20642,N_18873);
nor UO_2660 (O_2660,N_20537,N_22062);
nor UO_2661 (O_2661,N_24396,N_22506);
or UO_2662 (O_2662,N_23396,N_20060);
xnor UO_2663 (O_2663,N_18892,N_21116);
or UO_2664 (O_2664,N_23170,N_23275);
xnor UO_2665 (O_2665,N_24297,N_20129);
or UO_2666 (O_2666,N_22177,N_23227);
or UO_2667 (O_2667,N_21842,N_20597);
and UO_2668 (O_2668,N_23639,N_24721);
or UO_2669 (O_2669,N_19664,N_18790);
and UO_2670 (O_2670,N_20314,N_23195);
nor UO_2671 (O_2671,N_20069,N_20856);
nor UO_2672 (O_2672,N_24503,N_19774);
and UO_2673 (O_2673,N_19374,N_20021);
nand UO_2674 (O_2674,N_21192,N_20357);
or UO_2675 (O_2675,N_18932,N_20569);
or UO_2676 (O_2676,N_18841,N_22510);
and UO_2677 (O_2677,N_22291,N_22833);
nand UO_2678 (O_2678,N_19983,N_23961);
xnor UO_2679 (O_2679,N_19642,N_21593);
nand UO_2680 (O_2680,N_24391,N_23234);
and UO_2681 (O_2681,N_21821,N_19973);
and UO_2682 (O_2682,N_19335,N_23669);
xor UO_2683 (O_2683,N_21530,N_23390);
xor UO_2684 (O_2684,N_21944,N_24538);
or UO_2685 (O_2685,N_22641,N_21213);
or UO_2686 (O_2686,N_22451,N_18867);
and UO_2687 (O_2687,N_21906,N_24848);
nand UO_2688 (O_2688,N_21878,N_21190);
nand UO_2689 (O_2689,N_22045,N_20511);
xnor UO_2690 (O_2690,N_23286,N_24457);
nand UO_2691 (O_2691,N_19032,N_20949);
nor UO_2692 (O_2692,N_20618,N_24658);
nor UO_2693 (O_2693,N_21304,N_20998);
and UO_2694 (O_2694,N_19816,N_21286);
nand UO_2695 (O_2695,N_24661,N_20936);
nand UO_2696 (O_2696,N_22850,N_19684);
nor UO_2697 (O_2697,N_23236,N_18813);
nor UO_2698 (O_2698,N_21220,N_21405);
nor UO_2699 (O_2699,N_21635,N_19991);
nor UO_2700 (O_2700,N_21061,N_21458);
xor UO_2701 (O_2701,N_21241,N_20497);
nand UO_2702 (O_2702,N_19253,N_23294);
xor UO_2703 (O_2703,N_23014,N_24383);
xor UO_2704 (O_2704,N_24830,N_23900);
nor UO_2705 (O_2705,N_19419,N_20449);
or UO_2706 (O_2706,N_23992,N_21924);
and UO_2707 (O_2707,N_18933,N_24749);
nand UO_2708 (O_2708,N_19622,N_19063);
and UO_2709 (O_2709,N_23312,N_21443);
or UO_2710 (O_2710,N_19675,N_22043);
and UO_2711 (O_2711,N_22462,N_21499);
and UO_2712 (O_2712,N_22589,N_21323);
or UO_2713 (O_2713,N_20231,N_20645);
and UO_2714 (O_2714,N_22326,N_19105);
nand UO_2715 (O_2715,N_19284,N_24946);
and UO_2716 (O_2716,N_21778,N_21084);
and UO_2717 (O_2717,N_20044,N_22094);
nor UO_2718 (O_2718,N_22300,N_19402);
or UO_2719 (O_2719,N_20337,N_18786);
and UO_2720 (O_2720,N_23246,N_20933);
nor UO_2721 (O_2721,N_23648,N_22336);
nor UO_2722 (O_2722,N_23219,N_21695);
and UO_2723 (O_2723,N_19010,N_18877);
nor UO_2724 (O_2724,N_19182,N_19980);
nor UO_2725 (O_2725,N_19844,N_20774);
and UO_2726 (O_2726,N_22793,N_20707);
nor UO_2727 (O_2727,N_24502,N_19834);
and UO_2728 (O_2728,N_22561,N_24901);
xnor UO_2729 (O_2729,N_20915,N_24246);
and UO_2730 (O_2730,N_24728,N_20568);
or UO_2731 (O_2731,N_24529,N_24590);
and UO_2732 (O_2732,N_23373,N_24954);
xnor UO_2733 (O_2733,N_21125,N_20287);
nor UO_2734 (O_2734,N_21602,N_20488);
nand UO_2735 (O_2735,N_24339,N_20233);
and UO_2736 (O_2736,N_19201,N_24342);
or UO_2737 (O_2737,N_24182,N_20591);
and UO_2738 (O_2738,N_21175,N_20493);
nand UO_2739 (O_2739,N_24237,N_22128);
and UO_2740 (O_2740,N_22337,N_20686);
xor UO_2741 (O_2741,N_22044,N_19845);
nor UO_2742 (O_2742,N_19523,N_24212);
or UO_2743 (O_2743,N_19341,N_21658);
nand UO_2744 (O_2744,N_19812,N_21836);
nand UO_2745 (O_2745,N_21993,N_22745);
xor UO_2746 (O_2746,N_21662,N_21964);
nor UO_2747 (O_2747,N_21009,N_19538);
xor UO_2748 (O_2748,N_22519,N_21085);
nor UO_2749 (O_2749,N_18804,N_21500);
and UO_2750 (O_2750,N_22503,N_20201);
nand UO_2751 (O_2751,N_19064,N_23591);
and UO_2752 (O_2752,N_19594,N_20495);
xnor UO_2753 (O_2753,N_19042,N_22551);
and UO_2754 (O_2754,N_23916,N_19714);
nor UO_2755 (O_2755,N_22776,N_22125);
nand UO_2756 (O_2756,N_23612,N_21851);
and UO_2757 (O_2757,N_19180,N_20632);
and UO_2758 (O_2758,N_23671,N_24014);
nand UO_2759 (O_2759,N_20967,N_22698);
xnor UO_2760 (O_2760,N_24279,N_19125);
xnor UO_2761 (O_2761,N_21457,N_21209);
and UO_2762 (O_2762,N_23406,N_19130);
nand UO_2763 (O_2763,N_22489,N_20065);
nand UO_2764 (O_2764,N_21077,N_21705);
nand UO_2765 (O_2765,N_20143,N_19447);
xnor UO_2766 (O_2766,N_18788,N_24795);
xor UO_2767 (O_2767,N_22085,N_20113);
xnor UO_2768 (O_2768,N_22127,N_19488);
xor UO_2769 (O_2769,N_23870,N_19749);
and UO_2770 (O_2770,N_22475,N_21847);
or UO_2771 (O_2771,N_20997,N_23578);
xnor UO_2772 (O_2772,N_22461,N_21519);
xnor UO_2773 (O_2773,N_19252,N_23750);
nor UO_2774 (O_2774,N_19536,N_22915);
xnor UO_2775 (O_2775,N_24090,N_19229);
or UO_2776 (O_2776,N_23502,N_23051);
and UO_2777 (O_2777,N_19745,N_22562);
nand UO_2778 (O_2778,N_23738,N_21411);
or UO_2779 (O_2779,N_21239,N_20742);
nand UO_2780 (O_2780,N_22722,N_24873);
or UO_2781 (O_2781,N_23488,N_21627);
and UO_2782 (O_2782,N_21159,N_20971);
nand UO_2783 (O_2783,N_20765,N_21934);
nor UO_2784 (O_2784,N_21385,N_24543);
xor UO_2785 (O_2785,N_21165,N_24358);
and UO_2786 (O_2786,N_23693,N_20312);
and UO_2787 (O_2787,N_21666,N_21909);
xnor UO_2788 (O_2788,N_22823,N_21156);
or UO_2789 (O_2789,N_24335,N_21057);
nor UO_2790 (O_2790,N_19608,N_21606);
and UO_2791 (O_2791,N_24792,N_22205);
xor UO_2792 (O_2792,N_23013,N_22939);
or UO_2793 (O_2793,N_22197,N_22435);
nand UO_2794 (O_2794,N_24204,N_23965);
nand UO_2795 (O_2795,N_24582,N_20766);
and UO_2796 (O_2796,N_21364,N_22400);
and UO_2797 (O_2797,N_24459,N_21983);
and UO_2798 (O_2798,N_18862,N_20273);
nand UO_2799 (O_2799,N_23607,N_19802);
xor UO_2800 (O_2800,N_20397,N_21746);
nor UO_2801 (O_2801,N_21406,N_21982);
or UO_2802 (O_2802,N_21597,N_24717);
nand UO_2803 (O_2803,N_23114,N_24702);
xor UO_2804 (O_2804,N_20871,N_21929);
nor UO_2805 (O_2805,N_22147,N_19922);
nor UO_2806 (O_2806,N_19723,N_23482);
nand UO_2807 (O_2807,N_23994,N_21355);
and UO_2808 (O_2808,N_19514,N_22500);
nand UO_2809 (O_2809,N_22389,N_23191);
nor UO_2810 (O_2810,N_24780,N_24813);
xor UO_2811 (O_2811,N_21874,N_20402);
nor UO_2812 (O_2812,N_20834,N_22544);
and UO_2813 (O_2813,N_19235,N_21536);
and UO_2814 (O_2814,N_19988,N_20614);
or UO_2815 (O_2815,N_23535,N_23204);
and UO_2816 (O_2816,N_19120,N_21708);
xnor UO_2817 (O_2817,N_20931,N_19483);
nor UO_2818 (O_2818,N_23122,N_20395);
nor UO_2819 (O_2819,N_18853,N_19717);
nand UO_2820 (O_2820,N_21247,N_21167);
and UO_2821 (O_2821,N_22634,N_22464);
nor UO_2822 (O_2822,N_24124,N_21380);
and UO_2823 (O_2823,N_24485,N_18914);
xnor UO_2824 (O_2824,N_20830,N_22694);
nor UO_2825 (O_2825,N_22948,N_19478);
nor UO_2826 (O_2826,N_22615,N_23056);
nor UO_2827 (O_2827,N_23708,N_20323);
and UO_2828 (O_2828,N_21032,N_22066);
nand UO_2829 (O_2829,N_19892,N_20812);
nand UO_2830 (O_2830,N_22284,N_22651);
or UO_2831 (O_2831,N_21811,N_24606);
nand UO_2832 (O_2832,N_21040,N_24248);
nor UO_2833 (O_2833,N_24635,N_22822);
nand UO_2834 (O_2834,N_21466,N_20796);
nor UO_2835 (O_2835,N_19725,N_22924);
nor UO_2836 (O_2836,N_20426,N_22744);
nor UO_2837 (O_2837,N_18785,N_21545);
xor UO_2838 (O_2838,N_24553,N_21496);
xor UO_2839 (O_2839,N_20346,N_24149);
or UO_2840 (O_2840,N_18768,N_23235);
xnor UO_2841 (O_2841,N_23974,N_23228);
and UO_2842 (O_2842,N_19733,N_23999);
nand UO_2843 (O_2843,N_20576,N_23956);
and UO_2844 (O_2844,N_22889,N_20033);
nor UO_2845 (O_2845,N_22448,N_23206);
or UO_2846 (O_2846,N_22526,N_19197);
nand UO_2847 (O_2847,N_23043,N_20125);
and UO_2848 (O_2848,N_23789,N_20570);
nand UO_2849 (O_2849,N_23119,N_23450);
nand UO_2850 (O_2850,N_22848,N_22936);
and UO_2851 (O_2851,N_21767,N_22818);
and UO_2852 (O_2852,N_19746,N_19656);
and UO_2853 (O_2853,N_19899,N_23161);
xnor UO_2854 (O_2854,N_21757,N_21460);
nand UO_2855 (O_2855,N_24840,N_24086);
or UO_2856 (O_2856,N_20204,N_21600);
or UO_2857 (O_2857,N_20375,N_22232);
and UO_2858 (O_2858,N_19337,N_20052);
nor UO_2859 (O_2859,N_22427,N_23366);
and UO_2860 (O_2860,N_20329,N_21023);
or UO_2861 (O_2861,N_21196,N_22905);
or UO_2862 (O_2862,N_24713,N_24860);
nand UO_2863 (O_2863,N_21942,N_20135);
xor UO_2864 (O_2864,N_22287,N_20367);
nand UO_2865 (O_2865,N_19248,N_23523);
or UO_2866 (O_2866,N_19400,N_23452);
and UO_2867 (O_2867,N_20024,N_22373);
nand UO_2868 (O_2868,N_24189,N_21678);
nor UO_2869 (O_2869,N_22803,N_22460);
xor UO_2870 (O_2870,N_22666,N_22917);
xor UO_2871 (O_2871,N_24046,N_23757);
or UO_2872 (O_2872,N_21066,N_24201);
nand UO_2873 (O_2873,N_23842,N_18857);
xnor UO_2874 (O_2874,N_23995,N_19001);
and UO_2875 (O_2875,N_22512,N_24683);
or UO_2876 (O_2876,N_23412,N_21351);
or UO_2877 (O_2877,N_24872,N_21844);
or UO_2878 (O_2878,N_19088,N_20509);
xor UO_2879 (O_2879,N_22996,N_18925);
or UO_2880 (O_2880,N_21673,N_22916);
and UO_2881 (O_2881,N_20486,N_22108);
or UO_2882 (O_2882,N_23702,N_22398);
and UO_2883 (O_2883,N_19761,N_21730);
nor UO_2884 (O_2884,N_20843,N_22680);
nor UO_2885 (O_2885,N_23080,N_22175);
nand UO_2886 (O_2886,N_24979,N_24892);
nand UO_2887 (O_2887,N_21634,N_19825);
and UO_2888 (O_2888,N_21477,N_19971);
xor UO_2889 (O_2889,N_20762,N_21880);
xnor UO_2890 (O_2890,N_20523,N_21797);
xnor UO_2891 (O_2891,N_22202,N_22189);
nand UO_2892 (O_2892,N_24343,N_22377);
or UO_2893 (O_2893,N_19439,N_24224);
nand UO_2894 (O_2894,N_24233,N_21265);
xnor UO_2895 (O_2895,N_23263,N_20118);
or UO_2896 (O_2896,N_21235,N_21119);
xnor UO_2897 (O_2897,N_23342,N_21999);
nand UO_2898 (O_2898,N_23430,N_20202);
xor UO_2899 (O_2899,N_22740,N_19752);
nor UO_2900 (O_2900,N_21227,N_18888);
xnor UO_2901 (O_2901,N_20324,N_23222);
nand UO_2902 (O_2902,N_24460,N_20891);
or UO_2903 (O_2903,N_23105,N_21573);
xnor UO_2904 (O_2904,N_19444,N_21686);
nand UO_2905 (O_2905,N_23506,N_23968);
and UO_2906 (O_2906,N_21488,N_19117);
and UO_2907 (O_2907,N_19422,N_21195);
nor UO_2908 (O_2908,N_23674,N_22294);
nand UO_2909 (O_2909,N_23310,N_22244);
or UO_2910 (O_2910,N_24344,N_21587);
and UO_2911 (O_2911,N_19058,N_23058);
nand UO_2912 (O_2912,N_23537,N_20563);
nand UO_2913 (O_2913,N_22302,N_19198);
xor UO_2914 (O_2914,N_23201,N_24512);
nor UO_2915 (O_2915,N_22019,N_20637);
or UO_2916 (O_2916,N_21622,N_21305);
nand UO_2917 (O_2917,N_19639,N_19231);
nand UO_2918 (O_2918,N_23762,N_22583);
or UO_2919 (O_2919,N_21715,N_23584);
nand UO_2920 (O_2920,N_24585,N_23520);
nor UO_2921 (O_2921,N_24510,N_18922);
and UO_2922 (O_2922,N_21473,N_22538);
nand UO_2923 (O_2923,N_21685,N_20010);
xor UO_2924 (O_2924,N_22922,N_20663);
and UO_2925 (O_2925,N_21672,N_24107);
xnor UO_2926 (O_2926,N_24509,N_23868);
nand UO_2927 (O_2927,N_24612,N_21992);
or UO_2928 (O_2928,N_24141,N_24200);
and UO_2929 (O_2929,N_20538,N_22951);
or UO_2930 (O_2930,N_23290,N_21390);
nor UO_2931 (O_2931,N_21407,N_20504);
nand UO_2932 (O_2932,N_24465,N_23836);
nand UO_2933 (O_2933,N_22201,N_24594);
or UO_2934 (O_2934,N_19530,N_18935);
or UO_2935 (O_2935,N_24262,N_22322);
nor UO_2936 (O_2936,N_22967,N_21926);
nand UO_2937 (O_2937,N_22842,N_21129);
nand UO_2938 (O_2938,N_21100,N_24956);
and UO_2939 (O_2939,N_19178,N_22488);
and UO_2940 (O_2940,N_20466,N_24138);
nand UO_2941 (O_2941,N_24720,N_21454);
nand UO_2942 (O_2942,N_22706,N_21144);
or UO_2943 (O_2943,N_24471,N_19710);
or UO_2944 (O_2944,N_24698,N_19869);
nor UO_2945 (O_2945,N_20373,N_22241);
nand UO_2946 (O_2946,N_21464,N_22409);
nor UO_2947 (O_2947,N_24093,N_20378);
xor UO_2948 (O_2948,N_23087,N_22430);
and UO_2949 (O_2949,N_20188,N_23476);
or UO_2950 (O_2950,N_19242,N_19734);
nor UO_2951 (O_2951,N_21510,N_19808);
nand UO_2952 (O_2952,N_24511,N_24015);
or UO_2953 (O_2953,N_20377,N_23519);
or UO_2954 (O_2954,N_21269,N_19258);
or UO_2955 (O_2955,N_19277,N_19497);
or UO_2956 (O_2956,N_23076,N_20002);
xnor UO_2957 (O_2957,N_22182,N_22868);
and UO_2958 (O_2958,N_20096,N_19381);
nand UO_2959 (O_2959,N_18855,N_22701);
and UO_2960 (O_2960,N_20261,N_21709);
or UO_2961 (O_2961,N_23491,N_20144);
nor UO_2962 (O_2962,N_20111,N_21056);
nor UO_2963 (O_2963,N_21528,N_19545);
or UO_2964 (O_2964,N_21892,N_23772);
nor UO_2965 (O_2965,N_20670,N_20920);
nor UO_2966 (O_2966,N_19789,N_19903);
or UO_2967 (O_2967,N_20651,N_19602);
and UO_2968 (O_2968,N_19629,N_20748);
and UO_2969 (O_2969,N_22865,N_19247);
and UO_2970 (O_2970,N_21613,N_24166);
or UO_2971 (O_2971,N_24567,N_21509);
and UO_2972 (O_2972,N_24627,N_19100);
nand UO_2973 (O_2973,N_19773,N_19521);
nor UO_2974 (O_2974,N_19850,N_21632);
xor UO_2975 (O_2975,N_18986,N_23036);
or UO_2976 (O_2976,N_20207,N_24588);
or UO_2977 (O_2977,N_22626,N_24057);
nand UO_2978 (O_2978,N_20300,N_22534);
xor UO_2979 (O_2979,N_24349,N_19660);
and UO_2980 (O_2980,N_23716,N_24825);
nand UO_2981 (O_2981,N_23969,N_21428);
nand UO_2982 (O_2982,N_22119,N_22986);
and UO_2983 (O_2983,N_19950,N_21128);
nor UO_2984 (O_2984,N_24703,N_24113);
xnor UO_2985 (O_2985,N_20136,N_18970);
nor UO_2986 (O_2986,N_22608,N_18982);
nor UO_2987 (O_2987,N_24807,N_21823);
or UO_2988 (O_2988,N_20827,N_22662);
xor UO_2989 (O_2989,N_20514,N_23071);
nor UO_2990 (O_2990,N_23567,N_23319);
xnor UO_2991 (O_2991,N_23796,N_18992);
nor UO_2992 (O_2992,N_19880,N_20034);
nand UO_2993 (O_2993,N_21671,N_24944);
nor UO_2994 (O_2994,N_19854,N_20086);
and UO_2995 (O_2995,N_22575,N_24879);
or UO_2996 (O_2996,N_21287,N_23168);
nor UO_2997 (O_2997,N_21515,N_23061);
nor UO_2998 (O_2998,N_22998,N_18819);
and UO_2999 (O_2999,N_20882,N_24712);
endmodule