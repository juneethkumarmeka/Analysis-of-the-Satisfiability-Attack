module basic_500_3000_500_4_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_488,In_121);
nand U1 (N_1,In_169,In_325);
or U2 (N_2,In_25,In_156);
nor U3 (N_3,In_129,In_238);
or U4 (N_4,In_187,In_143);
nand U5 (N_5,In_321,In_343);
or U6 (N_6,In_80,In_46);
nor U7 (N_7,In_190,In_381);
nand U8 (N_8,In_105,In_295);
nand U9 (N_9,In_222,In_8);
and U10 (N_10,In_366,In_140);
and U11 (N_11,In_342,In_130);
nand U12 (N_12,In_337,In_82);
or U13 (N_13,In_123,In_193);
nand U14 (N_14,In_77,In_76);
and U15 (N_15,In_47,In_252);
nand U16 (N_16,In_137,In_67);
nand U17 (N_17,In_410,In_29);
nor U18 (N_18,In_91,In_486);
nand U19 (N_19,In_172,In_469);
and U20 (N_20,In_346,In_303);
or U21 (N_21,In_332,In_145);
nand U22 (N_22,In_429,In_306);
nand U23 (N_23,In_18,In_63);
nand U24 (N_24,In_377,In_356);
nand U25 (N_25,In_363,In_95);
nor U26 (N_26,In_480,In_307);
or U27 (N_27,In_414,In_4);
nor U28 (N_28,In_92,In_371);
and U29 (N_29,In_352,In_225);
or U30 (N_30,In_370,In_173);
nand U31 (N_31,In_39,In_289);
nand U32 (N_32,In_440,In_167);
and U33 (N_33,In_28,In_24);
nand U34 (N_34,In_115,In_174);
nor U35 (N_35,In_208,In_90);
nor U36 (N_36,In_402,In_361);
or U37 (N_37,In_396,In_400);
and U38 (N_38,In_58,In_125);
nand U39 (N_39,In_186,In_434);
or U40 (N_40,In_360,In_498);
and U41 (N_41,In_312,In_481);
or U42 (N_42,In_443,In_375);
and U43 (N_43,In_459,In_170);
and U44 (N_44,In_326,In_231);
nor U45 (N_45,In_13,In_280);
or U46 (N_46,In_255,In_73);
nor U47 (N_47,In_185,In_53);
nand U48 (N_48,In_59,In_286);
xor U49 (N_49,In_355,In_165);
nor U50 (N_50,In_250,In_86);
or U51 (N_51,In_97,In_249);
nor U52 (N_52,In_499,In_229);
nor U53 (N_53,In_308,In_446);
or U54 (N_54,In_248,In_142);
and U55 (N_55,In_38,In_221);
and U56 (N_56,In_344,In_114);
and U57 (N_57,In_52,In_495);
xor U58 (N_58,In_405,In_292);
and U59 (N_59,In_372,In_262);
or U60 (N_60,In_196,In_61);
or U61 (N_61,In_263,In_107);
nand U62 (N_62,In_171,In_69);
and U63 (N_63,In_224,In_1);
nand U64 (N_64,In_180,In_94);
or U65 (N_65,In_37,In_198);
or U66 (N_66,In_78,In_467);
and U67 (N_67,In_23,In_425);
nand U68 (N_68,In_132,In_213);
or U69 (N_69,In_124,In_436);
or U70 (N_70,In_181,In_462);
nor U71 (N_71,In_113,In_475);
nand U72 (N_72,In_157,In_182);
and U73 (N_73,In_484,In_333);
or U74 (N_74,In_444,In_164);
or U75 (N_75,In_272,In_409);
or U76 (N_76,In_463,In_12);
or U77 (N_77,In_168,In_7);
and U78 (N_78,In_100,In_131);
or U79 (N_79,In_179,In_406);
and U80 (N_80,In_454,In_240);
and U81 (N_81,In_88,In_184);
nor U82 (N_82,In_258,In_228);
nand U83 (N_83,In_83,In_247);
nand U84 (N_84,In_387,In_87);
or U85 (N_85,In_353,In_296);
and U86 (N_86,In_2,In_139);
nand U87 (N_87,In_192,In_122);
nand U88 (N_88,In_5,In_141);
and U89 (N_89,In_188,In_49);
nor U90 (N_90,In_146,In_389);
nand U91 (N_91,In_232,In_220);
and U92 (N_92,In_259,In_70);
and U93 (N_93,In_490,In_93);
or U94 (N_94,In_417,In_199);
nor U95 (N_95,In_471,In_494);
or U96 (N_96,In_383,In_104);
nor U97 (N_97,In_176,In_466);
or U98 (N_98,In_393,In_474);
nor U99 (N_99,In_233,In_230);
and U100 (N_100,In_470,In_430);
nor U101 (N_101,In_17,In_246);
and U102 (N_102,In_278,In_281);
nand U103 (N_103,In_439,In_210);
and U104 (N_104,In_20,In_460);
or U105 (N_105,In_437,In_345);
nand U106 (N_106,In_461,In_398);
and U107 (N_107,In_253,In_98);
and U108 (N_108,In_66,In_21);
and U109 (N_109,In_215,In_458);
and U110 (N_110,In_265,In_314);
nor U111 (N_111,In_261,In_364);
nor U112 (N_112,In_223,In_476);
nand U113 (N_113,In_413,In_403);
or U114 (N_114,In_111,In_497);
nor U115 (N_115,In_424,In_448);
or U116 (N_116,In_19,In_478);
nor U117 (N_117,In_160,In_175);
nand U118 (N_118,In_154,In_420);
nor U119 (N_119,In_34,In_358);
nand U120 (N_120,In_316,In_482);
and U121 (N_121,In_84,In_242);
nand U122 (N_122,In_9,In_43);
or U123 (N_123,In_136,In_309);
and U124 (N_124,In_384,In_149);
or U125 (N_125,In_219,In_178);
nor U126 (N_126,In_71,In_218);
and U127 (N_127,In_202,In_365);
nor U128 (N_128,In_291,In_10);
or U129 (N_129,In_338,In_26);
nand U130 (N_130,In_112,In_269);
or U131 (N_131,In_340,In_305);
or U132 (N_132,In_323,In_45);
or U133 (N_133,In_422,In_382);
or U134 (N_134,In_464,In_85);
nand U135 (N_135,In_334,In_260);
and U136 (N_136,In_27,In_126);
or U137 (N_137,In_290,In_216);
and U138 (N_138,In_110,In_177);
or U139 (N_139,In_450,In_395);
and U140 (N_140,In_391,In_330);
and U141 (N_141,In_133,In_319);
or U142 (N_142,In_11,In_419);
nor U143 (N_143,In_407,In_380);
xor U144 (N_144,In_431,In_89);
nor U145 (N_145,In_99,In_270);
nand U146 (N_146,In_282,In_349);
and U147 (N_147,In_206,In_368);
and U148 (N_148,In_150,In_264);
nand U149 (N_149,In_339,In_350);
and U150 (N_150,In_3,In_376);
xor U151 (N_151,In_204,In_418);
nor U152 (N_152,In_435,In_159);
nand U153 (N_153,In_135,In_217);
and U154 (N_154,In_166,In_60);
or U155 (N_155,In_211,In_318);
and U156 (N_156,In_310,In_268);
or U157 (N_157,In_447,In_254);
and U158 (N_158,In_416,In_277);
or U159 (N_159,In_485,In_279);
or U160 (N_160,In_134,In_108);
and U161 (N_161,In_492,In_191);
nor U162 (N_162,In_283,In_327);
and U163 (N_163,In_341,In_120);
nand U164 (N_164,In_144,In_465);
and U165 (N_165,In_235,In_241);
or U166 (N_166,In_412,In_385);
nand U167 (N_167,In_234,In_449);
and U168 (N_168,In_392,In_496);
nand U169 (N_169,In_62,In_489);
and U170 (N_170,In_452,In_36);
or U171 (N_171,In_151,In_483);
and U172 (N_172,In_399,In_74);
nor U173 (N_173,In_251,In_32);
or U174 (N_174,In_72,In_479);
or U175 (N_175,In_294,In_347);
or U176 (N_176,In_455,In_293);
or U177 (N_177,In_138,In_408);
and U178 (N_178,In_109,In_390);
or U179 (N_179,In_359,In_96);
and U180 (N_180,In_378,In_31);
and U181 (N_181,In_456,In_423);
nor U182 (N_182,In_68,In_183);
and U183 (N_183,In_275,In_54);
or U184 (N_184,In_304,In_298);
nor U185 (N_185,In_51,In_106);
nand U186 (N_186,In_212,In_427);
nand U187 (N_187,In_320,In_55);
and U188 (N_188,In_276,In_155);
and U189 (N_189,In_153,In_16);
or U190 (N_190,In_297,In_64);
and U191 (N_191,In_14,In_421);
or U192 (N_192,In_491,In_236);
nand U193 (N_193,In_267,In_301);
nor U194 (N_194,In_493,In_324);
nand U195 (N_195,In_311,In_40);
or U196 (N_196,In_243,In_33);
or U197 (N_197,In_457,In_237);
and U198 (N_198,In_101,In_57);
and U199 (N_199,In_411,In_453);
or U200 (N_200,In_300,In_487);
nor U201 (N_201,In_473,In_103);
or U202 (N_202,In_207,In_79);
and U203 (N_203,In_257,In_317);
and U204 (N_204,In_335,In_328);
nor U205 (N_205,In_362,In_438);
or U206 (N_206,In_441,In_41);
and U207 (N_207,In_200,In_329);
or U208 (N_208,In_245,In_432);
nor U209 (N_209,In_472,In_256);
and U210 (N_210,In_147,In_285);
or U211 (N_211,In_6,In_374);
nand U212 (N_212,In_117,In_428);
nand U213 (N_213,In_394,In_477);
nand U214 (N_214,In_152,In_426);
or U215 (N_215,In_48,In_22);
nor U216 (N_216,In_161,In_373);
and U217 (N_217,In_433,In_442);
and U218 (N_218,In_336,In_331);
nor U219 (N_219,In_401,In_201);
nor U220 (N_220,In_205,In_367);
nor U221 (N_221,In_386,In_30);
or U222 (N_222,In_445,In_351);
or U223 (N_223,In_379,In_128);
nand U224 (N_224,In_163,In_119);
nor U225 (N_225,In_209,In_451);
nor U226 (N_226,In_322,In_197);
nor U227 (N_227,In_288,In_65);
or U228 (N_228,In_227,In_189);
nor U229 (N_229,In_302,In_15);
nor U230 (N_230,In_75,In_195);
or U231 (N_231,In_203,In_287);
nor U232 (N_232,In_273,In_194);
nand U233 (N_233,In_274,In_404);
or U234 (N_234,In_35,In_239);
nor U235 (N_235,In_397,In_369);
nand U236 (N_236,In_468,In_388);
nor U237 (N_237,In_271,In_56);
or U238 (N_238,In_162,In_0);
or U239 (N_239,In_158,In_354);
or U240 (N_240,In_226,In_313);
or U241 (N_241,In_127,In_116);
nor U242 (N_242,In_44,In_284);
nor U243 (N_243,In_357,In_42);
nand U244 (N_244,In_148,In_348);
and U245 (N_245,In_118,In_315);
or U246 (N_246,In_299,In_266);
nand U247 (N_247,In_214,In_102);
and U248 (N_248,In_415,In_81);
and U249 (N_249,In_50,In_244);
and U250 (N_250,In_471,In_484);
and U251 (N_251,In_125,In_2);
and U252 (N_252,In_321,In_476);
nor U253 (N_253,In_299,In_41);
nand U254 (N_254,In_241,In_31);
and U255 (N_255,In_64,In_264);
nand U256 (N_256,In_134,In_302);
nor U257 (N_257,In_305,In_150);
xor U258 (N_258,In_219,In_56);
nand U259 (N_259,In_154,In_31);
or U260 (N_260,In_403,In_465);
nor U261 (N_261,In_274,In_54);
xor U262 (N_262,In_110,In_435);
or U263 (N_263,In_437,In_176);
nand U264 (N_264,In_410,In_316);
or U265 (N_265,In_444,In_438);
or U266 (N_266,In_373,In_471);
nor U267 (N_267,In_250,In_283);
nor U268 (N_268,In_446,In_327);
nand U269 (N_269,In_400,In_344);
and U270 (N_270,In_228,In_115);
nor U271 (N_271,In_396,In_381);
nand U272 (N_272,In_242,In_48);
nand U273 (N_273,In_94,In_370);
nor U274 (N_274,In_103,In_201);
or U275 (N_275,In_78,In_496);
nor U276 (N_276,In_70,In_361);
nor U277 (N_277,In_23,In_236);
and U278 (N_278,In_426,In_284);
and U279 (N_279,In_81,In_347);
nand U280 (N_280,In_230,In_184);
nand U281 (N_281,In_14,In_349);
nand U282 (N_282,In_247,In_285);
and U283 (N_283,In_429,In_466);
nor U284 (N_284,In_189,In_129);
and U285 (N_285,In_169,In_375);
or U286 (N_286,In_21,In_210);
or U287 (N_287,In_265,In_215);
nor U288 (N_288,In_382,In_387);
and U289 (N_289,In_376,In_253);
and U290 (N_290,In_127,In_297);
or U291 (N_291,In_156,In_229);
or U292 (N_292,In_94,In_420);
nor U293 (N_293,In_422,In_380);
nor U294 (N_294,In_35,In_364);
nand U295 (N_295,In_439,In_402);
and U296 (N_296,In_37,In_178);
or U297 (N_297,In_400,In_207);
or U298 (N_298,In_116,In_477);
and U299 (N_299,In_253,In_374);
nor U300 (N_300,In_205,In_397);
and U301 (N_301,In_172,In_240);
nand U302 (N_302,In_200,In_330);
and U303 (N_303,In_442,In_167);
and U304 (N_304,In_485,In_184);
or U305 (N_305,In_121,In_176);
or U306 (N_306,In_138,In_35);
and U307 (N_307,In_347,In_175);
nor U308 (N_308,In_102,In_496);
nor U309 (N_309,In_220,In_150);
or U310 (N_310,In_75,In_370);
and U311 (N_311,In_165,In_447);
and U312 (N_312,In_312,In_397);
nand U313 (N_313,In_190,In_82);
nand U314 (N_314,In_181,In_342);
nor U315 (N_315,In_22,In_333);
or U316 (N_316,In_111,In_211);
nand U317 (N_317,In_383,In_442);
nand U318 (N_318,In_291,In_454);
and U319 (N_319,In_358,In_422);
and U320 (N_320,In_76,In_270);
nand U321 (N_321,In_93,In_411);
nor U322 (N_322,In_121,In_295);
nor U323 (N_323,In_293,In_92);
nor U324 (N_324,In_192,In_38);
or U325 (N_325,In_250,In_111);
nor U326 (N_326,In_337,In_493);
and U327 (N_327,In_95,In_16);
or U328 (N_328,In_287,In_12);
or U329 (N_329,In_458,In_113);
or U330 (N_330,In_425,In_410);
and U331 (N_331,In_160,In_372);
nand U332 (N_332,In_485,In_395);
nand U333 (N_333,In_453,In_288);
and U334 (N_334,In_350,In_299);
nand U335 (N_335,In_444,In_206);
nand U336 (N_336,In_125,In_199);
nand U337 (N_337,In_116,In_498);
or U338 (N_338,In_63,In_369);
or U339 (N_339,In_154,In_367);
nand U340 (N_340,In_279,In_224);
and U341 (N_341,In_325,In_432);
or U342 (N_342,In_144,In_470);
and U343 (N_343,In_119,In_228);
or U344 (N_344,In_165,In_47);
and U345 (N_345,In_184,In_477);
nor U346 (N_346,In_13,In_60);
or U347 (N_347,In_145,In_403);
nor U348 (N_348,In_26,In_349);
nand U349 (N_349,In_465,In_463);
and U350 (N_350,In_445,In_89);
and U351 (N_351,In_386,In_225);
nor U352 (N_352,In_417,In_432);
or U353 (N_353,In_111,In_53);
or U354 (N_354,In_172,In_115);
nor U355 (N_355,In_246,In_188);
nor U356 (N_356,In_160,In_453);
nor U357 (N_357,In_410,In_186);
nand U358 (N_358,In_86,In_55);
or U359 (N_359,In_317,In_226);
or U360 (N_360,In_92,In_107);
nand U361 (N_361,In_287,In_322);
and U362 (N_362,In_211,In_200);
and U363 (N_363,In_95,In_280);
or U364 (N_364,In_441,In_57);
or U365 (N_365,In_72,In_386);
nand U366 (N_366,In_235,In_211);
or U367 (N_367,In_122,In_252);
and U368 (N_368,In_290,In_31);
or U369 (N_369,In_232,In_471);
or U370 (N_370,In_128,In_33);
nand U371 (N_371,In_103,In_209);
nor U372 (N_372,In_258,In_289);
or U373 (N_373,In_12,In_382);
or U374 (N_374,In_261,In_191);
nand U375 (N_375,In_130,In_168);
or U376 (N_376,In_480,In_17);
and U377 (N_377,In_131,In_122);
or U378 (N_378,In_470,In_104);
and U379 (N_379,In_332,In_4);
or U380 (N_380,In_215,In_461);
nand U381 (N_381,In_358,In_175);
and U382 (N_382,In_171,In_354);
nand U383 (N_383,In_475,In_437);
or U384 (N_384,In_28,In_55);
nor U385 (N_385,In_148,In_306);
nor U386 (N_386,In_146,In_128);
nor U387 (N_387,In_22,In_89);
and U388 (N_388,In_48,In_404);
nor U389 (N_389,In_444,In_218);
nand U390 (N_390,In_82,In_51);
nor U391 (N_391,In_283,In_102);
and U392 (N_392,In_139,In_119);
or U393 (N_393,In_490,In_41);
or U394 (N_394,In_203,In_189);
nand U395 (N_395,In_454,In_118);
nor U396 (N_396,In_315,In_26);
nand U397 (N_397,In_407,In_302);
or U398 (N_398,In_28,In_161);
nand U399 (N_399,In_350,In_244);
nor U400 (N_400,In_68,In_175);
nor U401 (N_401,In_476,In_14);
nand U402 (N_402,In_149,In_251);
nand U403 (N_403,In_195,In_133);
and U404 (N_404,In_338,In_44);
or U405 (N_405,In_204,In_427);
nor U406 (N_406,In_85,In_194);
and U407 (N_407,In_60,In_224);
nand U408 (N_408,In_401,In_386);
and U409 (N_409,In_199,In_105);
and U410 (N_410,In_179,In_226);
and U411 (N_411,In_68,In_11);
nand U412 (N_412,In_478,In_73);
and U413 (N_413,In_479,In_114);
and U414 (N_414,In_198,In_393);
or U415 (N_415,In_409,In_369);
nor U416 (N_416,In_496,In_379);
and U417 (N_417,In_191,In_189);
nor U418 (N_418,In_288,In_352);
and U419 (N_419,In_208,In_216);
or U420 (N_420,In_468,In_106);
nor U421 (N_421,In_108,In_150);
or U422 (N_422,In_345,In_26);
and U423 (N_423,In_110,In_211);
or U424 (N_424,In_369,In_331);
nand U425 (N_425,In_288,In_267);
nor U426 (N_426,In_384,In_365);
nand U427 (N_427,In_76,In_160);
and U428 (N_428,In_468,In_481);
nand U429 (N_429,In_34,In_174);
or U430 (N_430,In_411,In_122);
and U431 (N_431,In_137,In_169);
or U432 (N_432,In_208,In_286);
nor U433 (N_433,In_190,In_199);
nor U434 (N_434,In_38,In_417);
nand U435 (N_435,In_52,In_83);
or U436 (N_436,In_479,In_239);
nor U437 (N_437,In_380,In_480);
nor U438 (N_438,In_133,In_91);
or U439 (N_439,In_361,In_160);
nand U440 (N_440,In_76,In_17);
or U441 (N_441,In_374,In_454);
nor U442 (N_442,In_393,In_322);
nand U443 (N_443,In_280,In_119);
or U444 (N_444,In_448,In_52);
or U445 (N_445,In_67,In_367);
nand U446 (N_446,In_229,In_309);
nor U447 (N_447,In_266,In_202);
nand U448 (N_448,In_254,In_38);
nor U449 (N_449,In_342,In_173);
nor U450 (N_450,In_106,In_406);
nand U451 (N_451,In_251,In_305);
and U452 (N_452,In_421,In_141);
and U453 (N_453,In_114,In_80);
and U454 (N_454,In_209,In_114);
or U455 (N_455,In_298,In_8);
nor U456 (N_456,In_254,In_332);
and U457 (N_457,In_440,In_271);
nand U458 (N_458,In_289,In_404);
nand U459 (N_459,In_380,In_481);
nand U460 (N_460,In_70,In_323);
or U461 (N_461,In_126,In_202);
and U462 (N_462,In_16,In_397);
or U463 (N_463,In_267,In_238);
nor U464 (N_464,In_335,In_91);
nor U465 (N_465,In_9,In_427);
nand U466 (N_466,In_37,In_26);
or U467 (N_467,In_221,In_111);
nor U468 (N_468,In_184,In_52);
and U469 (N_469,In_90,In_79);
nand U470 (N_470,In_123,In_205);
and U471 (N_471,In_491,In_404);
nor U472 (N_472,In_27,In_85);
or U473 (N_473,In_46,In_367);
or U474 (N_474,In_179,In_396);
nor U475 (N_475,In_156,In_199);
and U476 (N_476,In_203,In_252);
nand U477 (N_477,In_68,In_343);
and U478 (N_478,In_323,In_173);
and U479 (N_479,In_333,In_133);
nor U480 (N_480,In_348,In_388);
or U481 (N_481,In_115,In_110);
and U482 (N_482,In_498,In_385);
nand U483 (N_483,In_171,In_178);
or U484 (N_484,In_217,In_41);
nor U485 (N_485,In_213,In_425);
and U486 (N_486,In_371,In_331);
nor U487 (N_487,In_223,In_215);
nand U488 (N_488,In_160,In_95);
nand U489 (N_489,In_453,In_174);
nand U490 (N_490,In_287,In_234);
nand U491 (N_491,In_80,In_308);
and U492 (N_492,In_26,In_108);
nor U493 (N_493,In_83,In_258);
and U494 (N_494,In_129,In_330);
or U495 (N_495,In_303,In_339);
or U496 (N_496,In_474,In_78);
or U497 (N_497,In_463,In_325);
nor U498 (N_498,In_280,In_482);
nor U499 (N_499,In_448,In_408);
or U500 (N_500,In_350,In_486);
or U501 (N_501,In_96,In_345);
nor U502 (N_502,In_350,In_259);
nor U503 (N_503,In_455,In_321);
nor U504 (N_504,In_370,In_120);
or U505 (N_505,In_369,In_9);
nand U506 (N_506,In_48,In_97);
or U507 (N_507,In_472,In_136);
or U508 (N_508,In_148,In_387);
and U509 (N_509,In_465,In_46);
nor U510 (N_510,In_88,In_275);
and U511 (N_511,In_262,In_425);
and U512 (N_512,In_144,In_238);
nand U513 (N_513,In_246,In_137);
nor U514 (N_514,In_39,In_88);
and U515 (N_515,In_247,In_121);
or U516 (N_516,In_84,In_478);
or U517 (N_517,In_17,In_107);
nor U518 (N_518,In_376,In_179);
nor U519 (N_519,In_84,In_188);
or U520 (N_520,In_438,In_473);
nor U521 (N_521,In_414,In_341);
nor U522 (N_522,In_191,In_286);
and U523 (N_523,In_447,In_406);
nand U524 (N_524,In_212,In_360);
nor U525 (N_525,In_314,In_281);
nor U526 (N_526,In_39,In_116);
nand U527 (N_527,In_455,In_357);
nor U528 (N_528,In_151,In_337);
and U529 (N_529,In_387,In_121);
and U530 (N_530,In_163,In_479);
nand U531 (N_531,In_215,In_96);
nand U532 (N_532,In_62,In_172);
or U533 (N_533,In_282,In_493);
nand U534 (N_534,In_231,In_382);
or U535 (N_535,In_188,In_110);
or U536 (N_536,In_182,In_380);
and U537 (N_537,In_335,In_413);
nand U538 (N_538,In_430,In_286);
nor U539 (N_539,In_252,In_107);
or U540 (N_540,In_497,In_48);
or U541 (N_541,In_308,In_77);
or U542 (N_542,In_307,In_344);
nor U543 (N_543,In_120,In_209);
nor U544 (N_544,In_155,In_272);
nand U545 (N_545,In_132,In_234);
and U546 (N_546,In_198,In_200);
or U547 (N_547,In_466,In_108);
nor U548 (N_548,In_312,In_284);
nand U549 (N_549,In_392,In_159);
nand U550 (N_550,In_185,In_418);
nor U551 (N_551,In_9,In_168);
nand U552 (N_552,In_480,In_329);
nand U553 (N_553,In_313,In_441);
or U554 (N_554,In_336,In_429);
and U555 (N_555,In_447,In_418);
or U556 (N_556,In_98,In_6);
nand U557 (N_557,In_383,In_403);
or U558 (N_558,In_435,In_302);
nor U559 (N_559,In_46,In_429);
or U560 (N_560,In_316,In_348);
or U561 (N_561,In_105,In_314);
nor U562 (N_562,In_338,In_234);
and U563 (N_563,In_395,In_76);
or U564 (N_564,In_471,In_12);
or U565 (N_565,In_463,In_480);
nand U566 (N_566,In_420,In_378);
nor U567 (N_567,In_438,In_13);
or U568 (N_568,In_96,In_17);
nand U569 (N_569,In_68,In_440);
and U570 (N_570,In_407,In_180);
nand U571 (N_571,In_401,In_296);
and U572 (N_572,In_203,In_231);
or U573 (N_573,In_114,In_348);
nand U574 (N_574,In_229,In_226);
and U575 (N_575,In_308,In_241);
nand U576 (N_576,In_46,In_190);
or U577 (N_577,In_147,In_201);
or U578 (N_578,In_3,In_392);
nand U579 (N_579,In_156,In_136);
or U580 (N_580,In_16,In_140);
nor U581 (N_581,In_69,In_382);
or U582 (N_582,In_354,In_229);
or U583 (N_583,In_325,In_91);
nor U584 (N_584,In_402,In_346);
nor U585 (N_585,In_429,In_71);
nand U586 (N_586,In_472,In_206);
nand U587 (N_587,In_40,In_140);
nor U588 (N_588,In_310,In_218);
or U589 (N_589,In_146,In_20);
xnor U590 (N_590,In_424,In_488);
nor U591 (N_591,In_19,In_134);
nand U592 (N_592,In_90,In_217);
or U593 (N_593,In_334,In_26);
or U594 (N_594,In_72,In_414);
or U595 (N_595,In_366,In_282);
or U596 (N_596,In_63,In_187);
nor U597 (N_597,In_179,In_105);
or U598 (N_598,In_223,In_264);
nor U599 (N_599,In_250,In_315);
and U600 (N_600,In_429,In_18);
nand U601 (N_601,In_47,In_495);
or U602 (N_602,In_346,In_1);
or U603 (N_603,In_420,In_232);
or U604 (N_604,In_496,In_267);
and U605 (N_605,In_460,In_353);
and U606 (N_606,In_398,In_4);
or U607 (N_607,In_136,In_298);
nor U608 (N_608,In_346,In_77);
and U609 (N_609,In_386,In_279);
nand U610 (N_610,In_349,In_152);
nand U611 (N_611,In_42,In_196);
nor U612 (N_612,In_329,In_308);
nor U613 (N_613,In_265,In_136);
nand U614 (N_614,In_278,In_96);
xnor U615 (N_615,In_447,In_217);
nand U616 (N_616,In_294,In_53);
or U617 (N_617,In_425,In_26);
xor U618 (N_618,In_179,In_378);
nor U619 (N_619,In_166,In_346);
and U620 (N_620,In_46,In_35);
xor U621 (N_621,In_442,In_51);
and U622 (N_622,In_430,In_267);
nand U623 (N_623,In_76,In_217);
and U624 (N_624,In_492,In_116);
nand U625 (N_625,In_211,In_462);
nor U626 (N_626,In_368,In_353);
and U627 (N_627,In_499,In_46);
or U628 (N_628,In_439,In_385);
nor U629 (N_629,In_73,In_409);
nand U630 (N_630,In_366,In_246);
or U631 (N_631,In_319,In_300);
or U632 (N_632,In_149,In_43);
nand U633 (N_633,In_403,In_134);
and U634 (N_634,In_40,In_342);
and U635 (N_635,In_127,In_362);
nand U636 (N_636,In_284,In_200);
or U637 (N_637,In_72,In_5);
or U638 (N_638,In_59,In_201);
nor U639 (N_639,In_497,In_182);
or U640 (N_640,In_330,In_236);
or U641 (N_641,In_245,In_236);
nand U642 (N_642,In_90,In_159);
or U643 (N_643,In_216,In_106);
nand U644 (N_644,In_42,In_88);
and U645 (N_645,In_247,In_289);
nor U646 (N_646,In_400,In_373);
and U647 (N_647,In_29,In_55);
or U648 (N_648,In_361,In_335);
nand U649 (N_649,In_465,In_272);
nand U650 (N_650,In_493,In_469);
nor U651 (N_651,In_437,In_324);
nand U652 (N_652,In_340,In_18);
or U653 (N_653,In_259,In_399);
nand U654 (N_654,In_53,In_171);
or U655 (N_655,In_69,In_107);
or U656 (N_656,In_4,In_361);
and U657 (N_657,In_203,In_202);
or U658 (N_658,In_465,In_285);
nand U659 (N_659,In_371,In_324);
or U660 (N_660,In_405,In_304);
nand U661 (N_661,In_11,In_58);
nand U662 (N_662,In_147,In_171);
nand U663 (N_663,In_332,In_484);
and U664 (N_664,In_28,In_316);
and U665 (N_665,In_325,In_464);
or U666 (N_666,In_139,In_168);
nand U667 (N_667,In_490,In_388);
nand U668 (N_668,In_378,In_106);
and U669 (N_669,In_338,In_239);
nand U670 (N_670,In_61,In_241);
and U671 (N_671,In_497,In_151);
nor U672 (N_672,In_171,In_345);
or U673 (N_673,In_316,In_457);
nor U674 (N_674,In_342,In_167);
nand U675 (N_675,In_431,In_41);
nand U676 (N_676,In_65,In_28);
and U677 (N_677,In_101,In_498);
nand U678 (N_678,In_482,In_492);
or U679 (N_679,In_27,In_53);
nor U680 (N_680,In_130,In_142);
nand U681 (N_681,In_188,In_264);
or U682 (N_682,In_92,In_199);
nand U683 (N_683,In_308,In_382);
nor U684 (N_684,In_102,In_247);
nand U685 (N_685,In_355,In_473);
nor U686 (N_686,In_160,In_60);
and U687 (N_687,In_152,In_116);
and U688 (N_688,In_112,In_366);
or U689 (N_689,In_376,In_37);
and U690 (N_690,In_178,In_197);
nor U691 (N_691,In_315,In_280);
and U692 (N_692,In_313,In_142);
nor U693 (N_693,In_480,In_159);
nor U694 (N_694,In_389,In_180);
nor U695 (N_695,In_463,In_193);
nand U696 (N_696,In_193,In_25);
or U697 (N_697,In_41,In_78);
nand U698 (N_698,In_387,In_79);
nor U699 (N_699,In_372,In_66);
or U700 (N_700,In_72,In_176);
nor U701 (N_701,In_462,In_465);
or U702 (N_702,In_97,In_88);
nand U703 (N_703,In_317,In_394);
nand U704 (N_704,In_22,In_360);
or U705 (N_705,In_116,In_493);
nand U706 (N_706,In_357,In_456);
nor U707 (N_707,In_293,In_83);
and U708 (N_708,In_260,In_37);
nand U709 (N_709,In_408,In_58);
and U710 (N_710,In_257,In_494);
or U711 (N_711,In_370,In_294);
nor U712 (N_712,In_31,In_230);
nor U713 (N_713,In_96,In_372);
nor U714 (N_714,In_402,In_38);
nand U715 (N_715,In_291,In_387);
or U716 (N_716,In_391,In_435);
nor U717 (N_717,In_276,In_348);
and U718 (N_718,In_237,In_144);
nor U719 (N_719,In_128,In_370);
or U720 (N_720,In_14,In_133);
and U721 (N_721,In_39,In_211);
nor U722 (N_722,In_395,In_166);
and U723 (N_723,In_364,In_318);
nand U724 (N_724,In_37,In_484);
nand U725 (N_725,In_103,In_385);
nor U726 (N_726,In_450,In_284);
and U727 (N_727,In_208,In_8);
nand U728 (N_728,In_100,In_490);
or U729 (N_729,In_36,In_330);
or U730 (N_730,In_24,In_397);
xnor U731 (N_731,In_72,In_348);
and U732 (N_732,In_260,In_163);
and U733 (N_733,In_460,In_37);
nand U734 (N_734,In_197,In_299);
nor U735 (N_735,In_250,In_176);
nor U736 (N_736,In_346,In_209);
nor U737 (N_737,In_74,In_2);
nand U738 (N_738,In_302,In_376);
and U739 (N_739,In_252,In_75);
nand U740 (N_740,In_55,In_418);
nand U741 (N_741,In_240,In_210);
nand U742 (N_742,In_344,In_54);
nand U743 (N_743,In_364,In_293);
nand U744 (N_744,In_436,In_274);
or U745 (N_745,In_442,In_5);
nor U746 (N_746,In_148,In_374);
and U747 (N_747,In_470,In_257);
nor U748 (N_748,In_473,In_481);
and U749 (N_749,In_268,In_329);
and U750 (N_750,N_587,N_480);
nand U751 (N_751,N_546,N_652);
nand U752 (N_752,N_594,N_644);
and U753 (N_753,N_54,N_595);
and U754 (N_754,N_110,N_305);
and U755 (N_755,N_465,N_673);
nor U756 (N_756,N_473,N_560);
or U757 (N_757,N_374,N_33);
or U758 (N_758,N_552,N_17);
and U759 (N_759,N_405,N_498);
nand U760 (N_760,N_212,N_703);
nor U761 (N_761,N_461,N_640);
nor U762 (N_762,N_302,N_194);
and U763 (N_763,N_271,N_419);
or U764 (N_764,N_626,N_399);
and U765 (N_765,N_157,N_295);
and U766 (N_766,N_620,N_651);
nand U767 (N_767,N_232,N_493);
and U768 (N_768,N_311,N_439);
or U769 (N_769,N_347,N_240);
nand U770 (N_770,N_579,N_230);
nor U771 (N_771,N_713,N_359);
nand U772 (N_772,N_237,N_401);
nor U773 (N_773,N_430,N_127);
and U774 (N_774,N_734,N_443);
nor U775 (N_775,N_450,N_203);
and U776 (N_776,N_60,N_691);
nand U777 (N_777,N_433,N_675);
or U778 (N_778,N_529,N_187);
nand U779 (N_779,N_446,N_61);
nand U780 (N_780,N_536,N_234);
and U781 (N_781,N_534,N_638);
nand U782 (N_782,N_109,N_325);
nand U783 (N_783,N_338,N_490);
nor U784 (N_784,N_396,N_455);
nand U785 (N_785,N_719,N_600);
and U786 (N_786,N_254,N_70);
and U787 (N_787,N_161,N_226);
nor U788 (N_788,N_133,N_126);
nand U789 (N_789,N_647,N_50);
nor U790 (N_790,N_561,N_591);
and U791 (N_791,N_417,N_721);
nor U792 (N_792,N_192,N_298);
xnor U793 (N_793,N_138,N_225);
nor U794 (N_794,N_294,N_505);
nand U795 (N_795,N_142,N_738);
xor U796 (N_796,N_603,N_467);
and U797 (N_797,N_264,N_55);
or U798 (N_798,N_684,N_735);
or U799 (N_799,N_167,N_631);
nor U800 (N_800,N_458,N_736);
nor U801 (N_801,N_181,N_261);
nor U802 (N_802,N_266,N_436);
and U803 (N_803,N_395,N_71);
nand U804 (N_804,N_674,N_14);
nand U805 (N_805,N_507,N_427);
nor U806 (N_806,N_425,N_743);
nor U807 (N_807,N_72,N_292);
or U808 (N_808,N_80,N_550);
or U809 (N_809,N_658,N_313);
nor U810 (N_810,N_376,N_654);
nand U811 (N_811,N_366,N_402);
or U812 (N_812,N_469,N_216);
nor U813 (N_813,N_680,N_285);
nor U814 (N_814,N_682,N_702);
nor U815 (N_815,N_79,N_58);
or U816 (N_816,N_189,N_362);
and U817 (N_817,N_547,N_116);
nor U818 (N_818,N_501,N_532);
nand U819 (N_819,N_13,N_643);
nand U820 (N_820,N_385,N_291);
nor U821 (N_821,N_9,N_416);
and U822 (N_822,N_340,N_179);
nand U823 (N_823,N_98,N_256);
nand U824 (N_824,N_356,N_155);
nand U825 (N_825,N_645,N_514);
and U826 (N_826,N_4,N_343);
nand U827 (N_827,N_668,N_77);
nand U828 (N_828,N_633,N_278);
nand U829 (N_829,N_479,N_213);
nand U830 (N_830,N_308,N_48);
nor U831 (N_831,N_492,N_306);
and U832 (N_832,N_732,N_500);
or U833 (N_833,N_22,N_464);
or U834 (N_834,N_460,N_342);
and U835 (N_835,N_276,N_693);
and U836 (N_836,N_391,N_201);
nor U837 (N_837,N_564,N_335);
or U838 (N_838,N_265,N_319);
or U839 (N_839,N_130,N_330);
or U840 (N_840,N_349,N_437);
or U841 (N_841,N_383,N_290);
nand U842 (N_842,N_584,N_745);
nor U843 (N_843,N_68,N_695);
nand U844 (N_844,N_169,N_5);
nand U845 (N_845,N_255,N_683);
nand U846 (N_846,N_530,N_243);
or U847 (N_847,N_44,N_105);
nor U848 (N_848,N_217,N_337);
or U849 (N_849,N_336,N_281);
nand U850 (N_850,N_678,N_456);
and U851 (N_851,N_36,N_400);
nand U852 (N_852,N_82,N_275);
or U853 (N_853,N_388,N_528);
and U854 (N_854,N_608,N_152);
nor U855 (N_855,N_519,N_568);
nand U856 (N_856,N_510,N_559);
or U857 (N_857,N_164,N_12);
or U858 (N_858,N_576,N_139);
or U859 (N_859,N_454,N_51);
and U860 (N_860,N_613,N_410);
and U861 (N_861,N_483,N_392);
nand U862 (N_862,N_270,N_182);
nand U863 (N_863,N_669,N_300);
or U864 (N_864,N_453,N_512);
or U865 (N_865,N_227,N_90);
or U866 (N_866,N_304,N_318);
or U867 (N_867,N_257,N_357);
and U868 (N_868,N_485,N_279);
nand U869 (N_869,N_346,N_46);
and U870 (N_870,N_516,N_370);
nor U871 (N_871,N_160,N_100);
nand U872 (N_872,N_601,N_665);
or U873 (N_873,N_34,N_351);
and U874 (N_874,N_59,N_146);
and U875 (N_875,N_361,N_156);
or U876 (N_876,N_555,N_153);
nor U877 (N_877,N_476,N_365);
nor U878 (N_878,N_566,N_296);
or U879 (N_879,N_438,N_421);
and U880 (N_880,N_150,N_329);
nand U881 (N_881,N_168,N_462);
and U882 (N_882,N_605,N_679);
and U883 (N_883,N_162,N_714);
or U884 (N_884,N_563,N_517);
nand U885 (N_885,N_727,N_185);
nor U886 (N_886,N_208,N_586);
and U887 (N_887,N_94,N_316);
or U888 (N_888,N_685,N_73);
nor U889 (N_889,N_544,N_681);
nand U890 (N_890,N_19,N_432);
or U891 (N_891,N_689,N_6);
nand U892 (N_892,N_409,N_214);
or U893 (N_893,N_672,N_659);
nor U894 (N_894,N_250,N_163);
nor U895 (N_895,N_621,N_398);
nand U896 (N_896,N_287,N_572);
nor U897 (N_897,N_288,N_140);
nand U898 (N_898,N_597,N_725);
or U899 (N_899,N_692,N_364);
nand U900 (N_900,N_487,N_24);
and U901 (N_901,N_634,N_260);
nor U902 (N_902,N_125,N_667);
and U903 (N_903,N_380,N_372);
nor U904 (N_904,N_43,N_656);
nand U905 (N_905,N_429,N_128);
or U906 (N_906,N_627,N_67);
and U907 (N_907,N_89,N_615);
and U908 (N_908,N_120,N_671);
nand U909 (N_909,N_573,N_56);
nand U910 (N_910,N_562,N_657);
and U911 (N_911,N_404,N_539);
or U912 (N_912,N_245,N_108);
nor U913 (N_913,N_611,N_134);
and U914 (N_914,N_556,N_258);
nand U915 (N_915,N_145,N_687);
nor U916 (N_916,N_466,N_333);
nand U917 (N_917,N_497,N_81);
nor U918 (N_918,N_37,N_717);
nand U919 (N_919,N_583,N_88);
nand U920 (N_920,N_307,N_733);
and U921 (N_921,N_614,N_151);
nand U922 (N_922,N_377,N_589);
and U923 (N_923,N_277,N_701);
nand U924 (N_924,N_321,N_696);
or U925 (N_925,N_641,N_707);
and U926 (N_926,N_47,N_314);
nor U927 (N_927,N_440,N_414);
or U928 (N_928,N_570,N_622);
or U929 (N_929,N_368,N_222);
xor U930 (N_930,N_180,N_578);
or U931 (N_931,N_171,N_147);
nand U932 (N_932,N_303,N_8);
nand U933 (N_933,N_229,N_623);
nor U934 (N_934,N_25,N_286);
and U935 (N_935,N_706,N_273);
or U936 (N_936,N_252,N_353);
and U937 (N_937,N_551,N_495);
or U938 (N_938,N_75,N_619);
nand U939 (N_939,N_653,N_575);
nor U940 (N_940,N_720,N_382);
nand U941 (N_941,N_535,N_580);
and U942 (N_942,N_363,N_259);
nand U943 (N_943,N_747,N_11);
nand U944 (N_944,N_341,N_457);
nand U945 (N_945,N_543,N_241);
nand U946 (N_946,N_741,N_170);
nand U947 (N_947,N_195,N_65);
or U948 (N_948,N_749,N_159);
and U949 (N_949,N_708,N_522);
nor U950 (N_950,N_709,N_740);
or U951 (N_951,N_328,N_371);
nor U952 (N_952,N_135,N_577);
nor U953 (N_953,N_729,N_7);
and U954 (N_954,N_215,N_26);
or U955 (N_955,N_165,N_21);
xnor U956 (N_956,N_426,N_269);
nand U957 (N_957,N_315,N_3);
or U958 (N_958,N_716,N_62);
and U959 (N_959,N_228,N_10);
or U960 (N_960,N_344,N_205);
and U961 (N_961,N_445,N_297);
nor U962 (N_962,N_57,N_557);
and U963 (N_963,N_553,N_78);
and U964 (N_964,N_32,N_686);
nor U965 (N_965,N_690,N_397);
nand U966 (N_966,N_642,N_183);
and U967 (N_967,N_103,N_334);
nor U968 (N_968,N_301,N_69);
and U969 (N_969,N_637,N_122);
and U970 (N_970,N_206,N_246);
nand U971 (N_971,N_431,N_124);
nor U972 (N_972,N_384,N_123);
or U973 (N_973,N_558,N_705);
or U974 (N_974,N_381,N_742);
nand U975 (N_975,N_172,N_518);
and U976 (N_976,N_548,N_710);
nor U977 (N_977,N_74,N_210);
nand U978 (N_978,N_119,N_604);
and U979 (N_979,N_188,N_0);
or U980 (N_980,N_309,N_64);
nor U981 (N_981,N_111,N_20);
nand U982 (N_982,N_268,N_525);
or U983 (N_983,N_567,N_610);
nor U984 (N_984,N_209,N_428);
nand U985 (N_985,N_470,N_662);
nor U986 (N_986,N_324,N_317);
and U987 (N_987,N_85,N_617);
or U988 (N_988,N_84,N_92);
and U989 (N_989,N_549,N_28);
nor U990 (N_990,N_632,N_718);
and U991 (N_991,N_554,N_694);
and U992 (N_992,N_731,N_724);
and U993 (N_993,N_219,N_722);
or U994 (N_994,N_412,N_523);
and U995 (N_995,N_129,N_393);
nor U996 (N_996,N_38,N_373);
nor U997 (N_997,N_249,N_166);
xnor U998 (N_998,N_660,N_477);
or U999 (N_999,N_655,N_96);
nor U1000 (N_1000,N_199,N_16);
or U1001 (N_1001,N_251,N_451);
nor U1002 (N_1002,N_101,N_66);
and U1003 (N_1003,N_191,N_262);
and U1004 (N_1004,N_282,N_233);
or U1005 (N_1005,N_650,N_49);
or U1006 (N_1006,N_508,N_35);
or U1007 (N_1007,N_102,N_141);
nor U1008 (N_1008,N_114,N_326);
or U1009 (N_1009,N_15,N_198);
and U1010 (N_1010,N_97,N_178);
and U1011 (N_1011,N_283,N_231);
and U1012 (N_1012,N_533,N_585);
nor U1013 (N_1013,N_131,N_593);
nor U1014 (N_1014,N_503,N_609);
nand U1015 (N_1015,N_41,N_158);
nor U1016 (N_1016,N_661,N_521);
and U1017 (N_1017,N_423,N_87);
nor U1018 (N_1018,N_253,N_352);
or U1019 (N_1019,N_137,N_442);
or U1020 (N_1020,N_86,N_220);
nand U1021 (N_1021,N_176,N_379);
nor U1022 (N_1022,N_284,N_739);
or U1023 (N_1023,N_29,N_630);
or U1024 (N_1024,N_18,N_737);
nor U1025 (N_1025,N_569,N_389);
nand U1026 (N_1026,N_320,N_360);
nor U1027 (N_1027,N_504,N_527);
nor U1028 (N_1028,N_53,N_649);
nand U1029 (N_1029,N_452,N_390);
nor U1030 (N_1030,N_113,N_76);
nand U1031 (N_1031,N_602,N_267);
and U1032 (N_1032,N_310,N_515);
nand U1033 (N_1033,N_697,N_420);
nand U1034 (N_1034,N_545,N_486);
nand U1035 (N_1035,N_132,N_418);
and U1036 (N_1036,N_99,N_39);
nand U1037 (N_1037,N_629,N_511);
nand U1038 (N_1038,N_524,N_531);
and U1039 (N_1039,N_475,N_244);
nor U1040 (N_1040,N_596,N_348);
and U1041 (N_1041,N_538,N_403);
nor U1042 (N_1042,N_327,N_463);
or U1043 (N_1043,N_663,N_144);
and U1044 (N_1044,N_293,N_699);
nand U1045 (N_1045,N_136,N_369);
or U1046 (N_1046,N_339,N_407);
or U1047 (N_1047,N_491,N_599);
nand U1048 (N_1048,N_715,N_197);
and U1049 (N_1049,N_506,N_173);
nand U1050 (N_1050,N_223,N_143);
nand U1051 (N_1051,N_274,N_424);
or U1052 (N_1052,N_435,N_280);
nor U1053 (N_1053,N_204,N_323);
and U1054 (N_1054,N_648,N_31);
nor U1055 (N_1055,N_496,N_526);
or U1056 (N_1056,N_242,N_289);
and U1057 (N_1057,N_408,N_40);
nand U1058 (N_1058,N_509,N_200);
and U1059 (N_1059,N_387,N_482);
nand U1060 (N_1060,N_574,N_484);
nor U1061 (N_1061,N_236,N_481);
nand U1062 (N_1062,N_441,N_666);
or U1063 (N_1063,N_639,N_263);
nand U1064 (N_1064,N_646,N_444);
and U1065 (N_1065,N_121,N_375);
nor U1066 (N_1066,N_540,N_471);
and U1067 (N_1067,N_30,N_625);
or U1068 (N_1068,N_186,N_499);
nor U1069 (N_1069,N_571,N_618);
or U1070 (N_1070,N_744,N_202);
or U1071 (N_1071,N_582,N_196);
and U1072 (N_1072,N_193,N_728);
nand U1073 (N_1073,N_238,N_345);
or U1074 (N_1074,N_184,N_502);
nand U1075 (N_1075,N_2,N_358);
nor U1076 (N_1076,N_494,N_434);
or U1077 (N_1077,N_478,N_449);
or U1078 (N_1078,N_676,N_332);
nor U1079 (N_1079,N_354,N_748);
nand U1080 (N_1080,N_588,N_207);
and U1081 (N_1081,N_248,N_247);
nand U1082 (N_1082,N_664,N_322);
and U1083 (N_1083,N_624,N_91);
nand U1084 (N_1084,N_175,N_590);
nand U1085 (N_1085,N_474,N_711);
nor U1086 (N_1086,N_415,N_211);
xnor U1087 (N_1087,N_468,N_537);
or U1088 (N_1088,N_355,N_106);
nand U1089 (N_1089,N_350,N_149);
nor U1090 (N_1090,N_117,N_312);
nor U1091 (N_1091,N_63,N_541);
nor U1092 (N_1092,N_386,N_598);
and U1093 (N_1093,N_635,N_628);
nand U1094 (N_1094,N_112,N_606);
nand U1095 (N_1095,N_726,N_93);
and U1096 (N_1096,N_1,N_612);
nand U1097 (N_1097,N_177,N_406);
and U1098 (N_1098,N_730,N_218);
or U1099 (N_1099,N_712,N_174);
nor U1100 (N_1100,N_224,N_704);
and U1101 (N_1101,N_27,N_95);
nor U1102 (N_1102,N_513,N_723);
and U1103 (N_1103,N_239,N_104);
or U1104 (N_1104,N_698,N_592);
or U1105 (N_1105,N_190,N_115);
and U1106 (N_1106,N_272,N_154);
nand U1107 (N_1107,N_459,N_367);
nand U1108 (N_1108,N_565,N_378);
nand U1109 (N_1109,N_472,N_23);
or U1110 (N_1110,N_235,N_148);
and U1111 (N_1111,N_746,N_688);
and U1112 (N_1112,N_488,N_299);
nand U1113 (N_1113,N_677,N_700);
or U1114 (N_1114,N_616,N_394);
nand U1115 (N_1115,N_448,N_581);
nand U1116 (N_1116,N_83,N_42);
or U1117 (N_1117,N_413,N_542);
or U1118 (N_1118,N_447,N_607);
nand U1119 (N_1119,N_520,N_411);
and U1120 (N_1120,N_489,N_422);
nor U1121 (N_1121,N_221,N_670);
and U1122 (N_1122,N_45,N_107);
nand U1123 (N_1123,N_331,N_636);
or U1124 (N_1124,N_52,N_118);
and U1125 (N_1125,N_243,N_134);
or U1126 (N_1126,N_626,N_114);
or U1127 (N_1127,N_404,N_233);
nor U1128 (N_1128,N_369,N_633);
nand U1129 (N_1129,N_357,N_128);
nor U1130 (N_1130,N_295,N_495);
nand U1131 (N_1131,N_40,N_201);
nand U1132 (N_1132,N_738,N_745);
nor U1133 (N_1133,N_500,N_577);
nand U1134 (N_1134,N_491,N_360);
nor U1135 (N_1135,N_722,N_658);
and U1136 (N_1136,N_694,N_38);
or U1137 (N_1137,N_374,N_616);
nor U1138 (N_1138,N_50,N_641);
or U1139 (N_1139,N_662,N_635);
nor U1140 (N_1140,N_720,N_126);
nand U1141 (N_1141,N_527,N_40);
or U1142 (N_1142,N_153,N_441);
or U1143 (N_1143,N_2,N_735);
nor U1144 (N_1144,N_475,N_268);
and U1145 (N_1145,N_85,N_296);
xor U1146 (N_1146,N_260,N_329);
nor U1147 (N_1147,N_738,N_388);
and U1148 (N_1148,N_60,N_649);
nand U1149 (N_1149,N_478,N_639);
nor U1150 (N_1150,N_420,N_459);
and U1151 (N_1151,N_432,N_190);
and U1152 (N_1152,N_18,N_340);
nor U1153 (N_1153,N_576,N_62);
nor U1154 (N_1154,N_198,N_246);
nand U1155 (N_1155,N_309,N_657);
xnor U1156 (N_1156,N_423,N_521);
xnor U1157 (N_1157,N_83,N_358);
or U1158 (N_1158,N_12,N_126);
nor U1159 (N_1159,N_91,N_666);
nand U1160 (N_1160,N_506,N_687);
nand U1161 (N_1161,N_583,N_590);
or U1162 (N_1162,N_233,N_639);
and U1163 (N_1163,N_275,N_492);
and U1164 (N_1164,N_171,N_609);
or U1165 (N_1165,N_193,N_503);
and U1166 (N_1166,N_581,N_403);
and U1167 (N_1167,N_112,N_627);
nand U1168 (N_1168,N_347,N_582);
or U1169 (N_1169,N_701,N_749);
or U1170 (N_1170,N_610,N_463);
and U1171 (N_1171,N_14,N_589);
nand U1172 (N_1172,N_401,N_726);
or U1173 (N_1173,N_682,N_93);
and U1174 (N_1174,N_502,N_270);
nand U1175 (N_1175,N_204,N_12);
or U1176 (N_1176,N_485,N_31);
and U1177 (N_1177,N_667,N_607);
nand U1178 (N_1178,N_650,N_100);
nor U1179 (N_1179,N_414,N_201);
or U1180 (N_1180,N_449,N_9);
nand U1181 (N_1181,N_175,N_138);
nand U1182 (N_1182,N_133,N_502);
nor U1183 (N_1183,N_68,N_471);
nand U1184 (N_1184,N_517,N_690);
or U1185 (N_1185,N_123,N_356);
nand U1186 (N_1186,N_202,N_312);
or U1187 (N_1187,N_541,N_24);
nand U1188 (N_1188,N_19,N_343);
nor U1189 (N_1189,N_215,N_361);
nand U1190 (N_1190,N_289,N_420);
or U1191 (N_1191,N_315,N_507);
nor U1192 (N_1192,N_508,N_320);
and U1193 (N_1193,N_539,N_154);
nor U1194 (N_1194,N_705,N_139);
xnor U1195 (N_1195,N_129,N_477);
and U1196 (N_1196,N_678,N_144);
or U1197 (N_1197,N_410,N_281);
nor U1198 (N_1198,N_425,N_577);
nor U1199 (N_1199,N_588,N_704);
or U1200 (N_1200,N_504,N_418);
or U1201 (N_1201,N_288,N_737);
and U1202 (N_1202,N_52,N_367);
nand U1203 (N_1203,N_63,N_51);
or U1204 (N_1204,N_192,N_278);
nor U1205 (N_1205,N_465,N_375);
nor U1206 (N_1206,N_493,N_62);
nand U1207 (N_1207,N_749,N_194);
nand U1208 (N_1208,N_588,N_550);
nand U1209 (N_1209,N_68,N_513);
nor U1210 (N_1210,N_194,N_83);
or U1211 (N_1211,N_547,N_660);
and U1212 (N_1212,N_177,N_101);
nand U1213 (N_1213,N_407,N_323);
or U1214 (N_1214,N_288,N_12);
nand U1215 (N_1215,N_201,N_307);
and U1216 (N_1216,N_592,N_733);
or U1217 (N_1217,N_477,N_161);
nand U1218 (N_1218,N_286,N_574);
and U1219 (N_1219,N_662,N_104);
nand U1220 (N_1220,N_747,N_53);
nand U1221 (N_1221,N_700,N_348);
or U1222 (N_1222,N_451,N_268);
nor U1223 (N_1223,N_505,N_212);
and U1224 (N_1224,N_401,N_559);
nand U1225 (N_1225,N_43,N_664);
or U1226 (N_1226,N_713,N_235);
nand U1227 (N_1227,N_625,N_577);
and U1228 (N_1228,N_731,N_319);
nor U1229 (N_1229,N_27,N_475);
or U1230 (N_1230,N_218,N_358);
nor U1231 (N_1231,N_203,N_221);
and U1232 (N_1232,N_246,N_257);
nor U1233 (N_1233,N_421,N_63);
nand U1234 (N_1234,N_672,N_159);
nor U1235 (N_1235,N_406,N_529);
nand U1236 (N_1236,N_747,N_656);
or U1237 (N_1237,N_241,N_652);
nand U1238 (N_1238,N_218,N_204);
or U1239 (N_1239,N_221,N_216);
nor U1240 (N_1240,N_321,N_675);
nor U1241 (N_1241,N_587,N_591);
nand U1242 (N_1242,N_386,N_24);
nor U1243 (N_1243,N_454,N_381);
nand U1244 (N_1244,N_382,N_526);
xor U1245 (N_1245,N_736,N_397);
or U1246 (N_1246,N_92,N_285);
nor U1247 (N_1247,N_447,N_496);
and U1248 (N_1248,N_299,N_10);
and U1249 (N_1249,N_676,N_649);
and U1250 (N_1250,N_92,N_659);
and U1251 (N_1251,N_301,N_698);
and U1252 (N_1252,N_17,N_656);
and U1253 (N_1253,N_708,N_232);
or U1254 (N_1254,N_201,N_739);
or U1255 (N_1255,N_408,N_435);
nand U1256 (N_1256,N_173,N_672);
or U1257 (N_1257,N_40,N_696);
or U1258 (N_1258,N_424,N_588);
nand U1259 (N_1259,N_265,N_293);
nor U1260 (N_1260,N_452,N_6);
and U1261 (N_1261,N_377,N_365);
nand U1262 (N_1262,N_1,N_23);
nor U1263 (N_1263,N_64,N_552);
and U1264 (N_1264,N_651,N_363);
nand U1265 (N_1265,N_423,N_24);
nand U1266 (N_1266,N_12,N_605);
nand U1267 (N_1267,N_604,N_401);
and U1268 (N_1268,N_67,N_734);
nand U1269 (N_1269,N_62,N_140);
nor U1270 (N_1270,N_59,N_680);
or U1271 (N_1271,N_64,N_234);
nor U1272 (N_1272,N_741,N_63);
or U1273 (N_1273,N_22,N_71);
nand U1274 (N_1274,N_232,N_280);
and U1275 (N_1275,N_72,N_563);
or U1276 (N_1276,N_676,N_232);
or U1277 (N_1277,N_400,N_388);
and U1278 (N_1278,N_303,N_452);
or U1279 (N_1279,N_144,N_64);
or U1280 (N_1280,N_343,N_235);
nand U1281 (N_1281,N_439,N_88);
nor U1282 (N_1282,N_154,N_491);
or U1283 (N_1283,N_36,N_415);
and U1284 (N_1284,N_74,N_496);
nor U1285 (N_1285,N_107,N_455);
nand U1286 (N_1286,N_582,N_225);
nor U1287 (N_1287,N_367,N_282);
nor U1288 (N_1288,N_468,N_287);
nor U1289 (N_1289,N_284,N_451);
nor U1290 (N_1290,N_568,N_581);
and U1291 (N_1291,N_123,N_70);
and U1292 (N_1292,N_687,N_238);
or U1293 (N_1293,N_669,N_107);
or U1294 (N_1294,N_569,N_563);
nand U1295 (N_1295,N_374,N_562);
or U1296 (N_1296,N_654,N_228);
and U1297 (N_1297,N_245,N_566);
nand U1298 (N_1298,N_572,N_531);
or U1299 (N_1299,N_595,N_301);
nand U1300 (N_1300,N_547,N_523);
nand U1301 (N_1301,N_197,N_393);
nand U1302 (N_1302,N_659,N_176);
nor U1303 (N_1303,N_176,N_691);
or U1304 (N_1304,N_306,N_638);
and U1305 (N_1305,N_57,N_46);
xor U1306 (N_1306,N_496,N_576);
nand U1307 (N_1307,N_516,N_519);
and U1308 (N_1308,N_499,N_578);
nor U1309 (N_1309,N_733,N_197);
and U1310 (N_1310,N_675,N_600);
nor U1311 (N_1311,N_258,N_722);
or U1312 (N_1312,N_306,N_484);
nand U1313 (N_1313,N_705,N_568);
nand U1314 (N_1314,N_32,N_64);
and U1315 (N_1315,N_572,N_698);
nor U1316 (N_1316,N_52,N_321);
xor U1317 (N_1317,N_400,N_556);
nor U1318 (N_1318,N_744,N_229);
or U1319 (N_1319,N_98,N_584);
nand U1320 (N_1320,N_455,N_130);
or U1321 (N_1321,N_213,N_207);
and U1322 (N_1322,N_638,N_616);
nor U1323 (N_1323,N_459,N_548);
nand U1324 (N_1324,N_44,N_457);
and U1325 (N_1325,N_195,N_386);
nor U1326 (N_1326,N_608,N_368);
and U1327 (N_1327,N_484,N_232);
and U1328 (N_1328,N_101,N_337);
nor U1329 (N_1329,N_437,N_533);
or U1330 (N_1330,N_669,N_464);
nand U1331 (N_1331,N_262,N_342);
and U1332 (N_1332,N_710,N_305);
nor U1333 (N_1333,N_352,N_477);
or U1334 (N_1334,N_357,N_660);
or U1335 (N_1335,N_293,N_134);
or U1336 (N_1336,N_340,N_676);
or U1337 (N_1337,N_691,N_213);
nand U1338 (N_1338,N_566,N_278);
or U1339 (N_1339,N_106,N_72);
nand U1340 (N_1340,N_511,N_496);
nand U1341 (N_1341,N_640,N_197);
nand U1342 (N_1342,N_211,N_706);
nor U1343 (N_1343,N_460,N_569);
or U1344 (N_1344,N_195,N_685);
and U1345 (N_1345,N_339,N_270);
nor U1346 (N_1346,N_201,N_270);
or U1347 (N_1347,N_131,N_171);
nor U1348 (N_1348,N_51,N_379);
nand U1349 (N_1349,N_582,N_28);
or U1350 (N_1350,N_120,N_443);
and U1351 (N_1351,N_532,N_293);
and U1352 (N_1352,N_13,N_247);
nand U1353 (N_1353,N_4,N_203);
and U1354 (N_1354,N_349,N_111);
and U1355 (N_1355,N_185,N_95);
nor U1356 (N_1356,N_104,N_374);
xor U1357 (N_1357,N_261,N_746);
and U1358 (N_1358,N_464,N_449);
nor U1359 (N_1359,N_171,N_660);
or U1360 (N_1360,N_709,N_176);
or U1361 (N_1361,N_635,N_622);
and U1362 (N_1362,N_157,N_266);
and U1363 (N_1363,N_280,N_63);
nor U1364 (N_1364,N_449,N_51);
or U1365 (N_1365,N_684,N_545);
or U1366 (N_1366,N_579,N_728);
or U1367 (N_1367,N_88,N_126);
and U1368 (N_1368,N_671,N_548);
and U1369 (N_1369,N_419,N_693);
nor U1370 (N_1370,N_126,N_172);
nor U1371 (N_1371,N_362,N_696);
nand U1372 (N_1372,N_561,N_427);
nor U1373 (N_1373,N_613,N_296);
and U1374 (N_1374,N_406,N_98);
or U1375 (N_1375,N_385,N_36);
nor U1376 (N_1376,N_439,N_173);
and U1377 (N_1377,N_292,N_731);
nand U1378 (N_1378,N_215,N_528);
or U1379 (N_1379,N_272,N_183);
nor U1380 (N_1380,N_115,N_285);
nand U1381 (N_1381,N_113,N_14);
nand U1382 (N_1382,N_201,N_625);
and U1383 (N_1383,N_711,N_130);
nand U1384 (N_1384,N_353,N_640);
nand U1385 (N_1385,N_181,N_63);
nand U1386 (N_1386,N_562,N_14);
or U1387 (N_1387,N_373,N_639);
nor U1388 (N_1388,N_0,N_301);
nand U1389 (N_1389,N_518,N_199);
or U1390 (N_1390,N_311,N_669);
and U1391 (N_1391,N_23,N_642);
or U1392 (N_1392,N_451,N_28);
and U1393 (N_1393,N_306,N_412);
nand U1394 (N_1394,N_323,N_616);
and U1395 (N_1395,N_270,N_374);
nand U1396 (N_1396,N_674,N_60);
or U1397 (N_1397,N_152,N_79);
or U1398 (N_1398,N_741,N_236);
nand U1399 (N_1399,N_702,N_110);
nand U1400 (N_1400,N_361,N_419);
nor U1401 (N_1401,N_638,N_218);
and U1402 (N_1402,N_51,N_721);
nand U1403 (N_1403,N_195,N_557);
nor U1404 (N_1404,N_569,N_390);
and U1405 (N_1405,N_99,N_205);
or U1406 (N_1406,N_169,N_45);
or U1407 (N_1407,N_735,N_525);
and U1408 (N_1408,N_390,N_159);
and U1409 (N_1409,N_612,N_566);
or U1410 (N_1410,N_610,N_411);
nand U1411 (N_1411,N_438,N_84);
and U1412 (N_1412,N_451,N_228);
and U1413 (N_1413,N_577,N_523);
nand U1414 (N_1414,N_86,N_174);
or U1415 (N_1415,N_98,N_269);
and U1416 (N_1416,N_64,N_8);
nand U1417 (N_1417,N_716,N_506);
nor U1418 (N_1418,N_690,N_6);
nand U1419 (N_1419,N_38,N_73);
or U1420 (N_1420,N_6,N_613);
or U1421 (N_1421,N_52,N_271);
nand U1422 (N_1422,N_602,N_143);
nor U1423 (N_1423,N_546,N_534);
nor U1424 (N_1424,N_594,N_598);
nor U1425 (N_1425,N_317,N_510);
or U1426 (N_1426,N_280,N_41);
or U1427 (N_1427,N_337,N_184);
or U1428 (N_1428,N_53,N_504);
and U1429 (N_1429,N_404,N_622);
nor U1430 (N_1430,N_267,N_575);
and U1431 (N_1431,N_125,N_392);
or U1432 (N_1432,N_579,N_389);
nand U1433 (N_1433,N_334,N_243);
or U1434 (N_1434,N_197,N_111);
nor U1435 (N_1435,N_220,N_639);
nor U1436 (N_1436,N_53,N_312);
nand U1437 (N_1437,N_339,N_621);
and U1438 (N_1438,N_24,N_295);
or U1439 (N_1439,N_425,N_578);
or U1440 (N_1440,N_362,N_250);
nor U1441 (N_1441,N_149,N_74);
or U1442 (N_1442,N_178,N_410);
nand U1443 (N_1443,N_657,N_84);
and U1444 (N_1444,N_383,N_334);
nor U1445 (N_1445,N_662,N_361);
and U1446 (N_1446,N_697,N_385);
or U1447 (N_1447,N_136,N_228);
nand U1448 (N_1448,N_238,N_52);
and U1449 (N_1449,N_173,N_470);
and U1450 (N_1450,N_725,N_570);
nor U1451 (N_1451,N_396,N_568);
or U1452 (N_1452,N_283,N_719);
nand U1453 (N_1453,N_12,N_359);
or U1454 (N_1454,N_488,N_265);
nand U1455 (N_1455,N_687,N_51);
nor U1456 (N_1456,N_613,N_645);
or U1457 (N_1457,N_463,N_723);
and U1458 (N_1458,N_314,N_705);
and U1459 (N_1459,N_131,N_34);
nor U1460 (N_1460,N_292,N_218);
nand U1461 (N_1461,N_329,N_537);
nor U1462 (N_1462,N_203,N_574);
and U1463 (N_1463,N_48,N_258);
nor U1464 (N_1464,N_724,N_425);
nand U1465 (N_1465,N_643,N_729);
or U1466 (N_1466,N_728,N_317);
nand U1467 (N_1467,N_690,N_703);
or U1468 (N_1468,N_240,N_253);
and U1469 (N_1469,N_624,N_110);
or U1470 (N_1470,N_138,N_587);
and U1471 (N_1471,N_108,N_665);
nand U1472 (N_1472,N_282,N_330);
or U1473 (N_1473,N_480,N_305);
or U1474 (N_1474,N_99,N_660);
and U1475 (N_1475,N_530,N_201);
or U1476 (N_1476,N_345,N_561);
nand U1477 (N_1477,N_647,N_709);
nand U1478 (N_1478,N_111,N_72);
nor U1479 (N_1479,N_425,N_466);
nor U1480 (N_1480,N_31,N_432);
nand U1481 (N_1481,N_33,N_362);
or U1482 (N_1482,N_720,N_305);
or U1483 (N_1483,N_614,N_432);
or U1484 (N_1484,N_142,N_416);
nand U1485 (N_1485,N_204,N_64);
nor U1486 (N_1486,N_709,N_82);
nand U1487 (N_1487,N_444,N_471);
nand U1488 (N_1488,N_589,N_562);
and U1489 (N_1489,N_682,N_599);
and U1490 (N_1490,N_201,N_368);
or U1491 (N_1491,N_609,N_507);
nor U1492 (N_1492,N_675,N_123);
nand U1493 (N_1493,N_570,N_740);
or U1494 (N_1494,N_185,N_167);
nor U1495 (N_1495,N_327,N_1);
nand U1496 (N_1496,N_717,N_124);
nor U1497 (N_1497,N_374,N_310);
and U1498 (N_1498,N_92,N_407);
or U1499 (N_1499,N_519,N_258);
nor U1500 (N_1500,N_1112,N_1209);
nand U1501 (N_1501,N_1361,N_933);
or U1502 (N_1502,N_925,N_1492);
nand U1503 (N_1503,N_1034,N_1074);
nor U1504 (N_1504,N_1077,N_1351);
or U1505 (N_1505,N_777,N_1494);
or U1506 (N_1506,N_1484,N_1315);
nand U1507 (N_1507,N_1240,N_1460);
and U1508 (N_1508,N_815,N_1142);
nor U1509 (N_1509,N_1357,N_1038);
and U1510 (N_1510,N_888,N_1427);
or U1511 (N_1511,N_1172,N_904);
nand U1512 (N_1512,N_1375,N_1325);
and U1513 (N_1513,N_1115,N_958);
or U1514 (N_1514,N_882,N_1407);
nor U1515 (N_1515,N_1064,N_808);
nand U1516 (N_1516,N_985,N_922);
or U1517 (N_1517,N_1195,N_1014);
or U1518 (N_1518,N_1045,N_1436);
nor U1519 (N_1519,N_874,N_1071);
nand U1520 (N_1520,N_964,N_960);
or U1521 (N_1521,N_1400,N_1477);
or U1522 (N_1522,N_1211,N_1030);
nand U1523 (N_1523,N_1449,N_896);
nor U1524 (N_1524,N_990,N_1300);
or U1525 (N_1525,N_1339,N_956);
or U1526 (N_1526,N_914,N_982);
nand U1527 (N_1527,N_1164,N_1466);
nor U1528 (N_1528,N_943,N_1213);
or U1529 (N_1529,N_1270,N_861);
nand U1530 (N_1530,N_1148,N_1403);
nor U1531 (N_1531,N_1323,N_1496);
nor U1532 (N_1532,N_1473,N_879);
or U1533 (N_1533,N_1435,N_1157);
nand U1534 (N_1534,N_1425,N_1192);
or U1535 (N_1535,N_1495,N_767);
nor U1536 (N_1536,N_1346,N_760);
and U1537 (N_1537,N_1061,N_1440);
or U1538 (N_1538,N_1016,N_1200);
or U1539 (N_1539,N_1311,N_868);
nor U1540 (N_1540,N_847,N_932);
nand U1541 (N_1541,N_1131,N_970);
nand U1542 (N_1542,N_974,N_1010);
nand U1543 (N_1543,N_934,N_1120);
nor U1544 (N_1544,N_1432,N_1210);
nand U1545 (N_1545,N_949,N_1220);
nor U1546 (N_1546,N_1146,N_794);
nor U1547 (N_1547,N_1415,N_1006);
and U1548 (N_1548,N_776,N_1292);
and U1549 (N_1549,N_1499,N_1469);
nand U1550 (N_1550,N_1025,N_961);
or U1551 (N_1551,N_1453,N_1019);
or U1552 (N_1552,N_871,N_848);
or U1553 (N_1553,N_1481,N_1281);
and U1554 (N_1554,N_762,N_911);
nor U1555 (N_1555,N_792,N_1386);
and U1556 (N_1556,N_787,N_1486);
nor U1557 (N_1557,N_1321,N_1332);
and U1558 (N_1558,N_814,N_1297);
and U1559 (N_1559,N_1276,N_1185);
or U1560 (N_1560,N_862,N_1135);
nand U1561 (N_1561,N_757,N_1116);
and U1562 (N_1562,N_953,N_1405);
nand U1563 (N_1563,N_1046,N_1450);
nor U1564 (N_1564,N_1150,N_1479);
nor U1565 (N_1565,N_1387,N_1416);
nand U1566 (N_1566,N_1483,N_1487);
xnor U1567 (N_1567,N_1129,N_1409);
nand U1568 (N_1568,N_1255,N_889);
nand U1569 (N_1569,N_969,N_1385);
nand U1570 (N_1570,N_1250,N_1137);
nand U1571 (N_1571,N_995,N_986);
and U1572 (N_1572,N_1284,N_1169);
nand U1573 (N_1573,N_1491,N_860);
or U1574 (N_1574,N_863,N_1467);
or U1575 (N_1575,N_805,N_1028);
or U1576 (N_1576,N_1293,N_1207);
and U1577 (N_1577,N_1406,N_906);
or U1578 (N_1578,N_1048,N_1335);
and U1579 (N_1579,N_1099,N_1160);
and U1580 (N_1580,N_920,N_946);
nor U1581 (N_1581,N_1431,N_1272);
nand U1582 (N_1582,N_786,N_1227);
or U1583 (N_1583,N_916,N_1102);
or U1584 (N_1584,N_1373,N_1404);
or U1585 (N_1585,N_1318,N_1352);
and U1586 (N_1586,N_826,N_765);
and U1587 (N_1587,N_793,N_1362);
nand U1588 (N_1588,N_1041,N_820);
or U1589 (N_1589,N_1419,N_1094);
nor U1590 (N_1590,N_1465,N_796);
or U1591 (N_1591,N_1412,N_1100);
nor U1592 (N_1592,N_1127,N_1333);
nor U1593 (N_1593,N_1394,N_756);
or U1594 (N_1594,N_1219,N_1012);
nand U1595 (N_1595,N_1475,N_1249);
nor U1596 (N_1596,N_1269,N_1065);
and U1597 (N_1597,N_1290,N_1152);
nor U1598 (N_1598,N_901,N_1086);
and U1599 (N_1599,N_893,N_1130);
or U1600 (N_1600,N_1391,N_1277);
or U1601 (N_1601,N_1085,N_1295);
and U1602 (N_1602,N_1162,N_1205);
or U1603 (N_1603,N_1196,N_799);
nand U1604 (N_1604,N_1263,N_1447);
nand U1605 (N_1605,N_1165,N_1398);
and U1606 (N_1606,N_1091,N_1093);
nand U1607 (N_1607,N_1124,N_1376);
nor U1608 (N_1608,N_837,N_1066);
and U1609 (N_1609,N_1215,N_1001);
and U1610 (N_1610,N_1326,N_1155);
nor U1611 (N_1611,N_1004,N_780);
nand U1612 (N_1612,N_1364,N_1365);
nand U1613 (N_1613,N_1265,N_1374);
and U1614 (N_1614,N_918,N_929);
nor U1615 (N_1615,N_1348,N_910);
nand U1616 (N_1616,N_1360,N_905);
nor U1617 (N_1617,N_1083,N_1147);
or U1618 (N_1618,N_1478,N_1134);
and U1619 (N_1619,N_994,N_1096);
nand U1620 (N_1620,N_790,N_887);
or U1621 (N_1621,N_839,N_761);
or U1622 (N_1622,N_1214,N_1232);
or U1623 (N_1623,N_923,N_819);
or U1624 (N_1624,N_1109,N_1050);
or U1625 (N_1625,N_1183,N_1203);
or U1626 (N_1626,N_1345,N_1336);
and U1627 (N_1627,N_1382,N_962);
nor U1628 (N_1628,N_1184,N_886);
xor U1629 (N_1629,N_1383,N_816);
or U1630 (N_1630,N_1231,N_997);
and U1631 (N_1631,N_1344,N_784);
nor U1632 (N_1632,N_1397,N_857);
and U1633 (N_1633,N_927,N_967);
or U1634 (N_1634,N_1088,N_1461);
nor U1635 (N_1635,N_821,N_753);
and U1636 (N_1636,N_832,N_1328);
nor U1637 (N_1637,N_1110,N_989);
nor U1638 (N_1638,N_800,N_754);
and U1639 (N_1639,N_1390,N_1138);
and U1640 (N_1640,N_1218,N_1118);
or U1641 (N_1641,N_951,N_1191);
and U1642 (N_1642,N_1471,N_883);
xnor U1643 (N_1643,N_766,N_1414);
or U1644 (N_1644,N_877,N_843);
and U1645 (N_1645,N_1437,N_1101);
or U1646 (N_1646,N_1489,N_1455);
or U1647 (N_1647,N_1485,N_1125);
or U1648 (N_1648,N_865,N_1291);
and U1649 (N_1649,N_1171,N_1056);
nor U1650 (N_1650,N_1395,N_1243);
and U1651 (N_1651,N_1279,N_836);
or U1652 (N_1652,N_1474,N_1079);
nand U1653 (N_1653,N_1384,N_1178);
and U1654 (N_1654,N_1410,N_1123);
nand U1655 (N_1655,N_1128,N_1354);
and U1656 (N_1656,N_919,N_957);
nand U1657 (N_1657,N_1229,N_789);
and U1658 (N_1658,N_824,N_1073);
or U1659 (N_1659,N_1188,N_1081);
and U1660 (N_1660,N_1228,N_1298);
or U1661 (N_1661,N_1040,N_1262);
nor U1662 (N_1662,N_1458,N_779);
and U1663 (N_1663,N_885,N_1241);
nand U1664 (N_1664,N_1063,N_1433);
nor U1665 (N_1665,N_1245,N_1417);
and U1666 (N_1666,N_1076,N_1342);
nor U1667 (N_1667,N_952,N_1158);
nand U1668 (N_1668,N_1426,N_1133);
nand U1669 (N_1669,N_1264,N_1173);
or U1670 (N_1670,N_1121,N_1015);
and U1671 (N_1671,N_1170,N_1089);
or U1672 (N_1672,N_1441,N_813);
or U1673 (N_1673,N_1057,N_1259);
and U1674 (N_1674,N_1381,N_1055);
or U1675 (N_1675,N_1206,N_1039);
nand U1676 (N_1676,N_1472,N_1468);
xor U1677 (N_1677,N_1343,N_1108);
nand U1678 (N_1678,N_954,N_1371);
nor U1679 (N_1679,N_1197,N_998);
nor U1680 (N_1680,N_1372,N_1226);
nand U1681 (N_1681,N_1018,N_1166);
nand U1682 (N_1682,N_1363,N_1238);
or U1683 (N_1683,N_1418,N_1256);
or U1684 (N_1684,N_856,N_1430);
nand U1685 (N_1685,N_1009,N_1463);
or U1686 (N_1686,N_781,N_1498);
or U1687 (N_1687,N_1003,N_1182);
nand U1688 (N_1688,N_1257,N_1180);
and U1689 (N_1689,N_936,N_1072);
and U1690 (N_1690,N_1296,N_1439);
nor U1691 (N_1691,N_999,N_921);
nand U1692 (N_1692,N_768,N_890);
nor U1693 (N_1693,N_850,N_944);
nor U1694 (N_1694,N_1026,N_1049);
and U1695 (N_1695,N_1189,N_1023);
nand U1696 (N_1696,N_976,N_900);
nor U1697 (N_1697,N_1198,N_1080);
nor U1698 (N_1698,N_1271,N_1070);
or U1699 (N_1699,N_1275,N_1451);
and U1700 (N_1700,N_1389,N_1338);
nand U1701 (N_1701,N_924,N_898);
or U1702 (N_1702,N_1031,N_1236);
or U1703 (N_1703,N_977,N_1052);
or U1704 (N_1704,N_908,N_915);
xor U1705 (N_1705,N_913,N_1267);
nor U1706 (N_1706,N_1244,N_1482);
or U1707 (N_1707,N_869,N_1078);
or U1708 (N_1708,N_912,N_897);
nand U1709 (N_1709,N_867,N_759);
nor U1710 (N_1710,N_1201,N_1266);
nand U1711 (N_1711,N_1208,N_1017);
or U1712 (N_1712,N_1497,N_1286);
nand U1713 (N_1713,N_1320,N_1358);
nor U1714 (N_1714,N_1204,N_1002);
nand U1715 (N_1715,N_1119,N_1105);
or U1716 (N_1716,N_834,N_1153);
nand U1717 (N_1717,N_1175,N_1464);
nand U1718 (N_1718,N_1177,N_1225);
and U1719 (N_1719,N_981,N_846);
and U1720 (N_1720,N_1082,N_1420);
and U1721 (N_1721,N_1370,N_1047);
and U1722 (N_1722,N_769,N_1429);
nor U1723 (N_1723,N_1239,N_1424);
nor U1724 (N_1724,N_764,N_1434);
nand U1725 (N_1725,N_1330,N_1037);
or U1726 (N_1726,N_1104,N_1036);
nor U1727 (N_1727,N_978,N_975);
nand U1728 (N_1728,N_941,N_1285);
and U1729 (N_1729,N_1470,N_1107);
and U1730 (N_1730,N_1313,N_1062);
or U1731 (N_1731,N_963,N_1233);
or U1732 (N_1732,N_845,N_798);
or U1733 (N_1733,N_947,N_1139);
nor U1734 (N_1734,N_835,N_1307);
or U1735 (N_1735,N_1457,N_945);
and U1736 (N_1736,N_875,N_1349);
nand U1737 (N_1737,N_1174,N_1042);
or U1738 (N_1738,N_1117,N_1401);
nand U1739 (N_1739,N_881,N_1221);
nand U1740 (N_1740,N_849,N_852);
nor U1741 (N_1741,N_1008,N_965);
nand U1742 (N_1742,N_1179,N_1033);
nor U1743 (N_1743,N_1224,N_822);
and U1744 (N_1744,N_1258,N_755);
or U1745 (N_1745,N_1377,N_1024);
and U1746 (N_1746,N_903,N_1248);
nand U1747 (N_1747,N_1319,N_1278);
and U1748 (N_1748,N_1329,N_1480);
or U1749 (N_1749,N_894,N_872);
nor U1750 (N_1750,N_1168,N_983);
nand U1751 (N_1751,N_1011,N_907);
nand U1752 (N_1752,N_892,N_1421);
and U1753 (N_1753,N_1044,N_1163);
nor U1754 (N_1754,N_1299,N_1212);
or U1755 (N_1755,N_831,N_859);
nor U1756 (N_1756,N_1246,N_1490);
and U1757 (N_1757,N_1443,N_1359);
and U1758 (N_1758,N_1438,N_1442);
nand U1759 (N_1759,N_854,N_1058);
or U1760 (N_1760,N_1428,N_763);
nor U1761 (N_1761,N_1223,N_1251);
and U1762 (N_1762,N_1310,N_926);
nand U1763 (N_1763,N_1303,N_771);
nor U1764 (N_1764,N_770,N_1022);
or U1765 (N_1765,N_1067,N_1476);
and U1766 (N_1766,N_1393,N_1446);
or U1767 (N_1767,N_1273,N_1156);
nor U1768 (N_1768,N_1230,N_1388);
nand U1769 (N_1769,N_1422,N_1347);
and U1770 (N_1770,N_1305,N_1316);
and U1771 (N_1771,N_1253,N_778);
or U1772 (N_1772,N_1114,N_1402);
or U1773 (N_1773,N_1304,N_1268);
or U1774 (N_1774,N_806,N_1282);
and U1775 (N_1775,N_1029,N_1252);
and U1776 (N_1776,N_1366,N_750);
and U1777 (N_1777,N_909,N_1322);
nand U1778 (N_1778,N_1314,N_1217);
and U1779 (N_1779,N_984,N_788);
nor U1780 (N_1780,N_1122,N_817);
and U1781 (N_1781,N_1098,N_818);
nand U1782 (N_1782,N_993,N_1260);
nor U1783 (N_1783,N_1126,N_1020);
or U1784 (N_1784,N_782,N_988);
and U1785 (N_1785,N_1035,N_855);
or U1786 (N_1786,N_758,N_1144);
and U1787 (N_1787,N_895,N_917);
nor U1788 (N_1788,N_785,N_1097);
nor U1789 (N_1789,N_942,N_1167);
nand U1790 (N_1790,N_841,N_1154);
nor U1791 (N_1791,N_1187,N_939);
and U1792 (N_1792,N_801,N_752);
or U1793 (N_1793,N_1069,N_1059);
nand U1794 (N_1794,N_804,N_1087);
or U1795 (N_1795,N_1222,N_1161);
or U1796 (N_1796,N_1176,N_1302);
nand U1797 (N_1797,N_1199,N_1095);
nand U1798 (N_1798,N_1151,N_991);
nand U1799 (N_1799,N_853,N_1235);
and U1800 (N_1800,N_840,N_992);
xor U1801 (N_1801,N_1350,N_823);
and U1802 (N_1802,N_1488,N_775);
and U1803 (N_1803,N_1092,N_1306);
nor U1804 (N_1804,N_1337,N_928);
or U1805 (N_1805,N_774,N_1053);
or U1806 (N_1806,N_803,N_1159);
nor U1807 (N_1807,N_1355,N_1448);
nand U1808 (N_1808,N_809,N_1324);
nor U1809 (N_1809,N_899,N_1423);
or U1810 (N_1810,N_1202,N_1021);
or U1811 (N_1811,N_1111,N_884);
nor U1812 (N_1812,N_1247,N_940);
nor U1813 (N_1813,N_966,N_935);
and U1814 (N_1814,N_1043,N_807);
nor U1815 (N_1815,N_783,N_1274);
and U1816 (N_1816,N_876,N_1294);
nand U1817 (N_1817,N_937,N_1216);
or U1818 (N_1818,N_1190,N_864);
or U1819 (N_1819,N_1186,N_1234);
nor U1820 (N_1820,N_1334,N_1367);
nor U1821 (N_1821,N_1288,N_870);
nor U1822 (N_1822,N_1301,N_1032);
nor U1823 (N_1823,N_1084,N_1369);
nand U1824 (N_1824,N_825,N_1075);
nand U1825 (N_1825,N_1140,N_1090);
or U1826 (N_1826,N_1051,N_1242);
nor U1827 (N_1827,N_1136,N_1413);
nand U1828 (N_1828,N_797,N_829);
or U1829 (N_1829,N_1327,N_858);
nor U1830 (N_1830,N_1459,N_878);
nor U1831 (N_1831,N_833,N_987);
nor U1832 (N_1832,N_1454,N_851);
nor U1833 (N_1833,N_1289,N_1309);
nand U1834 (N_1834,N_1194,N_968);
nor U1835 (N_1835,N_972,N_1380);
nor U1836 (N_1836,N_959,N_902);
nor U1837 (N_1837,N_1396,N_1143);
nor U1838 (N_1838,N_751,N_795);
and U1839 (N_1839,N_880,N_1340);
nand U1840 (N_1840,N_973,N_1054);
and U1841 (N_1841,N_1445,N_1149);
nand U1842 (N_1842,N_1379,N_996);
and U1843 (N_1843,N_1399,N_1005);
and U1844 (N_1844,N_950,N_979);
and U1845 (N_1845,N_1113,N_1287);
and U1846 (N_1846,N_1068,N_1411);
nor U1847 (N_1847,N_1331,N_1378);
nor U1848 (N_1848,N_1408,N_802);
or U1849 (N_1849,N_773,N_1462);
nand U1850 (N_1850,N_930,N_971);
nand U1851 (N_1851,N_1493,N_1254);
nor U1852 (N_1852,N_1237,N_1392);
and U1853 (N_1853,N_873,N_1283);
nor U1854 (N_1854,N_891,N_1353);
nor U1855 (N_1855,N_1456,N_866);
and U1856 (N_1856,N_1280,N_1141);
nor U1857 (N_1857,N_938,N_1356);
and U1858 (N_1858,N_772,N_1013);
or U1859 (N_1859,N_811,N_1060);
or U1860 (N_1860,N_830,N_828);
and U1861 (N_1861,N_1444,N_1181);
nor U1862 (N_1862,N_1027,N_980);
and U1863 (N_1863,N_1145,N_931);
nor U1864 (N_1864,N_1308,N_812);
or U1865 (N_1865,N_791,N_1132);
nand U1866 (N_1866,N_1341,N_1103);
and U1867 (N_1867,N_1312,N_827);
or U1868 (N_1868,N_955,N_1452);
or U1869 (N_1869,N_1193,N_1317);
or U1870 (N_1870,N_1106,N_842);
nand U1871 (N_1871,N_844,N_838);
nor U1872 (N_1872,N_1000,N_1007);
or U1873 (N_1873,N_810,N_948);
nand U1874 (N_1874,N_1261,N_1368);
or U1875 (N_1875,N_1096,N_870);
nor U1876 (N_1876,N_1498,N_1284);
nor U1877 (N_1877,N_1272,N_1007);
or U1878 (N_1878,N_1124,N_1299);
nand U1879 (N_1879,N_1366,N_1374);
nor U1880 (N_1880,N_900,N_971);
and U1881 (N_1881,N_1309,N_954);
and U1882 (N_1882,N_1261,N_807);
nand U1883 (N_1883,N_1289,N_1006);
nand U1884 (N_1884,N_1238,N_1020);
nor U1885 (N_1885,N_919,N_1021);
nor U1886 (N_1886,N_1150,N_1091);
and U1887 (N_1887,N_1014,N_774);
or U1888 (N_1888,N_1464,N_1185);
and U1889 (N_1889,N_945,N_895);
nand U1890 (N_1890,N_1098,N_1490);
and U1891 (N_1891,N_1380,N_762);
or U1892 (N_1892,N_1152,N_1383);
nor U1893 (N_1893,N_1297,N_1246);
nand U1894 (N_1894,N_1319,N_1432);
nor U1895 (N_1895,N_1249,N_839);
nor U1896 (N_1896,N_760,N_1040);
and U1897 (N_1897,N_1119,N_1123);
nand U1898 (N_1898,N_1060,N_860);
xor U1899 (N_1899,N_1164,N_1385);
and U1900 (N_1900,N_982,N_920);
and U1901 (N_1901,N_1366,N_1424);
nand U1902 (N_1902,N_755,N_958);
nor U1903 (N_1903,N_1142,N_990);
nand U1904 (N_1904,N_1240,N_1434);
nor U1905 (N_1905,N_767,N_1298);
nand U1906 (N_1906,N_872,N_1290);
nand U1907 (N_1907,N_1370,N_803);
or U1908 (N_1908,N_1486,N_1312);
and U1909 (N_1909,N_1328,N_1341);
and U1910 (N_1910,N_941,N_1136);
nor U1911 (N_1911,N_766,N_1040);
or U1912 (N_1912,N_1326,N_991);
nor U1913 (N_1913,N_816,N_1386);
nand U1914 (N_1914,N_1127,N_1033);
nor U1915 (N_1915,N_872,N_1251);
and U1916 (N_1916,N_1232,N_1060);
nor U1917 (N_1917,N_813,N_950);
or U1918 (N_1918,N_927,N_1101);
or U1919 (N_1919,N_944,N_978);
and U1920 (N_1920,N_1131,N_1263);
nand U1921 (N_1921,N_1182,N_974);
or U1922 (N_1922,N_1464,N_900);
or U1923 (N_1923,N_1246,N_1390);
nand U1924 (N_1924,N_1324,N_1001);
or U1925 (N_1925,N_797,N_934);
nor U1926 (N_1926,N_1491,N_1139);
nand U1927 (N_1927,N_762,N_978);
and U1928 (N_1928,N_1149,N_1196);
or U1929 (N_1929,N_922,N_885);
nand U1930 (N_1930,N_1391,N_1415);
and U1931 (N_1931,N_1205,N_827);
or U1932 (N_1932,N_1365,N_981);
nor U1933 (N_1933,N_1453,N_1243);
nor U1934 (N_1934,N_890,N_1162);
nand U1935 (N_1935,N_771,N_1400);
or U1936 (N_1936,N_1493,N_1469);
nand U1937 (N_1937,N_787,N_1261);
or U1938 (N_1938,N_1463,N_1049);
nor U1939 (N_1939,N_1280,N_1023);
nor U1940 (N_1940,N_1292,N_1319);
nor U1941 (N_1941,N_1064,N_1469);
nand U1942 (N_1942,N_1361,N_1371);
and U1943 (N_1943,N_1491,N_1296);
nand U1944 (N_1944,N_796,N_1169);
nand U1945 (N_1945,N_1129,N_1453);
nor U1946 (N_1946,N_1174,N_825);
nand U1947 (N_1947,N_935,N_944);
nand U1948 (N_1948,N_1441,N_1421);
and U1949 (N_1949,N_975,N_1100);
nand U1950 (N_1950,N_806,N_1048);
and U1951 (N_1951,N_1369,N_1009);
and U1952 (N_1952,N_1084,N_1251);
nor U1953 (N_1953,N_1309,N_853);
and U1954 (N_1954,N_765,N_1086);
nor U1955 (N_1955,N_1212,N_1369);
nor U1956 (N_1956,N_1065,N_1182);
and U1957 (N_1957,N_1344,N_920);
and U1958 (N_1958,N_1473,N_765);
and U1959 (N_1959,N_887,N_972);
and U1960 (N_1960,N_978,N_1424);
or U1961 (N_1961,N_867,N_1096);
or U1962 (N_1962,N_784,N_1303);
nand U1963 (N_1963,N_1455,N_955);
and U1964 (N_1964,N_1117,N_1409);
and U1965 (N_1965,N_1432,N_857);
and U1966 (N_1966,N_1296,N_992);
nand U1967 (N_1967,N_944,N_938);
nand U1968 (N_1968,N_791,N_1468);
nand U1969 (N_1969,N_1213,N_1250);
or U1970 (N_1970,N_816,N_1109);
or U1971 (N_1971,N_1214,N_1341);
nor U1972 (N_1972,N_1216,N_1297);
or U1973 (N_1973,N_858,N_1415);
nand U1974 (N_1974,N_1110,N_1031);
nor U1975 (N_1975,N_1496,N_1444);
nor U1976 (N_1976,N_908,N_1006);
nand U1977 (N_1977,N_1174,N_870);
nand U1978 (N_1978,N_844,N_1107);
nor U1979 (N_1979,N_1112,N_1102);
nand U1980 (N_1980,N_987,N_1299);
and U1981 (N_1981,N_809,N_1357);
nor U1982 (N_1982,N_1495,N_1053);
nor U1983 (N_1983,N_979,N_1074);
and U1984 (N_1984,N_1366,N_1092);
and U1985 (N_1985,N_1102,N_975);
nand U1986 (N_1986,N_1270,N_793);
xor U1987 (N_1987,N_856,N_1197);
or U1988 (N_1988,N_1408,N_1446);
or U1989 (N_1989,N_1313,N_920);
nor U1990 (N_1990,N_825,N_1300);
or U1991 (N_1991,N_905,N_1245);
nand U1992 (N_1992,N_1097,N_1151);
or U1993 (N_1993,N_1228,N_1451);
nand U1994 (N_1994,N_1123,N_1221);
and U1995 (N_1995,N_1372,N_1388);
and U1996 (N_1996,N_1396,N_1457);
and U1997 (N_1997,N_969,N_866);
and U1998 (N_1998,N_944,N_1322);
or U1999 (N_1999,N_1002,N_1231);
and U2000 (N_2000,N_1418,N_814);
or U2001 (N_2001,N_804,N_1458);
nand U2002 (N_2002,N_1205,N_781);
or U2003 (N_2003,N_1202,N_1112);
and U2004 (N_2004,N_1478,N_1372);
nor U2005 (N_2005,N_1109,N_1450);
or U2006 (N_2006,N_1117,N_778);
and U2007 (N_2007,N_1066,N_1273);
or U2008 (N_2008,N_946,N_1129);
nor U2009 (N_2009,N_987,N_953);
or U2010 (N_2010,N_781,N_997);
nand U2011 (N_2011,N_949,N_830);
nor U2012 (N_2012,N_789,N_1237);
and U2013 (N_2013,N_1243,N_940);
and U2014 (N_2014,N_1406,N_1195);
or U2015 (N_2015,N_798,N_1039);
or U2016 (N_2016,N_883,N_964);
nand U2017 (N_2017,N_970,N_1366);
nand U2018 (N_2018,N_1298,N_1258);
nand U2019 (N_2019,N_1378,N_1021);
nand U2020 (N_2020,N_1021,N_1292);
nor U2021 (N_2021,N_1098,N_1057);
or U2022 (N_2022,N_990,N_1313);
nor U2023 (N_2023,N_928,N_1036);
nor U2024 (N_2024,N_885,N_1423);
nand U2025 (N_2025,N_794,N_1490);
or U2026 (N_2026,N_1382,N_809);
or U2027 (N_2027,N_925,N_870);
or U2028 (N_2028,N_928,N_1358);
and U2029 (N_2029,N_1005,N_998);
or U2030 (N_2030,N_1424,N_774);
and U2031 (N_2031,N_1342,N_1307);
and U2032 (N_2032,N_835,N_1236);
or U2033 (N_2033,N_1396,N_897);
nand U2034 (N_2034,N_1495,N_1134);
nor U2035 (N_2035,N_910,N_1171);
nand U2036 (N_2036,N_927,N_891);
or U2037 (N_2037,N_1130,N_781);
or U2038 (N_2038,N_1185,N_1205);
nor U2039 (N_2039,N_1358,N_1306);
nor U2040 (N_2040,N_1476,N_1048);
nor U2041 (N_2041,N_1064,N_1059);
nor U2042 (N_2042,N_1068,N_984);
nand U2043 (N_2043,N_1105,N_1317);
or U2044 (N_2044,N_1037,N_1475);
or U2045 (N_2045,N_1203,N_1431);
nor U2046 (N_2046,N_1344,N_940);
or U2047 (N_2047,N_1183,N_1422);
and U2048 (N_2048,N_1046,N_835);
or U2049 (N_2049,N_795,N_867);
nor U2050 (N_2050,N_855,N_817);
nand U2051 (N_2051,N_1400,N_1263);
and U2052 (N_2052,N_1463,N_845);
nor U2053 (N_2053,N_1479,N_1294);
and U2054 (N_2054,N_1318,N_1048);
or U2055 (N_2055,N_882,N_1225);
or U2056 (N_2056,N_1491,N_1466);
nor U2057 (N_2057,N_1212,N_1478);
and U2058 (N_2058,N_1247,N_1131);
nand U2059 (N_2059,N_949,N_1038);
nor U2060 (N_2060,N_1157,N_786);
nand U2061 (N_2061,N_1268,N_1092);
nand U2062 (N_2062,N_1409,N_1464);
or U2063 (N_2063,N_1166,N_1217);
and U2064 (N_2064,N_879,N_1123);
nor U2065 (N_2065,N_1479,N_1458);
nand U2066 (N_2066,N_1173,N_1275);
and U2067 (N_2067,N_987,N_856);
nor U2068 (N_2068,N_1415,N_1293);
and U2069 (N_2069,N_787,N_1060);
or U2070 (N_2070,N_763,N_1444);
nor U2071 (N_2071,N_841,N_1281);
and U2072 (N_2072,N_1106,N_861);
or U2073 (N_2073,N_1148,N_1393);
nand U2074 (N_2074,N_915,N_1234);
and U2075 (N_2075,N_953,N_1121);
nand U2076 (N_2076,N_1258,N_1414);
or U2077 (N_2077,N_1224,N_872);
nand U2078 (N_2078,N_1040,N_1267);
nand U2079 (N_2079,N_1468,N_903);
or U2080 (N_2080,N_965,N_1329);
or U2081 (N_2081,N_888,N_1083);
and U2082 (N_2082,N_1437,N_1484);
and U2083 (N_2083,N_1335,N_1049);
nand U2084 (N_2084,N_791,N_1017);
nor U2085 (N_2085,N_955,N_1432);
and U2086 (N_2086,N_977,N_1032);
or U2087 (N_2087,N_1451,N_1215);
or U2088 (N_2088,N_1273,N_1163);
and U2089 (N_2089,N_1216,N_1325);
nor U2090 (N_2090,N_791,N_1061);
and U2091 (N_2091,N_977,N_1048);
nor U2092 (N_2092,N_1268,N_1376);
nor U2093 (N_2093,N_1486,N_1175);
nand U2094 (N_2094,N_893,N_1090);
nand U2095 (N_2095,N_1196,N_1361);
or U2096 (N_2096,N_1176,N_1473);
nor U2097 (N_2097,N_1071,N_1039);
and U2098 (N_2098,N_826,N_899);
nor U2099 (N_2099,N_982,N_959);
nor U2100 (N_2100,N_1118,N_1009);
nand U2101 (N_2101,N_1233,N_1276);
or U2102 (N_2102,N_877,N_1074);
or U2103 (N_2103,N_791,N_1469);
nor U2104 (N_2104,N_1201,N_804);
nor U2105 (N_2105,N_910,N_991);
nand U2106 (N_2106,N_1451,N_1329);
nor U2107 (N_2107,N_1123,N_834);
nand U2108 (N_2108,N_1294,N_1305);
nand U2109 (N_2109,N_1096,N_1288);
nor U2110 (N_2110,N_813,N_1493);
nor U2111 (N_2111,N_1407,N_959);
or U2112 (N_2112,N_1138,N_1245);
nor U2113 (N_2113,N_1319,N_1154);
nand U2114 (N_2114,N_927,N_1406);
nand U2115 (N_2115,N_1161,N_1233);
or U2116 (N_2116,N_1102,N_1488);
or U2117 (N_2117,N_1425,N_1139);
nor U2118 (N_2118,N_830,N_874);
and U2119 (N_2119,N_989,N_1121);
nor U2120 (N_2120,N_852,N_780);
nand U2121 (N_2121,N_1387,N_1447);
or U2122 (N_2122,N_1159,N_1279);
nor U2123 (N_2123,N_1007,N_1383);
and U2124 (N_2124,N_1444,N_840);
nor U2125 (N_2125,N_1145,N_813);
and U2126 (N_2126,N_935,N_936);
nor U2127 (N_2127,N_1387,N_1093);
or U2128 (N_2128,N_1196,N_1031);
and U2129 (N_2129,N_760,N_1173);
or U2130 (N_2130,N_760,N_1045);
and U2131 (N_2131,N_1225,N_1079);
nand U2132 (N_2132,N_1051,N_908);
or U2133 (N_2133,N_900,N_763);
or U2134 (N_2134,N_825,N_1387);
nand U2135 (N_2135,N_1309,N_1143);
nor U2136 (N_2136,N_1431,N_1489);
or U2137 (N_2137,N_971,N_973);
nand U2138 (N_2138,N_864,N_1124);
nand U2139 (N_2139,N_1257,N_1480);
or U2140 (N_2140,N_1341,N_796);
nand U2141 (N_2141,N_1105,N_1276);
nor U2142 (N_2142,N_1057,N_1490);
and U2143 (N_2143,N_1296,N_862);
and U2144 (N_2144,N_987,N_792);
and U2145 (N_2145,N_891,N_776);
and U2146 (N_2146,N_1135,N_1343);
nand U2147 (N_2147,N_1147,N_1070);
and U2148 (N_2148,N_925,N_812);
and U2149 (N_2149,N_951,N_919);
and U2150 (N_2150,N_1322,N_1206);
nor U2151 (N_2151,N_1189,N_1088);
nand U2152 (N_2152,N_1262,N_1234);
nand U2153 (N_2153,N_1372,N_1475);
and U2154 (N_2154,N_1313,N_976);
nor U2155 (N_2155,N_1387,N_800);
nand U2156 (N_2156,N_1310,N_1285);
nor U2157 (N_2157,N_1319,N_1297);
and U2158 (N_2158,N_829,N_795);
nand U2159 (N_2159,N_979,N_1316);
nand U2160 (N_2160,N_1382,N_821);
or U2161 (N_2161,N_1220,N_874);
nand U2162 (N_2162,N_1428,N_789);
nand U2163 (N_2163,N_1217,N_1247);
nor U2164 (N_2164,N_1105,N_1309);
or U2165 (N_2165,N_1099,N_1080);
or U2166 (N_2166,N_1396,N_1363);
or U2167 (N_2167,N_1290,N_1223);
nand U2168 (N_2168,N_850,N_1071);
and U2169 (N_2169,N_1079,N_1288);
nand U2170 (N_2170,N_912,N_1277);
and U2171 (N_2171,N_1016,N_1201);
or U2172 (N_2172,N_825,N_1027);
nor U2173 (N_2173,N_1285,N_1248);
nand U2174 (N_2174,N_925,N_1496);
nor U2175 (N_2175,N_988,N_1060);
or U2176 (N_2176,N_1037,N_1232);
or U2177 (N_2177,N_1417,N_1112);
and U2178 (N_2178,N_1443,N_1312);
or U2179 (N_2179,N_1074,N_1239);
and U2180 (N_2180,N_1051,N_862);
and U2181 (N_2181,N_916,N_1373);
and U2182 (N_2182,N_1459,N_780);
or U2183 (N_2183,N_1229,N_1013);
nand U2184 (N_2184,N_1383,N_1294);
and U2185 (N_2185,N_1407,N_1180);
nand U2186 (N_2186,N_1117,N_1152);
or U2187 (N_2187,N_1113,N_863);
or U2188 (N_2188,N_1440,N_1303);
nor U2189 (N_2189,N_991,N_796);
and U2190 (N_2190,N_850,N_931);
or U2191 (N_2191,N_1196,N_781);
nor U2192 (N_2192,N_1002,N_760);
nor U2193 (N_2193,N_823,N_910);
and U2194 (N_2194,N_994,N_1146);
and U2195 (N_2195,N_1195,N_779);
nor U2196 (N_2196,N_838,N_1307);
nor U2197 (N_2197,N_953,N_1305);
xor U2198 (N_2198,N_1442,N_953);
and U2199 (N_2199,N_781,N_1233);
and U2200 (N_2200,N_888,N_1241);
nand U2201 (N_2201,N_1145,N_1172);
xnor U2202 (N_2202,N_793,N_1359);
nor U2203 (N_2203,N_1173,N_1434);
or U2204 (N_2204,N_1309,N_1347);
nor U2205 (N_2205,N_1261,N_1461);
nand U2206 (N_2206,N_753,N_1342);
or U2207 (N_2207,N_846,N_1348);
nor U2208 (N_2208,N_1287,N_977);
and U2209 (N_2209,N_1258,N_1306);
or U2210 (N_2210,N_987,N_801);
nor U2211 (N_2211,N_802,N_1405);
nor U2212 (N_2212,N_1380,N_873);
nand U2213 (N_2213,N_870,N_1135);
and U2214 (N_2214,N_1385,N_1001);
or U2215 (N_2215,N_1166,N_1128);
nor U2216 (N_2216,N_1490,N_1207);
and U2217 (N_2217,N_1389,N_1175);
and U2218 (N_2218,N_1356,N_1488);
and U2219 (N_2219,N_1175,N_947);
or U2220 (N_2220,N_885,N_1382);
or U2221 (N_2221,N_1372,N_1415);
and U2222 (N_2222,N_781,N_1448);
or U2223 (N_2223,N_1262,N_862);
and U2224 (N_2224,N_1195,N_1024);
and U2225 (N_2225,N_989,N_797);
nand U2226 (N_2226,N_1078,N_1107);
nor U2227 (N_2227,N_1212,N_1161);
xor U2228 (N_2228,N_1392,N_769);
or U2229 (N_2229,N_1347,N_1278);
or U2230 (N_2230,N_1036,N_1300);
and U2231 (N_2231,N_1469,N_884);
and U2232 (N_2232,N_1064,N_783);
or U2233 (N_2233,N_1044,N_1272);
and U2234 (N_2234,N_1179,N_1160);
and U2235 (N_2235,N_1374,N_1492);
or U2236 (N_2236,N_1014,N_1455);
and U2237 (N_2237,N_1280,N_1042);
or U2238 (N_2238,N_1182,N_1397);
and U2239 (N_2239,N_1256,N_1172);
or U2240 (N_2240,N_1477,N_963);
nand U2241 (N_2241,N_1213,N_872);
nand U2242 (N_2242,N_802,N_842);
nor U2243 (N_2243,N_1411,N_1152);
nand U2244 (N_2244,N_1344,N_1243);
or U2245 (N_2245,N_942,N_1058);
or U2246 (N_2246,N_1245,N_1151);
nor U2247 (N_2247,N_1396,N_819);
or U2248 (N_2248,N_937,N_1243);
and U2249 (N_2249,N_1077,N_1235);
or U2250 (N_2250,N_2106,N_1999);
nor U2251 (N_2251,N_1760,N_1838);
or U2252 (N_2252,N_1706,N_2189);
nor U2253 (N_2253,N_2094,N_1744);
and U2254 (N_2254,N_1717,N_1572);
xor U2255 (N_2255,N_2028,N_1930);
nand U2256 (N_2256,N_2167,N_1877);
nand U2257 (N_2257,N_1563,N_2135);
and U2258 (N_2258,N_2101,N_1737);
or U2259 (N_2259,N_1536,N_1643);
or U2260 (N_2260,N_1668,N_1519);
and U2261 (N_2261,N_1538,N_1855);
nor U2262 (N_2262,N_1761,N_1607);
and U2263 (N_2263,N_1810,N_2129);
nand U2264 (N_2264,N_1879,N_1615);
or U2265 (N_2265,N_2116,N_1714);
nor U2266 (N_2266,N_2209,N_2126);
nand U2267 (N_2267,N_2032,N_1638);
nand U2268 (N_2268,N_1500,N_2082);
nand U2269 (N_2269,N_1866,N_1790);
and U2270 (N_2270,N_2013,N_1829);
or U2271 (N_2271,N_1949,N_2067);
and U2272 (N_2272,N_1974,N_1680);
or U2273 (N_2273,N_1520,N_1653);
nor U2274 (N_2274,N_1694,N_1822);
nor U2275 (N_2275,N_2198,N_1891);
and U2276 (N_2276,N_2138,N_1530);
nand U2277 (N_2277,N_1881,N_1735);
nand U2278 (N_2278,N_1874,N_1675);
and U2279 (N_2279,N_1647,N_1656);
and U2280 (N_2280,N_2027,N_1590);
or U2281 (N_2281,N_1834,N_1780);
or U2282 (N_2282,N_2145,N_1669);
nand U2283 (N_2283,N_2016,N_2071);
nor U2284 (N_2284,N_2150,N_1682);
nor U2285 (N_2285,N_2085,N_1807);
and U2286 (N_2286,N_1942,N_1716);
nor U2287 (N_2287,N_2022,N_2151);
nor U2288 (N_2288,N_1920,N_1571);
and U2289 (N_2289,N_1599,N_1612);
xor U2290 (N_2290,N_2007,N_1894);
nand U2291 (N_2291,N_1733,N_1658);
and U2292 (N_2292,N_1922,N_1748);
or U2293 (N_2293,N_1973,N_1712);
and U2294 (N_2294,N_2225,N_1814);
or U2295 (N_2295,N_1606,N_1614);
nand U2296 (N_2296,N_2224,N_1932);
nor U2297 (N_2297,N_1642,N_1598);
or U2298 (N_2298,N_1856,N_2204);
or U2299 (N_2299,N_2235,N_1657);
or U2300 (N_2300,N_1763,N_1904);
nor U2301 (N_2301,N_1961,N_1788);
nor U2302 (N_2302,N_1512,N_1539);
nand U2303 (N_2303,N_1911,N_1965);
nand U2304 (N_2304,N_2112,N_2055);
nand U2305 (N_2305,N_1857,N_2045);
nor U2306 (N_2306,N_2023,N_1581);
and U2307 (N_2307,N_2088,N_1947);
and U2308 (N_2308,N_1799,N_1683);
nand U2309 (N_2309,N_1787,N_1910);
and U2310 (N_2310,N_1559,N_2195);
or U2311 (N_2311,N_2025,N_1805);
or U2312 (N_2312,N_1724,N_1764);
nor U2313 (N_2313,N_1871,N_1673);
nor U2314 (N_2314,N_2118,N_1986);
xnor U2315 (N_2315,N_1943,N_1725);
and U2316 (N_2316,N_2048,N_1644);
and U2317 (N_2317,N_2131,N_1765);
nor U2318 (N_2318,N_1975,N_1603);
and U2319 (N_2319,N_1864,N_1586);
and U2320 (N_2320,N_1867,N_2015);
and U2321 (N_2321,N_1854,N_1844);
or U2322 (N_2322,N_1645,N_2220);
nor U2323 (N_2323,N_1613,N_1742);
or U2324 (N_2324,N_1508,N_2169);
nor U2325 (N_2325,N_2218,N_1623);
or U2326 (N_2326,N_1621,N_1897);
or U2327 (N_2327,N_1575,N_1823);
and U2328 (N_2328,N_1831,N_2184);
xnor U2329 (N_2329,N_1749,N_1596);
nand U2330 (N_2330,N_1727,N_1704);
nor U2331 (N_2331,N_1967,N_2115);
nand U2332 (N_2332,N_2199,N_2047);
nor U2333 (N_2333,N_1789,N_2190);
nand U2334 (N_2334,N_1962,N_1913);
nand U2335 (N_2335,N_1858,N_1954);
and U2336 (N_2336,N_2057,N_1970);
nor U2337 (N_2337,N_1531,N_2114);
nand U2338 (N_2338,N_1779,N_2091);
nand U2339 (N_2339,N_2104,N_1522);
or U2340 (N_2340,N_1501,N_1887);
or U2341 (N_2341,N_2072,N_1718);
nand U2342 (N_2342,N_1688,N_1702);
nand U2343 (N_2343,N_1795,N_1602);
and U2344 (N_2344,N_1786,N_1849);
nor U2345 (N_2345,N_1580,N_1859);
nor U2346 (N_2346,N_2246,N_2083);
nor U2347 (N_2347,N_1915,N_1529);
and U2348 (N_2348,N_1958,N_1720);
nor U2349 (N_2349,N_2039,N_2242);
nand U2350 (N_2350,N_1811,N_2044);
nor U2351 (N_2351,N_1593,N_2056);
or U2352 (N_2352,N_2130,N_1983);
and U2353 (N_2353,N_1626,N_1755);
nor U2354 (N_2354,N_1848,N_1818);
and U2355 (N_2355,N_1729,N_1561);
and U2356 (N_2356,N_2205,N_1558);
and U2357 (N_2357,N_1707,N_1698);
nor U2358 (N_2358,N_2035,N_1541);
nand U2359 (N_2359,N_2000,N_1711);
or U2360 (N_2360,N_2139,N_1825);
nand U2361 (N_2361,N_2086,N_2160);
or U2362 (N_2362,N_2233,N_1762);
nor U2363 (N_2363,N_2073,N_2049);
xor U2364 (N_2364,N_1641,N_2024);
nand U2365 (N_2365,N_2146,N_2148);
and U2366 (N_2366,N_1952,N_1792);
nor U2367 (N_2367,N_1994,N_1595);
nand U2368 (N_2368,N_1671,N_2058);
nand U2369 (N_2369,N_1991,N_1842);
nand U2370 (N_2370,N_1525,N_1701);
or U2371 (N_2371,N_2120,N_2134);
nand U2372 (N_2372,N_1912,N_2002);
nor U2373 (N_2373,N_1752,N_2046);
nand U2374 (N_2374,N_1837,N_1797);
nor U2375 (N_2375,N_1544,N_2176);
nor U2376 (N_2376,N_1997,N_1537);
or U2377 (N_2377,N_1921,N_2125);
nand U2378 (N_2378,N_2227,N_2143);
nor U2379 (N_2379,N_1532,N_2226);
and U2380 (N_2380,N_2201,N_2231);
or U2381 (N_2381,N_2156,N_1776);
nand U2382 (N_2382,N_1995,N_2163);
and U2383 (N_2383,N_1827,N_1906);
nor U2384 (N_2384,N_1568,N_1747);
nor U2385 (N_2385,N_2200,N_2228);
and U2386 (N_2386,N_1664,N_1988);
nor U2387 (N_2387,N_2078,N_1506);
or U2388 (N_2388,N_1772,N_1916);
and U2389 (N_2389,N_1778,N_1959);
or U2390 (N_2390,N_2215,N_1660);
or U2391 (N_2391,N_1869,N_1710);
nand U2392 (N_2392,N_1734,N_2018);
nand U2393 (N_2393,N_1739,N_2140);
or U2394 (N_2394,N_1515,N_1627);
nor U2395 (N_2395,N_1969,N_2216);
nand U2396 (N_2396,N_2026,N_1582);
or U2397 (N_2397,N_1608,N_1819);
and U2398 (N_2398,N_1948,N_1862);
nand U2399 (N_2399,N_2004,N_1803);
and U2400 (N_2400,N_1721,N_2191);
and U2401 (N_2401,N_1557,N_1631);
nand U2402 (N_2402,N_2095,N_2068);
nor U2403 (N_2403,N_1513,N_1726);
nor U2404 (N_2404,N_2113,N_1655);
nand U2405 (N_2405,N_2092,N_1567);
and U2406 (N_2406,N_1960,N_2149);
nand U2407 (N_2407,N_1956,N_1985);
or U2408 (N_2408,N_1528,N_2075);
and U2409 (N_2409,N_1774,N_2234);
and U2410 (N_2410,N_2108,N_1800);
or U2411 (N_2411,N_1944,N_1992);
and U2412 (N_2412,N_2237,N_1950);
or U2413 (N_2413,N_1663,N_2232);
or U2414 (N_2414,N_2196,N_1628);
or U2415 (N_2415,N_1941,N_2171);
nand U2416 (N_2416,N_1928,N_1521);
and U2417 (N_2417,N_2157,N_2051);
and U2418 (N_2418,N_1903,N_1900);
and U2419 (N_2419,N_1611,N_2203);
nand U2420 (N_2420,N_1868,N_1832);
nor U2421 (N_2421,N_2074,N_1979);
or U2422 (N_2422,N_1955,N_1684);
or U2423 (N_2423,N_1546,N_2192);
nor U2424 (N_2424,N_1987,N_1890);
and U2425 (N_2425,N_1968,N_1951);
and U2426 (N_2426,N_1886,N_1732);
or U2427 (N_2427,N_2170,N_1873);
or U2428 (N_2428,N_2248,N_1980);
or U2429 (N_2429,N_1649,N_1610);
and U2430 (N_2430,N_2168,N_1750);
nor U2431 (N_2431,N_1622,N_2179);
nand U2432 (N_2432,N_1978,N_1852);
nor U2433 (N_2433,N_1888,N_1933);
or U2434 (N_2434,N_1518,N_1667);
nor U2435 (N_2435,N_2202,N_1882);
or U2436 (N_2436,N_2152,N_1579);
or U2437 (N_2437,N_2065,N_1830);
or U2438 (N_2438,N_1545,N_1836);
nand U2439 (N_2439,N_1594,N_1556);
nand U2440 (N_2440,N_1976,N_1796);
and U2441 (N_2441,N_2102,N_2037);
nand U2442 (N_2442,N_2137,N_1619);
and U2443 (N_2443,N_2211,N_1835);
and U2444 (N_2444,N_2177,N_2142);
and U2445 (N_2445,N_1768,N_1700);
nor U2446 (N_2446,N_2033,N_1632);
nand U2447 (N_2447,N_1981,N_1597);
nor U2448 (N_2448,N_2063,N_1826);
nand U2449 (N_2449,N_1821,N_2119);
or U2450 (N_2450,N_1996,N_1770);
or U2451 (N_2451,N_1926,N_1816);
or U2452 (N_2452,N_1804,N_2001);
or U2453 (N_2453,N_1989,N_2124);
nor U2454 (N_2454,N_1679,N_2080);
or U2455 (N_2455,N_1570,N_1865);
nand U2456 (N_2456,N_2011,N_1773);
nor U2457 (N_2457,N_2123,N_1901);
nor U2458 (N_2458,N_2188,N_2197);
or U2459 (N_2459,N_1708,N_1808);
nand U2460 (N_2460,N_2219,N_1629);
and U2461 (N_2461,N_1802,N_1990);
and U2462 (N_2462,N_1840,N_1939);
nand U2463 (N_2463,N_2081,N_1691);
nand U2464 (N_2464,N_1534,N_2208);
nand U2465 (N_2465,N_1713,N_1757);
nor U2466 (N_2466,N_1678,N_1977);
nand U2467 (N_2467,N_1782,N_1817);
nor U2468 (N_2468,N_2052,N_2110);
nor U2469 (N_2469,N_1535,N_1845);
nor U2470 (N_2470,N_2008,N_2229);
nand U2471 (N_2471,N_2042,N_1919);
nand U2472 (N_2472,N_1692,N_1934);
nand U2473 (N_2473,N_1651,N_1553);
xor U2474 (N_2474,N_1516,N_1741);
nand U2475 (N_2475,N_1982,N_1935);
nor U2476 (N_2476,N_1524,N_1861);
or U2477 (N_2477,N_1895,N_2147);
and U2478 (N_2478,N_1775,N_1709);
nand U2479 (N_2479,N_1847,N_2247);
nor U2480 (N_2480,N_1543,N_1870);
or U2481 (N_2481,N_2061,N_2241);
or U2482 (N_2482,N_2165,N_2133);
nand U2483 (N_2483,N_2117,N_2240);
and U2484 (N_2484,N_2207,N_2193);
and U2485 (N_2485,N_2183,N_1555);
nand U2486 (N_2486,N_1853,N_2021);
xnor U2487 (N_2487,N_1578,N_2030);
nor U2488 (N_2488,N_2214,N_1533);
nand U2489 (N_2489,N_2144,N_1504);
or U2490 (N_2490,N_2164,N_1938);
or U2491 (N_2491,N_2069,N_1617);
and U2492 (N_2492,N_1604,N_2019);
or U2493 (N_2493,N_1601,N_1646);
or U2494 (N_2494,N_1918,N_1892);
nor U2495 (N_2495,N_2161,N_2238);
nand U2496 (N_2496,N_1662,N_1514);
nor U2497 (N_2497,N_2187,N_2141);
and U2498 (N_2498,N_1542,N_2173);
or U2499 (N_2499,N_1640,N_1931);
and U2500 (N_2500,N_2111,N_2159);
and U2501 (N_2501,N_2174,N_1589);
and U2502 (N_2502,N_1588,N_1730);
and U2503 (N_2503,N_1677,N_1562);
or U2504 (N_2504,N_1722,N_2090);
nand U2505 (N_2505,N_1794,N_2212);
nand U2506 (N_2506,N_2185,N_2121);
and U2507 (N_2507,N_2038,N_2132);
nor U2508 (N_2508,N_1812,N_1957);
nand U2509 (N_2509,N_1509,N_1876);
nand U2510 (N_2510,N_1899,N_2103);
nand U2511 (N_2511,N_1851,N_1753);
and U2512 (N_2512,N_1907,N_1585);
and U2513 (N_2513,N_2079,N_1674);
nand U2514 (N_2514,N_1652,N_2105);
nor U2515 (N_2515,N_1884,N_1693);
or U2516 (N_2516,N_2017,N_1548);
nand U2517 (N_2517,N_1863,N_2006);
nor U2518 (N_2518,N_1905,N_1909);
nand U2519 (N_2519,N_2206,N_1550);
nor U2520 (N_2520,N_1654,N_1695);
or U2521 (N_2521,N_2100,N_2236);
nand U2522 (N_2522,N_2036,N_1502);
or U2523 (N_2523,N_1777,N_1699);
and U2524 (N_2524,N_1625,N_1785);
or U2525 (N_2525,N_2158,N_1806);
nor U2526 (N_2526,N_1728,N_2230);
and U2527 (N_2527,N_2050,N_2180);
nor U2528 (N_2528,N_1738,N_2244);
nand U2529 (N_2529,N_2054,N_2098);
and U2530 (N_2530,N_2223,N_1689);
or U2531 (N_2531,N_2003,N_2239);
or U2532 (N_2532,N_2043,N_1756);
nand U2533 (N_2533,N_1705,N_1843);
and U2534 (N_2534,N_2222,N_1551);
nand U2535 (N_2535,N_1624,N_2099);
nand U2536 (N_2536,N_1784,N_2153);
xnor U2537 (N_2537,N_1526,N_1924);
or U2538 (N_2538,N_1583,N_1577);
and U2539 (N_2539,N_1875,N_1883);
nand U2540 (N_2540,N_2213,N_1659);
and U2541 (N_2541,N_1860,N_1833);
or U2542 (N_2542,N_2062,N_1940);
and U2543 (N_2543,N_1573,N_1552);
nand U2544 (N_2544,N_2076,N_1540);
or U2545 (N_2545,N_2009,N_1605);
nand U2546 (N_2546,N_1511,N_1554);
and U2547 (N_2547,N_1549,N_1839);
xor U2548 (N_2548,N_2128,N_1998);
nand U2549 (N_2549,N_2066,N_1685);
nor U2550 (N_2550,N_1743,N_1609);
nor U2551 (N_2551,N_1681,N_1719);
and U2552 (N_2552,N_2181,N_1616);
nor U2553 (N_2553,N_1824,N_1759);
nor U2554 (N_2554,N_1769,N_2154);
or U2555 (N_2555,N_1953,N_1591);
and U2556 (N_2556,N_2186,N_2107);
nor U2557 (N_2557,N_1766,N_1600);
or U2558 (N_2558,N_1569,N_1963);
or U2559 (N_2559,N_2182,N_1564);
nor U2560 (N_2560,N_2029,N_1917);
or U2561 (N_2561,N_1898,N_1925);
nor U2562 (N_2562,N_1620,N_1813);
or U2563 (N_2563,N_2059,N_1731);
nor U2564 (N_2564,N_1723,N_1793);
or U2565 (N_2565,N_1809,N_2041);
and U2566 (N_2566,N_2245,N_1878);
nor U2567 (N_2567,N_1984,N_2221);
or U2568 (N_2568,N_1560,N_2217);
nor U2569 (N_2569,N_1828,N_1503);
nand U2570 (N_2570,N_1880,N_1736);
or U2571 (N_2571,N_1574,N_1885);
nor U2572 (N_2572,N_1676,N_1771);
nor U2573 (N_2573,N_2053,N_1791);
or U2574 (N_2574,N_2175,N_1686);
nand U2575 (N_2575,N_1715,N_2194);
nand U2576 (N_2576,N_1618,N_2210);
nor U2577 (N_2577,N_1566,N_1576);
and U2578 (N_2578,N_2136,N_2155);
or U2579 (N_2579,N_1889,N_1507);
and U2580 (N_2580,N_1665,N_1767);
nor U2581 (N_2581,N_1637,N_2040);
and U2582 (N_2582,N_1820,N_2014);
and U2583 (N_2583,N_1697,N_1636);
nand U2584 (N_2584,N_2166,N_2089);
and U2585 (N_2585,N_1745,N_2077);
nand U2586 (N_2586,N_1815,N_1633);
or U2587 (N_2587,N_2084,N_1672);
nand U2588 (N_2588,N_1972,N_1929);
and U2589 (N_2589,N_2178,N_1893);
and U2590 (N_2590,N_1639,N_1592);
nor U2591 (N_2591,N_1850,N_2012);
or U2592 (N_2592,N_1971,N_1510);
nand U2593 (N_2593,N_2060,N_1666);
nand U2594 (N_2594,N_1758,N_1740);
nand U2595 (N_2595,N_2096,N_2172);
and U2596 (N_2596,N_1584,N_2243);
nand U2597 (N_2597,N_2034,N_1547);
and U2598 (N_2598,N_2249,N_1801);
nand U2599 (N_2599,N_1517,N_1670);
nand U2600 (N_2600,N_1798,N_2093);
or U2601 (N_2601,N_1993,N_1946);
nand U2602 (N_2602,N_1937,N_1696);
nor U2603 (N_2603,N_2010,N_1690);
or U2604 (N_2604,N_2070,N_1650);
nor U2605 (N_2605,N_2127,N_1914);
and U2606 (N_2606,N_1902,N_1523);
nor U2607 (N_2607,N_1565,N_1505);
and U2608 (N_2608,N_1841,N_1754);
and U2609 (N_2609,N_1927,N_1896);
or U2610 (N_2610,N_2020,N_1687);
nor U2611 (N_2611,N_1781,N_2064);
or U2612 (N_2612,N_1648,N_2122);
nor U2613 (N_2613,N_1703,N_1964);
or U2614 (N_2614,N_1527,N_2109);
nor U2615 (N_2615,N_1945,N_1846);
and U2616 (N_2616,N_1630,N_1746);
or U2617 (N_2617,N_1908,N_2097);
and U2618 (N_2618,N_1936,N_1783);
and U2619 (N_2619,N_1587,N_1661);
nand U2620 (N_2620,N_2005,N_1872);
and U2621 (N_2621,N_1634,N_1751);
or U2622 (N_2622,N_2162,N_2087);
nor U2623 (N_2623,N_1923,N_1635);
nor U2624 (N_2624,N_1966,N_2031);
and U2625 (N_2625,N_2222,N_1642);
or U2626 (N_2626,N_1544,N_1545);
and U2627 (N_2627,N_1651,N_2221);
or U2628 (N_2628,N_2031,N_1533);
nand U2629 (N_2629,N_2183,N_1892);
nand U2630 (N_2630,N_2068,N_1768);
and U2631 (N_2631,N_2007,N_1912);
and U2632 (N_2632,N_1657,N_1509);
nand U2633 (N_2633,N_2108,N_1900);
nand U2634 (N_2634,N_2127,N_2050);
or U2635 (N_2635,N_1641,N_1621);
nor U2636 (N_2636,N_1588,N_1781);
and U2637 (N_2637,N_2016,N_1782);
nand U2638 (N_2638,N_1523,N_1872);
and U2639 (N_2639,N_1578,N_1570);
nand U2640 (N_2640,N_2209,N_1540);
and U2641 (N_2641,N_1959,N_1857);
and U2642 (N_2642,N_1918,N_1509);
xor U2643 (N_2643,N_1727,N_1719);
or U2644 (N_2644,N_1981,N_1781);
or U2645 (N_2645,N_1858,N_1935);
nand U2646 (N_2646,N_2006,N_2173);
nor U2647 (N_2647,N_1611,N_2097);
and U2648 (N_2648,N_1970,N_1560);
and U2649 (N_2649,N_1733,N_2089);
nand U2650 (N_2650,N_1921,N_1674);
nand U2651 (N_2651,N_1815,N_1779);
and U2652 (N_2652,N_2133,N_1732);
nor U2653 (N_2653,N_1775,N_2074);
and U2654 (N_2654,N_1649,N_1599);
nand U2655 (N_2655,N_1877,N_1598);
nand U2656 (N_2656,N_1630,N_1970);
nor U2657 (N_2657,N_1835,N_1834);
or U2658 (N_2658,N_2182,N_1599);
nor U2659 (N_2659,N_1963,N_1748);
nor U2660 (N_2660,N_1694,N_1898);
nor U2661 (N_2661,N_2247,N_1848);
nor U2662 (N_2662,N_1862,N_1732);
and U2663 (N_2663,N_1905,N_2046);
or U2664 (N_2664,N_2030,N_1975);
and U2665 (N_2665,N_1738,N_1773);
nand U2666 (N_2666,N_2176,N_2114);
nor U2667 (N_2667,N_1858,N_1742);
nor U2668 (N_2668,N_2163,N_2089);
or U2669 (N_2669,N_2213,N_1501);
or U2670 (N_2670,N_1629,N_2155);
nand U2671 (N_2671,N_1657,N_2199);
or U2672 (N_2672,N_1718,N_2220);
nor U2673 (N_2673,N_1865,N_1510);
nand U2674 (N_2674,N_1894,N_1856);
or U2675 (N_2675,N_1849,N_1881);
and U2676 (N_2676,N_1809,N_1575);
and U2677 (N_2677,N_2170,N_1548);
and U2678 (N_2678,N_2195,N_2081);
or U2679 (N_2679,N_2059,N_1950);
nor U2680 (N_2680,N_1764,N_1772);
nor U2681 (N_2681,N_2198,N_2176);
xor U2682 (N_2682,N_1762,N_2242);
nand U2683 (N_2683,N_1893,N_1612);
nand U2684 (N_2684,N_1934,N_2086);
and U2685 (N_2685,N_1793,N_2182);
nor U2686 (N_2686,N_1870,N_1592);
and U2687 (N_2687,N_2242,N_1940);
nor U2688 (N_2688,N_1964,N_2055);
nand U2689 (N_2689,N_1711,N_1827);
and U2690 (N_2690,N_1730,N_2164);
nor U2691 (N_2691,N_1915,N_1627);
nor U2692 (N_2692,N_2014,N_1531);
or U2693 (N_2693,N_1842,N_1851);
and U2694 (N_2694,N_1803,N_2238);
nand U2695 (N_2695,N_2081,N_2199);
and U2696 (N_2696,N_2023,N_1572);
or U2697 (N_2697,N_1950,N_2123);
and U2698 (N_2698,N_1954,N_2087);
or U2699 (N_2699,N_1779,N_2101);
nand U2700 (N_2700,N_2200,N_2030);
nor U2701 (N_2701,N_1543,N_2144);
and U2702 (N_2702,N_1544,N_2012);
and U2703 (N_2703,N_1513,N_1728);
or U2704 (N_2704,N_2018,N_1521);
nand U2705 (N_2705,N_2156,N_1740);
and U2706 (N_2706,N_2143,N_1920);
nand U2707 (N_2707,N_1935,N_2058);
or U2708 (N_2708,N_1600,N_1996);
nor U2709 (N_2709,N_2025,N_1736);
nor U2710 (N_2710,N_1889,N_1979);
nor U2711 (N_2711,N_1561,N_1903);
and U2712 (N_2712,N_2155,N_2227);
nand U2713 (N_2713,N_2074,N_1657);
and U2714 (N_2714,N_1697,N_1802);
nor U2715 (N_2715,N_1532,N_1948);
or U2716 (N_2716,N_1924,N_1575);
and U2717 (N_2717,N_1838,N_2018);
or U2718 (N_2718,N_1695,N_1741);
nand U2719 (N_2719,N_1795,N_1580);
and U2720 (N_2720,N_1594,N_1522);
nor U2721 (N_2721,N_2137,N_2106);
or U2722 (N_2722,N_1559,N_2191);
nand U2723 (N_2723,N_2046,N_1636);
and U2724 (N_2724,N_2104,N_2158);
or U2725 (N_2725,N_1535,N_1545);
nor U2726 (N_2726,N_1695,N_1909);
and U2727 (N_2727,N_2060,N_1608);
nor U2728 (N_2728,N_1790,N_1599);
nand U2729 (N_2729,N_2027,N_2213);
nand U2730 (N_2730,N_1570,N_1600);
and U2731 (N_2731,N_2216,N_1712);
nand U2732 (N_2732,N_1930,N_2128);
or U2733 (N_2733,N_2037,N_1646);
and U2734 (N_2734,N_1594,N_1615);
xnor U2735 (N_2735,N_1526,N_1918);
and U2736 (N_2736,N_2238,N_1632);
nor U2737 (N_2737,N_1876,N_1685);
or U2738 (N_2738,N_2193,N_1817);
nand U2739 (N_2739,N_1717,N_2084);
and U2740 (N_2740,N_2072,N_1656);
nand U2741 (N_2741,N_1841,N_2248);
and U2742 (N_2742,N_2041,N_1727);
or U2743 (N_2743,N_2093,N_1657);
nor U2744 (N_2744,N_2155,N_1697);
or U2745 (N_2745,N_1871,N_1895);
or U2746 (N_2746,N_1606,N_2063);
nor U2747 (N_2747,N_1704,N_1802);
nor U2748 (N_2748,N_1854,N_1745);
and U2749 (N_2749,N_1765,N_1660);
and U2750 (N_2750,N_1521,N_1895);
and U2751 (N_2751,N_1904,N_2061);
or U2752 (N_2752,N_2237,N_1710);
or U2753 (N_2753,N_1589,N_1996);
and U2754 (N_2754,N_2150,N_1881);
and U2755 (N_2755,N_2131,N_1788);
nor U2756 (N_2756,N_1965,N_2030);
and U2757 (N_2757,N_1996,N_1637);
and U2758 (N_2758,N_1526,N_1997);
and U2759 (N_2759,N_2235,N_1638);
nand U2760 (N_2760,N_2210,N_1816);
nand U2761 (N_2761,N_2245,N_1679);
xnor U2762 (N_2762,N_2086,N_2185);
and U2763 (N_2763,N_1770,N_2066);
nand U2764 (N_2764,N_1926,N_1571);
and U2765 (N_2765,N_1971,N_1587);
and U2766 (N_2766,N_1640,N_2021);
nand U2767 (N_2767,N_1545,N_1738);
nor U2768 (N_2768,N_2215,N_2225);
nor U2769 (N_2769,N_1950,N_1845);
and U2770 (N_2770,N_2225,N_1978);
nor U2771 (N_2771,N_1872,N_1828);
and U2772 (N_2772,N_1765,N_2095);
or U2773 (N_2773,N_1727,N_1658);
and U2774 (N_2774,N_2079,N_2224);
or U2775 (N_2775,N_1821,N_1894);
nor U2776 (N_2776,N_2000,N_2207);
and U2777 (N_2777,N_1698,N_1711);
nor U2778 (N_2778,N_2054,N_1802);
nand U2779 (N_2779,N_2108,N_1723);
nor U2780 (N_2780,N_1962,N_2144);
and U2781 (N_2781,N_1948,N_1646);
nand U2782 (N_2782,N_1739,N_2053);
nand U2783 (N_2783,N_1973,N_1568);
or U2784 (N_2784,N_1838,N_1733);
or U2785 (N_2785,N_1942,N_1784);
and U2786 (N_2786,N_1548,N_2197);
and U2787 (N_2787,N_2107,N_2219);
or U2788 (N_2788,N_1604,N_1686);
nand U2789 (N_2789,N_1594,N_2041);
nand U2790 (N_2790,N_1990,N_2070);
or U2791 (N_2791,N_1672,N_2242);
nand U2792 (N_2792,N_1983,N_2152);
nor U2793 (N_2793,N_2069,N_1966);
nor U2794 (N_2794,N_1788,N_1884);
nand U2795 (N_2795,N_2106,N_1562);
and U2796 (N_2796,N_1580,N_1565);
nand U2797 (N_2797,N_1512,N_1773);
nand U2798 (N_2798,N_2127,N_2076);
or U2799 (N_2799,N_1617,N_2116);
or U2800 (N_2800,N_2202,N_2109);
nor U2801 (N_2801,N_2060,N_2133);
and U2802 (N_2802,N_1899,N_2040);
or U2803 (N_2803,N_2069,N_1714);
nor U2804 (N_2804,N_2001,N_1757);
or U2805 (N_2805,N_2027,N_1866);
nand U2806 (N_2806,N_2224,N_2204);
and U2807 (N_2807,N_2105,N_1827);
or U2808 (N_2808,N_2082,N_1640);
nor U2809 (N_2809,N_2185,N_1561);
or U2810 (N_2810,N_2015,N_1703);
nor U2811 (N_2811,N_1670,N_1613);
nor U2812 (N_2812,N_1999,N_2108);
or U2813 (N_2813,N_1989,N_2231);
xnor U2814 (N_2814,N_1767,N_2213);
and U2815 (N_2815,N_1835,N_1598);
nor U2816 (N_2816,N_1615,N_2189);
and U2817 (N_2817,N_1668,N_1620);
nor U2818 (N_2818,N_2205,N_1893);
or U2819 (N_2819,N_1729,N_1648);
or U2820 (N_2820,N_2046,N_1510);
nor U2821 (N_2821,N_2086,N_2000);
or U2822 (N_2822,N_1584,N_1968);
nand U2823 (N_2823,N_1695,N_1899);
and U2824 (N_2824,N_1879,N_1869);
nor U2825 (N_2825,N_1546,N_2238);
nand U2826 (N_2826,N_1606,N_2115);
nand U2827 (N_2827,N_1618,N_1778);
and U2828 (N_2828,N_2027,N_1990);
nor U2829 (N_2829,N_1670,N_2036);
nor U2830 (N_2830,N_1629,N_1635);
nor U2831 (N_2831,N_1826,N_1759);
nand U2832 (N_2832,N_2181,N_2170);
and U2833 (N_2833,N_1647,N_1661);
or U2834 (N_2834,N_1783,N_1691);
or U2835 (N_2835,N_2181,N_1702);
nand U2836 (N_2836,N_1785,N_2072);
nand U2837 (N_2837,N_1883,N_1873);
nor U2838 (N_2838,N_1813,N_1830);
nor U2839 (N_2839,N_2132,N_1823);
and U2840 (N_2840,N_2185,N_1792);
nand U2841 (N_2841,N_1530,N_1825);
and U2842 (N_2842,N_2111,N_1896);
or U2843 (N_2843,N_2155,N_1972);
or U2844 (N_2844,N_1960,N_2064);
nand U2845 (N_2845,N_1904,N_1600);
and U2846 (N_2846,N_1722,N_1559);
nor U2847 (N_2847,N_1584,N_1949);
nand U2848 (N_2848,N_1761,N_1733);
nand U2849 (N_2849,N_2074,N_2005);
nand U2850 (N_2850,N_1524,N_2201);
and U2851 (N_2851,N_1609,N_2245);
and U2852 (N_2852,N_1673,N_2128);
nor U2853 (N_2853,N_2086,N_1824);
nand U2854 (N_2854,N_1951,N_1840);
or U2855 (N_2855,N_2193,N_2127);
or U2856 (N_2856,N_1538,N_1974);
or U2857 (N_2857,N_1926,N_1563);
nand U2858 (N_2858,N_2228,N_1573);
or U2859 (N_2859,N_1570,N_1924);
and U2860 (N_2860,N_1552,N_1900);
xnor U2861 (N_2861,N_1614,N_1936);
and U2862 (N_2862,N_1908,N_2208);
and U2863 (N_2863,N_2158,N_1671);
and U2864 (N_2864,N_2034,N_1583);
and U2865 (N_2865,N_2117,N_2043);
nand U2866 (N_2866,N_1999,N_1597);
and U2867 (N_2867,N_1743,N_1582);
nand U2868 (N_2868,N_2083,N_1893);
nand U2869 (N_2869,N_2220,N_1746);
nor U2870 (N_2870,N_1624,N_1602);
and U2871 (N_2871,N_1863,N_1723);
and U2872 (N_2872,N_1809,N_2176);
and U2873 (N_2873,N_1928,N_1719);
and U2874 (N_2874,N_1947,N_1601);
nor U2875 (N_2875,N_1835,N_2038);
and U2876 (N_2876,N_2210,N_1967);
and U2877 (N_2877,N_2031,N_2003);
nor U2878 (N_2878,N_1849,N_1680);
and U2879 (N_2879,N_1965,N_1715);
nand U2880 (N_2880,N_1580,N_1568);
xnor U2881 (N_2881,N_1702,N_2001);
and U2882 (N_2882,N_2010,N_1978);
nor U2883 (N_2883,N_1877,N_1890);
nand U2884 (N_2884,N_1681,N_1808);
nand U2885 (N_2885,N_2162,N_1633);
nand U2886 (N_2886,N_1854,N_1605);
or U2887 (N_2887,N_2075,N_2024);
nor U2888 (N_2888,N_1600,N_2231);
and U2889 (N_2889,N_2022,N_1816);
and U2890 (N_2890,N_1963,N_2210);
and U2891 (N_2891,N_1861,N_2210);
nand U2892 (N_2892,N_1962,N_2006);
and U2893 (N_2893,N_2150,N_1717);
nand U2894 (N_2894,N_1838,N_1626);
or U2895 (N_2895,N_2202,N_2203);
nand U2896 (N_2896,N_1530,N_1817);
nor U2897 (N_2897,N_1580,N_1889);
nand U2898 (N_2898,N_1965,N_2115);
or U2899 (N_2899,N_1574,N_1954);
nor U2900 (N_2900,N_1757,N_1663);
or U2901 (N_2901,N_1529,N_1534);
and U2902 (N_2902,N_1744,N_1642);
nand U2903 (N_2903,N_2162,N_1715);
and U2904 (N_2904,N_1577,N_1604);
or U2905 (N_2905,N_1735,N_1579);
or U2906 (N_2906,N_1978,N_1596);
nor U2907 (N_2907,N_1605,N_2050);
nand U2908 (N_2908,N_2035,N_1708);
nor U2909 (N_2909,N_2094,N_1819);
nor U2910 (N_2910,N_2157,N_1735);
or U2911 (N_2911,N_1932,N_1775);
and U2912 (N_2912,N_1844,N_1550);
nor U2913 (N_2913,N_1741,N_1910);
or U2914 (N_2914,N_1990,N_1772);
and U2915 (N_2915,N_2038,N_1528);
or U2916 (N_2916,N_1506,N_1676);
nor U2917 (N_2917,N_1892,N_1765);
and U2918 (N_2918,N_1964,N_1741);
and U2919 (N_2919,N_2053,N_2095);
or U2920 (N_2920,N_2107,N_2240);
and U2921 (N_2921,N_1865,N_1726);
nor U2922 (N_2922,N_1717,N_1569);
and U2923 (N_2923,N_1712,N_1747);
nor U2924 (N_2924,N_2105,N_1574);
nand U2925 (N_2925,N_1769,N_2113);
nand U2926 (N_2926,N_2234,N_2124);
nor U2927 (N_2927,N_1691,N_1832);
nand U2928 (N_2928,N_1704,N_1987);
nand U2929 (N_2929,N_1819,N_1590);
nand U2930 (N_2930,N_1992,N_1975);
nand U2931 (N_2931,N_1670,N_1739);
and U2932 (N_2932,N_2017,N_2050);
nand U2933 (N_2933,N_1619,N_2113);
nor U2934 (N_2934,N_1950,N_1571);
and U2935 (N_2935,N_1687,N_1679);
nand U2936 (N_2936,N_1813,N_1695);
and U2937 (N_2937,N_2190,N_1815);
nor U2938 (N_2938,N_1977,N_2102);
and U2939 (N_2939,N_1910,N_2150);
and U2940 (N_2940,N_1619,N_1518);
and U2941 (N_2941,N_1855,N_1836);
nand U2942 (N_2942,N_2220,N_1976);
nor U2943 (N_2943,N_1880,N_2193);
and U2944 (N_2944,N_1909,N_1625);
or U2945 (N_2945,N_1725,N_1782);
nor U2946 (N_2946,N_1919,N_1789);
nor U2947 (N_2947,N_2245,N_1731);
nor U2948 (N_2948,N_2155,N_2147);
xor U2949 (N_2949,N_1815,N_2187);
or U2950 (N_2950,N_1757,N_1959);
nor U2951 (N_2951,N_1695,N_1661);
or U2952 (N_2952,N_1704,N_1619);
or U2953 (N_2953,N_1951,N_1640);
and U2954 (N_2954,N_1502,N_1859);
nand U2955 (N_2955,N_2208,N_1540);
or U2956 (N_2956,N_2016,N_1851);
or U2957 (N_2957,N_1997,N_1890);
and U2958 (N_2958,N_2124,N_2088);
nor U2959 (N_2959,N_1663,N_1683);
and U2960 (N_2960,N_2075,N_2126);
nand U2961 (N_2961,N_1654,N_2123);
or U2962 (N_2962,N_2174,N_2002);
and U2963 (N_2963,N_1940,N_2102);
nand U2964 (N_2964,N_1598,N_1660);
and U2965 (N_2965,N_2243,N_1781);
nor U2966 (N_2966,N_1960,N_1547);
and U2967 (N_2967,N_2128,N_2243);
nand U2968 (N_2968,N_1993,N_1767);
nand U2969 (N_2969,N_1856,N_1553);
nand U2970 (N_2970,N_2153,N_1777);
or U2971 (N_2971,N_1694,N_1745);
and U2972 (N_2972,N_2064,N_1819);
nand U2973 (N_2973,N_1983,N_2198);
or U2974 (N_2974,N_1719,N_1633);
nor U2975 (N_2975,N_1726,N_2112);
xor U2976 (N_2976,N_2173,N_1622);
nand U2977 (N_2977,N_1953,N_1721);
and U2978 (N_2978,N_2101,N_2227);
nor U2979 (N_2979,N_2040,N_1748);
or U2980 (N_2980,N_1568,N_1546);
xor U2981 (N_2981,N_1835,N_1785);
nand U2982 (N_2982,N_1658,N_2249);
nor U2983 (N_2983,N_1616,N_2163);
nor U2984 (N_2984,N_1879,N_2015);
nand U2985 (N_2985,N_1550,N_1667);
and U2986 (N_2986,N_2192,N_1562);
nor U2987 (N_2987,N_1940,N_1631);
nor U2988 (N_2988,N_1644,N_1679);
or U2989 (N_2989,N_1874,N_1633);
or U2990 (N_2990,N_1634,N_1960);
nor U2991 (N_2991,N_1566,N_2187);
or U2992 (N_2992,N_2122,N_1639);
and U2993 (N_2993,N_1656,N_2108);
and U2994 (N_2994,N_2144,N_1850);
nand U2995 (N_2995,N_2088,N_1734);
nand U2996 (N_2996,N_1940,N_2034);
nand U2997 (N_2997,N_1651,N_1630);
and U2998 (N_2998,N_2143,N_1945);
and U2999 (N_2999,N_1581,N_1511);
and UO_0 (O_0,N_2771,N_2668);
and UO_1 (O_1,N_2405,N_2568);
nor UO_2 (O_2,N_2303,N_2586);
and UO_3 (O_3,N_2814,N_2307);
nor UO_4 (O_4,N_2394,N_2609);
nand UO_5 (O_5,N_2426,N_2382);
nor UO_6 (O_6,N_2437,N_2756);
nor UO_7 (O_7,N_2862,N_2272);
and UO_8 (O_8,N_2885,N_2353);
nand UO_9 (O_9,N_2493,N_2963);
or UO_10 (O_10,N_2517,N_2552);
nand UO_11 (O_11,N_2624,N_2514);
nand UO_12 (O_12,N_2314,N_2306);
or UO_13 (O_13,N_2560,N_2444);
nor UO_14 (O_14,N_2789,N_2978);
nor UO_15 (O_15,N_2572,N_2258);
xor UO_16 (O_16,N_2599,N_2810);
nor UO_17 (O_17,N_2754,N_2906);
or UO_18 (O_18,N_2799,N_2470);
nand UO_19 (O_19,N_2429,N_2705);
nor UO_20 (O_20,N_2686,N_2519);
nand UO_21 (O_21,N_2784,N_2373);
nor UO_22 (O_22,N_2701,N_2850);
and UO_23 (O_23,N_2466,N_2261);
nor UO_24 (O_24,N_2853,N_2869);
and UO_25 (O_25,N_2908,N_2494);
and UO_26 (O_26,N_2366,N_2865);
or UO_27 (O_27,N_2372,N_2492);
or UO_28 (O_28,N_2635,N_2331);
or UO_29 (O_29,N_2846,N_2495);
nand UO_30 (O_30,N_2556,N_2914);
nand UO_31 (O_31,N_2293,N_2581);
nand UO_32 (O_32,N_2699,N_2950);
nor UO_33 (O_33,N_2792,N_2652);
nor UO_34 (O_34,N_2297,N_2641);
and UO_35 (O_35,N_2897,N_2743);
nor UO_36 (O_36,N_2421,N_2887);
or UO_37 (O_37,N_2540,N_2286);
nand UO_38 (O_38,N_2974,N_2323);
nor UO_39 (O_39,N_2377,N_2413);
nand UO_40 (O_40,N_2951,N_2453);
nor UO_41 (O_41,N_2940,N_2656);
nor UO_42 (O_42,N_2833,N_2925);
and UO_43 (O_43,N_2773,N_2555);
nor UO_44 (O_44,N_2937,N_2956);
or UO_45 (O_45,N_2481,N_2328);
nand UO_46 (O_46,N_2681,N_2881);
nand UO_47 (O_47,N_2562,N_2325);
or UO_48 (O_48,N_2612,N_2276);
nand UO_49 (O_49,N_2619,N_2473);
and UO_50 (O_50,N_2785,N_2991);
nand UO_51 (O_51,N_2278,N_2574);
and UO_52 (O_52,N_2528,N_2874);
nand UO_53 (O_53,N_2938,N_2883);
nand UO_54 (O_54,N_2875,N_2888);
and UO_55 (O_55,N_2873,N_2456);
nand UO_56 (O_56,N_2904,N_2428);
nor UO_57 (O_57,N_2847,N_2305);
nor UO_58 (O_58,N_2500,N_2797);
or UO_59 (O_59,N_2858,N_2917);
nand UO_60 (O_60,N_2597,N_2700);
nor UO_61 (O_61,N_2588,N_2291);
or UO_62 (O_62,N_2840,N_2545);
nor UO_63 (O_63,N_2804,N_2318);
nor UO_64 (O_64,N_2651,N_2300);
and UO_65 (O_65,N_2465,N_2987);
nor UO_66 (O_66,N_2871,N_2665);
or UO_67 (O_67,N_2482,N_2851);
or UO_68 (O_68,N_2768,N_2455);
or UO_69 (O_69,N_2687,N_2721);
and UO_70 (O_70,N_2460,N_2928);
nor UO_71 (O_71,N_2905,N_2817);
nor UO_72 (O_72,N_2359,N_2504);
nor UO_73 (O_73,N_2923,N_2330);
and UO_74 (O_74,N_2884,N_2393);
nor UO_75 (O_75,N_2296,N_2876);
nand UO_76 (O_76,N_2315,N_2713);
nand UO_77 (O_77,N_2600,N_2707);
nor UO_78 (O_78,N_2692,N_2622);
or UO_79 (O_79,N_2658,N_2302);
nand UO_80 (O_80,N_2724,N_2759);
nor UO_81 (O_81,N_2535,N_2605);
and UO_82 (O_82,N_2774,N_2832);
or UO_83 (O_83,N_2835,N_2412);
nor UO_84 (O_84,N_2990,N_2601);
nor UO_85 (O_85,N_2549,N_2625);
nor UO_86 (O_86,N_2866,N_2653);
nor UO_87 (O_87,N_2538,N_2354);
or UO_88 (O_88,N_2253,N_2631);
and UO_89 (O_89,N_2578,N_2844);
and UO_90 (O_90,N_2396,N_2526);
or UO_91 (O_91,N_2746,N_2387);
nand UO_92 (O_92,N_2423,N_2585);
nand UO_93 (O_93,N_2436,N_2731);
nor UO_94 (O_94,N_2663,N_2335);
nor UO_95 (O_95,N_2899,N_2469);
or UO_96 (O_96,N_2269,N_2410);
nand UO_97 (O_97,N_2918,N_2669);
and UO_98 (O_98,N_2606,N_2638);
nand UO_99 (O_99,N_2979,N_2758);
nand UO_100 (O_100,N_2486,N_2666);
or UO_101 (O_101,N_2803,N_2988);
nand UO_102 (O_102,N_2634,N_2621);
nand UO_103 (O_103,N_2725,N_2348);
xnor UO_104 (O_104,N_2563,N_2801);
or UO_105 (O_105,N_2843,N_2831);
nor UO_106 (O_106,N_2970,N_2676);
nand UO_107 (O_107,N_2854,N_2339);
or UO_108 (O_108,N_2936,N_2818);
nor UO_109 (O_109,N_2714,N_2274);
or UO_110 (O_110,N_2878,N_2298);
nor UO_111 (O_111,N_2525,N_2824);
and UO_112 (O_112,N_2781,N_2934);
nand UO_113 (O_113,N_2659,N_2633);
or UO_114 (O_114,N_2886,N_2271);
nor UO_115 (O_115,N_2367,N_2856);
and UO_116 (O_116,N_2948,N_2288);
nand UO_117 (O_117,N_2523,N_2900);
nand UO_118 (O_118,N_2501,N_2356);
nor UO_119 (O_119,N_2975,N_2484);
nor UO_120 (O_120,N_2769,N_2966);
and UO_121 (O_121,N_2476,N_2439);
nor UO_122 (O_122,N_2573,N_2349);
or UO_123 (O_123,N_2608,N_2332);
nand UO_124 (O_124,N_2971,N_2507);
nand UO_125 (O_125,N_2326,N_2986);
or UO_126 (O_126,N_2941,N_2596);
nand UO_127 (O_127,N_2648,N_2842);
or UO_128 (O_128,N_2409,N_2960);
nor UO_129 (O_129,N_2637,N_2374);
and UO_130 (O_130,N_2702,N_2380);
or UO_131 (O_131,N_2644,N_2610);
or UO_132 (O_132,N_2931,N_2965);
and UO_133 (O_133,N_2613,N_2683);
and UO_134 (O_134,N_2593,N_2390);
nand UO_135 (O_135,N_2491,N_2776);
and UO_136 (O_136,N_2712,N_2358);
or UO_137 (O_137,N_2877,N_2760);
or UO_138 (O_138,N_2317,N_2431);
or UO_139 (O_139,N_2901,N_2259);
nand UO_140 (O_140,N_2250,N_2787);
or UO_141 (O_141,N_2312,N_2376);
nor UO_142 (O_142,N_2567,N_2996);
nor UO_143 (O_143,N_2282,N_2468);
or UO_144 (O_144,N_2639,N_2920);
or UO_145 (O_145,N_2320,N_2660);
nor UO_146 (O_146,N_2794,N_2509);
or UO_147 (O_147,N_2662,N_2350);
and UO_148 (O_148,N_2748,N_2790);
and UO_149 (O_149,N_2984,N_2632);
nor UO_150 (O_150,N_2365,N_2755);
or UO_151 (O_151,N_2694,N_2547);
xnor UO_152 (O_152,N_2689,N_2848);
nor UO_153 (O_153,N_2459,N_2706);
nand UO_154 (O_154,N_2999,N_2506);
nor UO_155 (O_155,N_2434,N_2762);
nor UO_156 (O_156,N_2252,N_2375);
nand UO_157 (O_157,N_2337,N_2441);
nand UO_158 (O_158,N_2451,N_2417);
nor UO_159 (O_159,N_2565,N_2998);
nand UO_160 (O_160,N_2402,N_2723);
nand UO_161 (O_161,N_2825,N_2779);
nor UO_162 (O_162,N_2962,N_2418);
nand UO_163 (O_163,N_2642,N_2811);
nor UO_164 (O_164,N_2682,N_2602);
and UO_165 (O_165,N_2497,N_2362);
and UO_166 (O_166,N_2364,N_2968);
and UO_167 (O_167,N_2577,N_2343);
and UO_168 (O_168,N_2793,N_2630);
or UO_169 (O_169,N_2932,N_2520);
nand UO_170 (O_170,N_2595,N_2916);
nor UO_171 (O_171,N_2802,N_2720);
nor UO_172 (O_172,N_2718,N_2935);
or UO_173 (O_173,N_2989,N_2284);
nor UO_174 (O_174,N_2691,N_2281);
nor UO_175 (O_175,N_2620,N_2379);
nand UO_176 (O_176,N_2628,N_2564);
or UO_177 (O_177,N_2255,N_2598);
nand UO_178 (O_178,N_2921,N_2403);
nor UO_179 (O_179,N_2942,N_2452);
and UO_180 (O_180,N_2747,N_2430);
nor UO_181 (O_181,N_2679,N_2744);
or UO_182 (O_182,N_2959,N_2708);
nor UO_183 (O_183,N_2254,N_2684);
and UO_184 (O_184,N_2667,N_2741);
nor UO_185 (O_185,N_2615,N_2378);
or UO_186 (O_186,N_2344,N_2280);
nand UO_187 (O_187,N_2961,N_2477);
nor UO_188 (O_188,N_2313,N_2438);
and UO_189 (O_189,N_2397,N_2419);
and UO_190 (O_190,N_2454,N_2551);
nand UO_191 (O_191,N_2443,N_2321);
or UO_192 (O_192,N_2503,N_2995);
nand UO_193 (O_193,N_2894,N_2767);
nor UO_194 (O_194,N_2765,N_2386);
or UO_195 (O_195,N_2912,N_2704);
nor UO_196 (O_196,N_2299,N_2442);
or UO_197 (O_197,N_2953,N_2745);
nand UO_198 (O_198,N_2715,N_2532);
nor UO_199 (O_199,N_2902,N_2757);
nor UO_200 (O_200,N_2536,N_2910);
nor UO_201 (O_201,N_2636,N_2827);
nand UO_202 (O_202,N_2327,N_2279);
or UO_203 (O_203,N_2558,N_2262);
and UO_204 (O_204,N_2485,N_2550);
nand UO_205 (O_205,N_2414,N_2777);
and UO_206 (O_206,N_2450,N_2997);
xnor UO_207 (O_207,N_2457,N_2859);
or UO_208 (O_208,N_2929,N_2533);
or UO_209 (O_209,N_2571,N_2993);
and UO_210 (O_210,N_2719,N_2816);
nor UO_211 (O_211,N_2487,N_2717);
nor UO_212 (O_212,N_2710,N_2983);
and UO_213 (O_213,N_2919,N_2675);
xor UO_214 (O_214,N_2289,N_2643);
and UO_215 (O_215,N_2994,N_2815);
nor UO_216 (O_216,N_2408,N_2582);
nor UO_217 (O_217,N_2370,N_2614);
and UO_218 (O_218,N_2892,N_2273);
nand UO_219 (O_219,N_2890,N_2406);
nand UO_220 (O_220,N_2478,N_2664);
nor UO_221 (O_221,N_2333,N_2310);
and UO_222 (O_222,N_2945,N_2969);
nand UO_223 (O_223,N_2727,N_2680);
nand UO_224 (O_224,N_2909,N_2957);
nor UO_225 (O_225,N_2579,N_2295);
nand UO_226 (O_226,N_2864,N_2576);
nand UO_227 (O_227,N_2780,N_2355);
nor UO_228 (O_228,N_2911,N_2496);
and UO_229 (O_229,N_2251,N_2674);
nor UO_230 (O_230,N_2357,N_2806);
and UO_231 (O_231,N_2889,N_2839);
nor UO_232 (O_232,N_2980,N_2823);
nor UO_233 (O_233,N_2294,N_2308);
and UO_234 (O_234,N_2471,N_2479);
and UO_235 (O_235,N_2537,N_2316);
nor UO_236 (O_236,N_2837,N_2527);
nand UO_237 (O_237,N_2617,N_2860);
and UO_238 (O_238,N_2753,N_2750);
or UO_239 (O_239,N_2924,N_2590);
nor UO_240 (O_240,N_2480,N_2285);
or UO_241 (O_241,N_2764,N_2435);
and UO_242 (O_242,N_2913,N_2381);
nor UO_243 (O_243,N_2543,N_2783);
and UO_244 (O_244,N_2260,N_2982);
and UO_245 (O_245,N_2518,N_2268);
and UO_246 (O_246,N_2618,N_2734);
and UO_247 (O_247,N_2770,N_2407);
or UO_248 (O_248,N_2392,N_2872);
or UO_249 (O_249,N_2541,N_2311);
or UO_250 (O_250,N_2627,N_2739);
nand UO_251 (O_251,N_2670,N_2967);
and UO_252 (O_252,N_2368,N_2855);
nand UO_253 (O_253,N_2742,N_2616);
or UO_254 (O_254,N_2510,N_2726);
nor UO_255 (O_255,N_2677,N_2861);
nor UO_256 (O_256,N_2287,N_2645);
and UO_257 (O_257,N_2398,N_2657);
and UO_258 (O_258,N_2829,N_2626);
nand UO_259 (O_259,N_2733,N_2880);
or UO_260 (O_260,N_2594,N_2907);
and UO_261 (O_261,N_2334,N_2788);
or UO_262 (O_262,N_2973,N_2432);
and UO_263 (O_263,N_2265,N_2369);
and UO_264 (O_264,N_2304,N_2384);
or UO_265 (O_265,N_2964,N_2290);
nand UO_266 (O_266,N_2530,N_2542);
or UO_267 (O_267,N_2508,N_2363);
nand UO_268 (O_268,N_2654,N_2342);
nor UO_269 (O_269,N_2834,N_2433);
nor UO_270 (O_270,N_2729,N_2711);
nand UO_271 (O_271,N_2749,N_2474);
and UO_272 (O_272,N_2821,N_2944);
nand UO_273 (O_273,N_2766,N_2352);
or UO_274 (O_274,N_2943,N_2399);
and UO_275 (O_275,N_2926,N_2604);
or UO_276 (O_276,N_2270,N_2778);
nand UO_277 (O_277,N_2895,N_2800);
nor UO_278 (O_278,N_2868,N_2425);
and UO_279 (O_279,N_2752,N_2322);
nor UO_280 (O_280,N_2420,N_2830);
nand UO_281 (O_281,N_2650,N_2611);
nand UO_282 (O_282,N_2688,N_2805);
and UO_283 (O_283,N_2673,N_2548);
or UO_284 (O_284,N_2782,N_2267);
nor UO_285 (O_285,N_2703,N_2857);
or UO_286 (O_286,N_2347,N_2440);
or UO_287 (O_287,N_2820,N_2661);
nand UO_288 (O_288,N_2575,N_2685);
nand UO_289 (O_289,N_2791,N_2695);
and UO_290 (O_290,N_2461,N_2922);
nand UO_291 (O_291,N_2587,N_2388);
or UO_292 (O_292,N_2896,N_2882);
and UO_293 (O_293,N_2512,N_2730);
nand UO_294 (O_294,N_2401,N_2505);
and UO_295 (O_295,N_2709,N_2400);
and UO_296 (O_296,N_2483,N_2716);
and UO_297 (O_297,N_2553,N_2319);
nand UO_298 (O_298,N_2580,N_2891);
nor UO_299 (O_299,N_2589,N_2972);
and UO_300 (O_300,N_2488,N_2849);
nand UO_301 (O_301,N_2371,N_2499);
nand UO_302 (O_302,N_2826,N_2649);
and UO_303 (O_303,N_2389,N_2534);
or UO_304 (O_304,N_2690,N_2722);
nand UO_305 (O_305,N_2728,N_2809);
or UO_306 (O_306,N_2863,N_2698);
and UO_307 (O_307,N_2329,N_2772);
or UO_308 (O_308,N_2592,N_2795);
and UO_309 (O_309,N_2822,N_2529);
and UO_310 (O_310,N_2345,N_2395);
nand UO_311 (O_311,N_2531,N_2458);
or UO_312 (O_312,N_2415,N_2445);
and UO_313 (O_313,N_2257,N_2893);
nand UO_314 (O_314,N_2557,N_2502);
nor UO_315 (O_315,N_2336,N_2775);
and UO_316 (O_316,N_2671,N_2561);
nor UO_317 (O_317,N_2277,N_2603);
or UO_318 (O_318,N_2761,N_2447);
nand UO_319 (O_319,N_2584,N_2448);
or UO_320 (O_320,N_2647,N_2607);
and UO_321 (O_321,N_2696,N_2786);
nor UO_322 (O_322,N_2513,N_2411);
and UO_323 (O_323,N_2836,N_2736);
nand UO_324 (O_324,N_2903,N_2841);
and UO_325 (O_325,N_2958,N_2977);
nor UO_326 (O_326,N_2404,N_2655);
or UO_327 (O_327,N_2292,N_2732);
and UO_328 (O_328,N_2475,N_2522);
nor UO_329 (O_329,N_2751,N_2283);
nor UO_330 (O_330,N_2340,N_2898);
or UO_331 (O_331,N_2763,N_2351);
and UO_332 (O_332,N_2424,N_2985);
or UO_333 (O_333,N_2828,N_2385);
or UO_334 (O_334,N_2264,N_2955);
xor UO_335 (O_335,N_2427,N_2852);
nand UO_336 (O_336,N_2697,N_2338);
nor UO_337 (O_337,N_2933,N_2813);
or UO_338 (O_338,N_2490,N_2623);
nand UO_339 (O_339,N_2256,N_2693);
or UO_340 (O_340,N_2583,N_2266);
nor UO_341 (O_341,N_2566,N_2383);
nor UO_342 (O_342,N_2838,N_2646);
nor UO_343 (O_343,N_2489,N_2498);
and UO_344 (O_344,N_2879,N_2808);
nor UO_345 (O_345,N_2446,N_2546);
nor UO_346 (O_346,N_2467,N_2361);
and UO_347 (O_347,N_2915,N_2629);
or UO_348 (O_348,N_2867,N_2992);
nand UO_349 (O_349,N_2570,N_2949);
or UO_350 (O_350,N_2870,N_2927);
and UO_351 (O_351,N_2740,N_2516);
nand UO_352 (O_352,N_2341,N_2524);
nand UO_353 (O_353,N_2569,N_2952);
nand UO_354 (O_354,N_2554,N_2263);
or UO_355 (O_355,N_2798,N_2735);
nor UO_356 (O_356,N_2309,N_2930);
nand UO_357 (O_357,N_2464,N_2812);
xnor UO_358 (O_358,N_2449,N_2796);
nor UO_359 (O_359,N_2515,N_2737);
or UO_360 (O_360,N_2391,N_2640);
nand UO_361 (O_361,N_2939,N_2511);
and UO_362 (O_362,N_2807,N_2416);
or UO_363 (O_363,N_2678,N_2463);
and UO_364 (O_364,N_2301,N_2462);
and UO_365 (O_365,N_2521,N_2324);
and UO_366 (O_366,N_2981,N_2360);
xnor UO_367 (O_367,N_2947,N_2672);
or UO_368 (O_368,N_2544,N_2559);
and UO_369 (O_369,N_2346,N_2954);
and UO_370 (O_370,N_2976,N_2422);
nor UO_371 (O_371,N_2539,N_2946);
or UO_372 (O_372,N_2738,N_2275);
or UO_373 (O_373,N_2591,N_2472);
and UO_374 (O_374,N_2845,N_2819);
nand UO_375 (O_375,N_2664,N_2763);
or UO_376 (O_376,N_2346,N_2631);
nand UO_377 (O_377,N_2727,N_2861);
nor UO_378 (O_378,N_2726,N_2669);
or UO_379 (O_379,N_2401,N_2534);
or UO_380 (O_380,N_2662,N_2978);
nor UO_381 (O_381,N_2664,N_2830);
or UO_382 (O_382,N_2973,N_2319);
and UO_383 (O_383,N_2901,N_2848);
xnor UO_384 (O_384,N_2789,N_2812);
and UO_385 (O_385,N_2578,N_2355);
and UO_386 (O_386,N_2878,N_2260);
and UO_387 (O_387,N_2497,N_2492);
nor UO_388 (O_388,N_2880,N_2813);
and UO_389 (O_389,N_2499,N_2297);
or UO_390 (O_390,N_2824,N_2398);
nand UO_391 (O_391,N_2925,N_2745);
or UO_392 (O_392,N_2741,N_2797);
or UO_393 (O_393,N_2956,N_2256);
and UO_394 (O_394,N_2550,N_2335);
nor UO_395 (O_395,N_2498,N_2346);
nor UO_396 (O_396,N_2827,N_2520);
nand UO_397 (O_397,N_2389,N_2575);
and UO_398 (O_398,N_2681,N_2532);
nand UO_399 (O_399,N_2713,N_2535);
or UO_400 (O_400,N_2464,N_2404);
nand UO_401 (O_401,N_2342,N_2450);
nand UO_402 (O_402,N_2993,N_2391);
or UO_403 (O_403,N_2310,N_2965);
and UO_404 (O_404,N_2677,N_2631);
nand UO_405 (O_405,N_2669,N_2349);
nand UO_406 (O_406,N_2874,N_2667);
nand UO_407 (O_407,N_2283,N_2397);
nor UO_408 (O_408,N_2598,N_2330);
nor UO_409 (O_409,N_2661,N_2912);
and UO_410 (O_410,N_2549,N_2386);
nor UO_411 (O_411,N_2362,N_2591);
or UO_412 (O_412,N_2860,N_2283);
nor UO_413 (O_413,N_2544,N_2665);
nor UO_414 (O_414,N_2435,N_2880);
or UO_415 (O_415,N_2545,N_2526);
or UO_416 (O_416,N_2713,N_2783);
nor UO_417 (O_417,N_2632,N_2377);
or UO_418 (O_418,N_2606,N_2747);
or UO_419 (O_419,N_2729,N_2888);
and UO_420 (O_420,N_2607,N_2564);
or UO_421 (O_421,N_2656,N_2382);
or UO_422 (O_422,N_2356,N_2665);
nand UO_423 (O_423,N_2949,N_2284);
or UO_424 (O_424,N_2931,N_2846);
nor UO_425 (O_425,N_2576,N_2543);
or UO_426 (O_426,N_2458,N_2313);
nor UO_427 (O_427,N_2650,N_2797);
nand UO_428 (O_428,N_2768,N_2425);
or UO_429 (O_429,N_2387,N_2964);
nor UO_430 (O_430,N_2934,N_2253);
or UO_431 (O_431,N_2778,N_2929);
xnor UO_432 (O_432,N_2671,N_2482);
nor UO_433 (O_433,N_2364,N_2396);
or UO_434 (O_434,N_2868,N_2565);
nand UO_435 (O_435,N_2382,N_2581);
nand UO_436 (O_436,N_2313,N_2790);
and UO_437 (O_437,N_2798,N_2877);
and UO_438 (O_438,N_2463,N_2628);
nor UO_439 (O_439,N_2972,N_2367);
nand UO_440 (O_440,N_2436,N_2730);
or UO_441 (O_441,N_2703,N_2731);
or UO_442 (O_442,N_2436,N_2658);
and UO_443 (O_443,N_2347,N_2744);
and UO_444 (O_444,N_2536,N_2749);
or UO_445 (O_445,N_2652,N_2257);
nand UO_446 (O_446,N_2457,N_2336);
or UO_447 (O_447,N_2427,N_2501);
and UO_448 (O_448,N_2339,N_2660);
and UO_449 (O_449,N_2802,N_2651);
nand UO_450 (O_450,N_2548,N_2508);
and UO_451 (O_451,N_2983,N_2664);
and UO_452 (O_452,N_2273,N_2496);
or UO_453 (O_453,N_2569,N_2324);
nand UO_454 (O_454,N_2304,N_2464);
nand UO_455 (O_455,N_2551,N_2388);
and UO_456 (O_456,N_2266,N_2513);
xor UO_457 (O_457,N_2624,N_2251);
or UO_458 (O_458,N_2488,N_2582);
nor UO_459 (O_459,N_2750,N_2777);
nor UO_460 (O_460,N_2772,N_2581);
and UO_461 (O_461,N_2259,N_2620);
or UO_462 (O_462,N_2775,N_2511);
and UO_463 (O_463,N_2505,N_2717);
nor UO_464 (O_464,N_2848,N_2874);
nor UO_465 (O_465,N_2852,N_2842);
or UO_466 (O_466,N_2333,N_2705);
nand UO_467 (O_467,N_2673,N_2555);
and UO_468 (O_468,N_2283,N_2774);
nand UO_469 (O_469,N_2346,N_2381);
nand UO_470 (O_470,N_2419,N_2996);
nor UO_471 (O_471,N_2703,N_2333);
nor UO_472 (O_472,N_2968,N_2717);
and UO_473 (O_473,N_2286,N_2952);
or UO_474 (O_474,N_2748,N_2609);
or UO_475 (O_475,N_2987,N_2738);
nor UO_476 (O_476,N_2781,N_2269);
and UO_477 (O_477,N_2853,N_2872);
or UO_478 (O_478,N_2327,N_2566);
nand UO_479 (O_479,N_2648,N_2448);
nor UO_480 (O_480,N_2809,N_2262);
nand UO_481 (O_481,N_2833,N_2252);
or UO_482 (O_482,N_2703,N_2752);
and UO_483 (O_483,N_2739,N_2456);
nand UO_484 (O_484,N_2759,N_2508);
or UO_485 (O_485,N_2807,N_2310);
nand UO_486 (O_486,N_2908,N_2623);
xor UO_487 (O_487,N_2294,N_2883);
or UO_488 (O_488,N_2793,N_2551);
nor UO_489 (O_489,N_2795,N_2562);
nand UO_490 (O_490,N_2443,N_2656);
nand UO_491 (O_491,N_2557,N_2548);
or UO_492 (O_492,N_2518,N_2755);
nor UO_493 (O_493,N_2576,N_2446);
nor UO_494 (O_494,N_2995,N_2824);
nor UO_495 (O_495,N_2379,N_2376);
nor UO_496 (O_496,N_2942,N_2955);
xnor UO_497 (O_497,N_2325,N_2263);
or UO_498 (O_498,N_2985,N_2854);
and UO_499 (O_499,N_2446,N_2772);
endmodule