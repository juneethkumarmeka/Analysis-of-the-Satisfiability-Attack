module basic_750_5000_1000_5_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_15,In_118);
nor U1 (N_1,In_164,In_219);
nand U2 (N_2,In_6,In_155);
nor U3 (N_3,In_480,In_721);
or U4 (N_4,In_166,In_553);
and U5 (N_5,In_59,In_695);
and U6 (N_6,In_134,In_530);
and U7 (N_7,In_541,In_549);
and U8 (N_8,In_489,In_653);
and U9 (N_9,In_637,In_552);
or U10 (N_10,In_399,In_42);
and U11 (N_11,In_660,In_383);
nand U12 (N_12,In_335,In_570);
and U13 (N_13,In_439,In_318);
or U14 (N_14,In_72,In_131);
and U15 (N_15,In_438,In_370);
nand U16 (N_16,In_427,In_581);
nand U17 (N_17,In_182,In_706);
and U18 (N_18,In_665,In_705);
or U19 (N_19,In_57,In_266);
and U20 (N_20,In_731,In_436);
xnor U21 (N_21,In_623,In_395);
or U22 (N_22,In_109,In_607);
nand U23 (N_23,In_286,In_49);
nor U24 (N_24,In_401,In_160);
nand U25 (N_25,In_75,In_478);
nor U26 (N_26,In_260,In_17);
nand U27 (N_27,In_594,In_415);
and U28 (N_28,In_545,In_672);
or U29 (N_29,In_363,In_408);
and U30 (N_30,In_741,In_384);
nand U31 (N_31,In_38,In_218);
nand U32 (N_32,In_104,In_224);
or U33 (N_33,In_678,In_176);
or U34 (N_34,In_681,In_40);
or U35 (N_35,In_112,In_19);
or U36 (N_36,In_454,In_471);
or U37 (N_37,In_126,In_125);
nor U38 (N_38,In_61,In_511);
nor U39 (N_39,In_371,In_196);
nor U40 (N_40,In_127,In_12);
or U41 (N_41,In_357,In_734);
or U42 (N_42,In_240,In_246);
nor U43 (N_43,In_597,In_696);
and U44 (N_44,In_114,In_729);
and U45 (N_45,In_404,In_199);
nor U46 (N_46,In_239,In_270);
and U47 (N_47,In_373,In_668);
nand U48 (N_48,In_650,In_120);
or U49 (N_49,In_567,In_647);
and U50 (N_50,In_157,In_303);
or U51 (N_51,In_66,In_736);
nor U52 (N_52,In_187,In_361);
nor U53 (N_53,In_58,In_600);
and U54 (N_54,In_711,In_391);
or U55 (N_55,In_381,In_732);
and U56 (N_56,In_22,In_161);
nand U57 (N_57,In_100,In_130);
nand U58 (N_58,In_586,In_669);
and U59 (N_59,In_618,In_228);
and U60 (N_60,In_205,In_296);
and U61 (N_61,In_188,In_382);
nand U62 (N_62,In_119,In_251);
or U63 (N_63,In_298,In_25);
nand U64 (N_64,In_128,In_414);
or U65 (N_65,In_186,In_516);
or U66 (N_66,In_314,In_233);
or U67 (N_67,In_204,In_247);
nor U68 (N_68,In_483,In_649);
nor U69 (N_69,In_368,In_9);
nor U70 (N_70,In_619,In_47);
and U71 (N_71,In_577,In_501);
or U72 (N_72,In_611,In_238);
and U73 (N_73,In_662,In_437);
or U74 (N_74,In_10,In_542);
and U75 (N_75,In_200,In_379);
or U76 (N_76,In_201,In_525);
or U77 (N_77,In_275,In_617);
and U78 (N_78,In_496,In_304);
or U79 (N_79,In_277,In_95);
and U80 (N_80,In_630,In_282);
or U81 (N_81,In_26,In_31);
or U82 (N_82,In_728,In_641);
nor U83 (N_83,In_343,In_624);
or U84 (N_84,In_227,In_253);
nor U85 (N_85,In_74,In_595);
nand U86 (N_86,In_244,In_132);
and U87 (N_87,In_505,In_432);
nand U88 (N_88,In_94,In_550);
nor U89 (N_89,In_488,In_431);
and U90 (N_90,In_389,In_689);
nor U91 (N_91,In_338,In_529);
or U92 (N_92,In_537,In_472);
and U93 (N_93,In_674,In_329);
nand U94 (N_94,In_297,In_78);
nand U95 (N_95,In_36,In_710);
and U96 (N_96,In_321,In_216);
nor U97 (N_97,In_378,In_601);
nor U98 (N_98,In_326,In_101);
nand U99 (N_99,In_687,In_453);
or U100 (N_100,In_485,In_707);
nor U101 (N_101,In_733,In_392);
and U102 (N_102,In_573,In_7);
and U103 (N_103,In_463,In_613);
or U104 (N_104,In_446,In_517);
nor U105 (N_105,In_367,In_85);
and U106 (N_106,In_425,In_614);
or U107 (N_107,In_195,In_281);
or U108 (N_108,In_102,In_83);
nand U109 (N_109,In_461,In_450);
and U110 (N_110,In_465,In_261);
nor U111 (N_111,In_434,In_346);
xnor U112 (N_112,In_521,In_352);
or U113 (N_113,In_725,In_234);
nand U114 (N_114,In_143,In_492);
nor U115 (N_115,In_150,In_295);
nor U116 (N_116,In_257,In_158);
nand U117 (N_117,In_460,In_443);
nand U118 (N_118,In_355,In_359);
nor U119 (N_119,In_703,In_46);
nand U120 (N_120,In_691,In_615);
and U121 (N_121,In_274,In_646);
or U122 (N_122,In_299,In_591);
and U123 (N_123,In_675,In_123);
nor U124 (N_124,In_583,In_593);
or U125 (N_125,In_533,In_612);
and U126 (N_126,In_51,In_466);
nor U127 (N_127,In_688,In_590);
xor U128 (N_128,In_458,In_555);
and U129 (N_129,In_148,In_663);
nor U130 (N_130,In_291,In_154);
nand U131 (N_131,In_642,In_579);
and U132 (N_132,In_474,In_279);
nor U133 (N_133,In_121,In_53);
nand U134 (N_134,In_177,In_440);
nor U135 (N_135,In_560,In_667);
nand U136 (N_136,In_745,In_726);
nand U137 (N_137,In_347,In_727);
nand U138 (N_138,In_174,In_226);
or U139 (N_139,In_410,In_147);
nor U140 (N_140,In_167,In_657);
and U141 (N_141,In_222,In_34);
nor U142 (N_142,In_494,In_290);
or U143 (N_143,In_500,In_551);
nand U144 (N_144,In_353,In_620);
or U145 (N_145,In_292,In_634);
nand U146 (N_146,In_628,In_207);
nor U147 (N_147,In_548,In_142);
or U148 (N_148,In_162,In_68);
nand U149 (N_149,In_151,In_563);
and U150 (N_150,In_429,In_445);
or U151 (N_151,In_189,In_518);
nand U152 (N_152,In_423,In_71);
nand U153 (N_153,In_522,In_481);
nand U154 (N_154,In_639,In_97);
nor U155 (N_155,In_743,In_340);
xor U156 (N_156,In_385,In_449);
nand U157 (N_157,In_258,In_564);
and U158 (N_158,In_310,In_106);
nor U159 (N_159,In_682,In_193);
or U160 (N_160,In_271,In_333);
nor U161 (N_161,In_676,In_141);
nor U162 (N_162,In_576,In_293);
nor U163 (N_163,In_625,In_67);
nand U164 (N_164,In_362,In_602);
and U165 (N_165,In_209,In_418);
nor U166 (N_166,In_635,In_116);
nand U167 (N_167,In_287,In_405);
xnor U168 (N_168,In_2,In_64);
and U169 (N_169,In_21,In_210);
nor U170 (N_170,In_580,In_543);
nand U171 (N_171,In_35,In_722);
or U172 (N_172,In_319,In_532);
nor U173 (N_173,In_73,In_428);
nand U174 (N_174,In_37,In_629);
or U175 (N_175,In_221,In_502);
or U176 (N_176,In_81,In_197);
nand U177 (N_177,In_477,In_360);
and U178 (N_178,In_544,In_685);
and U179 (N_179,In_90,In_351);
nand U180 (N_180,In_719,In_495);
nand U181 (N_181,In_23,In_237);
nor U182 (N_182,In_337,In_411);
or U183 (N_183,In_235,In_365);
nand U184 (N_184,In_376,In_616);
nand U185 (N_185,In_582,In_331);
nor U186 (N_186,In_179,In_265);
nor U187 (N_187,In_124,In_185);
and U188 (N_188,In_394,In_11);
nand U189 (N_189,In_349,In_413);
or U190 (N_190,In_144,In_621);
nor U191 (N_191,In_43,In_467);
nand U192 (N_192,In_571,In_504);
and U193 (N_193,In_14,In_172);
nand U194 (N_194,In_269,In_278);
or U195 (N_195,In_165,In_178);
nand U196 (N_196,In_89,In_402);
nor U197 (N_197,In_744,In_609);
or U198 (N_198,In_574,In_441);
nand U199 (N_199,In_203,In_473);
nand U200 (N_200,In_198,In_538);
nor U201 (N_201,In_739,In_54);
nand U202 (N_202,In_354,In_153);
and U203 (N_203,In_698,In_747);
nand U204 (N_204,In_273,In_330);
nand U205 (N_205,In_372,In_208);
and U206 (N_206,In_444,In_152);
and U207 (N_207,In_554,In_626);
or U208 (N_208,In_515,In_490);
or U209 (N_209,In_704,In_190);
or U210 (N_210,In_417,In_430);
and U211 (N_211,In_531,In_254);
and U212 (N_212,In_631,In_249);
nand U213 (N_213,In_173,In_60);
and U214 (N_214,In_566,In_724);
xor U215 (N_215,In_644,In_746);
nand U216 (N_216,In_175,In_1);
nor U217 (N_217,In_223,In_4);
nor U218 (N_218,In_715,In_252);
nor U219 (N_219,In_403,In_217);
or U220 (N_220,In_632,In_28);
or U221 (N_221,In_108,In_699);
and U222 (N_222,In_526,In_700);
and U223 (N_223,In_32,In_105);
nor U224 (N_224,In_103,In_345);
nor U225 (N_225,In_540,In_679);
nand U226 (N_226,In_146,In_211);
nand U227 (N_227,In_284,In_457);
or U228 (N_228,In_328,In_697);
xor U229 (N_229,In_55,In_643);
and U230 (N_230,In_486,In_497);
nor U231 (N_231,In_742,In_470);
and U232 (N_232,In_191,In_264);
and U233 (N_233,In_670,In_740);
nand U234 (N_234,In_92,In_712);
nand U235 (N_235,In_137,In_556);
nor U236 (N_236,In_588,In_433);
nand U237 (N_237,In_462,In_451);
or U238 (N_238,In_348,In_212);
or U239 (N_239,In_256,In_325);
nand U240 (N_240,In_48,In_70);
and U241 (N_241,In_435,In_133);
or U242 (N_242,In_311,In_547);
or U243 (N_243,In_163,In_350);
nand U244 (N_244,In_263,In_476);
or U245 (N_245,In_168,In_589);
or U246 (N_246,In_342,In_499);
nand U247 (N_247,In_568,In_230);
or U248 (N_248,In_398,In_673);
nand U249 (N_249,In_416,In_693);
nor U250 (N_250,In_135,In_664);
nor U251 (N_251,In_181,In_327);
and U252 (N_252,In_107,In_259);
nand U253 (N_253,In_307,In_484);
nand U254 (N_254,In_80,In_692);
or U255 (N_255,In_468,In_701);
nor U256 (N_256,In_183,In_113);
and U257 (N_257,In_312,In_690);
nor U258 (N_258,In_339,In_420);
nand U259 (N_259,In_336,In_622);
and U260 (N_260,In_585,In_86);
nor U261 (N_261,In_27,In_317);
or U262 (N_262,In_656,In_575);
or U263 (N_263,In_122,In_598);
nand U264 (N_264,In_214,In_714);
or U265 (N_265,In_396,In_375);
nor U266 (N_266,In_510,In_145);
and U267 (N_267,In_289,In_422);
nand U268 (N_268,In_76,In_559);
and U269 (N_269,In_636,In_33);
nor U270 (N_270,In_301,In_400);
nand U271 (N_271,In_694,In_442);
nand U272 (N_272,In_652,In_18);
nand U273 (N_273,In_140,In_651);
or U274 (N_274,In_3,In_412);
nand U275 (N_275,In_369,In_677);
nor U276 (N_276,In_39,In_661);
nand U277 (N_277,In_308,In_65);
and U278 (N_278,In_98,In_730);
nand U279 (N_279,In_606,In_503);
or U280 (N_280,In_52,In_524);
nand U281 (N_281,In_332,In_184);
and U282 (N_282,In_749,In_487);
nor U283 (N_283,In_684,In_215);
and U284 (N_284,In_393,In_519);
nor U285 (N_285,In_305,In_464);
or U286 (N_286,In_170,In_84);
xor U287 (N_287,In_565,In_720);
nand U288 (N_288,In_507,In_283);
and U289 (N_289,In_654,In_316);
and U290 (N_290,In_262,In_324);
nor U291 (N_291,In_236,In_180);
nand U292 (N_292,In_229,In_272);
nor U293 (N_293,In_91,In_280);
or U294 (N_294,In_666,In_426);
nand U295 (N_295,In_479,In_421);
or U296 (N_296,In_309,In_633);
and U297 (N_297,In_220,In_285);
nor U298 (N_298,In_323,In_225);
and U299 (N_299,In_605,In_294);
nand U300 (N_300,In_0,In_386);
and U301 (N_301,In_527,In_380);
or U302 (N_302,In_96,In_202);
nand U303 (N_303,In_717,In_129);
or U304 (N_304,In_138,In_206);
and U305 (N_305,In_93,In_723);
nand U306 (N_306,In_718,In_232);
nor U307 (N_307,In_514,In_534);
and U308 (N_308,In_456,In_77);
or U309 (N_309,In_627,In_546);
nor U310 (N_310,In_506,In_115);
or U311 (N_311,In_409,In_62);
and U312 (N_312,In_455,In_557);
nor U313 (N_313,In_493,In_508);
or U314 (N_314,In_610,In_388);
nand U315 (N_315,In_110,In_50);
nand U316 (N_316,In_709,In_599);
nor U317 (N_317,In_248,In_671);
and U318 (N_318,In_406,In_587);
nand U319 (N_319,In_315,In_255);
nor U320 (N_320,In_366,In_159);
and U321 (N_321,In_659,In_447);
nand U322 (N_322,In_169,In_16);
and U323 (N_323,In_267,In_302);
nand U324 (N_324,In_592,In_686);
nand U325 (N_325,In_117,In_63);
and U326 (N_326,In_300,In_523);
nor U327 (N_327,In_419,In_658);
nand U328 (N_328,In_341,In_748);
nor U329 (N_329,In_29,In_578);
or U330 (N_330,In_475,In_82);
or U331 (N_331,In_374,In_241);
or U332 (N_332,In_528,In_390);
nand U333 (N_333,In_24,In_99);
and U334 (N_334,In_604,In_572);
nand U335 (N_335,In_156,In_88);
and U336 (N_336,In_469,In_306);
or U337 (N_337,In_87,In_680);
nand U338 (N_338,In_708,In_231);
or U339 (N_339,In_171,In_387);
nor U340 (N_340,In_520,In_448);
nand U341 (N_341,In_79,In_30);
nand U342 (N_342,In_640,In_111);
nand U343 (N_343,In_737,In_13);
nor U344 (N_344,In_320,In_364);
and U345 (N_345,In_44,In_648);
nand U346 (N_346,In_558,In_322);
or U347 (N_347,In_713,In_344);
nand U348 (N_348,In_192,In_243);
and U349 (N_349,In_288,In_513);
nor U350 (N_350,In_569,In_397);
or U351 (N_351,In_452,In_149);
and U352 (N_352,In_738,In_407);
nor U353 (N_353,In_655,In_535);
and U354 (N_354,In_213,In_356);
nor U355 (N_355,In_334,In_735);
nand U356 (N_356,In_509,In_377);
nand U357 (N_357,In_45,In_245);
nor U358 (N_358,In_512,In_5);
nor U359 (N_359,In_358,In_608);
and U360 (N_360,In_584,In_41);
nand U361 (N_361,In_603,In_562);
nand U362 (N_362,In_498,In_491);
or U363 (N_363,In_139,In_20);
nor U364 (N_364,In_638,In_683);
and U365 (N_365,In_702,In_313);
or U366 (N_366,In_56,In_561);
nor U367 (N_367,In_69,In_276);
and U368 (N_368,In_645,In_536);
nor U369 (N_369,In_250,In_268);
nor U370 (N_370,In_242,In_482);
nor U371 (N_371,In_194,In_596);
nand U372 (N_372,In_136,In_424);
nand U373 (N_373,In_539,In_716);
nor U374 (N_374,In_459,In_8);
nand U375 (N_375,In_113,In_39);
and U376 (N_376,In_585,In_168);
nand U377 (N_377,In_700,In_737);
nand U378 (N_378,In_653,In_612);
nor U379 (N_379,In_324,In_99);
nor U380 (N_380,In_279,In_29);
or U381 (N_381,In_406,In_523);
and U382 (N_382,In_472,In_263);
nand U383 (N_383,In_251,In_320);
nand U384 (N_384,In_699,In_711);
nand U385 (N_385,In_616,In_38);
nor U386 (N_386,In_395,In_487);
and U387 (N_387,In_479,In_557);
nor U388 (N_388,In_748,In_589);
nor U389 (N_389,In_452,In_449);
nor U390 (N_390,In_667,In_18);
and U391 (N_391,In_110,In_447);
nand U392 (N_392,In_628,In_327);
nor U393 (N_393,In_345,In_478);
nand U394 (N_394,In_601,In_347);
or U395 (N_395,In_445,In_598);
nor U396 (N_396,In_312,In_391);
nand U397 (N_397,In_660,In_39);
or U398 (N_398,In_476,In_150);
or U399 (N_399,In_530,In_684);
nand U400 (N_400,In_182,In_71);
or U401 (N_401,In_168,In_139);
nor U402 (N_402,In_346,In_56);
nor U403 (N_403,In_117,In_362);
and U404 (N_404,In_637,In_697);
nand U405 (N_405,In_717,In_320);
nand U406 (N_406,In_140,In_669);
or U407 (N_407,In_324,In_383);
nor U408 (N_408,In_459,In_132);
and U409 (N_409,In_206,In_584);
and U410 (N_410,In_416,In_400);
or U411 (N_411,In_167,In_405);
nand U412 (N_412,In_211,In_638);
nand U413 (N_413,In_582,In_516);
nand U414 (N_414,In_303,In_530);
nor U415 (N_415,In_185,In_396);
and U416 (N_416,In_60,In_148);
and U417 (N_417,In_29,In_487);
nor U418 (N_418,In_668,In_602);
and U419 (N_419,In_509,In_85);
and U420 (N_420,In_84,In_21);
nand U421 (N_421,In_407,In_514);
or U422 (N_422,In_742,In_198);
nand U423 (N_423,In_243,In_186);
and U424 (N_424,In_241,In_252);
and U425 (N_425,In_567,In_45);
or U426 (N_426,In_634,In_548);
and U427 (N_427,In_112,In_346);
nand U428 (N_428,In_541,In_1);
nor U429 (N_429,In_205,In_347);
nand U430 (N_430,In_659,In_150);
or U431 (N_431,In_345,In_328);
and U432 (N_432,In_2,In_265);
nor U433 (N_433,In_137,In_724);
nor U434 (N_434,In_710,In_102);
and U435 (N_435,In_746,In_563);
nor U436 (N_436,In_52,In_322);
nand U437 (N_437,In_729,In_317);
or U438 (N_438,In_346,In_113);
nor U439 (N_439,In_473,In_716);
and U440 (N_440,In_44,In_292);
nor U441 (N_441,In_537,In_556);
nand U442 (N_442,In_322,In_1);
nand U443 (N_443,In_327,In_621);
nand U444 (N_444,In_280,In_634);
or U445 (N_445,In_703,In_696);
or U446 (N_446,In_696,In_399);
and U447 (N_447,In_276,In_697);
nor U448 (N_448,In_337,In_435);
or U449 (N_449,In_179,In_32);
nor U450 (N_450,In_460,In_414);
nor U451 (N_451,In_256,In_354);
nand U452 (N_452,In_458,In_338);
or U453 (N_453,In_713,In_237);
nor U454 (N_454,In_179,In_35);
nand U455 (N_455,In_58,In_387);
xor U456 (N_456,In_454,In_504);
nor U457 (N_457,In_135,In_590);
nor U458 (N_458,In_710,In_212);
nor U459 (N_459,In_506,In_26);
and U460 (N_460,In_257,In_289);
nor U461 (N_461,In_492,In_296);
and U462 (N_462,In_390,In_251);
or U463 (N_463,In_616,In_550);
nand U464 (N_464,In_243,In_674);
or U465 (N_465,In_479,In_122);
nor U466 (N_466,In_348,In_682);
and U467 (N_467,In_620,In_278);
nand U468 (N_468,In_89,In_227);
and U469 (N_469,In_500,In_166);
nor U470 (N_470,In_71,In_235);
nand U471 (N_471,In_280,In_35);
and U472 (N_472,In_366,In_260);
and U473 (N_473,In_469,In_474);
nand U474 (N_474,In_82,In_345);
and U475 (N_475,In_387,In_532);
and U476 (N_476,In_189,In_433);
and U477 (N_477,In_120,In_334);
and U478 (N_478,In_25,In_377);
nand U479 (N_479,In_216,In_499);
or U480 (N_480,In_380,In_667);
nand U481 (N_481,In_73,In_384);
nand U482 (N_482,In_594,In_252);
and U483 (N_483,In_674,In_700);
nor U484 (N_484,In_237,In_602);
nor U485 (N_485,In_115,In_517);
nand U486 (N_486,In_730,In_60);
and U487 (N_487,In_13,In_486);
and U488 (N_488,In_608,In_159);
nor U489 (N_489,In_651,In_76);
and U490 (N_490,In_271,In_63);
nand U491 (N_491,In_710,In_585);
or U492 (N_492,In_111,In_738);
and U493 (N_493,In_686,In_671);
nor U494 (N_494,In_584,In_453);
nor U495 (N_495,In_595,In_176);
and U496 (N_496,In_532,In_481);
or U497 (N_497,In_543,In_682);
or U498 (N_498,In_399,In_637);
or U499 (N_499,In_655,In_7);
or U500 (N_500,In_158,In_146);
and U501 (N_501,In_288,In_591);
and U502 (N_502,In_402,In_228);
nand U503 (N_503,In_655,In_741);
nand U504 (N_504,In_376,In_59);
nor U505 (N_505,In_251,In_23);
and U506 (N_506,In_95,In_243);
or U507 (N_507,In_735,In_728);
nand U508 (N_508,In_370,In_220);
nor U509 (N_509,In_299,In_142);
nor U510 (N_510,In_479,In_260);
nand U511 (N_511,In_441,In_533);
and U512 (N_512,In_61,In_651);
nand U513 (N_513,In_501,In_54);
nand U514 (N_514,In_214,In_549);
nor U515 (N_515,In_362,In_431);
or U516 (N_516,In_84,In_575);
nand U517 (N_517,In_60,In_635);
nand U518 (N_518,In_84,In_608);
and U519 (N_519,In_580,In_272);
nand U520 (N_520,In_130,In_327);
nor U521 (N_521,In_345,In_367);
nand U522 (N_522,In_576,In_534);
and U523 (N_523,In_551,In_0);
nor U524 (N_524,In_153,In_712);
or U525 (N_525,In_208,In_31);
and U526 (N_526,In_715,In_241);
or U527 (N_527,In_510,In_308);
or U528 (N_528,In_356,In_604);
nor U529 (N_529,In_657,In_638);
nor U530 (N_530,In_287,In_305);
nand U531 (N_531,In_180,In_111);
or U532 (N_532,In_518,In_181);
nor U533 (N_533,In_293,In_301);
nand U534 (N_534,In_490,In_367);
nand U535 (N_535,In_527,In_72);
or U536 (N_536,In_672,In_153);
or U537 (N_537,In_107,In_140);
nand U538 (N_538,In_723,In_150);
nor U539 (N_539,In_407,In_646);
and U540 (N_540,In_151,In_308);
and U541 (N_541,In_729,In_542);
nand U542 (N_542,In_265,In_500);
or U543 (N_543,In_668,In_402);
nand U544 (N_544,In_6,In_215);
and U545 (N_545,In_343,In_231);
nand U546 (N_546,In_201,In_80);
and U547 (N_547,In_455,In_241);
nand U548 (N_548,In_354,In_599);
nor U549 (N_549,In_656,In_480);
nor U550 (N_550,In_749,In_72);
nand U551 (N_551,In_701,In_722);
and U552 (N_552,In_174,In_319);
nor U553 (N_553,In_506,In_148);
nand U554 (N_554,In_331,In_294);
nand U555 (N_555,In_76,In_463);
or U556 (N_556,In_593,In_349);
nand U557 (N_557,In_517,In_158);
and U558 (N_558,In_215,In_694);
nand U559 (N_559,In_502,In_372);
and U560 (N_560,In_594,In_37);
or U561 (N_561,In_233,In_136);
nand U562 (N_562,In_183,In_203);
nor U563 (N_563,In_70,In_735);
and U564 (N_564,In_337,In_485);
or U565 (N_565,In_596,In_351);
nor U566 (N_566,In_677,In_331);
and U567 (N_567,In_146,In_350);
or U568 (N_568,In_559,In_118);
nor U569 (N_569,In_429,In_277);
nand U570 (N_570,In_470,In_28);
and U571 (N_571,In_614,In_137);
nand U572 (N_572,In_446,In_500);
or U573 (N_573,In_450,In_327);
or U574 (N_574,In_10,In_737);
nor U575 (N_575,In_568,In_712);
nand U576 (N_576,In_21,In_606);
or U577 (N_577,In_673,In_119);
and U578 (N_578,In_360,In_625);
nand U579 (N_579,In_519,In_120);
nand U580 (N_580,In_353,In_686);
nand U581 (N_581,In_152,In_263);
or U582 (N_582,In_58,In_339);
nor U583 (N_583,In_556,In_590);
nand U584 (N_584,In_434,In_749);
nor U585 (N_585,In_356,In_18);
nand U586 (N_586,In_147,In_743);
nor U587 (N_587,In_647,In_671);
or U588 (N_588,In_117,In_409);
or U589 (N_589,In_344,In_635);
or U590 (N_590,In_58,In_118);
nand U591 (N_591,In_657,In_533);
nor U592 (N_592,In_563,In_149);
nand U593 (N_593,In_458,In_577);
or U594 (N_594,In_636,In_132);
or U595 (N_595,In_22,In_472);
and U596 (N_596,In_658,In_21);
and U597 (N_597,In_392,In_168);
nand U598 (N_598,In_471,In_97);
xnor U599 (N_599,In_458,In_143);
or U600 (N_600,In_248,In_92);
nand U601 (N_601,In_231,In_475);
or U602 (N_602,In_198,In_506);
nor U603 (N_603,In_430,In_656);
nand U604 (N_604,In_661,In_234);
and U605 (N_605,In_547,In_611);
and U606 (N_606,In_233,In_741);
or U607 (N_607,In_566,In_288);
nand U608 (N_608,In_688,In_21);
nor U609 (N_609,In_630,In_705);
or U610 (N_610,In_28,In_318);
nor U611 (N_611,In_497,In_741);
or U612 (N_612,In_495,In_342);
and U613 (N_613,In_342,In_373);
or U614 (N_614,In_428,In_71);
or U615 (N_615,In_423,In_471);
nand U616 (N_616,In_571,In_384);
and U617 (N_617,In_87,In_358);
or U618 (N_618,In_55,In_338);
nor U619 (N_619,In_92,In_532);
or U620 (N_620,In_340,In_480);
nand U621 (N_621,In_209,In_740);
nor U622 (N_622,In_223,In_520);
nand U623 (N_623,In_731,In_172);
nand U624 (N_624,In_279,In_240);
nor U625 (N_625,In_625,In_318);
and U626 (N_626,In_743,In_356);
nand U627 (N_627,In_659,In_492);
nand U628 (N_628,In_184,In_670);
or U629 (N_629,In_529,In_643);
and U630 (N_630,In_129,In_302);
and U631 (N_631,In_728,In_447);
or U632 (N_632,In_318,In_176);
nand U633 (N_633,In_569,In_26);
or U634 (N_634,In_2,In_435);
nand U635 (N_635,In_73,In_210);
and U636 (N_636,In_640,In_666);
nand U637 (N_637,In_503,In_32);
or U638 (N_638,In_292,In_335);
nor U639 (N_639,In_325,In_14);
and U640 (N_640,In_481,In_730);
and U641 (N_641,In_518,In_342);
nor U642 (N_642,In_262,In_398);
or U643 (N_643,In_213,In_134);
or U644 (N_644,In_111,In_15);
or U645 (N_645,In_264,In_31);
nor U646 (N_646,In_480,In_273);
nor U647 (N_647,In_569,In_599);
and U648 (N_648,In_81,In_170);
and U649 (N_649,In_636,In_677);
nor U650 (N_650,In_302,In_469);
nor U651 (N_651,In_264,In_382);
nand U652 (N_652,In_597,In_674);
or U653 (N_653,In_258,In_272);
nand U654 (N_654,In_609,In_161);
nand U655 (N_655,In_562,In_299);
nor U656 (N_656,In_580,In_115);
and U657 (N_657,In_367,In_22);
nand U658 (N_658,In_371,In_7);
nand U659 (N_659,In_715,In_37);
nor U660 (N_660,In_435,In_50);
or U661 (N_661,In_212,In_315);
nor U662 (N_662,In_126,In_230);
or U663 (N_663,In_556,In_622);
nor U664 (N_664,In_105,In_127);
nand U665 (N_665,In_192,In_155);
or U666 (N_666,In_112,In_622);
and U667 (N_667,In_24,In_191);
nor U668 (N_668,In_476,In_571);
or U669 (N_669,In_281,In_548);
and U670 (N_670,In_430,In_674);
nor U671 (N_671,In_106,In_312);
or U672 (N_672,In_405,In_217);
and U673 (N_673,In_489,In_14);
nand U674 (N_674,In_360,In_672);
xor U675 (N_675,In_170,In_167);
and U676 (N_676,In_693,In_533);
nor U677 (N_677,In_560,In_142);
or U678 (N_678,In_130,In_433);
or U679 (N_679,In_723,In_466);
xnor U680 (N_680,In_403,In_320);
nor U681 (N_681,In_523,In_723);
or U682 (N_682,In_4,In_44);
and U683 (N_683,In_470,In_522);
and U684 (N_684,In_123,In_390);
or U685 (N_685,In_664,In_206);
and U686 (N_686,In_564,In_32);
or U687 (N_687,In_257,In_365);
nor U688 (N_688,In_66,In_361);
nor U689 (N_689,In_225,In_324);
nor U690 (N_690,In_245,In_451);
nor U691 (N_691,In_504,In_333);
and U692 (N_692,In_448,In_219);
nor U693 (N_693,In_129,In_726);
nor U694 (N_694,In_474,In_446);
nand U695 (N_695,In_489,In_565);
and U696 (N_696,In_423,In_501);
and U697 (N_697,In_182,In_322);
nor U698 (N_698,In_41,In_475);
or U699 (N_699,In_382,In_508);
and U700 (N_700,In_572,In_57);
or U701 (N_701,In_306,In_71);
or U702 (N_702,In_564,In_329);
nand U703 (N_703,In_619,In_86);
xor U704 (N_704,In_360,In_511);
and U705 (N_705,In_412,In_532);
and U706 (N_706,In_413,In_251);
nand U707 (N_707,In_682,In_327);
nand U708 (N_708,In_551,In_358);
or U709 (N_709,In_614,In_250);
nand U710 (N_710,In_648,In_152);
and U711 (N_711,In_415,In_493);
nor U712 (N_712,In_55,In_349);
or U713 (N_713,In_692,In_275);
nand U714 (N_714,In_528,In_384);
or U715 (N_715,In_613,In_488);
or U716 (N_716,In_171,In_528);
or U717 (N_717,In_546,In_693);
xnor U718 (N_718,In_71,In_434);
nor U719 (N_719,In_742,In_39);
nand U720 (N_720,In_666,In_4);
or U721 (N_721,In_604,In_685);
or U722 (N_722,In_728,In_136);
and U723 (N_723,In_399,In_436);
and U724 (N_724,In_550,In_486);
and U725 (N_725,In_77,In_482);
nand U726 (N_726,In_473,In_592);
and U727 (N_727,In_126,In_485);
and U728 (N_728,In_614,In_339);
and U729 (N_729,In_616,In_41);
or U730 (N_730,In_339,In_106);
or U731 (N_731,In_56,In_163);
or U732 (N_732,In_561,In_462);
or U733 (N_733,In_79,In_501);
nor U734 (N_734,In_320,In_559);
or U735 (N_735,In_44,In_567);
or U736 (N_736,In_298,In_733);
or U737 (N_737,In_503,In_626);
and U738 (N_738,In_193,In_388);
and U739 (N_739,In_493,In_543);
and U740 (N_740,In_324,In_646);
and U741 (N_741,In_182,In_342);
or U742 (N_742,In_118,In_685);
or U743 (N_743,In_513,In_294);
and U744 (N_744,In_242,In_625);
nor U745 (N_745,In_268,In_387);
or U746 (N_746,In_99,In_450);
and U747 (N_747,In_481,In_187);
nor U748 (N_748,In_50,In_520);
and U749 (N_749,In_171,In_39);
and U750 (N_750,In_569,In_310);
and U751 (N_751,In_118,In_289);
and U752 (N_752,In_567,In_317);
or U753 (N_753,In_152,In_1);
nor U754 (N_754,In_38,In_219);
nor U755 (N_755,In_196,In_582);
and U756 (N_756,In_262,In_514);
or U757 (N_757,In_478,In_118);
nand U758 (N_758,In_613,In_493);
nand U759 (N_759,In_325,In_608);
or U760 (N_760,In_645,In_660);
nor U761 (N_761,In_702,In_244);
xnor U762 (N_762,In_263,In_23);
and U763 (N_763,In_399,In_543);
and U764 (N_764,In_157,In_110);
and U765 (N_765,In_280,In_702);
nand U766 (N_766,In_518,In_354);
and U767 (N_767,In_648,In_569);
xor U768 (N_768,In_632,In_366);
nor U769 (N_769,In_351,In_479);
or U770 (N_770,In_709,In_727);
or U771 (N_771,In_478,In_330);
nor U772 (N_772,In_732,In_668);
nor U773 (N_773,In_243,In_9);
xnor U774 (N_774,In_388,In_734);
nor U775 (N_775,In_331,In_136);
xnor U776 (N_776,In_638,In_10);
nand U777 (N_777,In_726,In_735);
or U778 (N_778,In_676,In_231);
nor U779 (N_779,In_682,In_347);
nand U780 (N_780,In_345,In_242);
nor U781 (N_781,In_741,In_499);
and U782 (N_782,In_651,In_362);
xnor U783 (N_783,In_632,In_497);
nor U784 (N_784,In_253,In_107);
and U785 (N_785,In_405,In_389);
and U786 (N_786,In_707,In_526);
or U787 (N_787,In_188,In_489);
or U788 (N_788,In_208,In_132);
nand U789 (N_789,In_657,In_649);
nand U790 (N_790,In_471,In_72);
nand U791 (N_791,In_468,In_188);
nand U792 (N_792,In_632,In_693);
nand U793 (N_793,In_269,In_338);
or U794 (N_794,In_265,In_704);
and U795 (N_795,In_161,In_68);
or U796 (N_796,In_265,In_391);
nor U797 (N_797,In_324,In_617);
nand U798 (N_798,In_173,In_614);
or U799 (N_799,In_241,In_144);
and U800 (N_800,In_570,In_84);
nor U801 (N_801,In_719,In_83);
nor U802 (N_802,In_321,In_167);
nand U803 (N_803,In_91,In_162);
and U804 (N_804,In_625,In_147);
and U805 (N_805,In_662,In_633);
nand U806 (N_806,In_604,In_446);
and U807 (N_807,In_485,In_275);
or U808 (N_808,In_170,In_159);
nor U809 (N_809,In_33,In_53);
or U810 (N_810,In_29,In_332);
nor U811 (N_811,In_21,In_667);
or U812 (N_812,In_235,In_731);
nor U813 (N_813,In_267,In_578);
nor U814 (N_814,In_276,In_580);
or U815 (N_815,In_416,In_527);
nor U816 (N_816,In_459,In_83);
nor U817 (N_817,In_190,In_407);
nand U818 (N_818,In_437,In_283);
and U819 (N_819,In_255,In_551);
or U820 (N_820,In_543,In_18);
or U821 (N_821,In_709,In_414);
nand U822 (N_822,In_404,In_616);
and U823 (N_823,In_398,In_386);
nor U824 (N_824,In_258,In_306);
nor U825 (N_825,In_319,In_163);
and U826 (N_826,In_501,In_342);
nor U827 (N_827,In_596,In_696);
and U828 (N_828,In_230,In_668);
nand U829 (N_829,In_86,In_317);
nand U830 (N_830,In_160,In_70);
and U831 (N_831,In_339,In_252);
or U832 (N_832,In_732,In_742);
nand U833 (N_833,In_713,In_334);
nor U834 (N_834,In_162,In_571);
nand U835 (N_835,In_282,In_397);
and U836 (N_836,In_306,In_159);
nor U837 (N_837,In_45,In_655);
or U838 (N_838,In_647,In_477);
or U839 (N_839,In_174,In_743);
and U840 (N_840,In_169,In_298);
nand U841 (N_841,In_283,In_489);
nand U842 (N_842,In_63,In_541);
and U843 (N_843,In_658,In_457);
and U844 (N_844,In_380,In_506);
nand U845 (N_845,In_164,In_186);
nand U846 (N_846,In_676,In_468);
nand U847 (N_847,In_269,In_66);
nor U848 (N_848,In_700,In_218);
nor U849 (N_849,In_716,In_32);
nand U850 (N_850,In_201,In_570);
or U851 (N_851,In_641,In_392);
nand U852 (N_852,In_600,In_23);
nand U853 (N_853,In_139,In_70);
nor U854 (N_854,In_85,In_73);
nor U855 (N_855,In_408,In_484);
and U856 (N_856,In_97,In_190);
nor U857 (N_857,In_158,In_251);
nand U858 (N_858,In_294,In_474);
nor U859 (N_859,In_207,In_483);
and U860 (N_860,In_580,In_74);
or U861 (N_861,In_728,In_101);
nand U862 (N_862,In_566,In_64);
or U863 (N_863,In_367,In_666);
and U864 (N_864,In_498,In_421);
nand U865 (N_865,In_57,In_571);
or U866 (N_866,In_252,In_204);
nand U867 (N_867,In_55,In_276);
or U868 (N_868,In_45,In_256);
nor U869 (N_869,In_70,In_471);
and U870 (N_870,In_406,In_14);
and U871 (N_871,In_733,In_127);
nor U872 (N_872,In_626,In_467);
and U873 (N_873,In_598,In_561);
xnor U874 (N_874,In_137,In_28);
nand U875 (N_875,In_424,In_606);
nor U876 (N_876,In_644,In_40);
nand U877 (N_877,In_238,In_655);
and U878 (N_878,In_535,In_656);
or U879 (N_879,In_129,In_518);
nand U880 (N_880,In_40,In_115);
nor U881 (N_881,In_396,In_287);
and U882 (N_882,In_88,In_393);
nor U883 (N_883,In_212,In_432);
and U884 (N_884,In_518,In_361);
and U885 (N_885,In_583,In_318);
nand U886 (N_886,In_112,In_492);
nand U887 (N_887,In_568,In_574);
and U888 (N_888,In_684,In_592);
nand U889 (N_889,In_420,In_390);
nor U890 (N_890,In_336,In_94);
and U891 (N_891,In_705,In_603);
nand U892 (N_892,In_163,In_605);
and U893 (N_893,In_289,In_732);
and U894 (N_894,In_619,In_498);
and U895 (N_895,In_440,In_195);
nor U896 (N_896,In_444,In_683);
nand U897 (N_897,In_502,In_104);
and U898 (N_898,In_232,In_280);
and U899 (N_899,In_529,In_600);
and U900 (N_900,In_259,In_46);
nor U901 (N_901,In_660,In_100);
xnor U902 (N_902,In_312,In_205);
and U903 (N_903,In_432,In_337);
nor U904 (N_904,In_587,In_698);
or U905 (N_905,In_167,In_516);
and U906 (N_906,In_281,In_285);
or U907 (N_907,In_720,In_39);
and U908 (N_908,In_523,In_369);
nor U909 (N_909,In_452,In_540);
nor U910 (N_910,In_155,In_385);
and U911 (N_911,In_747,In_325);
or U912 (N_912,In_491,In_146);
or U913 (N_913,In_537,In_372);
xnor U914 (N_914,In_16,In_375);
nor U915 (N_915,In_744,In_601);
or U916 (N_916,In_192,In_642);
or U917 (N_917,In_624,In_186);
and U918 (N_918,In_127,In_391);
nand U919 (N_919,In_433,In_497);
or U920 (N_920,In_58,In_547);
and U921 (N_921,In_376,In_575);
and U922 (N_922,In_155,In_185);
nor U923 (N_923,In_42,In_146);
nand U924 (N_924,In_235,In_452);
nor U925 (N_925,In_93,In_675);
nand U926 (N_926,In_748,In_746);
and U927 (N_927,In_203,In_670);
or U928 (N_928,In_465,In_406);
and U929 (N_929,In_442,In_632);
nand U930 (N_930,In_340,In_21);
nand U931 (N_931,In_725,In_210);
nor U932 (N_932,In_627,In_186);
or U933 (N_933,In_603,In_422);
and U934 (N_934,In_493,In_51);
nor U935 (N_935,In_368,In_147);
or U936 (N_936,In_66,In_56);
or U937 (N_937,In_693,In_547);
or U938 (N_938,In_50,In_648);
or U939 (N_939,In_730,In_385);
nor U940 (N_940,In_271,In_385);
and U941 (N_941,In_576,In_340);
and U942 (N_942,In_264,In_278);
nor U943 (N_943,In_251,In_66);
nor U944 (N_944,In_583,In_569);
and U945 (N_945,In_58,In_670);
nor U946 (N_946,In_337,In_180);
or U947 (N_947,In_518,In_475);
and U948 (N_948,In_315,In_454);
nor U949 (N_949,In_376,In_370);
and U950 (N_950,In_655,In_549);
and U951 (N_951,In_12,In_482);
or U952 (N_952,In_88,In_93);
or U953 (N_953,In_302,In_404);
nand U954 (N_954,In_608,In_682);
or U955 (N_955,In_279,In_58);
nand U956 (N_956,In_289,In_260);
nor U957 (N_957,In_138,In_282);
or U958 (N_958,In_258,In_608);
nand U959 (N_959,In_616,In_654);
and U960 (N_960,In_137,In_416);
and U961 (N_961,In_433,In_328);
and U962 (N_962,In_173,In_570);
nor U963 (N_963,In_4,In_364);
and U964 (N_964,In_8,In_224);
and U965 (N_965,In_465,In_450);
nor U966 (N_966,In_413,In_506);
or U967 (N_967,In_478,In_233);
nor U968 (N_968,In_220,In_420);
or U969 (N_969,In_612,In_125);
nand U970 (N_970,In_571,In_195);
or U971 (N_971,In_4,In_74);
nand U972 (N_972,In_276,In_508);
and U973 (N_973,In_532,In_638);
nor U974 (N_974,In_35,In_20);
or U975 (N_975,In_305,In_430);
and U976 (N_976,In_699,In_163);
nand U977 (N_977,In_294,In_681);
and U978 (N_978,In_167,In_83);
or U979 (N_979,In_598,In_335);
or U980 (N_980,In_699,In_606);
or U981 (N_981,In_309,In_519);
and U982 (N_982,In_70,In_250);
xor U983 (N_983,In_567,In_160);
or U984 (N_984,In_362,In_175);
or U985 (N_985,In_729,In_123);
and U986 (N_986,In_625,In_95);
and U987 (N_987,In_732,In_336);
nand U988 (N_988,In_741,In_557);
nand U989 (N_989,In_627,In_404);
and U990 (N_990,In_648,In_689);
or U991 (N_991,In_383,In_521);
or U992 (N_992,In_285,In_625);
nor U993 (N_993,In_263,In_178);
nor U994 (N_994,In_503,In_413);
or U995 (N_995,In_48,In_329);
and U996 (N_996,In_215,In_586);
nor U997 (N_997,In_710,In_63);
and U998 (N_998,In_444,In_670);
or U999 (N_999,In_568,In_348);
or U1000 (N_1000,N_326,N_797);
nor U1001 (N_1001,N_397,N_337);
nor U1002 (N_1002,N_327,N_615);
nor U1003 (N_1003,N_446,N_883);
and U1004 (N_1004,N_567,N_284);
or U1005 (N_1005,N_86,N_831);
nand U1006 (N_1006,N_993,N_694);
or U1007 (N_1007,N_483,N_991);
nand U1008 (N_1008,N_411,N_714);
and U1009 (N_1009,N_51,N_468);
or U1010 (N_1010,N_642,N_335);
nand U1011 (N_1011,N_627,N_646);
or U1012 (N_1012,N_471,N_179);
and U1013 (N_1013,N_971,N_949);
nand U1014 (N_1014,N_453,N_955);
nand U1015 (N_1015,N_67,N_792);
nor U1016 (N_1016,N_681,N_264);
nand U1017 (N_1017,N_999,N_666);
and U1018 (N_1018,N_703,N_366);
or U1019 (N_1019,N_550,N_813);
or U1020 (N_1020,N_18,N_473);
nand U1021 (N_1021,N_157,N_426);
and U1022 (N_1022,N_93,N_131);
or U1023 (N_1023,N_99,N_6);
nor U1024 (N_1024,N_21,N_440);
and U1025 (N_1025,N_391,N_387);
nor U1026 (N_1026,N_619,N_765);
nand U1027 (N_1027,N_838,N_719);
and U1028 (N_1028,N_522,N_811);
and U1029 (N_1029,N_960,N_401);
nand U1030 (N_1030,N_526,N_28);
and U1031 (N_1031,N_353,N_136);
nand U1032 (N_1032,N_94,N_854);
nor U1033 (N_1033,N_599,N_501);
or U1034 (N_1034,N_965,N_520);
nand U1035 (N_1035,N_71,N_66);
nor U1036 (N_1036,N_866,N_978);
nor U1037 (N_1037,N_377,N_727);
nor U1038 (N_1038,N_995,N_459);
or U1039 (N_1039,N_92,N_114);
nor U1040 (N_1040,N_500,N_258);
or U1041 (N_1041,N_879,N_144);
nor U1042 (N_1042,N_205,N_894);
nor U1043 (N_1043,N_100,N_7);
nand U1044 (N_1044,N_933,N_887);
nand U1045 (N_1045,N_858,N_50);
nor U1046 (N_1046,N_649,N_328);
nor U1047 (N_1047,N_232,N_187);
nand U1048 (N_1048,N_689,N_862);
nor U1049 (N_1049,N_231,N_472);
and U1050 (N_1050,N_45,N_677);
nor U1051 (N_1051,N_17,N_768);
nand U1052 (N_1052,N_660,N_134);
nor U1053 (N_1053,N_626,N_464);
or U1054 (N_1054,N_530,N_569);
nand U1055 (N_1055,N_771,N_850);
nand U1056 (N_1056,N_315,N_442);
or U1057 (N_1057,N_773,N_899);
and U1058 (N_1058,N_103,N_751);
nor U1059 (N_1059,N_113,N_209);
nand U1060 (N_1060,N_212,N_553);
nor U1061 (N_1061,N_102,N_10);
and U1062 (N_1062,N_273,N_980);
or U1063 (N_1063,N_312,N_2);
or U1064 (N_1064,N_23,N_47);
or U1065 (N_1065,N_480,N_156);
nor U1066 (N_1066,N_348,N_913);
and U1067 (N_1067,N_705,N_695);
or U1068 (N_1068,N_554,N_128);
and U1069 (N_1069,N_656,N_430);
nor U1070 (N_1070,N_537,N_730);
or U1071 (N_1071,N_623,N_979);
and U1072 (N_1072,N_531,N_837);
nand U1073 (N_1073,N_517,N_344);
nand U1074 (N_1074,N_11,N_732);
and U1075 (N_1075,N_295,N_593);
nand U1076 (N_1076,N_684,N_829);
and U1077 (N_1077,N_701,N_183);
or U1078 (N_1078,N_217,N_132);
and U1079 (N_1079,N_953,N_814);
or U1080 (N_1080,N_952,N_781);
and U1081 (N_1081,N_549,N_355);
or U1082 (N_1082,N_221,N_223);
and U1083 (N_1083,N_824,N_449);
nand U1084 (N_1084,N_659,N_279);
or U1085 (N_1085,N_467,N_566);
or U1086 (N_1086,N_929,N_175);
nor U1087 (N_1087,N_176,N_213);
and U1088 (N_1088,N_84,N_91);
nor U1089 (N_1089,N_774,N_177);
or U1090 (N_1090,N_383,N_769);
nand U1091 (N_1091,N_20,N_380);
nor U1092 (N_1092,N_3,N_402);
nor U1093 (N_1093,N_885,N_72);
and U1094 (N_1094,N_687,N_713);
and U1095 (N_1095,N_535,N_462);
nand U1096 (N_1096,N_195,N_29);
nor U1097 (N_1097,N_547,N_492);
nand U1098 (N_1098,N_789,N_634);
nor U1099 (N_1099,N_403,N_149);
or U1100 (N_1100,N_637,N_386);
or U1101 (N_1101,N_470,N_924);
or U1102 (N_1102,N_935,N_834);
nor U1103 (N_1103,N_55,N_880);
and U1104 (N_1104,N_840,N_428);
nor U1105 (N_1105,N_692,N_388);
nor U1106 (N_1106,N_643,N_297);
nand U1107 (N_1107,N_307,N_350);
nand U1108 (N_1108,N_267,N_389);
or U1109 (N_1109,N_153,N_243);
or U1110 (N_1110,N_305,N_256);
or U1111 (N_1111,N_359,N_529);
nor U1112 (N_1112,N_252,N_787);
and U1113 (N_1113,N_145,N_25);
nand U1114 (N_1114,N_966,N_658);
nor U1115 (N_1115,N_793,N_393);
and U1116 (N_1116,N_786,N_720);
and U1117 (N_1117,N_191,N_673);
nor U1118 (N_1118,N_998,N_609);
or U1119 (N_1119,N_400,N_877);
and U1120 (N_1120,N_320,N_461);
nor U1121 (N_1121,N_667,N_89);
nand U1122 (N_1122,N_543,N_541);
or U1123 (N_1123,N_715,N_976);
nor U1124 (N_1124,N_192,N_909);
or U1125 (N_1125,N_63,N_747);
nand U1126 (N_1126,N_9,N_122);
and U1127 (N_1127,N_802,N_404);
nor U1128 (N_1128,N_398,N_882);
nand U1129 (N_1129,N_240,N_417);
nand U1130 (N_1130,N_488,N_85);
or U1131 (N_1131,N_260,N_38);
and U1132 (N_1132,N_836,N_281);
and U1133 (N_1133,N_286,N_928);
or U1134 (N_1134,N_853,N_280);
and U1135 (N_1135,N_572,N_871);
nor U1136 (N_1136,N_598,N_839);
xor U1137 (N_1137,N_448,N_241);
or U1138 (N_1138,N_653,N_324);
nand U1139 (N_1139,N_206,N_641);
nor U1140 (N_1140,N_861,N_395);
and U1141 (N_1141,N_819,N_557);
and U1142 (N_1142,N_251,N_319);
nand U1143 (N_1143,N_437,N_515);
or U1144 (N_1144,N_847,N_772);
and U1145 (N_1145,N_538,N_675);
nand U1146 (N_1146,N_717,N_982);
nor U1147 (N_1147,N_498,N_788);
nor U1148 (N_1148,N_146,N_601);
or U1149 (N_1149,N_565,N_941);
nand U1150 (N_1150,N_575,N_578);
nor U1151 (N_1151,N_101,N_372);
nand U1152 (N_1152,N_19,N_345);
nor U1153 (N_1153,N_314,N_943);
nor U1154 (N_1154,N_974,N_680);
and U1155 (N_1155,N_794,N_670);
or U1156 (N_1156,N_382,N_934);
nor U1157 (N_1157,N_548,N_561);
nor U1158 (N_1158,N_203,N_210);
or U1159 (N_1159,N_621,N_672);
nor U1160 (N_1160,N_64,N_215);
and U1161 (N_1161,N_186,N_560);
and U1162 (N_1162,N_5,N_647);
nand U1163 (N_1163,N_800,N_571);
and U1164 (N_1164,N_607,N_140);
nor U1165 (N_1165,N_945,N_964);
nor U1166 (N_1166,N_590,N_151);
or U1167 (N_1167,N_616,N_475);
or U1168 (N_1168,N_117,N_988);
and U1169 (N_1169,N_235,N_617);
nand U1170 (N_1170,N_851,N_583);
or U1171 (N_1171,N_37,N_639);
nor U1172 (N_1172,N_52,N_920);
nand U1173 (N_1173,N_779,N_484);
or U1174 (N_1174,N_247,N_669);
and U1175 (N_1175,N_174,N_518);
nor U1176 (N_1176,N_584,N_152);
nor U1177 (N_1177,N_527,N_271);
nand U1178 (N_1178,N_302,N_166);
or U1179 (N_1179,N_61,N_586);
nor U1180 (N_1180,N_644,N_849);
or U1181 (N_1181,N_226,N_276);
nand U1182 (N_1182,N_904,N_13);
nand U1183 (N_1183,N_168,N_313);
nand U1184 (N_1184,N_334,N_80);
or U1185 (N_1185,N_233,N_514);
nand U1186 (N_1186,N_88,N_375);
and U1187 (N_1187,N_27,N_494);
and U1188 (N_1188,N_546,N_886);
and U1189 (N_1189,N_754,N_652);
and U1190 (N_1190,N_390,N_524);
nand U1191 (N_1191,N_722,N_507);
and U1192 (N_1192,N_936,N_568);
nor U1193 (N_1193,N_265,N_758);
or U1194 (N_1194,N_482,N_620);
nand U1195 (N_1195,N_463,N_984);
nor U1196 (N_1196,N_97,N_511);
and U1197 (N_1197,N_458,N_229);
nand U1198 (N_1198,N_989,N_762);
and U1199 (N_1199,N_436,N_782);
or U1200 (N_1200,N_288,N_98);
or U1201 (N_1201,N_962,N_664);
nor U1202 (N_1202,N_413,N_182);
or U1203 (N_1203,N_870,N_30);
nand U1204 (N_1204,N_912,N_107);
and U1205 (N_1205,N_476,N_594);
and U1206 (N_1206,N_369,N_981);
nor U1207 (N_1207,N_190,N_384);
nor U1208 (N_1208,N_255,N_169);
nor U1209 (N_1209,N_650,N_60);
nor U1210 (N_1210,N_333,N_282);
nor U1211 (N_1211,N_491,N_330);
nor U1212 (N_1212,N_946,N_274);
nor U1213 (N_1213,N_15,N_211);
nand U1214 (N_1214,N_683,N_542);
or U1215 (N_1215,N_582,N_490);
or U1216 (N_1216,N_311,N_833);
or U1217 (N_1217,N_825,N_749);
xor U1218 (N_1218,N_285,N_361);
and U1219 (N_1219,N_58,N_42);
nor U1220 (N_1220,N_801,N_668);
and U1221 (N_1221,N_931,N_706);
nor U1222 (N_1222,N_775,N_505);
nor U1223 (N_1223,N_611,N_742);
nor U1224 (N_1224,N_126,N_671);
nand U1225 (N_1225,N_306,N_465);
or U1226 (N_1226,N_352,N_194);
and U1227 (N_1227,N_59,N_865);
or U1228 (N_1228,N_248,N_351);
nor U1229 (N_1229,N_0,N_910);
and U1230 (N_1230,N_693,N_605);
nor U1231 (N_1231,N_696,N_452);
and U1232 (N_1232,N_164,N_208);
and U1233 (N_1233,N_112,N_418);
or U1234 (N_1234,N_34,N_489);
or U1235 (N_1235,N_610,N_767);
and U1236 (N_1236,N_371,N_301);
nand U1237 (N_1237,N_405,N_784);
nor U1238 (N_1238,N_394,N_581);
or U1239 (N_1239,N_44,N_678);
nand U1240 (N_1240,N_227,N_648);
or U1241 (N_1241,N_43,N_421);
and U1242 (N_1242,N_602,N_911);
and U1243 (N_1243,N_821,N_869);
nand U1244 (N_1244,N_368,N_597);
nand U1245 (N_1245,N_26,N_396);
nand U1246 (N_1246,N_777,N_143);
or U1247 (N_1247,N_835,N_874);
nor U1248 (N_1248,N_392,N_329);
or U1249 (N_1249,N_937,N_996);
nand U1250 (N_1250,N_116,N_662);
nor U1251 (N_1251,N_622,N_291);
nand U1252 (N_1252,N_173,N_625);
nor U1253 (N_1253,N_890,N_354);
or U1254 (N_1254,N_545,N_65);
nor U1255 (N_1255,N_796,N_133);
or U1256 (N_1256,N_932,N_339);
or U1257 (N_1257,N_70,N_457);
nor U1258 (N_1258,N_534,N_532);
nor U1259 (N_1259,N_69,N_275);
nor U1260 (N_1260,N_105,N_414);
or U1261 (N_1261,N_77,N_555);
nand U1262 (N_1262,N_444,N_363);
nor U1263 (N_1263,N_709,N_863);
nand U1264 (N_1264,N_519,N_24);
nand U1265 (N_1265,N_528,N_939);
or U1266 (N_1266,N_573,N_129);
and U1267 (N_1267,N_419,N_270);
and U1268 (N_1268,N_33,N_655);
or U1269 (N_1269,N_737,N_299);
nor U1270 (N_1270,N_663,N_525);
or U1271 (N_1271,N_272,N_188);
or U1272 (N_1272,N_111,N_635);
nor U1273 (N_1273,N_222,N_921);
nand U1274 (N_1274,N_540,N_466);
nand U1275 (N_1275,N_234,N_138);
nor U1276 (N_1276,N_53,N_916);
or U1277 (N_1277,N_806,N_172);
and U1278 (N_1278,N_496,N_987);
nor U1279 (N_1279,N_917,N_477);
or U1280 (N_1280,N_373,N_410);
nand U1281 (N_1281,N_367,N_218);
or U1282 (N_1282,N_805,N_115);
nor U1283 (N_1283,N_125,N_764);
or U1284 (N_1284,N_592,N_385);
nand U1285 (N_1285,N_985,N_87);
and U1286 (N_1286,N_603,N_219);
nor U1287 (N_1287,N_926,N_596);
or U1288 (N_1288,N_556,N_406);
and U1289 (N_1289,N_481,N_803);
or U1290 (N_1290,N_278,N_124);
nor U1291 (N_1291,N_283,N_898);
nand U1292 (N_1292,N_559,N_293);
nor U1293 (N_1293,N_576,N_159);
or U1294 (N_1294,N_432,N_558);
xor U1295 (N_1295,N_628,N_588);
xor U1296 (N_1296,N_262,N_127);
or U1297 (N_1297,N_901,N_657);
and U1298 (N_1298,N_225,N_726);
nand U1299 (N_1299,N_755,N_171);
nor U1300 (N_1300,N_249,N_407);
nand U1301 (N_1301,N_748,N_508);
nand U1302 (N_1302,N_358,N_318);
nor U1303 (N_1303,N_947,N_416);
nor U1304 (N_1304,N_679,N_296);
and U1305 (N_1305,N_848,N_736);
nand U1306 (N_1306,N_298,N_940);
nor U1307 (N_1307,N_544,N_474);
nand U1308 (N_1308,N_81,N_346);
or U1309 (N_1309,N_728,N_257);
or U1310 (N_1310,N_253,N_763);
nand U1311 (N_1311,N_563,N_486);
and U1312 (N_1312,N_614,N_76);
and U1313 (N_1313,N_704,N_741);
nor U1314 (N_1314,N_927,N_859);
and U1315 (N_1315,N_710,N_820);
and U1316 (N_1316,N_365,N_423);
or U1317 (N_1317,N_948,N_493);
nand U1318 (N_1318,N_739,N_14);
nand U1319 (N_1319,N_973,N_503);
or U1320 (N_1320,N_56,N_332);
and U1321 (N_1321,N_236,N_487);
nor U1322 (N_1322,N_110,N_746);
and U1323 (N_1323,N_817,N_155);
and U1324 (N_1324,N_198,N_54);
and U1325 (N_1325,N_857,N_700);
nor U1326 (N_1326,N_431,N_31);
nor U1327 (N_1327,N_591,N_983);
nor U1328 (N_1328,N_433,N_816);
nand U1329 (N_1329,N_150,N_686);
nand U1330 (N_1330,N_629,N_364);
nand U1331 (N_1331,N_734,N_896);
nor U1332 (N_1332,N_950,N_304);
and U1333 (N_1333,N_676,N_161);
or U1334 (N_1334,N_277,N_577);
nor U1335 (N_1335,N_712,N_897);
and U1336 (N_1336,N_261,N_310);
and U1337 (N_1337,N_914,N_180);
nand U1338 (N_1338,N_731,N_562);
or U1339 (N_1339,N_994,N_197);
nand U1340 (N_1340,N_908,N_992);
and U1341 (N_1341,N_269,N_756);
and U1342 (N_1342,N_699,N_323);
and U1343 (N_1343,N_809,N_83);
nand U1344 (N_1344,N_986,N_972);
and U1345 (N_1345,N_944,N_82);
and U1346 (N_1346,N_918,N_743);
or U1347 (N_1347,N_199,N_753);
nor U1348 (N_1348,N_162,N_200);
and U1349 (N_1349,N_178,N_967);
xnor U1350 (N_1350,N_435,N_903);
nor U1351 (N_1351,N_815,N_340);
nor U1352 (N_1352,N_303,N_420);
nor U1353 (N_1353,N_504,N_970);
and U1354 (N_1354,N_141,N_422);
nor U1355 (N_1355,N_266,N_32);
nor U1356 (N_1356,N_872,N_638);
and U1357 (N_1357,N_895,N_954);
and U1358 (N_1358,N_580,N_427);
nor U1359 (N_1359,N_938,N_73);
nor U1360 (N_1360,N_68,N_119);
and U1361 (N_1361,N_708,N_724);
and U1362 (N_1362,N_875,N_244);
nor U1363 (N_1363,N_370,N_163);
nor U1364 (N_1364,N_90,N_977);
and U1365 (N_1365,N_864,N_968);
or U1366 (N_1366,N_881,N_893);
or U1367 (N_1367,N_798,N_376);
or U1368 (N_1368,N_104,N_711);
and U1369 (N_1369,N_841,N_95);
or U1370 (N_1370,N_624,N_828);
nor U1371 (N_1371,N_795,N_661);
nor U1372 (N_1372,N_1,N_79);
nor U1373 (N_1373,N_922,N_915);
nand U1374 (N_1374,N_723,N_204);
nor U1375 (N_1375,N_441,N_439);
nor U1376 (N_1376,N_612,N_536);
and U1377 (N_1377,N_469,N_189);
nor U1378 (N_1378,N_900,N_147);
or U1379 (N_1379,N_654,N_499);
or U1380 (N_1380,N_842,N_287);
or U1381 (N_1381,N_259,N_497);
or U1382 (N_1382,N_832,N_878);
and U1383 (N_1383,N_357,N_292);
nand U1384 (N_1384,N_740,N_160);
or U1385 (N_1385,N_845,N_956);
nand U1386 (N_1386,N_135,N_347);
or U1387 (N_1387,N_242,N_509);
nor U1388 (N_1388,N_716,N_108);
xnor U1389 (N_1389,N_207,N_343);
nor U1390 (N_1390,N_826,N_906);
and U1391 (N_1391,N_379,N_889);
nand U1392 (N_1392,N_139,N_856);
and U1393 (N_1393,N_109,N_807);
or U1394 (N_1394,N_697,N_338);
nor U1395 (N_1395,N_516,N_49);
nand U1396 (N_1396,N_925,N_137);
or U1397 (N_1397,N_760,N_969);
nand U1398 (N_1398,N_636,N_237);
nor U1399 (N_1399,N_429,N_4);
nor U1400 (N_1400,N_818,N_785);
nor U1401 (N_1401,N_513,N_224);
nor U1402 (N_1402,N_214,N_674);
nand U1403 (N_1403,N_378,N_263);
nor U1404 (N_1404,N_812,N_778);
nor U1405 (N_1405,N_951,N_239);
or U1406 (N_1406,N_539,N_963);
or U1407 (N_1407,N_595,N_827);
or U1408 (N_1408,N_40,N_184);
nand U1409 (N_1409,N_632,N_574);
nor U1410 (N_1410,N_451,N_640);
nor U1411 (N_1411,N_645,N_254);
nand U1412 (N_1412,N_852,N_822);
nand U1413 (N_1413,N_733,N_551);
nand U1414 (N_1414,N_246,N_447);
nand U1415 (N_1415,N_485,N_454);
nand U1416 (N_1416,N_185,N_399);
xor U1417 (N_1417,N_478,N_957);
and U1418 (N_1418,N_691,N_961);
and U1419 (N_1419,N_325,N_631);
and U1420 (N_1420,N_589,N_290);
and U1421 (N_1421,N_445,N_876);
or U1422 (N_1422,N_342,N_606);
nand U1423 (N_1423,N_721,N_682);
nand U1424 (N_1424,N_118,N_362);
or U1425 (N_1425,N_181,N_250);
nor U1426 (N_1426,N_230,N_321);
nor U1427 (N_1427,N_62,N_780);
and U1428 (N_1428,N_201,N_506);
or U1429 (N_1429,N_245,N_142);
nor U1430 (N_1430,N_381,N_804);
or U1431 (N_1431,N_823,N_349);
nand U1432 (N_1432,N_867,N_46);
or U1433 (N_1433,N_570,N_356);
nor U1434 (N_1434,N_608,N_873);
or U1435 (N_1435,N_604,N_630);
and U1436 (N_1436,N_322,N_438);
or U1437 (N_1437,N_930,N_39);
nor U1438 (N_1438,N_220,N_512);
nand U1439 (N_1439,N_336,N_759);
or U1440 (N_1440,N_533,N_702);
and U1441 (N_1441,N_331,N_860);
and U1442 (N_1442,N_341,N_975);
nor U1443 (N_1443,N_434,N_868);
and U1444 (N_1444,N_425,N_300);
nand U1445 (N_1445,N_735,N_238);
or U1446 (N_1446,N_923,N_106);
nand U1447 (N_1447,N_317,N_729);
and U1448 (N_1448,N_587,N_744);
nand U1449 (N_1449,N_997,N_718);
nor U1450 (N_1450,N_202,N_665);
or U1451 (N_1451,N_750,N_552);
or U1452 (N_1452,N_57,N_690);
and U1453 (N_1453,N_855,N_450);
or U1454 (N_1454,N_770,N_745);
nor U1455 (N_1455,N_844,N_830);
nor U1456 (N_1456,N_791,N_959);
xor U1457 (N_1457,N_167,N_651);
and U1458 (N_1458,N_48,N_309);
nand U1459 (N_1459,N_752,N_409);
xnor U1460 (N_1460,N_74,N_698);
or U1461 (N_1461,N_600,N_158);
nor U1462 (N_1462,N_902,N_685);
or U1463 (N_1463,N_810,N_585);
or U1464 (N_1464,N_130,N_907);
and U1465 (N_1465,N_766,N_120);
nand U1466 (N_1466,N_360,N_165);
nor U1467 (N_1467,N_564,N_148);
nand U1468 (N_1468,N_884,N_846);
and U1469 (N_1469,N_41,N_123);
nand U1470 (N_1470,N_502,N_216);
nand U1471 (N_1471,N_843,N_308);
nor U1472 (N_1472,N_268,N_415);
or U1473 (N_1473,N_289,N_8);
nor U1474 (N_1474,N_294,N_75);
and U1475 (N_1475,N_193,N_613);
and U1476 (N_1476,N_688,N_990);
nand U1477 (N_1477,N_412,N_761);
nand U1478 (N_1478,N_408,N_776);
nand U1479 (N_1479,N_170,N_78);
xnor U1480 (N_1480,N_374,N_460);
or U1481 (N_1481,N_799,N_443);
nor U1482 (N_1482,N_228,N_783);
nor U1483 (N_1483,N_942,N_808);
and U1484 (N_1484,N_96,N_35);
or U1485 (N_1485,N_16,N_757);
nand U1486 (N_1486,N_790,N_479);
and U1487 (N_1487,N_633,N_456);
and U1488 (N_1488,N_905,N_424);
nor U1489 (N_1489,N_22,N_12);
nand U1490 (N_1490,N_725,N_958);
nand U1491 (N_1491,N_121,N_738);
and U1492 (N_1492,N_618,N_892);
nand U1493 (N_1493,N_919,N_316);
and U1494 (N_1494,N_888,N_891);
or U1495 (N_1495,N_154,N_495);
nor U1496 (N_1496,N_523,N_707);
nand U1497 (N_1497,N_196,N_36);
or U1498 (N_1498,N_510,N_579);
and U1499 (N_1499,N_455,N_521);
and U1500 (N_1500,N_601,N_996);
nor U1501 (N_1501,N_44,N_516);
nor U1502 (N_1502,N_678,N_668);
nor U1503 (N_1503,N_957,N_279);
or U1504 (N_1504,N_524,N_223);
and U1505 (N_1505,N_981,N_491);
or U1506 (N_1506,N_794,N_592);
nand U1507 (N_1507,N_812,N_229);
nand U1508 (N_1508,N_538,N_762);
nor U1509 (N_1509,N_521,N_403);
nand U1510 (N_1510,N_214,N_338);
and U1511 (N_1511,N_315,N_840);
nand U1512 (N_1512,N_772,N_353);
and U1513 (N_1513,N_27,N_647);
nor U1514 (N_1514,N_392,N_641);
nor U1515 (N_1515,N_172,N_718);
nor U1516 (N_1516,N_562,N_230);
nand U1517 (N_1517,N_27,N_759);
nor U1518 (N_1518,N_531,N_113);
or U1519 (N_1519,N_268,N_830);
nor U1520 (N_1520,N_790,N_617);
or U1521 (N_1521,N_549,N_287);
nor U1522 (N_1522,N_598,N_648);
nor U1523 (N_1523,N_504,N_300);
nand U1524 (N_1524,N_168,N_591);
and U1525 (N_1525,N_630,N_784);
or U1526 (N_1526,N_854,N_600);
or U1527 (N_1527,N_787,N_261);
or U1528 (N_1528,N_909,N_496);
nor U1529 (N_1529,N_565,N_269);
or U1530 (N_1530,N_67,N_944);
nor U1531 (N_1531,N_465,N_959);
nor U1532 (N_1532,N_522,N_301);
nand U1533 (N_1533,N_203,N_534);
nand U1534 (N_1534,N_441,N_876);
and U1535 (N_1535,N_682,N_978);
nand U1536 (N_1536,N_935,N_640);
nand U1537 (N_1537,N_557,N_991);
and U1538 (N_1538,N_473,N_259);
or U1539 (N_1539,N_972,N_133);
nor U1540 (N_1540,N_883,N_630);
or U1541 (N_1541,N_541,N_366);
nand U1542 (N_1542,N_451,N_380);
nor U1543 (N_1543,N_389,N_827);
and U1544 (N_1544,N_132,N_722);
nor U1545 (N_1545,N_271,N_45);
nor U1546 (N_1546,N_279,N_623);
and U1547 (N_1547,N_252,N_809);
nor U1548 (N_1548,N_788,N_105);
nand U1549 (N_1549,N_855,N_431);
and U1550 (N_1550,N_501,N_691);
or U1551 (N_1551,N_234,N_722);
nor U1552 (N_1552,N_330,N_301);
nand U1553 (N_1553,N_353,N_769);
or U1554 (N_1554,N_433,N_748);
or U1555 (N_1555,N_513,N_191);
nor U1556 (N_1556,N_758,N_203);
or U1557 (N_1557,N_281,N_976);
nor U1558 (N_1558,N_182,N_12);
nand U1559 (N_1559,N_694,N_278);
nand U1560 (N_1560,N_551,N_421);
and U1561 (N_1561,N_936,N_898);
or U1562 (N_1562,N_638,N_253);
nor U1563 (N_1563,N_862,N_915);
and U1564 (N_1564,N_563,N_131);
nand U1565 (N_1565,N_63,N_219);
nand U1566 (N_1566,N_385,N_942);
or U1567 (N_1567,N_593,N_312);
nor U1568 (N_1568,N_691,N_529);
nand U1569 (N_1569,N_798,N_48);
nor U1570 (N_1570,N_774,N_426);
and U1571 (N_1571,N_476,N_312);
nor U1572 (N_1572,N_250,N_505);
and U1573 (N_1573,N_444,N_435);
nand U1574 (N_1574,N_456,N_919);
or U1575 (N_1575,N_36,N_429);
nor U1576 (N_1576,N_430,N_687);
and U1577 (N_1577,N_189,N_186);
nand U1578 (N_1578,N_503,N_409);
and U1579 (N_1579,N_753,N_604);
nor U1580 (N_1580,N_988,N_31);
nand U1581 (N_1581,N_562,N_938);
and U1582 (N_1582,N_402,N_459);
nor U1583 (N_1583,N_444,N_101);
or U1584 (N_1584,N_258,N_856);
nor U1585 (N_1585,N_999,N_348);
nor U1586 (N_1586,N_640,N_767);
and U1587 (N_1587,N_649,N_295);
or U1588 (N_1588,N_885,N_645);
and U1589 (N_1589,N_424,N_356);
nand U1590 (N_1590,N_765,N_723);
or U1591 (N_1591,N_226,N_465);
and U1592 (N_1592,N_176,N_757);
or U1593 (N_1593,N_586,N_308);
and U1594 (N_1594,N_628,N_340);
nand U1595 (N_1595,N_418,N_57);
or U1596 (N_1596,N_531,N_155);
nand U1597 (N_1597,N_714,N_632);
or U1598 (N_1598,N_630,N_124);
nand U1599 (N_1599,N_954,N_15);
nor U1600 (N_1600,N_410,N_91);
nand U1601 (N_1601,N_708,N_505);
nand U1602 (N_1602,N_251,N_363);
or U1603 (N_1603,N_583,N_711);
nor U1604 (N_1604,N_290,N_998);
and U1605 (N_1605,N_797,N_159);
nor U1606 (N_1606,N_434,N_114);
nand U1607 (N_1607,N_270,N_843);
nor U1608 (N_1608,N_358,N_84);
nand U1609 (N_1609,N_415,N_596);
and U1610 (N_1610,N_97,N_619);
or U1611 (N_1611,N_589,N_524);
and U1612 (N_1612,N_310,N_263);
nor U1613 (N_1613,N_966,N_801);
and U1614 (N_1614,N_954,N_860);
nor U1615 (N_1615,N_595,N_708);
nor U1616 (N_1616,N_550,N_963);
and U1617 (N_1617,N_371,N_198);
nor U1618 (N_1618,N_306,N_36);
or U1619 (N_1619,N_744,N_295);
and U1620 (N_1620,N_843,N_356);
nor U1621 (N_1621,N_331,N_562);
and U1622 (N_1622,N_574,N_430);
and U1623 (N_1623,N_417,N_95);
and U1624 (N_1624,N_19,N_577);
nand U1625 (N_1625,N_710,N_333);
nor U1626 (N_1626,N_203,N_739);
nor U1627 (N_1627,N_975,N_318);
or U1628 (N_1628,N_910,N_698);
nor U1629 (N_1629,N_659,N_87);
or U1630 (N_1630,N_87,N_482);
and U1631 (N_1631,N_450,N_820);
nor U1632 (N_1632,N_265,N_620);
xor U1633 (N_1633,N_308,N_367);
and U1634 (N_1634,N_50,N_439);
nand U1635 (N_1635,N_259,N_12);
nor U1636 (N_1636,N_29,N_787);
nand U1637 (N_1637,N_204,N_993);
nand U1638 (N_1638,N_47,N_438);
nand U1639 (N_1639,N_617,N_351);
or U1640 (N_1640,N_59,N_168);
nor U1641 (N_1641,N_106,N_857);
and U1642 (N_1642,N_897,N_804);
and U1643 (N_1643,N_963,N_155);
or U1644 (N_1644,N_521,N_752);
nand U1645 (N_1645,N_564,N_823);
or U1646 (N_1646,N_116,N_9);
nor U1647 (N_1647,N_589,N_997);
nand U1648 (N_1648,N_928,N_883);
or U1649 (N_1649,N_198,N_703);
nor U1650 (N_1650,N_746,N_369);
nand U1651 (N_1651,N_516,N_763);
and U1652 (N_1652,N_221,N_17);
or U1653 (N_1653,N_806,N_241);
or U1654 (N_1654,N_395,N_321);
or U1655 (N_1655,N_561,N_113);
and U1656 (N_1656,N_328,N_251);
nor U1657 (N_1657,N_983,N_773);
and U1658 (N_1658,N_245,N_5);
and U1659 (N_1659,N_192,N_231);
or U1660 (N_1660,N_423,N_65);
nand U1661 (N_1661,N_741,N_651);
and U1662 (N_1662,N_890,N_258);
and U1663 (N_1663,N_555,N_530);
or U1664 (N_1664,N_222,N_128);
nand U1665 (N_1665,N_332,N_662);
and U1666 (N_1666,N_826,N_334);
and U1667 (N_1667,N_114,N_837);
or U1668 (N_1668,N_593,N_546);
nor U1669 (N_1669,N_91,N_650);
nor U1670 (N_1670,N_870,N_787);
nand U1671 (N_1671,N_215,N_118);
or U1672 (N_1672,N_485,N_947);
and U1673 (N_1673,N_916,N_131);
and U1674 (N_1674,N_800,N_132);
or U1675 (N_1675,N_521,N_330);
or U1676 (N_1676,N_557,N_288);
nor U1677 (N_1677,N_498,N_938);
nand U1678 (N_1678,N_152,N_504);
and U1679 (N_1679,N_47,N_874);
nand U1680 (N_1680,N_140,N_435);
nand U1681 (N_1681,N_812,N_627);
nand U1682 (N_1682,N_0,N_10);
nand U1683 (N_1683,N_96,N_864);
nand U1684 (N_1684,N_327,N_640);
nor U1685 (N_1685,N_78,N_184);
nor U1686 (N_1686,N_761,N_9);
or U1687 (N_1687,N_496,N_479);
or U1688 (N_1688,N_415,N_930);
nand U1689 (N_1689,N_314,N_106);
or U1690 (N_1690,N_82,N_235);
nor U1691 (N_1691,N_608,N_278);
nor U1692 (N_1692,N_755,N_330);
nor U1693 (N_1693,N_383,N_850);
nand U1694 (N_1694,N_937,N_822);
nor U1695 (N_1695,N_798,N_270);
nor U1696 (N_1696,N_667,N_97);
and U1697 (N_1697,N_777,N_556);
nor U1698 (N_1698,N_601,N_220);
nand U1699 (N_1699,N_669,N_627);
nand U1700 (N_1700,N_699,N_547);
nor U1701 (N_1701,N_740,N_42);
nand U1702 (N_1702,N_185,N_734);
or U1703 (N_1703,N_218,N_8);
nor U1704 (N_1704,N_901,N_331);
nor U1705 (N_1705,N_397,N_888);
or U1706 (N_1706,N_934,N_610);
xnor U1707 (N_1707,N_666,N_719);
nand U1708 (N_1708,N_743,N_74);
and U1709 (N_1709,N_362,N_636);
nor U1710 (N_1710,N_318,N_189);
or U1711 (N_1711,N_698,N_562);
or U1712 (N_1712,N_782,N_809);
and U1713 (N_1713,N_498,N_117);
or U1714 (N_1714,N_318,N_699);
nand U1715 (N_1715,N_620,N_776);
nand U1716 (N_1716,N_14,N_722);
nand U1717 (N_1717,N_779,N_569);
and U1718 (N_1718,N_40,N_333);
nor U1719 (N_1719,N_446,N_521);
xor U1720 (N_1720,N_471,N_291);
and U1721 (N_1721,N_261,N_530);
nand U1722 (N_1722,N_296,N_779);
and U1723 (N_1723,N_907,N_41);
nor U1724 (N_1724,N_569,N_870);
nand U1725 (N_1725,N_738,N_329);
and U1726 (N_1726,N_924,N_442);
and U1727 (N_1727,N_474,N_966);
or U1728 (N_1728,N_298,N_931);
or U1729 (N_1729,N_836,N_344);
nand U1730 (N_1730,N_417,N_184);
nand U1731 (N_1731,N_351,N_900);
nor U1732 (N_1732,N_40,N_322);
nor U1733 (N_1733,N_345,N_35);
nand U1734 (N_1734,N_549,N_290);
nand U1735 (N_1735,N_236,N_798);
nor U1736 (N_1736,N_920,N_906);
and U1737 (N_1737,N_587,N_254);
nand U1738 (N_1738,N_339,N_707);
nor U1739 (N_1739,N_564,N_351);
or U1740 (N_1740,N_3,N_182);
or U1741 (N_1741,N_120,N_883);
nor U1742 (N_1742,N_86,N_82);
nand U1743 (N_1743,N_556,N_306);
and U1744 (N_1744,N_180,N_793);
nand U1745 (N_1745,N_892,N_656);
nor U1746 (N_1746,N_19,N_392);
nor U1747 (N_1747,N_844,N_352);
nor U1748 (N_1748,N_734,N_735);
or U1749 (N_1749,N_510,N_41);
nand U1750 (N_1750,N_128,N_944);
and U1751 (N_1751,N_29,N_174);
nor U1752 (N_1752,N_98,N_212);
and U1753 (N_1753,N_933,N_808);
nor U1754 (N_1754,N_290,N_966);
and U1755 (N_1755,N_512,N_103);
nor U1756 (N_1756,N_445,N_262);
nand U1757 (N_1757,N_638,N_704);
nor U1758 (N_1758,N_636,N_527);
nor U1759 (N_1759,N_791,N_474);
nand U1760 (N_1760,N_220,N_746);
or U1761 (N_1761,N_426,N_860);
or U1762 (N_1762,N_221,N_170);
and U1763 (N_1763,N_917,N_787);
and U1764 (N_1764,N_548,N_287);
nor U1765 (N_1765,N_275,N_595);
and U1766 (N_1766,N_753,N_282);
or U1767 (N_1767,N_304,N_332);
nand U1768 (N_1768,N_243,N_759);
nand U1769 (N_1769,N_893,N_777);
and U1770 (N_1770,N_750,N_83);
nand U1771 (N_1771,N_268,N_248);
or U1772 (N_1772,N_656,N_531);
nand U1773 (N_1773,N_979,N_795);
and U1774 (N_1774,N_704,N_548);
nand U1775 (N_1775,N_577,N_842);
nor U1776 (N_1776,N_18,N_189);
and U1777 (N_1777,N_969,N_961);
and U1778 (N_1778,N_96,N_221);
nor U1779 (N_1779,N_244,N_841);
nand U1780 (N_1780,N_300,N_768);
or U1781 (N_1781,N_941,N_763);
or U1782 (N_1782,N_125,N_11);
nor U1783 (N_1783,N_62,N_953);
nor U1784 (N_1784,N_884,N_612);
or U1785 (N_1785,N_769,N_746);
and U1786 (N_1786,N_849,N_512);
and U1787 (N_1787,N_479,N_457);
or U1788 (N_1788,N_143,N_938);
or U1789 (N_1789,N_283,N_186);
or U1790 (N_1790,N_50,N_628);
xnor U1791 (N_1791,N_560,N_35);
or U1792 (N_1792,N_35,N_989);
or U1793 (N_1793,N_175,N_252);
nor U1794 (N_1794,N_33,N_140);
xor U1795 (N_1795,N_527,N_723);
nand U1796 (N_1796,N_196,N_105);
or U1797 (N_1797,N_561,N_542);
or U1798 (N_1798,N_792,N_178);
or U1799 (N_1799,N_348,N_168);
nand U1800 (N_1800,N_903,N_503);
nand U1801 (N_1801,N_694,N_553);
nor U1802 (N_1802,N_234,N_980);
and U1803 (N_1803,N_559,N_410);
nor U1804 (N_1804,N_816,N_308);
and U1805 (N_1805,N_470,N_145);
and U1806 (N_1806,N_805,N_781);
nand U1807 (N_1807,N_2,N_162);
nor U1808 (N_1808,N_523,N_870);
nor U1809 (N_1809,N_918,N_275);
and U1810 (N_1810,N_680,N_638);
nand U1811 (N_1811,N_967,N_232);
nor U1812 (N_1812,N_738,N_466);
or U1813 (N_1813,N_271,N_587);
nor U1814 (N_1814,N_67,N_814);
nor U1815 (N_1815,N_207,N_832);
nor U1816 (N_1816,N_235,N_189);
nor U1817 (N_1817,N_718,N_943);
nor U1818 (N_1818,N_152,N_53);
and U1819 (N_1819,N_458,N_746);
or U1820 (N_1820,N_738,N_185);
and U1821 (N_1821,N_939,N_868);
nand U1822 (N_1822,N_298,N_988);
or U1823 (N_1823,N_663,N_957);
nand U1824 (N_1824,N_58,N_429);
nor U1825 (N_1825,N_610,N_99);
or U1826 (N_1826,N_961,N_985);
nand U1827 (N_1827,N_713,N_322);
or U1828 (N_1828,N_298,N_366);
nand U1829 (N_1829,N_643,N_411);
nor U1830 (N_1830,N_147,N_291);
and U1831 (N_1831,N_447,N_973);
nor U1832 (N_1832,N_804,N_888);
nor U1833 (N_1833,N_523,N_472);
and U1834 (N_1834,N_776,N_302);
and U1835 (N_1835,N_84,N_401);
and U1836 (N_1836,N_664,N_954);
or U1837 (N_1837,N_523,N_422);
nand U1838 (N_1838,N_984,N_974);
nand U1839 (N_1839,N_359,N_299);
nand U1840 (N_1840,N_265,N_801);
nand U1841 (N_1841,N_538,N_801);
and U1842 (N_1842,N_180,N_670);
nor U1843 (N_1843,N_565,N_106);
nor U1844 (N_1844,N_163,N_965);
and U1845 (N_1845,N_561,N_346);
nor U1846 (N_1846,N_896,N_517);
nand U1847 (N_1847,N_503,N_147);
and U1848 (N_1848,N_175,N_893);
nor U1849 (N_1849,N_804,N_211);
or U1850 (N_1850,N_49,N_576);
nor U1851 (N_1851,N_257,N_56);
and U1852 (N_1852,N_360,N_961);
nor U1853 (N_1853,N_458,N_66);
nor U1854 (N_1854,N_680,N_933);
or U1855 (N_1855,N_418,N_542);
and U1856 (N_1856,N_391,N_317);
or U1857 (N_1857,N_244,N_822);
or U1858 (N_1858,N_924,N_743);
and U1859 (N_1859,N_700,N_697);
or U1860 (N_1860,N_890,N_364);
or U1861 (N_1861,N_85,N_109);
and U1862 (N_1862,N_440,N_210);
nand U1863 (N_1863,N_973,N_232);
or U1864 (N_1864,N_525,N_226);
nand U1865 (N_1865,N_328,N_370);
or U1866 (N_1866,N_133,N_390);
and U1867 (N_1867,N_122,N_5);
nor U1868 (N_1868,N_627,N_833);
or U1869 (N_1869,N_407,N_707);
nor U1870 (N_1870,N_432,N_476);
nor U1871 (N_1871,N_596,N_441);
nor U1872 (N_1872,N_471,N_369);
nor U1873 (N_1873,N_745,N_367);
or U1874 (N_1874,N_944,N_338);
and U1875 (N_1875,N_396,N_535);
nor U1876 (N_1876,N_954,N_103);
or U1877 (N_1877,N_273,N_81);
and U1878 (N_1878,N_636,N_931);
nand U1879 (N_1879,N_903,N_266);
or U1880 (N_1880,N_930,N_289);
nand U1881 (N_1881,N_77,N_946);
nor U1882 (N_1882,N_954,N_566);
or U1883 (N_1883,N_257,N_120);
xor U1884 (N_1884,N_161,N_741);
nor U1885 (N_1885,N_598,N_659);
and U1886 (N_1886,N_984,N_263);
nor U1887 (N_1887,N_730,N_258);
nor U1888 (N_1888,N_495,N_552);
or U1889 (N_1889,N_323,N_139);
nor U1890 (N_1890,N_995,N_788);
nand U1891 (N_1891,N_477,N_411);
nand U1892 (N_1892,N_682,N_691);
nor U1893 (N_1893,N_664,N_335);
nand U1894 (N_1894,N_180,N_443);
or U1895 (N_1895,N_921,N_563);
and U1896 (N_1896,N_875,N_307);
and U1897 (N_1897,N_39,N_444);
or U1898 (N_1898,N_822,N_235);
and U1899 (N_1899,N_839,N_629);
nand U1900 (N_1900,N_332,N_166);
and U1901 (N_1901,N_898,N_747);
or U1902 (N_1902,N_316,N_956);
and U1903 (N_1903,N_873,N_779);
or U1904 (N_1904,N_897,N_765);
nor U1905 (N_1905,N_403,N_429);
nand U1906 (N_1906,N_437,N_24);
nor U1907 (N_1907,N_565,N_485);
or U1908 (N_1908,N_680,N_1);
nand U1909 (N_1909,N_846,N_457);
and U1910 (N_1910,N_745,N_356);
and U1911 (N_1911,N_380,N_822);
and U1912 (N_1912,N_477,N_130);
and U1913 (N_1913,N_37,N_943);
or U1914 (N_1914,N_889,N_91);
nor U1915 (N_1915,N_133,N_536);
or U1916 (N_1916,N_517,N_295);
nand U1917 (N_1917,N_953,N_882);
nand U1918 (N_1918,N_495,N_796);
nand U1919 (N_1919,N_727,N_484);
nand U1920 (N_1920,N_177,N_206);
nor U1921 (N_1921,N_341,N_700);
and U1922 (N_1922,N_803,N_27);
nor U1923 (N_1923,N_24,N_718);
or U1924 (N_1924,N_638,N_355);
and U1925 (N_1925,N_604,N_134);
and U1926 (N_1926,N_268,N_658);
or U1927 (N_1927,N_557,N_364);
nor U1928 (N_1928,N_135,N_486);
or U1929 (N_1929,N_66,N_408);
nor U1930 (N_1930,N_290,N_620);
nor U1931 (N_1931,N_301,N_977);
and U1932 (N_1932,N_659,N_738);
nand U1933 (N_1933,N_582,N_985);
or U1934 (N_1934,N_48,N_258);
nand U1935 (N_1935,N_565,N_196);
xnor U1936 (N_1936,N_799,N_234);
nand U1937 (N_1937,N_863,N_411);
and U1938 (N_1938,N_743,N_911);
or U1939 (N_1939,N_259,N_616);
or U1940 (N_1940,N_757,N_907);
xor U1941 (N_1941,N_25,N_482);
nor U1942 (N_1942,N_547,N_178);
and U1943 (N_1943,N_649,N_182);
nand U1944 (N_1944,N_649,N_64);
or U1945 (N_1945,N_734,N_51);
or U1946 (N_1946,N_111,N_949);
and U1947 (N_1947,N_966,N_436);
xnor U1948 (N_1948,N_618,N_21);
or U1949 (N_1949,N_97,N_287);
nand U1950 (N_1950,N_745,N_663);
and U1951 (N_1951,N_579,N_571);
and U1952 (N_1952,N_643,N_177);
nor U1953 (N_1953,N_512,N_699);
or U1954 (N_1954,N_732,N_862);
nand U1955 (N_1955,N_837,N_888);
and U1956 (N_1956,N_643,N_732);
nor U1957 (N_1957,N_151,N_167);
nor U1958 (N_1958,N_968,N_548);
nand U1959 (N_1959,N_11,N_407);
nand U1960 (N_1960,N_706,N_500);
and U1961 (N_1961,N_675,N_364);
nand U1962 (N_1962,N_197,N_382);
and U1963 (N_1963,N_278,N_659);
and U1964 (N_1964,N_833,N_683);
nand U1965 (N_1965,N_560,N_61);
or U1966 (N_1966,N_450,N_38);
nor U1967 (N_1967,N_698,N_389);
or U1968 (N_1968,N_616,N_778);
nand U1969 (N_1969,N_477,N_553);
nor U1970 (N_1970,N_2,N_85);
nor U1971 (N_1971,N_142,N_552);
nor U1972 (N_1972,N_513,N_655);
nand U1973 (N_1973,N_4,N_262);
nor U1974 (N_1974,N_864,N_899);
and U1975 (N_1975,N_627,N_713);
and U1976 (N_1976,N_196,N_949);
nand U1977 (N_1977,N_451,N_249);
or U1978 (N_1978,N_318,N_143);
nand U1979 (N_1979,N_173,N_54);
or U1980 (N_1980,N_227,N_145);
xnor U1981 (N_1981,N_910,N_322);
nand U1982 (N_1982,N_641,N_866);
and U1983 (N_1983,N_798,N_134);
and U1984 (N_1984,N_972,N_503);
nor U1985 (N_1985,N_534,N_674);
and U1986 (N_1986,N_275,N_775);
or U1987 (N_1987,N_200,N_364);
nor U1988 (N_1988,N_391,N_750);
nor U1989 (N_1989,N_362,N_250);
nand U1990 (N_1990,N_621,N_407);
nand U1991 (N_1991,N_386,N_197);
or U1992 (N_1992,N_274,N_683);
nor U1993 (N_1993,N_269,N_981);
nand U1994 (N_1994,N_383,N_736);
or U1995 (N_1995,N_268,N_812);
and U1996 (N_1996,N_307,N_13);
nor U1997 (N_1997,N_119,N_162);
or U1998 (N_1998,N_898,N_123);
nand U1999 (N_1999,N_687,N_389);
or U2000 (N_2000,N_1986,N_1588);
nand U2001 (N_2001,N_1943,N_1562);
and U2002 (N_2002,N_1001,N_1063);
nand U2003 (N_2003,N_1507,N_1208);
or U2004 (N_2004,N_1372,N_1849);
and U2005 (N_2005,N_1904,N_1133);
or U2006 (N_2006,N_1613,N_1534);
nor U2007 (N_2007,N_1308,N_1352);
and U2008 (N_2008,N_1920,N_1688);
and U2009 (N_2009,N_1483,N_1855);
nor U2010 (N_2010,N_1791,N_1443);
and U2011 (N_2011,N_1994,N_1912);
nand U2012 (N_2012,N_1865,N_1579);
and U2013 (N_2013,N_1632,N_1415);
and U2014 (N_2014,N_1827,N_1875);
or U2015 (N_2015,N_1664,N_1864);
nor U2016 (N_2016,N_1332,N_1874);
or U2017 (N_2017,N_1614,N_1626);
nand U2018 (N_2018,N_1342,N_1597);
and U2019 (N_2019,N_1709,N_1438);
nand U2020 (N_2020,N_1427,N_1319);
and U2021 (N_2021,N_1363,N_1704);
or U2022 (N_2022,N_1120,N_1168);
or U2023 (N_2023,N_1173,N_1093);
nand U2024 (N_2024,N_1247,N_1464);
nor U2025 (N_2025,N_1650,N_1333);
or U2026 (N_2026,N_1795,N_1387);
or U2027 (N_2027,N_1863,N_1091);
or U2028 (N_2028,N_1019,N_1422);
or U2029 (N_2029,N_1498,N_1869);
or U2030 (N_2030,N_1105,N_1288);
or U2031 (N_2031,N_1757,N_1343);
or U2032 (N_2032,N_1354,N_1011);
or U2033 (N_2033,N_1031,N_1548);
nor U2034 (N_2034,N_1639,N_1222);
or U2035 (N_2035,N_1634,N_1574);
nand U2036 (N_2036,N_1264,N_1382);
and U2037 (N_2037,N_1385,N_1151);
and U2038 (N_2038,N_1403,N_1881);
nand U2039 (N_2039,N_1494,N_1629);
and U2040 (N_2040,N_1199,N_1822);
or U2041 (N_2041,N_1648,N_1367);
or U2042 (N_2042,N_1457,N_1254);
or U2043 (N_2043,N_1416,N_1197);
nand U2044 (N_2044,N_1395,N_1733);
nand U2045 (N_2045,N_1122,N_1779);
nand U2046 (N_2046,N_1041,N_1542);
nor U2047 (N_2047,N_1998,N_1182);
nand U2048 (N_2048,N_1274,N_1771);
nor U2049 (N_2049,N_1490,N_1453);
nor U2050 (N_2050,N_1877,N_1889);
nand U2051 (N_2051,N_1447,N_1318);
and U2052 (N_2052,N_1742,N_1831);
nor U2053 (N_2053,N_1720,N_1564);
nor U2054 (N_2054,N_1880,N_1040);
and U2055 (N_2055,N_1708,N_1723);
nor U2056 (N_2056,N_1409,N_1240);
nand U2057 (N_2057,N_1551,N_1493);
nor U2058 (N_2058,N_1200,N_1108);
and U2059 (N_2059,N_1316,N_1546);
nand U2060 (N_2060,N_1687,N_1901);
or U2061 (N_2061,N_1056,N_1995);
nand U2062 (N_2062,N_1171,N_1336);
nor U2063 (N_2063,N_1769,N_1295);
and U2064 (N_2064,N_1472,N_1426);
and U2065 (N_2065,N_1839,N_1030);
nor U2066 (N_2066,N_1203,N_1965);
nand U2067 (N_2067,N_1149,N_1898);
nor U2068 (N_2068,N_1775,N_1469);
nor U2069 (N_2069,N_1711,N_1068);
and U2070 (N_2070,N_1530,N_1259);
nor U2071 (N_2071,N_1911,N_1045);
nor U2072 (N_2072,N_1279,N_1265);
nor U2073 (N_2073,N_1862,N_1619);
and U2074 (N_2074,N_1136,N_1408);
or U2075 (N_2075,N_1992,N_1519);
or U2076 (N_2076,N_1402,N_1028);
and U2077 (N_2077,N_1275,N_1824);
or U2078 (N_2078,N_1516,N_1923);
nor U2079 (N_2079,N_1698,N_1523);
xnor U2080 (N_2080,N_1356,N_1162);
nor U2081 (N_2081,N_1599,N_1303);
nand U2082 (N_2082,N_1902,N_1896);
nand U2083 (N_2083,N_1370,N_1014);
nor U2084 (N_2084,N_1592,N_1398);
and U2085 (N_2085,N_1432,N_1962);
or U2086 (N_2086,N_1907,N_1241);
and U2087 (N_2087,N_1248,N_1331);
or U2088 (N_2088,N_1966,N_1861);
and U2089 (N_2089,N_1581,N_1334);
and U2090 (N_2090,N_1643,N_1048);
or U2091 (N_2091,N_1079,N_1100);
and U2092 (N_2092,N_1677,N_1654);
nor U2093 (N_2093,N_1411,N_1990);
or U2094 (N_2094,N_1537,N_1955);
or U2095 (N_2095,N_1550,N_1859);
nor U2096 (N_2096,N_1139,N_1852);
or U2097 (N_2097,N_1716,N_1140);
nor U2098 (N_2098,N_1231,N_1695);
nand U2099 (N_2099,N_1391,N_1702);
and U2100 (N_2100,N_1773,N_1157);
or U2101 (N_2101,N_1021,N_1183);
nand U2102 (N_2102,N_1871,N_1662);
nand U2103 (N_2103,N_1484,N_1908);
nand U2104 (N_2104,N_1125,N_1009);
and U2105 (N_2105,N_1557,N_1997);
or U2106 (N_2106,N_1207,N_1917);
nor U2107 (N_2107,N_1718,N_1536);
nand U2108 (N_2108,N_1987,N_1508);
or U2109 (N_2109,N_1217,N_1324);
nand U2110 (N_2110,N_1413,N_1095);
and U2111 (N_2111,N_1057,N_1892);
and U2112 (N_2112,N_1476,N_1958);
or U2113 (N_2113,N_1186,N_1355);
and U2114 (N_2114,N_1518,N_1475);
and U2115 (N_2115,N_1833,N_1710);
nor U2116 (N_2116,N_1243,N_1299);
or U2117 (N_2117,N_1442,N_1660);
and U2118 (N_2118,N_1107,N_1142);
and U2119 (N_2119,N_1276,N_1287);
and U2120 (N_2120,N_1237,N_1364);
and U2121 (N_2121,N_1081,N_1608);
xnor U2122 (N_2122,N_1641,N_1749);
and U2123 (N_2123,N_1073,N_1346);
nand U2124 (N_2124,N_1857,N_1329);
nor U2125 (N_2125,N_1780,N_1492);
or U2126 (N_2126,N_1089,N_1510);
and U2127 (N_2127,N_1585,N_1435);
and U2128 (N_2128,N_1478,N_1460);
nand U2129 (N_2129,N_1134,N_1979);
and U2130 (N_2130,N_1307,N_1218);
or U2131 (N_2131,N_1956,N_1948);
nor U2132 (N_2132,N_1394,N_1129);
xnor U2133 (N_2133,N_1777,N_1281);
nand U2134 (N_2134,N_1529,N_1651);
nand U2135 (N_2135,N_1971,N_1233);
nand U2136 (N_2136,N_1357,N_1396);
nor U2137 (N_2137,N_1817,N_1646);
or U2138 (N_2138,N_1512,N_1383);
and U2139 (N_2139,N_1211,N_1052);
nand U2140 (N_2140,N_1148,N_1730);
nand U2141 (N_2141,N_1844,N_1375);
and U2142 (N_2142,N_1503,N_1114);
xnor U2143 (N_2143,N_1999,N_1910);
and U2144 (N_2144,N_1843,N_1188);
and U2145 (N_2145,N_1527,N_1541);
and U2146 (N_2146,N_1658,N_1797);
or U2147 (N_2147,N_1804,N_1419);
and U2148 (N_2148,N_1158,N_1528);
or U2149 (N_2149,N_1604,N_1689);
or U2150 (N_2150,N_1553,N_1027);
nor U2151 (N_2151,N_1595,N_1765);
and U2152 (N_2152,N_1128,N_1339);
or U2153 (N_2153,N_1668,N_1781);
and U2154 (N_2154,N_1373,N_1576);
nand U2155 (N_2155,N_1325,N_1894);
and U2156 (N_2156,N_1437,N_1786);
or U2157 (N_2157,N_1851,N_1468);
and U2158 (N_2158,N_1180,N_1906);
nand U2159 (N_2159,N_1913,N_1025);
or U2160 (N_2160,N_1818,N_1347);
nand U2161 (N_2161,N_1082,N_1473);
or U2162 (N_2162,N_1885,N_1868);
or U2163 (N_2163,N_1296,N_1722);
nand U2164 (N_2164,N_1944,N_1927);
or U2165 (N_2165,N_1676,N_1117);
or U2166 (N_2166,N_1834,N_1763);
nand U2167 (N_2167,N_1344,N_1263);
nor U2168 (N_2168,N_1219,N_1666);
nand U2169 (N_2169,N_1671,N_1480);
nand U2170 (N_2170,N_1060,N_1617);
or U2171 (N_2171,N_1399,N_1178);
nor U2172 (N_2172,N_1793,N_1456);
or U2173 (N_2173,N_1450,N_1338);
or U2174 (N_2174,N_1882,N_1116);
nand U2175 (N_2175,N_1828,N_1072);
and U2176 (N_2176,N_1055,N_1008);
nor U2177 (N_2177,N_1462,N_1854);
or U2178 (N_2178,N_1729,N_1177);
nand U2179 (N_2179,N_1627,N_1230);
nand U2180 (N_2180,N_1803,N_1522);
and U2181 (N_2181,N_1262,N_1061);
or U2182 (N_2182,N_1739,N_1431);
and U2183 (N_2183,N_1034,N_1505);
nand U2184 (N_2184,N_1813,N_1270);
nand U2185 (N_2185,N_1015,N_1572);
nor U2186 (N_2186,N_1830,N_1097);
nand U2187 (N_2187,N_1502,N_1423);
nand U2188 (N_2188,N_1558,N_1821);
or U2189 (N_2189,N_1705,N_1315);
nand U2190 (N_2190,N_1993,N_1606);
and U2191 (N_2191,N_1421,N_1937);
or U2192 (N_2192,N_1414,N_1637);
nand U2193 (N_2193,N_1837,N_1206);
nor U2194 (N_2194,N_1916,N_1560);
and U2195 (N_2195,N_1286,N_1446);
and U2196 (N_2196,N_1044,N_1888);
and U2197 (N_2197,N_1486,N_1135);
or U2198 (N_2198,N_1376,N_1064);
nand U2199 (N_2199,N_1582,N_1531);
nor U2200 (N_2200,N_1022,N_1360);
nor U2201 (N_2201,N_1080,N_1578);
or U2202 (N_2202,N_1684,N_1312);
or U2203 (N_2203,N_1846,N_1016);
nand U2204 (N_2204,N_1938,N_1043);
nor U2205 (N_2205,N_1776,N_1841);
nand U2206 (N_2206,N_1945,N_1147);
or U2207 (N_2207,N_1330,N_1591);
nand U2208 (N_2208,N_1113,N_1098);
nand U2209 (N_2209,N_1046,N_1732);
or U2210 (N_2210,N_1561,N_1485);
and U2211 (N_2211,N_1320,N_1566);
nor U2212 (N_2212,N_1584,N_1215);
nor U2213 (N_2213,N_1974,N_1002);
nand U2214 (N_2214,N_1118,N_1767);
nor U2215 (N_2215,N_1682,N_1198);
or U2216 (N_2216,N_1221,N_1154);
nand U2217 (N_2217,N_1701,N_1670);
or U2218 (N_2218,N_1418,N_1146);
and U2219 (N_2219,N_1176,N_1615);
and U2220 (N_2220,N_1895,N_1351);
and U2221 (N_2221,N_1448,N_1466);
nand U2222 (N_2222,N_1850,N_1463);
and U2223 (N_2223,N_1870,N_1878);
nor U2224 (N_2224,N_1526,N_1305);
nor U2225 (N_2225,N_1227,N_1808);
nand U2226 (N_2226,N_1939,N_1205);
nor U2227 (N_2227,N_1083,N_1238);
nor U2228 (N_2228,N_1616,N_1514);
nor U2229 (N_2229,N_1903,N_1700);
nor U2230 (N_2230,N_1369,N_1618);
nor U2231 (N_2231,N_1397,N_1761);
or U2232 (N_2232,N_1007,N_1005);
nand U2233 (N_2233,N_1829,N_1890);
or U2234 (N_2234,N_1388,N_1989);
or U2235 (N_2235,N_1038,N_1380);
nand U2236 (N_2236,N_1362,N_1268);
nand U2237 (N_2237,N_1488,N_1544);
nor U2238 (N_2238,N_1524,N_1814);
or U2239 (N_2239,N_1066,N_1681);
nor U2240 (N_2240,N_1065,N_1153);
nand U2241 (N_2241,N_1379,N_1212);
and U2242 (N_2242,N_1745,N_1800);
nand U2243 (N_2243,N_1326,N_1214);
and U2244 (N_2244,N_1954,N_1792);
and U2245 (N_2245,N_1253,N_1980);
and U2246 (N_2246,N_1897,N_1036);
nand U2247 (N_2247,N_1915,N_1412);
nor U2248 (N_2248,N_1246,N_1690);
or U2249 (N_2249,N_1328,N_1420);
nand U2250 (N_2250,N_1549,N_1109);
and U2251 (N_2251,N_1131,N_1925);
nand U2252 (N_2252,N_1663,N_1235);
or U2253 (N_2253,N_1481,N_1587);
xnor U2254 (N_2254,N_1784,N_1598);
nand U2255 (N_2255,N_1714,N_1406);
nor U2256 (N_2256,N_1694,N_1764);
and U2257 (N_2257,N_1630,N_1145);
and U2258 (N_2258,N_1170,N_1759);
nor U2259 (N_2259,N_1282,N_1758);
nor U2260 (N_2260,N_1174,N_1216);
nand U2261 (N_2261,N_1750,N_1094);
or U2262 (N_2262,N_1244,N_1589);
nor U2263 (N_2263,N_1126,N_1285);
and U2264 (N_2264,N_1751,N_1899);
and U2265 (N_2265,N_1744,N_1278);
or U2266 (N_2266,N_1461,N_1725);
nand U2267 (N_2267,N_1922,N_1790);
and U2268 (N_2268,N_1085,N_1189);
nor U2269 (N_2269,N_1020,N_1436);
and U2270 (N_2270,N_1185,N_1289);
nor U2271 (N_2271,N_1787,N_1161);
or U2272 (N_2272,N_1590,N_1389);
or U2273 (N_2273,N_1166,N_1191);
and U2274 (N_2274,N_1042,N_1930);
and U2275 (N_2275,N_1873,N_1187);
and U2276 (N_2276,N_1283,N_1740);
or U2277 (N_2277,N_1856,N_1292);
and U2278 (N_2278,N_1770,N_1565);
and U2279 (N_2279,N_1968,N_1430);
nor U2280 (N_2280,N_1074,N_1736);
nand U2281 (N_2281,N_1201,N_1569);
nor U2282 (N_2282,N_1543,N_1459);
nand U2283 (N_2283,N_1547,N_1410);
or U2284 (N_2284,N_1812,N_1699);
or U2285 (N_2285,N_1636,N_1953);
nand U2286 (N_2286,N_1455,N_1961);
and U2287 (N_2287,N_1096,N_1424);
nand U2288 (N_2288,N_1600,N_1631);
or U2289 (N_2289,N_1479,N_1605);
and U2290 (N_2290,N_1719,N_1353);
nor U2291 (N_2291,N_1257,N_1006);
and U2292 (N_2292,N_1612,N_1921);
or U2293 (N_2293,N_1900,N_1224);
nand U2294 (N_2294,N_1284,N_1314);
or U2295 (N_2295,N_1973,N_1876);
nand U2296 (N_2296,N_1032,N_1638);
nand U2297 (N_2297,N_1748,N_1054);
or U2298 (N_2298,N_1559,N_1349);
xnor U2299 (N_2299,N_1358,N_1746);
and U2300 (N_2300,N_1620,N_1807);
nor U2301 (N_2301,N_1384,N_1076);
nand U2302 (N_2302,N_1940,N_1290);
and U2303 (N_2303,N_1607,N_1236);
or U2304 (N_2304,N_1712,N_1350);
or U2305 (N_2305,N_1445,N_1267);
or U2306 (N_2306,N_1070,N_1838);
nor U2307 (N_2307,N_1103,N_1220);
nor U2308 (N_2308,N_1778,N_1556);
and U2309 (N_2309,N_1169,N_1836);
nand U2310 (N_2310,N_1024,N_1306);
nor U2311 (N_2311,N_1728,N_1652);
xnor U2312 (N_2312,N_1743,N_1121);
or U2313 (N_2313,N_1371,N_1381);
or U2314 (N_2314,N_1321,N_1947);
nor U2315 (N_2315,N_1449,N_1842);
or U2316 (N_2316,N_1084,N_1210);
nand U2317 (N_2317,N_1573,N_1322);
or U2318 (N_2318,N_1884,N_1672);
nand U2319 (N_2319,N_1348,N_1075);
nor U2320 (N_2320,N_1327,N_1539);
nor U2321 (N_2321,N_1951,N_1984);
nand U2322 (N_2322,N_1825,N_1713);
nand U2323 (N_2323,N_1949,N_1458);
or U2324 (N_2324,N_1752,N_1345);
or U2325 (N_2325,N_1101,N_1640);
and U2326 (N_2326,N_1088,N_1794);
and U2327 (N_2327,N_1934,N_1840);
or U2328 (N_2328,N_1872,N_1832);
or U2329 (N_2329,N_1209,N_1192);
nor U2330 (N_2330,N_1071,N_1035);
nand U2331 (N_2331,N_1686,N_1960);
and U2332 (N_2332,N_1946,N_1806);
and U2333 (N_2333,N_1820,N_1610);
and U2334 (N_2334,N_1933,N_1496);
and U2335 (N_2335,N_1138,N_1175);
nor U2336 (N_2336,N_1935,N_1970);
nor U2337 (N_2337,N_1050,N_1981);
and U2338 (N_2338,N_1132,N_1853);
nor U2339 (N_2339,N_1417,N_1633);
nor U2340 (N_2340,N_1390,N_1179);
nand U2341 (N_2341,N_1517,N_1404);
nor U2342 (N_2342,N_1622,N_1540);
or U2343 (N_2343,N_1644,N_1297);
and U2344 (N_2344,N_1674,N_1317);
and U2345 (N_2345,N_1195,N_1809);
or U2346 (N_2346,N_1232,N_1805);
or U2347 (N_2347,N_1500,N_1159);
nor U2348 (N_2348,N_1996,N_1796);
nand U2349 (N_2349,N_1801,N_1256);
or U2350 (N_2350,N_1515,N_1069);
nor U2351 (N_2351,N_1571,N_1225);
or U2352 (N_2352,N_1474,N_1340);
or U2353 (N_2353,N_1033,N_1647);
and U2354 (N_2354,N_1623,N_1665);
nor U2355 (N_2355,N_1172,N_1621);
and U2356 (N_2356,N_1789,N_1680);
nor U2357 (N_2357,N_1501,N_1545);
nand U2358 (N_2358,N_1451,N_1452);
xor U2359 (N_2359,N_1957,N_1150);
and U2360 (N_2360,N_1444,N_1428);
nor U2361 (N_2361,N_1625,N_1819);
and U2362 (N_2362,N_1657,N_1762);
nand U2363 (N_2363,N_1706,N_1504);
nand U2364 (N_2364,N_1051,N_1988);
and U2365 (N_2365,N_1931,N_1703);
and U2366 (N_2366,N_1491,N_1609);
and U2367 (N_2367,N_1577,N_1249);
and U2368 (N_2368,N_1715,N_1659);
or U2369 (N_2369,N_1642,N_1405);
or U2370 (N_2370,N_1985,N_1099);
nor U2371 (N_2371,N_1747,N_1766);
nor U2372 (N_2372,N_1799,N_1977);
or U2373 (N_2373,N_1835,N_1104);
and U2374 (N_2374,N_1772,N_1774);
or U2375 (N_2375,N_1982,N_1513);
nand U2376 (N_2376,N_1506,N_1090);
or U2377 (N_2377,N_1628,N_1509);
nor U2378 (N_2378,N_1738,N_1086);
or U2379 (N_2379,N_1735,N_1969);
and U2380 (N_2380,N_1310,N_1039);
nand U2381 (N_2381,N_1123,N_1141);
nor U2382 (N_2382,N_1683,N_1811);
and U2383 (N_2383,N_1078,N_1783);
and U2384 (N_2384,N_1959,N_1401);
or U2385 (N_2385,N_1092,N_1026);
nor U2386 (N_2386,N_1049,N_1361);
nor U2387 (N_2387,N_1721,N_1497);
or U2388 (N_2388,N_1731,N_1229);
and U2389 (N_2389,N_1127,N_1798);
nand U2390 (N_2390,N_1929,N_1313);
or U2391 (N_2391,N_1685,N_1656);
nor U2392 (N_2392,N_1645,N_1887);
or U2393 (N_2393,N_1300,N_1675);
nand U2394 (N_2394,N_1741,N_1053);
and U2395 (N_2395,N_1905,N_1234);
nor U2396 (N_2396,N_1782,N_1879);
and U2397 (N_2397,N_1860,N_1261);
nand U2398 (N_2398,N_1193,N_1359);
and U2399 (N_2399,N_1983,N_1568);
nor U2400 (N_2400,N_1909,N_1555);
nor U2401 (N_2401,N_1823,N_1487);
or U2402 (N_2402,N_1304,N_1593);
and U2403 (N_2403,N_1155,N_1810);
or U2404 (N_2404,N_1273,N_1693);
or U2405 (N_2405,N_1272,N_1277);
or U2406 (N_2406,N_1112,N_1223);
and U2407 (N_2407,N_1309,N_1583);
nand U2408 (N_2408,N_1047,N_1724);
or U2409 (N_2409,N_1816,N_1124);
or U2410 (N_2410,N_1298,N_1950);
and U2411 (N_2411,N_1554,N_1470);
and U2412 (N_2412,N_1611,N_1691);
or U2413 (N_2413,N_1269,N_1137);
xnor U2414 (N_2414,N_1365,N_1378);
nor U2415 (N_2415,N_1533,N_1737);
and U2416 (N_2416,N_1848,N_1266);
nand U2417 (N_2417,N_1110,N_1111);
xor U2418 (N_2418,N_1707,N_1717);
nand U2419 (N_2419,N_1067,N_1521);
nand U2420 (N_2420,N_1335,N_1003);
nor U2421 (N_2421,N_1760,N_1919);
or U2422 (N_2422,N_1570,N_1144);
nor U2423 (N_2423,N_1004,N_1013);
nor U2424 (N_2424,N_1926,N_1425);
nor U2425 (N_2425,N_1826,N_1802);
or U2426 (N_2426,N_1156,N_1433);
and U2427 (N_2427,N_1883,N_1673);
and U2428 (N_2428,N_1018,N_1858);
and U2429 (N_2429,N_1062,N_1037);
nand U2430 (N_2430,N_1678,N_1184);
nor U2431 (N_2431,N_1785,N_1552);
or U2432 (N_2432,N_1251,N_1441);
nor U2433 (N_2433,N_1252,N_1190);
and U2434 (N_2434,N_1495,N_1963);
or U2435 (N_2435,N_1392,N_1194);
nor U2436 (N_2436,N_1454,N_1258);
nor U2437 (N_2437,N_1538,N_1368);
nor U2438 (N_2438,N_1181,N_1087);
nor U2439 (N_2439,N_1239,N_1115);
nand U2440 (N_2440,N_1978,N_1753);
and U2441 (N_2441,N_1815,N_1012);
and U2442 (N_2442,N_1482,N_1160);
or U2443 (N_2443,N_1059,N_1649);
and U2444 (N_2444,N_1429,N_1291);
or U2445 (N_2445,N_1499,N_1102);
nor U2446 (N_2446,N_1596,N_1374);
and U2447 (N_2447,N_1972,N_1580);
or U2448 (N_2448,N_1563,N_1280);
and U2449 (N_2449,N_1029,N_1866);
and U2450 (N_2450,N_1669,N_1726);
and U2451 (N_2451,N_1928,N_1655);
nor U2452 (N_2452,N_1077,N_1377);
or U2453 (N_2453,N_1471,N_1967);
or U2454 (N_2454,N_1696,N_1106);
or U2455 (N_2455,N_1727,N_1601);
nand U2456 (N_2456,N_1964,N_1603);
nand U2457 (N_2457,N_1535,N_1010);
nand U2458 (N_2458,N_1271,N_1692);
and U2459 (N_2459,N_1337,N_1952);
and U2460 (N_2460,N_1886,N_1366);
and U2461 (N_2461,N_1932,N_1301);
nand U2462 (N_2462,N_1341,N_1386);
or U2463 (N_2463,N_1661,N_1697);
nor U2464 (N_2464,N_1393,N_1255);
nor U2465 (N_2465,N_1893,N_1196);
and U2466 (N_2466,N_1250,N_1294);
and U2467 (N_2467,N_1130,N_1311);
and U2468 (N_2468,N_1755,N_1204);
xor U2469 (N_2469,N_1143,N_1768);
or U2470 (N_2470,N_1164,N_1594);
or U2471 (N_2471,N_1602,N_1293);
nor U2472 (N_2472,N_1942,N_1400);
or U2473 (N_2473,N_1754,N_1936);
and U2474 (N_2474,N_1023,N_1058);
nor U2475 (N_2475,N_1918,N_1467);
nand U2476 (N_2476,N_1653,N_1323);
or U2477 (N_2477,N_1788,N_1152);
nor U2478 (N_2478,N_1465,N_1017);
or U2479 (N_2479,N_1213,N_1202);
and U2480 (N_2480,N_1407,N_1260);
nor U2481 (N_2481,N_1489,N_1439);
or U2482 (N_2482,N_1756,N_1242);
nor U2483 (N_2483,N_1167,N_1586);
and U2484 (N_2484,N_1867,N_1532);
or U2485 (N_2485,N_1976,N_1163);
nor U2486 (N_2486,N_1525,N_1575);
and U2487 (N_2487,N_1511,N_1477);
nor U2488 (N_2488,N_1520,N_1226);
nand U2489 (N_2489,N_1119,N_1302);
nand U2490 (N_2490,N_1667,N_1679);
and U2491 (N_2491,N_1000,N_1165);
nand U2492 (N_2492,N_1434,N_1845);
nor U2493 (N_2493,N_1975,N_1624);
or U2494 (N_2494,N_1228,N_1941);
or U2495 (N_2495,N_1635,N_1245);
and U2496 (N_2496,N_1440,N_1567);
and U2497 (N_2497,N_1991,N_1924);
and U2498 (N_2498,N_1734,N_1891);
and U2499 (N_2499,N_1914,N_1847);
nor U2500 (N_2500,N_1279,N_1517);
and U2501 (N_2501,N_1265,N_1360);
or U2502 (N_2502,N_1940,N_1395);
nand U2503 (N_2503,N_1863,N_1274);
nor U2504 (N_2504,N_1083,N_1585);
nand U2505 (N_2505,N_1074,N_1601);
nand U2506 (N_2506,N_1143,N_1886);
nor U2507 (N_2507,N_1385,N_1350);
or U2508 (N_2508,N_1317,N_1514);
or U2509 (N_2509,N_1395,N_1530);
xor U2510 (N_2510,N_1779,N_1552);
nor U2511 (N_2511,N_1003,N_1062);
nor U2512 (N_2512,N_1760,N_1841);
or U2513 (N_2513,N_1489,N_1125);
or U2514 (N_2514,N_1232,N_1081);
nand U2515 (N_2515,N_1115,N_1728);
nor U2516 (N_2516,N_1809,N_1554);
nand U2517 (N_2517,N_1194,N_1891);
nand U2518 (N_2518,N_1328,N_1695);
xnor U2519 (N_2519,N_1158,N_1060);
nand U2520 (N_2520,N_1809,N_1650);
or U2521 (N_2521,N_1549,N_1741);
and U2522 (N_2522,N_1886,N_1000);
or U2523 (N_2523,N_1341,N_1626);
and U2524 (N_2524,N_1805,N_1733);
nand U2525 (N_2525,N_1413,N_1724);
nor U2526 (N_2526,N_1001,N_1513);
nor U2527 (N_2527,N_1845,N_1294);
and U2528 (N_2528,N_1734,N_1224);
nor U2529 (N_2529,N_1520,N_1538);
or U2530 (N_2530,N_1723,N_1063);
or U2531 (N_2531,N_1735,N_1504);
nor U2532 (N_2532,N_1671,N_1069);
nand U2533 (N_2533,N_1637,N_1116);
or U2534 (N_2534,N_1846,N_1778);
nand U2535 (N_2535,N_1035,N_1960);
or U2536 (N_2536,N_1050,N_1118);
or U2537 (N_2537,N_1104,N_1977);
nand U2538 (N_2538,N_1881,N_1713);
nand U2539 (N_2539,N_1218,N_1254);
and U2540 (N_2540,N_1002,N_1493);
nand U2541 (N_2541,N_1077,N_1700);
and U2542 (N_2542,N_1363,N_1003);
nor U2543 (N_2543,N_1354,N_1846);
or U2544 (N_2544,N_1785,N_1902);
nand U2545 (N_2545,N_1508,N_1432);
nand U2546 (N_2546,N_1903,N_1312);
and U2547 (N_2547,N_1758,N_1138);
nand U2548 (N_2548,N_1076,N_1085);
nand U2549 (N_2549,N_1706,N_1982);
nand U2550 (N_2550,N_1761,N_1224);
and U2551 (N_2551,N_1077,N_1932);
or U2552 (N_2552,N_1382,N_1553);
and U2553 (N_2553,N_1528,N_1492);
nand U2554 (N_2554,N_1989,N_1571);
and U2555 (N_2555,N_1983,N_1870);
xor U2556 (N_2556,N_1758,N_1650);
nor U2557 (N_2557,N_1597,N_1381);
nand U2558 (N_2558,N_1168,N_1386);
or U2559 (N_2559,N_1946,N_1966);
nor U2560 (N_2560,N_1949,N_1707);
and U2561 (N_2561,N_1656,N_1217);
or U2562 (N_2562,N_1837,N_1864);
nand U2563 (N_2563,N_1900,N_1523);
or U2564 (N_2564,N_1986,N_1584);
nand U2565 (N_2565,N_1223,N_1012);
nand U2566 (N_2566,N_1617,N_1226);
nor U2567 (N_2567,N_1409,N_1590);
and U2568 (N_2568,N_1044,N_1251);
or U2569 (N_2569,N_1855,N_1937);
nor U2570 (N_2570,N_1440,N_1134);
nand U2571 (N_2571,N_1978,N_1494);
or U2572 (N_2572,N_1559,N_1199);
and U2573 (N_2573,N_1598,N_1730);
and U2574 (N_2574,N_1889,N_1680);
and U2575 (N_2575,N_1400,N_1527);
or U2576 (N_2576,N_1988,N_1671);
nand U2577 (N_2577,N_1139,N_1372);
nor U2578 (N_2578,N_1127,N_1873);
and U2579 (N_2579,N_1399,N_1580);
nor U2580 (N_2580,N_1292,N_1551);
nand U2581 (N_2581,N_1653,N_1881);
or U2582 (N_2582,N_1121,N_1017);
nand U2583 (N_2583,N_1927,N_1347);
and U2584 (N_2584,N_1924,N_1870);
xnor U2585 (N_2585,N_1695,N_1451);
or U2586 (N_2586,N_1222,N_1598);
nor U2587 (N_2587,N_1186,N_1734);
nor U2588 (N_2588,N_1786,N_1563);
or U2589 (N_2589,N_1630,N_1097);
and U2590 (N_2590,N_1952,N_1598);
and U2591 (N_2591,N_1615,N_1581);
and U2592 (N_2592,N_1147,N_1289);
nand U2593 (N_2593,N_1743,N_1701);
and U2594 (N_2594,N_1800,N_1644);
and U2595 (N_2595,N_1436,N_1800);
and U2596 (N_2596,N_1550,N_1535);
xor U2597 (N_2597,N_1676,N_1819);
nor U2598 (N_2598,N_1240,N_1681);
and U2599 (N_2599,N_1779,N_1200);
nand U2600 (N_2600,N_1432,N_1976);
and U2601 (N_2601,N_1726,N_1487);
or U2602 (N_2602,N_1414,N_1532);
nand U2603 (N_2603,N_1066,N_1780);
nor U2604 (N_2604,N_1100,N_1483);
or U2605 (N_2605,N_1798,N_1781);
or U2606 (N_2606,N_1402,N_1958);
nor U2607 (N_2607,N_1112,N_1049);
and U2608 (N_2608,N_1993,N_1359);
nor U2609 (N_2609,N_1099,N_1605);
nor U2610 (N_2610,N_1212,N_1055);
nand U2611 (N_2611,N_1538,N_1880);
or U2612 (N_2612,N_1555,N_1375);
or U2613 (N_2613,N_1291,N_1668);
and U2614 (N_2614,N_1096,N_1848);
nor U2615 (N_2615,N_1537,N_1820);
nor U2616 (N_2616,N_1370,N_1063);
and U2617 (N_2617,N_1691,N_1081);
and U2618 (N_2618,N_1957,N_1631);
nand U2619 (N_2619,N_1406,N_1340);
nand U2620 (N_2620,N_1509,N_1958);
nand U2621 (N_2621,N_1300,N_1445);
nand U2622 (N_2622,N_1817,N_1909);
nor U2623 (N_2623,N_1473,N_1938);
nand U2624 (N_2624,N_1528,N_1938);
nand U2625 (N_2625,N_1818,N_1664);
and U2626 (N_2626,N_1566,N_1451);
nor U2627 (N_2627,N_1470,N_1764);
and U2628 (N_2628,N_1563,N_1074);
or U2629 (N_2629,N_1737,N_1049);
nand U2630 (N_2630,N_1223,N_1162);
nand U2631 (N_2631,N_1081,N_1252);
nor U2632 (N_2632,N_1203,N_1888);
xor U2633 (N_2633,N_1792,N_1315);
nor U2634 (N_2634,N_1694,N_1677);
nand U2635 (N_2635,N_1078,N_1909);
or U2636 (N_2636,N_1250,N_1203);
nor U2637 (N_2637,N_1421,N_1983);
and U2638 (N_2638,N_1057,N_1472);
nor U2639 (N_2639,N_1166,N_1726);
and U2640 (N_2640,N_1913,N_1972);
and U2641 (N_2641,N_1378,N_1507);
nand U2642 (N_2642,N_1434,N_1360);
nand U2643 (N_2643,N_1370,N_1906);
nand U2644 (N_2644,N_1294,N_1173);
or U2645 (N_2645,N_1147,N_1813);
nor U2646 (N_2646,N_1720,N_1935);
nand U2647 (N_2647,N_1499,N_1618);
or U2648 (N_2648,N_1941,N_1902);
and U2649 (N_2649,N_1048,N_1461);
nand U2650 (N_2650,N_1549,N_1949);
nor U2651 (N_2651,N_1937,N_1310);
or U2652 (N_2652,N_1210,N_1773);
or U2653 (N_2653,N_1374,N_1932);
or U2654 (N_2654,N_1066,N_1908);
or U2655 (N_2655,N_1872,N_1926);
and U2656 (N_2656,N_1514,N_1904);
nand U2657 (N_2657,N_1512,N_1286);
nor U2658 (N_2658,N_1341,N_1101);
nand U2659 (N_2659,N_1092,N_1605);
nor U2660 (N_2660,N_1395,N_1259);
nor U2661 (N_2661,N_1882,N_1816);
nor U2662 (N_2662,N_1677,N_1408);
or U2663 (N_2663,N_1977,N_1942);
and U2664 (N_2664,N_1431,N_1958);
and U2665 (N_2665,N_1751,N_1370);
nor U2666 (N_2666,N_1213,N_1304);
or U2667 (N_2667,N_1088,N_1816);
or U2668 (N_2668,N_1371,N_1958);
nand U2669 (N_2669,N_1268,N_1861);
nand U2670 (N_2670,N_1227,N_1634);
and U2671 (N_2671,N_1860,N_1191);
nand U2672 (N_2672,N_1179,N_1799);
nor U2673 (N_2673,N_1372,N_1802);
nor U2674 (N_2674,N_1572,N_1319);
nand U2675 (N_2675,N_1962,N_1128);
and U2676 (N_2676,N_1755,N_1885);
xor U2677 (N_2677,N_1410,N_1367);
nand U2678 (N_2678,N_1479,N_1091);
nor U2679 (N_2679,N_1693,N_1745);
nor U2680 (N_2680,N_1942,N_1859);
or U2681 (N_2681,N_1968,N_1516);
and U2682 (N_2682,N_1747,N_1791);
nand U2683 (N_2683,N_1469,N_1004);
nor U2684 (N_2684,N_1825,N_1542);
and U2685 (N_2685,N_1403,N_1178);
nand U2686 (N_2686,N_1621,N_1351);
nor U2687 (N_2687,N_1577,N_1098);
nand U2688 (N_2688,N_1171,N_1580);
and U2689 (N_2689,N_1526,N_1952);
nand U2690 (N_2690,N_1419,N_1563);
nor U2691 (N_2691,N_1480,N_1730);
nand U2692 (N_2692,N_1298,N_1207);
or U2693 (N_2693,N_1490,N_1424);
nand U2694 (N_2694,N_1278,N_1386);
or U2695 (N_2695,N_1928,N_1649);
or U2696 (N_2696,N_1196,N_1420);
nand U2697 (N_2697,N_1947,N_1551);
and U2698 (N_2698,N_1784,N_1188);
nand U2699 (N_2699,N_1583,N_1828);
nor U2700 (N_2700,N_1437,N_1900);
nor U2701 (N_2701,N_1552,N_1237);
and U2702 (N_2702,N_1587,N_1836);
or U2703 (N_2703,N_1164,N_1746);
nor U2704 (N_2704,N_1514,N_1984);
nand U2705 (N_2705,N_1520,N_1096);
or U2706 (N_2706,N_1747,N_1495);
xnor U2707 (N_2707,N_1163,N_1337);
or U2708 (N_2708,N_1083,N_1213);
nor U2709 (N_2709,N_1520,N_1193);
nor U2710 (N_2710,N_1706,N_1987);
and U2711 (N_2711,N_1536,N_1114);
and U2712 (N_2712,N_1987,N_1144);
nand U2713 (N_2713,N_1884,N_1239);
nor U2714 (N_2714,N_1138,N_1787);
nor U2715 (N_2715,N_1278,N_1799);
or U2716 (N_2716,N_1978,N_1327);
nand U2717 (N_2717,N_1839,N_1202);
nor U2718 (N_2718,N_1112,N_1106);
nor U2719 (N_2719,N_1483,N_1118);
and U2720 (N_2720,N_1454,N_1120);
and U2721 (N_2721,N_1578,N_1092);
nor U2722 (N_2722,N_1992,N_1295);
nand U2723 (N_2723,N_1602,N_1861);
or U2724 (N_2724,N_1044,N_1905);
and U2725 (N_2725,N_1776,N_1938);
nand U2726 (N_2726,N_1883,N_1429);
and U2727 (N_2727,N_1947,N_1699);
and U2728 (N_2728,N_1491,N_1380);
and U2729 (N_2729,N_1356,N_1794);
nor U2730 (N_2730,N_1529,N_1821);
or U2731 (N_2731,N_1821,N_1358);
and U2732 (N_2732,N_1239,N_1768);
or U2733 (N_2733,N_1640,N_1937);
and U2734 (N_2734,N_1613,N_1064);
and U2735 (N_2735,N_1623,N_1622);
nand U2736 (N_2736,N_1739,N_1906);
nand U2737 (N_2737,N_1324,N_1413);
nor U2738 (N_2738,N_1767,N_1380);
or U2739 (N_2739,N_1410,N_1920);
nor U2740 (N_2740,N_1087,N_1853);
nand U2741 (N_2741,N_1448,N_1147);
nor U2742 (N_2742,N_1909,N_1412);
nor U2743 (N_2743,N_1204,N_1641);
and U2744 (N_2744,N_1190,N_1069);
and U2745 (N_2745,N_1925,N_1732);
and U2746 (N_2746,N_1978,N_1207);
nor U2747 (N_2747,N_1907,N_1242);
and U2748 (N_2748,N_1661,N_1087);
or U2749 (N_2749,N_1746,N_1968);
or U2750 (N_2750,N_1301,N_1779);
nand U2751 (N_2751,N_1493,N_1460);
and U2752 (N_2752,N_1384,N_1498);
or U2753 (N_2753,N_1040,N_1227);
or U2754 (N_2754,N_1891,N_1100);
or U2755 (N_2755,N_1243,N_1460);
and U2756 (N_2756,N_1526,N_1268);
and U2757 (N_2757,N_1176,N_1070);
nor U2758 (N_2758,N_1946,N_1526);
nand U2759 (N_2759,N_1296,N_1857);
and U2760 (N_2760,N_1111,N_1465);
and U2761 (N_2761,N_1098,N_1084);
and U2762 (N_2762,N_1251,N_1045);
or U2763 (N_2763,N_1157,N_1028);
or U2764 (N_2764,N_1260,N_1072);
or U2765 (N_2765,N_1571,N_1912);
nor U2766 (N_2766,N_1334,N_1136);
and U2767 (N_2767,N_1595,N_1956);
nand U2768 (N_2768,N_1915,N_1391);
or U2769 (N_2769,N_1654,N_1386);
and U2770 (N_2770,N_1177,N_1642);
nand U2771 (N_2771,N_1063,N_1685);
nor U2772 (N_2772,N_1592,N_1401);
and U2773 (N_2773,N_1860,N_1414);
nor U2774 (N_2774,N_1957,N_1781);
and U2775 (N_2775,N_1542,N_1577);
or U2776 (N_2776,N_1785,N_1931);
or U2777 (N_2777,N_1809,N_1626);
and U2778 (N_2778,N_1066,N_1719);
nor U2779 (N_2779,N_1626,N_1328);
and U2780 (N_2780,N_1973,N_1535);
and U2781 (N_2781,N_1998,N_1691);
and U2782 (N_2782,N_1998,N_1027);
and U2783 (N_2783,N_1017,N_1727);
or U2784 (N_2784,N_1528,N_1249);
nand U2785 (N_2785,N_1881,N_1598);
and U2786 (N_2786,N_1265,N_1460);
or U2787 (N_2787,N_1025,N_1238);
nor U2788 (N_2788,N_1577,N_1672);
nand U2789 (N_2789,N_1174,N_1898);
and U2790 (N_2790,N_1373,N_1366);
nand U2791 (N_2791,N_1560,N_1190);
and U2792 (N_2792,N_1929,N_1540);
and U2793 (N_2793,N_1914,N_1325);
nand U2794 (N_2794,N_1986,N_1617);
or U2795 (N_2795,N_1162,N_1002);
or U2796 (N_2796,N_1264,N_1151);
nor U2797 (N_2797,N_1406,N_1136);
nor U2798 (N_2798,N_1202,N_1783);
or U2799 (N_2799,N_1583,N_1026);
and U2800 (N_2800,N_1728,N_1619);
nand U2801 (N_2801,N_1795,N_1223);
nor U2802 (N_2802,N_1034,N_1798);
nor U2803 (N_2803,N_1195,N_1555);
nor U2804 (N_2804,N_1036,N_1102);
nand U2805 (N_2805,N_1777,N_1019);
nor U2806 (N_2806,N_1238,N_1296);
and U2807 (N_2807,N_1244,N_1359);
nor U2808 (N_2808,N_1849,N_1126);
and U2809 (N_2809,N_1137,N_1458);
or U2810 (N_2810,N_1839,N_1947);
or U2811 (N_2811,N_1395,N_1362);
or U2812 (N_2812,N_1755,N_1212);
or U2813 (N_2813,N_1529,N_1783);
and U2814 (N_2814,N_1411,N_1270);
and U2815 (N_2815,N_1780,N_1650);
or U2816 (N_2816,N_1064,N_1107);
nand U2817 (N_2817,N_1664,N_1011);
nor U2818 (N_2818,N_1858,N_1921);
or U2819 (N_2819,N_1312,N_1304);
nor U2820 (N_2820,N_1126,N_1516);
nand U2821 (N_2821,N_1568,N_1219);
nor U2822 (N_2822,N_1450,N_1798);
and U2823 (N_2823,N_1632,N_1794);
and U2824 (N_2824,N_1995,N_1786);
or U2825 (N_2825,N_1559,N_1044);
nor U2826 (N_2826,N_1506,N_1593);
nand U2827 (N_2827,N_1133,N_1769);
or U2828 (N_2828,N_1329,N_1096);
nor U2829 (N_2829,N_1100,N_1395);
nand U2830 (N_2830,N_1851,N_1767);
nand U2831 (N_2831,N_1527,N_1473);
or U2832 (N_2832,N_1730,N_1669);
nor U2833 (N_2833,N_1112,N_1327);
nand U2834 (N_2834,N_1707,N_1612);
or U2835 (N_2835,N_1246,N_1617);
nand U2836 (N_2836,N_1650,N_1112);
and U2837 (N_2837,N_1145,N_1850);
nor U2838 (N_2838,N_1867,N_1808);
and U2839 (N_2839,N_1439,N_1414);
or U2840 (N_2840,N_1314,N_1461);
nor U2841 (N_2841,N_1998,N_1678);
and U2842 (N_2842,N_1724,N_1711);
or U2843 (N_2843,N_1875,N_1898);
nor U2844 (N_2844,N_1232,N_1873);
nand U2845 (N_2845,N_1458,N_1425);
or U2846 (N_2846,N_1692,N_1673);
nor U2847 (N_2847,N_1668,N_1213);
nor U2848 (N_2848,N_1052,N_1416);
and U2849 (N_2849,N_1980,N_1701);
nand U2850 (N_2850,N_1201,N_1097);
nor U2851 (N_2851,N_1695,N_1286);
and U2852 (N_2852,N_1191,N_1344);
and U2853 (N_2853,N_1807,N_1574);
or U2854 (N_2854,N_1151,N_1074);
or U2855 (N_2855,N_1054,N_1500);
and U2856 (N_2856,N_1570,N_1391);
or U2857 (N_2857,N_1280,N_1640);
and U2858 (N_2858,N_1855,N_1431);
nor U2859 (N_2859,N_1792,N_1191);
or U2860 (N_2860,N_1837,N_1820);
nand U2861 (N_2861,N_1511,N_1061);
nor U2862 (N_2862,N_1747,N_1371);
nor U2863 (N_2863,N_1466,N_1670);
or U2864 (N_2864,N_1895,N_1103);
nor U2865 (N_2865,N_1684,N_1174);
and U2866 (N_2866,N_1573,N_1209);
or U2867 (N_2867,N_1801,N_1481);
nand U2868 (N_2868,N_1628,N_1160);
nand U2869 (N_2869,N_1437,N_1932);
or U2870 (N_2870,N_1678,N_1837);
and U2871 (N_2871,N_1264,N_1031);
nor U2872 (N_2872,N_1590,N_1470);
nand U2873 (N_2873,N_1181,N_1481);
or U2874 (N_2874,N_1432,N_1456);
nor U2875 (N_2875,N_1293,N_1895);
nor U2876 (N_2876,N_1027,N_1540);
or U2877 (N_2877,N_1331,N_1864);
or U2878 (N_2878,N_1699,N_1392);
nand U2879 (N_2879,N_1709,N_1784);
nand U2880 (N_2880,N_1844,N_1970);
and U2881 (N_2881,N_1771,N_1999);
and U2882 (N_2882,N_1619,N_1347);
nor U2883 (N_2883,N_1276,N_1990);
nand U2884 (N_2884,N_1822,N_1952);
nand U2885 (N_2885,N_1441,N_1217);
and U2886 (N_2886,N_1334,N_1605);
or U2887 (N_2887,N_1699,N_1865);
or U2888 (N_2888,N_1065,N_1679);
or U2889 (N_2889,N_1660,N_1111);
or U2890 (N_2890,N_1511,N_1957);
nand U2891 (N_2891,N_1012,N_1082);
or U2892 (N_2892,N_1744,N_1639);
and U2893 (N_2893,N_1414,N_1715);
nor U2894 (N_2894,N_1944,N_1148);
and U2895 (N_2895,N_1714,N_1624);
nand U2896 (N_2896,N_1146,N_1896);
and U2897 (N_2897,N_1309,N_1132);
nand U2898 (N_2898,N_1086,N_1298);
and U2899 (N_2899,N_1425,N_1526);
and U2900 (N_2900,N_1518,N_1164);
nor U2901 (N_2901,N_1633,N_1459);
xnor U2902 (N_2902,N_1262,N_1606);
and U2903 (N_2903,N_1490,N_1980);
xor U2904 (N_2904,N_1313,N_1772);
and U2905 (N_2905,N_1170,N_1459);
and U2906 (N_2906,N_1938,N_1245);
nand U2907 (N_2907,N_1640,N_1746);
or U2908 (N_2908,N_1506,N_1771);
and U2909 (N_2909,N_1806,N_1664);
nor U2910 (N_2910,N_1411,N_1572);
xnor U2911 (N_2911,N_1489,N_1410);
nand U2912 (N_2912,N_1182,N_1084);
xor U2913 (N_2913,N_1883,N_1576);
nor U2914 (N_2914,N_1667,N_1527);
or U2915 (N_2915,N_1960,N_1034);
and U2916 (N_2916,N_1589,N_1227);
nand U2917 (N_2917,N_1621,N_1374);
or U2918 (N_2918,N_1973,N_1369);
nor U2919 (N_2919,N_1568,N_1617);
nor U2920 (N_2920,N_1433,N_1612);
nand U2921 (N_2921,N_1753,N_1410);
or U2922 (N_2922,N_1679,N_1458);
or U2923 (N_2923,N_1282,N_1445);
xor U2924 (N_2924,N_1307,N_1004);
and U2925 (N_2925,N_1838,N_1970);
and U2926 (N_2926,N_1515,N_1006);
or U2927 (N_2927,N_1536,N_1963);
nand U2928 (N_2928,N_1670,N_1023);
nand U2929 (N_2929,N_1217,N_1759);
nor U2930 (N_2930,N_1339,N_1876);
and U2931 (N_2931,N_1758,N_1700);
nor U2932 (N_2932,N_1694,N_1540);
nand U2933 (N_2933,N_1702,N_1197);
and U2934 (N_2934,N_1268,N_1269);
and U2935 (N_2935,N_1953,N_1369);
and U2936 (N_2936,N_1175,N_1349);
or U2937 (N_2937,N_1766,N_1265);
nand U2938 (N_2938,N_1822,N_1824);
and U2939 (N_2939,N_1168,N_1006);
or U2940 (N_2940,N_1483,N_1633);
nor U2941 (N_2941,N_1651,N_1642);
nor U2942 (N_2942,N_1198,N_1416);
nand U2943 (N_2943,N_1195,N_1679);
nand U2944 (N_2944,N_1751,N_1434);
nand U2945 (N_2945,N_1878,N_1533);
nor U2946 (N_2946,N_1101,N_1775);
and U2947 (N_2947,N_1247,N_1032);
nor U2948 (N_2948,N_1673,N_1817);
nand U2949 (N_2949,N_1012,N_1475);
nor U2950 (N_2950,N_1794,N_1790);
and U2951 (N_2951,N_1723,N_1430);
or U2952 (N_2952,N_1384,N_1089);
nor U2953 (N_2953,N_1065,N_1182);
and U2954 (N_2954,N_1848,N_1658);
or U2955 (N_2955,N_1839,N_1287);
nand U2956 (N_2956,N_1039,N_1299);
or U2957 (N_2957,N_1042,N_1528);
nor U2958 (N_2958,N_1141,N_1530);
nor U2959 (N_2959,N_1359,N_1439);
nand U2960 (N_2960,N_1068,N_1153);
or U2961 (N_2961,N_1947,N_1757);
and U2962 (N_2962,N_1944,N_1075);
nand U2963 (N_2963,N_1427,N_1363);
nand U2964 (N_2964,N_1232,N_1249);
nand U2965 (N_2965,N_1845,N_1646);
nand U2966 (N_2966,N_1281,N_1862);
nand U2967 (N_2967,N_1537,N_1787);
and U2968 (N_2968,N_1784,N_1337);
and U2969 (N_2969,N_1728,N_1848);
and U2970 (N_2970,N_1756,N_1971);
nor U2971 (N_2971,N_1872,N_1484);
nor U2972 (N_2972,N_1094,N_1242);
nor U2973 (N_2973,N_1408,N_1304);
and U2974 (N_2974,N_1428,N_1902);
and U2975 (N_2975,N_1380,N_1841);
nand U2976 (N_2976,N_1475,N_1728);
or U2977 (N_2977,N_1392,N_1906);
and U2978 (N_2978,N_1982,N_1797);
or U2979 (N_2979,N_1828,N_1019);
or U2980 (N_2980,N_1453,N_1874);
and U2981 (N_2981,N_1426,N_1972);
and U2982 (N_2982,N_1941,N_1772);
or U2983 (N_2983,N_1480,N_1412);
and U2984 (N_2984,N_1657,N_1976);
and U2985 (N_2985,N_1295,N_1915);
and U2986 (N_2986,N_1305,N_1796);
nor U2987 (N_2987,N_1007,N_1439);
and U2988 (N_2988,N_1978,N_1615);
nand U2989 (N_2989,N_1405,N_1737);
or U2990 (N_2990,N_1434,N_1146);
nand U2991 (N_2991,N_1641,N_1711);
or U2992 (N_2992,N_1826,N_1751);
nand U2993 (N_2993,N_1744,N_1835);
and U2994 (N_2994,N_1061,N_1890);
nand U2995 (N_2995,N_1175,N_1001);
nand U2996 (N_2996,N_1803,N_1455);
and U2997 (N_2997,N_1415,N_1660);
nand U2998 (N_2998,N_1389,N_1539);
nor U2999 (N_2999,N_1275,N_1500);
nand U3000 (N_3000,N_2318,N_2263);
nand U3001 (N_3001,N_2904,N_2385);
nor U3002 (N_3002,N_2211,N_2028);
nand U3003 (N_3003,N_2353,N_2450);
or U3004 (N_3004,N_2189,N_2221);
and U3005 (N_3005,N_2215,N_2696);
nand U3006 (N_3006,N_2614,N_2136);
nand U3007 (N_3007,N_2245,N_2514);
nor U3008 (N_3008,N_2827,N_2980);
nand U3009 (N_3009,N_2192,N_2570);
or U3010 (N_3010,N_2493,N_2368);
xor U3011 (N_3011,N_2947,N_2473);
or U3012 (N_3012,N_2411,N_2715);
nor U3013 (N_3013,N_2174,N_2400);
or U3014 (N_3014,N_2191,N_2195);
nor U3015 (N_3015,N_2084,N_2374);
nor U3016 (N_3016,N_2573,N_2212);
and U3017 (N_3017,N_2319,N_2496);
and U3018 (N_3018,N_2394,N_2405);
nor U3019 (N_3019,N_2160,N_2476);
nand U3020 (N_3020,N_2105,N_2659);
and U3021 (N_3021,N_2726,N_2973);
or U3022 (N_3022,N_2623,N_2092);
and U3023 (N_3023,N_2046,N_2963);
and U3024 (N_3024,N_2009,N_2870);
nand U3025 (N_3025,N_2333,N_2860);
and U3026 (N_3026,N_2356,N_2499);
nor U3027 (N_3027,N_2054,N_2932);
and U3028 (N_3028,N_2812,N_2579);
nor U3029 (N_3029,N_2455,N_2223);
and U3030 (N_3030,N_2267,N_2996);
xnor U3031 (N_3031,N_2995,N_2924);
nand U3032 (N_3032,N_2808,N_2561);
nand U3033 (N_3033,N_2178,N_2705);
or U3034 (N_3034,N_2361,N_2880);
or U3035 (N_3035,N_2372,N_2020);
or U3036 (N_3036,N_2422,N_2509);
nand U3037 (N_3037,N_2882,N_2930);
nand U3038 (N_3038,N_2261,N_2923);
and U3039 (N_3039,N_2384,N_2665);
or U3040 (N_3040,N_2065,N_2822);
nor U3041 (N_3041,N_2584,N_2828);
or U3042 (N_3042,N_2453,N_2586);
nor U3043 (N_3043,N_2602,N_2551);
nand U3044 (N_3044,N_2644,N_2108);
and U3045 (N_3045,N_2007,N_2064);
nor U3046 (N_3046,N_2554,N_2595);
xor U3047 (N_3047,N_2658,N_2596);
nand U3048 (N_3048,N_2617,N_2480);
or U3049 (N_3049,N_2601,N_2866);
nor U3050 (N_3050,N_2387,N_2537);
or U3051 (N_3051,N_2100,N_2327);
and U3052 (N_3052,N_2734,N_2910);
and U3053 (N_3053,N_2430,N_2180);
nand U3054 (N_3054,N_2317,N_2343);
nand U3055 (N_3055,N_2226,N_2477);
and U3056 (N_3056,N_2764,N_2663);
nor U3057 (N_3057,N_2116,N_2294);
or U3058 (N_3058,N_2351,N_2655);
nand U3059 (N_3059,N_2578,N_2867);
and U3060 (N_3060,N_2155,N_2194);
and U3061 (N_3061,N_2110,N_2558);
and U3062 (N_3062,N_2058,N_2909);
or U3063 (N_3063,N_2606,N_2287);
nand U3064 (N_3064,N_2919,N_2720);
nor U3065 (N_3065,N_2711,N_2671);
nand U3066 (N_3066,N_2692,N_2086);
nor U3067 (N_3067,N_2814,N_2145);
xnor U3068 (N_3068,N_2627,N_2396);
and U3069 (N_3069,N_2684,N_2024);
nor U3070 (N_3070,N_2251,N_2774);
and U3071 (N_3071,N_2890,N_2953);
nand U3072 (N_3072,N_2414,N_2666);
nand U3073 (N_3073,N_2399,N_2798);
and U3074 (N_3074,N_2735,N_2202);
and U3075 (N_3075,N_2725,N_2817);
and U3076 (N_3076,N_2304,N_2795);
or U3077 (N_3077,N_2687,N_2161);
nor U3078 (N_3078,N_2971,N_2714);
nand U3079 (N_3079,N_2873,N_2470);
and U3080 (N_3080,N_2299,N_2442);
nor U3081 (N_3081,N_2184,N_2707);
nand U3082 (N_3082,N_2522,N_2447);
or U3083 (N_3083,N_2926,N_2111);
and U3084 (N_3084,N_2106,N_2605);
nor U3085 (N_3085,N_2029,N_2902);
nor U3086 (N_3086,N_2490,N_2373);
or U3087 (N_3087,N_2213,N_2790);
nor U3088 (N_3088,N_2330,N_2437);
nor U3089 (N_3089,N_2062,N_2527);
and U3090 (N_3090,N_2694,N_2102);
nand U3091 (N_3091,N_2320,N_2047);
and U3092 (N_3092,N_2367,N_2463);
or U3093 (N_3093,N_2598,N_2557);
nand U3094 (N_3094,N_2364,N_2646);
nor U3095 (N_3095,N_2335,N_2744);
nor U3096 (N_3096,N_2885,N_2495);
or U3097 (N_3097,N_2901,N_2457);
nor U3098 (N_3098,N_2234,N_2154);
and U3099 (N_3099,N_2847,N_2152);
or U3100 (N_3100,N_2432,N_2148);
nand U3101 (N_3101,N_2849,N_2197);
or U3102 (N_3102,N_2994,N_2324);
nor U3103 (N_3103,N_2289,N_2278);
nor U3104 (N_3104,N_2440,N_2162);
and U3105 (N_3105,N_2260,N_2295);
nand U3106 (N_3106,N_2042,N_2780);
nor U3107 (N_3107,N_2560,N_2546);
and U3108 (N_3108,N_2378,N_2507);
and U3109 (N_3109,N_2183,N_2445);
and U3110 (N_3110,N_2826,N_2208);
nand U3111 (N_3111,N_2163,N_2231);
nor U3112 (N_3112,N_2738,N_2946);
nor U3113 (N_3113,N_2066,N_2695);
nand U3114 (N_3114,N_2533,N_2887);
and U3115 (N_3115,N_2079,N_2217);
and U3116 (N_3116,N_2563,N_2959);
and U3117 (N_3117,N_2371,N_2182);
nor U3118 (N_3118,N_2369,N_2270);
nor U3119 (N_3119,N_2977,N_2392);
or U3120 (N_3120,N_2346,N_2265);
nor U3121 (N_3121,N_2697,N_2002);
nor U3122 (N_3122,N_2503,N_2017);
or U3123 (N_3123,N_2168,N_2094);
nor U3124 (N_3124,N_2326,N_2843);
and U3125 (N_3125,N_2088,N_2433);
nor U3126 (N_3126,N_2719,N_2500);
and U3127 (N_3127,N_2815,N_2417);
nor U3128 (N_3128,N_2583,N_2948);
nor U3129 (N_3129,N_2104,N_2908);
nor U3130 (N_3130,N_2489,N_2199);
and U3131 (N_3131,N_2669,N_2166);
nor U3132 (N_3132,N_2892,N_2524);
nor U3133 (N_3133,N_2954,N_2481);
and U3134 (N_3134,N_2772,N_2135);
nor U3135 (N_3135,N_2675,N_2733);
or U3136 (N_3136,N_2091,N_2019);
nand U3137 (N_3137,N_2139,N_2298);
or U3138 (N_3138,N_2642,N_2253);
nor U3139 (N_3139,N_2545,N_2159);
nand U3140 (N_3140,N_2210,N_2142);
or U3141 (N_3141,N_2051,N_2750);
or U3142 (N_3142,N_2539,N_2006);
nand U3143 (N_3143,N_2264,N_2991);
nand U3144 (N_3144,N_2087,N_2126);
and U3145 (N_3145,N_2616,N_2363);
nand U3146 (N_3146,N_2760,N_2407);
or U3147 (N_3147,N_2775,N_2138);
or U3148 (N_3148,N_2370,N_2275);
nor U3149 (N_3149,N_2763,N_2296);
nor U3150 (N_3150,N_2460,N_2582);
nor U3151 (N_3151,N_2331,N_2678);
nand U3152 (N_3152,N_2300,N_2063);
or U3153 (N_3153,N_2703,N_2864);
or U3154 (N_3154,N_2724,N_2742);
and U3155 (N_3155,N_2905,N_2376);
nor U3156 (N_3156,N_2525,N_2248);
nand U3157 (N_3157,N_2884,N_2032);
and U3158 (N_3158,N_2801,N_2841);
nand U3159 (N_3159,N_2033,N_2409);
nor U3160 (N_3160,N_2342,N_2876);
or U3161 (N_3161,N_2730,N_2421);
nand U3162 (N_3162,N_2836,N_2941);
nand U3163 (N_3163,N_2482,N_2016);
or U3164 (N_3164,N_2768,N_2117);
or U3165 (N_3165,N_2829,N_2577);
nor U3166 (N_3166,N_2955,N_2816);
nand U3167 (N_3167,N_2528,N_2740);
or U3168 (N_3168,N_2165,N_2201);
nor U3169 (N_3169,N_2676,N_2049);
nor U3170 (N_3170,N_2259,N_2030);
nor U3171 (N_3171,N_2842,N_2284);
nand U3172 (N_3172,N_2280,N_2428);
or U3173 (N_3173,N_2523,N_2747);
nand U3174 (N_3174,N_2920,N_2293);
nand U3175 (N_3175,N_2788,N_2095);
or U3176 (N_3176,N_2938,N_2940);
nor U3177 (N_3177,N_2505,N_2756);
and U3178 (N_3178,N_2883,N_2521);
nand U3179 (N_3179,N_2365,N_2393);
nor U3180 (N_3180,N_2518,N_2000);
nor U3181 (N_3181,N_2581,N_2519);
nand U3182 (N_3182,N_2220,N_2746);
and U3183 (N_3183,N_2475,N_2618);
or U3184 (N_3184,N_2246,N_2027);
nor U3185 (N_3185,N_2322,N_2691);
or U3186 (N_3186,N_2629,N_2609);
or U3187 (N_3187,N_2585,N_2262);
nor U3188 (N_3188,N_2674,N_2636);
nand U3189 (N_3189,N_2188,N_2698);
nand U3190 (N_3190,N_2778,N_2472);
and U3191 (N_3191,N_2757,N_2965);
and U3192 (N_3192,N_2978,N_2983);
nand U3193 (N_3193,N_2562,N_2288);
or U3194 (N_3194,N_2532,N_2244);
and U3195 (N_3195,N_2951,N_2358);
and U3196 (N_3196,N_2332,N_2127);
nor U3197 (N_3197,N_2818,N_2269);
or U3198 (N_3198,N_2881,N_2310);
nor U3199 (N_3199,N_2968,N_2530);
and U3200 (N_3200,N_2039,N_2120);
nor U3201 (N_3201,N_2654,N_2918);
nor U3202 (N_3202,N_2336,N_2990);
nand U3203 (N_3203,N_2101,N_2803);
or U3204 (N_3204,N_2141,N_2035);
nor U3205 (N_3205,N_2787,N_2082);
or U3206 (N_3206,N_2534,N_2593);
nor U3207 (N_3207,N_2282,N_2809);
nand U3208 (N_3208,N_2594,N_2693);
nand U3209 (N_3209,N_2034,N_2588);
or U3210 (N_3210,N_2179,N_2660);
or U3211 (N_3211,N_2540,N_2751);
or U3212 (N_3212,N_2429,N_2567);
nor U3213 (N_3213,N_2709,N_2648);
nand U3214 (N_3214,N_2877,N_2786);
nor U3215 (N_3215,N_2799,N_2680);
or U3216 (N_3216,N_2410,N_2230);
nor U3217 (N_3217,N_2468,N_2115);
and U3218 (N_3218,N_2303,N_2633);
nand U3219 (N_3219,N_2690,N_2053);
xor U3220 (N_3220,N_2541,N_2498);
and U3221 (N_3221,N_2899,N_2982);
and U3222 (N_3222,N_2435,N_2869);
nor U3223 (N_3223,N_2825,N_2339);
and U3224 (N_3224,N_2257,N_2390);
or U3225 (N_3225,N_2664,N_2471);
nor U3226 (N_3226,N_2717,N_2357);
or U3227 (N_3227,N_2382,N_2837);
or U3228 (N_3228,N_2914,N_2173);
nor U3229 (N_3229,N_2931,N_2792);
nand U3230 (N_3230,N_2640,N_2060);
and U3231 (N_3231,N_2713,N_2439);
or U3232 (N_3232,N_2626,N_2635);
nor U3233 (N_3233,N_2939,N_2279);
nand U3234 (N_3234,N_2743,N_2689);
nor U3235 (N_3235,N_2891,N_2085);
nor U3236 (N_3236,N_2894,N_2458);
nand U3237 (N_3237,N_2972,N_2340);
and U3238 (N_3238,N_2526,N_2942);
or U3239 (N_3239,N_2395,N_2144);
xnor U3240 (N_3240,N_2441,N_2607);
nor U3241 (N_3241,N_2992,N_2250);
and U3242 (N_3242,N_2728,N_2896);
and U3243 (N_3243,N_2121,N_2164);
nand U3244 (N_3244,N_2542,N_2677);
or U3245 (N_3245,N_2716,N_2590);
or U3246 (N_3246,N_2113,N_2846);
and U3247 (N_3247,N_2611,N_2258);
nand U3248 (N_3248,N_2078,N_2469);
nand U3249 (N_3249,N_2456,N_2181);
or U3250 (N_3250,N_2190,N_2454);
or U3251 (N_3251,N_2810,N_2097);
nand U3252 (N_3252,N_2535,N_2416);
nor U3253 (N_3253,N_2449,N_2451);
and U3254 (N_3254,N_2037,N_2425);
and U3255 (N_3255,N_2576,N_2137);
nor U3256 (N_3256,N_2015,N_2388);
and U3257 (N_3257,N_2124,N_2966);
nor U3258 (N_3258,N_2794,N_2071);
nand U3259 (N_3259,N_2132,N_2315);
and U3260 (N_3260,N_2819,N_2737);
and U3261 (N_3261,N_2222,N_2712);
nand U3262 (N_3262,N_2538,N_2824);
and U3263 (N_3263,N_2831,N_2083);
nand U3264 (N_3264,N_2272,N_2653);
and U3265 (N_3265,N_2987,N_2797);
nand U3266 (N_3266,N_2804,N_2699);
nand U3267 (N_3267,N_2861,N_2397);
nand U3268 (N_3268,N_2549,N_2249);
nand U3269 (N_3269,N_2044,N_2520);
and U3270 (N_3270,N_2625,N_2292);
nand U3271 (N_3271,N_2359,N_2076);
nor U3272 (N_3272,N_2599,N_2912);
or U3273 (N_3273,N_2515,N_2306);
and U3274 (N_3274,N_2309,N_2484);
nor U3275 (N_3275,N_2005,N_2872);
nand U3276 (N_3276,N_2855,N_2638);
and U3277 (N_3277,N_2650,N_2186);
nor U3278 (N_3278,N_2830,N_2402);
and U3279 (N_3279,N_2207,N_2014);
or U3280 (N_3280,N_2377,N_2949);
and U3281 (N_3281,N_2237,N_2858);
nand U3282 (N_3282,N_2957,N_2070);
or U3283 (N_3283,N_2045,N_2158);
nand U3284 (N_3284,N_2820,N_2945);
nand U3285 (N_3285,N_2723,N_2851);
or U3286 (N_3286,N_2893,N_2771);
nand U3287 (N_3287,N_2185,N_2950);
and U3288 (N_3288,N_2967,N_2565);
xnor U3289 (N_3289,N_2485,N_2813);
and U3290 (N_3290,N_2718,N_2895);
nor U3291 (N_3291,N_2604,N_2206);
nor U3292 (N_3292,N_2052,N_2219);
nor U3293 (N_3293,N_2401,N_2436);
nand U3294 (N_3294,N_2307,N_2238);
or U3295 (N_3295,N_2352,N_2273);
nand U3296 (N_3296,N_2670,N_2090);
or U3297 (N_3297,N_2301,N_2026);
and U3298 (N_3298,N_2103,N_2886);
nor U3299 (N_3299,N_2479,N_2125);
or U3300 (N_3300,N_2752,N_2023);
nor U3301 (N_3301,N_2871,N_2898);
nor U3302 (N_3302,N_2235,N_2140);
nor U3303 (N_3303,N_2112,N_2512);
xor U3304 (N_3304,N_2610,N_2175);
or U3305 (N_3305,N_2960,N_2840);
nand U3306 (N_3306,N_2214,N_2917);
and U3307 (N_3307,N_2419,N_2721);
or U3308 (N_3308,N_2759,N_2956);
nand U3309 (N_3309,N_2061,N_2398);
nand U3310 (N_3310,N_2031,N_2271);
nand U3311 (N_3311,N_2227,N_2631);
nand U3312 (N_3312,N_2854,N_2494);
nand U3313 (N_3313,N_2232,N_2732);
nand U3314 (N_3314,N_2193,N_2661);
nor U3315 (N_3315,N_2254,N_2438);
nor U3316 (N_3316,N_2935,N_2649);
or U3317 (N_3317,N_2683,N_2150);
and U3318 (N_3318,N_2970,N_2986);
and U3319 (N_3319,N_2443,N_2900);
nand U3320 (N_3320,N_2952,N_2555);
xnor U3321 (N_3321,N_2656,N_2915);
nand U3322 (N_3322,N_2888,N_2998);
nand U3323 (N_3323,N_2704,N_2408);
or U3324 (N_3324,N_2040,N_2928);
nand U3325 (N_3325,N_2123,N_2838);
nand U3326 (N_3326,N_2686,N_2338);
or U3327 (N_3327,N_2706,N_2427);
and U3328 (N_3328,N_2767,N_2879);
or U3329 (N_3329,N_2412,N_2615);
and U3330 (N_3330,N_2488,N_2321);
or U3331 (N_3331,N_2647,N_2681);
or U3332 (N_3332,N_2073,N_2431);
and U3333 (N_3333,N_2391,N_2710);
or U3334 (N_3334,N_2256,N_2969);
nand U3335 (N_3335,N_2510,N_2651);
nand U3336 (N_3336,N_2922,N_2785);
or U3337 (N_3337,N_2807,N_2462);
or U3338 (N_3338,N_2722,N_2630);
nand U3339 (N_3339,N_2620,N_2652);
and U3340 (N_3340,N_2621,N_2057);
and U3341 (N_3341,N_2056,N_2921);
nand U3342 (N_3342,N_2461,N_2467);
nor U3343 (N_3343,N_2513,N_2613);
nor U3344 (N_3344,N_2552,N_2823);
nand U3345 (N_3345,N_2380,N_2571);
or U3346 (N_3346,N_2362,N_2913);
and U3347 (N_3347,N_2048,N_2933);
nor U3348 (N_3348,N_2003,N_2069);
and U3349 (N_3349,N_2021,N_2536);
nor U3350 (N_3350,N_2997,N_2118);
nand U3351 (N_3351,N_2502,N_2354);
nor U3352 (N_3352,N_2308,N_2143);
or U3353 (N_3353,N_2753,N_2059);
xnor U3354 (N_3354,N_2283,N_2559);
or U3355 (N_3355,N_2679,N_2853);
nor U3356 (N_3356,N_2239,N_2404);
and U3357 (N_3357,N_2682,N_2013);
and U3358 (N_3358,N_2848,N_2156);
and U3359 (N_3359,N_2700,N_2964);
nand U3360 (N_3360,N_2255,N_2415);
or U3361 (N_3361,N_2575,N_2897);
and U3362 (N_3362,N_2464,N_2975);
nor U3363 (N_3363,N_2564,N_2889);
or U3364 (N_3364,N_2566,N_2381);
or U3365 (N_3365,N_2360,N_2770);
and U3366 (N_3366,N_2739,N_2018);
or U3367 (N_3367,N_2348,N_2600);
or U3368 (N_3368,N_2478,N_2266);
and U3369 (N_3369,N_2857,N_2688);
nor U3370 (N_3370,N_2568,N_2247);
nor U3371 (N_3371,N_2313,N_2286);
and U3372 (N_3372,N_2001,N_2749);
nand U3373 (N_3373,N_2821,N_2741);
nand U3374 (N_3374,N_2011,N_2218);
or U3375 (N_3375,N_2762,N_2334);
nor U3376 (N_3376,N_2448,N_2999);
nand U3377 (N_3377,N_2727,N_2597);
nor U3378 (N_3378,N_2171,N_2934);
nand U3379 (N_3379,N_2129,N_2167);
nor U3380 (N_3380,N_2784,N_2268);
nand U3381 (N_3381,N_2022,N_2375);
nand U3382 (N_3382,N_2632,N_2242);
and U3383 (N_3383,N_2157,N_2107);
nor U3384 (N_3384,N_2349,N_2589);
nand U3385 (N_3385,N_2662,N_2834);
or U3386 (N_3386,N_2311,N_2444);
nand U3387 (N_3387,N_2765,N_2119);
or U3388 (N_3388,N_2731,N_2592);
and U3389 (N_3389,N_2976,N_2093);
or U3390 (N_3390,N_2233,N_2203);
and U3391 (N_3391,N_2929,N_2151);
or U3392 (N_3392,N_2859,N_2702);
or U3393 (N_3393,N_2243,N_2755);
xnor U3394 (N_3394,N_2511,N_2745);
nand U3395 (N_3395,N_2989,N_2641);
xor U3396 (N_3396,N_2529,N_2010);
nor U3397 (N_3397,N_2645,N_2835);
nor U3398 (N_3398,N_2216,N_2506);
or U3399 (N_3399,N_2769,N_2277);
nor U3400 (N_3400,N_2802,N_2783);
xnor U3401 (N_3401,N_2036,N_2122);
or U3402 (N_3402,N_2608,N_2133);
and U3403 (N_3403,N_2228,N_2386);
nor U3404 (N_3404,N_2782,N_2556);
or U3405 (N_3405,N_2043,N_2067);
or U3406 (N_3406,N_2572,N_2668);
and U3407 (N_3407,N_2096,N_2341);
nor U3408 (N_3408,N_2544,N_2981);
nor U3409 (N_3409,N_2205,N_2177);
or U3410 (N_3410,N_2172,N_2789);
and U3411 (N_3411,N_2038,N_2350);
nor U3412 (N_3412,N_2302,N_2281);
nor U3413 (N_3413,N_2548,N_2791);
nand U3414 (N_3414,N_2553,N_2196);
nor U3415 (N_3415,N_2209,N_2850);
nor U3416 (N_3416,N_2793,N_2875);
and U3417 (N_3417,N_2673,N_2974);
nand U3418 (N_3418,N_2466,N_2345);
or U3419 (N_3419,N_2314,N_2634);
nor U3420 (N_3420,N_2114,N_2420);
and U3421 (N_3421,N_2657,N_2988);
nand U3422 (N_3422,N_2543,N_2291);
nor U3423 (N_3423,N_2487,N_2832);
or U3424 (N_3424,N_2225,N_2916);
and U3425 (N_3425,N_2619,N_2497);
nor U3426 (N_3426,N_2501,N_2077);
nand U3427 (N_3427,N_2531,N_2580);
nand U3428 (N_3428,N_2406,N_2591);
and U3429 (N_3429,N_2492,N_2587);
nor U3430 (N_3430,N_2628,N_2486);
or U3431 (N_3431,N_2758,N_2459);
nand U3432 (N_3432,N_2383,N_2491);
and U3433 (N_3433,N_2779,N_2911);
or U3434 (N_3434,N_2347,N_2622);
or U3435 (N_3435,N_2241,N_2041);
nor U3436 (N_3436,N_2639,N_2252);
or U3437 (N_3437,N_2569,N_2483);
and U3438 (N_3438,N_2961,N_2907);
nor U3439 (N_3439,N_2081,N_2413);
or U3440 (N_3440,N_2147,N_2080);
and U3441 (N_3441,N_2766,N_2574);
or U3442 (N_3442,N_2344,N_2637);
or U3443 (N_3443,N_2329,N_2776);
and U3444 (N_3444,N_2603,N_2856);
nand U3445 (N_3445,N_2229,N_2075);
and U3446 (N_3446,N_2833,N_2985);
and U3447 (N_3447,N_2379,N_2134);
nor U3448 (N_3448,N_2805,N_2130);
and U3449 (N_3449,N_2773,N_2153);
nand U3450 (N_3450,N_2781,N_2424);
nor U3451 (N_3451,N_2099,N_2811);
and U3452 (N_3452,N_2806,N_2906);
nor U3453 (N_3453,N_2878,N_2667);
and U3454 (N_3454,N_2672,N_2925);
nand U3455 (N_3455,N_2012,N_2055);
nor U3456 (N_3456,N_2170,N_2474);
and U3457 (N_3457,N_2403,N_2204);
and U3458 (N_3458,N_2297,N_2927);
or U3459 (N_3459,N_2944,N_2426);
nor U3460 (N_3460,N_2937,N_2285);
or U3461 (N_3461,N_2050,N_2187);
or U3462 (N_3462,N_2550,N_2305);
nor U3463 (N_3463,N_2962,N_2852);
and U3464 (N_3464,N_2748,N_2423);
or U3465 (N_3465,N_2612,N_2072);
or U3466 (N_3466,N_2936,N_2979);
nor U3467 (N_3467,N_2736,N_2290);
nor U3468 (N_3468,N_2276,N_2754);
nand U3469 (N_3469,N_2224,N_2337);
nand U3470 (N_3470,N_2729,N_2993);
nand U3471 (N_3471,N_2389,N_2068);
nor U3472 (N_3472,N_2169,N_2465);
or U3473 (N_3473,N_2312,N_2874);
and U3474 (N_3474,N_2236,N_2547);
nand U3475 (N_3475,N_2761,N_2328);
nand U3476 (N_3476,N_2089,N_2074);
or U3477 (N_3477,N_2323,N_2366);
and U3478 (N_3478,N_2903,N_2685);
nor U3479 (N_3479,N_2198,N_2516);
or U3480 (N_3480,N_2839,N_2098);
or U3481 (N_3481,N_2862,N_2504);
nor U3482 (N_3482,N_2240,N_2128);
and U3483 (N_3483,N_2109,N_2517);
nand U3484 (N_3484,N_2025,N_2418);
nor U3485 (N_3485,N_2316,N_2146);
nor U3486 (N_3486,N_2865,N_2446);
and U3487 (N_3487,N_2796,N_2984);
and U3488 (N_3488,N_2643,N_2200);
or U3489 (N_3489,N_2452,N_2701);
xnor U3490 (N_3490,N_2434,N_2863);
xnor U3491 (N_3491,N_2800,N_2844);
or U3492 (N_3492,N_2624,N_2274);
nor U3493 (N_3493,N_2355,N_2176);
and U3494 (N_3494,N_2868,N_2131);
nor U3495 (N_3495,N_2508,N_2777);
nand U3496 (N_3496,N_2958,N_2004);
nor U3497 (N_3497,N_2325,N_2845);
nand U3498 (N_3498,N_2708,N_2943);
nand U3499 (N_3499,N_2149,N_2008);
nand U3500 (N_3500,N_2089,N_2615);
nand U3501 (N_3501,N_2476,N_2980);
nand U3502 (N_3502,N_2259,N_2233);
and U3503 (N_3503,N_2731,N_2478);
nor U3504 (N_3504,N_2587,N_2826);
nand U3505 (N_3505,N_2464,N_2810);
or U3506 (N_3506,N_2789,N_2680);
and U3507 (N_3507,N_2549,N_2201);
or U3508 (N_3508,N_2548,N_2647);
nor U3509 (N_3509,N_2393,N_2463);
nor U3510 (N_3510,N_2682,N_2441);
or U3511 (N_3511,N_2126,N_2437);
and U3512 (N_3512,N_2231,N_2169);
or U3513 (N_3513,N_2130,N_2559);
nor U3514 (N_3514,N_2381,N_2236);
nor U3515 (N_3515,N_2701,N_2511);
and U3516 (N_3516,N_2886,N_2915);
or U3517 (N_3517,N_2895,N_2068);
nand U3518 (N_3518,N_2146,N_2602);
and U3519 (N_3519,N_2263,N_2856);
nand U3520 (N_3520,N_2452,N_2991);
nor U3521 (N_3521,N_2887,N_2464);
or U3522 (N_3522,N_2476,N_2354);
nand U3523 (N_3523,N_2928,N_2948);
or U3524 (N_3524,N_2107,N_2462);
or U3525 (N_3525,N_2044,N_2346);
nor U3526 (N_3526,N_2933,N_2262);
or U3527 (N_3527,N_2326,N_2084);
and U3528 (N_3528,N_2520,N_2658);
and U3529 (N_3529,N_2616,N_2473);
nand U3530 (N_3530,N_2242,N_2062);
or U3531 (N_3531,N_2638,N_2273);
and U3532 (N_3532,N_2927,N_2765);
or U3533 (N_3533,N_2096,N_2739);
nand U3534 (N_3534,N_2768,N_2637);
or U3535 (N_3535,N_2316,N_2053);
and U3536 (N_3536,N_2125,N_2601);
and U3537 (N_3537,N_2548,N_2645);
and U3538 (N_3538,N_2676,N_2170);
nand U3539 (N_3539,N_2540,N_2040);
nor U3540 (N_3540,N_2657,N_2809);
or U3541 (N_3541,N_2265,N_2985);
and U3542 (N_3542,N_2114,N_2513);
nand U3543 (N_3543,N_2493,N_2794);
nand U3544 (N_3544,N_2278,N_2993);
and U3545 (N_3545,N_2242,N_2401);
and U3546 (N_3546,N_2403,N_2634);
nand U3547 (N_3547,N_2049,N_2379);
and U3548 (N_3548,N_2019,N_2353);
or U3549 (N_3549,N_2421,N_2680);
nor U3550 (N_3550,N_2221,N_2413);
and U3551 (N_3551,N_2953,N_2738);
nor U3552 (N_3552,N_2027,N_2071);
or U3553 (N_3553,N_2923,N_2099);
and U3554 (N_3554,N_2376,N_2441);
or U3555 (N_3555,N_2825,N_2377);
nand U3556 (N_3556,N_2003,N_2807);
nand U3557 (N_3557,N_2287,N_2362);
and U3558 (N_3558,N_2173,N_2747);
nor U3559 (N_3559,N_2779,N_2003);
nor U3560 (N_3560,N_2217,N_2988);
nand U3561 (N_3561,N_2912,N_2390);
nor U3562 (N_3562,N_2832,N_2748);
nand U3563 (N_3563,N_2492,N_2516);
nor U3564 (N_3564,N_2086,N_2586);
nand U3565 (N_3565,N_2739,N_2848);
and U3566 (N_3566,N_2150,N_2215);
or U3567 (N_3567,N_2734,N_2536);
nor U3568 (N_3568,N_2986,N_2423);
or U3569 (N_3569,N_2654,N_2813);
or U3570 (N_3570,N_2140,N_2448);
nand U3571 (N_3571,N_2884,N_2870);
nor U3572 (N_3572,N_2704,N_2885);
nor U3573 (N_3573,N_2300,N_2995);
and U3574 (N_3574,N_2341,N_2814);
nor U3575 (N_3575,N_2415,N_2565);
or U3576 (N_3576,N_2303,N_2305);
and U3577 (N_3577,N_2315,N_2548);
or U3578 (N_3578,N_2351,N_2370);
nand U3579 (N_3579,N_2081,N_2986);
nand U3580 (N_3580,N_2443,N_2445);
or U3581 (N_3581,N_2268,N_2375);
and U3582 (N_3582,N_2796,N_2920);
xor U3583 (N_3583,N_2308,N_2598);
nand U3584 (N_3584,N_2248,N_2043);
nand U3585 (N_3585,N_2666,N_2958);
nor U3586 (N_3586,N_2322,N_2422);
or U3587 (N_3587,N_2544,N_2367);
and U3588 (N_3588,N_2683,N_2501);
nor U3589 (N_3589,N_2889,N_2178);
and U3590 (N_3590,N_2860,N_2671);
or U3591 (N_3591,N_2633,N_2710);
or U3592 (N_3592,N_2911,N_2520);
or U3593 (N_3593,N_2425,N_2502);
nor U3594 (N_3594,N_2999,N_2669);
nand U3595 (N_3595,N_2308,N_2311);
nand U3596 (N_3596,N_2644,N_2826);
nor U3597 (N_3597,N_2400,N_2623);
nand U3598 (N_3598,N_2745,N_2832);
and U3599 (N_3599,N_2470,N_2661);
or U3600 (N_3600,N_2869,N_2094);
nand U3601 (N_3601,N_2828,N_2771);
nor U3602 (N_3602,N_2713,N_2534);
or U3603 (N_3603,N_2720,N_2857);
xnor U3604 (N_3604,N_2751,N_2108);
and U3605 (N_3605,N_2605,N_2476);
or U3606 (N_3606,N_2597,N_2549);
and U3607 (N_3607,N_2863,N_2487);
and U3608 (N_3608,N_2629,N_2321);
or U3609 (N_3609,N_2717,N_2756);
nor U3610 (N_3610,N_2383,N_2322);
nand U3611 (N_3611,N_2441,N_2943);
or U3612 (N_3612,N_2591,N_2422);
and U3613 (N_3613,N_2191,N_2677);
and U3614 (N_3614,N_2965,N_2192);
and U3615 (N_3615,N_2452,N_2969);
or U3616 (N_3616,N_2099,N_2654);
nand U3617 (N_3617,N_2366,N_2866);
or U3618 (N_3618,N_2074,N_2018);
or U3619 (N_3619,N_2908,N_2377);
or U3620 (N_3620,N_2588,N_2153);
nor U3621 (N_3621,N_2010,N_2432);
nor U3622 (N_3622,N_2528,N_2048);
nor U3623 (N_3623,N_2063,N_2980);
and U3624 (N_3624,N_2588,N_2538);
or U3625 (N_3625,N_2386,N_2413);
nand U3626 (N_3626,N_2291,N_2027);
nor U3627 (N_3627,N_2414,N_2683);
nand U3628 (N_3628,N_2373,N_2074);
nor U3629 (N_3629,N_2432,N_2223);
nand U3630 (N_3630,N_2664,N_2807);
or U3631 (N_3631,N_2607,N_2586);
and U3632 (N_3632,N_2953,N_2923);
or U3633 (N_3633,N_2488,N_2482);
and U3634 (N_3634,N_2903,N_2630);
nand U3635 (N_3635,N_2687,N_2466);
and U3636 (N_3636,N_2312,N_2566);
nor U3637 (N_3637,N_2879,N_2727);
or U3638 (N_3638,N_2601,N_2411);
or U3639 (N_3639,N_2893,N_2196);
or U3640 (N_3640,N_2995,N_2933);
and U3641 (N_3641,N_2221,N_2669);
or U3642 (N_3642,N_2037,N_2359);
or U3643 (N_3643,N_2564,N_2406);
or U3644 (N_3644,N_2977,N_2197);
xnor U3645 (N_3645,N_2497,N_2635);
nand U3646 (N_3646,N_2142,N_2118);
or U3647 (N_3647,N_2506,N_2154);
or U3648 (N_3648,N_2572,N_2119);
nor U3649 (N_3649,N_2870,N_2343);
and U3650 (N_3650,N_2182,N_2817);
nand U3651 (N_3651,N_2465,N_2108);
nor U3652 (N_3652,N_2556,N_2293);
nand U3653 (N_3653,N_2570,N_2122);
nor U3654 (N_3654,N_2586,N_2135);
or U3655 (N_3655,N_2655,N_2512);
or U3656 (N_3656,N_2654,N_2306);
or U3657 (N_3657,N_2254,N_2585);
and U3658 (N_3658,N_2818,N_2980);
or U3659 (N_3659,N_2587,N_2250);
nand U3660 (N_3660,N_2594,N_2563);
nor U3661 (N_3661,N_2633,N_2389);
nand U3662 (N_3662,N_2392,N_2841);
nand U3663 (N_3663,N_2672,N_2583);
nor U3664 (N_3664,N_2794,N_2082);
or U3665 (N_3665,N_2046,N_2766);
nand U3666 (N_3666,N_2139,N_2159);
nand U3667 (N_3667,N_2279,N_2358);
nand U3668 (N_3668,N_2063,N_2570);
or U3669 (N_3669,N_2602,N_2776);
nor U3670 (N_3670,N_2373,N_2672);
nand U3671 (N_3671,N_2009,N_2040);
or U3672 (N_3672,N_2546,N_2231);
nand U3673 (N_3673,N_2558,N_2660);
or U3674 (N_3674,N_2978,N_2505);
or U3675 (N_3675,N_2418,N_2640);
and U3676 (N_3676,N_2417,N_2399);
and U3677 (N_3677,N_2193,N_2179);
nand U3678 (N_3678,N_2040,N_2565);
and U3679 (N_3679,N_2781,N_2494);
and U3680 (N_3680,N_2677,N_2654);
or U3681 (N_3681,N_2024,N_2762);
and U3682 (N_3682,N_2745,N_2016);
nand U3683 (N_3683,N_2624,N_2860);
xnor U3684 (N_3684,N_2898,N_2616);
nor U3685 (N_3685,N_2882,N_2307);
and U3686 (N_3686,N_2253,N_2786);
nand U3687 (N_3687,N_2461,N_2777);
nand U3688 (N_3688,N_2642,N_2431);
and U3689 (N_3689,N_2371,N_2967);
nor U3690 (N_3690,N_2254,N_2402);
nor U3691 (N_3691,N_2231,N_2748);
nand U3692 (N_3692,N_2989,N_2177);
and U3693 (N_3693,N_2540,N_2197);
or U3694 (N_3694,N_2019,N_2404);
nor U3695 (N_3695,N_2825,N_2156);
nand U3696 (N_3696,N_2235,N_2185);
or U3697 (N_3697,N_2258,N_2964);
nand U3698 (N_3698,N_2560,N_2034);
and U3699 (N_3699,N_2936,N_2393);
nand U3700 (N_3700,N_2694,N_2143);
and U3701 (N_3701,N_2498,N_2443);
or U3702 (N_3702,N_2611,N_2486);
nand U3703 (N_3703,N_2801,N_2891);
or U3704 (N_3704,N_2613,N_2828);
nand U3705 (N_3705,N_2027,N_2492);
nor U3706 (N_3706,N_2635,N_2164);
nand U3707 (N_3707,N_2476,N_2751);
or U3708 (N_3708,N_2310,N_2431);
or U3709 (N_3709,N_2392,N_2450);
and U3710 (N_3710,N_2440,N_2630);
and U3711 (N_3711,N_2103,N_2614);
and U3712 (N_3712,N_2068,N_2029);
nor U3713 (N_3713,N_2407,N_2665);
and U3714 (N_3714,N_2765,N_2869);
nor U3715 (N_3715,N_2285,N_2124);
nand U3716 (N_3716,N_2044,N_2762);
nor U3717 (N_3717,N_2655,N_2540);
or U3718 (N_3718,N_2643,N_2392);
nand U3719 (N_3719,N_2047,N_2689);
and U3720 (N_3720,N_2676,N_2212);
and U3721 (N_3721,N_2234,N_2386);
nor U3722 (N_3722,N_2428,N_2031);
nand U3723 (N_3723,N_2806,N_2131);
nand U3724 (N_3724,N_2430,N_2270);
nand U3725 (N_3725,N_2364,N_2084);
nand U3726 (N_3726,N_2865,N_2703);
nand U3727 (N_3727,N_2874,N_2278);
or U3728 (N_3728,N_2815,N_2903);
or U3729 (N_3729,N_2694,N_2322);
nor U3730 (N_3730,N_2589,N_2933);
nand U3731 (N_3731,N_2327,N_2132);
nor U3732 (N_3732,N_2712,N_2095);
nand U3733 (N_3733,N_2341,N_2446);
nor U3734 (N_3734,N_2585,N_2365);
nor U3735 (N_3735,N_2070,N_2098);
xor U3736 (N_3736,N_2605,N_2847);
or U3737 (N_3737,N_2749,N_2901);
nor U3738 (N_3738,N_2046,N_2747);
and U3739 (N_3739,N_2612,N_2642);
or U3740 (N_3740,N_2483,N_2780);
and U3741 (N_3741,N_2264,N_2903);
nand U3742 (N_3742,N_2499,N_2185);
nor U3743 (N_3743,N_2699,N_2519);
nand U3744 (N_3744,N_2232,N_2044);
and U3745 (N_3745,N_2992,N_2028);
or U3746 (N_3746,N_2988,N_2771);
and U3747 (N_3747,N_2360,N_2748);
xor U3748 (N_3748,N_2291,N_2166);
nand U3749 (N_3749,N_2750,N_2540);
or U3750 (N_3750,N_2876,N_2420);
nand U3751 (N_3751,N_2936,N_2739);
nand U3752 (N_3752,N_2692,N_2404);
nor U3753 (N_3753,N_2019,N_2236);
and U3754 (N_3754,N_2424,N_2473);
nand U3755 (N_3755,N_2913,N_2548);
or U3756 (N_3756,N_2037,N_2622);
nor U3757 (N_3757,N_2415,N_2707);
and U3758 (N_3758,N_2418,N_2502);
nor U3759 (N_3759,N_2943,N_2425);
or U3760 (N_3760,N_2125,N_2645);
nand U3761 (N_3761,N_2769,N_2616);
and U3762 (N_3762,N_2077,N_2376);
nor U3763 (N_3763,N_2777,N_2359);
nor U3764 (N_3764,N_2883,N_2934);
nand U3765 (N_3765,N_2401,N_2821);
and U3766 (N_3766,N_2365,N_2934);
and U3767 (N_3767,N_2020,N_2744);
nor U3768 (N_3768,N_2409,N_2192);
nor U3769 (N_3769,N_2601,N_2630);
or U3770 (N_3770,N_2335,N_2175);
or U3771 (N_3771,N_2956,N_2212);
nand U3772 (N_3772,N_2261,N_2768);
nand U3773 (N_3773,N_2158,N_2732);
and U3774 (N_3774,N_2631,N_2466);
or U3775 (N_3775,N_2398,N_2507);
and U3776 (N_3776,N_2468,N_2856);
and U3777 (N_3777,N_2261,N_2227);
nor U3778 (N_3778,N_2355,N_2425);
nor U3779 (N_3779,N_2755,N_2078);
and U3780 (N_3780,N_2377,N_2811);
nor U3781 (N_3781,N_2554,N_2880);
nor U3782 (N_3782,N_2055,N_2404);
and U3783 (N_3783,N_2647,N_2021);
or U3784 (N_3784,N_2028,N_2729);
nand U3785 (N_3785,N_2231,N_2955);
and U3786 (N_3786,N_2310,N_2036);
nand U3787 (N_3787,N_2422,N_2643);
and U3788 (N_3788,N_2547,N_2180);
nor U3789 (N_3789,N_2493,N_2744);
nand U3790 (N_3790,N_2780,N_2233);
nor U3791 (N_3791,N_2050,N_2265);
nand U3792 (N_3792,N_2067,N_2362);
nor U3793 (N_3793,N_2303,N_2150);
nor U3794 (N_3794,N_2016,N_2972);
nand U3795 (N_3795,N_2206,N_2184);
nor U3796 (N_3796,N_2722,N_2542);
nor U3797 (N_3797,N_2493,N_2951);
and U3798 (N_3798,N_2174,N_2026);
nand U3799 (N_3799,N_2934,N_2615);
or U3800 (N_3800,N_2668,N_2321);
and U3801 (N_3801,N_2983,N_2689);
or U3802 (N_3802,N_2312,N_2980);
and U3803 (N_3803,N_2172,N_2710);
or U3804 (N_3804,N_2476,N_2538);
nand U3805 (N_3805,N_2393,N_2160);
nand U3806 (N_3806,N_2880,N_2383);
nand U3807 (N_3807,N_2967,N_2681);
nand U3808 (N_3808,N_2274,N_2361);
nand U3809 (N_3809,N_2456,N_2890);
nor U3810 (N_3810,N_2265,N_2097);
nand U3811 (N_3811,N_2835,N_2092);
nor U3812 (N_3812,N_2826,N_2873);
and U3813 (N_3813,N_2749,N_2168);
or U3814 (N_3814,N_2702,N_2548);
or U3815 (N_3815,N_2365,N_2604);
or U3816 (N_3816,N_2910,N_2929);
nor U3817 (N_3817,N_2318,N_2025);
nor U3818 (N_3818,N_2813,N_2570);
and U3819 (N_3819,N_2404,N_2297);
nand U3820 (N_3820,N_2142,N_2127);
and U3821 (N_3821,N_2579,N_2555);
and U3822 (N_3822,N_2738,N_2734);
or U3823 (N_3823,N_2895,N_2079);
nor U3824 (N_3824,N_2025,N_2146);
nor U3825 (N_3825,N_2658,N_2562);
and U3826 (N_3826,N_2540,N_2365);
or U3827 (N_3827,N_2736,N_2375);
nand U3828 (N_3828,N_2063,N_2070);
xor U3829 (N_3829,N_2683,N_2956);
nor U3830 (N_3830,N_2418,N_2654);
or U3831 (N_3831,N_2955,N_2924);
or U3832 (N_3832,N_2658,N_2482);
and U3833 (N_3833,N_2864,N_2527);
nand U3834 (N_3834,N_2686,N_2769);
and U3835 (N_3835,N_2566,N_2286);
nand U3836 (N_3836,N_2142,N_2415);
nor U3837 (N_3837,N_2540,N_2651);
nand U3838 (N_3838,N_2555,N_2979);
or U3839 (N_3839,N_2772,N_2967);
nor U3840 (N_3840,N_2170,N_2287);
or U3841 (N_3841,N_2946,N_2604);
or U3842 (N_3842,N_2261,N_2851);
or U3843 (N_3843,N_2338,N_2852);
nor U3844 (N_3844,N_2497,N_2789);
nor U3845 (N_3845,N_2498,N_2737);
or U3846 (N_3846,N_2287,N_2391);
or U3847 (N_3847,N_2058,N_2223);
or U3848 (N_3848,N_2246,N_2842);
nand U3849 (N_3849,N_2872,N_2489);
and U3850 (N_3850,N_2499,N_2877);
or U3851 (N_3851,N_2668,N_2929);
and U3852 (N_3852,N_2612,N_2479);
or U3853 (N_3853,N_2873,N_2404);
and U3854 (N_3854,N_2783,N_2035);
or U3855 (N_3855,N_2677,N_2383);
and U3856 (N_3856,N_2383,N_2748);
and U3857 (N_3857,N_2023,N_2105);
and U3858 (N_3858,N_2026,N_2261);
or U3859 (N_3859,N_2456,N_2718);
nand U3860 (N_3860,N_2274,N_2685);
and U3861 (N_3861,N_2369,N_2275);
and U3862 (N_3862,N_2391,N_2193);
nor U3863 (N_3863,N_2797,N_2400);
or U3864 (N_3864,N_2138,N_2160);
nand U3865 (N_3865,N_2444,N_2423);
nor U3866 (N_3866,N_2413,N_2224);
and U3867 (N_3867,N_2082,N_2871);
nor U3868 (N_3868,N_2981,N_2267);
nor U3869 (N_3869,N_2254,N_2318);
and U3870 (N_3870,N_2372,N_2671);
nand U3871 (N_3871,N_2012,N_2123);
nand U3872 (N_3872,N_2215,N_2241);
or U3873 (N_3873,N_2947,N_2844);
nor U3874 (N_3874,N_2502,N_2944);
and U3875 (N_3875,N_2806,N_2963);
nand U3876 (N_3876,N_2607,N_2221);
nor U3877 (N_3877,N_2835,N_2988);
and U3878 (N_3878,N_2299,N_2726);
and U3879 (N_3879,N_2231,N_2107);
or U3880 (N_3880,N_2146,N_2902);
and U3881 (N_3881,N_2459,N_2300);
and U3882 (N_3882,N_2629,N_2330);
or U3883 (N_3883,N_2756,N_2858);
or U3884 (N_3884,N_2713,N_2484);
nand U3885 (N_3885,N_2143,N_2687);
or U3886 (N_3886,N_2814,N_2744);
nand U3887 (N_3887,N_2344,N_2310);
nor U3888 (N_3888,N_2191,N_2140);
and U3889 (N_3889,N_2526,N_2468);
or U3890 (N_3890,N_2271,N_2852);
or U3891 (N_3891,N_2822,N_2152);
or U3892 (N_3892,N_2509,N_2098);
or U3893 (N_3893,N_2188,N_2991);
and U3894 (N_3894,N_2278,N_2590);
and U3895 (N_3895,N_2415,N_2438);
nor U3896 (N_3896,N_2707,N_2369);
nand U3897 (N_3897,N_2779,N_2806);
nand U3898 (N_3898,N_2901,N_2874);
nor U3899 (N_3899,N_2102,N_2370);
and U3900 (N_3900,N_2382,N_2407);
and U3901 (N_3901,N_2934,N_2844);
nand U3902 (N_3902,N_2644,N_2385);
nand U3903 (N_3903,N_2639,N_2437);
or U3904 (N_3904,N_2328,N_2551);
nor U3905 (N_3905,N_2411,N_2852);
or U3906 (N_3906,N_2847,N_2045);
and U3907 (N_3907,N_2491,N_2072);
or U3908 (N_3908,N_2302,N_2688);
and U3909 (N_3909,N_2643,N_2906);
nand U3910 (N_3910,N_2493,N_2382);
and U3911 (N_3911,N_2916,N_2669);
nor U3912 (N_3912,N_2560,N_2471);
and U3913 (N_3913,N_2625,N_2542);
and U3914 (N_3914,N_2967,N_2407);
and U3915 (N_3915,N_2497,N_2946);
or U3916 (N_3916,N_2124,N_2661);
nand U3917 (N_3917,N_2877,N_2401);
and U3918 (N_3918,N_2929,N_2070);
nand U3919 (N_3919,N_2139,N_2277);
nor U3920 (N_3920,N_2280,N_2645);
or U3921 (N_3921,N_2005,N_2094);
nor U3922 (N_3922,N_2500,N_2746);
and U3923 (N_3923,N_2405,N_2917);
and U3924 (N_3924,N_2014,N_2858);
and U3925 (N_3925,N_2901,N_2054);
nand U3926 (N_3926,N_2627,N_2498);
and U3927 (N_3927,N_2846,N_2901);
nand U3928 (N_3928,N_2963,N_2055);
nor U3929 (N_3929,N_2762,N_2513);
and U3930 (N_3930,N_2184,N_2803);
nor U3931 (N_3931,N_2580,N_2071);
and U3932 (N_3932,N_2135,N_2870);
and U3933 (N_3933,N_2623,N_2214);
or U3934 (N_3934,N_2887,N_2473);
nor U3935 (N_3935,N_2216,N_2408);
nand U3936 (N_3936,N_2540,N_2159);
nand U3937 (N_3937,N_2683,N_2783);
nor U3938 (N_3938,N_2248,N_2392);
or U3939 (N_3939,N_2166,N_2753);
nand U3940 (N_3940,N_2853,N_2749);
or U3941 (N_3941,N_2934,N_2555);
nor U3942 (N_3942,N_2169,N_2485);
nand U3943 (N_3943,N_2339,N_2353);
nor U3944 (N_3944,N_2364,N_2240);
nor U3945 (N_3945,N_2059,N_2621);
and U3946 (N_3946,N_2195,N_2949);
or U3947 (N_3947,N_2604,N_2643);
or U3948 (N_3948,N_2933,N_2578);
nand U3949 (N_3949,N_2985,N_2155);
nor U3950 (N_3950,N_2428,N_2081);
or U3951 (N_3951,N_2116,N_2496);
xnor U3952 (N_3952,N_2411,N_2723);
nor U3953 (N_3953,N_2378,N_2538);
nor U3954 (N_3954,N_2621,N_2159);
nand U3955 (N_3955,N_2601,N_2085);
or U3956 (N_3956,N_2628,N_2640);
nor U3957 (N_3957,N_2045,N_2845);
or U3958 (N_3958,N_2874,N_2298);
and U3959 (N_3959,N_2491,N_2368);
nor U3960 (N_3960,N_2901,N_2960);
and U3961 (N_3961,N_2381,N_2680);
and U3962 (N_3962,N_2619,N_2836);
or U3963 (N_3963,N_2187,N_2485);
and U3964 (N_3964,N_2389,N_2924);
nand U3965 (N_3965,N_2189,N_2445);
xnor U3966 (N_3966,N_2564,N_2067);
nor U3967 (N_3967,N_2682,N_2539);
or U3968 (N_3968,N_2763,N_2121);
and U3969 (N_3969,N_2831,N_2893);
or U3970 (N_3970,N_2374,N_2627);
nor U3971 (N_3971,N_2010,N_2791);
or U3972 (N_3972,N_2943,N_2149);
nand U3973 (N_3973,N_2807,N_2132);
nor U3974 (N_3974,N_2396,N_2502);
and U3975 (N_3975,N_2318,N_2581);
and U3976 (N_3976,N_2797,N_2191);
and U3977 (N_3977,N_2044,N_2591);
and U3978 (N_3978,N_2071,N_2069);
nand U3979 (N_3979,N_2515,N_2839);
nor U3980 (N_3980,N_2335,N_2871);
and U3981 (N_3981,N_2316,N_2182);
and U3982 (N_3982,N_2051,N_2249);
nand U3983 (N_3983,N_2626,N_2566);
or U3984 (N_3984,N_2629,N_2106);
or U3985 (N_3985,N_2199,N_2636);
or U3986 (N_3986,N_2143,N_2106);
nand U3987 (N_3987,N_2691,N_2426);
or U3988 (N_3988,N_2734,N_2142);
nand U3989 (N_3989,N_2758,N_2515);
nand U3990 (N_3990,N_2925,N_2054);
and U3991 (N_3991,N_2207,N_2702);
and U3992 (N_3992,N_2250,N_2885);
nor U3993 (N_3993,N_2408,N_2286);
and U3994 (N_3994,N_2793,N_2509);
and U3995 (N_3995,N_2833,N_2476);
nand U3996 (N_3996,N_2252,N_2787);
or U3997 (N_3997,N_2864,N_2719);
nor U3998 (N_3998,N_2029,N_2534);
xor U3999 (N_3999,N_2099,N_2593);
or U4000 (N_4000,N_3768,N_3266);
and U4001 (N_4001,N_3316,N_3690);
or U4002 (N_4002,N_3815,N_3490);
and U4003 (N_4003,N_3094,N_3204);
or U4004 (N_4004,N_3485,N_3749);
and U4005 (N_4005,N_3072,N_3503);
nor U4006 (N_4006,N_3097,N_3767);
nor U4007 (N_4007,N_3748,N_3597);
and U4008 (N_4008,N_3525,N_3961);
or U4009 (N_4009,N_3776,N_3392);
and U4010 (N_4010,N_3856,N_3281);
nand U4011 (N_4011,N_3543,N_3186);
or U4012 (N_4012,N_3109,N_3249);
and U4013 (N_4013,N_3498,N_3360);
and U4014 (N_4014,N_3358,N_3104);
nor U4015 (N_4015,N_3982,N_3102);
nor U4016 (N_4016,N_3884,N_3053);
and U4017 (N_4017,N_3524,N_3783);
nor U4018 (N_4018,N_3279,N_3998);
nand U4019 (N_4019,N_3652,N_3636);
and U4020 (N_4020,N_3379,N_3665);
or U4021 (N_4021,N_3575,N_3523);
nand U4022 (N_4022,N_3054,N_3489);
nor U4023 (N_4023,N_3931,N_3194);
nand U4024 (N_4024,N_3635,N_3669);
nand U4025 (N_4025,N_3324,N_3828);
nand U4026 (N_4026,N_3165,N_3025);
xor U4027 (N_4027,N_3534,N_3391);
nor U4028 (N_4028,N_3091,N_3300);
or U4029 (N_4029,N_3552,N_3949);
and U4030 (N_4030,N_3028,N_3851);
nor U4031 (N_4031,N_3003,N_3133);
or U4032 (N_4032,N_3223,N_3466);
or U4033 (N_4033,N_3976,N_3247);
nor U4034 (N_4034,N_3447,N_3981);
nand U4035 (N_4035,N_3656,N_3637);
or U4036 (N_4036,N_3873,N_3208);
or U4037 (N_4037,N_3581,N_3607);
or U4038 (N_4038,N_3043,N_3566);
nor U4039 (N_4039,N_3340,N_3659);
nor U4040 (N_4040,N_3892,N_3839);
and U4041 (N_4041,N_3514,N_3101);
nand U4042 (N_4042,N_3163,N_3427);
nor U4043 (N_4043,N_3381,N_3793);
xnor U4044 (N_4044,N_3937,N_3331);
and U4045 (N_4045,N_3728,N_3911);
nand U4046 (N_4046,N_3154,N_3123);
and U4047 (N_4047,N_3402,N_3900);
nand U4048 (N_4048,N_3726,N_3598);
or U4049 (N_4049,N_3295,N_3416);
nor U4050 (N_4050,N_3445,N_3239);
or U4051 (N_4051,N_3022,N_3510);
nor U4052 (N_4052,N_3095,N_3067);
and U4053 (N_4053,N_3007,N_3390);
nor U4054 (N_4054,N_3867,N_3679);
or U4055 (N_4055,N_3940,N_3739);
or U4056 (N_4056,N_3076,N_3660);
and U4057 (N_4057,N_3676,N_3327);
nor U4058 (N_4058,N_3273,N_3755);
or U4059 (N_4059,N_3587,N_3782);
or U4060 (N_4060,N_3435,N_3549);
and U4061 (N_4061,N_3599,N_3866);
nand U4062 (N_4062,N_3137,N_3718);
and U4063 (N_4063,N_3181,N_3605);
or U4064 (N_4064,N_3522,N_3168);
or U4065 (N_4065,N_3332,N_3568);
or U4066 (N_4066,N_3688,N_3772);
and U4067 (N_4067,N_3974,N_3288);
or U4068 (N_4068,N_3929,N_3057);
or U4069 (N_4069,N_3009,N_3257);
or U4070 (N_4070,N_3084,N_3443);
or U4071 (N_4071,N_3662,N_3893);
nand U4072 (N_4072,N_3642,N_3989);
nor U4073 (N_4073,N_3225,N_3577);
and U4074 (N_4074,N_3167,N_3396);
nand U4075 (N_4075,N_3356,N_3500);
nor U4076 (N_4076,N_3362,N_3151);
or U4077 (N_4077,N_3326,N_3978);
and U4078 (N_4078,N_3719,N_3120);
and U4079 (N_4079,N_3244,N_3672);
and U4080 (N_4080,N_3980,N_3818);
and U4081 (N_4081,N_3945,N_3841);
nand U4082 (N_4082,N_3559,N_3730);
nand U4083 (N_4083,N_3077,N_3175);
and U4084 (N_4084,N_3188,N_3214);
nor U4085 (N_4085,N_3070,N_3738);
nor U4086 (N_4086,N_3148,N_3837);
nor U4087 (N_4087,N_3284,N_3130);
nand U4088 (N_4088,N_3275,N_3721);
nor U4089 (N_4089,N_3802,N_3126);
or U4090 (N_4090,N_3617,N_3897);
or U4091 (N_4091,N_3702,N_3848);
and U4092 (N_4092,N_3221,N_3859);
and U4093 (N_4093,N_3339,N_3852);
and U4094 (N_4094,N_3263,N_3840);
xnor U4095 (N_4095,N_3882,N_3086);
or U4096 (N_4096,N_3378,N_3769);
or U4097 (N_4097,N_3424,N_3143);
nor U4098 (N_4098,N_3232,N_3483);
and U4099 (N_4099,N_3805,N_3709);
or U4100 (N_4100,N_3042,N_3314);
nand U4101 (N_4101,N_3171,N_3253);
or U4102 (N_4102,N_3554,N_3680);
nand U4103 (N_4103,N_3363,N_3562);
and U4104 (N_4104,N_3212,N_3317);
nor U4105 (N_4105,N_3634,N_3527);
nand U4106 (N_4106,N_3272,N_3441);
nor U4107 (N_4107,N_3789,N_3894);
or U4108 (N_4108,N_3073,N_3477);
or U4109 (N_4109,N_3140,N_3589);
nor U4110 (N_4110,N_3842,N_3355);
or U4111 (N_4111,N_3712,N_3533);
nand U4112 (N_4112,N_3422,N_3908);
or U4113 (N_4113,N_3472,N_3521);
nor U4114 (N_4114,N_3011,N_3180);
or U4115 (N_4115,N_3258,N_3863);
nor U4116 (N_4116,N_3289,N_3520);
and U4117 (N_4117,N_3578,N_3325);
nor U4118 (N_4118,N_3750,N_3128);
and U4119 (N_4119,N_3613,N_3453);
and U4120 (N_4120,N_3467,N_3801);
nand U4121 (N_4121,N_3087,N_3798);
nor U4122 (N_4122,N_3686,N_3499);
nand U4123 (N_4123,N_3943,N_3517);
and U4124 (N_4124,N_3992,N_3038);
and U4125 (N_4125,N_3838,N_3746);
nand U4126 (N_4126,N_3707,N_3954);
nor U4127 (N_4127,N_3437,N_3752);
nor U4128 (N_4128,N_3546,N_3556);
or U4129 (N_4129,N_3021,N_3398);
nand U4130 (N_4130,N_3735,N_3705);
nor U4131 (N_4131,N_3890,N_3969);
or U4132 (N_4132,N_3925,N_3313);
and U4133 (N_4133,N_3991,N_3306);
nand U4134 (N_4134,N_3387,N_3280);
nor U4135 (N_4135,N_3600,N_3190);
nand U4136 (N_4136,N_3393,N_3995);
nor U4137 (N_4137,N_3569,N_3444);
nand U4138 (N_4138,N_3582,N_3920);
nor U4139 (N_4139,N_3315,N_3384);
and U4140 (N_4140,N_3117,N_3027);
or U4141 (N_4141,N_3891,N_3913);
or U4142 (N_4142,N_3111,N_3687);
xnor U4143 (N_4143,N_3810,N_3001);
nor U4144 (N_4144,N_3450,N_3501);
nor U4145 (N_4145,N_3159,N_3082);
or U4146 (N_4146,N_3189,N_3919);
nor U4147 (N_4147,N_3051,N_3946);
nor U4148 (N_4148,N_3385,N_3304);
nor U4149 (N_4149,N_3220,N_3196);
or U4150 (N_4150,N_3729,N_3256);
nand U4151 (N_4151,N_3080,N_3031);
nor U4152 (N_4152,N_3010,N_3723);
or U4153 (N_4153,N_3948,N_3651);
and U4154 (N_4154,N_3207,N_3865);
nand U4155 (N_4155,N_3098,N_3703);
or U4156 (N_4156,N_3507,N_3791);
nand U4157 (N_4157,N_3487,N_3732);
and U4158 (N_4158,N_3243,N_3184);
or U4159 (N_4159,N_3542,N_3796);
nand U4160 (N_4160,N_3335,N_3606);
and U4161 (N_4161,N_3622,N_3682);
nand U4162 (N_4162,N_3493,N_3696);
or U4163 (N_4163,N_3400,N_3129);
nor U4164 (N_4164,N_3661,N_3085);
and U4165 (N_4165,N_3537,N_3226);
and U4166 (N_4166,N_3431,N_3020);
and U4167 (N_4167,N_3238,N_3417);
and U4168 (N_4168,N_3629,N_3583);
or U4169 (N_4169,N_3348,N_3905);
or U4170 (N_4170,N_3736,N_3200);
nand U4171 (N_4171,N_3853,N_3264);
nand U4172 (N_4172,N_3799,N_3830);
nand U4173 (N_4173,N_3731,N_3904);
and U4174 (N_4174,N_3357,N_3887);
and U4175 (N_4175,N_3488,N_3172);
nor U4176 (N_4176,N_3017,N_3570);
nand U4177 (N_4177,N_3854,N_3177);
nand U4178 (N_4178,N_3685,N_3470);
nand U4179 (N_4179,N_3922,N_3386);
or U4180 (N_4180,N_3794,N_3322);
or U4181 (N_4181,N_3297,N_3650);
and U4182 (N_4182,N_3640,N_3733);
and U4183 (N_4183,N_3013,N_3855);
or U4184 (N_4184,N_3242,N_3780);
nand U4185 (N_4185,N_3278,N_3717);
nand U4186 (N_4186,N_3530,N_3601);
or U4187 (N_4187,N_3955,N_3683);
nor U4188 (N_4188,N_3869,N_3674);
or U4189 (N_4189,N_3142,N_3026);
nor U4190 (N_4190,N_3963,N_3847);
or U4191 (N_4191,N_3495,N_3055);
and U4192 (N_4192,N_3734,N_3135);
or U4193 (N_4193,N_3024,N_3347);
or U4194 (N_4194,N_3246,N_3762);
and U4195 (N_4195,N_3807,N_3408);
and U4196 (N_4196,N_3333,N_3996);
nand U4197 (N_4197,N_3164,N_3059);
nand U4198 (N_4198,N_3227,N_3824);
or U4199 (N_4199,N_3664,N_3078);
nand U4200 (N_4200,N_3228,N_3519);
nand U4201 (N_4201,N_3361,N_3213);
nand U4202 (N_4202,N_3106,N_3299);
nand U4203 (N_4203,N_3504,N_3502);
or U4204 (N_4204,N_3835,N_3404);
nand U4205 (N_4205,N_3083,N_3754);
nand U4206 (N_4206,N_3114,N_3667);
and U4207 (N_4207,N_3480,N_3455);
nor U4208 (N_4208,N_3241,N_3037);
or U4209 (N_4209,N_3074,N_3343);
nand U4210 (N_4210,N_3147,N_3250);
nor U4211 (N_4211,N_3236,N_3162);
nand U4212 (N_4212,N_3293,N_3321);
nand U4213 (N_4213,N_3302,N_3710);
nor U4214 (N_4214,N_3857,N_3486);
and U4215 (N_4215,N_3956,N_3876);
and U4216 (N_4216,N_3345,N_3359);
and U4217 (N_4217,N_3639,N_3591);
nor U4218 (N_4218,N_3697,N_3366);
nand U4219 (N_4219,N_3035,N_3459);
nand U4220 (N_4220,N_3458,N_3144);
nor U4221 (N_4221,N_3179,N_3428);
or U4222 (N_4222,N_3099,N_3370);
or U4223 (N_4223,N_3616,N_3215);
nor U4224 (N_4224,N_3950,N_3457);
nand U4225 (N_4225,N_3108,N_3131);
and U4226 (N_4226,N_3722,N_3328);
and U4227 (N_4227,N_3862,N_3463);
or U4228 (N_4228,N_3985,N_3883);
and U4229 (N_4229,N_3329,N_3045);
and U4230 (N_4230,N_3777,N_3720);
nand U4231 (N_4231,N_3182,N_3727);
or U4232 (N_4232,N_3944,N_3528);
nor U4233 (N_4233,N_3909,N_3896);
nand U4234 (N_4234,N_3513,N_3066);
nor U4235 (N_4235,N_3388,N_3806);
or U4236 (N_4236,N_3870,N_3678);
or U4237 (N_4237,N_3716,N_3382);
nor U4238 (N_4238,N_3973,N_3604);
or U4239 (N_4239,N_3555,N_3364);
nand U4240 (N_4240,N_3088,N_3438);
nor U4241 (N_4241,N_3254,N_3594);
and U4242 (N_4242,N_3781,N_3819);
and U4243 (N_4243,N_3018,N_3689);
and U4244 (N_4244,N_3354,N_3291);
nand U4245 (N_4245,N_3494,N_3574);
and U4246 (N_4246,N_3540,N_3432);
nor U4247 (N_4247,N_3874,N_3725);
nor U4248 (N_4248,N_3039,N_3516);
nor U4249 (N_4249,N_3561,N_3990);
nor U4250 (N_4250,N_3217,N_3849);
or U4251 (N_4251,N_3918,N_3033);
nor U4252 (N_4252,N_3063,N_3365);
nand U4253 (N_4253,N_3633,N_3004);
nand U4254 (N_4254,N_3994,N_3000);
nand U4255 (N_4255,N_3383,N_3609);
or U4256 (N_4256,N_3958,N_3751);
and U4257 (N_4257,N_3538,N_3786);
and U4258 (N_4258,N_3708,N_3089);
and U4259 (N_4259,N_3681,N_3529);
nand U4260 (N_4260,N_3409,N_3218);
nor U4261 (N_4261,N_3002,N_3627);
or U4262 (N_4262,N_3539,N_3462);
nand U4263 (N_4263,N_3713,N_3456);
and U4264 (N_4264,N_3090,N_3820);
and U4265 (N_4265,N_3049,N_3965);
or U4266 (N_4266,N_3939,N_3988);
nor U4267 (N_4267,N_3482,N_3337);
and U4268 (N_4268,N_3684,N_3198);
and U4269 (N_4269,N_3595,N_3704);
and U4270 (N_4270,N_3052,N_3132);
nor U4271 (N_4271,N_3774,N_3262);
nor U4272 (N_4272,N_3715,N_3760);
or U4273 (N_4273,N_3015,N_3816);
nand U4274 (N_4274,N_3967,N_3454);
nor U4275 (N_4275,N_3630,N_3100);
and U4276 (N_4276,N_3927,N_3953);
nand U4277 (N_4277,N_3394,N_3330);
or U4278 (N_4278,N_3193,N_3693);
and U4279 (N_4279,N_3375,N_3825);
nand U4280 (N_4280,N_3512,N_3368);
nor U4281 (N_4281,N_3195,N_3380);
or U4282 (N_4282,N_3334,N_3508);
or U4283 (N_4283,N_3603,N_3511);
and U4284 (N_4284,N_3237,N_3972);
nand U4285 (N_4285,N_3836,N_3319);
or U4286 (N_4286,N_3979,N_3014);
nand U4287 (N_4287,N_3858,N_3318);
or U4288 (N_4288,N_3222,N_3233);
nand U4289 (N_4289,N_3060,N_3871);
and U4290 (N_4290,N_3446,N_3833);
nor U4291 (N_4291,N_3743,N_3473);
and U4292 (N_4292,N_3229,N_3158);
nor U4293 (N_4293,N_3276,N_3023);
and U4294 (N_4294,N_3649,N_3753);
or U4295 (N_4295,N_3584,N_3923);
nand U4296 (N_4296,N_3658,N_3771);
or U4297 (N_4297,N_3641,N_3050);
or U4298 (N_4298,N_3397,N_3742);
nand U4299 (N_4299,N_3061,N_3252);
and U4300 (N_4300,N_3505,N_3115);
and U4301 (N_4301,N_3880,N_3251);
and U4302 (N_4302,N_3210,N_3235);
or U4303 (N_4303,N_3418,N_3934);
or U4304 (N_4304,N_3700,N_3271);
nand U4305 (N_4305,N_3535,N_3541);
nor U4306 (N_4306,N_3645,N_3763);
and U4307 (N_4307,N_3277,N_3558);
nand U4308 (N_4308,N_3079,N_3536);
nand U4309 (N_4309,N_3471,N_3832);
and U4310 (N_4310,N_3691,N_3030);
or U4311 (N_4311,N_3187,N_3987);
xor U4312 (N_4312,N_3610,N_3149);
and U4313 (N_4313,N_3040,N_3515);
nor U4314 (N_4314,N_3758,N_3206);
or U4315 (N_4315,N_3959,N_3579);
and U4316 (N_4316,N_3192,N_3618);
and U4317 (N_4317,N_3544,N_3770);
nand U4318 (N_4318,N_3248,N_3975);
or U4319 (N_4319,N_3756,N_3269);
nand U4320 (N_4320,N_3506,N_3576);
nor U4321 (N_4321,N_3788,N_3434);
or U4322 (N_4322,N_3823,N_3136);
and U4323 (N_4323,N_3166,N_3122);
nand U4324 (N_4324,N_3846,N_3353);
nor U4325 (N_4325,N_3008,N_3296);
nor U4326 (N_4326,N_3588,N_3006);
and U4327 (N_4327,N_3460,N_3898);
nand U4328 (N_4328,N_3121,N_3290);
and U4329 (N_4329,N_3230,N_3492);
or U4330 (N_4330,N_3942,N_3986);
nor U4331 (N_4331,N_3608,N_3046);
nor U4332 (N_4332,N_3968,N_3655);
nand U4333 (N_4333,N_3663,N_3829);
and U4334 (N_4334,N_3778,N_3551);
and U4335 (N_4335,N_3790,N_3211);
nor U4336 (N_4336,N_3984,N_3921);
nor U4337 (N_4337,N_3301,N_3845);
and U4338 (N_4338,N_3926,N_3139);
or U4339 (N_4339,N_3096,N_3917);
nor U4340 (N_4340,N_3265,N_3260);
or U4341 (N_4341,N_3952,N_3532);
or U4342 (N_4342,N_3903,N_3029);
and U4343 (N_4343,N_3351,N_3915);
nand U4344 (N_4344,N_3938,N_3877);
nor U4345 (N_4345,N_3653,N_3294);
and U4346 (N_4346,N_3930,N_3270);
nor U4347 (N_4347,N_3231,N_3881);
nor U4348 (N_4348,N_3071,N_3474);
nand U4349 (N_4349,N_3827,N_3107);
nor U4350 (N_4350,N_3421,N_3425);
nand U4351 (N_4351,N_3625,N_3668);
nand U4352 (N_4352,N_3548,N_3414);
nor U4353 (N_4353,N_3861,N_3626);
or U4354 (N_4354,N_3412,N_3119);
nand U4355 (N_4355,N_3047,N_3797);
or U4356 (N_4356,N_3803,N_3879);
nor U4357 (N_4357,N_3369,N_3932);
nor U4358 (N_4358,N_3936,N_3176);
or U4359 (N_4359,N_3062,N_3349);
nor U4360 (N_4360,N_3415,N_3912);
nand U4361 (N_4361,N_3563,N_3423);
or U4362 (N_4362,N_3478,N_3413);
nand U4363 (N_4363,N_3110,N_3309);
and U4364 (N_4364,N_3970,N_3401);
nor U4365 (N_4365,N_3906,N_3872);
and U4366 (N_4366,N_3469,N_3757);
and U4367 (N_4367,N_3560,N_3614);
and U4368 (N_4368,N_3878,N_3885);
nor U4369 (N_4369,N_3312,N_3962);
and U4370 (N_4370,N_3699,N_3307);
and U4371 (N_4371,N_3621,N_3916);
nand U4372 (N_4372,N_3161,N_3553);
nor U4373 (N_4373,N_3675,N_3202);
nor U4374 (N_4374,N_3886,N_3191);
or U4375 (N_4375,N_3285,N_3826);
xor U4376 (N_4376,N_3268,N_3644);
and U4377 (N_4377,N_3673,N_3411);
nand U4378 (N_4378,N_3367,N_3804);
nand U4379 (N_4379,N_3889,N_3150);
and U4380 (N_4380,N_3888,N_3138);
and U4381 (N_4381,N_3407,N_3596);
nor U4382 (N_4382,N_3283,N_3638);
and U4383 (N_4383,N_3765,N_3779);
nand U4384 (N_4384,N_3183,N_3311);
or U4385 (N_4385,N_3174,N_3924);
nand U4386 (N_4386,N_3844,N_3240);
nand U4387 (N_4387,N_3694,N_3695);
and U4388 (N_4388,N_3116,N_3267);
and U4389 (N_4389,N_3058,N_3547);
and U4390 (N_4390,N_3737,N_3395);
nand U4391 (N_4391,N_3479,N_3298);
nand U4392 (N_4392,N_3580,N_3773);
or U4393 (N_4393,N_3666,N_3376);
nor U4394 (N_4394,N_3817,N_3373);
or U4395 (N_4395,N_3744,N_3567);
and U4396 (N_4396,N_3624,N_3766);
nand U4397 (N_4397,N_3999,N_3813);
nand U4398 (N_4398,N_3775,N_3468);
or U4399 (N_4399,N_3628,N_3741);
and U4400 (N_4400,N_3205,N_3997);
or U4401 (N_4401,N_3914,N_3759);
or U4402 (N_4402,N_3406,N_3592);
xnor U4403 (N_4403,N_3935,N_3261);
or U4404 (N_4404,N_3016,N_3620);
or U4405 (N_4405,N_3372,N_3112);
or U4406 (N_4406,N_3118,N_3692);
nor U4407 (N_4407,N_3907,N_3899);
and U4408 (N_4408,N_3550,N_3127);
and U4409 (N_4409,N_3430,N_3611);
or U4410 (N_4410,N_3784,N_3185);
and U4411 (N_4411,N_3465,N_3259);
and U4412 (N_4412,N_3677,N_3448);
xnor U4413 (N_4413,N_3701,N_3808);
nor U4414 (N_4414,N_3064,N_3648);
nor U4415 (N_4415,N_3178,N_3497);
nand U4416 (N_4416,N_3305,N_3092);
nor U4417 (N_4417,N_3875,N_3654);
nor U4418 (N_4418,N_3436,N_3419);
and U4419 (N_4419,N_3103,N_3439);
nand U4420 (N_4420,N_3977,N_3706);
nor U4421 (N_4421,N_3152,N_3745);
or U4422 (N_4422,N_3747,N_3352);
nor U4423 (N_4423,N_3048,N_3590);
and U4424 (N_4424,N_3005,N_3141);
or U4425 (N_4425,N_3631,N_3812);
or U4426 (N_4426,N_3134,N_3336);
nand U4427 (N_4427,N_3951,N_3234);
nor U4428 (N_4428,N_3643,N_3377);
nor U4429 (N_4429,N_3405,N_3449);
and U4430 (N_4430,N_3093,N_3216);
or U4431 (N_4431,N_3971,N_3868);
or U4432 (N_4432,N_3557,N_3034);
or U4433 (N_4433,N_3787,N_3209);
nand U4434 (N_4434,N_3032,N_3203);
nand U4435 (N_4435,N_3410,N_3593);
nor U4436 (N_4436,N_3320,N_3573);
or U4437 (N_4437,N_3983,N_3632);
and U4438 (N_4438,N_3545,N_3081);
and U4439 (N_4439,N_3671,N_3509);
or U4440 (N_4440,N_3910,N_3044);
nor U4441 (N_4441,N_3160,N_3308);
or U4442 (N_4442,N_3036,N_3947);
and U4443 (N_4443,N_3440,N_3287);
or U4444 (N_4444,N_3255,N_3966);
nand U4445 (N_4445,N_3041,N_3346);
or U4446 (N_4446,N_3811,N_3399);
nor U4447 (N_4447,N_3341,N_3451);
or U4448 (N_4448,N_3714,N_3764);
or U4449 (N_4449,N_3792,N_3993);
nor U4450 (N_4450,N_3433,N_3461);
and U4451 (N_4451,N_3821,N_3481);
or U4452 (N_4452,N_3496,N_3429);
nand U4453 (N_4453,N_3199,N_3800);
or U4454 (N_4454,N_3012,N_3170);
nor U4455 (N_4455,N_3711,N_3420);
or U4456 (N_4456,N_3310,N_3657);
or U4457 (N_4457,N_3623,N_3350);
nand U4458 (N_4458,N_3476,N_3224);
or U4459 (N_4459,N_3785,N_3565);
and U4460 (N_4460,N_3901,N_3274);
nand U4461 (N_4461,N_3452,N_3518);
or U4462 (N_4462,N_3698,N_3146);
and U4463 (N_4463,N_3484,N_3615);
or U4464 (N_4464,N_3374,N_3612);
and U4465 (N_4465,N_3105,N_3850);
and U4466 (N_4466,N_3173,N_3860);
nor U4467 (N_4467,N_3303,N_3814);
and U4468 (N_4468,N_3075,N_3960);
nor U4469 (N_4469,N_3426,N_3201);
or U4470 (N_4470,N_3586,N_3124);
and U4471 (N_4471,N_3475,N_3902);
nor U4472 (N_4472,N_3155,N_3864);
and U4473 (N_4473,N_3571,N_3019);
or U4474 (N_4474,N_3156,N_3761);
nand U4475 (N_4475,N_3572,N_3068);
and U4476 (N_4476,N_3831,N_3442);
and U4477 (N_4477,N_3564,N_3125);
nand U4478 (N_4478,N_3403,N_3323);
or U4479 (N_4479,N_3670,N_3197);
nor U4480 (N_4480,N_3282,N_3342);
nand U4481 (N_4481,N_3113,N_3928);
and U4482 (N_4482,N_3585,N_3526);
nand U4483 (N_4483,N_3145,N_3809);
and U4484 (N_4484,N_3245,N_3895);
nor U4485 (N_4485,N_3371,N_3338);
nand U4486 (N_4486,N_3286,N_3619);
nor U4487 (N_4487,N_3933,N_3964);
and U4488 (N_4488,N_3834,N_3219);
and U4489 (N_4489,N_3724,N_3169);
and U4490 (N_4490,N_3389,N_3344);
or U4491 (N_4491,N_3531,N_3843);
nand U4492 (N_4492,N_3065,N_3647);
nor U4493 (N_4493,N_3153,N_3069);
nor U4494 (N_4494,N_3056,N_3740);
nor U4495 (N_4495,N_3602,N_3795);
nor U4496 (N_4496,N_3157,N_3646);
and U4497 (N_4497,N_3491,N_3292);
or U4498 (N_4498,N_3957,N_3822);
nand U4499 (N_4499,N_3464,N_3941);
nand U4500 (N_4500,N_3412,N_3816);
and U4501 (N_4501,N_3780,N_3622);
nand U4502 (N_4502,N_3072,N_3613);
nor U4503 (N_4503,N_3541,N_3133);
nor U4504 (N_4504,N_3267,N_3175);
nor U4505 (N_4505,N_3548,N_3604);
nand U4506 (N_4506,N_3320,N_3444);
nand U4507 (N_4507,N_3197,N_3734);
nand U4508 (N_4508,N_3510,N_3026);
nor U4509 (N_4509,N_3516,N_3648);
and U4510 (N_4510,N_3354,N_3023);
nor U4511 (N_4511,N_3862,N_3890);
nor U4512 (N_4512,N_3866,N_3615);
nor U4513 (N_4513,N_3548,N_3205);
or U4514 (N_4514,N_3398,N_3193);
and U4515 (N_4515,N_3933,N_3324);
or U4516 (N_4516,N_3934,N_3706);
or U4517 (N_4517,N_3392,N_3673);
nor U4518 (N_4518,N_3625,N_3065);
or U4519 (N_4519,N_3456,N_3515);
nand U4520 (N_4520,N_3849,N_3576);
and U4521 (N_4521,N_3469,N_3281);
and U4522 (N_4522,N_3136,N_3816);
or U4523 (N_4523,N_3422,N_3027);
or U4524 (N_4524,N_3215,N_3272);
and U4525 (N_4525,N_3291,N_3136);
nor U4526 (N_4526,N_3566,N_3049);
nor U4527 (N_4527,N_3033,N_3374);
nor U4528 (N_4528,N_3164,N_3944);
nor U4529 (N_4529,N_3173,N_3999);
and U4530 (N_4530,N_3463,N_3899);
or U4531 (N_4531,N_3792,N_3999);
and U4532 (N_4532,N_3859,N_3124);
and U4533 (N_4533,N_3081,N_3994);
or U4534 (N_4534,N_3948,N_3933);
nor U4535 (N_4535,N_3243,N_3460);
nor U4536 (N_4536,N_3183,N_3851);
nand U4537 (N_4537,N_3709,N_3990);
and U4538 (N_4538,N_3271,N_3813);
nand U4539 (N_4539,N_3086,N_3163);
and U4540 (N_4540,N_3678,N_3575);
or U4541 (N_4541,N_3755,N_3120);
or U4542 (N_4542,N_3914,N_3314);
or U4543 (N_4543,N_3646,N_3923);
or U4544 (N_4544,N_3908,N_3286);
or U4545 (N_4545,N_3306,N_3836);
nand U4546 (N_4546,N_3029,N_3922);
nor U4547 (N_4547,N_3174,N_3577);
nand U4548 (N_4548,N_3502,N_3035);
nand U4549 (N_4549,N_3137,N_3144);
and U4550 (N_4550,N_3009,N_3159);
and U4551 (N_4551,N_3687,N_3123);
and U4552 (N_4552,N_3256,N_3628);
nor U4553 (N_4553,N_3744,N_3707);
nor U4554 (N_4554,N_3124,N_3260);
nor U4555 (N_4555,N_3312,N_3020);
nand U4556 (N_4556,N_3339,N_3095);
nand U4557 (N_4557,N_3269,N_3466);
and U4558 (N_4558,N_3677,N_3484);
or U4559 (N_4559,N_3404,N_3668);
or U4560 (N_4560,N_3217,N_3072);
or U4561 (N_4561,N_3134,N_3988);
and U4562 (N_4562,N_3997,N_3003);
nor U4563 (N_4563,N_3134,N_3735);
and U4564 (N_4564,N_3512,N_3587);
and U4565 (N_4565,N_3850,N_3351);
nor U4566 (N_4566,N_3280,N_3707);
xor U4567 (N_4567,N_3282,N_3663);
or U4568 (N_4568,N_3833,N_3181);
nor U4569 (N_4569,N_3612,N_3253);
and U4570 (N_4570,N_3522,N_3263);
nand U4571 (N_4571,N_3208,N_3232);
and U4572 (N_4572,N_3581,N_3062);
nor U4573 (N_4573,N_3598,N_3559);
nand U4574 (N_4574,N_3132,N_3174);
nor U4575 (N_4575,N_3236,N_3747);
and U4576 (N_4576,N_3310,N_3134);
or U4577 (N_4577,N_3655,N_3709);
nand U4578 (N_4578,N_3627,N_3937);
nand U4579 (N_4579,N_3350,N_3008);
nand U4580 (N_4580,N_3533,N_3472);
or U4581 (N_4581,N_3564,N_3153);
or U4582 (N_4582,N_3117,N_3505);
and U4583 (N_4583,N_3363,N_3459);
or U4584 (N_4584,N_3577,N_3999);
nor U4585 (N_4585,N_3779,N_3253);
nand U4586 (N_4586,N_3316,N_3290);
nand U4587 (N_4587,N_3641,N_3440);
or U4588 (N_4588,N_3147,N_3680);
nand U4589 (N_4589,N_3992,N_3543);
nor U4590 (N_4590,N_3574,N_3472);
and U4591 (N_4591,N_3827,N_3477);
or U4592 (N_4592,N_3604,N_3417);
xnor U4593 (N_4593,N_3627,N_3661);
and U4594 (N_4594,N_3447,N_3584);
or U4595 (N_4595,N_3531,N_3155);
nor U4596 (N_4596,N_3291,N_3311);
and U4597 (N_4597,N_3538,N_3049);
and U4598 (N_4598,N_3169,N_3017);
nand U4599 (N_4599,N_3437,N_3461);
or U4600 (N_4600,N_3976,N_3735);
or U4601 (N_4601,N_3136,N_3988);
nor U4602 (N_4602,N_3984,N_3091);
nand U4603 (N_4603,N_3783,N_3096);
nand U4604 (N_4604,N_3143,N_3947);
or U4605 (N_4605,N_3334,N_3519);
nand U4606 (N_4606,N_3952,N_3934);
or U4607 (N_4607,N_3034,N_3259);
nor U4608 (N_4608,N_3632,N_3906);
or U4609 (N_4609,N_3698,N_3596);
and U4610 (N_4610,N_3564,N_3219);
nand U4611 (N_4611,N_3743,N_3069);
nand U4612 (N_4612,N_3213,N_3868);
and U4613 (N_4613,N_3832,N_3108);
nor U4614 (N_4614,N_3274,N_3599);
nand U4615 (N_4615,N_3543,N_3550);
and U4616 (N_4616,N_3643,N_3094);
or U4617 (N_4617,N_3992,N_3193);
nor U4618 (N_4618,N_3232,N_3429);
and U4619 (N_4619,N_3974,N_3999);
nand U4620 (N_4620,N_3995,N_3650);
or U4621 (N_4621,N_3968,N_3246);
nor U4622 (N_4622,N_3884,N_3753);
and U4623 (N_4623,N_3738,N_3319);
nor U4624 (N_4624,N_3726,N_3717);
or U4625 (N_4625,N_3890,N_3934);
nor U4626 (N_4626,N_3047,N_3363);
nor U4627 (N_4627,N_3434,N_3736);
or U4628 (N_4628,N_3921,N_3083);
nor U4629 (N_4629,N_3552,N_3061);
nand U4630 (N_4630,N_3370,N_3401);
or U4631 (N_4631,N_3956,N_3573);
or U4632 (N_4632,N_3566,N_3235);
nor U4633 (N_4633,N_3207,N_3161);
nor U4634 (N_4634,N_3820,N_3338);
nor U4635 (N_4635,N_3587,N_3615);
nor U4636 (N_4636,N_3292,N_3950);
nand U4637 (N_4637,N_3467,N_3815);
and U4638 (N_4638,N_3937,N_3779);
or U4639 (N_4639,N_3409,N_3130);
nor U4640 (N_4640,N_3241,N_3706);
or U4641 (N_4641,N_3240,N_3496);
or U4642 (N_4642,N_3330,N_3663);
xor U4643 (N_4643,N_3596,N_3609);
nor U4644 (N_4644,N_3260,N_3366);
nand U4645 (N_4645,N_3981,N_3627);
or U4646 (N_4646,N_3906,N_3707);
or U4647 (N_4647,N_3659,N_3108);
and U4648 (N_4648,N_3512,N_3963);
or U4649 (N_4649,N_3443,N_3387);
nand U4650 (N_4650,N_3522,N_3238);
and U4651 (N_4651,N_3266,N_3977);
nand U4652 (N_4652,N_3639,N_3069);
nor U4653 (N_4653,N_3292,N_3350);
and U4654 (N_4654,N_3727,N_3629);
nand U4655 (N_4655,N_3323,N_3956);
nor U4656 (N_4656,N_3723,N_3490);
and U4657 (N_4657,N_3133,N_3905);
nand U4658 (N_4658,N_3211,N_3471);
nor U4659 (N_4659,N_3022,N_3137);
and U4660 (N_4660,N_3903,N_3837);
and U4661 (N_4661,N_3170,N_3761);
nor U4662 (N_4662,N_3569,N_3087);
or U4663 (N_4663,N_3313,N_3051);
and U4664 (N_4664,N_3333,N_3662);
and U4665 (N_4665,N_3231,N_3563);
nor U4666 (N_4666,N_3939,N_3102);
nor U4667 (N_4667,N_3225,N_3698);
nand U4668 (N_4668,N_3808,N_3297);
and U4669 (N_4669,N_3393,N_3873);
nor U4670 (N_4670,N_3375,N_3100);
or U4671 (N_4671,N_3511,N_3918);
nor U4672 (N_4672,N_3907,N_3131);
nand U4673 (N_4673,N_3195,N_3389);
and U4674 (N_4674,N_3693,N_3252);
nand U4675 (N_4675,N_3050,N_3607);
or U4676 (N_4676,N_3193,N_3945);
nand U4677 (N_4677,N_3354,N_3500);
nand U4678 (N_4678,N_3873,N_3104);
nand U4679 (N_4679,N_3055,N_3810);
and U4680 (N_4680,N_3206,N_3663);
and U4681 (N_4681,N_3231,N_3591);
and U4682 (N_4682,N_3017,N_3041);
nor U4683 (N_4683,N_3989,N_3836);
nand U4684 (N_4684,N_3898,N_3310);
nor U4685 (N_4685,N_3532,N_3191);
nor U4686 (N_4686,N_3923,N_3408);
and U4687 (N_4687,N_3344,N_3763);
nand U4688 (N_4688,N_3059,N_3602);
or U4689 (N_4689,N_3884,N_3260);
nand U4690 (N_4690,N_3651,N_3405);
nor U4691 (N_4691,N_3884,N_3750);
or U4692 (N_4692,N_3854,N_3024);
and U4693 (N_4693,N_3643,N_3077);
and U4694 (N_4694,N_3743,N_3349);
and U4695 (N_4695,N_3033,N_3541);
nor U4696 (N_4696,N_3969,N_3161);
nor U4697 (N_4697,N_3136,N_3447);
and U4698 (N_4698,N_3374,N_3540);
or U4699 (N_4699,N_3205,N_3731);
nand U4700 (N_4700,N_3693,N_3681);
and U4701 (N_4701,N_3036,N_3355);
nand U4702 (N_4702,N_3755,N_3475);
and U4703 (N_4703,N_3218,N_3248);
nand U4704 (N_4704,N_3173,N_3127);
nand U4705 (N_4705,N_3495,N_3618);
and U4706 (N_4706,N_3737,N_3531);
nor U4707 (N_4707,N_3733,N_3562);
nand U4708 (N_4708,N_3517,N_3271);
and U4709 (N_4709,N_3876,N_3356);
nand U4710 (N_4710,N_3646,N_3302);
or U4711 (N_4711,N_3052,N_3826);
or U4712 (N_4712,N_3509,N_3534);
nor U4713 (N_4713,N_3606,N_3694);
or U4714 (N_4714,N_3392,N_3642);
or U4715 (N_4715,N_3831,N_3906);
or U4716 (N_4716,N_3628,N_3057);
nand U4717 (N_4717,N_3418,N_3128);
nand U4718 (N_4718,N_3793,N_3765);
and U4719 (N_4719,N_3811,N_3571);
and U4720 (N_4720,N_3342,N_3042);
nor U4721 (N_4721,N_3027,N_3663);
and U4722 (N_4722,N_3802,N_3012);
or U4723 (N_4723,N_3185,N_3178);
nand U4724 (N_4724,N_3694,N_3215);
and U4725 (N_4725,N_3838,N_3819);
or U4726 (N_4726,N_3419,N_3078);
nand U4727 (N_4727,N_3402,N_3031);
nor U4728 (N_4728,N_3547,N_3356);
xor U4729 (N_4729,N_3877,N_3802);
nand U4730 (N_4730,N_3207,N_3649);
nand U4731 (N_4731,N_3004,N_3866);
or U4732 (N_4732,N_3437,N_3082);
nor U4733 (N_4733,N_3183,N_3548);
and U4734 (N_4734,N_3041,N_3774);
nor U4735 (N_4735,N_3812,N_3313);
or U4736 (N_4736,N_3664,N_3946);
or U4737 (N_4737,N_3746,N_3144);
nor U4738 (N_4738,N_3858,N_3397);
nand U4739 (N_4739,N_3035,N_3182);
or U4740 (N_4740,N_3472,N_3074);
and U4741 (N_4741,N_3123,N_3448);
xnor U4742 (N_4742,N_3339,N_3667);
or U4743 (N_4743,N_3232,N_3871);
nor U4744 (N_4744,N_3301,N_3781);
and U4745 (N_4745,N_3256,N_3544);
nand U4746 (N_4746,N_3789,N_3327);
and U4747 (N_4747,N_3378,N_3599);
or U4748 (N_4748,N_3633,N_3245);
or U4749 (N_4749,N_3739,N_3553);
and U4750 (N_4750,N_3194,N_3736);
nor U4751 (N_4751,N_3854,N_3400);
nand U4752 (N_4752,N_3542,N_3055);
and U4753 (N_4753,N_3263,N_3124);
or U4754 (N_4754,N_3812,N_3471);
nand U4755 (N_4755,N_3404,N_3053);
nand U4756 (N_4756,N_3021,N_3800);
and U4757 (N_4757,N_3336,N_3287);
nor U4758 (N_4758,N_3597,N_3384);
nor U4759 (N_4759,N_3981,N_3463);
nor U4760 (N_4760,N_3132,N_3588);
nor U4761 (N_4761,N_3487,N_3907);
nand U4762 (N_4762,N_3534,N_3380);
or U4763 (N_4763,N_3441,N_3715);
nor U4764 (N_4764,N_3103,N_3912);
nand U4765 (N_4765,N_3124,N_3413);
nand U4766 (N_4766,N_3587,N_3088);
nor U4767 (N_4767,N_3873,N_3059);
nand U4768 (N_4768,N_3687,N_3770);
nand U4769 (N_4769,N_3611,N_3346);
nand U4770 (N_4770,N_3858,N_3708);
and U4771 (N_4771,N_3611,N_3037);
nand U4772 (N_4772,N_3225,N_3207);
nand U4773 (N_4773,N_3601,N_3478);
or U4774 (N_4774,N_3888,N_3998);
and U4775 (N_4775,N_3196,N_3644);
or U4776 (N_4776,N_3850,N_3752);
nand U4777 (N_4777,N_3387,N_3424);
and U4778 (N_4778,N_3061,N_3172);
and U4779 (N_4779,N_3612,N_3854);
nor U4780 (N_4780,N_3380,N_3703);
nand U4781 (N_4781,N_3125,N_3879);
nand U4782 (N_4782,N_3613,N_3773);
and U4783 (N_4783,N_3884,N_3550);
nor U4784 (N_4784,N_3163,N_3469);
or U4785 (N_4785,N_3640,N_3674);
nand U4786 (N_4786,N_3033,N_3830);
and U4787 (N_4787,N_3207,N_3972);
nand U4788 (N_4788,N_3443,N_3085);
nand U4789 (N_4789,N_3614,N_3424);
nand U4790 (N_4790,N_3389,N_3595);
nor U4791 (N_4791,N_3657,N_3955);
nand U4792 (N_4792,N_3845,N_3022);
nand U4793 (N_4793,N_3881,N_3902);
nor U4794 (N_4794,N_3681,N_3846);
or U4795 (N_4795,N_3327,N_3988);
and U4796 (N_4796,N_3725,N_3818);
nor U4797 (N_4797,N_3377,N_3504);
nand U4798 (N_4798,N_3596,N_3365);
xor U4799 (N_4799,N_3233,N_3132);
and U4800 (N_4800,N_3554,N_3778);
nor U4801 (N_4801,N_3294,N_3955);
nand U4802 (N_4802,N_3760,N_3291);
nor U4803 (N_4803,N_3938,N_3445);
nor U4804 (N_4804,N_3594,N_3330);
nor U4805 (N_4805,N_3557,N_3430);
xnor U4806 (N_4806,N_3457,N_3949);
nand U4807 (N_4807,N_3987,N_3520);
nor U4808 (N_4808,N_3875,N_3283);
or U4809 (N_4809,N_3189,N_3150);
nand U4810 (N_4810,N_3273,N_3530);
nand U4811 (N_4811,N_3600,N_3722);
nor U4812 (N_4812,N_3611,N_3229);
xnor U4813 (N_4813,N_3443,N_3919);
and U4814 (N_4814,N_3416,N_3359);
nor U4815 (N_4815,N_3173,N_3176);
or U4816 (N_4816,N_3758,N_3261);
and U4817 (N_4817,N_3250,N_3131);
nor U4818 (N_4818,N_3574,N_3092);
nand U4819 (N_4819,N_3372,N_3214);
nor U4820 (N_4820,N_3889,N_3102);
or U4821 (N_4821,N_3480,N_3456);
nor U4822 (N_4822,N_3137,N_3586);
nand U4823 (N_4823,N_3716,N_3411);
nor U4824 (N_4824,N_3682,N_3397);
nor U4825 (N_4825,N_3846,N_3859);
nor U4826 (N_4826,N_3509,N_3682);
or U4827 (N_4827,N_3971,N_3216);
nand U4828 (N_4828,N_3473,N_3954);
nand U4829 (N_4829,N_3304,N_3020);
and U4830 (N_4830,N_3051,N_3266);
or U4831 (N_4831,N_3024,N_3088);
nor U4832 (N_4832,N_3620,N_3823);
nand U4833 (N_4833,N_3382,N_3959);
and U4834 (N_4834,N_3624,N_3050);
nand U4835 (N_4835,N_3886,N_3255);
or U4836 (N_4836,N_3071,N_3964);
and U4837 (N_4837,N_3032,N_3904);
nand U4838 (N_4838,N_3910,N_3128);
and U4839 (N_4839,N_3829,N_3983);
nor U4840 (N_4840,N_3200,N_3158);
nand U4841 (N_4841,N_3637,N_3833);
or U4842 (N_4842,N_3620,N_3921);
or U4843 (N_4843,N_3342,N_3702);
nor U4844 (N_4844,N_3520,N_3039);
nand U4845 (N_4845,N_3810,N_3405);
and U4846 (N_4846,N_3223,N_3514);
nand U4847 (N_4847,N_3111,N_3852);
or U4848 (N_4848,N_3535,N_3886);
nand U4849 (N_4849,N_3310,N_3342);
or U4850 (N_4850,N_3273,N_3269);
and U4851 (N_4851,N_3447,N_3484);
nand U4852 (N_4852,N_3680,N_3454);
nor U4853 (N_4853,N_3856,N_3987);
or U4854 (N_4854,N_3726,N_3351);
or U4855 (N_4855,N_3459,N_3243);
or U4856 (N_4856,N_3066,N_3409);
or U4857 (N_4857,N_3624,N_3101);
and U4858 (N_4858,N_3672,N_3971);
or U4859 (N_4859,N_3153,N_3855);
or U4860 (N_4860,N_3797,N_3034);
and U4861 (N_4861,N_3809,N_3691);
or U4862 (N_4862,N_3689,N_3916);
nand U4863 (N_4863,N_3743,N_3715);
nand U4864 (N_4864,N_3271,N_3012);
and U4865 (N_4865,N_3735,N_3433);
or U4866 (N_4866,N_3269,N_3973);
nor U4867 (N_4867,N_3382,N_3738);
nand U4868 (N_4868,N_3930,N_3826);
nor U4869 (N_4869,N_3422,N_3187);
or U4870 (N_4870,N_3343,N_3387);
or U4871 (N_4871,N_3702,N_3399);
and U4872 (N_4872,N_3147,N_3341);
or U4873 (N_4873,N_3677,N_3511);
nand U4874 (N_4874,N_3450,N_3183);
nand U4875 (N_4875,N_3113,N_3340);
nand U4876 (N_4876,N_3368,N_3057);
and U4877 (N_4877,N_3649,N_3252);
and U4878 (N_4878,N_3544,N_3903);
nand U4879 (N_4879,N_3900,N_3406);
nand U4880 (N_4880,N_3108,N_3295);
nand U4881 (N_4881,N_3157,N_3748);
nand U4882 (N_4882,N_3648,N_3677);
or U4883 (N_4883,N_3131,N_3277);
and U4884 (N_4884,N_3817,N_3714);
or U4885 (N_4885,N_3091,N_3592);
and U4886 (N_4886,N_3106,N_3705);
and U4887 (N_4887,N_3345,N_3106);
nand U4888 (N_4888,N_3945,N_3153);
nor U4889 (N_4889,N_3873,N_3620);
or U4890 (N_4890,N_3991,N_3142);
or U4891 (N_4891,N_3761,N_3172);
nor U4892 (N_4892,N_3287,N_3180);
nor U4893 (N_4893,N_3079,N_3795);
or U4894 (N_4894,N_3973,N_3116);
or U4895 (N_4895,N_3813,N_3450);
or U4896 (N_4896,N_3151,N_3424);
nor U4897 (N_4897,N_3005,N_3506);
nor U4898 (N_4898,N_3383,N_3747);
nand U4899 (N_4899,N_3874,N_3698);
and U4900 (N_4900,N_3350,N_3386);
and U4901 (N_4901,N_3762,N_3842);
nor U4902 (N_4902,N_3540,N_3761);
nand U4903 (N_4903,N_3471,N_3487);
nor U4904 (N_4904,N_3576,N_3648);
nor U4905 (N_4905,N_3370,N_3158);
nor U4906 (N_4906,N_3027,N_3327);
nor U4907 (N_4907,N_3572,N_3909);
nand U4908 (N_4908,N_3609,N_3223);
or U4909 (N_4909,N_3595,N_3723);
nand U4910 (N_4910,N_3654,N_3140);
and U4911 (N_4911,N_3432,N_3196);
or U4912 (N_4912,N_3631,N_3888);
and U4913 (N_4913,N_3764,N_3439);
and U4914 (N_4914,N_3144,N_3658);
or U4915 (N_4915,N_3214,N_3554);
and U4916 (N_4916,N_3239,N_3391);
nand U4917 (N_4917,N_3522,N_3448);
and U4918 (N_4918,N_3710,N_3204);
nand U4919 (N_4919,N_3193,N_3817);
or U4920 (N_4920,N_3069,N_3517);
nor U4921 (N_4921,N_3548,N_3294);
and U4922 (N_4922,N_3909,N_3652);
nand U4923 (N_4923,N_3402,N_3910);
or U4924 (N_4924,N_3267,N_3752);
and U4925 (N_4925,N_3595,N_3850);
nor U4926 (N_4926,N_3285,N_3746);
nor U4927 (N_4927,N_3740,N_3892);
nand U4928 (N_4928,N_3361,N_3825);
or U4929 (N_4929,N_3564,N_3739);
nand U4930 (N_4930,N_3920,N_3439);
and U4931 (N_4931,N_3134,N_3614);
nor U4932 (N_4932,N_3232,N_3958);
nand U4933 (N_4933,N_3049,N_3379);
or U4934 (N_4934,N_3459,N_3851);
nand U4935 (N_4935,N_3569,N_3118);
nor U4936 (N_4936,N_3542,N_3983);
nor U4937 (N_4937,N_3972,N_3895);
nand U4938 (N_4938,N_3241,N_3696);
nor U4939 (N_4939,N_3050,N_3022);
and U4940 (N_4940,N_3648,N_3980);
or U4941 (N_4941,N_3149,N_3860);
or U4942 (N_4942,N_3802,N_3133);
nand U4943 (N_4943,N_3941,N_3168);
or U4944 (N_4944,N_3068,N_3841);
nor U4945 (N_4945,N_3491,N_3999);
nor U4946 (N_4946,N_3052,N_3717);
and U4947 (N_4947,N_3679,N_3838);
nand U4948 (N_4948,N_3644,N_3945);
nor U4949 (N_4949,N_3083,N_3606);
nand U4950 (N_4950,N_3143,N_3700);
and U4951 (N_4951,N_3709,N_3516);
nand U4952 (N_4952,N_3672,N_3886);
nand U4953 (N_4953,N_3749,N_3956);
and U4954 (N_4954,N_3846,N_3590);
and U4955 (N_4955,N_3508,N_3698);
nor U4956 (N_4956,N_3062,N_3662);
xnor U4957 (N_4957,N_3813,N_3840);
nand U4958 (N_4958,N_3591,N_3894);
or U4959 (N_4959,N_3805,N_3860);
or U4960 (N_4960,N_3638,N_3401);
nand U4961 (N_4961,N_3631,N_3526);
and U4962 (N_4962,N_3840,N_3514);
and U4963 (N_4963,N_3452,N_3040);
nor U4964 (N_4964,N_3847,N_3144);
and U4965 (N_4965,N_3374,N_3943);
nor U4966 (N_4966,N_3669,N_3287);
or U4967 (N_4967,N_3980,N_3081);
nor U4968 (N_4968,N_3055,N_3669);
and U4969 (N_4969,N_3735,N_3654);
nand U4970 (N_4970,N_3328,N_3908);
and U4971 (N_4971,N_3943,N_3826);
and U4972 (N_4972,N_3454,N_3091);
nand U4973 (N_4973,N_3211,N_3116);
or U4974 (N_4974,N_3657,N_3290);
or U4975 (N_4975,N_3070,N_3787);
nand U4976 (N_4976,N_3201,N_3322);
nor U4977 (N_4977,N_3070,N_3170);
nand U4978 (N_4978,N_3539,N_3427);
or U4979 (N_4979,N_3816,N_3876);
nand U4980 (N_4980,N_3170,N_3026);
nand U4981 (N_4981,N_3353,N_3346);
nand U4982 (N_4982,N_3516,N_3851);
nand U4983 (N_4983,N_3345,N_3621);
nand U4984 (N_4984,N_3017,N_3539);
nor U4985 (N_4985,N_3356,N_3312);
or U4986 (N_4986,N_3566,N_3575);
and U4987 (N_4987,N_3832,N_3506);
nor U4988 (N_4988,N_3969,N_3514);
and U4989 (N_4989,N_3620,N_3673);
or U4990 (N_4990,N_3193,N_3164);
nor U4991 (N_4991,N_3686,N_3547);
and U4992 (N_4992,N_3191,N_3282);
and U4993 (N_4993,N_3208,N_3202);
or U4994 (N_4994,N_3268,N_3518);
and U4995 (N_4995,N_3473,N_3601);
and U4996 (N_4996,N_3159,N_3785);
and U4997 (N_4997,N_3156,N_3567);
and U4998 (N_4998,N_3706,N_3198);
or U4999 (N_4999,N_3778,N_3826);
or UO_0 (O_0,N_4073,N_4704);
nand UO_1 (O_1,N_4927,N_4948);
or UO_2 (O_2,N_4468,N_4110);
nand UO_3 (O_3,N_4973,N_4819);
nand UO_4 (O_4,N_4232,N_4109);
nor UO_5 (O_5,N_4604,N_4367);
and UO_6 (O_6,N_4955,N_4675);
and UO_7 (O_7,N_4561,N_4104);
xnor UO_8 (O_8,N_4556,N_4080);
or UO_9 (O_9,N_4686,N_4546);
nor UO_10 (O_10,N_4303,N_4473);
and UO_11 (O_11,N_4424,N_4606);
or UO_12 (O_12,N_4373,N_4240);
nand UO_13 (O_13,N_4289,N_4952);
nor UO_14 (O_14,N_4827,N_4551);
or UO_15 (O_15,N_4800,N_4278);
and UO_16 (O_16,N_4884,N_4145);
and UO_17 (O_17,N_4463,N_4993);
nand UO_18 (O_18,N_4084,N_4797);
and UO_19 (O_19,N_4245,N_4485);
nand UO_20 (O_20,N_4881,N_4703);
nand UO_21 (O_21,N_4255,N_4740);
nor UO_22 (O_22,N_4030,N_4777);
nor UO_23 (O_23,N_4879,N_4862);
nor UO_24 (O_24,N_4090,N_4869);
nand UO_25 (O_25,N_4527,N_4118);
and UO_26 (O_26,N_4630,N_4048);
nand UO_27 (O_27,N_4554,N_4286);
or UO_28 (O_28,N_4691,N_4706);
nand UO_29 (O_29,N_4587,N_4886);
and UO_30 (O_30,N_4978,N_4380);
or UO_31 (O_31,N_4455,N_4078);
nand UO_32 (O_32,N_4493,N_4935);
and UO_33 (O_33,N_4169,N_4997);
nor UO_34 (O_34,N_4023,N_4020);
nor UO_35 (O_35,N_4343,N_4887);
or UO_36 (O_36,N_4427,N_4735);
and UO_37 (O_37,N_4235,N_4496);
nor UO_38 (O_38,N_4435,N_4847);
and UO_39 (O_39,N_4051,N_4059);
or UO_40 (O_40,N_4697,N_4752);
nand UO_41 (O_41,N_4215,N_4433);
and UO_42 (O_42,N_4345,N_4316);
and UO_43 (O_43,N_4195,N_4888);
nor UO_44 (O_44,N_4419,N_4854);
nand UO_45 (O_45,N_4996,N_4041);
or UO_46 (O_46,N_4189,N_4470);
nand UO_47 (O_47,N_4197,N_4635);
or UO_48 (O_48,N_4368,N_4313);
nor UO_49 (O_49,N_4115,N_4812);
and UO_50 (O_50,N_4096,N_4641);
nor UO_51 (O_51,N_4001,N_4160);
nand UO_52 (O_52,N_4707,N_4113);
and UO_53 (O_53,N_4227,N_4206);
nand UO_54 (O_54,N_4829,N_4762);
and UO_55 (O_55,N_4487,N_4922);
and UO_56 (O_56,N_4179,N_4914);
or UO_57 (O_57,N_4272,N_4324);
nand UO_58 (O_58,N_4678,N_4399);
nand UO_59 (O_59,N_4773,N_4045);
xnor UO_60 (O_60,N_4052,N_4792);
or UO_61 (O_61,N_4295,N_4397);
or UO_62 (O_62,N_4639,N_4943);
or UO_63 (O_63,N_4103,N_4122);
nor UO_64 (O_64,N_4055,N_4186);
and UO_65 (O_65,N_4178,N_4437);
nand UO_66 (O_66,N_4867,N_4076);
and UO_67 (O_67,N_4285,N_4002);
and UO_68 (O_68,N_4834,N_4067);
nor UO_69 (O_69,N_4921,N_4564);
or UO_70 (O_70,N_4199,N_4765);
nand UO_71 (O_71,N_4065,N_4168);
nor UO_72 (O_72,N_4591,N_4550);
or UO_73 (O_73,N_4007,N_4226);
or UO_74 (O_74,N_4649,N_4726);
nor UO_75 (O_75,N_4476,N_4071);
nand UO_76 (O_76,N_4617,N_4269);
or UO_77 (O_77,N_4183,N_4790);
nor UO_78 (O_78,N_4489,N_4063);
nand UO_79 (O_79,N_4018,N_4687);
nand UO_80 (O_80,N_4991,N_4577);
nand UO_81 (O_81,N_4840,N_4263);
or UO_82 (O_82,N_4594,N_4481);
nand UO_83 (O_83,N_4456,N_4393);
nand UO_84 (O_84,N_4961,N_4028);
nand UO_85 (O_85,N_4770,N_4552);
or UO_86 (O_86,N_4369,N_4563);
and UO_87 (O_87,N_4631,N_4816);
nand UO_88 (O_88,N_4629,N_4776);
or UO_89 (O_89,N_4513,N_4628);
or UO_90 (O_90,N_4663,N_4739);
and UO_91 (O_91,N_4533,N_4259);
and UO_92 (O_92,N_4971,N_4166);
and UO_93 (O_93,N_4785,N_4287);
nor UO_94 (O_94,N_4849,N_4781);
nand UO_95 (O_95,N_4085,N_4037);
and UO_96 (O_96,N_4842,N_4448);
and UO_97 (O_97,N_4086,N_4190);
nand UO_98 (O_98,N_4129,N_4667);
or UO_99 (O_99,N_4909,N_4980);
nand UO_100 (O_100,N_4831,N_4690);
and UO_101 (O_101,N_4852,N_4446);
or UO_102 (O_102,N_4817,N_4321);
and UO_103 (O_103,N_4810,N_4549);
nor UO_104 (O_104,N_4696,N_4214);
nand UO_105 (O_105,N_4748,N_4256);
nor UO_106 (O_106,N_4772,N_4273);
or UO_107 (O_107,N_4242,N_4469);
or UO_108 (O_108,N_4216,N_4536);
nand UO_109 (O_109,N_4276,N_4264);
or UO_110 (O_110,N_4353,N_4746);
and UO_111 (O_111,N_4106,N_4046);
nor UO_112 (O_112,N_4344,N_4454);
or UO_113 (O_113,N_4681,N_4260);
nor UO_114 (O_114,N_4648,N_4265);
nand UO_115 (O_115,N_4778,N_4389);
nor UO_116 (O_116,N_4666,N_4652);
and UO_117 (O_117,N_4580,N_4135);
and UO_118 (O_118,N_4172,N_4569);
nand UO_119 (O_119,N_4504,N_4105);
nor UO_120 (O_120,N_4205,N_4782);
and UO_121 (O_121,N_4501,N_4234);
and UO_122 (O_122,N_4458,N_4310);
nor UO_123 (O_123,N_4593,N_4089);
or UO_124 (O_124,N_4679,N_4671);
and UO_125 (O_125,N_4848,N_4567);
and UO_126 (O_126,N_4358,N_4668);
nor UO_127 (O_127,N_4420,N_4855);
nand UO_128 (O_128,N_4725,N_4412);
nor UO_129 (O_129,N_4656,N_4281);
nor UO_130 (O_130,N_4486,N_4787);
or UO_131 (O_131,N_4522,N_4669);
nand UO_132 (O_132,N_4994,N_4568);
or UO_133 (O_133,N_4043,N_4645);
nand UO_134 (O_134,N_4116,N_4676);
nor UO_135 (O_135,N_4429,N_4820);
and UO_136 (O_136,N_4187,N_4144);
and UO_137 (O_137,N_4282,N_4119);
nor UO_138 (O_138,N_4941,N_4066);
or UO_139 (O_139,N_4572,N_4155);
or UO_140 (O_140,N_4795,N_4123);
nand UO_141 (O_141,N_4574,N_4545);
and UO_142 (O_142,N_4062,N_4117);
or UO_143 (O_143,N_4813,N_4444);
nand UO_144 (O_144,N_4699,N_4526);
or UO_145 (O_145,N_4516,N_4718);
and UO_146 (O_146,N_4225,N_4127);
nand UO_147 (O_147,N_4902,N_4992);
nor UO_148 (O_148,N_4284,N_4844);
nor UO_149 (O_149,N_4490,N_4379);
or UO_150 (O_150,N_4859,N_4356);
nor UO_151 (O_151,N_4025,N_4908);
nand UO_152 (O_152,N_4453,N_4893);
and UO_153 (O_153,N_4158,N_4870);
or UO_154 (O_154,N_4904,N_4530);
nor UO_155 (O_155,N_4478,N_4767);
or UO_156 (O_156,N_4670,N_4161);
nand UO_157 (O_157,N_4081,N_4965);
and UO_158 (O_158,N_4911,N_4388);
or UO_159 (O_159,N_4708,N_4715);
or UO_160 (O_160,N_4452,N_4154);
or UO_161 (O_161,N_4775,N_4839);
or UO_162 (O_162,N_4900,N_4700);
nand UO_163 (O_163,N_4713,N_4638);
and UO_164 (O_164,N_4163,N_4498);
and UO_165 (O_165,N_4769,N_4520);
nand UO_166 (O_166,N_4222,N_4053);
and UO_167 (O_167,N_4985,N_4822);
nor UO_168 (O_168,N_4966,N_4525);
or UO_169 (O_169,N_4714,N_4874);
or UO_170 (O_170,N_4944,N_4381);
and UO_171 (O_171,N_4026,N_4083);
or UO_172 (O_172,N_4883,N_4658);
or UO_173 (O_173,N_4180,N_4885);
and UO_174 (O_174,N_4609,N_4832);
or UO_175 (O_175,N_4413,N_4040);
nand UO_176 (O_176,N_4302,N_4061);
nor UO_177 (O_177,N_4916,N_4167);
nand UO_178 (O_178,N_4695,N_4934);
nand UO_179 (O_179,N_4586,N_4531);
nor UO_180 (O_180,N_4688,N_4384);
or UO_181 (O_181,N_4833,N_4139);
and UO_182 (O_182,N_4625,N_4624);
and UO_183 (O_183,N_4120,N_4529);
nor UO_184 (O_184,N_4014,N_4091);
nand UO_185 (O_185,N_4156,N_4352);
and UO_186 (O_186,N_4431,N_4494);
nor UO_187 (O_187,N_4951,N_4508);
or UO_188 (O_188,N_4712,N_4818);
and UO_189 (O_189,N_4005,N_4464);
or UO_190 (O_190,N_4644,N_4406);
and UO_191 (O_191,N_4434,N_4836);
nand UO_192 (O_192,N_4796,N_4989);
and UO_193 (O_193,N_4191,N_4212);
or UO_194 (O_194,N_4990,N_4512);
nor UO_195 (O_195,N_4217,N_4233);
nor UO_196 (O_196,N_4607,N_4003);
nor UO_197 (O_197,N_4202,N_4684);
and UO_198 (O_198,N_4336,N_4049);
or UO_199 (O_199,N_4376,N_4643);
nand UO_200 (O_200,N_4959,N_4064);
xnor UO_201 (O_201,N_4890,N_4837);
or UO_202 (O_202,N_4148,N_4573);
nand UO_203 (O_203,N_4432,N_4857);
or UO_204 (O_204,N_4804,N_4791);
nand UO_205 (O_205,N_4057,N_4069);
nand UO_206 (O_206,N_4541,N_4540);
and UO_207 (O_207,N_4403,N_4502);
and UO_208 (O_208,N_4779,N_4015);
xnor UO_209 (O_209,N_4537,N_4034);
nor UO_210 (O_210,N_4876,N_4974);
or UO_211 (O_211,N_4351,N_4590);
nor UO_212 (O_212,N_4266,N_4548);
or UO_213 (O_213,N_4618,N_4484);
nor UO_214 (O_214,N_4111,N_4764);
or UO_215 (O_215,N_4292,N_4471);
nand UO_216 (O_216,N_4728,N_4661);
nor UO_217 (O_217,N_4450,N_4672);
and UO_218 (O_218,N_4133,N_4954);
nand UO_219 (O_219,N_4070,N_4491);
nand UO_220 (O_220,N_4280,N_4042);
nand UO_221 (O_221,N_4185,N_4000);
and UO_222 (O_222,N_4237,N_4325);
and UO_223 (O_223,N_4983,N_4438);
and UO_224 (O_224,N_4756,N_4760);
nor UO_225 (O_225,N_4755,N_4315);
nor UO_226 (O_226,N_4290,N_4033);
nor UO_227 (O_227,N_4171,N_4605);
and UO_228 (O_228,N_4979,N_4632);
and UO_229 (O_229,N_4142,N_4004);
and UO_230 (O_230,N_4655,N_4747);
and UO_231 (O_231,N_4309,N_4087);
nor UO_232 (O_232,N_4447,N_4017);
nand UO_233 (O_233,N_4132,N_4360);
or UO_234 (O_234,N_4730,N_4753);
and UO_235 (O_235,N_4441,N_4924);
nor UO_236 (O_236,N_4022,N_4794);
and UO_237 (O_237,N_4860,N_4068);
nor UO_238 (O_238,N_4864,N_4114);
and UO_239 (O_239,N_4333,N_4986);
nand UO_240 (O_240,N_4738,N_4174);
or UO_241 (O_241,N_4340,N_4268);
nand UO_242 (O_242,N_4600,N_4421);
nand UO_243 (O_243,N_4032,N_4492);
nor UO_244 (O_244,N_4724,N_4058);
nor UO_245 (O_245,N_4578,N_4535);
nand UO_246 (O_246,N_4377,N_4505);
nand UO_247 (O_247,N_4200,N_4694);
or UO_248 (O_248,N_4633,N_4056);
and UO_249 (O_249,N_4339,N_4942);
nor UO_250 (O_250,N_4383,N_4938);
nand UO_251 (O_251,N_4466,N_4560);
nand UO_252 (O_252,N_4400,N_4248);
nor UO_253 (O_253,N_4627,N_4774);
nand UO_254 (O_254,N_4024,N_4611);
nor UO_255 (O_255,N_4251,N_4683);
or UO_256 (O_256,N_4210,N_4363);
nand UO_257 (O_257,N_4912,N_4319);
nand UO_258 (O_258,N_4244,N_4744);
and UO_259 (O_259,N_4194,N_4228);
or UO_260 (O_260,N_4723,N_4647);
and UO_261 (O_261,N_4398,N_4653);
or UO_262 (O_262,N_4899,N_4897);
and UO_263 (O_263,N_4873,N_4177);
and UO_264 (O_264,N_4737,N_4483);
or UO_265 (O_265,N_4291,N_4461);
or UO_266 (O_266,N_4945,N_4918);
and UO_267 (O_267,N_4330,N_4112);
nor UO_268 (O_268,N_4875,N_4386);
nor UO_269 (O_269,N_4326,N_4359);
nor UO_270 (O_270,N_4761,N_4962);
nand UO_271 (O_271,N_4300,N_4253);
and UO_272 (O_272,N_4121,N_4603);
and UO_273 (O_273,N_4987,N_4793);
and UO_274 (O_274,N_4824,N_4650);
and UO_275 (O_275,N_4298,N_4246);
nand UO_276 (O_276,N_4141,N_4385);
or UO_277 (O_277,N_4662,N_4134);
and UO_278 (O_278,N_4750,N_4998);
nand UO_279 (O_279,N_4592,N_4868);
nor UO_280 (O_280,N_4387,N_4571);
or UO_281 (O_281,N_4125,N_4620);
and UO_282 (O_282,N_4510,N_4830);
nor UO_283 (O_283,N_4249,N_4414);
or UO_284 (O_284,N_4673,N_4853);
or UO_285 (O_285,N_4659,N_4338);
or UO_286 (O_286,N_4254,N_4891);
nand UO_287 (O_287,N_4108,N_4329);
nor UO_288 (O_288,N_4660,N_4674);
nand UO_289 (O_289,N_4162,N_4152);
nor UO_290 (O_290,N_4277,N_4140);
and UO_291 (O_291,N_4920,N_4150);
or UO_292 (O_292,N_4093,N_4882);
or UO_293 (O_293,N_4188,N_4733);
and UO_294 (O_294,N_4229,N_4518);
nand UO_295 (O_295,N_4362,N_4100);
and UO_296 (O_296,N_4601,N_4449);
nand UO_297 (O_297,N_4126,N_4936);
nor UO_298 (O_298,N_4239,N_4404);
nand UO_299 (O_299,N_4841,N_4088);
nor UO_300 (O_300,N_4274,N_4534);
nand UO_301 (O_301,N_4247,N_4223);
and UO_302 (O_302,N_4759,N_4230);
or UO_303 (O_303,N_4497,N_4612);
or UO_304 (O_304,N_4371,N_4375);
nor UO_305 (O_305,N_4192,N_4895);
and UO_306 (O_306,N_4843,N_4008);
nor UO_307 (O_307,N_4743,N_4422);
and UO_308 (O_308,N_4415,N_4558);
nand UO_309 (O_309,N_4271,N_4072);
or UO_310 (O_310,N_4250,N_4408);
nor UO_311 (O_311,N_4465,N_4858);
and UO_312 (O_312,N_4511,N_4950);
nor UO_313 (O_313,N_4296,N_4425);
or UO_314 (O_314,N_4780,N_4270);
nor UO_315 (O_315,N_4995,N_4917);
and UO_316 (O_316,N_4850,N_4693);
nor UO_317 (O_317,N_4811,N_4621);
or UO_318 (O_318,N_4401,N_4238);
and UO_319 (O_319,N_4975,N_4809);
nor UO_320 (O_320,N_4288,N_4877);
nand UO_321 (O_321,N_4430,N_4705);
nor UO_322 (O_322,N_4582,N_4933);
nor UO_323 (O_323,N_4038,N_4392);
nor UO_324 (O_324,N_4814,N_4821);
nand UO_325 (O_325,N_4521,N_4613);
nor UO_326 (O_326,N_4374,N_4736);
and UO_327 (O_327,N_4823,N_4299);
nor UO_328 (O_328,N_4312,N_4405);
nand UO_329 (O_329,N_4354,N_4749);
and UO_330 (O_330,N_4682,N_4539);
nor UO_331 (O_331,N_4306,N_4349);
nand UO_332 (O_332,N_4588,N_4204);
nand UO_333 (O_333,N_4929,N_4532);
nor UO_334 (O_334,N_4872,N_4193);
and UO_335 (O_335,N_4981,N_4845);
or UO_336 (O_336,N_4846,N_4283);
and UO_337 (O_337,N_4006,N_4826);
or UO_338 (O_338,N_4337,N_4634);
nor UO_339 (O_339,N_4716,N_4459);
nand UO_340 (O_340,N_4626,N_4495);
nand UO_341 (O_341,N_4013,N_4953);
or UO_342 (O_342,N_4925,N_4970);
nand UO_343 (O_343,N_4758,N_4428);
nor UO_344 (O_344,N_4865,N_4598);
nor UO_345 (O_345,N_4440,N_4642);
or UO_346 (O_346,N_4153,N_4131);
nor UO_347 (O_347,N_4010,N_4967);
nor UO_348 (O_348,N_4957,N_4903);
and UO_349 (O_349,N_4721,N_4964);
nand UO_350 (O_350,N_4701,N_4828);
nand UO_351 (O_351,N_4689,N_4182);
or UO_352 (O_352,N_4036,N_4317);
and UO_353 (O_353,N_4528,N_4341);
nand UO_354 (O_354,N_4878,N_4209);
nand UO_355 (O_355,N_4555,N_4236);
nand UO_356 (O_356,N_4301,N_4717);
nor UO_357 (O_357,N_4467,N_4047);
nand UO_358 (O_358,N_4307,N_4956);
nor UO_359 (O_359,N_4207,N_4297);
nor UO_360 (O_360,N_4364,N_4538);
nand UO_361 (O_361,N_4543,N_4729);
nand UO_362 (O_362,N_4101,N_4757);
nor UO_363 (O_363,N_4932,N_4547);
nor UO_364 (O_364,N_4479,N_4597);
or UO_365 (O_365,N_4789,N_4581);
nor UO_366 (O_366,N_4305,N_4963);
and UO_367 (O_367,N_4019,N_4542);
xnor UO_368 (O_368,N_4806,N_4808);
nand UO_369 (O_369,N_4871,N_4409);
and UO_370 (O_370,N_4734,N_4742);
and UO_371 (O_371,N_4799,N_4732);
nand UO_372 (O_372,N_4334,N_4984);
nand UO_373 (O_373,N_4097,N_4709);
nand UO_374 (O_374,N_4784,N_4391);
or UO_375 (O_375,N_4958,N_4027);
and UO_376 (O_376,N_4173,N_4651);
xor UO_377 (O_377,N_4436,N_4480);
and UO_378 (O_378,N_4031,N_4029);
nand UO_379 (O_379,N_4077,N_4976);
nor UO_380 (O_380,N_4896,N_4426);
nand UO_381 (O_381,N_4323,N_4930);
and UO_382 (O_382,N_4390,N_4610);
nor UO_383 (O_383,N_4722,N_4327);
and UO_384 (O_384,N_4318,N_4999);
nand UO_385 (O_385,N_4856,N_4788);
or UO_386 (O_386,N_4181,N_4589);
nand UO_387 (O_387,N_4157,N_4488);
nor UO_388 (O_388,N_4016,N_4137);
nand UO_389 (O_389,N_4901,N_4905);
xor UO_390 (O_390,N_4442,N_4275);
nand UO_391 (O_391,N_4915,N_4322);
and UO_392 (O_392,N_4913,N_4418);
or UO_393 (O_393,N_4880,N_4640);
and UO_394 (O_394,N_4124,N_4079);
nand UO_395 (O_395,N_4803,N_4243);
or UO_396 (O_396,N_4664,N_4894);
nand UO_397 (O_397,N_4128,N_4523);
nor UO_398 (O_398,N_4698,N_4009);
or UO_399 (O_399,N_4231,N_4960);
and UO_400 (O_400,N_4710,N_4863);
and UO_401 (O_401,N_4515,N_4372);
nor UO_402 (O_402,N_4092,N_4175);
and UO_403 (O_403,N_4050,N_4615);
and UO_404 (O_404,N_4939,N_4347);
nand UO_405 (O_405,N_4602,N_4482);
nand UO_406 (O_406,N_4802,N_4261);
and UO_407 (O_407,N_4098,N_4786);
nand UO_408 (O_408,N_4382,N_4075);
and UO_409 (O_409,N_4149,N_4176);
and UO_410 (O_410,N_4094,N_4570);
nor UO_411 (O_411,N_4074,N_4342);
xor UO_412 (O_412,N_4143,N_4328);
nor UO_413 (O_413,N_4907,N_4304);
nand UO_414 (O_414,N_4711,N_4614);
or UO_415 (O_415,N_4477,N_4553);
and UO_416 (O_416,N_4224,N_4107);
nor UO_417 (O_417,N_4320,N_4969);
or UO_418 (O_418,N_4208,N_4151);
nand UO_419 (O_419,N_4257,N_4350);
or UO_420 (O_420,N_4308,N_4460);
and UO_421 (O_421,N_4095,N_4928);
nand UO_422 (O_422,N_4102,N_4378);
nor UO_423 (O_423,N_4314,N_4475);
nand UO_424 (O_424,N_4294,N_4919);
nand UO_425 (O_425,N_4211,N_4584);
or UO_426 (O_426,N_4039,N_4396);
or UO_427 (O_427,N_4517,N_4851);
nand UO_428 (O_428,N_4727,N_4665);
nor UO_429 (O_429,N_4355,N_4439);
nand UO_430 (O_430,N_4366,N_4720);
and UO_431 (O_431,N_4576,N_4754);
xnor UO_432 (O_432,N_4219,N_4147);
and UO_433 (O_433,N_4771,N_4130);
nor UO_434 (O_434,N_4357,N_4361);
nor UO_435 (O_435,N_4861,N_4335);
xor UO_436 (O_436,N_4506,N_4262);
nand UO_437 (O_437,N_4346,N_4692);
or UO_438 (O_438,N_4623,N_4221);
or UO_439 (O_439,N_4203,N_4702);
or UO_440 (O_440,N_4462,N_4949);
nand UO_441 (O_441,N_4011,N_4348);
nor UO_442 (O_442,N_4599,N_4500);
or UO_443 (O_443,N_4198,N_4196);
or UO_444 (O_444,N_4566,N_4457);
and UO_445 (O_445,N_4411,N_4741);
and UO_446 (O_446,N_4972,N_4835);
nand UO_447 (O_447,N_4267,N_4519);
or UO_448 (O_448,N_4252,N_4258);
and UO_449 (O_449,N_4407,N_4751);
and UO_450 (O_450,N_4402,N_4499);
and UO_451 (O_451,N_4509,N_4923);
nor UO_452 (O_452,N_4798,N_4866);
nor UO_453 (O_453,N_4892,N_4562);
and UO_454 (O_454,N_4825,N_4745);
and UO_455 (O_455,N_4423,N_4218);
or UO_456 (O_456,N_4474,N_4146);
and UO_457 (O_457,N_4099,N_4054);
nand UO_458 (O_458,N_4763,N_4184);
and UO_459 (O_459,N_4165,N_4807);
and UO_460 (O_460,N_4138,N_4410);
and UO_461 (O_461,N_4926,N_4443);
nand UO_462 (O_462,N_4657,N_4279);
and UO_463 (O_463,N_4619,N_4680);
nor UO_464 (O_464,N_4596,N_4608);
or UO_465 (O_465,N_4685,N_4332);
nand UO_466 (O_466,N_4170,N_4012);
nand UO_467 (O_467,N_4331,N_4082);
or UO_468 (O_468,N_4898,N_4394);
or UO_469 (O_469,N_4977,N_4622);
nor UO_470 (O_470,N_4988,N_4937);
nand UO_471 (O_471,N_4768,N_4947);
nand UO_472 (O_472,N_4507,N_4293);
nand UO_473 (O_473,N_4946,N_4910);
or UO_474 (O_474,N_4940,N_4044);
nand UO_475 (O_475,N_4060,N_4164);
or UO_476 (O_476,N_4451,N_4637);
nand UO_477 (O_477,N_4136,N_4445);
nor UO_478 (O_478,N_4677,N_4766);
or UO_479 (O_479,N_4801,N_4503);
nor UO_480 (O_480,N_4815,N_4311);
and UO_481 (O_481,N_4035,N_4159);
or UO_482 (O_482,N_4579,N_4719);
nor UO_483 (O_483,N_4201,N_4583);
nor UO_484 (O_484,N_4417,N_4982);
nand UO_485 (O_485,N_4646,N_4731);
and UO_486 (O_486,N_4514,N_4931);
or UO_487 (O_487,N_4968,N_4220);
or UO_488 (O_488,N_4544,N_4370);
xor UO_489 (O_489,N_4636,N_4783);
and UO_490 (O_490,N_4416,N_4616);
nor UO_491 (O_491,N_4654,N_4557);
nand UO_492 (O_492,N_4524,N_4213);
and UO_493 (O_493,N_4241,N_4395);
or UO_494 (O_494,N_4575,N_4472);
nand UO_495 (O_495,N_4838,N_4559);
nor UO_496 (O_496,N_4365,N_4565);
nand UO_497 (O_497,N_4805,N_4906);
or UO_498 (O_498,N_4585,N_4889);
nor UO_499 (O_499,N_4595,N_4021);
nor UO_500 (O_500,N_4176,N_4847);
or UO_501 (O_501,N_4334,N_4410);
nand UO_502 (O_502,N_4855,N_4164);
nand UO_503 (O_503,N_4953,N_4403);
nor UO_504 (O_504,N_4615,N_4884);
nor UO_505 (O_505,N_4395,N_4415);
and UO_506 (O_506,N_4891,N_4802);
and UO_507 (O_507,N_4435,N_4017);
nand UO_508 (O_508,N_4995,N_4627);
nor UO_509 (O_509,N_4969,N_4656);
nand UO_510 (O_510,N_4684,N_4537);
nand UO_511 (O_511,N_4395,N_4291);
nor UO_512 (O_512,N_4707,N_4694);
nand UO_513 (O_513,N_4613,N_4689);
nor UO_514 (O_514,N_4798,N_4776);
nand UO_515 (O_515,N_4508,N_4460);
and UO_516 (O_516,N_4420,N_4246);
nand UO_517 (O_517,N_4889,N_4644);
nand UO_518 (O_518,N_4164,N_4650);
nor UO_519 (O_519,N_4884,N_4906);
or UO_520 (O_520,N_4908,N_4006);
and UO_521 (O_521,N_4350,N_4052);
or UO_522 (O_522,N_4063,N_4592);
nand UO_523 (O_523,N_4755,N_4459);
or UO_524 (O_524,N_4002,N_4221);
nor UO_525 (O_525,N_4120,N_4494);
and UO_526 (O_526,N_4921,N_4966);
and UO_527 (O_527,N_4494,N_4678);
or UO_528 (O_528,N_4547,N_4455);
nand UO_529 (O_529,N_4261,N_4636);
or UO_530 (O_530,N_4978,N_4822);
nor UO_531 (O_531,N_4282,N_4917);
and UO_532 (O_532,N_4573,N_4771);
or UO_533 (O_533,N_4231,N_4350);
nor UO_534 (O_534,N_4240,N_4731);
or UO_535 (O_535,N_4458,N_4640);
nor UO_536 (O_536,N_4879,N_4902);
nand UO_537 (O_537,N_4905,N_4149);
and UO_538 (O_538,N_4836,N_4456);
nor UO_539 (O_539,N_4577,N_4818);
nor UO_540 (O_540,N_4831,N_4877);
xor UO_541 (O_541,N_4045,N_4719);
or UO_542 (O_542,N_4023,N_4078);
and UO_543 (O_543,N_4069,N_4629);
nor UO_544 (O_544,N_4682,N_4575);
nand UO_545 (O_545,N_4252,N_4943);
nor UO_546 (O_546,N_4999,N_4566);
and UO_547 (O_547,N_4080,N_4256);
nand UO_548 (O_548,N_4283,N_4691);
and UO_549 (O_549,N_4173,N_4157);
nor UO_550 (O_550,N_4482,N_4101);
nor UO_551 (O_551,N_4539,N_4818);
or UO_552 (O_552,N_4900,N_4262);
nor UO_553 (O_553,N_4315,N_4959);
or UO_554 (O_554,N_4078,N_4943);
or UO_555 (O_555,N_4705,N_4933);
and UO_556 (O_556,N_4943,N_4126);
nor UO_557 (O_557,N_4199,N_4979);
or UO_558 (O_558,N_4042,N_4861);
or UO_559 (O_559,N_4737,N_4804);
or UO_560 (O_560,N_4060,N_4767);
and UO_561 (O_561,N_4275,N_4649);
nor UO_562 (O_562,N_4052,N_4761);
nand UO_563 (O_563,N_4490,N_4337);
and UO_564 (O_564,N_4914,N_4054);
or UO_565 (O_565,N_4513,N_4433);
nor UO_566 (O_566,N_4295,N_4502);
nor UO_567 (O_567,N_4236,N_4929);
nand UO_568 (O_568,N_4578,N_4031);
and UO_569 (O_569,N_4551,N_4014);
nand UO_570 (O_570,N_4891,N_4525);
nor UO_571 (O_571,N_4199,N_4714);
nor UO_572 (O_572,N_4607,N_4957);
and UO_573 (O_573,N_4057,N_4741);
nand UO_574 (O_574,N_4603,N_4228);
or UO_575 (O_575,N_4739,N_4799);
and UO_576 (O_576,N_4515,N_4782);
nor UO_577 (O_577,N_4486,N_4861);
nor UO_578 (O_578,N_4056,N_4086);
and UO_579 (O_579,N_4999,N_4591);
or UO_580 (O_580,N_4753,N_4520);
nand UO_581 (O_581,N_4937,N_4308);
nand UO_582 (O_582,N_4318,N_4911);
or UO_583 (O_583,N_4089,N_4991);
or UO_584 (O_584,N_4317,N_4505);
and UO_585 (O_585,N_4810,N_4953);
and UO_586 (O_586,N_4612,N_4413);
and UO_587 (O_587,N_4031,N_4813);
nor UO_588 (O_588,N_4106,N_4861);
and UO_589 (O_589,N_4835,N_4427);
or UO_590 (O_590,N_4987,N_4771);
nor UO_591 (O_591,N_4229,N_4782);
and UO_592 (O_592,N_4641,N_4415);
or UO_593 (O_593,N_4216,N_4497);
nor UO_594 (O_594,N_4204,N_4380);
nand UO_595 (O_595,N_4685,N_4506);
and UO_596 (O_596,N_4618,N_4794);
nor UO_597 (O_597,N_4090,N_4909);
nor UO_598 (O_598,N_4780,N_4785);
nor UO_599 (O_599,N_4408,N_4354);
nand UO_600 (O_600,N_4597,N_4077);
nor UO_601 (O_601,N_4293,N_4738);
nor UO_602 (O_602,N_4040,N_4336);
nand UO_603 (O_603,N_4459,N_4068);
nand UO_604 (O_604,N_4875,N_4766);
nand UO_605 (O_605,N_4630,N_4201);
nand UO_606 (O_606,N_4036,N_4292);
nand UO_607 (O_607,N_4886,N_4924);
or UO_608 (O_608,N_4981,N_4447);
nor UO_609 (O_609,N_4369,N_4777);
nand UO_610 (O_610,N_4306,N_4676);
nand UO_611 (O_611,N_4489,N_4638);
or UO_612 (O_612,N_4768,N_4898);
nor UO_613 (O_613,N_4208,N_4003);
or UO_614 (O_614,N_4994,N_4355);
and UO_615 (O_615,N_4296,N_4710);
or UO_616 (O_616,N_4034,N_4979);
nor UO_617 (O_617,N_4747,N_4656);
nor UO_618 (O_618,N_4764,N_4974);
nand UO_619 (O_619,N_4969,N_4978);
or UO_620 (O_620,N_4178,N_4527);
or UO_621 (O_621,N_4630,N_4591);
nand UO_622 (O_622,N_4326,N_4092);
and UO_623 (O_623,N_4962,N_4221);
nand UO_624 (O_624,N_4039,N_4772);
and UO_625 (O_625,N_4194,N_4575);
or UO_626 (O_626,N_4645,N_4922);
or UO_627 (O_627,N_4326,N_4869);
or UO_628 (O_628,N_4899,N_4519);
and UO_629 (O_629,N_4251,N_4853);
and UO_630 (O_630,N_4978,N_4538);
and UO_631 (O_631,N_4807,N_4856);
or UO_632 (O_632,N_4270,N_4737);
or UO_633 (O_633,N_4529,N_4492);
nor UO_634 (O_634,N_4985,N_4445);
xnor UO_635 (O_635,N_4866,N_4409);
or UO_636 (O_636,N_4312,N_4012);
nand UO_637 (O_637,N_4688,N_4342);
and UO_638 (O_638,N_4283,N_4276);
or UO_639 (O_639,N_4338,N_4243);
or UO_640 (O_640,N_4111,N_4945);
nand UO_641 (O_641,N_4312,N_4661);
nor UO_642 (O_642,N_4052,N_4995);
and UO_643 (O_643,N_4484,N_4812);
nand UO_644 (O_644,N_4592,N_4847);
or UO_645 (O_645,N_4775,N_4952);
xnor UO_646 (O_646,N_4477,N_4016);
nand UO_647 (O_647,N_4513,N_4833);
nand UO_648 (O_648,N_4133,N_4438);
and UO_649 (O_649,N_4106,N_4949);
nor UO_650 (O_650,N_4909,N_4601);
nor UO_651 (O_651,N_4658,N_4223);
or UO_652 (O_652,N_4895,N_4553);
or UO_653 (O_653,N_4702,N_4814);
or UO_654 (O_654,N_4407,N_4791);
nand UO_655 (O_655,N_4258,N_4846);
or UO_656 (O_656,N_4750,N_4409);
or UO_657 (O_657,N_4457,N_4237);
and UO_658 (O_658,N_4810,N_4256);
and UO_659 (O_659,N_4266,N_4192);
xnor UO_660 (O_660,N_4010,N_4663);
nand UO_661 (O_661,N_4597,N_4505);
nor UO_662 (O_662,N_4205,N_4893);
nand UO_663 (O_663,N_4045,N_4602);
nor UO_664 (O_664,N_4468,N_4661);
nor UO_665 (O_665,N_4146,N_4517);
nand UO_666 (O_666,N_4787,N_4130);
and UO_667 (O_667,N_4125,N_4370);
and UO_668 (O_668,N_4007,N_4442);
or UO_669 (O_669,N_4954,N_4174);
and UO_670 (O_670,N_4696,N_4857);
nand UO_671 (O_671,N_4600,N_4971);
and UO_672 (O_672,N_4887,N_4165);
nand UO_673 (O_673,N_4093,N_4684);
nand UO_674 (O_674,N_4891,N_4619);
and UO_675 (O_675,N_4268,N_4775);
nor UO_676 (O_676,N_4747,N_4319);
or UO_677 (O_677,N_4190,N_4019);
nor UO_678 (O_678,N_4943,N_4042);
nand UO_679 (O_679,N_4343,N_4620);
and UO_680 (O_680,N_4240,N_4712);
nor UO_681 (O_681,N_4494,N_4813);
nor UO_682 (O_682,N_4526,N_4755);
nor UO_683 (O_683,N_4729,N_4106);
or UO_684 (O_684,N_4885,N_4911);
nor UO_685 (O_685,N_4079,N_4399);
or UO_686 (O_686,N_4052,N_4263);
or UO_687 (O_687,N_4182,N_4342);
and UO_688 (O_688,N_4940,N_4366);
nand UO_689 (O_689,N_4417,N_4613);
or UO_690 (O_690,N_4104,N_4954);
or UO_691 (O_691,N_4173,N_4942);
nor UO_692 (O_692,N_4617,N_4173);
nand UO_693 (O_693,N_4139,N_4452);
and UO_694 (O_694,N_4316,N_4643);
nor UO_695 (O_695,N_4128,N_4161);
nor UO_696 (O_696,N_4177,N_4769);
or UO_697 (O_697,N_4287,N_4796);
or UO_698 (O_698,N_4762,N_4520);
and UO_699 (O_699,N_4624,N_4663);
nor UO_700 (O_700,N_4585,N_4483);
nor UO_701 (O_701,N_4981,N_4111);
and UO_702 (O_702,N_4539,N_4117);
nor UO_703 (O_703,N_4702,N_4173);
and UO_704 (O_704,N_4495,N_4888);
or UO_705 (O_705,N_4420,N_4298);
nor UO_706 (O_706,N_4084,N_4673);
and UO_707 (O_707,N_4463,N_4133);
nand UO_708 (O_708,N_4255,N_4314);
nand UO_709 (O_709,N_4507,N_4358);
nor UO_710 (O_710,N_4152,N_4064);
and UO_711 (O_711,N_4293,N_4443);
and UO_712 (O_712,N_4885,N_4969);
or UO_713 (O_713,N_4105,N_4506);
and UO_714 (O_714,N_4660,N_4576);
and UO_715 (O_715,N_4559,N_4223);
or UO_716 (O_716,N_4298,N_4381);
and UO_717 (O_717,N_4917,N_4252);
or UO_718 (O_718,N_4690,N_4055);
and UO_719 (O_719,N_4741,N_4716);
nand UO_720 (O_720,N_4580,N_4348);
nand UO_721 (O_721,N_4639,N_4502);
nand UO_722 (O_722,N_4198,N_4262);
and UO_723 (O_723,N_4023,N_4224);
or UO_724 (O_724,N_4627,N_4341);
nand UO_725 (O_725,N_4147,N_4822);
nor UO_726 (O_726,N_4871,N_4545);
and UO_727 (O_727,N_4354,N_4377);
nand UO_728 (O_728,N_4722,N_4888);
nand UO_729 (O_729,N_4356,N_4607);
or UO_730 (O_730,N_4688,N_4961);
nand UO_731 (O_731,N_4894,N_4288);
or UO_732 (O_732,N_4938,N_4930);
and UO_733 (O_733,N_4442,N_4947);
nor UO_734 (O_734,N_4811,N_4923);
and UO_735 (O_735,N_4972,N_4636);
nor UO_736 (O_736,N_4745,N_4620);
nor UO_737 (O_737,N_4896,N_4858);
or UO_738 (O_738,N_4234,N_4557);
nor UO_739 (O_739,N_4849,N_4809);
and UO_740 (O_740,N_4790,N_4537);
nand UO_741 (O_741,N_4394,N_4366);
or UO_742 (O_742,N_4543,N_4326);
and UO_743 (O_743,N_4938,N_4363);
or UO_744 (O_744,N_4132,N_4293);
and UO_745 (O_745,N_4691,N_4360);
or UO_746 (O_746,N_4466,N_4740);
or UO_747 (O_747,N_4531,N_4249);
nor UO_748 (O_748,N_4794,N_4933);
nand UO_749 (O_749,N_4055,N_4526);
nor UO_750 (O_750,N_4274,N_4000);
nand UO_751 (O_751,N_4946,N_4923);
nand UO_752 (O_752,N_4648,N_4154);
nand UO_753 (O_753,N_4076,N_4643);
nand UO_754 (O_754,N_4838,N_4633);
nor UO_755 (O_755,N_4350,N_4151);
nand UO_756 (O_756,N_4297,N_4079);
nand UO_757 (O_757,N_4721,N_4158);
nor UO_758 (O_758,N_4442,N_4266);
nand UO_759 (O_759,N_4615,N_4106);
nor UO_760 (O_760,N_4882,N_4503);
or UO_761 (O_761,N_4677,N_4668);
and UO_762 (O_762,N_4633,N_4003);
or UO_763 (O_763,N_4772,N_4087);
or UO_764 (O_764,N_4717,N_4400);
nand UO_765 (O_765,N_4268,N_4606);
and UO_766 (O_766,N_4076,N_4702);
or UO_767 (O_767,N_4903,N_4584);
or UO_768 (O_768,N_4209,N_4230);
nand UO_769 (O_769,N_4709,N_4265);
and UO_770 (O_770,N_4460,N_4431);
nor UO_771 (O_771,N_4225,N_4140);
or UO_772 (O_772,N_4635,N_4948);
nor UO_773 (O_773,N_4987,N_4246);
nand UO_774 (O_774,N_4245,N_4307);
or UO_775 (O_775,N_4418,N_4787);
or UO_776 (O_776,N_4639,N_4977);
nand UO_777 (O_777,N_4343,N_4118);
or UO_778 (O_778,N_4852,N_4921);
nor UO_779 (O_779,N_4914,N_4895);
and UO_780 (O_780,N_4284,N_4037);
and UO_781 (O_781,N_4737,N_4609);
or UO_782 (O_782,N_4790,N_4511);
nand UO_783 (O_783,N_4204,N_4645);
and UO_784 (O_784,N_4415,N_4202);
or UO_785 (O_785,N_4691,N_4622);
or UO_786 (O_786,N_4943,N_4670);
nand UO_787 (O_787,N_4740,N_4527);
xnor UO_788 (O_788,N_4087,N_4485);
or UO_789 (O_789,N_4979,N_4056);
nor UO_790 (O_790,N_4690,N_4977);
or UO_791 (O_791,N_4078,N_4712);
nand UO_792 (O_792,N_4389,N_4717);
and UO_793 (O_793,N_4461,N_4796);
nand UO_794 (O_794,N_4720,N_4779);
and UO_795 (O_795,N_4133,N_4630);
nand UO_796 (O_796,N_4570,N_4276);
or UO_797 (O_797,N_4392,N_4309);
nand UO_798 (O_798,N_4922,N_4523);
or UO_799 (O_799,N_4455,N_4783);
and UO_800 (O_800,N_4516,N_4657);
nand UO_801 (O_801,N_4522,N_4313);
and UO_802 (O_802,N_4424,N_4897);
and UO_803 (O_803,N_4397,N_4425);
and UO_804 (O_804,N_4934,N_4363);
nor UO_805 (O_805,N_4440,N_4308);
nor UO_806 (O_806,N_4712,N_4738);
or UO_807 (O_807,N_4242,N_4652);
nand UO_808 (O_808,N_4715,N_4166);
or UO_809 (O_809,N_4788,N_4482);
nor UO_810 (O_810,N_4551,N_4166);
nand UO_811 (O_811,N_4506,N_4484);
and UO_812 (O_812,N_4261,N_4718);
and UO_813 (O_813,N_4058,N_4585);
nor UO_814 (O_814,N_4205,N_4081);
or UO_815 (O_815,N_4558,N_4407);
nand UO_816 (O_816,N_4090,N_4521);
nand UO_817 (O_817,N_4406,N_4062);
nand UO_818 (O_818,N_4496,N_4272);
nand UO_819 (O_819,N_4024,N_4894);
nor UO_820 (O_820,N_4800,N_4807);
nand UO_821 (O_821,N_4771,N_4110);
nor UO_822 (O_822,N_4992,N_4526);
or UO_823 (O_823,N_4868,N_4744);
nor UO_824 (O_824,N_4429,N_4798);
and UO_825 (O_825,N_4139,N_4247);
or UO_826 (O_826,N_4882,N_4916);
and UO_827 (O_827,N_4712,N_4306);
and UO_828 (O_828,N_4738,N_4118);
nor UO_829 (O_829,N_4775,N_4982);
and UO_830 (O_830,N_4905,N_4203);
and UO_831 (O_831,N_4937,N_4568);
nand UO_832 (O_832,N_4801,N_4031);
and UO_833 (O_833,N_4257,N_4185);
or UO_834 (O_834,N_4513,N_4010);
nor UO_835 (O_835,N_4913,N_4864);
xor UO_836 (O_836,N_4091,N_4598);
nand UO_837 (O_837,N_4824,N_4995);
nand UO_838 (O_838,N_4726,N_4463);
and UO_839 (O_839,N_4511,N_4570);
or UO_840 (O_840,N_4238,N_4462);
nor UO_841 (O_841,N_4011,N_4404);
nor UO_842 (O_842,N_4484,N_4515);
and UO_843 (O_843,N_4089,N_4884);
nand UO_844 (O_844,N_4488,N_4803);
nor UO_845 (O_845,N_4379,N_4292);
nor UO_846 (O_846,N_4569,N_4428);
nor UO_847 (O_847,N_4063,N_4813);
nor UO_848 (O_848,N_4507,N_4142);
and UO_849 (O_849,N_4208,N_4966);
nor UO_850 (O_850,N_4909,N_4252);
nor UO_851 (O_851,N_4661,N_4531);
nand UO_852 (O_852,N_4640,N_4238);
nor UO_853 (O_853,N_4447,N_4610);
or UO_854 (O_854,N_4177,N_4547);
nand UO_855 (O_855,N_4434,N_4827);
nor UO_856 (O_856,N_4479,N_4239);
or UO_857 (O_857,N_4840,N_4386);
nor UO_858 (O_858,N_4234,N_4648);
and UO_859 (O_859,N_4828,N_4295);
nor UO_860 (O_860,N_4538,N_4554);
and UO_861 (O_861,N_4281,N_4907);
nand UO_862 (O_862,N_4969,N_4153);
or UO_863 (O_863,N_4869,N_4258);
nor UO_864 (O_864,N_4007,N_4616);
nand UO_865 (O_865,N_4664,N_4768);
nand UO_866 (O_866,N_4486,N_4673);
nand UO_867 (O_867,N_4602,N_4047);
nand UO_868 (O_868,N_4915,N_4088);
or UO_869 (O_869,N_4483,N_4615);
nand UO_870 (O_870,N_4383,N_4722);
nor UO_871 (O_871,N_4502,N_4539);
nor UO_872 (O_872,N_4025,N_4573);
nor UO_873 (O_873,N_4260,N_4253);
nor UO_874 (O_874,N_4993,N_4116);
nor UO_875 (O_875,N_4721,N_4890);
nand UO_876 (O_876,N_4019,N_4661);
nand UO_877 (O_877,N_4400,N_4741);
or UO_878 (O_878,N_4642,N_4825);
or UO_879 (O_879,N_4025,N_4397);
and UO_880 (O_880,N_4598,N_4776);
or UO_881 (O_881,N_4790,N_4747);
or UO_882 (O_882,N_4422,N_4389);
nand UO_883 (O_883,N_4383,N_4616);
or UO_884 (O_884,N_4649,N_4121);
nand UO_885 (O_885,N_4404,N_4551);
nand UO_886 (O_886,N_4558,N_4660);
nor UO_887 (O_887,N_4561,N_4446);
or UO_888 (O_888,N_4144,N_4679);
and UO_889 (O_889,N_4767,N_4607);
and UO_890 (O_890,N_4833,N_4300);
nor UO_891 (O_891,N_4372,N_4373);
nor UO_892 (O_892,N_4412,N_4527);
and UO_893 (O_893,N_4304,N_4667);
or UO_894 (O_894,N_4348,N_4462);
and UO_895 (O_895,N_4310,N_4794);
nor UO_896 (O_896,N_4465,N_4271);
nor UO_897 (O_897,N_4369,N_4733);
or UO_898 (O_898,N_4972,N_4626);
nor UO_899 (O_899,N_4142,N_4064);
or UO_900 (O_900,N_4641,N_4663);
and UO_901 (O_901,N_4391,N_4738);
nand UO_902 (O_902,N_4343,N_4836);
nand UO_903 (O_903,N_4007,N_4590);
xnor UO_904 (O_904,N_4538,N_4549);
and UO_905 (O_905,N_4810,N_4592);
and UO_906 (O_906,N_4282,N_4220);
and UO_907 (O_907,N_4755,N_4041);
nor UO_908 (O_908,N_4165,N_4248);
and UO_909 (O_909,N_4074,N_4191);
nor UO_910 (O_910,N_4734,N_4357);
or UO_911 (O_911,N_4183,N_4697);
nor UO_912 (O_912,N_4533,N_4330);
or UO_913 (O_913,N_4838,N_4808);
or UO_914 (O_914,N_4662,N_4836);
or UO_915 (O_915,N_4596,N_4155);
nor UO_916 (O_916,N_4216,N_4210);
or UO_917 (O_917,N_4330,N_4216);
and UO_918 (O_918,N_4696,N_4053);
nor UO_919 (O_919,N_4576,N_4144);
or UO_920 (O_920,N_4806,N_4797);
and UO_921 (O_921,N_4810,N_4430);
and UO_922 (O_922,N_4422,N_4567);
and UO_923 (O_923,N_4677,N_4616);
nor UO_924 (O_924,N_4078,N_4933);
nor UO_925 (O_925,N_4190,N_4257);
or UO_926 (O_926,N_4567,N_4530);
and UO_927 (O_927,N_4956,N_4105);
nor UO_928 (O_928,N_4840,N_4918);
nand UO_929 (O_929,N_4757,N_4907);
and UO_930 (O_930,N_4247,N_4502);
nor UO_931 (O_931,N_4909,N_4485);
nor UO_932 (O_932,N_4482,N_4622);
or UO_933 (O_933,N_4382,N_4319);
and UO_934 (O_934,N_4940,N_4041);
nand UO_935 (O_935,N_4627,N_4183);
or UO_936 (O_936,N_4855,N_4608);
nor UO_937 (O_937,N_4069,N_4186);
and UO_938 (O_938,N_4356,N_4821);
or UO_939 (O_939,N_4077,N_4901);
nand UO_940 (O_940,N_4560,N_4553);
nand UO_941 (O_941,N_4690,N_4287);
nor UO_942 (O_942,N_4516,N_4920);
or UO_943 (O_943,N_4722,N_4337);
and UO_944 (O_944,N_4658,N_4139);
nor UO_945 (O_945,N_4008,N_4243);
nor UO_946 (O_946,N_4127,N_4245);
or UO_947 (O_947,N_4754,N_4206);
or UO_948 (O_948,N_4588,N_4777);
nor UO_949 (O_949,N_4513,N_4592);
nand UO_950 (O_950,N_4101,N_4122);
or UO_951 (O_951,N_4760,N_4743);
nand UO_952 (O_952,N_4629,N_4318);
and UO_953 (O_953,N_4389,N_4163);
nor UO_954 (O_954,N_4092,N_4150);
and UO_955 (O_955,N_4619,N_4118);
nor UO_956 (O_956,N_4175,N_4734);
or UO_957 (O_957,N_4766,N_4936);
nor UO_958 (O_958,N_4882,N_4299);
or UO_959 (O_959,N_4350,N_4193);
or UO_960 (O_960,N_4090,N_4186);
nor UO_961 (O_961,N_4614,N_4177);
or UO_962 (O_962,N_4322,N_4185);
or UO_963 (O_963,N_4475,N_4819);
and UO_964 (O_964,N_4577,N_4407);
nor UO_965 (O_965,N_4275,N_4123);
nand UO_966 (O_966,N_4437,N_4285);
and UO_967 (O_967,N_4385,N_4550);
nand UO_968 (O_968,N_4190,N_4323);
or UO_969 (O_969,N_4358,N_4585);
or UO_970 (O_970,N_4887,N_4379);
and UO_971 (O_971,N_4208,N_4568);
and UO_972 (O_972,N_4716,N_4062);
nand UO_973 (O_973,N_4012,N_4741);
nand UO_974 (O_974,N_4115,N_4803);
or UO_975 (O_975,N_4896,N_4429);
nor UO_976 (O_976,N_4127,N_4531);
nor UO_977 (O_977,N_4253,N_4112);
and UO_978 (O_978,N_4475,N_4086);
or UO_979 (O_979,N_4368,N_4993);
or UO_980 (O_980,N_4165,N_4855);
and UO_981 (O_981,N_4098,N_4147);
or UO_982 (O_982,N_4137,N_4037);
or UO_983 (O_983,N_4291,N_4359);
nand UO_984 (O_984,N_4567,N_4464);
or UO_985 (O_985,N_4024,N_4431);
and UO_986 (O_986,N_4421,N_4428);
nor UO_987 (O_987,N_4389,N_4583);
nor UO_988 (O_988,N_4879,N_4458);
and UO_989 (O_989,N_4626,N_4697);
nor UO_990 (O_990,N_4533,N_4663);
or UO_991 (O_991,N_4633,N_4745);
or UO_992 (O_992,N_4352,N_4997);
or UO_993 (O_993,N_4766,N_4910);
nor UO_994 (O_994,N_4601,N_4925);
nor UO_995 (O_995,N_4040,N_4419);
and UO_996 (O_996,N_4569,N_4648);
and UO_997 (O_997,N_4633,N_4308);
and UO_998 (O_998,N_4039,N_4460);
or UO_999 (O_999,N_4639,N_4287);
endmodule