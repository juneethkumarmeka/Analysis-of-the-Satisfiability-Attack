module basic_750_5000_1000_25_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_28,In_101);
nor U1 (N_1,In_390,In_746);
or U2 (N_2,In_286,In_312);
xnor U3 (N_3,In_505,In_215);
nor U4 (N_4,In_375,In_659);
or U5 (N_5,In_330,In_747);
and U6 (N_6,In_151,In_598);
nor U7 (N_7,In_324,In_541);
or U8 (N_8,In_479,In_677);
nand U9 (N_9,In_601,In_696);
or U10 (N_10,In_449,In_511);
xnor U11 (N_11,In_251,In_535);
nor U12 (N_12,In_412,In_252);
or U13 (N_13,In_701,In_409);
nor U14 (N_14,In_315,In_456);
nor U15 (N_15,In_154,In_738);
or U16 (N_16,In_147,In_649);
xnor U17 (N_17,In_99,In_366);
nand U18 (N_18,In_407,In_382);
nor U19 (N_19,In_670,In_303);
and U20 (N_20,In_719,In_248);
or U21 (N_21,In_193,In_439);
nor U22 (N_22,In_727,In_432);
nand U23 (N_23,In_629,In_107);
nand U24 (N_24,In_219,In_437);
and U25 (N_25,In_524,In_499);
nand U26 (N_26,In_120,In_344);
and U27 (N_27,In_27,In_92);
or U28 (N_28,In_669,In_185);
and U29 (N_29,In_295,In_34);
xnor U30 (N_30,In_387,In_265);
nand U31 (N_31,In_273,In_357);
nor U32 (N_32,In_64,In_322);
nand U33 (N_33,In_373,In_9);
and U34 (N_34,In_579,In_229);
or U35 (N_35,In_413,In_451);
and U36 (N_36,In_143,In_411);
or U37 (N_37,In_179,In_171);
and U38 (N_38,In_586,In_492);
nand U39 (N_39,In_194,In_292);
nand U40 (N_40,In_381,In_630);
nand U41 (N_41,In_678,In_406);
nand U42 (N_42,In_686,In_305);
nand U43 (N_43,In_331,In_213);
and U44 (N_44,In_155,In_53);
or U45 (N_45,In_163,In_724);
nand U46 (N_46,In_7,In_567);
xnor U47 (N_47,In_580,In_323);
nor U48 (N_48,In_442,In_455);
and U49 (N_49,In_426,In_129);
and U50 (N_50,In_733,In_369);
and U51 (N_51,In_249,In_573);
or U52 (N_52,In_484,In_250);
and U53 (N_53,In_21,In_436);
xor U54 (N_54,In_658,In_632);
xor U55 (N_55,In_235,In_17);
nor U56 (N_56,In_731,In_201);
xor U57 (N_57,In_648,In_350);
nor U58 (N_58,In_198,In_278);
and U59 (N_59,In_145,In_564);
and U60 (N_60,In_207,In_48);
or U61 (N_61,In_689,In_142);
xnor U62 (N_62,In_540,In_467);
nand U63 (N_63,In_515,In_354);
nand U64 (N_64,In_539,In_279);
or U65 (N_65,In_110,In_512);
and U66 (N_66,In_137,In_584);
or U67 (N_67,In_135,In_531);
and U68 (N_68,In_404,In_58);
or U69 (N_69,In_55,In_191);
nor U70 (N_70,In_488,In_203);
nand U71 (N_71,In_594,In_370);
and U72 (N_72,In_304,In_87);
xnor U73 (N_73,In_743,In_418);
and U74 (N_74,In_386,In_236);
or U75 (N_75,In_617,In_328);
xor U76 (N_76,In_293,In_470);
nor U77 (N_77,In_52,In_321);
xor U78 (N_78,In_681,In_566);
nor U79 (N_79,In_359,In_486);
xor U80 (N_80,In_544,In_214);
xnor U81 (N_81,In_122,In_464);
and U82 (N_82,In_685,In_459);
nor U83 (N_83,In_634,In_656);
nor U84 (N_84,In_184,In_173);
or U85 (N_85,In_613,In_569);
nand U86 (N_86,In_161,In_337);
nor U87 (N_87,In_96,In_12);
or U88 (N_88,In_268,In_471);
nand U89 (N_89,In_523,In_644);
or U90 (N_90,In_698,In_410);
nand U91 (N_91,In_181,In_500);
xor U92 (N_92,In_454,In_542);
xnor U93 (N_93,In_647,In_425);
xor U94 (N_94,In_661,In_532);
and U95 (N_95,In_388,In_209);
and U96 (N_96,In_744,In_259);
and U97 (N_97,In_609,In_119);
xor U98 (N_98,In_98,In_57);
nor U99 (N_99,In_255,In_258);
and U100 (N_100,In_707,In_26);
or U101 (N_101,In_666,In_272);
and U102 (N_102,In_700,In_583);
nand U103 (N_103,In_285,In_671);
xor U104 (N_104,In_49,In_178);
and U105 (N_105,In_77,In_408);
xor U106 (N_106,In_296,In_559);
or U107 (N_107,In_317,In_25);
nand U108 (N_108,In_562,In_563);
or U109 (N_109,In_469,In_716);
xor U110 (N_110,In_231,In_428);
and U111 (N_111,In_614,In_624);
or U112 (N_112,In_402,In_551);
or U113 (N_113,In_503,In_38);
and U114 (N_114,In_189,In_74);
nor U115 (N_115,In_362,In_342);
nand U116 (N_116,In_336,In_391);
nor U117 (N_117,In_298,In_737);
or U118 (N_118,In_508,In_32);
nor U119 (N_119,In_473,In_620);
and U120 (N_120,In_663,In_282);
nor U121 (N_121,In_482,In_712);
xor U122 (N_122,In_177,In_11);
nor U123 (N_123,In_376,In_256);
nor U124 (N_124,In_146,In_734);
and U125 (N_125,In_104,In_16);
or U126 (N_126,In_24,In_489);
and U127 (N_127,In_434,In_622);
and U128 (N_128,In_684,In_136);
or U129 (N_129,In_90,In_314);
xor U130 (N_130,In_556,In_297);
or U131 (N_131,In_560,In_722);
and U132 (N_132,In_299,In_509);
nor U133 (N_133,In_550,In_596);
nor U134 (N_134,In_115,In_377);
nor U135 (N_135,In_218,In_160);
xnor U136 (N_136,In_385,In_233);
xor U137 (N_137,In_332,In_195);
nand U138 (N_138,In_54,In_168);
and U139 (N_139,In_497,In_623);
xor U140 (N_140,In_284,In_723);
nand U141 (N_141,In_138,In_513);
nand U142 (N_142,In_697,In_95);
nor U143 (N_143,In_237,In_414);
nor U144 (N_144,In_642,In_476);
or U145 (N_145,In_281,In_372);
or U146 (N_146,In_47,In_29);
and U147 (N_147,In_75,In_460);
xnor U148 (N_148,In_42,In_682);
nor U149 (N_149,In_525,In_130);
and U150 (N_150,In_275,In_326);
nand U151 (N_151,In_585,In_196);
xor U152 (N_152,In_529,In_234);
and U153 (N_153,In_393,In_157);
or U154 (N_154,In_520,In_263);
or U155 (N_155,In_557,In_483);
xor U156 (N_156,In_60,In_310);
and U157 (N_157,In_309,In_288);
and U158 (N_158,In_526,In_422);
nor U159 (N_159,In_444,In_496);
and U160 (N_160,In_687,In_695);
nand U161 (N_161,In_46,In_637);
nand U162 (N_162,In_748,In_175);
nand U163 (N_163,In_51,In_192);
xnor U164 (N_164,In_431,In_274);
nor U165 (N_165,In_23,In_225);
nor U166 (N_166,In_228,In_653);
and U167 (N_167,In_527,In_63);
or U168 (N_168,In_536,In_188);
nand U169 (N_169,In_170,In_453);
or U170 (N_170,In_302,In_243);
nor U171 (N_171,In_607,In_714);
xor U172 (N_172,In_144,In_223);
or U173 (N_173,In_35,In_635);
xnor U174 (N_174,In_472,In_591);
or U175 (N_175,In_577,In_18);
xor U176 (N_176,In_238,In_200);
nand U177 (N_177,In_334,In_291);
nand U178 (N_178,In_534,In_424);
or U179 (N_179,In_82,In_612);
nand U180 (N_180,In_216,In_461);
or U181 (N_181,In_389,In_668);
xnor U182 (N_182,In_679,In_240);
xor U183 (N_183,In_360,In_208);
xnor U184 (N_184,In_62,In_45);
nand U185 (N_185,In_589,In_169);
nor U186 (N_186,In_56,In_206);
nor U187 (N_187,In_106,In_39);
or U188 (N_188,In_131,In_538);
and U189 (N_189,In_61,In_545);
nand U190 (N_190,In_547,In_602);
and U191 (N_191,In_441,In_543);
nand U192 (N_192,In_19,In_380);
nor U193 (N_193,In_574,In_318);
and U194 (N_194,In_4,In_415);
nor U195 (N_195,In_537,In_148);
xnor U196 (N_196,In_108,In_552);
or U197 (N_197,In_133,In_14);
nor U198 (N_198,In_37,In_429);
nand U199 (N_199,In_313,In_43);
and U200 (N_200,In_260,N_16);
xnor U201 (N_201,In_205,In_735);
nor U202 (N_202,In_346,In_320);
or U203 (N_203,In_739,In_683);
and U204 (N_204,N_188,In_675);
or U205 (N_205,In_450,In_603);
nor U206 (N_206,In_266,In_162);
nand U207 (N_207,In_713,In_149);
or U208 (N_208,In_355,N_95);
and U209 (N_209,In_475,N_29);
or U210 (N_210,N_3,In_139);
xnor U211 (N_211,N_37,In_519);
and U212 (N_212,In_468,In_506);
and U213 (N_213,In_673,N_11);
and U214 (N_214,In_361,In_597);
or U215 (N_215,In_199,N_104);
and U216 (N_216,In_498,In_230);
nor U217 (N_217,N_64,In_638);
nand U218 (N_218,N_26,N_119);
or U219 (N_219,N_98,N_93);
nor U220 (N_220,In_561,N_73);
nor U221 (N_221,In_533,In_221);
xor U222 (N_222,N_142,In_246);
or U223 (N_223,N_53,N_149);
nand U224 (N_224,In_241,N_57);
nand U225 (N_225,In_174,N_152);
nor U226 (N_226,N_7,N_48);
nand U227 (N_227,N_132,N_179);
nor U228 (N_228,In_742,In_127);
or U229 (N_229,In_749,In_688);
or U230 (N_230,In_717,N_78);
nor U231 (N_231,In_572,N_153);
nor U232 (N_232,In_676,In_5);
or U233 (N_233,N_81,In_123);
xor U234 (N_234,In_31,In_319);
nand U235 (N_235,In_78,N_124);
xnor U236 (N_236,N_114,In_358);
or U237 (N_237,N_56,In_720);
xnor U238 (N_238,In_605,N_8);
nor U239 (N_239,N_150,In_244);
nor U240 (N_240,In_741,In_555);
and U241 (N_241,N_44,In_708);
nor U242 (N_242,In_399,N_143);
or U243 (N_243,In_491,N_67);
nor U244 (N_244,N_134,In_518);
xor U245 (N_245,In_264,In_71);
nand U246 (N_246,In_400,N_32);
nor U247 (N_247,In_277,In_433);
nand U248 (N_248,N_89,In_652);
xor U249 (N_249,In_481,N_110);
xor U250 (N_250,In_180,N_79);
xor U251 (N_251,In_384,N_109);
or U252 (N_252,In_2,In_655);
xnor U253 (N_253,In_116,In_628);
nor U254 (N_254,N_136,In_398);
or U255 (N_255,In_13,N_194);
xnor U256 (N_256,N_86,In_728);
nor U257 (N_257,In_50,In_553);
and U258 (N_258,In_97,In_72);
or U259 (N_259,In_445,N_61);
nor U260 (N_260,In_680,N_196);
nand U261 (N_261,In_570,In_36);
xor U262 (N_262,N_127,In_588);
nor U263 (N_263,N_58,N_173);
or U264 (N_264,In_480,In_262);
nor U265 (N_265,In_600,In_80);
nand U266 (N_266,N_113,In_639);
nor U267 (N_267,In_582,N_14);
nor U268 (N_268,In_117,In_67);
nor U269 (N_269,In_604,N_40);
nor U270 (N_270,In_186,N_105);
nor U271 (N_271,In_1,In_111);
xnor U272 (N_272,N_87,In_732);
and U273 (N_273,In_242,In_645);
and U274 (N_274,In_308,In_182);
and U275 (N_275,N_84,N_135);
or U276 (N_276,In_76,In_608);
nor U277 (N_277,N_51,In_294);
xor U278 (N_278,In_329,In_510);
and U279 (N_279,N_20,In_159);
xnor U280 (N_280,In_740,N_159);
nand U281 (N_281,In_516,In_643);
nor U282 (N_282,In_725,In_420);
xnor U283 (N_283,In_217,N_33);
and U284 (N_284,In_448,In_253);
and U285 (N_285,In_197,In_79);
nand U286 (N_286,N_195,In_507);
xor U287 (N_287,In_664,In_91);
nand U288 (N_288,In_709,N_122);
nor U289 (N_289,In_462,In_94);
or U290 (N_290,N_170,N_1);
nand U291 (N_291,N_137,N_35);
nor U292 (N_292,In_546,In_204);
nand U293 (N_293,N_103,In_554);
xor U294 (N_294,In_276,In_446);
xor U295 (N_295,N_72,In_417);
or U296 (N_296,N_0,N_148);
and U297 (N_297,In_68,N_155);
nor U298 (N_298,In_633,In_726);
or U299 (N_299,In_363,In_395);
nor U300 (N_300,In_704,In_226);
xnor U301 (N_301,In_494,In_153);
nand U302 (N_302,In_710,In_421);
nand U303 (N_303,In_347,In_333);
nor U304 (N_304,N_199,In_715);
or U305 (N_305,In_89,In_646);
xor U306 (N_306,In_477,N_123);
and U307 (N_307,In_718,In_581);
xor U308 (N_308,In_340,N_139);
nor U309 (N_309,In_311,N_128);
nor U310 (N_310,In_618,In_232);
xnor U311 (N_311,N_25,In_599);
and U312 (N_312,In_348,N_193);
nor U313 (N_313,N_18,N_23);
nor U314 (N_314,In_41,In_125);
nor U315 (N_315,In_44,N_138);
or U316 (N_316,N_118,In_345);
nand U317 (N_317,In_640,In_140);
and U318 (N_318,N_76,In_343);
and U319 (N_319,N_145,N_46);
and U320 (N_320,In_306,In_440);
xor U321 (N_321,In_269,In_548);
or U322 (N_322,N_39,N_83);
xnor U323 (N_323,In_365,N_182);
and U324 (N_324,In_183,N_175);
nor U325 (N_325,In_156,In_651);
xnor U326 (N_326,In_575,In_517);
or U327 (N_327,N_198,N_186);
and U328 (N_328,In_621,In_300);
or U329 (N_329,N_10,N_166);
nand U330 (N_330,In_691,In_374);
xnor U331 (N_331,In_325,N_162);
and U332 (N_332,N_187,In_222);
xor U333 (N_333,N_30,In_167);
nor U334 (N_334,In_416,In_352);
nor U335 (N_335,N_131,In_351);
nand U336 (N_336,N_191,N_94);
nand U337 (N_337,In_261,In_33);
xor U338 (N_338,In_383,In_290);
and U339 (N_339,N_157,N_34);
and U340 (N_340,In_430,N_185);
nand U341 (N_341,N_24,N_106);
nor U342 (N_342,In_474,In_619);
or U343 (N_343,N_88,In_88);
or U344 (N_344,In_280,In_493);
nand U345 (N_345,In_172,N_91);
and U346 (N_346,In_121,In_466);
xnor U347 (N_347,In_316,N_184);
or U348 (N_348,In_93,In_6);
and U349 (N_349,In_396,In_729);
nand U350 (N_350,In_401,In_327);
xor U351 (N_351,In_610,N_15);
nand U352 (N_352,In_502,In_165);
xor U353 (N_353,N_49,N_176);
nand U354 (N_354,In_118,In_341);
nor U355 (N_355,In_392,In_419);
and U356 (N_356,In_528,In_239);
nand U357 (N_357,N_52,In_487);
nor U358 (N_358,N_102,In_212);
or U359 (N_359,In_287,In_85);
and U360 (N_360,In_371,N_180);
or U361 (N_361,N_28,In_267);
and U362 (N_362,N_62,In_83);
and U363 (N_363,N_99,In_452);
or U364 (N_364,In_227,N_156);
nand U365 (N_365,In_356,In_611);
and U366 (N_366,In_627,In_86);
nor U367 (N_367,In_674,In_650);
nor U368 (N_368,In_592,N_144);
or U369 (N_369,N_181,N_147);
nand U370 (N_370,N_117,N_120);
or U371 (N_371,N_172,In_15);
nand U372 (N_372,In_378,N_41);
and U373 (N_373,In_565,N_130);
nor U374 (N_374,In_84,N_50);
or U375 (N_375,N_141,In_307);
or U376 (N_376,In_271,N_13);
nand U377 (N_377,N_190,In_730);
and U378 (N_378,N_160,In_124);
nor U379 (N_379,In_65,In_463);
xor U380 (N_380,In_69,In_672);
or U381 (N_381,N_177,In_736);
nand U382 (N_382,N_197,In_3);
xor U383 (N_383,In_0,In_103);
nand U384 (N_384,N_45,In_745);
or U385 (N_385,In_335,N_74);
and U386 (N_386,In_595,In_166);
xnor U387 (N_387,N_189,In_59);
xor U388 (N_388,In_132,N_68);
and U389 (N_389,N_17,N_192);
and U390 (N_390,N_96,In_721);
xnor U391 (N_391,In_641,In_447);
or U392 (N_392,N_6,In_30);
nand U393 (N_393,In_662,In_105);
and U394 (N_394,In_339,In_504);
or U395 (N_395,In_158,In_703);
xor U396 (N_396,In_73,In_66);
and U397 (N_397,In_522,In_134);
nand U398 (N_398,In_367,In_587);
nand U399 (N_399,In_220,In_435);
xnor U400 (N_400,N_247,N_213);
and U401 (N_401,N_374,N_360);
nor U402 (N_402,In_702,N_274);
and U403 (N_403,N_390,N_289);
or U404 (N_404,N_108,N_259);
nor U405 (N_405,N_126,N_281);
nand U406 (N_406,N_350,N_270);
nor U407 (N_407,N_101,In_202);
xor U408 (N_408,N_369,N_233);
xnor U409 (N_409,N_298,N_392);
nor U410 (N_410,N_288,N_262);
nand U411 (N_411,N_376,N_225);
or U412 (N_412,N_286,N_244);
nor U413 (N_413,N_293,In_458);
nand U414 (N_414,In_690,In_224);
or U415 (N_415,N_121,N_248);
nor U416 (N_416,N_69,N_336);
nand U417 (N_417,N_329,N_234);
or U418 (N_418,N_387,In_70);
xnor U419 (N_419,N_321,N_230);
xor U420 (N_420,N_22,In_660);
and U421 (N_421,In_164,In_465);
nor U422 (N_422,N_326,N_90);
or U423 (N_423,N_391,In_699);
nor U424 (N_424,N_375,In_289);
xnor U425 (N_425,N_224,N_171);
or U426 (N_426,N_211,N_165);
xor U427 (N_427,N_240,N_169);
nand U428 (N_428,N_163,In_657);
and U429 (N_429,N_364,N_303);
nor U430 (N_430,N_351,N_379);
nand U431 (N_431,N_82,N_272);
nor U432 (N_432,N_85,N_207);
nand U433 (N_433,N_317,In_247);
nor U434 (N_434,In_349,N_327);
nand U435 (N_435,N_19,N_43);
xnor U436 (N_436,N_276,N_358);
xnor U437 (N_437,In_338,N_280);
nand U438 (N_438,N_178,N_311);
and U439 (N_439,N_365,N_373);
nor U440 (N_440,N_381,In_20);
and U441 (N_441,N_284,N_278);
or U442 (N_442,N_54,N_164);
xor U443 (N_443,N_92,N_323);
nand U444 (N_444,N_218,N_314);
nand U445 (N_445,N_204,N_343);
and U446 (N_446,N_342,N_215);
or U447 (N_447,N_385,In_694);
or U448 (N_448,N_220,N_319);
nor U449 (N_449,N_97,N_330);
or U450 (N_450,N_290,N_217);
nand U451 (N_451,In_590,In_478);
xnor U452 (N_452,N_115,N_236);
and U453 (N_453,N_31,N_356);
xnor U454 (N_454,In_571,N_77);
nand U455 (N_455,N_202,In_353);
and U456 (N_456,N_313,N_151);
xor U457 (N_457,N_203,N_372);
nand U458 (N_458,N_209,In_457);
and U459 (N_459,N_335,N_252);
or U460 (N_460,In_100,N_378);
nor U461 (N_461,N_229,In_578);
nand U462 (N_462,N_370,In_113);
or U463 (N_463,In_254,In_283);
or U464 (N_464,In_576,N_133);
nand U465 (N_465,In_593,N_318);
xnor U466 (N_466,In_152,In_394);
and U467 (N_467,N_383,N_377);
or U468 (N_468,N_271,In_438);
or U469 (N_469,N_332,In_8);
xnor U470 (N_470,N_226,N_299);
xnor U471 (N_471,In_141,N_5);
or U472 (N_472,N_367,N_222);
or U473 (N_473,N_389,N_4);
xor U474 (N_474,N_251,N_346);
xnor U475 (N_475,In_403,N_65);
nand U476 (N_476,N_206,N_216);
and U477 (N_477,In_128,In_514);
nor U478 (N_478,N_107,N_129);
xor U479 (N_479,In_692,N_167);
and U480 (N_480,N_245,N_325);
xor U481 (N_481,N_399,In_615);
xnor U482 (N_482,N_349,N_296);
nand U483 (N_483,N_260,In_568);
and U484 (N_484,N_301,N_70);
nand U485 (N_485,N_305,N_256);
or U486 (N_486,N_306,In_530);
xnor U487 (N_487,N_221,N_297);
and U488 (N_488,N_388,In_190);
nand U489 (N_489,In_626,N_2);
nor U490 (N_490,In_81,N_295);
and U491 (N_491,N_111,N_268);
or U492 (N_492,In_636,In_705);
and U493 (N_493,N_357,In_427);
xnor U494 (N_494,N_380,N_300);
and U495 (N_495,N_397,N_38);
or U496 (N_496,N_183,In_405);
or U497 (N_497,N_324,N_12);
nand U498 (N_498,N_304,In_490);
nand U499 (N_499,In_558,N_361);
xnor U500 (N_500,N_214,In_423);
nor U501 (N_501,In_210,N_36);
nor U502 (N_502,N_75,N_125);
nor U503 (N_503,N_267,In_379);
xnor U504 (N_504,In_606,N_277);
and U505 (N_505,N_347,N_246);
nor U506 (N_506,N_161,N_243);
xnor U507 (N_507,N_258,N_116);
xnor U508 (N_508,N_352,N_261);
xnor U509 (N_509,N_359,In_654);
xor U510 (N_510,N_285,N_253);
and U511 (N_511,N_205,N_60);
and U512 (N_512,N_307,N_344);
xor U513 (N_513,N_283,N_47);
nand U514 (N_514,N_212,N_254);
and U515 (N_515,N_279,In_10);
and U516 (N_516,In_102,N_235);
nand U517 (N_517,N_241,In_257);
or U518 (N_518,N_328,N_263);
or U519 (N_519,In_187,N_264);
or U520 (N_520,In_495,N_396);
xor U521 (N_521,N_292,In_109);
nand U522 (N_522,In_397,In_150);
nor U523 (N_523,N_250,N_340);
nand U524 (N_524,N_368,In_501);
nand U525 (N_525,N_242,In_126);
nand U526 (N_526,N_228,N_322);
nand U527 (N_527,In_114,N_237);
and U528 (N_528,N_42,N_71);
xor U529 (N_529,N_231,N_80);
nand U530 (N_530,N_63,N_273);
nand U531 (N_531,N_227,In_706);
and U532 (N_532,N_238,N_366);
nor U533 (N_533,N_355,N_154);
or U534 (N_534,N_112,N_269);
and U535 (N_535,N_315,In_301);
xnor U536 (N_536,N_27,N_200);
xor U537 (N_537,N_282,N_210);
xor U538 (N_538,N_257,N_333);
nand U539 (N_539,N_208,N_393);
and U540 (N_540,N_232,N_266);
nand U541 (N_541,N_353,N_345);
nor U542 (N_542,In_40,N_339);
nand U543 (N_543,N_21,In_443);
or U544 (N_544,N_362,N_331);
nand U545 (N_545,N_100,N_287);
or U546 (N_546,N_337,N_354);
nor U547 (N_547,N_168,N_255);
or U548 (N_548,In_368,N_341);
nor U549 (N_549,In_625,N_9);
nand U550 (N_550,In_667,In_485);
xnor U551 (N_551,In_245,N_294);
nand U552 (N_552,In_521,N_158);
and U553 (N_553,N_398,In_631);
or U554 (N_554,N_384,In_22);
xor U555 (N_555,N_265,N_174);
and U556 (N_556,N_275,In_693);
xnor U557 (N_557,In_270,N_66);
and U558 (N_558,N_310,N_371);
nor U559 (N_559,In_549,N_395);
nor U560 (N_560,N_386,In_665);
xnor U561 (N_561,N_302,N_394);
and U562 (N_562,N_363,In_616);
or U563 (N_563,In_211,N_219);
nand U564 (N_564,In_176,N_146);
and U565 (N_565,In_711,In_364);
or U566 (N_566,N_348,N_55);
nand U567 (N_567,N_309,N_316);
and U568 (N_568,N_249,N_320);
xor U569 (N_569,N_201,N_308);
nor U570 (N_570,N_291,N_239);
and U571 (N_571,N_382,N_338);
nor U572 (N_572,N_223,N_334);
and U573 (N_573,N_140,In_112);
nand U574 (N_574,N_59,N_312);
nor U575 (N_575,In_211,In_112);
or U576 (N_576,In_126,In_397);
and U577 (N_577,N_80,N_214);
and U578 (N_578,N_398,N_174);
or U579 (N_579,In_112,N_158);
xnor U580 (N_580,N_171,N_387);
and U581 (N_581,In_631,N_280);
and U582 (N_582,In_112,N_281);
or U583 (N_583,N_295,N_335);
nand U584 (N_584,In_657,N_293);
nand U585 (N_585,N_351,N_385);
nor U586 (N_586,N_344,N_294);
xor U587 (N_587,In_224,N_22);
xor U588 (N_588,In_301,In_405);
or U589 (N_589,N_395,N_229);
and U590 (N_590,N_323,N_312);
or U591 (N_591,N_125,In_353);
xor U592 (N_592,N_225,In_485);
xor U593 (N_593,N_385,N_60);
nand U594 (N_594,N_126,N_265);
or U595 (N_595,N_364,N_222);
nor U596 (N_596,N_297,N_382);
nor U597 (N_597,In_397,In_247);
xor U598 (N_598,In_109,N_290);
and U599 (N_599,N_356,In_10);
and U600 (N_600,N_443,N_538);
nand U601 (N_601,N_556,N_473);
and U602 (N_602,N_433,N_578);
or U603 (N_603,N_497,N_533);
and U604 (N_604,N_498,N_494);
nor U605 (N_605,N_524,N_535);
nand U606 (N_606,N_579,N_424);
or U607 (N_607,N_594,N_401);
or U608 (N_608,N_503,N_515);
nor U609 (N_609,N_427,N_548);
xor U610 (N_610,N_451,N_508);
nand U611 (N_611,N_517,N_537);
nor U612 (N_612,N_452,N_575);
and U613 (N_613,N_410,N_532);
nor U614 (N_614,N_567,N_431);
or U615 (N_615,N_500,N_437);
and U616 (N_616,N_585,N_554);
nand U617 (N_617,N_423,N_471);
nand U618 (N_618,N_593,N_476);
nor U619 (N_619,N_408,N_597);
xnor U620 (N_620,N_481,N_445);
xnor U621 (N_621,N_463,N_415);
nor U622 (N_622,N_523,N_447);
or U623 (N_623,N_572,N_510);
and U624 (N_624,N_429,N_480);
nor U625 (N_625,N_436,N_435);
and U626 (N_626,N_495,N_422);
nand U627 (N_627,N_574,N_417);
nand U628 (N_628,N_441,N_465);
and U629 (N_629,N_453,N_553);
and U630 (N_630,N_490,N_496);
and U631 (N_631,N_582,N_565);
nor U632 (N_632,N_409,N_407);
or U633 (N_633,N_552,N_581);
or U634 (N_634,N_507,N_428);
or U635 (N_635,N_584,N_400);
or U636 (N_636,N_466,N_491);
or U637 (N_637,N_539,N_521);
and U638 (N_638,N_506,N_559);
and U639 (N_639,N_477,N_505);
and U640 (N_640,N_486,N_528);
xnor U641 (N_641,N_499,N_430);
xor U642 (N_642,N_446,N_432);
or U643 (N_643,N_545,N_529);
and U644 (N_644,N_444,N_599);
or U645 (N_645,N_542,N_464);
or U646 (N_646,N_595,N_440);
xnor U647 (N_647,N_478,N_461);
or U648 (N_648,N_544,N_531);
nand U649 (N_649,N_512,N_411);
nor U650 (N_650,N_536,N_406);
nand U651 (N_651,N_571,N_525);
or U652 (N_652,N_576,N_588);
nor U653 (N_653,N_566,N_475);
xor U654 (N_654,N_413,N_419);
nand U655 (N_655,N_509,N_470);
or U656 (N_656,N_418,N_561);
xnor U657 (N_657,N_540,N_558);
nor U658 (N_658,N_454,N_434);
or U659 (N_659,N_484,N_448);
nor U660 (N_660,N_560,N_442);
or U661 (N_661,N_522,N_569);
nor U662 (N_662,N_459,N_472);
nor U663 (N_663,N_489,N_402);
or U664 (N_664,N_449,N_483);
or U665 (N_665,N_577,N_564);
xnor U666 (N_666,N_421,N_511);
xnor U667 (N_667,N_412,N_462);
and U668 (N_668,N_426,N_530);
and U669 (N_669,N_439,N_557);
and U670 (N_670,N_546,N_555);
xnor U671 (N_671,N_457,N_455);
nand U672 (N_672,N_482,N_520);
or U673 (N_673,N_562,N_590);
or U674 (N_674,N_583,N_416);
or U675 (N_675,N_420,N_550);
or U676 (N_676,N_403,N_516);
and U677 (N_677,N_570,N_519);
and U678 (N_678,N_501,N_405);
nand U679 (N_679,N_547,N_596);
nor U680 (N_680,N_474,N_549);
nor U681 (N_681,N_504,N_527);
xnor U682 (N_682,N_450,N_580);
or U683 (N_683,N_493,N_438);
nor U684 (N_684,N_456,N_460);
xor U685 (N_685,N_587,N_414);
xor U686 (N_686,N_467,N_479);
nor U687 (N_687,N_518,N_589);
xnor U688 (N_688,N_573,N_468);
and U689 (N_689,N_485,N_568);
xnor U690 (N_690,N_425,N_543);
nor U691 (N_691,N_592,N_502);
xnor U692 (N_692,N_404,N_563);
nand U693 (N_693,N_586,N_598);
and U694 (N_694,N_541,N_492);
or U695 (N_695,N_526,N_591);
xor U696 (N_696,N_551,N_469);
xnor U697 (N_697,N_487,N_534);
nor U698 (N_698,N_514,N_458);
xor U699 (N_699,N_488,N_513);
xor U700 (N_700,N_515,N_528);
nand U701 (N_701,N_562,N_438);
xnor U702 (N_702,N_491,N_414);
nand U703 (N_703,N_545,N_434);
and U704 (N_704,N_514,N_497);
xnor U705 (N_705,N_467,N_590);
nor U706 (N_706,N_441,N_500);
xor U707 (N_707,N_524,N_413);
xnor U708 (N_708,N_530,N_445);
nor U709 (N_709,N_411,N_589);
nand U710 (N_710,N_500,N_552);
or U711 (N_711,N_419,N_412);
xor U712 (N_712,N_531,N_426);
nand U713 (N_713,N_545,N_413);
or U714 (N_714,N_543,N_570);
nand U715 (N_715,N_482,N_481);
xor U716 (N_716,N_405,N_429);
or U717 (N_717,N_477,N_446);
and U718 (N_718,N_524,N_464);
nor U719 (N_719,N_462,N_531);
nand U720 (N_720,N_411,N_448);
xor U721 (N_721,N_505,N_502);
xnor U722 (N_722,N_581,N_445);
nand U723 (N_723,N_414,N_453);
xnor U724 (N_724,N_429,N_582);
nand U725 (N_725,N_480,N_598);
xor U726 (N_726,N_597,N_455);
and U727 (N_727,N_584,N_575);
nor U728 (N_728,N_554,N_415);
or U729 (N_729,N_525,N_418);
nand U730 (N_730,N_509,N_514);
or U731 (N_731,N_439,N_406);
or U732 (N_732,N_427,N_492);
nand U733 (N_733,N_572,N_580);
nor U734 (N_734,N_416,N_465);
nor U735 (N_735,N_557,N_501);
nand U736 (N_736,N_564,N_581);
or U737 (N_737,N_433,N_477);
and U738 (N_738,N_526,N_483);
nand U739 (N_739,N_516,N_580);
or U740 (N_740,N_567,N_454);
xor U741 (N_741,N_535,N_420);
xnor U742 (N_742,N_449,N_537);
and U743 (N_743,N_594,N_436);
xor U744 (N_744,N_580,N_556);
nand U745 (N_745,N_424,N_574);
and U746 (N_746,N_431,N_529);
nand U747 (N_747,N_424,N_477);
and U748 (N_748,N_477,N_544);
nand U749 (N_749,N_532,N_480);
nor U750 (N_750,N_401,N_463);
nand U751 (N_751,N_477,N_441);
nand U752 (N_752,N_570,N_473);
nand U753 (N_753,N_488,N_556);
or U754 (N_754,N_538,N_541);
xnor U755 (N_755,N_488,N_451);
nand U756 (N_756,N_583,N_422);
xor U757 (N_757,N_485,N_480);
xor U758 (N_758,N_522,N_446);
xnor U759 (N_759,N_553,N_415);
or U760 (N_760,N_446,N_584);
nor U761 (N_761,N_554,N_425);
xor U762 (N_762,N_519,N_486);
xor U763 (N_763,N_450,N_508);
nand U764 (N_764,N_518,N_525);
or U765 (N_765,N_497,N_434);
or U766 (N_766,N_467,N_400);
nor U767 (N_767,N_520,N_503);
or U768 (N_768,N_469,N_431);
or U769 (N_769,N_440,N_426);
xnor U770 (N_770,N_550,N_500);
nor U771 (N_771,N_527,N_518);
nand U772 (N_772,N_566,N_580);
xnor U773 (N_773,N_540,N_433);
and U774 (N_774,N_538,N_537);
xor U775 (N_775,N_441,N_462);
xnor U776 (N_776,N_509,N_471);
nor U777 (N_777,N_404,N_516);
and U778 (N_778,N_495,N_573);
xor U779 (N_779,N_481,N_483);
nand U780 (N_780,N_598,N_487);
xnor U781 (N_781,N_444,N_462);
nor U782 (N_782,N_529,N_503);
and U783 (N_783,N_490,N_472);
xor U784 (N_784,N_560,N_404);
nor U785 (N_785,N_556,N_546);
nand U786 (N_786,N_402,N_553);
and U787 (N_787,N_497,N_474);
nand U788 (N_788,N_533,N_514);
nand U789 (N_789,N_502,N_445);
nand U790 (N_790,N_518,N_457);
nor U791 (N_791,N_452,N_502);
and U792 (N_792,N_458,N_484);
and U793 (N_793,N_403,N_537);
nand U794 (N_794,N_479,N_553);
and U795 (N_795,N_587,N_455);
and U796 (N_796,N_436,N_556);
xor U797 (N_797,N_559,N_513);
nor U798 (N_798,N_415,N_495);
nor U799 (N_799,N_442,N_579);
nor U800 (N_800,N_783,N_735);
nand U801 (N_801,N_630,N_770);
or U802 (N_802,N_754,N_622);
and U803 (N_803,N_767,N_733);
or U804 (N_804,N_796,N_711);
xnor U805 (N_805,N_680,N_659);
xnor U806 (N_806,N_746,N_647);
and U807 (N_807,N_641,N_776);
and U808 (N_808,N_696,N_632);
or U809 (N_809,N_657,N_759);
nand U810 (N_810,N_743,N_740);
nand U811 (N_811,N_737,N_683);
or U812 (N_812,N_753,N_712);
or U813 (N_813,N_721,N_701);
xor U814 (N_814,N_631,N_739);
nor U815 (N_815,N_706,N_797);
or U816 (N_816,N_663,N_628);
nor U817 (N_817,N_655,N_786);
or U818 (N_818,N_685,N_728);
or U819 (N_819,N_602,N_778);
and U820 (N_820,N_670,N_695);
and U821 (N_821,N_658,N_744);
nand U822 (N_822,N_763,N_742);
xnor U823 (N_823,N_722,N_620);
and U824 (N_824,N_633,N_629);
and U825 (N_825,N_707,N_784);
nor U826 (N_826,N_665,N_604);
nor U827 (N_827,N_757,N_718);
and U828 (N_828,N_668,N_758);
nor U829 (N_829,N_713,N_645);
xnor U830 (N_830,N_619,N_644);
nand U831 (N_831,N_724,N_760);
nor U832 (N_832,N_664,N_666);
or U833 (N_833,N_790,N_764);
nand U834 (N_834,N_719,N_667);
or U835 (N_835,N_799,N_793);
xor U836 (N_836,N_769,N_606);
nor U837 (N_837,N_725,N_714);
nor U838 (N_838,N_601,N_708);
or U839 (N_839,N_734,N_678);
xnor U840 (N_840,N_794,N_675);
xnor U841 (N_841,N_652,N_773);
and U842 (N_842,N_691,N_771);
nand U843 (N_843,N_747,N_600);
xnor U844 (N_844,N_603,N_736);
nor U845 (N_845,N_608,N_727);
or U846 (N_846,N_745,N_698);
nand U847 (N_847,N_792,N_661);
nor U848 (N_848,N_650,N_690);
nand U849 (N_849,N_723,N_779);
and U850 (N_850,N_774,N_654);
xnor U851 (N_851,N_781,N_780);
or U852 (N_852,N_677,N_703);
nor U853 (N_853,N_750,N_688);
nand U854 (N_854,N_689,N_626);
or U855 (N_855,N_787,N_611);
xnor U856 (N_856,N_791,N_637);
or U857 (N_857,N_612,N_738);
or U858 (N_858,N_653,N_648);
nand U859 (N_859,N_613,N_752);
xor U860 (N_860,N_642,N_762);
and U861 (N_861,N_682,N_662);
nor U862 (N_862,N_741,N_715);
xor U863 (N_863,N_704,N_636);
nand U864 (N_864,N_616,N_649);
xor U865 (N_865,N_765,N_673);
or U866 (N_866,N_614,N_639);
xor U867 (N_867,N_748,N_785);
nand U868 (N_868,N_635,N_699);
xor U869 (N_869,N_700,N_732);
nand U870 (N_870,N_756,N_795);
nor U871 (N_871,N_772,N_646);
xnor U872 (N_872,N_717,N_610);
and U873 (N_873,N_720,N_609);
nor U874 (N_874,N_615,N_694);
or U875 (N_875,N_782,N_618);
nand U876 (N_876,N_702,N_621);
xnor U877 (N_877,N_798,N_651);
xnor U878 (N_878,N_768,N_709);
xnor U879 (N_879,N_617,N_607);
or U880 (N_880,N_755,N_729);
nand U881 (N_881,N_766,N_624);
xor U882 (N_882,N_686,N_679);
nor U883 (N_883,N_643,N_692);
xor U884 (N_884,N_761,N_627);
nor U885 (N_885,N_669,N_705);
xnor U886 (N_886,N_605,N_681);
or U887 (N_887,N_726,N_623);
nand U888 (N_888,N_749,N_710);
nand U889 (N_889,N_638,N_716);
nor U890 (N_890,N_788,N_731);
xnor U891 (N_891,N_676,N_672);
nor U892 (N_892,N_671,N_789);
xnor U893 (N_893,N_684,N_730);
and U894 (N_894,N_751,N_634);
or U895 (N_895,N_625,N_660);
xor U896 (N_896,N_697,N_656);
nor U897 (N_897,N_777,N_775);
nor U898 (N_898,N_674,N_693);
nor U899 (N_899,N_640,N_687);
or U900 (N_900,N_759,N_721);
nor U901 (N_901,N_790,N_600);
nand U902 (N_902,N_753,N_685);
nor U903 (N_903,N_657,N_722);
xnor U904 (N_904,N_650,N_660);
nand U905 (N_905,N_764,N_612);
xnor U906 (N_906,N_637,N_638);
nand U907 (N_907,N_768,N_631);
xor U908 (N_908,N_672,N_602);
or U909 (N_909,N_703,N_741);
nand U910 (N_910,N_741,N_684);
xnor U911 (N_911,N_678,N_796);
nand U912 (N_912,N_750,N_631);
nor U913 (N_913,N_628,N_602);
xor U914 (N_914,N_695,N_786);
and U915 (N_915,N_658,N_751);
and U916 (N_916,N_629,N_728);
nand U917 (N_917,N_711,N_734);
xnor U918 (N_918,N_796,N_697);
xnor U919 (N_919,N_779,N_780);
nor U920 (N_920,N_751,N_769);
xnor U921 (N_921,N_786,N_761);
or U922 (N_922,N_638,N_693);
or U923 (N_923,N_783,N_797);
or U924 (N_924,N_769,N_651);
and U925 (N_925,N_734,N_752);
and U926 (N_926,N_717,N_753);
xor U927 (N_927,N_784,N_710);
or U928 (N_928,N_773,N_672);
and U929 (N_929,N_769,N_744);
nor U930 (N_930,N_754,N_686);
nor U931 (N_931,N_778,N_742);
nor U932 (N_932,N_664,N_629);
nor U933 (N_933,N_711,N_609);
nor U934 (N_934,N_610,N_711);
nand U935 (N_935,N_765,N_651);
and U936 (N_936,N_682,N_655);
nor U937 (N_937,N_673,N_799);
or U938 (N_938,N_691,N_723);
nand U939 (N_939,N_627,N_718);
or U940 (N_940,N_743,N_638);
nand U941 (N_941,N_791,N_695);
or U942 (N_942,N_675,N_789);
nor U943 (N_943,N_788,N_615);
xnor U944 (N_944,N_799,N_609);
or U945 (N_945,N_757,N_624);
nor U946 (N_946,N_786,N_728);
xor U947 (N_947,N_656,N_650);
nor U948 (N_948,N_656,N_776);
or U949 (N_949,N_726,N_647);
or U950 (N_950,N_682,N_737);
or U951 (N_951,N_723,N_618);
nor U952 (N_952,N_624,N_706);
nand U953 (N_953,N_636,N_623);
xor U954 (N_954,N_624,N_782);
nand U955 (N_955,N_756,N_760);
nand U956 (N_956,N_778,N_730);
xnor U957 (N_957,N_630,N_652);
and U958 (N_958,N_601,N_716);
and U959 (N_959,N_688,N_648);
nand U960 (N_960,N_604,N_781);
xnor U961 (N_961,N_673,N_658);
and U962 (N_962,N_756,N_792);
or U963 (N_963,N_794,N_765);
nor U964 (N_964,N_632,N_608);
xnor U965 (N_965,N_693,N_733);
and U966 (N_966,N_707,N_719);
and U967 (N_967,N_674,N_637);
nor U968 (N_968,N_624,N_653);
or U969 (N_969,N_708,N_695);
nand U970 (N_970,N_711,N_700);
or U971 (N_971,N_708,N_607);
xnor U972 (N_972,N_659,N_708);
nand U973 (N_973,N_707,N_745);
or U974 (N_974,N_790,N_683);
xnor U975 (N_975,N_730,N_692);
nor U976 (N_976,N_778,N_607);
and U977 (N_977,N_646,N_787);
xnor U978 (N_978,N_613,N_718);
nand U979 (N_979,N_780,N_653);
nand U980 (N_980,N_669,N_782);
nand U981 (N_981,N_744,N_792);
or U982 (N_982,N_674,N_785);
nand U983 (N_983,N_740,N_781);
or U984 (N_984,N_650,N_782);
nand U985 (N_985,N_639,N_788);
or U986 (N_986,N_755,N_757);
and U987 (N_987,N_785,N_760);
nand U988 (N_988,N_771,N_725);
and U989 (N_989,N_756,N_798);
xor U990 (N_990,N_656,N_633);
and U991 (N_991,N_648,N_607);
xor U992 (N_992,N_792,N_643);
xnor U993 (N_993,N_680,N_622);
nor U994 (N_994,N_648,N_604);
or U995 (N_995,N_654,N_786);
nand U996 (N_996,N_658,N_729);
or U997 (N_997,N_786,N_771);
or U998 (N_998,N_654,N_639);
nor U999 (N_999,N_776,N_775);
nand U1000 (N_1000,N_889,N_803);
nor U1001 (N_1001,N_818,N_858);
nand U1002 (N_1002,N_888,N_817);
nand U1003 (N_1003,N_808,N_993);
xnor U1004 (N_1004,N_978,N_981);
nand U1005 (N_1005,N_963,N_855);
or U1006 (N_1006,N_827,N_838);
nand U1007 (N_1007,N_813,N_931);
or U1008 (N_1008,N_939,N_955);
xor U1009 (N_1009,N_899,N_936);
or U1010 (N_1010,N_929,N_859);
nand U1011 (N_1011,N_850,N_924);
nand U1012 (N_1012,N_962,N_994);
or U1013 (N_1013,N_947,N_904);
xor U1014 (N_1014,N_999,N_917);
nand U1015 (N_1015,N_988,N_953);
or U1016 (N_1016,N_986,N_845);
or U1017 (N_1017,N_890,N_852);
xnor U1018 (N_1018,N_847,N_857);
nand U1019 (N_1019,N_842,N_892);
xor U1020 (N_1020,N_826,N_809);
or U1021 (N_1021,N_943,N_995);
nand U1022 (N_1022,N_912,N_985);
nand U1023 (N_1023,N_983,N_913);
nand U1024 (N_1024,N_844,N_928);
and U1025 (N_1025,N_834,N_841);
nor U1026 (N_1026,N_865,N_863);
and U1027 (N_1027,N_848,N_991);
or U1028 (N_1028,N_829,N_860);
or U1029 (N_1029,N_868,N_854);
xnor U1030 (N_1030,N_856,N_862);
and U1031 (N_1031,N_837,N_887);
nor U1032 (N_1032,N_902,N_949);
and U1033 (N_1033,N_935,N_875);
and U1034 (N_1034,N_934,N_884);
nand U1035 (N_1035,N_896,N_815);
xor U1036 (N_1036,N_940,N_980);
and U1037 (N_1037,N_982,N_825);
and U1038 (N_1038,N_846,N_926);
nand U1039 (N_1039,N_833,N_956);
nor U1040 (N_1040,N_977,N_918);
nor U1041 (N_1041,N_901,N_897);
or U1042 (N_1042,N_873,N_973);
nor U1043 (N_1043,N_882,N_861);
and U1044 (N_1044,N_804,N_972);
nand U1045 (N_1045,N_922,N_961);
nand U1046 (N_1046,N_911,N_971);
or U1047 (N_1047,N_945,N_946);
nand U1048 (N_1048,N_895,N_823);
and U1049 (N_1049,N_867,N_885);
nor U1050 (N_1050,N_828,N_941);
nor U1051 (N_1051,N_874,N_877);
and U1052 (N_1052,N_967,N_819);
and U1053 (N_1053,N_948,N_974);
and U1054 (N_1054,N_881,N_969);
nor U1055 (N_1055,N_959,N_814);
or U1056 (N_1056,N_965,N_851);
or U1057 (N_1057,N_968,N_822);
nor U1058 (N_1058,N_938,N_806);
or U1059 (N_1059,N_870,N_871);
and U1060 (N_1060,N_800,N_942);
xnor U1061 (N_1061,N_836,N_869);
nand U1062 (N_1062,N_970,N_883);
nor U1063 (N_1063,N_908,N_866);
or U1064 (N_1064,N_921,N_905);
and U1065 (N_1065,N_821,N_950);
nor U1066 (N_1066,N_954,N_960);
xor U1067 (N_1067,N_849,N_923);
or U1068 (N_1068,N_886,N_805);
nand U1069 (N_1069,N_906,N_996);
or U1070 (N_1070,N_932,N_900);
xnor U1071 (N_1071,N_878,N_964);
xor U1072 (N_1072,N_820,N_835);
or U1073 (N_1073,N_952,N_880);
nand U1074 (N_1074,N_801,N_990);
nor U1075 (N_1075,N_802,N_984);
xnor U1076 (N_1076,N_832,N_930);
xnor U1077 (N_1077,N_864,N_812);
or U1078 (N_1078,N_810,N_976);
xor U1079 (N_1079,N_987,N_891);
nand U1080 (N_1080,N_933,N_920);
nand U1081 (N_1081,N_903,N_915);
xor U1082 (N_1082,N_840,N_927);
or U1083 (N_1083,N_830,N_937);
xnor U1084 (N_1084,N_989,N_958);
xnor U1085 (N_1085,N_909,N_879);
xnor U1086 (N_1086,N_839,N_992);
xor U1087 (N_1087,N_919,N_944);
xor U1088 (N_1088,N_957,N_876);
and U1089 (N_1089,N_816,N_811);
nand U1090 (N_1090,N_951,N_898);
nor U1091 (N_1091,N_843,N_853);
and U1092 (N_1092,N_997,N_975);
or U1093 (N_1093,N_998,N_910);
nand U1094 (N_1094,N_916,N_979);
xor U1095 (N_1095,N_824,N_966);
xor U1096 (N_1096,N_831,N_807);
xor U1097 (N_1097,N_907,N_914);
xnor U1098 (N_1098,N_893,N_925);
xor U1099 (N_1099,N_894,N_872);
nor U1100 (N_1100,N_930,N_836);
xnor U1101 (N_1101,N_979,N_826);
and U1102 (N_1102,N_858,N_852);
xnor U1103 (N_1103,N_915,N_912);
and U1104 (N_1104,N_929,N_806);
and U1105 (N_1105,N_860,N_995);
xnor U1106 (N_1106,N_875,N_930);
or U1107 (N_1107,N_816,N_824);
nand U1108 (N_1108,N_845,N_919);
nand U1109 (N_1109,N_877,N_902);
xnor U1110 (N_1110,N_836,N_922);
nand U1111 (N_1111,N_982,N_850);
xor U1112 (N_1112,N_891,N_963);
xor U1113 (N_1113,N_911,N_885);
and U1114 (N_1114,N_879,N_928);
or U1115 (N_1115,N_974,N_899);
and U1116 (N_1116,N_834,N_890);
nand U1117 (N_1117,N_823,N_814);
nand U1118 (N_1118,N_920,N_812);
or U1119 (N_1119,N_960,N_813);
or U1120 (N_1120,N_898,N_901);
nor U1121 (N_1121,N_860,N_875);
nor U1122 (N_1122,N_950,N_968);
nor U1123 (N_1123,N_838,N_806);
nor U1124 (N_1124,N_887,N_868);
and U1125 (N_1125,N_968,N_883);
nand U1126 (N_1126,N_950,N_851);
and U1127 (N_1127,N_851,N_903);
nor U1128 (N_1128,N_984,N_846);
or U1129 (N_1129,N_924,N_973);
xnor U1130 (N_1130,N_854,N_949);
xnor U1131 (N_1131,N_939,N_907);
nor U1132 (N_1132,N_896,N_957);
nor U1133 (N_1133,N_893,N_926);
xnor U1134 (N_1134,N_852,N_968);
nor U1135 (N_1135,N_809,N_901);
nand U1136 (N_1136,N_931,N_993);
xnor U1137 (N_1137,N_845,N_824);
nand U1138 (N_1138,N_869,N_903);
nor U1139 (N_1139,N_838,N_968);
xnor U1140 (N_1140,N_962,N_807);
nor U1141 (N_1141,N_978,N_849);
or U1142 (N_1142,N_914,N_938);
nor U1143 (N_1143,N_854,N_927);
nor U1144 (N_1144,N_899,N_966);
xnor U1145 (N_1145,N_959,N_907);
xor U1146 (N_1146,N_991,N_983);
and U1147 (N_1147,N_862,N_997);
nor U1148 (N_1148,N_919,N_851);
nand U1149 (N_1149,N_825,N_890);
nor U1150 (N_1150,N_927,N_822);
nor U1151 (N_1151,N_843,N_833);
nand U1152 (N_1152,N_884,N_979);
nor U1153 (N_1153,N_999,N_957);
and U1154 (N_1154,N_894,N_975);
nand U1155 (N_1155,N_834,N_875);
and U1156 (N_1156,N_958,N_862);
or U1157 (N_1157,N_874,N_855);
xor U1158 (N_1158,N_895,N_908);
nor U1159 (N_1159,N_804,N_876);
xor U1160 (N_1160,N_844,N_874);
nor U1161 (N_1161,N_998,N_951);
xnor U1162 (N_1162,N_996,N_985);
nor U1163 (N_1163,N_911,N_831);
nor U1164 (N_1164,N_949,N_967);
xor U1165 (N_1165,N_941,N_836);
or U1166 (N_1166,N_886,N_912);
and U1167 (N_1167,N_926,N_875);
or U1168 (N_1168,N_920,N_852);
nand U1169 (N_1169,N_874,N_978);
nor U1170 (N_1170,N_986,N_827);
and U1171 (N_1171,N_900,N_822);
and U1172 (N_1172,N_874,N_800);
nand U1173 (N_1173,N_932,N_814);
nand U1174 (N_1174,N_963,N_832);
and U1175 (N_1175,N_851,N_866);
nand U1176 (N_1176,N_811,N_969);
nor U1177 (N_1177,N_919,N_913);
nand U1178 (N_1178,N_899,N_983);
xor U1179 (N_1179,N_851,N_893);
nor U1180 (N_1180,N_983,N_921);
nor U1181 (N_1181,N_943,N_887);
nand U1182 (N_1182,N_877,N_933);
nand U1183 (N_1183,N_941,N_877);
or U1184 (N_1184,N_885,N_869);
or U1185 (N_1185,N_915,N_997);
or U1186 (N_1186,N_873,N_995);
and U1187 (N_1187,N_965,N_815);
nand U1188 (N_1188,N_962,N_806);
and U1189 (N_1189,N_811,N_994);
nor U1190 (N_1190,N_838,N_948);
and U1191 (N_1191,N_839,N_993);
or U1192 (N_1192,N_986,N_916);
nor U1193 (N_1193,N_998,N_899);
xnor U1194 (N_1194,N_868,N_843);
nor U1195 (N_1195,N_902,N_926);
xor U1196 (N_1196,N_841,N_892);
xor U1197 (N_1197,N_835,N_849);
nor U1198 (N_1198,N_955,N_808);
and U1199 (N_1199,N_895,N_828);
xnor U1200 (N_1200,N_1032,N_1193);
and U1201 (N_1201,N_1077,N_1121);
and U1202 (N_1202,N_1008,N_1148);
nor U1203 (N_1203,N_1026,N_1183);
nand U1204 (N_1204,N_1015,N_1082);
xor U1205 (N_1205,N_1091,N_1150);
xor U1206 (N_1206,N_1034,N_1056);
and U1207 (N_1207,N_1162,N_1035);
or U1208 (N_1208,N_1063,N_1003);
or U1209 (N_1209,N_1068,N_1181);
and U1210 (N_1210,N_1112,N_1159);
or U1211 (N_1211,N_1095,N_1152);
xor U1212 (N_1212,N_1009,N_1149);
xor U1213 (N_1213,N_1027,N_1136);
xor U1214 (N_1214,N_1055,N_1129);
and U1215 (N_1215,N_1018,N_1065);
nor U1216 (N_1216,N_1040,N_1151);
nand U1217 (N_1217,N_1191,N_1021);
nand U1218 (N_1218,N_1146,N_1099);
nand U1219 (N_1219,N_1016,N_1156);
nor U1220 (N_1220,N_1022,N_1199);
xnor U1221 (N_1221,N_1154,N_1143);
or U1222 (N_1222,N_1005,N_1142);
nand U1223 (N_1223,N_1180,N_1103);
nor U1224 (N_1224,N_1002,N_1165);
xnor U1225 (N_1225,N_1036,N_1024);
or U1226 (N_1226,N_1107,N_1025);
or U1227 (N_1227,N_1189,N_1190);
nor U1228 (N_1228,N_1141,N_1088);
or U1229 (N_1229,N_1116,N_1147);
nand U1230 (N_1230,N_1120,N_1064);
nand U1231 (N_1231,N_1161,N_1131);
or U1232 (N_1232,N_1019,N_1124);
xnor U1233 (N_1233,N_1047,N_1145);
xor U1234 (N_1234,N_1080,N_1031);
nand U1235 (N_1235,N_1086,N_1113);
nand U1236 (N_1236,N_1188,N_1052);
xnor U1237 (N_1237,N_1172,N_1074);
nor U1238 (N_1238,N_1090,N_1184);
xor U1239 (N_1239,N_1072,N_1114);
xor U1240 (N_1240,N_1039,N_1109);
nand U1241 (N_1241,N_1071,N_1087);
and U1242 (N_1242,N_1157,N_1051);
and U1243 (N_1243,N_1057,N_1023);
nand U1244 (N_1244,N_1169,N_1198);
or U1245 (N_1245,N_1079,N_1028);
nand U1246 (N_1246,N_1158,N_1066);
xnor U1247 (N_1247,N_1128,N_1135);
xnor U1248 (N_1248,N_1166,N_1173);
and U1249 (N_1249,N_1105,N_1175);
xnor U1250 (N_1250,N_1139,N_1186);
and U1251 (N_1251,N_1177,N_1043);
and U1252 (N_1252,N_1012,N_1101);
nor U1253 (N_1253,N_1176,N_1178);
and U1254 (N_1254,N_1140,N_1168);
xor U1255 (N_1255,N_1060,N_1134);
nor U1256 (N_1256,N_1182,N_1167);
and U1257 (N_1257,N_1123,N_1118);
or U1258 (N_1258,N_1174,N_1075);
or U1259 (N_1259,N_1098,N_1010);
nand U1260 (N_1260,N_1069,N_1196);
nor U1261 (N_1261,N_1092,N_1104);
and U1262 (N_1262,N_1138,N_1119);
nor U1263 (N_1263,N_1062,N_1187);
xnor U1264 (N_1264,N_1106,N_1110);
xnor U1265 (N_1265,N_1179,N_1155);
and U1266 (N_1266,N_1042,N_1126);
and U1267 (N_1267,N_1073,N_1164);
nor U1268 (N_1268,N_1058,N_1011);
and U1269 (N_1269,N_1197,N_1050);
and U1270 (N_1270,N_1096,N_1102);
nand U1271 (N_1271,N_1001,N_1030);
nor U1272 (N_1272,N_1070,N_1033);
nor U1273 (N_1273,N_1194,N_1000);
nand U1274 (N_1274,N_1037,N_1017);
nand U1275 (N_1275,N_1130,N_1045);
or U1276 (N_1276,N_1100,N_1132);
nor U1277 (N_1277,N_1048,N_1163);
nand U1278 (N_1278,N_1171,N_1133);
xor U1279 (N_1279,N_1085,N_1144);
nand U1280 (N_1280,N_1038,N_1195);
xnor U1281 (N_1281,N_1125,N_1059);
nand U1282 (N_1282,N_1007,N_1004);
nor U1283 (N_1283,N_1094,N_1115);
nor U1284 (N_1284,N_1006,N_1046);
nor U1285 (N_1285,N_1067,N_1122);
nand U1286 (N_1286,N_1137,N_1097);
or U1287 (N_1287,N_1020,N_1081);
nor U1288 (N_1288,N_1054,N_1083);
or U1289 (N_1289,N_1061,N_1041);
nand U1290 (N_1290,N_1084,N_1117);
and U1291 (N_1291,N_1078,N_1049);
nor U1292 (N_1292,N_1153,N_1053);
xnor U1293 (N_1293,N_1013,N_1044);
and U1294 (N_1294,N_1160,N_1127);
xnor U1295 (N_1295,N_1108,N_1111);
xnor U1296 (N_1296,N_1192,N_1185);
nor U1297 (N_1297,N_1170,N_1089);
xnor U1298 (N_1298,N_1029,N_1076);
nor U1299 (N_1299,N_1093,N_1014);
nor U1300 (N_1300,N_1180,N_1104);
nor U1301 (N_1301,N_1031,N_1097);
nor U1302 (N_1302,N_1171,N_1090);
nand U1303 (N_1303,N_1190,N_1197);
and U1304 (N_1304,N_1028,N_1064);
xnor U1305 (N_1305,N_1178,N_1185);
nor U1306 (N_1306,N_1198,N_1086);
nor U1307 (N_1307,N_1124,N_1078);
xor U1308 (N_1308,N_1064,N_1003);
nand U1309 (N_1309,N_1164,N_1116);
xor U1310 (N_1310,N_1042,N_1111);
xor U1311 (N_1311,N_1167,N_1029);
and U1312 (N_1312,N_1117,N_1042);
nor U1313 (N_1313,N_1023,N_1015);
or U1314 (N_1314,N_1176,N_1022);
nand U1315 (N_1315,N_1118,N_1163);
nor U1316 (N_1316,N_1176,N_1155);
nand U1317 (N_1317,N_1122,N_1114);
and U1318 (N_1318,N_1054,N_1135);
and U1319 (N_1319,N_1004,N_1074);
and U1320 (N_1320,N_1165,N_1043);
or U1321 (N_1321,N_1137,N_1153);
xnor U1322 (N_1322,N_1098,N_1063);
nand U1323 (N_1323,N_1173,N_1021);
nand U1324 (N_1324,N_1117,N_1078);
or U1325 (N_1325,N_1142,N_1095);
nor U1326 (N_1326,N_1142,N_1103);
nand U1327 (N_1327,N_1048,N_1018);
nand U1328 (N_1328,N_1125,N_1110);
or U1329 (N_1329,N_1084,N_1193);
nand U1330 (N_1330,N_1070,N_1193);
nor U1331 (N_1331,N_1196,N_1159);
xor U1332 (N_1332,N_1103,N_1057);
xnor U1333 (N_1333,N_1090,N_1165);
or U1334 (N_1334,N_1062,N_1117);
and U1335 (N_1335,N_1161,N_1042);
and U1336 (N_1336,N_1121,N_1021);
or U1337 (N_1337,N_1132,N_1084);
xnor U1338 (N_1338,N_1016,N_1141);
xnor U1339 (N_1339,N_1046,N_1088);
nand U1340 (N_1340,N_1061,N_1006);
nand U1341 (N_1341,N_1069,N_1152);
nand U1342 (N_1342,N_1031,N_1002);
nor U1343 (N_1343,N_1032,N_1147);
xor U1344 (N_1344,N_1072,N_1058);
xor U1345 (N_1345,N_1125,N_1094);
or U1346 (N_1346,N_1014,N_1087);
or U1347 (N_1347,N_1120,N_1131);
and U1348 (N_1348,N_1196,N_1168);
nand U1349 (N_1349,N_1043,N_1187);
xnor U1350 (N_1350,N_1018,N_1041);
nand U1351 (N_1351,N_1094,N_1149);
xor U1352 (N_1352,N_1154,N_1102);
or U1353 (N_1353,N_1176,N_1118);
xnor U1354 (N_1354,N_1137,N_1015);
nand U1355 (N_1355,N_1190,N_1144);
nand U1356 (N_1356,N_1198,N_1136);
nand U1357 (N_1357,N_1138,N_1013);
nand U1358 (N_1358,N_1076,N_1183);
nand U1359 (N_1359,N_1115,N_1141);
and U1360 (N_1360,N_1013,N_1185);
and U1361 (N_1361,N_1040,N_1128);
or U1362 (N_1362,N_1000,N_1069);
nor U1363 (N_1363,N_1007,N_1077);
and U1364 (N_1364,N_1082,N_1061);
xnor U1365 (N_1365,N_1050,N_1022);
nand U1366 (N_1366,N_1112,N_1147);
xor U1367 (N_1367,N_1020,N_1100);
or U1368 (N_1368,N_1013,N_1104);
and U1369 (N_1369,N_1107,N_1055);
and U1370 (N_1370,N_1145,N_1069);
nand U1371 (N_1371,N_1143,N_1149);
nor U1372 (N_1372,N_1188,N_1173);
nor U1373 (N_1373,N_1194,N_1158);
and U1374 (N_1374,N_1003,N_1013);
xnor U1375 (N_1375,N_1039,N_1002);
or U1376 (N_1376,N_1039,N_1010);
xor U1377 (N_1377,N_1168,N_1099);
xor U1378 (N_1378,N_1167,N_1199);
xnor U1379 (N_1379,N_1193,N_1119);
and U1380 (N_1380,N_1014,N_1105);
xnor U1381 (N_1381,N_1162,N_1184);
nand U1382 (N_1382,N_1162,N_1101);
nand U1383 (N_1383,N_1043,N_1175);
xor U1384 (N_1384,N_1121,N_1199);
nand U1385 (N_1385,N_1193,N_1170);
nor U1386 (N_1386,N_1075,N_1084);
and U1387 (N_1387,N_1131,N_1000);
nand U1388 (N_1388,N_1193,N_1154);
nor U1389 (N_1389,N_1142,N_1061);
xnor U1390 (N_1390,N_1134,N_1000);
nor U1391 (N_1391,N_1059,N_1155);
xnor U1392 (N_1392,N_1031,N_1144);
nand U1393 (N_1393,N_1145,N_1112);
nor U1394 (N_1394,N_1133,N_1162);
nand U1395 (N_1395,N_1153,N_1004);
xnor U1396 (N_1396,N_1157,N_1048);
nand U1397 (N_1397,N_1125,N_1173);
nand U1398 (N_1398,N_1097,N_1198);
nand U1399 (N_1399,N_1092,N_1020);
and U1400 (N_1400,N_1360,N_1288);
nand U1401 (N_1401,N_1297,N_1320);
nor U1402 (N_1402,N_1394,N_1350);
or U1403 (N_1403,N_1237,N_1307);
xnor U1404 (N_1404,N_1382,N_1263);
nor U1405 (N_1405,N_1217,N_1223);
or U1406 (N_1406,N_1388,N_1353);
nand U1407 (N_1407,N_1399,N_1224);
nor U1408 (N_1408,N_1304,N_1232);
nand U1409 (N_1409,N_1257,N_1261);
nor U1410 (N_1410,N_1398,N_1367);
xnor U1411 (N_1411,N_1264,N_1219);
xor U1412 (N_1412,N_1317,N_1258);
xnor U1413 (N_1413,N_1332,N_1222);
xnor U1414 (N_1414,N_1236,N_1349);
nand U1415 (N_1415,N_1325,N_1283);
nand U1416 (N_1416,N_1213,N_1233);
nand U1417 (N_1417,N_1318,N_1313);
nor U1418 (N_1418,N_1384,N_1385);
nor U1419 (N_1419,N_1345,N_1253);
xor U1420 (N_1420,N_1206,N_1285);
or U1421 (N_1421,N_1259,N_1231);
nand U1422 (N_1422,N_1295,N_1269);
nand U1423 (N_1423,N_1234,N_1359);
xor U1424 (N_1424,N_1352,N_1267);
nor U1425 (N_1425,N_1372,N_1326);
nand U1426 (N_1426,N_1204,N_1312);
xnor U1427 (N_1427,N_1275,N_1230);
xor U1428 (N_1428,N_1272,N_1357);
xnor U1429 (N_1429,N_1362,N_1266);
xnor U1430 (N_1430,N_1247,N_1270);
and U1431 (N_1431,N_1205,N_1347);
or U1432 (N_1432,N_1211,N_1391);
xnor U1433 (N_1433,N_1355,N_1235);
or U1434 (N_1434,N_1280,N_1251);
nand U1435 (N_1435,N_1324,N_1208);
nand U1436 (N_1436,N_1358,N_1293);
nor U1437 (N_1437,N_1303,N_1308);
and U1438 (N_1438,N_1329,N_1323);
nand U1439 (N_1439,N_1338,N_1248);
nor U1440 (N_1440,N_1273,N_1225);
and U1441 (N_1441,N_1282,N_1389);
nor U1442 (N_1442,N_1207,N_1212);
and U1443 (N_1443,N_1256,N_1292);
nor U1444 (N_1444,N_1227,N_1340);
nor U1445 (N_1445,N_1226,N_1214);
xnor U1446 (N_1446,N_1315,N_1376);
nor U1447 (N_1447,N_1228,N_1316);
or U1448 (N_1448,N_1215,N_1243);
and U1449 (N_1449,N_1202,N_1311);
and U1450 (N_1450,N_1265,N_1250);
or U1451 (N_1451,N_1244,N_1374);
nor U1452 (N_1452,N_1271,N_1339);
xor U1453 (N_1453,N_1363,N_1284);
and U1454 (N_1454,N_1346,N_1242);
nand U1455 (N_1455,N_1369,N_1314);
xor U1456 (N_1456,N_1337,N_1302);
and U1457 (N_1457,N_1392,N_1305);
or U1458 (N_1458,N_1380,N_1245);
nand U1459 (N_1459,N_1368,N_1390);
xor U1460 (N_1460,N_1289,N_1383);
nand U1461 (N_1461,N_1336,N_1301);
or U1462 (N_1462,N_1278,N_1246);
nand U1463 (N_1463,N_1375,N_1218);
or U1464 (N_1464,N_1351,N_1331);
nor U1465 (N_1465,N_1354,N_1333);
and U1466 (N_1466,N_1309,N_1365);
and U1467 (N_1467,N_1238,N_1220);
nand U1468 (N_1468,N_1200,N_1387);
or U1469 (N_1469,N_1328,N_1341);
or U1470 (N_1470,N_1378,N_1310);
and U1471 (N_1471,N_1255,N_1348);
and U1472 (N_1472,N_1386,N_1286);
or U1473 (N_1473,N_1335,N_1277);
nor U1474 (N_1474,N_1299,N_1252);
or U1475 (N_1475,N_1327,N_1366);
or U1476 (N_1476,N_1322,N_1344);
and U1477 (N_1477,N_1210,N_1319);
and U1478 (N_1478,N_1396,N_1274);
nand U1479 (N_1479,N_1260,N_1300);
nand U1480 (N_1480,N_1379,N_1221);
or U1481 (N_1481,N_1241,N_1279);
nor U1482 (N_1482,N_1334,N_1262);
xnor U1483 (N_1483,N_1395,N_1281);
nor U1484 (N_1484,N_1373,N_1276);
or U1485 (N_1485,N_1249,N_1342);
or U1486 (N_1486,N_1209,N_1356);
and U1487 (N_1487,N_1296,N_1321);
xnor U1488 (N_1488,N_1294,N_1291);
and U1489 (N_1489,N_1290,N_1381);
or U1490 (N_1490,N_1239,N_1361);
and U1491 (N_1491,N_1306,N_1201);
xnor U1492 (N_1492,N_1203,N_1397);
nor U1493 (N_1493,N_1287,N_1370);
or U1494 (N_1494,N_1393,N_1343);
and U1495 (N_1495,N_1216,N_1268);
and U1496 (N_1496,N_1377,N_1330);
xnor U1497 (N_1497,N_1371,N_1298);
and U1498 (N_1498,N_1240,N_1254);
nand U1499 (N_1499,N_1229,N_1364);
xnor U1500 (N_1500,N_1254,N_1313);
nor U1501 (N_1501,N_1232,N_1202);
xor U1502 (N_1502,N_1389,N_1294);
nor U1503 (N_1503,N_1347,N_1372);
and U1504 (N_1504,N_1293,N_1207);
xor U1505 (N_1505,N_1306,N_1214);
xnor U1506 (N_1506,N_1207,N_1232);
or U1507 (N_1507,N_1334,N_1307);
and U1508 (N_1508,N_1227,N_1297);
and U1509 (N_1509,N_1382,N_1246);
xor U1510 (N_1510,N_1334,N_1212);
xnor U1511 (N_1511,N_1316,N_1330);
nor U1512 (N_1512,N_1394,N_1382);
xnor U1513 (N_1513,N_1274,N_1333);
xor U1514 (N_1514,N_1291,N_1323);
and U1515 (N_1515,N_1318,N_1208);
or U1516 (N_1516,N_1299,N_1357);
xnor U1517 (N_1517,N_1328,N_1387);
xnor U1518 (N_1518,N_1247,N_1337);
xor U1519 (N_1519,N_1312,N_1274);
or U1520 (N_1520,N_1292,N_1301);
xnor U1521 (N_1521,N_1251,N_1239);
or U1522 (N_1522,N_1225,N_1236);
nand U1523 (N_1523,N_1245,N_1241);
nand U1524 (N_1524,N_1390,N_1245);
nor U1525 (N_1525,N_1268,N_1379);
xor U1526 (N_1526,N_1226,N_1304);
xnor U1527 (N_1527,N_1300,N_1282);
and U1528 (N_1528,N_1274,N_1343);
nand U1529 (N_1529,N_1304,N_1270);
nand U1530 (N_1530,N_1318,N_1269);
nor U1531 (N_1531,N_1286,N_1377);
xnor U1532 (N_1532,N_1235,N_1350);
or U1533 (N_1533,N_1202,N_1331);
nand U1534 (N_1534,N_1223,N_1326);
and U1535 (N_1535,N_1353,N_1246);
or U1536 (N_1536,N_1346,N_1257);
and U1537 (N_1537,N_1381,N_1226);
xnor U1538 (N_1538,N_1397,N_1284);
or U1539 (N_1539,N_1207,N_1249);
xnor U1540 (N_1540,N_1263,N_1201);
xnor U1541 (N_1541,N_1361,N_1370);
or U1542 (N_1542,N_1245,N_1302);
or U1543 (N_1543,N_1307,N_1395);
or U1544 (N_1544,N_1281,N_1378);
nor U1545 (N_1545,N_1203,N_1355);
nor U1546 (N_1546,N_1376,N_1359);
nor U1547 (N_1547,N_1229,N_1251);
and U1548 (N_1548,N_1210,N_1289);
nor U1549 (N_1549,N_1396,N_1278);
or U1550 (N_1550,N_1376,N_1238);
or U1551 (N_1551,N_1249,N_1316);
or U1552 (N_1552,N_1383,N_1313);
nand U1553 (N_1553,N_1324,N_1381);
nand U1554 (N_1554,N_1285,N_1363);
and U1555 (N_1555,N_1343,N_1270);
xor U1556 (N_1556,N_1328,N_1318);
and U1557 (N_1557,N_1380,N_1355);
xnor U1558 (N_1558,N_1396,N_1389);
nor U1559 (N_1559,N_1223,N_1260);
or U1560 (N_1560,N_1326,N_1350);
xnor U1561 (N_1561,N_1258,N_1261);
and U1562 (N_1562,N_1221,N_1339);
and U1563 (N_1563,N_1290,N_1216);
or U1564 (N_1564,N_1240,N_1304);
nor U1565 (N_1565,N_1278,N_1277);
nor U1566 (N_1566,N_1222,N_1226);
nor U1567 (N_1567,N_1235,N_1289);
or U1568 (N_1568,N_1238,N_1319);
and U1569 (N_1569,N_1285,N_1346);
nor U1570 (N_1570,N_1306,N_1226);
nand U1571 (N_1571,N_1298,N_1360);
or U1572 (N_1572,N_1327,N_1256);
or U1573 (N_1573,N_1343,N_1332);
or U1574 (N_1574,N_1301,N_1282);
nand U1575 (N_1575,N_1364,N_1389);
and U1576 (N_1576,N_1236,N_1263);
nand U1577 (N_1577,N_1224,N_1391);
or U1578 (N_1578,N_1202,N_1373);
nand U1579 (N_1579,N_1343,N_1241);
nand U1580 (N_1580,N_1307,N_1390);
or U1581 (N_1581,N_1365,N_1282);
xor U1582 (N_1582,N_1340,N_1381);
xor U1583 (N_1583,N_1293,N_1333);
xnor U1584 (N_1584,N_1331,N_1312);
xnor U1585 (N_1585,N_1369,N_1206);
and U1586 (N_1586,N_1300,N_1339);
nand U1587 (N_1587,N_1287,N_1397);
nor U1588 (N_1588,N_1334,N_1345);
and U1589 (N_1589,N_1254,N_1300);
xnor U1590 (N_1590,N_1339,N_1328);
nand U1591 (N_1591,N_1334,N_1367);
nor U1592 (N_1592,N_1377,N_1291);
xnor U1593 (N_1593,N_1344,N_1281);
nand U1594 (N_1594,N_1258,N_1226);
and U1595 (N_1595,N_1243,N_1214);
and U1596 (N_1596,N_1337,N_1321);
xnor U1597 (N_1597,N_1257,N_1232);
xor U1598 (N_1598,N_1282,N_1246);
or U1599 (N_1599,N_1244,N_1306);
xor U1600 (N_1600,N_1417,N_1546);
nor U1601 (N_1601,N_1586,N_1593);
nand U1602 (N_1602,N_1486,N_1542);
and U1603 (N_1603,N_1495,N_1553);
nor U1604 (N_1604,N_1509,N_1535);
or U1605 (N_1605,N_1554,N_1468);
and U1606 (N_1606,N_1549,N_1424);
or U1607 (N_1607,N_1474,N_1513);
and U1608 (N_1608,N_1412,N_1415);
xor U1609 (N_1609,N_1505,N_1589);
nor U1610 (N_1610,N_1544,N_1472);
nand U1611 (N_1611,N_1539,N_1512);
xor U1612 (N_1612,N_1446,N_1431);
and U1613 (N_1613,N_1447,N_1471);
nand U1614 (N_1614,N_1518,N_1540);
or U1615 (N_1615,N_1462,N_1420);
or U1616 (N_1616,N_1499,N_1478);
and U1617 (N_1617,N_1436,N_1405);
xnor U1618 (N_1618,N_1489,N_1562);
or U1619 (N_1619,N_1584,N_1560);
nand U1620 (N_1620,N_1545,N_1402);
nor U1621 (N_1621,N_1506,N_1504);
xor U1622 (N_1622,N_1449,N_1527);
nor U1623 (N_1623,N_1592,N_1580);
or U1624 (N_1624,N_1414,N_1521);
nand U1625 (N_1625,N_1467,N_1524);
xnor U1626 (N_1626,N_1550,N_1531);
xnor U1627 (N_1627,N_1583,N_1522);
nor U1628 (N_1628,N_1451,N_1496);
nor U1629 (N_1629,N_1481,N_1422);
or U1630 (N_1630,N_1571,N_1557);
and U1631 (N_1631,N_1483,N_1438);
nor U1632 (N_1632,N_1595,N_1588);
xnor U1633 (N_1633,N_1514,N_1572);
xor U1634 (N_1634,N_1590,N_1458);
and U1635 (N_1635,N_1400,N_1536);
nand U1636 (N_1636,N_1575,N_1475);
nand U1637 (N_1637,N_1555,N_1587);
xor U1638 (N_1638,N_1455,N_1484);
xor U1639 (N_1639,N_1563,N_1480);
and U1640 (N_1640,N_1437,N_1517);
xnor U1641 (N_1641,N_1528,N_1461);
and U1642 (N_1642,N_1582,N_1444);
xnor U1643 (N_1643,N_1430,N_1538);
and U1644 (N_1644,N_1568,N_1429);
or U1645 (N_1645,N_1525,N_1526);
xnor U1646 (N_1646,N_1561,N_1511);
and U1647 (N_1647,N_1497,N_1532);
and U1648 (N_1648,N_1502,N_1441);
xor U1649 (N_1649,N_1594,N_1529);
xor U1650 (N_1650,N_1515,N_1564);
and U1651 (N_1651,N_1410,N_1547);
and U1652 (N_1652,N_1427,N_1534);
xnor U1653 (N_1653,N_1425,N_1465);
or U1654 (N_1654,N_1597,N_1477);
nor U1655 (N_1655,N_1408,N_1566);
nand U1656 (N_1656,N_1537,N_1579);
or U1657 (N_1657,N_1407,N_1570);
nand U1658 (N_1658,N_1473,N_1448);
nand U1659 (N_1659,N_1419,N_1490);
and U1660 (N_1660,N_1543,N_1574);
and U1661 (N_1661,N_1573,N_1432);
xnor U1662 (N_1662,N_1411,N_1533);
nand U1663 (N_1663,N_1459,N_1445);
nand U1664 (N_1664,N_1413,N_1463);
nand U1665 (N_1665,N_1498,N_1491);
or U1666 (N_1666,N_1460,N_1569);
xor U1667 (N_1667,N_1464,N_1428);
or U1668 (N_1668,N_1520,N_1403);
xor U1669 (N_1669,N_1482,N_1479);
and U1670 (N_1670,N_1501,N_1585);
xnor U1671 (N_1671,N_1510,N_1423);
or U1672 (N_1672,N_1488,N_1577);
nor U1673 (N_1673,N_1466,N_1552);
or U1674 (N_1674,N_1435,N_1406);
nor U1675 (N_1675,N_1456,N_1409);
nand U1676 (N_1676,N_1565,N_1401);
nor U1677 (N_1677,N_1433,N_1519);
nor U1678 (N_1678,N_1469,N_1452);
nand U1679 (N_1679,N_1598,N_1418);
xor U1680 (N_1680,N_1416,N_1476);
or U1681 (N_1681,N_1599,N_1440);
nand U1682 (N_1682,N_1442,N_1434);
nor U1683 (N_1683,N_1450,N_1404);
nor U1684 (N_1684,N_1487,N_1523);
nor U1685 (N_1685,N_1516,N_1508);
or U1686 (N_1686,N_1503,N_1485);
xor U1687 (N_1687,N_1530,N_1470);
and U1688 (N_1688,N_1500,N_1581);
or U1689 (N_1689,N_1457,N_1443);
or U1690 (N_1690,N_1421,N_1596);
nor U1691 (N_1691,N_1453,N_1558);
and U1692 (N_1692,N_1439,N_1576);
nor U1693 (N_1693,N_1559,N_1548);
or U1694 (N_1694,N_1567,N_1578);
or U1695 (N_1695,N_1556,N_1541);
xor U1696 (N_1696,N_1493,N_1492);
and U1697 (N_1697,N_1454,N_1494);
nor U1698 (N_1698,N_1507,N_1426);
and U1699 (N_1699,N_1591,N_1551);
or U1700 (N_1700,N_1504,N_1570);
and U1701 (N_1701,N_1421,N_1557);
and U1702 (N_1702,N_1547,N_1425);
and U1703 (N_1703,N_1537,N_1517);
nand U1704 (N_1704,N_1514,N_1559);
and U1705 (N_1705,N_1496,N_1572);
or U1706 (N_1706,N_1552,N_1531);
xor U1707 (N_1707,N_1557,N_1587);
and U1708 (N_1708,N_1402,N_1487);
nor U1709 (N_1709,N_1455,N_1501);
nand U1710 (N_1710,N_1523,N_1493);
and U1711 (N_1711,N_1431,N_1583);
nor U1712 (N_1712,N_1464,N_1415);
nand U1713 (N_1713,N_1596,N_1411);
nand U1714 (N_1714,N_1442,N_1556);
xnor U1715 (N_1715,N_1481,N_1556);
nor U1716 (N_1716,N_1540,N_1450);
nand U1717 (N_1717,N_1585,N_1535);
nor U1718 (N_1718,N_1535,N_1416);
xnor U1719 (N_1719,N_1422,N_1446);
nor U1720 (N_1720,N_1575,N_1471);
nor U1721 (N_1721,N_1424,N_1445);
xor U1722 (N_1722,N_1415,N_1501);
xnor U1723 (N_1723,N_1455,N_1497);
or U1724 (N_1724,N_1437,N_1490);
xnor U1725 (N_1725,N_1408,N_1517);
or U1726 (N_1726,N_1496,N_1524);
nor U1727 (N_1727,N_1442,N_1495);
or U1728 (N_1728,N_1401,N_1427);
nor U1729 (N_1729,N_1459,N_1537);
xor U1730 (N_1730,N_1523,N_1592);
nor U1731 (N_1731,N_1442,N_1486);
nand U1732 (N_1732,N_1536,N_1590);
or U1733 (N_1733,N_1468,N_1599);
nand U1734 (N_1734,N_1425,N_1439);
nand U1735 (N_1735,N_1535,N_1434);
nor U1736 (N_1736,N_1587,N_1556);
nor U1737 (N_1737,N_1521,N_1490);
nand U1738 (N_1738,N_1482,N_1597);
nand U1739 (N_1739,N_1461,N_1549);
nand U1740 (N_1740,N_1404,N_1521);
nand U1741 (N_1741,N_1501,N_1570);
nor U1742 (N_1742,N_1456,N_1497);
and U1743 (N_1743,N_1597,N_1476);
xnor U1744 (N_1744,N_1542,N_1511);
or U1745 (N_1745,N_1504,N_1404);
xnor U1746 (N_1746,N_1599,N_1497);
nor U1747 (N_1747,N_1501,N_1418);
nor U1748 (N_1748,N_1434,N_1532);
nor U1749 (N_1749,N_1565,N_1475);
nand U1750 (N_1750,N_1474,N_1485);
xor U1751 (N_1751,N_1572,N_1402);
xnor U1752 (N_1752,N_1404,N_1423);
nor U1753 (N_1753,N_1469,N_1556);
nand U1754 (N_1754,N_1488,N_1558);
and U1755 (N_1755,N_1550,N_1533);
and U1756 (N_1756,N_1574,N_1528);
xnor U1757 (N_1757,N_1460,N_1465);
and U1758 (N_1758,N_1586,N_1550);
xnor U1759 (N_1759,N_1424,N_1433);
and U1760 (N_1760,N_1456,N_1562);
nand U1761 (N_1761,N_1565,N_1420);
nor U1762 (N_1762,N_1524,N_1484);
nor U1763 (N_1763,N_1451,N_1596);
nand U1764 (N_1764,N_1504,N_1511);
nor U1765 (N_1765,N_1503,N_1424);
nor U1766 (N_1766,N_1592,N_1504);
or U1767 (N_1767,N_1535,N_1592);
nand U1768 (N_1768,N_1441,N_1508);
and U1769 (N_1769,N_1435,N_1482);
xnor U1770 (N_1770,N_1486,N_1437);
nor U1771 (N_1771,N_1593,N_1457);
and U1772 (N_1772,N_1577,N_1594);
nor U1773 (N_1773,N_1535,N_1574);
or U1774 (N_1774,N_1413,N_1506);
and U1775 (N_1775,N_1473,N_1414);
or U1776 (N_1776,N_1481,N_1585);
and U1777 (N_1777,N_1584,N_1410);
and U1778 (N_1778,N_1466,N_1477);
nand U1779 (N_1779,N_1560,N_1576);
or U1780 (N_1780,N_1440,N_1452);
xor U1781 (N_1781,N_1571,N_1560);
nand U1782 (N_1782,N_1578,N_1549);
xor U1783 (N_1783,N_1509,N_1456);
nor U1784 (N_1784,N_1448,N_1541);
nor U1785 (N_1785,N_1584,N_1596);
nor U1786 (N_1786,N_1485,N_1464);
nor U1787 (N_1787,N_1469,N_1533);
and U1788 (N_1788,N_1593,N_1501);
and U1789 (N_1789,N_1423,N_1528);
nand U1790 (N_1790,N_1437,N_1584);
and U1791 (N_1791,N_1468,N_1418);
or U1792 (N_1792,N_1447,N_1514);
or U1793 (N_1793,N_1552,N_1561);
or U1794 (N_1794,N_1526,N_1415);
nor U1795 (N_1795,N_1536,N_1526);
nand U1796 (N_1796,N_1446,N_1517);
or U1797 (N_1797,N_1558,N_1548);
nor U1798 (N_1798,N_1573,N_1542);
xnor U1799 (N_1799,N_1432,N_1479);
or U1800 (N_1800,N_1648,N_1661);
nand U1801 (N_1801,N_1692,N_1671);
and U1802 (N_1802,N_1741,N_1782);
or U1803 (N_1803,N_1652,N_1797);
nor U1804 (N_1804,N_1680,N_1754);
nor U1805 (N_1805,N_1767,N_1675);
xor U1806 (N_1806,N_1690,N_1721);
xnor U1807 (N_1807,N_1669,N_1704);
nand U1808 (N_1808,N_1683,N_1771);
or U1809 (N_1809,N_1733,N_1760);
or U1810 (N_1810,N_1738,N_1644);
and U1811 (N_1811,N_1616,N_1757);
nand U1812 (N_1812,N_1629,N_1613);
or U1813 (N_1813,N_1667,N_1612);
nand U1814 (N_1814,N_1676,N_1649);
or U1815 (N_1815,N_1748,N_1707);
and U1816 (N_1816,N_1663,N_1632);
nand U1817 (N_1817,N_1688,N_1702);
nand U1818 (N_1818,N_1665,N_1609);
nor U1819 (N_1819,N_1641,N_1745);
xor U1820 (N_1820,N_1716,N_1742);
or U1821 (N_1821,N_1780,N_1747);
nand U1822 (N_1822,N_1758,N_1701);
nand U1823 (N_1823,N_1793,N_1726);
and U1824 (N_1824,N_1600,N_1615);
xor U1825 (N_1825,N_1635,N_1769);
nand U1826 (N_1826,N_1603,N_1705);
nand U1827 (N_1827,N_1775,N_1684);
nand U1828 (N_1828,N_1651,N_1647);
and U1829 (N_1829,N_1777,N_1729);
xnor U1830 (N_1830,N_1677,N_1772);
xor U1831 (N_1831,N_1611,N_1620);
and U1832 (N_1832,N_1720,N_1781);
nor U1833 (N_1833,N_1714,N_1679);
and U1834 (N_1834,N_1696,N_1630);
nand U1835 (N_1835,N_1637,N_1786);
xnor U1836 (N_1836,N_1626,N_1792);
and U1837 (N_1837,N_1659,N_1619);
nor U1838 (N_1838,N_1674,N_1645);
xnor U1839 (N_1839,N_1617,N_1776);
xnor U1840 (N_1840,N_1666,N_1689);
and U1841 (N_1841,N_1799,N_1695);
nand U1842 (N_1842,N_1653,N_1761);
nand U1843 (N_1843,N_1606,N_1697);
and U1844 (N_1844,N_1788,N_1654);
nand U1845 (N_1845,N_1631,N_1766);
nor U1846 (N_1846,N_1715,N_1734);
xnor U1847 (N_1847,N_1610,N_1763);
nor U1848 (N_1848,N_1770,N_1795);
xnor U1849 (N_1849,N_1727,N_1672);
nor U1850 (N_1850,N_1650,N_1798);
and U1851 (N_1851,N_1700,N_1685);
and U1852 (N_1852,N_1622,N_1732);
or U1853 (N_1853,N_1655,N_1664);
nor U1854 (N_1854,N_1710,N_1794);
xnor U1855 (N_1855,N_1787,N_1625);
and U1856 (N_1856,N_1724,N_1633);
nor U1857 (N_1857,N_1642,N_1601);
xor U1858 (N_1858,N_1604,N_1627);
nand U1859 (N_1859,N_1686,N_1670);
nor U1860 (N_1860,N_1691,N_1737);
nor U1861 (N_1861,N_1711,N_1713);
xnor U1862 (N_1862,N_1759,N_1706);
nor U1863 (N_1863,N_1790,N_1608);
nand U1864 (N_1864,N_1657,N_1773);
nand U1865 (N_1865,N_1698,N_1719);
and U1866 (N_1866,N_1784,N_1658);
and U1867 (N_1867,N_1756,N_1739);
nand U1868 (N_1868,N_1694,N_1628);
xnor U1869 (N_1869,N_1646,N_1740);
or U1870 (N_1870,N_1774,N_1602);
nand U1871 (N_1871,N_1723,N_1725);
and U1872 (N_1872,N_1699,N_1750);
nor U1873 (N_1873,N_1722,N_1639);
nand U1874 (N_1874,N_1709,N_1623);
nand U1875 (N_1875,N_1668,N_1785);
xor U1876 (N_1876,N_1638,N_1783);
or U1877 (N_1877,N_1779,N_1681);
or U1878 (N_1878,N_1743,N_1703);
and U1879 (N_1879,N_1618,N_1662);
nand U1880 (N_1880,N_1728,N_1755);
nand U1881 (N_1881,N_1621,N_1765);
or U1882 (N_1882,N_1735,N_1643);
nor U1883 (N_1883,N_1640,N_1791);
nor U1884 (N_1884,N_1796,N_1789);
nor U1885 (N_1885,N_1634,N_1712);
nand U1886 (N_1886,N_1752,N_1607);
xnor U1887 (N_1887,N_1656,N_1693);
nor U1888 (N_1888,N_1731,N_1744);
nand U1889 (N_1889,N_1730,N_1768);
or U1890 (N_1890,N_1753,N_1736);
nand U1891 (N_1891,N_1678,N_1778);
xnor U1892 (N_1892,N_1614,N_1624);
nand U1893 (N_1893,N_1718,N_1749);
and U1894 (N_1894,N_1673,N_1636);
or U1895 (N_1895,N_1764,N_1746);
nand U1896 (N_1896,N_1708,N_1762);
xnor U1897 (N_1897,N_1682,N_1687);
or U1898 (N_1898,N_1717,N_1751);
xor U1899 (N_1899,N_1660,N_1605);
xor U1900 (N_1900,N_1644,N_1739);
or U1901 (N_1901,N_1717,N_1635);
nor U1902 (N_1902,N_1747,N_1621);
or U1903 (N_1903,N_1619,N_1636);
nor U1904 (N_1904,N_1723,N_1733);
or U1905 (N_1905,N_1766,N_1773);
nand U1906 (N_1906,N_1605,N_1699);
xor U1907 (N_1907,N_1662,N_1782);
or U1908 (N_1908,N_1768,N_1728);
or U1909 (N_1909,N_1779,N_1777);
nor U1910 (N_1910,N_1646,N_1705);
nand U1911 (N_1911,N_1710,N_1642);
or U1912 (N_1912,N_1693,N_1772);
nor U1913 (N_1913,N_1683,N_1689);
or U1914 (N_1914,N_1624,N_1660);
or U1915 (N_1915,N_1635,N_1797);
nor U1916 (N_1916,N_1623,N_1618);
or U1917 (N_1917,N_1756,N_1715);
and U1918 (N_1918,N_1666,N_1715);
nand U1919 (N_1919,N_1619,N_1692);
nand U1920 (N_1920,N_1669,N_1655);
or U1921 (N_1921,N_1749,N_1782);
nand U1922 (N_1922,N_1799,N_1640);
xnor U1923 (N_1923,N_1794,N_1670);
nand U1924 (N_1924,N_1774,N_1670);
and U1925 (N_1925,N_1778,N_1696);
and U1926 (N_1926,N_1678,N_1682);
or U1927 (N_1927,N_1609,N_1759);
nor U1928 (N_1928,N_1640,N_1645);
or U1929 (N_1929,N_1700,N_1733);
and U1930 (N_1930,N_1616,N_1738);
or U1931 (N_1931,N_1730,N_1799);
or U1932 (N_1932,N_1635,N_1727);
xor U1933 (N_1933,N_1684,N_1722);
nand U1934 (N_1934,N_1700,N_1669);
nor U1935 (N_1935,N_1703,N_1758);
nor U1936 (N_1936,N_1790,N_1769);
and U1937 (N_1937,N_1701,N_1714);
nor U1938 (N_1938,N_1719,N_1707);
or U1939 (N_1939,N_1654,N_1732);
xor U1940 (N_1940,N_1698,N_1679);
nor U1941 (N_1941,N_1691,N_1701);
and U1942 (N_1942,N_1758,N_1720);
nor U1943 (N_1943,N_1790,N_1742);
xnor U1944 (N_1944,N_1663,N_1638);
or U1945 (N_1945,N_1734,N_1602);
xor U1946 (N_1946,N_1776,N_1650);
or U1947 (N_1947,N_1734,N_1695);
or U1948 (N_1948,N_1667,N_1770);
xor U1949 (N_1949,N_1753,N_1796);
and U1950 (N_1950,N_1737,N_1649);
xor U1951 (N_1951,N_1679,N_1613);
and U1952 (N_1952,N_1706,N_1643);
and U1953 (N_1953,N_1626,N_1779);
xnor U1954 (N_1954,N_1674,N_1699);
nand U1955 (N_1955,N_1769,N_1632);
nand U1956 (N_1956,N_1792,N_1663);
or U1957 (N_1957,N_1656,N_1648);
and U1958 (N_1958,N_1621,N_1647);
nor U1959 (N_1959,N_1664,N_1707);
nor U1960 (N_1960,N_1728,N_1705);
nand U1961 (N_1961,N_1737,N_1741);
xnor U1962 (N_1962,N_1752,N_1750);
nor U1963 (N_1963,N_1681,N_1735);
xnor U1964 (N_1964,N_1766,N_1779);
xnor U1965 (N_1965,N_1635,N_1763);
xnor U1966 (N_1966,N_1777,N_1788);
nor U1967 (N_1967,N_1682,N_1775);
nor U1968 (N_1968,N_1640,N_1704);
and U1969 (N_1969,N_1618,N_1768);
xor U1970 (N_1970,N_1775,N_1608);
and U1971 (N_1971,N_1602,N_1725);
xnor U1972 (N_1972,N_1764,N_1771);
and U1973 (N_1973,N_1723,N_1668);
xnor U1974 (N_1974,N_1670,N_1691);
nand U1975 (N_1975,N_1648,N_1629);
or U1976 (N_1976,N_1646,N_1649);
and U1977 (N_1977,N_1669,N_1749);
and U1978 (N_1978,N_1604,N_1632);
nand U1979 (N_1979,N_1636,N_1755);
nand U1980 (N_1980,N_1788,N_1642);
nor U1981 (N_1981,N_1725,N_1662);
nand U1982 (N_1982,N_1615,N_1783);
or U1983 (N_1983,N_1796,N_1763);
or U1984 (N_1984,N_1736,N_1798);
nor U1985 (N_1985,N_1652,N_1669);
nand U1986 (N_1986,N_1686,N_1758);
xnor U1987 (N_1987,N_1629,N_1763);
and U1988 (N_1988,N_1695,N_1786);
and U1989 (N_1989,N_1772,N_1672);
or U1990 (N_1990,N_1675,N_1672);
and U1991 (N_1991,N_1774,N_1753);
or U1992 (N_1992,N_1797,N_1665);
and U1993 (N_1993,N_1631,N_1703);
xor U1994 (N_1994,N_1628,N_1639);
xnor U1995 (N_1995,N_1696,N_1644);
or U1996 (N_1996,N_1777,N_1750);
and U1997 (N_1997,N_1629,N_1636);
and U1998 (N_1998,N_1772,N_1644);
and U1999 (N_1999,N_1653,N_1697);
and U2000 (N_2000,N_1939,N_1845);
nand U2001 (N_2001,N_1811,N_1827);
or U2002 (N_2002,N_1975,N_1821);
or U2003 (N_2003,N_1829,N_1808);
and U2004 (N_2004,N_1819,N_1922);
or U2005 (N_2005,N_1871,N_1978);
xor U2006 (N_2006,N_1935,N_1900);
and U2007 (N_2007,N_1942,N_1914);
nand U2008 (N_2008,N_1875,N_1846);
nand U2009 (N_2009,N_1886,N_1999);
and U2010 (N_2010,N_1849,N_1833);
or U2011 (N_2011,N_1817,N_1854);
nand U2012 (N_2012,N_1948,N_1988);
and U2013 (N_2013,N_1934,N_1953);
xor U2014 (N_2014,N_1822,N_1993);
nand U2015 (N_2015,N_1860,N_1866);
or U2016 (N_2016,N_1800,N_1840);
or U2017 (N_2017,N_1940,N_1887);
nor U2018 (N_2018,N_1925,N_1931);
nor U2019 (N_2019,N_1927,N_1893);
or U2020 (N_2020,N_1895,N_1873);
nor U2021 (N_2021,N_1965,N_1937);
nand U2022 (N_2022,N_1888,N_1992);
xor U2023 (N_2023,N_1933,N_1859);
xor U2024 (N_2024,N_1944,N_1844);
or U2025 (N_2025,N_1928,N_1809);
and U2026 (N_2026,N_1987,N_1929);
xnor U2027 (N_2027,N_1810,N_1986);
xor U2028 (N_2028,N_1878,N_1853);
or U2029 (N_2029,N_1801,N_1973);
nand U2030 (N_2030,N_1976,N_1982);
or U2031 (N_2031,N_1995,N_1924);
or U2032 (N_2032,N_1950,N_1818);
nand U2033 (N_2033,N_1949,N_1857);
and U2034 (N_2034,N_1936,N_1960);
nand U2035 (N_2035,N_1861,N_1864);
nor U2036 (N_2036,N_1852,N_1957);
or U2037 (N_2037,N_1983,N_1923);
or U2038 (N_2038,N_1867,N_1991);
and U2039 (N_2039,N_1904,N_1890);
xnor U2040 (N_2040,N_1843,N_1915);
nor U2041 (N_2041,N_1903,N_1917);
or U2042 (N_2042,N_1894,N_1825);
and U2043 (N_2043,N_1896,N_1932);
or U2044 (N_2044,N_1838,N_1902);
and U2045 (N_2045,N_1961,N_1828);
nand U2046 (N_2046,N_1850,N_1981);
xor U2047 (N_2047,N_1984,N_1967);
and U2048 (N_2048,N_1803,N_1964);
or U2049 (N_2049,N_1834,N_1898);
or U2050 (N_2050,N_1974,N_1905);
and U2051 (N_2051,N_1835,N_1969);
xnor U2052 (N_2052,N_1814,N_1979);
xor U2053 (N_2053,N_1812,N_1862);
nand U2054 (N_2054,N_1881,N_1804);
nand U2055 (N_2055,N_1816,N_1868);
nor U2056 (N_2056,N_1882,N_1968);
or U2057 (N_2057,N_1963,N_1997);
nand U2058 (N_2058,N_1947,N_1863);
nand U2059 (N_2059,N_1971,N_1912);
and U2060 (N_2060,N_1842,N_1848);
or U2061 (N_2061,N_1989,N_1901);
xor U2062 (N_2062,N_1869,N_1891);
and U2063 (N_2063,N_1907,N_1972);
xor U2064 (N_2064,N_1906,N_1830);
or U2065 (N_2065,N_1856,N_1880);
or U2066 (N_2066,N_1956,N_1938);
or U2067 (N_2067,N_1883,N_1836);
or U2068 (N_2068,N_1897,N_1892);
or U2069 (N_2069,N_1865,N_1823);
xor U2070 (N_2070,N_1824,N_1977);
nand U2071 (N_2071,N_1955,N_1885);
and U2072 (N_2072,N_1998,N_1980);
nor U2073 (N_2073,N_1879,N_1826);
nor U2074 (N_2074,N_1806,N_1921);
nor U2075 (N_2075,N_1908,N_1877);
nor U2076 (N_2076,N_1899,N_1832);
nand U2077 (N_2077,N_1910,N_1911);
and U2078 (N_2078,N_1994,N_1954);
nand U2079 (N_2079,N_1966,N_1847);
nand U2080 (N_2080,N_1920,N_1841);
and U2081 (N_2081,N_1951,N_1874);
nor U2082 (N_2082,N_1959,N_1805);
nor U2083 (N_2083,N_1962,N_1985);
and U2084 (N_2084,N_1970,N_1839);
and U2085 (N_2085,N_1884,N_1941);
or U2086 (N_2086,N_1946,N_1952);
nor U2087 (N_2087,N_1807,N_1870);
or U2088 (N_2088,N_1918,N_1837);
and U2089 (N_2089,N_1919,N_1916);
nand U2090 (N_2090,N_1820,N_1876);
xor U2091 (N_2091,N_1872,N_1990);
xnor U2092 (N_2092,N_1930,N_1831);
and U2093 (N_2093,N_1855,N_1926);
and U2094 (N_2094,N_1958,N_1815);
or U2095 (N_2095,N_1858,N_1945);
and U2096 (N_2096,N_1913,N_1813);
xor U2097 (N_2097,N_1889,N_1909);
xor U2098 (N_2098,N_1802,N_1851);
nor U2099 (N_2099,N_1943,N_1996);
nor U2100 (N_2100,N_1871,N_1903);
nor U2101 (N_2101,N_1888,N_1959);
or U2102 (N_2102,N_1816,N_1801);
xnor U2103 (N_2103,N_1839,N_1991);
and U2104 (N_2104,N_1828,N_1974);
and U2105 (N_2105,N_1958,N_1828);
and U2106 (N_2106,N_1805,N_1860);
nand U2107 (N_2107,N_1841,N_1822);
nor U2108 (N_2108,N_1929,N_1923);
or U2109 (N_2109,N_1824,N_1860);
xor U2110 (N_2110,N_1937,N_1946);
and U2111 (N_2111,N_1944,N_1975);
and U2112 (N_2112,N_1905,N_1978);
nor U2113 (N_2113,N_1996,N_1892);
nand U2114 (N_2114,N_1956,N_1918);
xor U2115 (N_2115,N_1905,N_1909);
and U2116 (N_2116,N_1897,N_1948);
nand U2117 (N_2117,N_1923,N_1955);
nor U2118 (N_2118,N_1986,N_1980);
or U2119 (N_2119,N_1868,N_1971);
and U2120 (N_2120,N_1980,N_1999);
and U2121 (N_2121,N_1912,N_1934);
nor U2122 (N_2122,N_1993,N_1980);
or U2123 (N_2123,N_1993,N_1850);
or U2124 (N_2124,N_1803,N_1817);
and U2125 (N_2125,N_1952,N_1971);
or U2126 (N_2126,N_1900,N_1875);
or U2127 (N_2127,N_1995,N_1986);
and U2128 (N_2128,N_1984,N_1953);
or U2129 (N_2129,N_1883,N_1908);
nand U2130 (N_2130,N_1902,N_1952);
or U2131 (N_2131,N_1941,N_1870);
nor U2132 (N_2132,N_1863,N_1927);
or U2133 (N_2133,N_1839,N_1978);
or U2134 (N_2134,N_1880,N_1903);
xor U2135 (N_2135,N_1856,N_1818);
nor U2136 (N_2136,N_1846,N_1809);
nand U2137 (N_2137,N_1858,N_1833);
nand U2138 (N_2138,N_1937,N_1927);
or U2139 (N_2139,N_1867,N_1843);
or U2140 (N_2140,N_1953,N_1857);
or U2141 (N_2141,N_1981,N_1886);
xor U2142 (N_2142,N_1894,N_1823);
nor U2143 (N_2143,N_1805,N_1957);
xor U2144 (N_2144,N_1819,N_1889);
nand U2145 (N_2145,N_1893,N_1915);
xor U2146 (N_2146,N_1995,N_1835);
or U2147 (N_2147,N_1877,N_1915);
xor U2148 (N_2148,N_1861,N_1893);
nand U2149 (N_2149,N_1968,N_1811);
nor U2150 (N_2150,N_1881,N_1956);
xnor U2151 (N_2151,N_1921,N_1960);
nand U2152 (N_2152,N_1852,N_1960);
and U2153 (N_2153,N_1942,N_1911);
xor U2154 (N_2154,N_1957,N_1815);
or U2155 (N_2155,N_1988,N_1890);
nand U2156 (N_2156,N_1958,N_1812);
and U2157 (N_2157,N_1914,N_1904);
xor U2158 (N_2158,N_1859,N_1912);
and U2159 (N_2159,N_1845,N_1811);
or U2160 (N_2160,N_1882,N_1916);
nor U2161 (N_2161,N_1821,N_1980);
nand U2162 (N_2162,N_1834,N_1942);
nand U2163 (N_2163,N_1976,N_1996);
nor U2164 (N_2164,N_1865,N_1852);
and U2165 (N_2165,N_1850,N_1866);
nand U2166 (N_2166,N_1840,N_1848);
nand U2167 (N_2167,N_1876,N_1951);
nand U2168 (N_2168,N_1926,N_1986);
nand U2169 (N_2169,N_1971,N_1833);
or U2170 (N_2170,N_1836,N_1991);
or U2171 (N_2171,N_1922,N_1970);
xnor U2172 (N_2172,N_1876,N_1865);
xnor U2173 (N_2173,N_1959,N_1950);
or U2174 (N_2174,N_1820,N_1814);
xnor U2175 (N_2175,N_1860,N_1914);
or U2176 (N_2176,N_1827,N_1913);
nor U2177 (N_2177,N_1915,N_1818);
nand U2178 (N_2178,N_1908,N_1962);
xor U2179 (N_2179,N_1931,N_1836);
xnor U2180 (N_2180,N_1815,N_1821);
nor U2181 (N_2181,N_1912,N_1901);
nand U2182 (N_2182,N_1803,N_1845);
xor U2183 (N_2183,N_1866,N_1984);
or U2184 (N_2184,N_1929,N_1934);
or U2185 (N_2185,N_1892,N_1841);
nor U2186 (N_2186,N_1804,N_1832);
nor U2187 (N_2187,N_1961,N_1951);
nand U2188 (N_2188,N_1822,N_1942);
xnor U2189 (N_2189,N_1816,N_1866);
nand U2190 (N_2190,N_1847,N_1954);
nand U2191 (N_2191,N_1889,N_1836);
xor U2192 (N_2192,N_1841,N_1838);
nor U2193 (N_2193,N_1892,N_1914);
and U2194 (N_2194,N_1874,N_1857);
nor U2195 (N_2195,N_1996,N_1932);
xnor U2196 (N_2196,N_1853,N_1973);
xor U2197 (N_2197,N_1935,N_1819);
or U2198 (N_2198,N_1964,N_1990);
nor U2199 (N_2199,N_1874,N_1903);
or U2200 (N_2200,N_2124,N_2047);
or U2201 (N_2201,N_2165,N_2161);
xor U2202 (N_2202,N_2160,N_2090);
xor U2203 (N_2203,N_2108,N_2075);
or U2204 (N_2204,N_2032,N_2175);
nand U2205 (N_2205,N_2120,N_2051);
xor U2206 (N_2206,N_2187,N_2083);
nor U2207 (N_2207,N_2025,N_2041);
nand U2208 (N_2208,N_2196,N_2049);
nor U2209 (N_2209,N_2168,N_2106);
nand U2210 (N_2210,N_2194,N_2154);
nor U2211 (N_2211,N_2156,N_2101);
xor U2212 (N_2212,N_2105,N_2012);
or U2213 (N_2213,N_2043,N_2074);
or U2214 (N_2214,N_2065,N_2005);
nor U2215 (N_2215,N_2006,N_2086);
nand U2216 (N_2216,N_2099,N_2092);
and U2217 (N_2217,N_2126,N_2023);
nand U2218 (N_2218,N_2185,N_2153);
nor U2219 (N_2219,N_2027,N_2002);
nand U2220 (N_2220,N_2113,N_2037);
nor U2221 (N_2221,N_2088,N_2157);
or U2222 (N_2222,N_2193,N_2102);
xor U2223 (N_2223,N_2089,N_2095);
or U2224 (N_2224,N_2014,N_2176);
nand U2225 (N_2225,N_2056,N_2174);
or U2226 (N_2226,N_2036,N_2140);
or U2227 (N_2227,N_2183,N_2149);
nor U2228 (N_2228,N_2058,N_2097);
nor U2229 (N_2229,N_2003,N_2136);
or U2230 (N_2230,N_2080,N_2163);
and U2231 (N_2231,N_2019,N_2135);
and U2232 (N_2232,N_2181,N_2122);
xor U2233 (N_2233,N_2143,N_2031);
nor U2234 (N_2234,N_2068,N_2020);
nor U2235 (N_2235,N_2029,N_2033);
nand U2236 (N_2236,N_2178,N_2133);
nor U2237 (N_2237,N_2064,N_2171);
and U2238 (N_2238,N_2050,N_2035);
nor U2239 (N_2239,N_2008,N_2100);
nand U2240 (N_2240,N_2017,N_2131);
nand U2241 (N_2241,N_2054,N_2169);
or U2242 (N_2242,N_2162,N_2167);
and U2243 (N_2243,N_2158,N_2070);
or U2244 (N_2244,N_2172,N_2018);
nand U2245 (N_2245,N_2159,N_2059);
and U2246 (N_2246,N_2192,N_2057);
xnor U2247 (N_2247,N_2094,N_2053);
nor U2248 (N_2248,N_2128,N_2186);
xnor U2249 (N_2249,N_2114,N_2016);
or U2250 (N_2250,N_2085,N_2145);
nand U2251 (N_2251,N_2132,N_2039);
nand U2252 (N_2252,N_2180,N_2141);
nand U2253 (N_2253,N_2111,N_2123);
xnor U2254 (N_2254,N_2028,N_2125);
and U2255 (N_2255,N_2142,N_2103);
or U2256 (N_2256,N_2166,N_2188);
and U2257 (N_2257,N_2021,N_2079);
or U2258 (N_2258,N_2138,N_2081);
nand U2259 (N_2259,N_2015,N_2170);
or U2260 (N_2260,N_2030,N_2129);
nor U2261 (N_2261,N_2066,N_2110);
nand U2262 (N_2262,N_2010,N_2067);
xnor U2263 (N_2263,N_2034,N_2026);
nand U2264 (N_2264,N_2115,N_2062);
xnor U2265 (N_2265,N_2073,N_2177);
and U2266 (N_2266,N_2118,N_2011);
nand U2267 (N_2267,N_2179,N_2184);
or U2268 (N_2268,N_2093,N_2084);
nor U2269 (N_2269,N_2147,N_2013);
and U2270 (N_2270,N_2148,N_2121);
nor U2271 (N_2271,N_2063,N_2048);
or U2272 (N_2272,N_2190,N_2040);
and U2273 (N_2273,N_2001,N_2127);
or U2274 (N_2274,N_2134,N_2137);
or U2275 (N_2275,N_2055,N_2022);
nand U2276 (N_2276,N_2197,N_2139);
or U2277 (N_2277,N_2038,N_2109);
xor U2278 (N_2278,N_2116,N_2046);
xor U2279 (N_2279,N_2069,N_2182);
xnor U2280 (N_2280,N_2007,N_2042);
xor U2281 (N_2281,N_2198,N_2146);
and U2282 (N_2282,N_2045,N_2199);
nor U2283 (N_2283,N_2060,N_2000);
and U2284 (N_2284,N_2117,N_2155);
and U2285 (N_2285,N_2152,N_2151);
nor U2286 (N_2286,N_2173,N_2130);
nor U2287 (N_2287,N_2091,N_2189);
xnor U2288 (N_2288,N_2061,N_2024);
and U2289 (N_2289,N_2071,N_2112);
and U2290 (N_2290,N_2104,N_2004);
nand U2291 (N_2291,N_2119,N_2195);
xor U2292 (N_2292,N_2107,N_2164);
xor U2293 (N_2293,N_2144,N_2096);
nand U2294 (N_2294,N_2044,N_2087);
xnor U2295 (N_2295,N_2098,N_2078);
xor U2296 (N_2296,N_2191,N_2009);
and U2297 (N_2297,N_2077,N_2082);
nand U2298 (N_2298,N_2076,N_2150);
nand U2299 (N_2299,N_2072,N_2052);
and U2300 (N_2300,N_2047,N_2084);
and U2301 (N_2301,N_2102,N_2106);
or U2302 (N_2302,N_2170,N_2177);
and U2303 (N_2303,N_2054,N_2047);
xor U2304 (N_2304,N_2189,N_2021);
nor U2305 (N_2305,N_2107,N_2034);
or U2306 (N_2306,N_2007,N_2043);
nor U2307 (N_2307,N_2180,N_2121);
nor U2308 (N_2308,N_2052,N_2117);
or U2309 (N_2309,N_2162,N_2065);
nor U2310 (N_2310,N_2164,N_2004);
nor U2311 (N_2311,N_2089,N_2139);
nor U2312 (N_2312,N_2057,N_2020);
and U2313 (N_2313,N_2183,N_2057);
nand U2314 (N_2314,N_2034,N_2041);
or U2315 (N_2315,N_2174,N_2039);
or U2316 (N_2316,N_2111,N_2197);
nor U2317 (N_2317,N_2146,N_2180);
xor U2318 (N_2318,N_2079,N_2108);
nor U2319 (N_2319,N_2169,N_2093);
nor U2320 (N_2320,N_2035,N_2051);
or U2321 (N_2321,N_2058,N_2099);
nand U2322 (N_2322,N_2016,N_2040);
nand U2323 (N_2323,N_2042,N_2097);
nor U2324 (N_2324,N_2091,N_2151);
or U2325 (N_2325,N_2060,N_2039);
or U2326 (N_2326,N_2075,N_2092);
nand U2327 (N_2327,N_2073,N_2175);
and U2328 (N_2328,N_2183,N_2100);
nand U2329 (N_2329,N_2158,N_2100);
or U2330 (N_2330,N_2038,N_2120);
nor U2331 (N_2331,N_2146,N_2097);
or U2332 (N_2332,N_2017,N_2049);
nor U2333 (N_2333,N_2027,N_2070);
xnor U2334 (N_2334,N_2038,N_2158);
nor U2335 (N_2335,N_2185,N_2027);
nor U2336 (N_2336,N_2118,N_2002);
and U2337 (N_2337,N_2150,N_2159);
and U2338 (N_2338,N_2050,N_2013);
nand U2339 (N_2339,N_2092,N_2195);
xor U2340 (N_2340,N_2076,N_2191);
and U2341 (N_2341,N_2164,N_2003);
nand U2342 (N_2342,N_2159,N_2011);
and U2343 (N_2343,N_2015,N_2038);
and U2344 (N_2344,N_2139,N_2081);
and U2345 (N_2345,N_2008,N_2120);
and U2346 (N_2346,N_2115,N_2015);
nand U2347 (N_2347,N_2078,N_2122);
nand U2348 (N_2348,N_2130,N_2155);
nand U2349 (N_2349,N_2000,N_2196);
and U2350 (N_2350,N_2018,N_2198);
xnor U2351 (N_2351,N_2140,N_2064);
and U2352 (N_2352,N_2018,N_2054);
nor U2353 (N_2353,N_2085,N_2164);
and U2354 (N_2354,N_2194,N_2089);
or U2355 (N_2355,N_2166,N_2184);
or U2356 (N_2356,N_2023,N_2174);
and U2357 (N_2357,N_2160,N_2072);
nor U2358 (N_2358,N_2077,N_2098);
xnor U2359 (N_2359,N_2106,N_2050);
nor U2360 (N_2360,N_2001,N_2046);
xor U2361 (N_2361,N_2016,N_2127);
and U2362 (N_2362,N_2099,N_2065);
nand U2363 (N_2363,N_2129,N_2118);
or U2364 (N_2364,N_2070,N_2084);
nor U2365 (N_2365,N_2065,N_2166);
or U2366 (N_2366,N_2148,N_2056);
nand U2367 (N_2367,N_2033,N_2114);
nor U2368 (N_2368,N_2082,N_2182);
xor U2369 (N_2369,N_2047,N_2153);
nor U2370 (N_2370,N_2071,N_2188);
nand U2371 (N_2371,N_2110,N_2093);
xnor U2372 (N_2372,N_2071,N_2168);
nor U2373 (N_2373,N_2018,N_2100);
nor U2374 (N_2374,N_2030,N_2184);
or U2375 (N_2375,N_2100,N_2122);
and U2376 (N_2376,N_2091,N_2161);
nor U2377 (N_2377,N_2005,N_2034);
nand U2378 (N_2378,N_2190,N_2025);
xnor U2379 (N_2379,N_2033,N_2086);
nor U2380 (N_2380,N_2199,N_2114);
and U2381 (N_2381,N_2181,N_2090);
nor U2382 (N_2382,N_2066,N_2008);
xor U2383 (N_2383,N_2029,N_2146);
nor U2384 (N_2384,N_2195,N_2124);
xor U2385 (N_2385,N_2150,N_2132);
and U2386 (N_2386,N_2022,N_2160);
nor U2387 (N_2387,N_2068,N_2186);
nor U2388 (N_2388,N_2024,N_2145);
nand U2389 (N_2389,N_2158,N_2036);
nand U2390 (N_2390,N_2146,N_2091);
nand U2391 (N_2391,N_2138,N_2096);
or U2392 (N_2392,N_2076,N_2138);
nor U2393 (N_2393,N_2091,N_2028);
nand U2394 (N_2394,N_2034,N_2066);
and U2395 (N_2395,N_2049,N_2047);
and U2396 (N_2396,N_2081,N_2141);
or U2397 (N_2397,N_2003,N_2085);
nand U2398 (N_2398,N_2182,N_2060);
or U2399 (N_2399,N_2093,N_2182);
nor U2400 (N_2400,N_2348,N_2259);
nand U2401 (N_2401,N_2264,N_2272);
nand U2402 (N_2402,N_2286,N_2334);
nor U2403 (N_2403,N_2281,N_2352);
nand U2404 (N_2404,N_2224,N_2282);
xnor U2405 (N_2405,N_2253,N_2318);
nor U2406 (N_2406,N_2205,N_2262);
nand U2407 (N_2407,N_2364,N_2233);
nor U2408 (N_2408,N_2368,N_2301);
xor U2409 (N_2409,N_2375,N_2290);
or U2410 (N_2410,N_2372,N_2227);
nand U2411 (N_2411,N_2351,N_2344);
xor U2412 (N_2412,N_2346,N_2267);
or U2413 (N_2413,N_2353,N_2223);
and U2414 (N_2414,N_2232,N_2280);
xor U2415 (N_2415,N_2278,N_2356);
or U2416 (N_2416,N_2250,N_2381);
nor U2417 (N_2417,N_2366,N_2332);
or U2418 (N_2418,N_2222,N_2207);
nor U2419 (N_2419,N_2247,N_2221);
nor U2420 (N_2420,N_2374,N_2265);
or U2421 (N_2421,N_2220,N_2339);
or U2422 (N_2422,N_2300,N_2395);
nand U2423 (N_2423,N_2306,N_2303);
and U2424 (N_2424,N_2333,N_2311);
or U2425 (N_2425,N_2392,N_2327);
and U2426 (N_2426,N_2313,N_2373);
xnor U2427 (N_2427,N_2336,N_2218);
xor U2428 (N_2428,N_2248,N_2217);
nor U2429 (N_2429,N_2277,N_2316);
or U2430 (N_2430,N_2341,N_2256);
or U2431 (N_2431,N_2230,N_2245);
nand U2432 (N_2432,N_2254,N_2208);
or U2433 (N_2433,N_2321,N_2200);
or U2434 (N_2434,N_2291,N_2236);
and U2435 (N_2435,N_2314,N_2297);
or U2436 (N_2436,N_2292,N_2362);
or U2437 (N_2437,N_2210,N_2289);
nand U2438 (N_2438,N_2389,N_2363);
and U2439 (N_2439,N_2355,N_2325);
and U2440 (N_2440,N_2243,N_2257);
or U2441 (N_2441,N_2237,N_2231);
and U2442 (N_2442,N_2386,N_2331);
xor U2443 (N_2443,N_2305,N_2310);
and U2444 (N_2444,N_2229,N_2338);
xnor U2445 (N_2445,N_2328,N_2273);
or U2446 (N_2446,N_2387,N_2228);
nor U2447 (N_2447,N_2226,N_2371);
nand U2448 (N_2448,N_2343,N_2238);
and U2449 (N_2449,N_2370,N_2379);
or U2450 (N_2450,N_2399,N_2326);
xor U2451 (N_2451,N_2234,N_2271);
and U2452 (N_2452,N_2279,N_2347);
or U2453 (N_2453,N_2377,N_2394);
nor U2454 (N_2454,N_2295,N_2274);
or U2455 (N_2455,N_2376,N_2276);
or U2456 (N_2456,N_2261,N_2391);
xnor U2457 (N_2457,N_2342,N_2294);
nor U2458 (N_2458,N_2393,N_2358);
or U2459 (N_2459,N_2367,N_2382);
or U2460 (N_2460,N_2241,N_2266);
nor U2461 (N_2461,N_2213,N_2369);
or U2462 (N_2462,N_2307,N_2350);
or U2463 (N_2463,N_2255,N_2219);
xnor U2464 (N_2464,N_2203,N_2361);
xor U2465 (N_2465,N_2252,N_2225);
or U2466 (N_2466,N_2340,N_2304);
xnor U2467 (N_2467,N_2202,N_2345);
or U2468 (N_2468,N_2324,N_2283);
or U2469 (N_2469,N_2335,N_2204);
or U2470 (N_2470,N_2296,N_2285);
and U2471 (N_2471,N_2337,N_2322);
xor U2472 (N_2472,N_2260,N_2206);
nand U2473 (N_2473,N_2214,N_2378);
nand U2474 (N_2474,N_2329,N_2349);
xor U2475 (N_2475,N_2211,N_2287);
nor U2476 (N_2476,N_2235,N_2383);
xnor U2477 (N_2477,N_2201,N_2396);
nor U2478 (N_2478,N_2309,N_2330);
nor U2479 (N_2479,N_2216,N_2388);
or U2480 (N_2480,N_2319,N_2357);
nand U2481 (N_2481,N_2284,N_2385);
and U2482 (N_2482,N_2270,N_2354);
xnor U2483 (N_2483,N_2258,N_2268);
or U2484 (N_2484,N_2323,N_2293);
xnor U2485 (N_2485,N_2299,N_2397);
nor U2486 (N_2486,N_2251,N_2269);
or U2487 (N_2487,N_2390,N_2244);
nand U2488 (N_2488,N_2302,N_2288);
nand U2489 (N_2489,N_2263,N_2240);
nand U2490 (N_2490,N_2365,N_2242);
xnor U2491 (N_2491,N_2315,N_2360);
or U2492 (N_2492,N_2275,N_2308);
xnor U2493 (N_2493,N_2320,N_2359);
nor U2494 (N_2494,N_2249,N_2215);
and U2495 (N_2495,N_2212,N_2298);
nand U2496 (N_2496,N_2317,N_2239);
and U2497 (N_2497,N_2398,N_2246);
and U2498 (N_2498,N_2384,N_2380);
and U2499 (N_2499,N_2312,N_2209);
xnor U2500 (N_2500,N_2375,N_2255);
or U2501 (N_2501,N_2245,N_2349);
xnor U2502 (N_2502,N_2204,N_2373);
xor U2503 (N_2503,N_2258,N_2341);
or U2504 (N_2504,N_2337,N_2257);
or U2505 (N_2505,N_2333,N_2232);
nand U2506 (N_2506,N_2319,N_2276);
xnor U2507 (N_2507,N_2368,N_2366);
or U2508 (N_2508,N_2256,N_2367);
or U2509 (N_2509,N_2297,N_2328);
nand U2510 (N_2510,N_2244,N_2235);
nand U2511 (N_2511,N_2234,N_2245);
nand U2512 (N_2512,N_2398,N_2314);
xnor U2513 (N_2513,N_2216,N_2366);
and U2514 (N_2514,N_2359,N_2324);
and U2515 (N_2515,N_2246,N_2340);
xor U2516 (N_2516,N_2392,N_2263);
or U2517 (N_2517,N_2250,N_2371);
xnor U2518 (N_2518,N_2322,N_2233);
nand U2519 (N_2519,N_2378,N_2305);
nand U2520 (N_2520,N_2237,N_2352);
xnor U2521 (N_2521,N_2220,N_2376);
xor U2522 (N_2522,N_2204,N_2365);
and U2523 (N_2523,N_2278,N_2373);
nand U2524 (N_2524,N_2305,N_2391);
xor U2525 (N_2525,N_2204,N_2338);
nand U2526 (N_2526,N_2236,N_2315);
and U2527 (N_2527,N_2291,N_2285);
nand U2528 (N_2528,N_2282,N_2375);
xor U2529 (N_2529,N_2235,N_2377);
and U2530 (N_2530,N_2310,N_2263);
and U2531 (N_2531,N_2200,N_2345);
or U2532 (N_2532,N_2280,N_2206);
and U2533 (N_2533,N_2233,N_2256);
xor U2534 (N_2534,N_2329,N_2234);
nand U2535 (N_2535,N_2308,N_2390);
nand U2536 (N_2536,N_2320,N_2303);
and U2537 (N_2537,N_2399,N_2376);
xor U2538 (N_2538,N_2300,N_2314);
nand U2539 (N_2539,N_2369,N_2340);
and U2540 (N_2540,N_2327,N_2202);
and U2541 (N_2541,N_2316,N_2370);
xnor U2542 (N_2542,N_2305,N_2280);
or U2543 (N_2543,N_2395,N_2313);
xnor U2544 (N_2544,N_2204,N_2397);
or U2545 (N_2545,N_2387,N_2287);
or U2546 (N_2546,N_2243,N_2322);
nand U2547 (N_2547,N_2263,N_2377);
nand U2548 (N_2548,N_2215,N_2351);
nor U2549 (N_2549,N_2310,N_2362);
and U2550 (N_2550,N_2270,N_2221);
nand U2551 (N_2551,N_2221,N_2248);
xor U2552 (N_2552,N_2306,N_2339);
or U2553 (N_2553,N_2312,N_2314);
and U2554 (N_2554,N_2323,N_2328);
xor U2555 (N_2555,N_2327,N_2269);
nor U2556 (N_2556,N_2392,N_2386);
nor U2557 (N_2557,N_2391,N_2332);
or U2558 (N_2558,N_2295,N_2368);
or U2559 (N_2559,N_2253,N_2290);
and U2560 (N_2560,N_2221,N_2202);
and U2561 (N_2561,N_2390,N_2267);
or U2562 (N_2562,N_2299,N_2320);
xnor U2563 (N_2563,N_2242,N_2233);
xnor U2564 (N_2564,N_2383,N_2331);
nand U2565 (N_2565,N_2347,N_2271);
nor U2566 (N_2566,N_2203,N_2314);
xnor U2567 (N_2567,N_2346,N_2351);
or U2568 (N_2568,N_2221,N_2364);
or U2569 (N_2569,N_2246,N_2375);
nor U2570 (N_2570,N_2290,N_2222);
nand U2571 (N_2571,N_2268,N_2256);
xnor U2572 (N_2572,N_2246,N_2362);
xnor U2573 (N_2573,N_2387,N_2308);
and U2574 (N_2574,N_2398,N_2274);
xor U2575 (N_2575,N_2246,N_2343);
nand U2576 (N_2576,N_2371,N_2339);
xor U2577 (N_2577,N_2319,N_2390);
or U2578 (N_2578,N_2370,N_2296);
nor U2579 (N_2579,N_2372,N_2397);
and U2580 (N_2580,N_2377,N_2218);
and U2581 (N_2581,N_2222,N_2354);
nand U2582 (N_2582,N_2289,N_2281);
nor U2583 (N_2583,N_2343,N_2253);
and U2584 (N_2584,N_2281,N_2378);
xor U2585 (N_2585,N_2342,N_2322);
or U2586 (N_2586,N_2281,N_2288);
and U2587 (N_2587,N_2331,N_2286);
nor U2588 (N_2588,N_2328,N_2379);
xor U2589 (N_2589,N_2375,N_2223);
and U2590 (N_2590,N_2319,N_2226);
and U2591 (N_2591,N_2257,N_2284);
xor U2592 (N_2592,N_2389,N_2207);
nand U2593 (N_2593,N_2208,N_2242);
or U2594 (N_2594,N_2266,N_2251);
xor U2595 (N_2595,N_2393,N_2266);
nor U2596 (N_2596,N_2234,N_2238);
nand U2597 (N_2597,N_2250,N_2358);
and U2598 (N_2598,N_2370,N_2371);
nand U2599 (N_2599,N_2387,N_2334);
nand U2600 (N_2600,N_2524,N_2476);
xor U2601 (N_2601,N_2409,N_2456);
xnor U2602 (N_2602,N_2463,N_2418);
or U2603 (N_2603,N_2427,N_2421);
or U2604 (N_2604,N_2501,N_2483);
or U2605 (N_2605,N_2438,N_2484);
nor U2606 (N_2606,N_2434,N_2569);
or U2607 (N_2607,N_2440,N_2413);
and U2608 (N_2608,N_2449,N_2444);
nor U2609 (N_2609,N_2402,N_2499);
and U2610 (N_2610,N_2515,N_2598);
nor U2611 (N_2611,N_2417,N_2491);
nand U2612 (N_2612,N_2532,N_2591);
or U2613 (N_2613,N_2586,N_2445);
and U2614 (N_2614,N_2511,N_2459);
or U2615 (N_2615,N_2480,N_2432);
and U2616 (N_2616,N_2527,N_2549);
nor U2617 (N_2617,N_2462,N_2588);
and U2618 (N_2618,N_2519,N_2468);
and U2619 (N_2619,N_2494,N_2576);
or U2620 (N_2620,N_2573,N_2428);
and U2621 (N_2621,N_2521,N_2536);
or U2622 (N_2622,N_2448,N_2408);
or U2623 (N_2623,N_2572,N_2570);
and U2624 (N_2624,N_2506,N_2564);
xnor U2625 (N_2625,N_2581,N_2488);
nand U2626 (N_2626,N_2555,N_2400);
nor U2627 (N_2627,N_2443,N_2481);
and U2628 (N_2628,N_2487,N_2457);
xor U2629 (N_2629,N_2404,N_2552);
and U2630 (N_2630,N_2561,N_2442);
and U2631 (N_2631,N_2577,N_2550);
and U2632 (N_2632,N_2420,N_2568);
xor U2633 (N_2633,N_2415,N_2574);
and U2634 (N_2634,N_2493,N_2419);
nand U2635 (N_2635,N_2525,N_2430);
xnor U2636 (N_2636,N_2410,N_2567);
or U2637 (N_2637,N_2472,N_2575);
nor U2638 (N_2638,N_2422,N_2513);
xnor U2639 (N_2639,N_2553,N_2489);
and U2640 (N_2640,N_2450,N_2474);
nand U2641 (N_2641,N_2497,N_2473);
nor U2642 (N_2642,N_2543,N_2403);
or U2643 (N_2643,N_2423,N_2534);
nand U2644 (N_2644,N_2451,N_2594);
nand U2645 (N_2645,N_2469,N_2454);
nor U2646 (N_2646,N_2538,N_2530);
xor U2647 (N_2647,N_2475,N_2437);
nor U2648 (N_2648,N_2563,N_2592);
and U2649 (N_2649,N_2426,N_2556);
nor U2650 (N_2650,N_2495,N_2528);
or U2651 (N_2651,N_2508,N_2464);
nor U2652 (N_2652,N_2590,N_2560);
or U2653 (N_2653,N_2504,N_2579);
xnor U2654 (N_2654,N_2401,N_2535);
or U2655 (N_2655,N_2565,N_2412);
nor U2656 (N_2656,N_2599,N_2554);
nor U2657 (N_2657,N_2562,N_2539);
nor U2658 (N_2658,N_2496,N_2416);
nor U2659 (N_2659,N_2405,N_2447);
xnor U2660 (N_2660,N_2471,N_2557);
nor U2661 (N_2661,N_2465,N_2542);
nand U2662 (N_2662,N_2595,N_2478);
nand U2663 (N_2663,N_2516,N_2458);
xnor U2664 (N_2664,N_2584,N_2551);
nor U2665 (N_2665,N_2514,N_2547);
and U2666 (N_2666,N_2507,N_2452);
nor U2667 (N_2667,N_2531,N_2414);
nor U2668 (N_2668,N_2509,N_2441);
xnor U2669 (N_2669,N_2593,N_2470);
xnor U2670 (N_2670,N_2425,N_2461);
xor U2671 (N_2671,N_2518,N_2503);
and U2672 (N_2672,N_2431,N_2540);
xor U2673 (N_2673,N_2566,N_2429);
and U2674 (N_2674,N_2545,N_2436);
nand U2675 (N_2675,N_2485,N_2477);
or U2676 (N_2676,N_2479,N_2580);
xnor U2677 (N_2677,N_2541,N_2407);
or U2678 (N_2678,N_2498,N_2435);
or U2679 (N_2679,N_2433,N_2529);
nand U2680 (N_2680,N_2596,N_2411);
and U2681 (N_2681,N_2466,N_2585);
nor U2682 (N_2682,N_2486,N_2523);
nand U2683 (N_2683,N_2510,N_2597);
xnor U2684 (N_2684,N_2546,N_2548);
nand U2685 (N_2685,N_2455,N_2533);
or U2686 (N_2686,N_2439,N_2558);
xnor U2687 (N_2687,N_2453,N_2424);
nand U2688 (N_2688,N_2490,N_2406);
or U2689 (N_2689,N_2589,N_2446);
nor U2690 (N_2690,N_2505,N_2500);
xor U2691 (N_2691,N_2517,N_2537);
and U2692 (N_2692,N_2492,N_2544);
or U2693 (N_2693,N_2571,N_2526);
or U2694 (N_2694,N_2583,N_2582);
and U2695 (N_2695,N_2587,N_2467);
nand U2696 (N_2696,N_2578,N_2460);
and U2697 (N_2697,N_2482,N_2522);
nand U2698 (N_2698,N_2559,N_2502);
nand U2699 (N_2699,N_2520,N_2512);
nor U2700 (N_2700,N_2546,N_2496);
xnor U2701 (N_2701,N_2400,N_2413);
nor U2702 (N_2702,N_2589,N_2425);
or U2703 (N_2703,N_2452,N_2491);
and U2704 (N_2704,N_2451,N_2589);
nand U2705 (N_2705,N_2578,N_2568);
nor U2706 (N_2706,N_2527,N_2555);
xnor U2707 (N_2707,N_2474,N_2425);
nor U2708 (N_2708,N_2474,N_2563);
nand U2709 (N_2709,N_2497,N_2431);
nor U2710 (N_2710,N_2413,N_2436);
or U2711 (N_2711,N_2559,N_2578);
or U2712 (N_2712,N_2446,N_2510);
nor U2713 (N_2713,N_2549,N_2555);
xor U2714 (N_2714,N_2544,N_2528);
nand U2715 (N_2715,N_2507,N_2455);
nor U2716 (N_2716,N_2555,N_2481);
xor U2717 (N_2717,N_2518,N_2587);
nor U2718 (N_2718,N_2546,N_2420);
nor U2719 (N_2719,N_2504,N_2427);
nand U2720 (N_2720,N_2519,N_2450);
or U2721 (N_2721,N_2472,N_2406);
or U2722 (N_2722,N_2415,N_2473);
and U2723 (N_2723,N_2582,N_2408);
and U2724 (N_2724,N_2413,N_2471);
or U2725 (N_2725,N_2410,N_2514);
xnor U2726 (N_2726,N_2480,N_2497);
and U2727 (N_2727,N_2524,N_2465);
and U2728 (N_2728,N_2457,N_2437);
nand U2729 (N_2729,N_2477,N_2535);
and U2730 (N_2730,N_2562,N_2583);
nand U2731 (N_2731,N_2415,N_2520);
nand U2732 (N_2732,N_2574,N_2478);
or U2733 (N_2733,N_2449,N_2487);
or U2734 (N_2734,N_2455,N_2585);
nand U2735 (N_2735,N_2572,N_2450);
nand U2736 (N_2736,N_2577,N_2484);
xor U2737 (N_2737,N_2467,N_2454);
or U2738 (N_2738,N_2561,N_2407);
nor U2739 (N_2739,N_2432,N_2512);
xnor U2740 (N_2740,N_2493,N_2536);
and U2741 (N_2741,N_2574,N_2463);
xnor U2742 (N_2742,N_2534,N_2539);
nand U2743 (N_2743,N_2539,N_2451);
nand U2744 (N_2744,N_2477,N_2482);
or U2745 (N_2745,N_2577,N_2414);
nand U2746 (N_2746,N_2524,N_2571);
nor U2747 (N_2747,N_2423,N_2480);
xnor U2748 (N_2748,N_2471,N_2553);
nand U2749 (N_2749,N_2580,N_2474);
or U2750 (N_2750,N_2564,N_2524);
or U2751 (N_2751,N_2594,N_2563);
and U2752 (N_2752,N_2589,N_2405);
xnor U2753 (N_2753,N_2462,N_2503);
nand U2754 (N_2754,N_2570,N_2442);
and U2755 (N_2755,N_2408,N_2477);
nor U2756 (N_2756,N_2550,N_2574);
or U2757 (N_2757,N_2499,N_2451);
xor U2758 (N_2758,N_2591,N_2491);
xnor U2759 (N_2759,N_2566,N_2486);
and U2760 (N_2760,N_2529,N_2455);
and U2761 (N_2761,N_2430,N_2413);
nor U2762 (N_2762,N_2568,N_2436);
nor U2763 (N_2763,N_2436,N_2519);
nor U2764 (N_2764,N_2483,N_2457);
nor U2765 (N_2765,N_2473,N_2457);
xnor U2766 (N_2766,N_2420,N_2431);
or U2767 (N_2767,N_2434,N_2420);
xnor U2768 (N_2768,N_2540,N_2524);
xor U2769 (N_2769,N_2430,N_2445);
and U2770 (N_2770,N_2585,N_2506);
xnor U2771 (N_2771,N_2414,N_2505);
and U2772 (N_2772,N_2504,N_2487);
nor U2773 (N_2773,N_2579,N_2417);
and U2774 (N_2774,N_2579,N_2557);
and U2775 (N_2775,N_2563,N_2401);
nand U2776 (N_2776,N_2421,N_2446);
xor U2777 (N_2777,N_2487,N_2570);
nand U2778 (N_2778,N_2413,N_2485);
xnor U2779 (N_2779,N_2449,N_2535);
and U2780 (N_2780,N_2497,N_2468);
and U2781 (N_2781,N_2565,N_2575);
nor U2782 (N_2782,N_2584,N_2498);
xor U2783 (N_2783,N_2469,N_2566);
nand U2784 (N_2784,N_2524,N_2451);
nor U2785 (N_2785,N_2471,N_2430);
xnor U2786 (N_2786,N_2554,N_2574);
xor U2787 (N_2787,N_2567,N_2576);
and U2788 (N_2788,N_2424,N_2507);
nand U2789 (N_2789,N_2433,N_2552);
nor U2790 (N_2790,N_2416,N_2434);
nand U2791 (N_2791,N_2551,N_2527);
nor U2792 (N_2792,N_2554,N_2566);
or U2793 (N_2793,N_2509,N_2469);
nor U2794 (N_2794,N_2599,N_2484);
xnor U2795 (N_2795,N_2493,N_2503);
nand U2796 (N_2796,N_2516,N_2589);
nand U2797 (N_2797,N_2533,N_2440);
nand U2798 (N_2798,N_2455,N_2406);
nor U2799 (N_2799,N_2476,N_2561);
or U2800 (N_2800,N_2607,N_2699);
and U2801 (N_2801,N_2730,N_2705);
xor U2802 (N_2802,N_2748,N_2639);
or U2803 (N_2803,N_2709,N_2773);
or U2804 (N_2804,N_2728,N_2767);
and U2805 (N_2805,N_2660,N_2678);
nand U2806 (N_2806,N_2628,N_2691);
and U2807 (N_2807,N_2724,N_2722);
and U2808 (N_2808,N_2743,N_2623);
xnor U2809 (N_2809,N_2617,N_2631);
or U2810 (N_2810,N_2761,N_2770);
and U2811 (N_2811,N_2784,N_2642);
xnor U2812 (N_2812,N_2675,N_2774);
nand U2813 (N_2813,N_2794,N_2653);
xor U2814 (N_2814,N_2788,N_2713);
and U2815 (N_2815,N_2791,N_2654);
or U2816 (N_2816,N_2651,N_2627);
xor U2817 (N_2817,N_2674,N_2746);
or U2818 (N_2818,N_2650,N_2666);
xnor U2819 (N_2819,N_2669,N_2710);
nor U2820 (N_2820,N_2734,N_2630);
xor U2821 (N_2821,N_2667,N_2649);
xor U2822 (N_2822,N_2723,N_2759);
and U2823 (N_2823,N_2616,N_2643);
xnor U2824 (N_2824,N_2740,N_2779);
xnor U2825 (N_2825,N_2640,N_2638);
and U2826 (N_2826,N_2768,N_2787);
xnor U2827 (N_2827,N_2704,N_2727);
or U2828 (N_2828,N_2644,N_2656);
nand U2829 (N_2829,N_2696,N_2612);
or U2830 (N_2830,N_2742,N_2756);
xor U2831 (N_2831,N_2698,N_2786);
nor U2832 (N_2832,N_2738,N_2782);
nor U2833 (N_2833,N_2717,N_2732);
nor U2834 (N_2834,N_2697,N_2751);
xnor U2835 (N_2835,N_2601,N_2676);
and U2836 (N_2836,N_2690,N_2673);
nor U2837 (N_2837,N_2702,N_2711);
nand U2838 (N_2838,N_2677,N_2797);
nor U2839 (N_2839,N_2778,N_2629);
nor U2840 (N_2840,N_2754,N_2661);
nand U2841 (N_2841,N_2795,N_2634);
nor U2842 (N_2842,N_2610,N_2684);
and U2843 (N_2843,N_2613,N_2671);
or U2844 (N_2844,N_2731,N_2775);
or U2845 (N_2845,N_2659,N_2622);
xor U2846 (N_2846,N_2752,N_2672);
and U2847 (N_2847,N_2689,N_2688);
or U2848 (N_2848,N_2753,N_2658);
or U2849 (N_2849,N_2633,N_2685);
nor U2850 (N_2850,N_2632,N_2686);
nand U2851 (N_2851,N_2765,N_2747);
or U2852 (N_2852,N_2799,N_2624);
xnor U2853 (N_2853,N_2663,N_2647);
or U2854 (N_2854,N_2721,N_2655);
or U2855 (N_2855,N_2750,N_2762);
or U2856 (N_2856,N_2680,N_2602);
nand U2857 (N_2857,N_2668,N_2605);
nand U2858 (N_2858,N_2785,N_2700);
and U2859 (N_2859,N_2720,N_2687);
xor U2860 (N_2860,N_2789,N_2703);
and U2861 (N_2861,N_2739,N_2763);
or U2862 (N_2862,N_2606,N_2708);
xnor U2863 (N_2863,N_2764,N_2614);
and U2864 (N_2864,N_2693,N_2776);
nor U2865 (N_2865,N_2760,N_2652);
xor U2866 (N_2866,N_2603,N_2745);
xnor U2867 (N_2867,N_2625,N_2783);
and U2868 (N_2868,N_2604,N_2657);
or U2869 (N_2869,N_2611,N_2718);
and U2870 (N_2870,N_2757,N_2772);
nor U2871 (N_2871,N_2679,N_2769);
xnor U2872 (N_2872,N_2758,N_2798);
nor U2873 (N_2873,N_2744,N_2635);
nand U2874 (N_2874,N_2646,N_2790);
or U2875 (N_2875,N_2792,N_2636);
and U2876 (N_2876,N_2637,N_2777);
nor U2877 (N_2877,N_2715,N_2620);
nand U2878 (N_2878,N_2692,N_2716);
nand U2879 (N_2879,N_2741,N_2619);
nor U2880 (N_2880,N_2707,N_2755);
or U2881 (N_2881,N_2695,N_2683);
or U2882 (N_2882,N_2621,N_2670);
nor U2883 (N_2883,N_2706,N_2771);
or U2884 (N_2884,N_2648,N_2736);
nand U2885 (N_2885,N_2645,N_2626);
and U2886 (N_2886,N_2609,N_2793);
xor U2887 (N_2887,N_2681,N_2796);
xor U2888 (N_2888,N_2600,N_2729);
and U2889 (N_2889,N_2714,N_2781);
and U2890 (N_2890,N_2608,N_2725);
and U2891 (N_2891,N_2719,N_2665);
or U2892 (N_2892,N_2712,N_2780);
and U2893 (N_2893,N_2749,N_2701);
xnor U2894 (N_2894,N_2662,N_2726);
or U2895 (N_2895,N_2641,N_2735);
xnor U2896 (N_2896,N_2694,N_2733);
xnor U2897 (N_2897,N_2664,N_2737);
nor U2898 (N_2898,N_2618,N_2682);
xor U2899 (N_2899,N_2766,N_2615);
or U2900 (N_2900,N_2732,N_2634);
nand U2901 (N_2901,N_2627,N_2701);
and U2902 (N_2902,N_2749,N_2765);
or U2903 (N_2903,N_2655,N_2691);
xor U2904 (N_2904,N_2755,N_2682);
nand U2905 (N_2905,N_2708,N_2636);
nand U2906 (N_2906,N_2776,N_2684);
or U2907 (N_2907,N_2737,N_2774);
nand U2908 (N_2908,N_2643,N_2751);
nand U2909 (N_2909,N_2653,N_2665);
nor U2910 (N_2910,N_2664,N_2650);
or U2911 (N_2911,N_2787,N_2627);
nor U2912 (N_2912,N_2701,N_2664);
xnor U2913 (N_2913,N_2781,N_2791);
nand U2914 (N_2914,N_2795,N_2759);
and U2915 (N_2915,N_2611,N_2681);
xor U2916 (N_2916,N_2646,N_2771);
nand U2917 (N_2917,N_2782,N_2629);
or U2918 (N_2918,N_2638,N_2634);
and U2919 (N_2919,N_2666,N_2784);
or U2920 (N_2920,N_2614,N_2661);
xnor U2921 (N_2921,N_2672,N_2635);
nor U2922 (N_2922,N_2787,N_2625);
and U2923 (N_2923,N_2782,N_2692);
xor U2924 (N_2924,N_2676,N_2657);
or U2925 (N_2925,N_2636,N_2640);
and U2926 (N_2926,N_2748,N_2693);
xnor U2927 (N_2927,N_2643,N_2648);
xnor U2928 (N_2928,N_2677,N_2746);
or U2929 (N_2929,N_2736,N_2735);
xnor U2930 (N_2930,N_2657,N_2627);
nor U2931 (N_2931,N_2625,N_2718);
nor U2932 (N_2932,N_2722,N_2707);
xor U2933 (N_2933,N_2712,N_2677);
nand U2934 (N_2934,N_2716,N_2700);
xnor U2935 (N_2935,N_2643,N_2667);
or U2936 (N_2936,N_2605,N_2699);
nor U2937 (N_2937,N_2731,N_2626);
xnor U2938 (N_2938,N_2731,N_2718);
and U2939 (N_2939,N_2611,N_2749);
nand U2940 (N_2940,N_2643,N_2765);
and U2941 (N_2941,N_2751,N_2687);
or U2942 (N_2942,N_2758,N_2613);
and U2943 (N_2943,N_2697,N_2609);
xnor U2944 (N_2944,N_2607,N_2769);
or U2945 (N_2945,N_2711,N_2793);
nor U2946 (N_2946,N_2770,N_2607);
nand U2947 (N_2947,N_2628,N_2695);
nand U2948 (N_2948,N_2606,N_2735);
nor U2949 (N_2949,N_2751,N_2665);
or U2950 (N_2950,N_2617,N_2694);
nor U2951 (N_2951,N_2676,N_2710);
xnor U2952 (N_2952,N_2715,N_2784);
or U2953 (N_2953,N_2637,N_2683);
nand U2954 (N_2954,N_2771,N_2675);
nand U2955 (N_2955,N_2738,N_2727);
or U2956 (N_2956,N_2725,N_2799);
nor U2957 (N_2957,N_2608,N_2797);
xnor U2958 (N_2958,N_2604,N_2610);
xnor U2959 (N_2959,N_2680,N_2778);
nand U2960 (N_2960,N_2687,N_2703);
nand U2961 (N_2961,N_2763,N_2622);
and U2962 (N_2962,N_2713,N_2652);
and U2963 (N_2963,N_2799,N_2762);
nand U2964 (N_2964,N_2630,N_2779);
nor U2965 (N_2965,N_2733,N_2611);
nor U2966 (N_2966,N_2728,N_2684);
and U2967 (N_2967,N_2794,N_2783);
nand U2968 (N_2968,N_2724,N_2729);
or U2969 (N_2969,N_2790,N_2744);
or U2970 (N_2970,N_2643,N_2748);
and U2971 (N_2971,N_2661,N_2746);
nor U2972 (N_2972,N_2793,N_2612);
xnor U2973 (N_2973,N_2666,N_2703);
nor U2974 (N_2974,N_2600,N_2713);
xor U2975 (N_2975,N_2638,N_2677);
or U2976 (N_2976,N_2619,N_2660);
nand U2977 (N_2977,N_2621,N_2626);
and U2978 (N_2978,N_2621,N_2683);
and U2979 (N_2979,N_2719,N_2621);
and U2980 (N_2980,N_2723,N_2658);
nand U2981 (N_2981,N_2667,N_2732);
nor U2982 (N_2982,N_2784,N_2609);
and U2983 (N_2983,N_2790,N_2727);
nand U2984 (N_2984,N_2748,N_2753);
and U2985 (N_2985,N_2619,N_2787);
and U2986 (N_2986,N_2728,N_2754);
xor U2987 (N_2987,N_2731,N_2673);
and U2988 (N_2988,N_2725,N_2679);
and U2989 (N_2989,N_2789,N_2644);
or U2990 (N_2990,N_2604,N_2647);
nor U2991 (N_2991,N_2608,N_2721);
nor U2992 (N_2992,N_2650,N_2752);
nor U2993 (N_2993,N_2764,N_2702);
nand U2994 (N_2994,N_2645,N_2683);
nor U2995 (N_2995,N_2726,N_2722);
nand U2996 (N_2996,N_2773,N_2687);
and U2997 (N_2997,N_2605,N_2711);
nand U2998 (N_2998,N_2639,N_2737);
or U2999 (N_2999,N_2713,N_2702);
nand U3000 (N_3000,N_2915,N_2905);
nand U3001 (N_3001,N_2963,N_2892);
and U3002 (N_3002,N_2827,N_2847);
nor U3003 (N_3003,N_2875,N_2816);
nand U3004 (N_3004,N_2973,N_2840);
and U3005 (N_3005,N_2933,N_2980);
nand U3006 (N_3006,N_2971,N_2969);
and U3007 (N_3007,N_2812,N_2898);
or U3008 (N_3008,N_2859,N_2948);
nand U3009 (N_3009,N_2917,N_2823);
xnor U3010 (N_3010,N_2852,N_2965);
and U3011 (N_3011,N_2834,N_2990);
nand U3012 (N_3012,N_2931,N_2818);
or U3013 (N_3013,N_2983,N_2943);
and U3014 (N_3014,N_2803,N_2841);
nor U3015 (N_3015,N_2825,N_2872);
or U3016 (N_3016,N_2815,N_2853);
and U3017 (N_3017,N_2813,N_2972);
or U3018 (N_3018,N_2977,N_2838);
or U3019 (N_3019,N_2919,N_2927);
xnor U3020 (N_3020,N_2966,N_2949);
nand U3021 (N_3021,N_2806,N_2817);
and U3022 (N_3022,N_2962,N_2833);
and U3023 (N_3023,N_2975,N_2878);
nand U3024 (N_3024,N_2887,N_2894);
and U3025 (N_3025,N_2928,N_2809);
nor U3026 (N_3026,N_2985,N_2830);
xnor U3027 (N_3027,N_2924,N_2925);
xor U3028 (N_3028,N_2907,N_2845);
xnor U3029 (N_3029,N_2856,N_2921);
xor U3030 (N_3030,N_2916,N_2828);
or U3031 (N_3031,N_2993,N_2886);
or U3032 (N_3032,N_2920,N_2984);
nand U3033 (N_3033,N_2820,N_2836);
xor U3034 (N_3034,N_2938,N_2883);
or U3035 (N_3035,N_2944,N_2979);
and U3036 (N_3036,N_2939,N_2992);
xor U3037 (N_3037,N_2987,N_2849);
nor U3038 (N_3038,N_2868,N_2865);
nor U3039 (N_3039,N_2964,N_2897);
xor U3040 (N_3040,N_2810,N_2801);
xor U3041 (N_3041,N_2957,N_2857);
nand U3042 (N_3042,N_2945,N_2884);
and U3043 (N_3043,N_2807,N_2991);
xnor U3044 (N_3044,N_2954,N_2903);
and U3045 (N_3045,N_2960,N_2824);
xnor U3046 (N_3046,N_2906,N_2871);
nand U3047 (N_3047,N_2958,N_2974);
or U3048 (N_3048,N_2864,N_2885);
or U3049 (N_3049,N_2863,N_2937);
xor U3050 (N_3050,N_2837,N_2842);
nor U3051 (N_3051,N_2829,N_2870);
and U3052 (N_3052,N_2940,N_2831);
nand U3053 (N_3053,N_2844,N_2851);
and U3054 (N_3054,N_2946,N_2981);
xor U3055 (N_3055,N_2934,N_2876);
nor U3056 (N_3056,N_2880,N_2997);
or U3057 (N_3057,N_2947,N_2846);
nand U3058 (N_3058,N_2848,N_2976);
and U3059 (N_3059,N_2843,N_2996);
or U3060 (N_3060,N_2832,N_2804);
or U3061 (N_3061,N_2821,N_2978);
and U3062 (N_3062,N_2814,N_2802);
nor U3063 (N_3063,N_2936,N_2929);
or U3064 (N_3064,N_2900,N_2970);
and U3065 (N_3065,N_2994,N_2890);
and U3066 (N_3066,N_2858,N_2882);
and U3067 (N_3067,N_2896,N_2942);
nand U3068 (N_3068,N_2909,N_2999);
nand U3069 (N_3069,N_2826,N_2855);
or U3070 (N_3070,N_2891,N_2986);
xnor U3071 (N_3071,N_2959,N_2881);
xnor U3072 (N_3072,N_2901,N_2950);
xnor U3073 (N_3073,N_2819,N_2953);
and U3074 (N_3074,N_2808,N_2822);
nand U3075 (N_3075,N_2873,N_2926);
nand U3076 (N_3076,N_2805,N_2918);
xor U3077 (N_3077,N_2913,N_2968);
nand U3078 (N_3078,N_2862,N_2951);
and U3079 (N_3079,N_2860,N_2995);
and U3080 (N_3080,N_2893,N_2982);
xnor U3081 (N_3081,N_2952,N_2861);
xnor U3082 (N_3082,N_2889,N_2922);
and U3083 (N_3083,N_2961,N_2955);
or U3084 (N_3084,N_2989,N_2895);
xor U3085 (N_3085,N_2888,N_2850);
or U3086 (N_3086,N_2941,N_2879);
nor U3087 (N_3087,N_2854,N_2835);
and U3088 (N_3088,N_2967,N_2811);
nand U3089 (N_3089,N_2800,N_2932);
or U3090 (N_3090,N_2904,N_2923);
nor U3091 (N_3091,N_2908,N_2914);
nand U3092 (N_3092,N_2910,N_2912);
xnor U3093 (N_3093,N_2911,N_2867);
and U3094 (N_3094,N_2902,N_2988);
nand U3095 (N_3095,N_2839,N_2866);
or U3096 (N_3096,N_2869,N_2956);
or U3097 (N_3097,N_2935,N_2930);
or U3098 (N_3098,N_2899,N_2877);
xnor U3099 (N_3099,N_2998,N_2874);
and U3100 (N_3100,N_2885,N_2935);
nand U3101 (N_3101,N_2837,N_2979);
nor U3102 (N_3102,N_2979,N_2949);
and U3103 (N_3103,N_2817,N_2884);
or U3104 (N_3104,N_2990,N_2903);
and U3105 (N_3105,N_2832,N_2935);
nor U3106 (N_3106,N_2994,N_2816);
xor U3107 (N_3107,N_2995,N_2910);
nor U3108 (N_3108,N_2901,N_2878);
or U3109 (N_3109,N_2963,N_2851);
nand U3110 (N_3110,N_2975,N_2966);
and U3111 (N_3111,N_2958,N_2806);
xor U3112 (N_3112,N_2968,N_2879);
or U3113 (N_3113,N_2883,N_2966);
nand U3114 (N_3114,N_2912,N_2828);
or U3115 (N_3115,N_2973,N_2941);
xnor U3116 (N_3116,N_2975,N_2863);
xnor U3117 (N_3117,N_2918,N_2870);
and U3118 (N_3118,N_2946,N_2831);
xor U3119 (N_3119,N_2956,N_2939);
nand U3120 (N_3120,N_2924,N_2824);
or U3121 (N_3121,N_2892,N_2979);
nand U3122 (N_3122,N_2830,N_2896);
and U3123 (N_3123,N_2991,N_2914);
or U3124 (N_3124,N_2980,N_2880);
nor U3125 (N_3125,N_2843,N_2880);
xor U3126 (N_3126,N_2973,N_2989);
nand U3127 (N_3127,N_2827,N_2876);
or U3128 (N_3128,N_2901,N_2938);
nor U3129 (N_3129,N_2990,N_2897);
and U3130 (N_3130,N_2993,N_2848);
and U3131 (N_3131,N_2941,N_2810);
nand U3132 (N_3132,N_2863,N_2980);
and U3133 (N_3133,N_2835,N_2828);
xnor U3134 (N_3134,N_2863,N_2957);
or U3135 (N_3135,N_2926,N_2962);
or U3136 (N_3136,N_2858,N_2921);
or U3137 (N_3137,N_2988,N_2955);
xnor U3138 (N_3138,N_2881,N_2873);
nor U3139 (N_3139,N_2953,N_2829);
xor U3140 (N_3140,N_2955,N_2936);
and U3141 (N_3141,N_2922,N_2849);
xnor U3142 (N_3142,N_2896,N_2884);
and U3143 (N_3143,N_2897,N_2893);
nand U3144 (N_3144,N_2819,N_2861);
nor U3145 (N_3145,N_2901,N_2908);
or U3146 (N_3146,N_2866,N_2854);
nand U3147 (N_3147,N_2982,N_2831);
nand U3148 (N_3148,N_2896,N_2900);
and U3149 (N_3149,N_2880,N_2987);
xor U3150 (N_3150,N_2845,N_2851);
or U3151 (N_3151,N_2860,N_2881);
nor U3152 (N_3152,N_2880,N_2833);
xor U3153 (N_3153,N_2806,N_2811);
nor U3154 (N_3154,N_2931,N_2886);
and U3155 (N_3155,N_2956,N_2813);
xor U3156 (N_3156,N_2947,N_2912);
and U3157 (N_3157,N_2878,N_2857);
and U3158 (N_3158,N_2825,N_2875);
or U3159 (N_3159,N_2980,N_2814);
and U3160 (N_3160,N_2860,N_2867);
and U3161 (N_3161,N_2945,N_2812);
nor U3162 (N_3162,N_2966,N_2963);
and U3163 (N_3163,N_2979,N_2911);
xor U3164 (N_3164,N_2960,N_2803);
xor U3165 (N_3165,N_2948,N_2914);
nor U3166 (N_3166,N_2947,N_2875);
and U3167 (N_3167,N_2842,N_2990);
nand U3168 (N_3168,N_2841,N_2984);
or U3169 (N_3169,N_2987,N_2924);
nor U3170 (N_3170,N_2826,N_2829);
or U3171 (N_3171,N_2849,N_2865);
nand U3172 (N_3172,N_2950,N_2918);
xnor U3173 (N_3173,N_2810,N_2940);
and U3174 (N_3174,N_2965,N_2844);
xnor U3175 (N_3175,N_2982,N_2872);
xor U3176 (N_3176,N_2846,N_2845);
or U3177 (N_3177,N_2991,N_2943);
nor U3178 (N_3178,N_2932,N_2898);
and U3179 (N_3179,N_2803,N_2866);
nand U3180 (N_3180,N_2900,N_2876);
or U3181 (N_3181,N_2992,N_2931);
and U3182 (N_3182,N_2970,N_2901);
or U3183 (N_3183,N_2828,N_2906);
xor U3184 (N_3184,N_2955,N_2817);
or U3185 (N_3185,N_2821,N_2950);
nand U3186 (N_3186,N_2963,N_2845);
and U3187 (N_3187,N_2902,N_2804);
xnor U3188 (N_3188,N_2882,N_2836);
and U3189 (N_3189,N_2876,N_2821);
nand U3190 (N_3190,N_2843,N_2865);
and U3191 (N_3191,N_2968,N_2902);
and U3192 (N_3192,N_2873,N_2839);
nor U3193 (N_3193,N_2894,N_2906);
xor U3194 (N_3194,N_2838,N_2809);
xnor U3195 (N_3195,N_2932,N_2856);
or U3196 (N_3196,N_2879,N_2931);
or U3197 (N_3197,N_2912,N_2888);
xnor U3198 (N_3198,N_2897,N_2853);
or U3199 (N_3199,N_2876,N_2984);
or U3200 (N_3200,N_3165,N_3187);
nand U3201 (N_3201,N_3199,N_3119);
and U3202 (N_3202,N_3190,N_3186);
nand U3203 (N_3203,N_3167,N_3157);
xnor U3204 (N_3204,N_3063,N_3064);
nand U3205 (N_3205,N_3024,N_3079);
or U3206 (N_3206,N_3098,N_3151);
nand U3207 (N_3207,N_3074,N_3182);
nand U3208 (N_3208,N_3137,N_3006);
and U3209 (N_3209,N_3128,N_3011);
or U3210 (N_3210,N_3188,N_3016);
or U3211 (N_3211,N_3070,N_3061);
or U3212 (N_3212,N_3097,N_3022);
nand U3213 (N_3213,N_3082,N_3116);
or U3214 (N_3214,N_3034,N_3036);
nor U3215 (N_3215,N_3126,N_3004);
xor U3216 (N_3216,N_3175,N_3107);
or U3217 (N_3217,N_3065,N_3035);
nand U3218 (N_3218,N_3140,N_3158);
or U3219 (N_3219,N_3087,N_3124);
and U3220 (N_3220,N_3030,N_3010);
nand U3221 (N_3221,N_3162,N_3046);
nand U3222 (N_3222,N_3135,N_3147);
nor U3223 (N_3223,N_3038,N_3060);
nor U3224 (N_3224,N_3133,N_3156);
nand U3225 (N_3225,N_3054,N_3141);
nand U3226 (N_3226,N_3027,N_3000);
nor U3227 (N_3227,N_3076,N_3152);
or U3228 (N_3228,N_3192,N_3042);
and U3229 (N_3229,N_3005,N_3078);
xor U3230 (N_3230,N_3127,N_3026);
xnor U3231 (N_3231,N_3108,N_3164);
or U3232 (N_3232,N_3149,N_3049);
or U3233 (N_3233,N_3183,N_3168);
xnor U3234 (N_3234,N_3166,N_3086);
nand U3235 (N_3235,N_3075,N_3068);
nand U3236 (N_3236,N_3113,N_3132);
xor U3237 (N_3237,N_3172,N_3053);
or U3238 (N_3238,N_3146,N_3171);
or U3239 (N_3239,N_3109,N_3072);
xnor U3240 (N_3240,N_3160,N_3032);
xor U3241 (N_3241,N_3015,N_3031);
or U3242 (N_3242,N_3002,N_3196);
nand U3243 (N_3243,N_3048,N_3033);
and U3244 (N_3244,N_3096,N_3134);
nand U3245 (N_3245,N_3008,N_3111);
or U3246 (N_3246,N_3122,N_3067);
and U3247 (N_3247,N_3003,N_3130);
xnor U3248 (N_3248,N_3178,N_3050);
and U3249 (N_3249,N_3012,N_3103);
xnor U3250 (N_3250,N_3173,N_3161);
or U3251 (N_3251,N_3155,N_3117);
or U3252 (N_3252,N_3084,N_3057);
or U3253 (N_3253,N_3145,N_3189);
nor U3254 (N_3254,N_3052,N_3069);
or U3255 (N_3255,N_3013,N_3150);
nor U3256 (N_3256,N_3019,N_3176);
and U3257 (N_3257,N_3174,N_3101);
or U3258 (N_3258,N_3081,N_3062);
xor U3259 (N_3259,N_3138,N_3184);
xnor U3260 (N_3260,N_3073,N_3179);
nor U3261 (N_3261,N_3077,N_3115);
and U3262 (N_3262,N_3023,N_3114);
or U3263 (N_3263,N_3106,N_3009);
or U3264 (N_3264,N_3043,N_3102);
nor U3265 (N_3265,N_3112,N_3058);
nor U3266 (N_3266,N_3018,N_3191);
and U3267 (N_3267,N_3085,N_3039);
xnor U3268 (N_3268,N_3001,N_3025);
xor U3269 (N_3269,N_3080,N_3159);
nor U3270 (N_3270,N_3154,N_3088);
nor U3271 (N_3271,N_3095,N_3195);
xnor U3272 (N_3272,N_3047,N_3041);
nand U3273 (N_3273,N_3180,N_3017);
nand U3274 (N_3274,N_3177,N_3100);
xnor U3275 (N_3275,N_3198,N_3092);
or U3276 (N_3276,N_3037,N_3121);
and U3277 (N_3277,N_3056,N_3044);
nor U3278 (N_3278,N_3083,N_3129);
nor U3279 (N_3279,N_3125,N_3029);
xor U3280 (N_3280,N_3139,N_3194);
nand U3281 (N_3281,N_3144,N_3163);
or U3282 (N_3282,N_3120,N_3094);
nor U3283 (N_3283,N_3153,N_3020);
xnor U3284 (N_3284,N_3169,N_3007);
or U3285 (N_3285,N_3197,N_3028);
xor U3286 (N_3286,N_3066,N_3123);
nand U3287 (N_3287,N_3105,N_3143);
xnor U3288 (N_3288,N_3142,N_3014);
xor U3289 (N_3289,N_3131,N_3110);
and U3290 (N_3290,N_3090,N_3181);
xnor U3291 (N_3291,N_3136,N_3021);
nand U3292 (N_3292,N_3104,N_3099);
nand U3293 (N_3293,N_3093,N_3091);
nand U3294 (N_3294,N_3118,N_3170);
xnor U3295 (N_3295,N_3051,N_3040);
or U3296 (N_3296,N_3045,N_3148);
nor U3297 (N_3297,N_3193,N_3071);
and U3298 (N_3298,N_3059,N_3089);
xor U3299 (N_3299,N_3185,N_3055);
xnor U3300 (N_3300,N_3159,N_3072);
nand U3301 (N_3301,N_3159,N_3172);
and U3302 (N_3302,N_3014,N_3184);
or U3303 (N_3303,N_3048,N_3098);
nand U3304 (N_3304,N_3107,N_3055);
and U3305 (N_3305,N_3075,N_3188);
nor U3306 (N_3306,N_3017,N_3015);
nand U3307 (N_3307,N_3198,N_3171);
or U3308 (N_3308,N_3047,N_3036);
nor U3309 (N_3309,N_3098,N_3009);
nand U3310 (N_3310,N_3084,N_3070);
or U3311 (N_3311,N_3162,N_3031);
nand U3312 (N_3312,N_3179,N_3122);
and U3313 (N_3313,N_3126,N_3036);
nand U3314 (N_3314,N_3123,N_3036);
or U3315 (N_3315,N_3198,N_3022);
and U3316 (N_3316,N_3182,N_3020);
xor U3317 (N_3317,N_3055,N_3171);
nand U3318 (N_3318,N_3177,N_3111);
xnor U3319 (N_3319,N_3093,N_3117);
or U3320 (N_3320,N_3169,N_3013);
xnor U3321 (N_3321,N_3120,N_3130);
nor U3322 (N_3322,N_3122,N_3177);
xnor U3323 (N_3323,N_3130,N_3044);
and U3324 (N_3324,N_3102,N_3130);
xnor U3325 (N_3325,N_3164,N_3029);
nand U3326 (N_3326,N_3170,N_3133);
nor U3327 (N_3327,N_3157,N_3037);
and U3328 (N_3328,N_3094,N_3066);
and U3329 (N_3329,N_3175,N_3170);
nand U3330 (N_3330,N_3087,N_3028);
nand U3331 (N_3331,N_3131,N_3135);
and U3332 (N_3332,N_3084,N_3171);
and U3333 (N_3333,N_3133,N_3185);
nand U3334 (N_3334,N_3008,N_3089);
or U3335 (N_3335,N_3128,N_3138);
nand U3336 (N_3336,N_3097,N_3135);
or U3337 (N_3337,N_3131,N_3173);
and U3338 (N_3338,N_3016,N_3096);
or U3339 (N_3339,N_3167,N_3029);
nand U3340 (N_3340,N_3106,N_3157);
nor U3341 (N_3341,N_3074,N_3195);
and U3342 (N_3342,N_3060,N_3055);
nand U3343 (N_3343,N_3033,N_3139);
nor U3344 (N_3344,N_3130,N_3132);
xor U3345 (N_3345,N_3166,N_3147);
nand U3346 (N_3346,N_3101,N_3055);
xor U3347 (N_3347,N_3104,N_3180);
nor U3348 (N_3348,N_3109,N_3147);
nor U3349 (N_3349,N_3088,N_3175);
and U3350 (N_3350,N_3094,N_3130);
nor U3351 (N_3351,N_3174,N_3063);
xor U3352 (N_3352,N_3059,N_3002);
nand U3353 (N_3353,N_3159,N_3019);
nand U3354 (N_3354,N_3197,N_3180);
or U3355 (N_3355,N_3086,N_3071);
and U3356 (N_3356,N_3102,N_3047);
xnor U3357 (N_3357,N_3096,N_3061);
nand U3358 (N_3358,N_3097,N_3198);
nor U3359 (N_3359,N_3014,N_3036);
and U3360 (N_3360,N_3162,N_3178);
nand U3361 (N_3361,N_3086,N_3147);
nand U3362 (N_3362,N_3152,N_3151);
and U3363 (N_3363,N_3029,N_3094);
and U3364 (N_3364,N_3021,N_3105);
xor U3365 (N_3365,N_3092,N_3118);
and U3366 (N_3366,N_3112,N_3080);
and U3367 (N_3367,N_3193,N_3043);
nor U3368 (N_3368,N_3106,N_3056);
nand U3369 (N_3369,N_3158,N_3105);
nand U3370 (N_3370,N_3023,N_3153);
nand U3371 (N_3371,N_3084,N_3027);
nand U3372 (N_3372,N_3022,N_3160);
xnor U3373 (N_3373,N_3106,N_3122);
nor U3374 (N_3374,N_3058,N_3104);
nand U3375 (N_3375,N_3096,N_3179);
and U3376 (N_3376,N_3050,N_3185);
and U3377 (N_3377,N_3098,N_3089);
nor U3378 (N_3378,N_3019,N_3175);
nor U3379 (N_3379,N_3069,N_3061);
or U3380 (N_3380,N_3095,N_3109);
xor U3381 (N_3381,N_3095,N_3184);
nand U3382 (N_3382,N_3095,N_3106);
or U3383 (N_3383,N_3027,N_3157);
xnor U3384 (N_3384,N_3180,N_3096);
nor U3385 (N_3385,N_3082,N_3141);
nor U3386 (N_3386,N_3169,N_3128);
nor U3387 (N_3387,N_3123,N_3115);
or U3388 (N_3388,N_3096,N_3045);
nor U3389 (N_3389,N_3007,N_3109);
xor U3390 (N_3390,N_3192,N_3163);
and U3391 (N_3391,N_3154,N_3056);
or U3392 (N_3392,N_3192,N_3065);
xnor U3393 (N_3393,N_3045,N_3092);
xnor U3394 (N_3394,N_3063,N_3124);
nand U3395 (N_3395,N_3042,N_3044);
or U3396 (N_3396,N_3031,N_3087);
xnor U3397 (N_3397,N_3002,N_3178);
or U3398 (N_3398,N_3098,N_3034);
or U3399 (N_3399,N_3056,N_3164);
or U3400 (N_3400,N_3346,N_3378);
xnor U3401 (N_3401,N_3303,N_3365);
and U3402 (N_3402,N_3265,N_3398);
or U3403 (N_3403,N_3231,N_3310);
nor U3404 (N_3404,N_3308,N_3257);
and U3405 (N_3405,N_3215,N_3301);
xor U3406 (N_3406,N_3361,N_3382);
nand U3407 (N_3407,N_3349,N_3355);
nand U3408 (N_3408,N_3274,N_3395);
nor U3409 (N_3409,N_3287,N_3386);
or U3410 (N_3410,N_3311,N_3352);
and U3411 (N_3411,N_3342,N_3250);
xor U3412 (N_3412,N_3363,N_3201);
nor U3413 (N_3413,N_3279,N_3339);
nand U3414 (N_3414,N_3390,N_3353);
or U3415 (N_3415,N_3391,N_3240);
or U3416 (N_3416,N_3324,N_3221);
nor U3417 (N_3417,N_3229,N_3242);
and U3418 (N_3418,N_3225,N_3297);
or U3419 (N_3419,N_3243,N_3389);
xnor U3420 (N_3420,N_3347,N_3233);
nand U3421 (N_3421,N_3348,N_3202);
nand U3422 (N_3422,N_3337,N_3368);
or U3423 (N_3423,N_3372,N_3359);
nor U3424 (N_3424,N_3338,N_3350);
and U3425 (N_3425,N_3374,N_3321);
and U3426 (N_3426,N_3330,N_3376);
xnor U3427 (N_3427,N_3313,N_3219);
xor U3428 (N_3428,N_3369,N_3200);
or U3429 (N_3429,N_3248,N_3232);
nand U3430 (N_3430,N_3203,N_3305);
xor U3431 (N_3431,N_3283,N_3314);
or U3432 (N_3432,N_3299,N_3227);
nor U3433 (N_3433,N_3332,N_3343);
xor U3434 (N_3434,N_3317,N_3312);
xor U3435 (N_3435,N_3328,N_3370);
nand U3436 (N_3436,N_3254,N_3394);
or U3437 (N_3437,N_3286,N_3244);
or U3438 (N_3438,N_3335,N_3341);
nor U3439 (N_3439,N_3375,N_3280);
nand U3440 (N_3440,N_3253,N_3298);
xor U3441 (N_3441,N_3371,N_3320);
xor U3442 (N_3442,N_3327,N_3387);
or U3443 (N_3443,N_3292,N_3396);
or U3444 (N_3444,N_3304,N_3360);
xnor U3445 (N_3445,N_3358,N_3211);
nand U3446 (N_3446,N_3293,N_3294);
and U3447 (N_3447,N_3362,N_3307);
xnor U3448 (N_3448,N_3256,N_3315);
nand U3449 (N_3449,N_3384,N_3246);
and U3450 (N_3450,N_3356,N_3273);
xnor U3451 (N_3451,N_3357,N_3354);
nor U3452 (N_3452,N_3380,N_3345);
nand U3453 (N_3453,N_3290,N_3278);
nand U3454 (N_3454,N_3270,N_3210);
nand U3455 (N_3455,N_3269,N_3319);
xor U3456 (N_3456,N_3262,N_3222);
xnor U3457 (N_3457,N_3245,N_3306);
xor U3458 (N_3458,N_3255,N_3223);
nand U3459 (N_3459,N_3318,N_3272);
nand U3460 (N_3460,N_3238,N_3351);
and U3461 (N_3461,N_3316,N_3309);
nor U3462 (N_3462,N_3209,N_3331);
nor U3463 (N_3463,N_3336,N_3251);
or U3464 (N_3464,N_3226,N_3289);
nor U3465 (N_3465,N_3224,N_3241);
or U3466 (N_3466,N_3367,N_3260);
xnor U3467 (N_3467,N_3259,N_3267);
or U3468 (N_3468,N_3385,N_3239);
nand U3469 (N_3469,N_3217,N_3266);
nand U3470 (N_3470,N_3276,N_3268);
nand U3471 (N_3471,N_3291,N_3206);
xnor U3472 (N_3472,N_3261,N_3373);
and U3473 (N_3473,N_3204,N_3235);
and U3474 (N_3474,N_3399,N_3284);
nand U3475 (N_3475,N_3230,N_3205);
nand U3476 (N_3476,N_3302,N_3282);
and U3477 (N_3477,N_3300,N_3296);
nand U3478 (N_3478,N_3264,N_3249);
nor U3479 (N_3479,N_3218,N_3397);
and U3480 (N_3480,N_3285,N_3393);
nand U3481 (N_3481,N_3392,N_3258);
nor U3482 (N_3482,N_3252,N_3237);
or U3483 (N_3483,N_3220,N_3340);
nand U3484 (N_3484,N_3377,N_3247);
nand U3485 (N_3485,N_3383,N_3213);
nand U3486 (N_3486,N_3212,N_3275);
nor U3487 (N_3487,N_3234,N_3381);
and U3488 (N_3488,N_3322,N_3288);
nor U3489 (N_3489,N_3326,N_3333);
nand U3490 (N_3490,N_3329,N_3323);
nor U3491 (N_3491,N_3208,N_3281);
nor U3492 (N_3492,N_3344,N_3295);
or U3493 (N_3493,N_3216,N_3379);
and U3494 (N_3494,N_3325,N_3271);
xnor U3495 (N_3495,N_3207,N_3214);
and U3496 (N_3496,N_3334,N_3228);
nand U3497 (N_3497,N_3236,N_3263);
nor U3498 (N_3498,N_3366,N_3277);
and U3499 (N_3499,N_3388,N_3364);
or U3500 (N_3500,N_3393,N_3311);
xnor U3501 (N_3501,N_3255,N_3374);
nor U3502 (N_3502,N_3377,N_3237);
and U3503 (N_3503,N_3219,N_3384);
or U3504 (N_3504,N_3348,N_3248);
or U3505 (N_3505,N_3301,N_3281);
nand U3506 (N_3506,N_3221,N_3280);
and U3507 (N_3507,N_3261,N_3322);
xnor U3508 (N_3508,N_3312,N_3295);
nor U3509 (N_3509,N_3349,N_3218);
and U3510 (N_3510,N_3231,N_3393);
nand U3511 (N_3511,N_3280,N_3274);
xor U3512 (N_3512,N_3389,N_3324);
and U3513 (N_3513,N_3203,N_3389);
nand U3514 (N_3514,N_3300,N_3267);
and U3515 (N_3515,N_3314,N_3326);
or U3516 (N_3516,N_3385,N_3362);
xor U3517 (N_3517,N_3234,N_3202);
nor U3518 (N_3518,N_3330,N_3368);
nand U3519 (N_3519,N_3351,N_3333);
or U3520 (N_3520,N_3300,N_3313);
or U3521 (N_3521,N_3252,N_3310);
and U3522 (N_3522,N_3383,N_3354);
nand U3523 (N_3523,N_3279,N_3343);
nand U3524 (N_3524,N_3292,N_3397);
and U3525 (N_3525,N_3203,N_3382);
nor U3526 (N_3526,N_3267,N_3394);
and U3527 (N_3527,N_3258,N_3293);
xor U3528 (N_3528,N_3282,N_3313);
or U3529 (N_3529,N_3225,N_3382);
or U3530 (N_3530,N_3342,N_3273);
and U3531 (N_3531,N_3280,N_3247);
nor U3532 (N_3532,N_3382,N_3216);
or U3533 (N_3533,N_3395,N_3365);
or U3534 (N_3534,N_3367,N_3299);
and U3535 (N_3535,N_3339,N_3277);
and U3536 (N_3536,N_3298,N_3279);
nand U3537 (N_3537,N_3247,N_3329);
nor U3538 (N_3538,N_3250,N_3226);
and U3539 (N_3539,N_3235,N_3381);
nor U3540 (N_3540,N_3365,N_3263);
xor U3541 (N_3541,N_3349,N_3279);
and U3542 (N_3542,N_3340,N_3297);
nor U3543 (N_3543,N_3315,N_3224);
xnor U3544 (N_3544,N_3376,N_3265);
or U3545 (N_3545,N_3306,N_3334);
nor U3546 (N_3546,N_3326,N_3290);
nor U3547 (N_3547,N_3306,N_3282);
nor U3548 (N_3548,N_3207,N_3290);
xnor U3549 (N_3549,N_3306,N_3353);
or U3550 (N_3550,N_3306,N_3325);
or U3551 (N_3551,N_3352,N_3244);
nor U3552 (N_3552,N_3312,N_3373);
and U3553 (N_3553,N_3266,N_3265);
nor U3554 (N_3554,N_3205,N_3378);
xor U3555 (N_3555,N_3240,N_3265);
nor U3556 (N_3556,N_3304,N_3284);
and U3557 (N_3557,N_3323,N_3285);
nand U3558 (N_3558,N_3295,N_3358);
nor U3559 (N_3559,N_3239,N_3272);
nor U3560 (N_3560,N_3356,N_3249);
nand U3561 (N_3561,N_3206,N_3256);
nand U3562 (N_3562,N_3205,N_3393);
xnor U3563 (N_3563,N_3206,N_3204);
nor U3564 (N_3564,N_3313,N_3340);
nor U3565 (N_3565,N_3390,N_3310);
or U3566 (N_3566,N_3274,N_3296);
xor U3567 (N_3567,N_3297,N_3398);
xor U3568 (N_3568,N_3222,N_3216);
nor U3569 (N_3569,N_3237,N_3301);
and U3570 (N_3570,N_3295,N_3309);
and U3571 (N_3571,N_3315,N_3353);
and U3572 (N_3572,N_3252,N_3245);
or U3573 (N_3573,N_3222,N_3325);
or U3574 (N_3574,N_3282,N_3255);
or U3575 (N_3575,N_3331,N_3268);
nor U3576 (N_3576,N_3232,N_3309);
nand U3577 (N_3577,N_3214,N_3255);
or U3578 (N_3578,N_3314,N_3393);
or U3579 (N_3579,N_3347,N_3294);
nor U3580 (N_3580,N_3202,N_3246);
and U3581 (N_3581,N_3282,N_3275);
and U3582 (N_3582,N_3344,N_3329);
xnor U3583 (N_3583,N_3291,N_3361);
nand U3584 (N_3584,N_3368,N_3329);
nor U3585 (N_3585,N_3201,N_3252);
xor U3586 (N_3586,N_3306,N_3390);
and U3587 (N_3587,N_3209,N_3338);
or U3588 (N_3588,N_3327,N_3399);
nor U3589 (N_3589,N_3389,N_3296);
nand U3590 (N_3590,N_3350,N_3340);
nand U3591 (N_3591,N_3246,N_3286);
xnor U3592 (N_3592,N_3351,N_3347);
xnor U3593 (N_3593,N_3210,N_3291);
xor U3594 (N_3594,N_3232,N_3325);
or U3595 (N_3595,N_3291,N_3328);
nand U3596 (N_3596,N_3347,N_3339);
or U3597 (N_3597,N_3305,N_3249);
xnor U3598 (N_3598,N_3294,N_3217);
nand U3599 (N_3599,N_3356,N_3354);
xor U3600 (N_3600,N_3490,N_3525);
and U3601 (N_3601,N_3410,N_3509);
and U3602 (N_3602,N_3598,N_3495);
nor U3603 (N_3603,N_3431,N_3506);
or U3604 (N_3604,N_3422,N_3404);
nand U3605 (N_3605,N_3500,N_3520);
nand U3606 (N_3606,N_3524,N_3430);
xor U3607 (N_3607,N_3539,N_3538);
and U3608 (N_3608,N_3573,N_3474);
xnor U3609 (N_3609,N_3467,N_3477);
xnor U3610 (N_3610,N_3435,N_3546);
nor U3611 (N_3611,N_3476,N_3478);
nor U3612 (N_3612,N_3522,N_3423);
xor U3613 (N_3613,N_3559,N_3465);
nor U3614 (N_3614,N_3479,N_3408);
and U3615 (N_3615,N_3554,N_3584);
and U3616 (N_3616,N_3441,N_3402);
nor U3617 (N_3617,N_3472,N_3446);
xnor U3618 (N_3618,N_3510,N_3449);
nand U3619 (N_3619,N_3557,N_3492);
or U3620 (N_3620,N_3458,N_3594);
or U3621 (N_3621,N_3590,N_3589);
nand U3622 (N_3622,N_3537,N_3420);
xor U3623 (N_3623,N_3534,N_3542);
xnor U3624 (N_3624,N_3596,N_3443);
xor U3625 (N_3625,N_3580,N_3550);
and U3626 (N_3626,N_3581,N_3595);
and U3627 (N_3627,N_3496,N_3591);
nor U3628 (N_3628,N_3560,N_3406);
nand U3629 (N_3629,N_3526,N_3501);
or U3630 (N_3630,N_3517,N_3483);
or U3631 (N_3631,N_3558,N_3475);
xnor U3632 (N_3632,N_3400,N_3444);
nand U3633 (N_3633,N_3574,N_3487);
nand U3634 (N_3634,N_3507,N_3555);
nand U3635 (N_3635,N_3486,N_3417);
nand U3636 (N_3636,N_3535,N_3582);
nor U3637 (N_3637,N_3459,N_3513);
or U3638 (N_3638,N_3418,N_3426);
and U3639 (N_3639,N_3461,N_3586);
and U3640 (N_3640,N_3516,N_3540);
nand U3641 (N_3641,N_3434,N_3532);
and U3642 (N_3642,N_3407,N_3429);
nor U3643 (N_3643,N_3599,N_3549);
nand U3644 (N_3644,N_3468,N_3497);
nor U3645 (N_3645,N_3489,N_3587);
or U3646 (N_3646,N_3447,N_3541);
nor U3647 (N_3647,N_3412,N_3445);
nor U3648 (N_3648,N_3533,N_3564);
nand U3649 (N_3649,N_3428,N_3421);
nand U3650 (N_3650,N_3480,N_3503);
nand U3651 (N_3651,N_3519,N_3515);
nand U3652 (N_3652,N_3473,N_3561);
and U3653 (N_3653,N_3504,N_3572);
and U3654 (N_3654,N_3547,N_3579);
xnor U3655 (N_3655,N_3405,N_3482);
or U3656 (N_3656,N_3512,N_3562);
or U3657 (N_3657,N_3401,N_3457);
xnor U3658 (N_3658,N_3494,N_3593);
nand U3659 (N_3659,N_3552,N_3568);
nand U3660 (N_3660,N_3569,N_3553);
xnor U3661 (N_3661,N_3585,N_3448);
and U3662 (N_3662,N_3577,N_3518);
xnor U3663 (N_3663,N_3466,N_3427);
or U3664 (N_3664,N_3565,N_3484);
nor U3665 (N_3665,N_3460,N_3511);
and U3666 (N_3666,N_3415,N_3491);
and U3667 (N_3667,N_3536,N_3551);
and U3668 (N_3668,N_3416,N_3563);
nand U3669 (N_3669,N_3471,N_3424);
and U3670 (N_3670,N_3481,N_3456);
nor U3671 (N_3671,N_3493,N_3442);
nand U3672 (N_3672,N_3588,N_3543);
or U3673 (N_3673,N_3440,N_3498);
or U3674 (N_3674,N_3425,N_3502);
or U3675 (N_3675,N_3462,N_3527);
nor U3676 (N_3676,N_3545,N_3451);
xnor U3677 (N_3677,N_3469,N_3544);
or U3678 (N_3678,N_3488,N_3433);
nand U3679 (N_3679,N_3578,N_3531);
or U3680 (N_3680,N_3530,N_3499);
nor U3681 (N_3681,N_3528,N_3514);
or U3682 (N_3682,N_3597,N_3566);
nor U3683 (N_3683,N_3529,N_3485);
and U3684 (N_3684,N_3432,N_3438);
nor U3685 (N_3685,N_3414,N_3521);
xor U3686 (N_3686,N_3437,N_3413);
nor U3687 (N_3687,N_3453,N_3403);
or U3688 (N_3688,N_3576,N_3455);
nand U3689 (N_3689,N_3463,N_3452);
xnor U3690 (N_3690,N_3411,N_3450);
nand U3691 (N_3691,N_3439,N_3464);
nor U3692 (N_3692,N_3454,N_3436);
xor U3693 (N_3693,N_3567,N_3575);
nor U3694 (N_3694,N_3571,N_3548);
and U3695 (N_3695,N_3556,N_3419);
or U3696 (N_3696,N_3470,N_3505);
and U3697 (N_3697,N_3508,N_3583);
xnor U3698 (N_3698,N_3409,N_3592);
or U3699 (N_3699,N_3523,N_3570);
or U3700 (N_3700,N_3445,N_3437);
xor U3701 (N_3701,N_3577,N_3539);
and U3702 (N_3702,N_3437,N_3540);
nand U3703 (N_3703,N_3537,N_3524);
and U3704 (N_3704,N_3401,N_3449);
xor U3705 (N_3705,N_3546,N_3429);
nor U3706 (N_3706,N_3519,N_3547);
and U3707 (N_3707,N_3449,N_3525);
nor U3708 (N_3708,N_3426,N_3573);
or U3709 (N_3709,N_3494,N_3477);
and U3710 (N_3710,N_3505,N_3568);
nor U3711 (N_3711,N_3493,N_3431);
or U3712 (N_3712,N_3442,N_3418);
xor U3713 (N_3713,N_3505,N_3493);
xor U3714 (N_3714,N_3544,N_3555);
and U3715 (N_3715,N_3492,N_3530);
nand U3716 (N_3716,N_3424,N_3520);
nand U3717 (N_3717,N_3432,N_3412);
nand U3718 (N_3718,N_3541,N_3519);
nor U3719 (N_3719,N_3513,N_3458);
and U3720 (N_3720,N_3593,N_3441);
xor U3721 (N_3721,N_3582,N_3546);
and U3722 (N_3722,N_3596,N_3472);
or U3723 (N_3723,N_3494,N_3474);
nand U3724 (N_3724,N_3577,N_3415);
nor U3725 (N_3725,N_3512,N_3411);
xor U3726 (N_3726,N_3421,N_3426);
and U3727 (N_3727,N_3533,N_3531);
xor U3728 (N_3728,N_3485,N_3530);
nor U3729 (N_3729,N_3459,N_3564);
and U3730 (N_3730,N_3408,N_3461);
nand U3731 (N_3731,N_3516,N_3565);
and U3732 (N_3732,N_3566,N_3569);
nor U3733 (N_3733,N_3593,N_3472);
or U3734 (N_3734,N_3490,N_3411);
xnor U3735 (N_3735,N_3518,N_3401);
or U3736 (N_3736,N_3522,N_3550);
or U3737 (N_3737,N_3500,N_3545);
and U3738 (N_3738,N_3491,N_3599);
nor U3739 (N_3739,N_3595,N_3580);
xor U3740 (N_3740,N_3425,N_3446);
and U3741 (N_3741,N_3446,N_3522);
nand U3742 (N_3742,N_3564,N_3499);
nand U3743 (N_3743,N_3547,N_3558);
and U3744 (N_3744,N_3444,N_3439);
xnor U3745 (N_3745,N_3558,N_3430);
or U3746 (N_3746,N_3528,N_3535);
nor U3747 (N_3747,N_3516,N_3492);
xnor U3748 (N_3748,N_3578,N_3427);
xor U3749 (N_3749,N_3568,N_3565);
and U3750 (N_3750,N_3580,N_3402);
and U3751 (N_3751,N_3484,N_3492);
and U3752 (N_3752,N_3540,N_3490);
nand U3753 (N_3753,N_3550,N_3446);
nor U3754 (N_3754,N_3435,N_3480);
and U3755 (N_3755,N_3507,N_3471);
xor U3756 (N_3756,N_3473,N_3569);
xor U3757 (N_3757,N_3480,N_3411);
xnor U3758 (N_3758,N_3494,N_3512);
nand U3759 (N_3759,N_3504,N_3578);
or U3760 (N_3760,N_3477,N_3559);
xnor U3761 (N_3761,N_3562,N_3566);
nor U3762 (N_3762,N_3571,N_3498);
nand U3763 (N_3763,N_3581,N_3525);
and U3764 (N_3764,N_3573,N_3488);
xor U3765 (N_3765,N_3573,N_3445);
and U3766 (N_3766,N_3501,N_3417);
xor U3767 (N_3767,N_3466,N_3557);
xnor U3768 (N_3768,N_3532,N_3492);
and U3769 (N_3769,N_3420,N_3440);
or U3770 (N_3770,N_3532,N_3523);
and U3771 (N_3771,N_3409,N_3400);
and U3772 (N_3772,N_3417,N_3567);
nor U3773 (N_3773,N_3595,N_3499);
and U3774 (N_3774,N_3401,N_3592);
and U3775 (N_3775,N_3485,N_3467);
nor U3776 (N_3776,N_3473,N_3404);
and U3777 (N_3777,N_3426,N_3515);
nor U3778 (N_3778,N_3446,N_3481);
and U3779 (N_3779,N_3470,N_3525);
and U3780 (N_3780,N_3535,N_3487);
and U3781 (N_3781,N_3438,N_3417);
or U3782 (N_3782,N_3466,N_3485);
and U3783 (N_3783,N_3471,N_3591);
and U3784 (N_3784,N_3565,N_3444);
xor U3785 (N_3785,N_3456,N_3493);
or U3786 (N_3786,N_3552,N_3525);
nand U3787 (N_3787,N_3406,N_3531);
or U3788 (N_3788,N_3465,N_3591);
nand U3789 (N_3789,N_3478,N_3412);
nand U3790 (N_3790,N_3535,N_3558);
and U3791 (N_3791,N_3563,N_3560);
or U3792 (N_3792,N_3544,N_3421);
or U3793 (N_3793,N_3517,N_3571);
xor U3794 (N_3794,N_3402,N_3460);
xnor U3795 (N_3795,N_3517,N_3521);
nand U3796 (N_3796,N_3535,N_3443);
nand U3797 (N_3797,N_3591,N_3573);
and U3798 (N_3798,N_3556,N_3499);
or U3799 (N_3799,N_3563,N_3562);
and U3800 (N_3800,N_3766,N_3734);
nor U3801 (N_3801,N_3602,N_3746);
xnor U3802 (N_3802,N_3639,N_3617);
and U3803 (N_3803,N_3744,N_3687);
nand U3804 (N_3804,N_3729,N_3783);
and U3805 (N_3805,N_3647,N_3613);
or U3806 (N_3806,N_3761,N_3793);
and U3807 (N_3807,N_3656,N_3653);
or U3808 (N_3808,N_3696,N_3784);
nor U3809 (N_3809,N_3620,N_3727);
or U3810 (N_3810,N_3694,N_3777);
or U3811 (N_3811,N_3608,N_3663);
xor U3812 (N_3812,N_3673,N_3711);
xor U3813 (N_3813,N_3782,N_3741);
xor U3814 (N_3814,N_3728,N_3720);
nor U3815 (N_3815,N_3691,N_3632);
nor U3816 (N_3816,N_3775,N_3719);
nor U3817 (N_3817,N_3684,N_3667);
nand U3818 (N_3818,N_3699,N_3718);
nor U3819 (N_3819,N_3792,N_3754);
nand U3820 (N_3820,N_3797,N_3747);
nand U3821 (N_3821,N_3676,N_3655);
nor U3822 (N_3822,N_3654,N_3689);
nor U3823 (N_3823,N_3674,N_3749);
nand U3824 (N_3824,N_3764,N_3758);
xnor U3825 (N_3825,N_3600,N_3681);
xnor U3826 (N_3826,N_3604,N_3651);
nand U3827 (N_3827,N_3737,N_3657);
nand U3828 (N_3828,N_3751,N_3779);
xnor U3829 (N_3829,N_3706,N_3607);
nor U3830 (N_3830,N_3714,N_3743);
nand U3831 (N_3831,N_3759,N_3622);
and U3832 (N_3832,N_3789,N_3643);
or U3833 (N_3833,N_3703,N_3650);
or U3834 (N_3834,N_3715,N_3753);
xor U3835 (N_3835,N_3740,N_3637);
and U3836 (N_3836,N_3675,N_3610);
nand U3837 (N_3837,N_3660,N_3710);
or U3838 (N_3838,N_3733,N_3672);
or U3839 (N_3839,N_3773,N_3688);
nand U3840 (N_3840,N_3732,N_3636);
nand U3841 (N_3841,N_3736,N_3788);
or U3842 (N_3842,N_3731,N_3722);
xor U3843 (N_3843,N_3644,N_3770);
nor U3844 (N_3844,N_3790,N_3614);
nand U3845 (N_3845,N_3631,N_3763);
xor U3846 (N_3846,N_3630,N_3625);
or U3847 (N_3847,N_3616,N_3685);
or U3848 (N_3848,N_3641,N_3690);
nand U3849 (N_3849,N_3767,N_3799);
nand U3850 (N_3850,N_3633,N_3772);
xor U3851 (N_3851,N_3785,N_3635);
nor U3852 (N_3852,N_3760,N_3756);
or U3853 (N_3853,N_3748,N_3683);
nand U3854 (N_3854,N_3662,N_3723);
or U3855 (N_3855,N_3626,N_3665);
nor U3856 (N_3856,N_3709,N_3750);
nand U3857 (N_3857,N_3780,N_3730);
nor U3858 (N_3858,N_3752,N_3671);
nand U3859 (N_3859,N_3680,N_3678);
nor U3860 (N_3860,N_3682,N_3794);
nand U3861 (N_3861,N_3717,N_3716);
nor U3862 (N_3862,N_3796,N_3670);
xor U3863 (N_3863,N_3742,N_3726);
and U3864 (N_3864,N_3781,N_3621);
nor U3865 (N_3865,N_3755,N_3798);
or U3866 (N_3866,N_3679,N_3700);
xnor U3867 (N_3867,N_3795,N_3661);
or U3868 (N_3868,N_3762,N_3629);
and U3869 (N_3869,N_3765,N_3768);
and U3870 (N_3870,N_3771,N_3738);
xnor U3871 (N_3871,N_3618,N_3669);
nand U3872 (N_3872,N_3692,N_3739);
and U3873 (N_3873,N_3712,N_3615);
nor U3874 (N_3874,N_3713,N_3778);
nand U3875 (N_3875,N_3638,N_3724);
nand U3876 (N_3876,N_3708,N_3704);
or U3877 (N_3877,N_3611,N_3686);
or U3878 (N_3878,N_3666,N_3645);
xnor U3879 (N_3879,N_3725,N_3701);
nor U3880 (N_3880,N_3745,N_3609);
nand U3881 (N_3881,N_3702,N_3627);
or U3882 (N_3882,N_3791,N_3658);
and U3883 (N_3883,N_3640,N_3769);
nand U3884 (N_3884,N_3659,N_3735);
and U3885 (N_3885,N_3646,N_3757);
xor U3886 (N_3886,N_3787,N_3786);
and U3887 (N_3887,N_3695,N_3668);
xnor U3888 (N_3888,N_3612,N_3605);
or U3889 (N_3889,N_3619,N_3624);
xnor U3890 (N_3890,N_3677,N_3606);
nand U3891 (N_3891,N_3634,N_3721);
nand U3892 (N_3892,N_3649,N_3705);
nand U3893 (N_3893,N_3776,N_3601);
nor U3894 (N_3894,N_3642,N_3707);
nand U3895 (N_3895,N_3698,N_3774);
or U3896 (N_3896,N_3693,N_3628);
and U3897 (N_3897,N_3623,N_3652);
and U3898 (N_3898,N_3697,N_3648);
xor U3899 (N_3899,N_3664,N_3603);
nand U3900 (N_3900,N_3635,N_3673);
nand U3901 (N_3901,N_3625,N_3644);
nand U3902 (N_3902,N_3709,N_3726);
nand U3903 (N_3903,N_3600,N_3740);
xor U3904 (N_3904,N_3702,N_3717);
xor U3905 (N_3905,N_3709,N_3680);
xor U3906 (N_3906,N_3791,N_3752);
and U3907 (N_3907,N_3781,N_3714);
or U3908 (N_3908,N_3642,N_3684);
nand U3909 (N_3909,N_3767,N_3772);
nor U3910 (N_3910,N_3634,N_3607);
nand U3911 (N_3911,N_3622,N_3787);
xor U3912 (N_3912,N_3790,N_3759);
and U3913 (N_3913,N_3711,N_3627);
nor U3914 (N_3914,N_3661,N_3797);
nand U3915 (N_3915,N_3703,N_3630);
and U3916 (N_3916,N_3772,N_3687);
xor U3917 (N_3917,N_3624,N_3788);
nand U3918 (N_3918,N_3710,N_3636);
xor U3919 (N_3919,N_3655,N_3725);
or U3920 (N_3920,N_3600,N_3799);
nand U3921 (N_3921,N_3723,N_3620);
or U3922 (N_3922,N_3728,N_3724);
nand U3923 (N_3923,N_3685,N_3633);
nand U3924 (N_3924,N_3617,N_3647);
or U3925 (N_3925,N_3695,N_3641);
nand U3926 (N_3926,N_3679,N_3790);
and U3927 (N_3927,N_3769,N_3783);
nor U3928 (N_3928,N_3640,N_3721);
nand U3929 (N_3929,N_3665,N_3786);
or U3930 (N_3930,N_3713,N_3731);
xor U3931 (N_3931,N_3655,N_3636);
nand U3932 (N_3932,N_3752,N_3761);
nor U3933 (N_3933,N_3735,N_3639);
xnor U3934 (N_3934,N_3789,N_3719);
nor U3935 (N_3935,N_3734,N_3790);
nor U3936 (N_3936,N_3643,N_3767);
or U3937 (N_3937,N_3773,N_3649);
nand U3938 (N_3938,N_3793,N_3769);
nand U3939 (N_3939,N_3667,N_3789);
or U3940 (N_3940,N_3641,N_3775);
or U3941 (N_3941,N_3642,N_3659);
nor U3942 (N_3942,N_3623,N_3799);
and U3943 (N_3943,N_3741,N_3680);
or U3944 (N_3944,N_3631,N_3665);
nor U3945 (N_3945,N_3612,N_3792);
nor U3946 (N_3946,N_3682,N_3676);
nand U3947 (N_3947,N_3721,N_3605);
or U3948 (N_3948,N_3725,N_3732);
and U3949 (N_3949,N_3619,N_3792);
nand U3950 (N_3950,N_3746,N_3714);
nand U3951 (N_3951,N_3630,N_3600);
nand U3952 (N_3952,N_3725,N_3727);
or U3953 (N_3953,N_3775,N_3750);
and U3954 (N_3954,N_3604,N_3768);
xnor U3955 (N_3955,N_3760,N_3617);
and U3956 (N_3956,N_3604,N_3608);
nor U3957 (N_3957,N_3668,N_3683);
xor U3958 (N_3958,N_3648,N_3662);
xnor U3959 (N_3959,N_3646,N_3653);
or U3960 (N_3960,N_3764,N_3627);
nor U3961 (N_3961,N_3792,N_3613);
nand U3962 (N_3962,N_3683,N_3792);
or U3963 (N_3963,N_3665,N_3624);
or U3964 (N_3964,N_3792,N_3776);
or U3965 (N_3965,N_3636,N_3717);
xnor U3966 (N_3966,N_3702,N_3672);
nand U3967 (N_3967,N_3672,N_3784);
nand U3968 (N_3968,N_3662,N_3795);
xor U3969 (N_3969,N_3666,N_3711);
nor U3970 (N_3970,N_3750,N_3724);
xor U3971 (N_3971,N_3723,N_3792);
or U3972 (N_3972,N_3626,N_3755);
and U3973 (N_3973,N_3740,N_3755);
nand U3974 (N_3974,N_3664,N_3712);
xnor U3975 (N_3975,N_3615,N_3718);
nor U3976 (N_3976,N_3754,N_3659);
or U3977 (N_3977,N_3771,N_3656);
nor U3978 (N_3978,N_3720,N_3779);
nor U3979 (N_3979,N_3733,N_3671);
nor U3980 (N_3980,N_3636,N_3762);
or U3981 (N_3981,N_3711,N_3756);
or U3982 (N_3982,N_3627,N_3758);
or U3983 (N_3983,N_3643,N_3741);
xnor U3984 (N_3984,N_3638,N_3709);
and U3985 (N_3985,N_3797,N_3649);
nand U3986 (N_3986,N_3742,N_3738);
nor U3987 (N_3987,N_3604,N_3741);
nor U3988 (N_3988,N_3735,N_3720);
nor U3989 (N_3989,N_3670,N_3777);
and U3990 (N_3990,N_3711,N_3606);
nor U3991 (N_3991,N_3768,N_3712);
xor U3992 (N_3992,N_3655,N_3621);
xnor U3993 (N_3993,N_3652,N_3710);
xor U3994 (N_3994,N_3669,N_3652);
nor U3995 (N_3995,N_3696,N_3781);
xnor U3996 (N_3996,N_3730,N_3754);
xor U3997 (N_3997,N_3635,N_3630);
xnor U3998 (N_3998,N_3782,N_3763);
xor U3999 (N_3999,N_3756,N_3765);
nor U4000 (N_4000,N_3865,N_3950);
or U4001 (N_4001,N_3901,N_3947);
nor U4002 (N_4002,N_3908,N_3927);
or U4003 (N_4003,N_3864,N_3866);
nor U4004 (N_4004,N_3831,N_3931);
nor U4005 (N_4005,N_3982,N_3938);
xnor U4006 (N_4006,N_3909,N_3890);
nand U4007 (N_4007,N_3948,N_3945);
nor U4008 (N_4008,N_3887,N_3895);
nor U4009 (N_4009,N_3924,N_3983);
and U4010 (N_4010,N_3834,N_3861);
and U4011 (N_4011,N_3906,N_3801);
or U4012 (N_4012,N_3886,N_3943);
xnor U4013 (N_4013,N_3879,N_3874);
xor U4014 (N_4014,N_3851,N_3921);
and U4015 (N_4015,N_3941,N_3899);
xnor U4016 (N_4016,N_3936,N_3920);
nand U4017 (N_4017,N_3842,N_3970);
nor U4018 (N_4018,N_3824,N_3823);
xor U4019 (N_4019,N_3848,N_3857);
nor U4020 (N_4020,N_3869,N_3986);
or U4021 (N_4021,N_3944,N_3872);
and U4022 (N_4022,N_3889,N_3868);
and U4023 (N_4023,N_3997,N_3891);
and U4024 (N_4024,N_3978,N_3998);
and U4025 (N_4025,N_3989,N_3979);
nor U4026 (N_4026,N_3856,N_3883);
xnor U4027 (N_4027,N_3835,N_3917);
and U4028 (N_4028,N_3934,N_3907);
and U4029 (N_4029,N_3905,N_3830);
and U4030 (N_4030,N_3845,N_3987);
nor U4031 (N_4031,N_3815,N_3802);
nor U4032 (N_4032,N_3993,N_3942);
nor U4033 (N_4033,N_3820,N_3980);
and U4034 (N_4034,N_3958,N_3962);
xnor U4035 (N_4035,N_3839,N_3892);
nand U4036 (N_4036,N_3984,N_3885);
nor U4037 (N_4037,N_3976,N_3898);
or U4038 (N_4038,N_3825,N_3849);
or U4039 (N_4039,N_3952,N_3928);
nor U4040 (N_4040,N_3903,N_3914);
nand U4041 (N_4041,N_3965,N_3822);
xnor U4042 (N_4042,N_3964,N_3996);
and U4043 (N_4043,N_3813,N_3946);
nor U4044 (N_4044,N_3951,N_3988);
and U4045 (N_4045,N_3841,N_3949);
nand U4046 (N_4046,N_3873,N_3860);
nand U4047 (N_4047,N_3992,N_3811);
nor U4048 (N_4048,N_3960,N_3884);
nand U4049 (N_4049,N_3910,N_3990);
nor U4050 (N_4050,N_3827,N_3816);
xor U4051 (N_4051,N_3821,N_3863);
nor U4052 (N_4052,N_3806,N_3922);
nor U4053 (N_4053,N_3878,N_3862);
and U4054 (N_4054,N_3858,N_3955);
nand U4055 (N_4055,N_3853,N_3888);
or U4056 (N_4056,N_3926,N_3840);
or U4057 (N_4057,N_3995,N_3912);
nand U4058 (N_4058,N_3900,N_3854);
or U4059 (N_4059,N_3867,N_3800);
or U4060 (N_4060,N_3843,N_3870);
and U4061 (N_4061,N_3894,N_3953);
xnor U4062 (N_4062,N_3919,N_3836);
nand U4063 (N_4063,N_3959,N_3805);
and U4064 (N_4064,N_3932,N_3880);
xor U4065 (N_4065,N_3975,N_3994);
or U4066 (N_4066,N_3810,N_3833);
or U4067 (N_4067,N_3913,N_3881);
nor U4068 (N_4068,N_3882,N_3846);
and U4069 (N_4069,N_3859,N_3916);
and U4070 (N_4070,N_3929,N_3966);
nor U4071 (N_4071,N_3818,N_3902);
xnor U4072 (N_4072,N_3933,N_3939);
nand U4073 (N_4073,N_3808,N_3829);
nor U4074 (N_4074,N_3855,N_3973);
and U4075 (N_4075,N_3968,N_3875);
and U4076 (N_4076,N_3850,N_3918);
and U4077 (N_4077,N_3972,N_3826);
and U4078 (N_4078,N_3961,N_3925);
nor U4079 (N_4079,N_3803,N_3935);
xnor U4080 (N_4080,N_3915,N_3974);
xor U4081 (N_4081,N_3963,N_3871);
nor U4082 (N_4082,N_3911,N_3957);
nor U4083 (N_4083,N_3847,N_3940);
nor U4084 (N_4084,N_3991,N_3828);
or U4085 (N_4085,N_3930,N_3852);
nand U4086 (N_4086,N_3904,N_3923);
nand U4087 (N_4087,N_3937,N_3876);
or U4088 (N_4088,N_3804,N_3999);
nand U4089 (N_4089,N_3954,N_3832);
nor U4090 (N_4090,N_3814,N_3893);
or U4091 (N_4091,N_3812,N_3971);
and U4092 (N_4092,N_3844,N_3956);
and U4093 (N_4093,N_3981,N_3819);
nor U4094 (N_4094,N_3897,N_3877);
nor U4095 (N_4095,N_3837,N_3809);
xor U4096 (N_4096,N_3967,N_3817);
or U4097 (N_4097,N_3985,N_3807);
nor U4098 (N_4098,N_3838,N_3896);
nor U4099 (N_4099,N_3969,N_3977);
and U4100 (N_4100,N_3968,N_3808);
nor U4101 (N_4101,N_3955,N_3884);
and U4102 (N_4102,N_3833,N_3912);
and U4103 (N_4103,N_3970,N_3813);
or U4104 (N_4104,N_3840,N_3807);
and U4105 (N_4105,N_3845,N_3814);
and U4106 (N_4106,N_3934,N_3855);
nor U4107 (N_4107,N_3840,N_3866);
nor U4108 (N_4108,N_3931,N_3939);
and U4109 (N_4109,N_3923,N_3896);
nand U4110 (N_4110,N_3805,N_3811);
nand U4111 (N_4111,N_3874,N_3930);
and U4112 (N_4112,N_3901,N_3928);
and U4113 (N_4113,N_3907,N_3896);
xnor U4114 (N_4114,N_3916,N_3899);
or U4115 (N_4115,N_3984,N_3830);
xnor U4116 (N_4116,N_3957,N_3819);
and U4117 (N_4117,N_3856,N_3934);
nor U4118 (N_4118,N_3985,N_3949);
or U4119 (N_4119,N_3894,N_3969);
nor U4120 (N_4120,N_3988,N_3838);
nand U4121 (N_4121,N_3993,N_3983);
nor U4122 (N_4122,N_3934,N_3860);
or U4123 (N_4123,N_3888,N_3933);
xnor U4124 (N_4124,N_3888,N_3823);
and U4125 (N_4125,N_3882,N_3899);
nand U4126 (N_4126,N_3957,N_3961);
nor U4127 (N_4127,N_3900,N_3828);
nor U4128 (N_4128,N_3886,N_3961);
xor U4129 (N_4129,N_3878,N_3843);
nor U4130 (N_4130,N_3982,N_3875);
and U4131 (N_4131,N_3974,N_3848);
and U4132 (N_4132,N_3886,N_3858);
and U4133 (N_4133,N_3847,N_3852);
nor U4134 (N_4134,N_3805,N_3847);
and U4135 (N_4135,N_3888,N_3909);
and U4136 (N_4136,N_3982,N_3991);
nand U4137 (N_4137,N_3890,N_3836);
xnor U4138 (N_4138,N_3841,N_3895);
nor U4139 (N_4139,N_3899,N_3906);
or U4140 (N_4140,N_3870,N_3844);
nand U4141 (N_4141,N_3979,N_3984);
nand U4142 (N_4142,N_3866,N_3958);
xor U4143 (N_4143,N_3847,N_3811);
or U4144 (N_4144,N_3867,N_3834);
nor U4145 (N_4145,N_3992,N_3978);
or U4146 (N_4146,N_3889,N_3846);
or U4147 (N_4147,N_3906,N_3861);
xnor U4148 (N_4148,N_3940,N_3865);
nand U4149 (N_4149,N_3869,N_3827);
nor U4150 (N_4150,N_3999,N_3918);
xor U4151 (N_4151,N_3819,N_3837);
nand U4152 (N_4152,N_3883,N_3859);
or U4153 (N_4153,N_3869,N_3862);
and U4154 (N_4154,N_3865,N_3920);
nand U4155 (N_4155,N_3983,N_3887);
or U4156 (N_4156,N_3826,N_3892);
or U4157 (N_4157,N_3877,N_3863);
nand U4158 (N_4158,N_3860,N_3970);
and U4159 (N_4159,N_3914,N_3808);
xnor U4160 (N_4160,N_3966,N_3985);
and U4161 (N_4161,N_3810,N_3947);
nor U4162 (N_4162,N_3869,N_3924);
and U4163 (N_4163,N_3804,N_3831);
xnor U4164 (N_4164,N_3949,N_3911);
or U4165 (N_4165,N_3823,N_3843);
nor U4166 (N_4166,N_3908,N_3896);
or U4167 (N_4167,N_3986,N_3964);
nor U4168 (N_4168,N_3960,N_3842);
nor U4169 (N_4169,N_3926,N_3814);
xnor U4170 (N_4170,N_3991,N_3987);
nand U4171 (N_4171,N_3870,N_3863);
and U4172 (N_4172,N_3813,N_3888);
and U4173 (N_4173,N_3936,N_3930);
xnor U4174 (N_4174,N_3902,N_3800);
nor U4175 (N_4175,N_3823,N_3913);
and U4176 (N_4176,N_3806,N_3921);
nor U4177 (N_4177,N_3857,N_3902);
nor U4178 (N_4178,N_3824,N_3810);
or U4179 (N_4179,N_3880,N_3804);
and U4180 (N_4180,N_3939,N_3823);
and U4181 (N_4181,N_3983,N_3874);
xor U4182 (N_4182,N_3944,N_3992);
nor U4183 (N_4183,N_3842,N_3893);
nand U4184 (N_4184,N_3958,N_3983);
or U4185 (N_4185,N_3865,N_3986);
or U4186 (N_4186,N_3908,N_3924);
and U4187 (N_4187,N_3969,N_3961);
nand U4188 (N_4188,N_3947,N_3912);
xor U4189 (N_4189,N_3910,N_3839);
xnor U4190 (N_4190,N_3813,N_3885);
nor U4191 (N_4191,N_3907,N_3972);
and U4192 (N_4192,N_3802,N_3990);
nor U4193 (N_4193,N_3814,N_3962);
and U4194 (N_4194,N_3877,N_3987);
xor U4195 (N_4195,N_3811,N_3841);
nor U4196 (N_4196,N_3981,N_3973);
nor U4197 (N_4197,N_3985,N_3880);
nand U4198 (N_4198,N_3908,N_3930);
and U4199 (N_4199,N_3936,N_3889);
nand U4200 (N_4200,N_4144,N_4100);
or U4201 (N_4201,N_4102,N_4186);
nor U4202 (N_4202,N_4106,N_4179);
xnor U4203 (N_4203,N_4030,N_4156);
nor U4204 (N_4204,N_4183,N_4173);
xor U4205 (N_4205,N_4066,N_4035);
xor U4206 (N_4206,N_4111,N_4010);
nand U4207 (N_4207,N_4161,N_4051);
and U4208 (N_4208,N_4145,N_4047);
or U4209 (N_4209,N_4184,N_4107);
nor U4210 (N_4210,N_4089,N_4048);
or U4211 (N_4211,N_4121,N_4068);
xnor U4212 (N_4212,N_4151,N_4056);
and U4213 (N_4213,N_4191,N_4170);
or U4214 (N_4214,N_4165,N_4076);
nor U4215 (N_4215,N_4028,N_4070);
or U4216 (N_4216,N_4124,N_4116);
nor U4217 (N_4217,N_4109,N_4013);
or U4218 (N_4218,N_4099,N_4069);
nand U4219 (N_4219,N_4163,N_4188);
or U4220 (N_4220,N_4172,N_4060);
nand U4221 (N_4221,N_4079,N_4101);
or U4222 (N_4222,N_4143,N_4132);
and U4223 (N_4223,N_4136,N_4192);
xor U4224 (N_4224,N_4095,N_4131);
nand U4225 (N_4225,N_4159,N_4112);
or U4226 (N_4226,N_4037,N_4190);
and U4227 (N_4227,N_4018,N_4004);
nor U4228 (N_4228,N_4193,N_4171);
or U4229 (N_4229,N_4093,N_4091);
nand U4230 (N_4230,N_4046,N_4085);
or U4231 (N_4231,N_4067,N_4092);
xnor U4232 (N_4232,N_4141,N_4140);
nor U4233 (N_4233,N_4155,N_4084);
nor U4234 (N_4234,N_4023,N_4036);
or U4235 (N_4235,N_4119,N_4133);
nand U4236 (N_4236,N_4038,N_4104);
nand U4237 (N_4237,N_4098,N_4164);
and U4238 (N_4238,N_4025,N_4187);
nor U4239 (N_4239,N_4117,N_4158);
nand U4240 (N_4240,N_4041,N_4057);
and U4241 (N_4241,N_4105,N_4115);
or U4242 (N_4242,N_4130,N_4003);
nor U4243 (N_4243,N_4021,N_4162);
nor U4244 (N_4244,N_4148,N_4113);
and U4245 (N_4245,N_4011,N_4050);
xnor U4246 (N_4246,N_4014,N_4149);
nand U4247 (N_4247,N_4078,N_4139);
and U4248 (N_4248,N_4077,N_4012);
nand U4249 (N_4249,N_4182,N_4080);
nand U4250 (N_4250,N_4033,N_4005);
xor U4251 (N_4251,N_4065,N_4020);
or U4252 (N_4252,N_4052,N_4034);
nand U4253 (N_4253,N_4062,N_4063);
xnor U4254 (N_4254,N_4044,N_4160);
and U4255 (N_4255,N_4198,N_4194);
nand U4256 (N_4256,N_4032,N_4088);
or U4257 (N_4257,N_4097,N_4167);
and U4258 (N_4258,N_4015,N_4000);
and U4259 (N_4259,N_4040,N_4189);
or U4260 (N_4260,N_4053,N_4103);
nand U4261 (N_4261,N_4006,N_4042);
and U4262 (N_4262,N_4195,N_4175);
and U4263 (N_4263,N_4169,N_4031);
xor U4264 (N_4264,N_4166,N_4196);
or U4265 (N_4265,N_4045,N_4094);
xnor U4266 (N_4266,N_4026,N_4123);
or U4267 (N_4267,N_4152,N_4081);
or U4268 (N_4268,N_4174,N_4009);
nand U4269 (N_4269,N_4134,N_4049);
nor U4270 (N_4270,N_4017,N_4180);
or U4271 (N_4271,N_4146,N_4157);
nor U4272 (N_4272,N_4126,N_4122);
nand U4273 (N_4273,N_4022,N_4058);
xnor U4274 (N_4274,N_4142,N_4127);
and U4275 (N_4275,N_4001,N_4168);
or U4276 (N_4276,N_4073,N_4199);
nand U4277 (N_4277,N_4007,N_4181);
nor U4278 (N_4278,N_4064,N_4128);
or U4279 (N_4279,N_4086,N_4090);
or U4280 (N_4280,N_4054,N_4008);
nand U4281 (N_4281,N_4072,N_4153);
nand U4282 (N_4282,N_4096,N_4074);
or U4283 (N_4283,N_4083,N_4129);
nor U4284 (N_4284,N_4125,N_4137);
nand U4285 (N_4285,N_4027,N_4138);
nor U4286 (N_4286,N_4178,N_4135);
and U4287 (N_4287,N_4087,N_4002);
nor U4288 (N_4288,N_4029,N_4176);
or U4289 (N_4289,N_4147,N_4150);
and U4290 (N_4290,N_4059,N_4154);
xnor U4291 (N_4291,N_4071,N_4024);
xnor U4292 (N_4292,N_4019,N_4082);
or U4293 (N_4293,N_4120,N_4043);
xor U4294 (N_4294,N_4197,N_4016);
nor U4295 (N_4295,N_4108,N_4118);
nor U4296 (N_4296,N_4075,N_4110);
nand U4297 (N_4297,N_4177,N_4055);
xnor U4298 (N_4298,N_4114,N_4061);
xnor U4299 (N_4299,N_4039,N_4185);
xor U4300 (N_4300,N_4052,N_4191);
or U4301 (N_4301,N_4109,N_4049);
or U4302 (N_4302,N_4043,N_4170);
nand U4303 (N_4303,N_4063,N_4130);
or U4304 (N_4304,N_4054,N_4070);
xnor U4305 (N_4305,N_4060,N_4155);
nand U4306 (N_4306,N_4009,N_4124);
nor U4307 (N_4307,N_4042,N_4199);
nor U4308 (N_4308,N_4080,N_4001);
xor U4309 (N_4309,N_4057,N_4009);
xnor U4310 (N_4310,N_4075,N_4123);
nand U4311 (N_4311,N_4158,N_4044);
and U4312 (N_4312,N_4094,N_4006);
xor U4313 (N_4313,N_4115,N_4020);
and U4314 (N_4314,N_4116,N_4140);
nor U4315 (N_4315,N_4038,N_4056);
nor U4316 (N_4316,N_4019,N_4120);
xor U4317 (N_4317,N_4138,N_4012);
or U4318 (N_4318,N_4042,N_4174);
nand U4319 (N_4319,N_4021,N_4174);
xor U4320 (N_4320,N_4087,N_4101);
or U4321 (N_4321,N_4086,N_4093);
xnor U4322 (N_4322,N_4187,N_4199);
or U4323 (N_4323,N_4173,N_4119);
and U4324 (N_4324,N_4059,N_4029);
nor U4325 (N_4325,N_4098,N_4133);
nor U4326 (N_4326,N_4128,N_4193);
nand U4327 (N_4327,N_4061,N_4199);
and U4328 (N_4328,N_4064,N_4196);
xor U4329 (N_4329,N_4147,N_4071);
nor U4330 (N_4330,N_4129,N_4074);
nor U4331 (N_4331,N_4191,N_4066);
xnor U4332 (N_4332,N_4056,N_4130);
nor U4333 (N_4333,N_4190,N_4176);
and U4334 (N_4334,N_4041,N_4026);
nor U4335 (N_4335,N_4077,N_4088);
or U4336 (N_4336,N_4017,N_4004);
or U4337 (N_4337,N_4196,N_4105);
nor U4338 (N_4338,N_4135,N_4072);
nor U4339 (N_4339,N_4000,N_4063);
nor U4340 (N_4340,N_4197,N_4191);
or U4341 (N_4341,N_4043,N_4108);
or U4342 (N_4342,N_4169,N_4136);
nor U4343 (N_4343,N_4054,N_4017);
xor U4344 (N_4344,N_4010,N_4020);
or U4345 (N_4345,N_4010,N_4152);
nor U4346 (N_4346,N_4023,N_4109);
xor U4347 (N_4347,N_4134,N_4181);
xor U4348 (N_4348,N_4170,N_4069);
and U4349 (N_4349,N_4003,N_4018);
and U4350 (N_4350,N_4012,N_4126);
nor U4351 (N_4351,N_4055,N_4057);
nor U4352 (N_4352,N_4176,N_4089);
xor U4353 (N_4353,N_4139,N_4120);
nor U4354 (N_4354,N_4061,N_4155);
xnor U4355 (N_4355,N_4122,N_4190);
or U4356 (N_4356,N_4173,N_4040);
nand U4357 (N_4357,N_4112,N_4179);
xnor U4358 (N_4358,N_4088,N_4047);
and U4359 (N_4359,N_4138,N_4090);
or U4360 (N_4360,N_4020,N_4046);
xnor U4361 (N_4361,N_4042,N_4194);
xor U4362 (N_4362,N_4141,N_4184);
or U4363 (N_4363,N_4002,N_4129);
xor U4364 (N_4364,N_4148,N_4057);
and U4365 (N_4365,N_4118,N_4163);
nand U4366 (N_4366,N_4020,N_4087);
nor U4367 (N_4367,N_4093,N_4152);
xor U4368 (N_4368,N_4108,N_4197);
nand U4369 (N_4369,N_4156,N_4074);
nor U4370 (N_4370,N_4052,N_4068);
or U4371 (N_4371,N_4027,N_4187);
nor U4372 (N_4372,N_4070,N_4036);
xor U4373 (N_4373,N_4109,N_4123);
or U4374 (N_4374,N_4198,N_4108);
xor U4375 (N_4375,N_4066,N_4048);
nand U4376 (N_4376,N_4028,N_4175);
or U4377 (N_4377,N_4100,N_4199);
xnor U4378 (N_4378,N_4187,N_4101);
nor U4379 (N_4379,N_4001,N_4109);
or U4380 (N_4380,N_4125,N_4194);
nor U4381 (N_4381,N_4007,N_4187);
nor U4382 (N_4382,N_4051,N_4041);
and U4383 (N_4383,N_4093,N_4197);
and U4384 (N_4384,N_4090,N_4049);
xnor U4385 (N_4385,N_4049,N_4048);
or U4386 (N_4386,N_4160,N_4156);
and U4387 (N_4387,N_4143,N_4020);
nor U4388 (N_4388,N_4048,N_4095);
nand U4389 (N_4389,N_4002,N_4165);
nor U4390 (N_4390,N_4004,N_4005);
or U4391 (N_4391,N_4102,N_4020);
nand U4392 (N_4392,N_4178,N_4091);
and U4393 (N_4393,N_4095,N_4077);
and U4394 (N_4394,N_4084,N_4042);
or U4395 (N_4395,N_4044,N_4191);
and U4396 (N_4396,N_4076,N_4065);
and U4397 (N_4397,N_4023,N_4187);
xor U4398 (N_4398,N_4093,N_4004);
and U4399 (N_4399,N_4020,N_4180);
xnor U4400 (N_4400,N_4310,N_4272);
xor U4401 (N_4401,N_4372,N_4356);
and U4402 (N_4402,N_4298,N_4379);
nand U4403 (N_4403,N_4375,N_4271);
nor U4404 (N_4404,N_4318,N_4207);
or U4405 (N_4405,N_4225,N_4315);
nor U4406 (N_4406,N_4327,N_4282);
nor U4407 (N_4407,N_4306,N_4369);
xor U4408 (N_4408,N_4246,N_4389);
nor U4409 (N_4409,N_4312,N_4200);
xnor U4410 (N_4410,N_4233,N_4365);
or U4411 (N_4411,N_4337,N_4242);
and U4412 (N_4412,N_4270,N_4274);
or U4413 (N_4413,N_4206,N_4221);
nor U4414 (N_4414,N_4304,N_4319);
nor U4415 (N_4415,N_4366,N_4278);
nor U4416 (N_4416,N_4300,N_4215);
and U4417 (N_4417,N_4394,N_4224);
or U4418 (N_4418,N_4349,N_4360);
nor U4419 (N_4419,N_4383,N_4218);
or U4420 (N_4420,N_4330,N_4211);
nand U4421 (N_4421,N_4364,N_4236);
xor U4422 (N_4422,N_4230,N_4223);
nand U4423 (N_4423,N_4397,N_4249);
nand U4424 (N_4424,N_4244,N_4261);
xnor U4425 (N_4425,N_4228,N_4232);
and U4426 (N_4426,N_4205,N_4212);
nand U4427 (N_4427,N_4324,N_4339);
nor U4428 (N_4428,N_4226,N_4220);
nor U4429 (N_4429,N_4255,N_4276);
xor U4430 (N_4430,N_4243,N_4346);
or U4431 (N_4431,N_4374,N_4381);
xor U4432 (N_4432,N_4229,N_4257);
nand U4433 (N_4433,N_4378,N_4260);
xor U4434 (N_4434,N_4256,N_4214);
nand U4435 (N_4435,N_4347,N_4286);
xor U4436 (N_4436,N_4317,N_4362);
nand U4437 (N_4437,N_4336,N_4253);
nor U4438 (N_4438,N_4333,N_4338);
or U4439 (N_4439,N_4329,N_4250);
or U4440 (N_4440,N_4398,N_4380);
nand U4441 (N_4441,N_4263,N_4309);
nor U4442 (N_4442,N_4284,N_4393);
nand U4443 (N_4443,N_4252,N_4370);
nand U4444 (N_4444,N_4351,N_4291);
or U4445 (N_4445,N_4285,N_4363);
or U4446 (N_4446,N_4384,N_4386);
and U4447 (N_4447,N_4332,N_4245);
nand U4448 (N_4448,N_4316,N_4296);
nor U4449 (N_4449,N_4281,N_4340);
and U4450 (N_4450,N_4395,N_4288);
and U4451 (N_4451,N_4368,N_4361);
or U4452 (N_4452,N_4292,N_4358);
xor U4453 (N_4453,N_4202,N_4203);
or U4454 (N_4454,N_4267,N_4287);
xor U4455 (N_4455,N_4264,N_4385);
and U4456 (N_4456,N_4280,N_4305);
or U4457 (N_4457,N_4396,N_4247);
and U4458 (N_4458,N_4266,N_4313);
nand U4459 (N_4459,N_4290,N_4234);
and U4460 (N_4460,N_4320,N_4325);
nor U4461 (N_4461,N_4314,N_4399);
or U4462 (N_4462,N_4342,N_4219);
and U4463 (N_4463,N_4302,N_4345);
and U4464 (N_4464,N_4373,N_4299);
nand U4465 (N_4465,N_4268,N_4311);
nor U4466 (N_4466,N_4273,N_4210);
or U4467 (N_4467,N_4390,N_4307);
xnor U4468 (N_4468,N_4295,N_4275);
xnor U4469 (N_4469,N_4344,N_4334);
xnor U4470 (N_4470,N_4382,N_4297);
xor U4471 (N_4471,N_4239,N_4227);
nand U4472 (N_4472,N_4354,N_4277);
nand U4473 (N_4473,N_4248,N_4240);
nor U4474 (N_4474,N_4387,N_4237);
xnor U4475 (N_4475,N_4204,N_4231);
and U4476 (N_4476,N_4391,N_4303);
nand U4477 (N_4477,N_4376,N_4321);
xnor U4478 (N_4478,N_4359,N_4353);
nor U4479 (N_4479,N_4259,N_4367);
nor U4480 (N_4480,N_4283,N_4258);
xor U4481 (N_4481,N_4254,N_4357);
nor U4482 (N_4482,N_4350,N_4328);
xor U4483 (N_4483,N_4326,N_4377);
nand U4484 (N_4484,N_4269,N_4343);
xor U4485 (N_4485,N_4322,N_4348);
nand U4486 (N_4486,N_4235,N_4352);
and U4487 (N_4487,N_4341,N_4262);
nor U4488 (N_4488,N_4371,N_4301);
nand U4489 (N_4489,N_4289,N_4238);
nand U4490 (N_4490,N_4335,N_4388);
xor U4491 (N_4491,N_4294,N_4208);
nor U4492 (N_4492,N_4293,N_4217);
nand U4493 (N_4493,N_4209,N_4392);
nand U4494 (N_4494,N_4323,N_4308);
and U4495 (N_4495,N_4279,N_4201);
xor U4496 (N_4496,N_4213,N_4251);
xnor U4497 (N_4497,N_4222,N_4355);
xor U4498 (N_4498,N_4241,N_4265);
or U4499 (N_4499,N_4331,N_4216);
or U4500 (N_4500,N_4395,N_4289);
xor U4501 (N_4501,N_4264,N_4331);
and U4502 (N_4502,N_4382,N_4361);
xor U4503 (N_4503,N_4275,N_4243);
xnor U4504 (N_4504,N_4399,N_4274);
nand U4505 (N_4505,N_4341,N_4229);
nand U4506 (N_4506,N_4271,N_4361);
and U4507 (N_4507,N_4276,N_4220);
and U4508 (N_4508,N_4318,N_4213);
or U4509 (N_4509,N_4338,N_4367);
xnor U4510 (N_4510,N_4303,N_4234);
and U4511 (N_4511,N_4218,N_4275);
or U4512 (N_4512,N_4383,N_4242);
or U4513 (N_4513,N_4379,N_4382);
xor U4514 (N_4514,N_4247,N_4348);
or U4515 (N_4515,N_4238,N_4219);
nor U4516 (N_4516,N_4281,N_4275);
nand U4517 (N_4517,N_4275,N_4240);
and U4518 (N_4518,N_4381,N_4211);
nor U4519 (N_4519,N_4208,N_4392);
xnor U4520 (N_4520,N_4322,N_4203);
or U4521 (N_4521,N_4361,N_4373);
or U4522 (N_4522,N_4319,N_4268);
nand U4523 (N_4523,N_4243,N_4228);
xnor U4524 (N_4524,N_4278,N_4289);
and U4525 (N_4525,N_4350,N_4211);
nand U4526 (N_4526,N_4367,N_4322);
nor U4527 (N_4527,N_4383,N_4361);
xnor U4528 (N_4528,N_4256,N_4210);
and U4529 (N_4529,N_4280,N_4292);
nor U4530 (N_4530,N_4265,N_4395);
or U4531 (N_4531,N_4282,N_4203);
nand U4532 (N_4532,N_4343,N_4294);
nor U4533 (N_4533,N_4373,N_4242);
or U4534 (N_4534,N_4321,N_4312);
nor U4535 (N_4535,N_4382,N_4233);
or U4536 (N_4536,N_4316,N_4380);
nand U4537 (N_4537,N_4293,N_4351);
and U4538 (N_4538,N_4324,N_4332);
nor U4539 (N_4539,N_4310,N_4355);
nor U4540 (N_4540,N_4222,N_4336);
nand U4541 (N_4541,N_4247,N_4288);
nand U4542 (N_4542,N_4366,N_4215);
xor U4543 (N_4543,N_4337,N_4355);
nand U4544 (N_4544,N_4217,N_4247);
xor U4545 (N_4545,N_4218,N_4235);
and U4546 (N_4546,N_4307,N_4372);
xnor U4547 (N_4547,N_4360,N_4202);
and U4548 (N_4548,N_4395,N_4316);
xnor U4549 (N_4549,N_4319,N_4353);
and U4550 (N_4550,N_4247,N_4284);
or U4551 (N_4551,N_4272,N_4362);
nand U4552 (N_4552,N_4358,N_4263);
xor U4553 (N_4553,N_4312,N_4238);
and U4554 (N_4554,N_4396,N_4289);
nor U4555 (N_4555,N_4377,N_4347);
or U4556 (N_4556,N_4302,N_4277);
nand U4557 (N_4557,N_4237,N_4222);
and U4558 (N_4558,N_4343,N_4256);
nor U4559 (N_4559,N_4329,N_4276);
nand U4560 (N_4560,N_4253,N_4307);
nand U4561 (N_4561,N_4200,N_4257);
or U4562 (N_4562,N_4316,N_4394);
nand U4563 (N_4563,N_4322,N_4337);
xor U4564 (N_4564,N_4343,N_4360);
and U4565 (N_4565,N_4366,N_4275);
nor U4566 (N_4566,N_4363,N_4304);
or U4567 (N_4567,N_4244,N_4365);
nor U4568 (N_4568,N_4302,N_4294);
and U4569 (N_4569,N_4243,N_4237);
nor U4570 (N_4570,N_4220,N_4384);
or U4571 (N_4571,N_4269,N_4389);
and U4572 (N_4572,N_4262,N_4293);
or U4573 (N_4573,N_4294,N_4289);
nand U4574 (N_4574,N_4343,N_4295);
nor U4575 (N_4575,N_4338,N_4324);
xnor U4576 (N_4576,N_4297,N_4255);
or U4577 (N_4577,N_4398,N_4230);
and U4578 (N_4578,N_4376,N_4255);
and U4579 (N_4579,N_4347,N_4202);
or U4580 (N_4580,N_4295,N_4290);
nor U4581 (N_4581,N_4372,N_4256);
and U4582 (N_4582,N_4225,N_4397);
nand U4583 (N_4583,N_4386,N_4200);
xnor U4584 (N_4584,N_4252,N_4294);
xnor U4585 (N_4585,N_4290,N_4246);
nor U4586 (N_4586,N_4348,N_4277);
and U4587 (N_4587,N_4396,N_4293);
xor U4588 (N_4588,N_4215,N_4393);
xor U4589 (N_4589,N_4286,N_4302);
xor U4590 (N_4590,N_4298,N_4386);
or U4591 (N_4591,N_4304,N_4331);
nand U4592 (N_4592,N_4358,N_4377);
nor U4593 (N_4593,N_4225,N_4255);
xor U4594 (N_4594,N_4249,N_4291);
or U4595 (N_4595,N_4332,N_4381);
and U4596 (N_4596,N_4350,N_4391);
and U4597 (N_4597,N_4288,N_4353);
and U4598 (N_4598,N_4282,N_4224);
nand U4599 (N_4599,N_4258,N_4271);
or U4600 (N_4600,N_4460,N_4546);
and U4601 (N_4601,N_4569,N_4597);
nand U4602 (N_4602,N_4455,N_4561);
nor U4603 (N_4603,N_4403,N_4563);
nand U4604 (N_4604,N_4473,N_4431);
nand U4605 (N_4605,N_4535,N_4556);
or U4606 (N_4606,N_4517,N_4558);
or U4607 (N_4607,N_4492,N_4594);
xnor U4608 (N_4608,N_4401,N_4576);
xor U4609 (N_4609,N_4598,N_4539);
nor U4610 (N_4610,N_4588,N_4466);
or U4611 (N_4611,N_4452,N_4545);
xor U4612 (N_4612,N_4554,N_4549);
or U4613 (N_4613,N_4409,N_4418);
xor U4614 (N_4614,N_4481,N_4439);
xor U4615 (N_4615,N_4447,N_4463);
nor U4616 (N_4616,N_4415,N_4562);
or U4617 (N_4617,N_4474,N_4578);
nand U4618 (N_4618,N_4440,N_4541);
xnor U4619 (N_4619,N_4408,N_4570);
nand U4620 (N_4620,N_4519,N_4437);
xor U4621 (N_4621,N_4567,N_4504);
and U4622 (N_4622,N_4582,N_4461);
nand U4623 (N_4623,N_4585,N_4464);
nor U4624 (N_4624,N_4498,N_4433);
and U4625 (N_4625,N_4574,N_4420);
nand U4626 (N_4626,N_4407,N_4599);
nand U4627 (N_4627,N_4497,N_4413);
nand U4628 (N_4628,N_4500,N_4448);
xor U4629 (N_4629,N_4451,N_4553);
or U4630 (N_4630,N_4518,N_4577);
nand U4631 (N_4631,N_4469,N_4538);
or U4632 (N_4632,N_4506,N_4482);
and U4633 (N_4633,N_4446,N_4485);
and U4634 (N_4634,N_4540,N_4527);
and U4635 (N_4635,N_4572,N_4470);
and U4636 (N_4636,N_4445,N_4551);
nor U4637 (N_4637,N_4471,N_4559);
xor U4638 (N_4638,N_4525,N_4425);
xor U4639 (N_4639,N_4421,N_4457);
and U4640 (N_4640,N_4489,N_4596);
or U4641 (N_4641,N_4580,N_4534);
and U4642 (N_4642,N_4552,N_4502);
nand U4643 (N_4643,N_4548,N_4565);
xor U4644 (N_4644,N_4479,N_4417);
xnor U4645 (N_4645,N_4579,N_4442);
nor U4646 (N_4646,N_4483,N_4543);
or U4647 (N_4647,N_4514,N_4512);
nand U4648 (N_4648,N_4501,N_4505);
xor U4649 (N_4649,N_4449,N_4520);
nand U4650 (N_4650,N_4402,N_4476);
and U4651 (N_4651,N_4499,N_4532);
nor U4652 (N_4652,N_4443,N_4522);
nand U4653 (N_4653,N_4586,N_4595);
xnor U4654 (N_4654,N_4516,N_4468);
nor U4655 (N_4655,N_4557,N_4591);
or U4656 (N_4656,N_4515,N_4491);
or U4657 (N_4657,N_4494,N_4587);
nand U4658 (N_4658,N_4475,N_4495);
and U4659 (N_4659,N_4426,N_4486);
or U4660 (N_4660,N_4513,N_4584);
nand U4661 (N_4661,N_4509,N_4480);
nor U4662 (N_4662,N_4568,N_4530);
xor U4663 (N_4663,N_4478,N_4493);
nand U4664 (N_4664,N_4444,N_4547);
xor U4665 (N_4665,N_4537,N_4529);
and U4666 (N_4666,N_4593,N_4412);
nor U4667 (N_4667,N_4472,N_4428);
nor U4668 (N_4668,N_4508,N_4467);
and U4669 (N_4669,N_4410,N_4462);
nand U4670 (N_4670,N_4555,N_4432);
nor U4671 (N_4671,N_4458,N_4414);
xor U4672 (N_4672,N_4422,N_4583);
nor U4673 (N_4673,N_4424,N_4400);
nand U4674 (N_4674,N_4484,N_4465);
nand U4675 (N_4675,N_4573,N_4434);
and U4676 (N_4676,N_4416,N_4427);
xnor U4677 (N_4677,N_4450,N_4487);
nor U4678 (N_4678,N_4566,N_4454);
xnor U4679 (N_4679,N_4477,N_4571);
nor U4680 (N_4680,N_4503,N_4581);
nand U4681 (N_4681,N_4523,N_4592);
or U4682 (N_4682,N_4542,N_4423);
nand U4683 (N_4683,N_4575,N_4430);
xnor U4684 (N_4684,N_4550,N_4405);
and U4685 (N_4685,N_4590,N_4438);
nand U4686 (N_4686,N_4536,N_4526);
xnor U4687 (N_4687,N_4453,N_4411);
xnor U4688 (N_4688,N_4436,N_4528);
or U4689 (N_4689,N_4406,N_4435);
xor U4690 (N_4690,N_4496,N_4589);
nor U4691 (N_4691,N_4490,N_4524);
xnor U4692 (N_4692,N_4521,N_4511);
xor U4693 (N_4693,N_4533,N_4456);
or U4694 (N_4694,N_4560,N_4510);
and U4695 (N_4695,N_4507,N_4441);
nor U4696 (N_4696,N_4564,N_4429);
xor U4697 (N_4697,N_4459,N_4544);
and U4698 (N_4698,N_4404,N_4531);
xnor U4699 (N_4699,N_4488,N_4419);
nand U4700 (N_4700,N_4402,N_4454);
xor U4701 (N_4701,N_4481,N_4591);
and U4702 (N_4702,N_4408,N_4459);
nor U4703 (N_4703,N_4593,N_4503);
xor U4704 (N_4704,N_4558,N_4521);
and U4705 (N_4705,N_4493,N_4479);
nand U4706 (N_4706,N_4549,N_4578);
nor U4707 (N_4707,N_4584,N_4594);
or U4708 (N_4708,N_4457,N_4405);
or U4709 (N_4709,N_4577,N_4537);
nor U4710 (N_4710,N_4594,N_4590);
nand U4711 (N_4711,N_4561,N_4548);
nor U4712 (N_4712,N_4516,N_4579);
nand U4713 (N_4713,N_4511,N_4464);
nor U4714 (N_4714,N_4529,N_4469);
nand U4715 (N_4715,N_4507,N_4573);
xnor U4716 (N_4716,N_4453,N_4501);
xnor U4717 (N_4717,N_4527,N_4457);
nor U4718 (N_4718,N_4493,N_4465);
nand U4719 (N_4719,N_4487,N_4416);
xnor U4720 (N_4720,N_4460,N_4456);
xor U4721 (N_4721,N_4416,N_4534);
nor U4722 (N_4722,N_4494,N_4569);
and U4723 (N_4723,N_4516,N_4493);
nor U4724 (N_4724,N_4482,N_4438);
and U4725 (N_4725,N_4407,N_4403);
nor U4726 (N_4726,N_4554,N_4498);
xnor U4727 (N_4727,N_4431,N_4576);
and U4728 (N_4728,N_4558,N_4483);
nand U4729 (N_4729,N_4459,N_4415);
or U4730 (N_4730,N_4564,N_4596);
nand U4731 (N_4731,N_4483,N_4449);
or U4732 (N_4732,N_4492,N_4431);
or U4733 (N_4733,N_4564,N_4414);
and U4734 (N_4734,N_4585,N_4417);
nor U4735 (N_4735,N_4585,N_4578);
nor U4736 (N_4736,N_4567,N_4460);
or U4737 (N_4737,N_4491,N_4585);
xor U4738 (N_4738,N_4522,N_4470);
and U4739 (N_4739,N_4484,N_4565);
nor U4740 (N_4740,N_4520,N_4535);
xnor U4741 (N_4741,N_4540,N_4569);
and U4742 (N_4742,N_4503,N_4552);
and U4743 (N_4743,N_4491,N_4510);
or U4744 (N_4744,N_4439,N_4445);
nand U4745 (N_4745,N_4599,N_4553);
nand U4746 (N_4746,N_4433,N_4520);
nor U4747 (N_4747,N_4494,N_4506);
or U4748 (N_4748,N_4484,N_4499);
nor U4749 (N_4749,N_4456,N_4595);
or U4750 (N_4750,N_4553,N_4598);
and U4751 (N_4751,N_4532,N_4546);
nand U4752 (N_4752,N_4481,N_4538);
xnor U4753 (N_4753,N_4477,N_4577);
or U4754 (N_4754,N_4504,N_4404);
xor U4755 (N_4755,N_4542,N_4433);
nand U4756 (N_4756,N_4466,N_4457);
and U4757 (N_4757,N_4483,N_4451);
or U4758 (N_4758,N_4507,N_4439);
nand U4759 (N_4759,N_4460,N_4411);
xor U4760 (N_4760,N_4565,N_4438);
xnor U4761 (N_4761,N_4531,N_4516);
nor U4762 (N_4762,N_4525,N_4567);
nand U4763 (N_4763,N_4578,N_4406);
xor U4764 (N_4764,N_4559,N_4482);
nand U4765 (N_4765,N_4505,N_4455);
xor U4766 (N_4766,N_4537,N_4570);
nand U4767 (N_4767,N_4525,N_4486);
nand U4768 (N_4768,N_4583,N_4494);
or U4769 (N_4769,N_4590,N_4597);
nor U4770 (N_4770,N_4568,N_4493);
and U4771 (N_4771,N_4560,N_4548);
xor U4772 (N_4772,N_4415,N_4467);
nand U4773 (N_4773,N_4589,N_4463);
xor U4774 (N_4774,N_4515,N_4484);
xor U4775 (N_4775,N_4548,N_4502);
xor U4776 (N_4776,N_4442,N_4535);
xor U4777 (N_4777,N_4485,N_4426);
nand U4778 (N_4778,N_4569,N_4584);
nor U4779 (N_4779,N_4500,N_4478);
nor U4780 (N_4780,N_4418,N_4508);
nor U4781 (N_4781,N_4468,N_4537);
xnor U4782 (N_4782,N_4423,N_4526);
xnor U4783 (N_4783,N_4496,N_4508);
xnor U4784 (N_4784,N_4560,N_4432);
or U4785 (N_4785,N_4507,N_4590);
xor U4786 (N_4786,N_4516,N_4577);
nand U4787 (N_4787,N_4481,N_4529);
nor U4788 (N_4788,N_4455,N_4494);
xnor U4789 (N_4789,N_4503,N_4473);
xor U4790 (N_4790,N_4421,N_4551);
or U4791 (N_4791,N_4577,N_4487);
nand U4792 (N_4792,N_4412,N_4434);
nor U4793 (N_4793,N_4505,N_4422);
or U4794 (N_4794,N_4599,N_4572);
xnor U4795 (N_4795,N_4420,N_4540);
nand U4796 (N_4796,N_4585,N_4423);
xor U4797 (N_4797,N_4569,N_4513);
or U4798 (N_4798,N_4520,N_4461);
xnor U4799 (N_4799,N_4573,N_4460);
nand U4800 (N_4800,N_4637,N_4686);
xnor U4801 (N_4801,N_4702,N_4701);
nand U4802 (N_4802,N_4730,N_4692);
and U4803 (N_4803,N_4768,N_4688);
nand U4804 (N_4804,N_4611,N_4790);
or U4805 (N_4805,N_4799,N_4678);
and U4806 (N_4806,N_4605,N_4650);
nor U4807 (N_4807,N_4662,N_4759);
or U4808 (N_4808,N_4608,N_4663);
or U4809 (N_4809,N_4647,N_4723);
or U4810 (N_4810,N_4665,N_4752);
or U4811 (N_4811,N_4739,N_4771);
or U4812 (N_4812,N_4689,N_4656);
xor U4813 (N_4813,N_4666,N_4726);
nand U4814 (N_4814,N_4753,N_4755);
xnor U4815 (N_4815,N_4792,N_4785);
nand U4816 (N_4816,N_4738,N_4777);
and U4817 (N_4817,N_4672,N_4798);
nand U4818 (N_4818,N_4668,N_4643);
nor U4819 (N_4819,N_4646,N_4619);
nor U4820 (N_4820,N_4722,N_4659);
or U4821 (N_4821,N_4747,N_4660);
xnor U4822 (N_4822,N_4710,N_4763);
nand U4823 (N_4823,N_4622,N_4602);
nand U4824 (N_4824,N_4626,N_4742);
or U4825 (N_4825,N_4717,N_4741);
and U4826 (N_4826,N_4667,N_4708);
and U4827 (N_4827,N_4709,N_4704);
and U4828 (N_4828,N_4703,N_4766);
and U4829 (N_4829,N_4729,N_4633);
xnor U4830 (N_4830,N_4700,N_4671);
and U4831 (N_4831,N_4630,N_4731);
xnor U4832 (N_4832,N_4705,N_4744);
nor U4833 (N_4833,N_4774,N_4749);
nor U4834 (N_4834,N_4684,N_4603);
xor U4835 (N_4835,N_4788,N_4736);
xor U4836 (N_4836,N_4694,N_4740);
or U4837 (N_4837,N_4748,N_4649);
nand U4838 (N_4838,N_4779,N_4743);
nand U4839 (N_4839,N_4795,N_4712);
and U4840 (N_4840,N_4679,N_4655);
nand U4841 (N_4841,N_4651,N_4609);
nand U4842 (N_4842,N_4685,N_4797);
xor U4843 (N_4843,N_4786,N_4783);
xor U4844 (N_4844,N_4762,N_4617);
nand U4845 (N_4845,N_4628,N_4727);
xnor U4846 (N_4846,N_4769,N_4773);
xnor U4847 (N_4847,N_4789,N_4653);
or U4848 (N_4848,N_4697,N_4606);
or U4849 (N_4849,N_4765,N_4756);
or U4850 (N_4850,N_4751,N_4796);
or U4851 (N_4851,N_4680,N_4782);
and U4852 (N_4852,N_4794,N_4623);
and U4853 (N_4853,N_4616,N_4724);
and U4854 (N_4854,N_4698,N_4600);
nand U4855 (N_4855,N_4683,N_4677);
xnor U4856 (N_4856,N_4776,N_4640);
or U4857 (N_4857,N_4604,N_4601);
xor U4858 (N_4858,N_4661,N_4781);
nor U4859 (N_4859,N_4775,N_4618);
nor U4860 (N_4860,N_4784,N_4607);
and U4861 (N_4861,N_4673,N_4787);
nand U4862 (N_4862,N_4714,N_4636);
xnor U4863 (N_4863,N_4715,N_4706);
and U4864 (N_4864,N_4691,N_4631);
nor U4865 (N_4865,N_4681,N_4718);
xor U4866 (N_4866,N_4629,N_4674);
and U4867 (N_4867,N_4757,N_4652);
nand U4868 (N_4868,N_4638,N_4657);
xnor U4869 (N_4869,N_4615,N_4733);
nor U4870 (N_4870,N_4620,N_4645);
or U4871 (N_4871,N_4707,N_4670);
nand U4872 (N_4872,N_4719,N_4693);
nand U4873 (N_4873,N_4634,N_4641);
nand U4874 (N_4874,N_4760,N_4627);
nor U4875 (N_4875,N_4713,N_4612);
nor U4876 (N_4876,N_4761,N_4772);
and U4877 (N_4877,N_4676,N_4732);
nor U4878 (N_4878,N_4754,N_4621);
nand U4879 (N_4879,N_4664,N_4658);
nor U4880 (N_4880,N_4734,N_4745);
xor U4881 (N_4881,N_4711,N_4764);
and U4882 (N_4882,N_4725,N_4654);
or U4883 (N_4883,N_4635,N_4675);
nor U4884 (N_4884,N_4610,N_4791);
and U4885 (N_4885,N_4778,N_4687);
or U4886 (N_4886,N_4728,N_4699);
nand U4887 (N_4887,N_4669,N_4746);
xnor U4888 (N_4888,N_4624,N_4735);
xnor U4889 (N_4889,N_4767,N_4682);
xor U4890 (N_4890,N_4716,N_4690);
nand U4891 (N_4891,N_4613,N_4614);
and U4892 (N_4892,N_4770,N_4758);
nand U4893 (N_4893,N_4780,N_4737);
or U4894 (N_4894,N_4720,N_4695);
or U4895 (N_4895,N_4632,N_4625);
xnor U4896 (N_4896,N_4721,N_4639);
or U4897 (N_4897,N_4648,N_4793);
or U4898 (N_4898,N_4644,N_4750);
and U4899 (N_4899,N_4642,N_4696);
or U4900 (N_4900,N_4629,N_4648);
and U4901 (N_4901,N_4727,N_4751);
nor U4902 (N_4902,N_4735,N_4728);
nand U4903 (N_4903,N_4701,N_4761);
or U4904 (N_4904,N_4629,N_4657);
and U4905 (N_4905,N_4735,N_4769);
nor U4906 (N_4906,N_4683,N_4796);
and U4907 (N_4907,N_4757,N_4751);
and U4908 (N_4908,N_4605,N_4665);
or U4909 (N_4909,N_4607,N_4698);
or U4910 (N_4910,N_4672,N_4754);
xnor U4911 (N_4911,N_4608,N_4781);
and U4912 (N_4912,N_4773,N_4602);
nor U4913 (N_4913,N_4772,N_4780);
xnor U4914 (N_4914,N_4667,N_4775);
xnor U4915 (N_4915,N_4774,N_4753);
nand U4916 (N_4916,N_4619,N_4715);
nand U4917 (N_4917,N_4672,N_4729);
nor U4918 (N_4918,N_4634,N_4685);
and U4919 (N_4919,N_4791,N_4671);
xor U4920 (N_4920,N_4727,N_4622);
nand U4921 (N_4921,N_4762,N_4612);
or U4922 (N_4922,N_4615,N_4713);
nor U4923 (N_4923,N_4724,N_4749);
xor U4924 (N_4924,N_4604,N_4652);
nand U4925 (N_4925,N_4736,N_4785);
xor U4926 (N_4926,N_4662,N_4797);
nand U4927 (N_4927,N_4719,N_4779);
nand U4928 (N_4928,N_4629,N_4792);
xor U4929 (N_4929,N_4639,N_4710);
xnor U4930 (N_4930,N_4626,N_4736);
or U4931 (N_4931,N_4619,N_4747);
or U4932 (N_4932,N_4665,N_4742);
or U4933 (N_4933,N_4743,N_4782);
and U4934 (N_4934,N_4639,N_4793);
xnor U4935 (N_4935,N_4614,N_4746);
nand U4936 (N_4936,N_4672,N_4715);
or U4937 (N_4937,N_4734,N_4794);
nor U4938 (N_4938,N_4688,N_4712);
nor U4939 (N_4939,N_4751,N_4724);
or U4940 (N_4940,N_4744,N_4631);
nor U4941 (N_4941,N_4719,N_4708);
xor U4942 (N_4942,N_4772,N_4654);
and U4943 (N_4943,N_4706,N_4746);
nor U4944 (N_4944,N_4645,N_4778);
or U4945 (N_4945,N_4763,N_4722);
nor U4946 (N_4946,N_4684,N_4655);
and U4947 (N_4947,N_4673,N_4661);
and U4948 (N_4948,N_4601,N_4760);
or U4949 (N_4949,N_4736,N_4731);
xor U4950 (N_4950,N_4689,N_4605);
and U4951 (N_4951,N_4708,N_4745);
and U4952 (N_4952,N_4653,N_4717);
nor U4953 (N_4953,N_4667,N_4668);
nand U4954 (N_4954,N_4624,N_4614);
nand U4955 (N_4955,N_4710,N_4684);
nor U4956 (N_4956,N_4727,N_4790);
xor U4957 (N_4957,N_4717,N_4633);
nor U4958 (N_4958,N_4642,N_4607);
and U4959 (N_4959,N_4635,N_4763);
nor U4960 (N_4960,N_4773,N_4709);
nand U4961 (N_4961,N_4672,N_4668);
or U4962 (N_4962,N_4739,N_4795);
xor U4963 (N_4963,N_4688,N_4764);
nand U4964 (N_4964,N_4632,N_4697);
nor U4965 (N_4965,N_4763,N_4717);
nand U4966 (N_4966,N_4614,N_4652);
xnor U4967 (N_4967,N_4666,N_4719);
and U4968 (N_4968,N_4668,N_4790);
nand U4969 (N_4969,N_4762,N_4784);
or U4970 (N_4970,N_4607,N_4794);
nand U4971 (N_4971,N_4656,N_4766);
and U4972 (N_4972,N_4663,N_4669);
nor U4973 (N_4973,N_4741,N_4634);
xnor U4974 (N_4974,N_4739,N_4774);
xor U4975 (N_4975,N_4608,N_4667);
nand U4976 (N_4976,N_4612,N_4674);
and U4977 (N_4977,N_4762,N_4724);
and U4978 (N_4978,N_4778,N_4697);
xor U4979 (N_4979,N_4676,N_4674);
xor U4980 (N_4980,N_4737,N_4636);
and U4981 (N_4981,N_4649,N_4629);
xnor U4982 (N_4982,N_4751,N_4686);
or U4983 (N_4983,N_4711,N_4644);
or U4984 (N_4984,N_4651,N_4600);
nor U4985 (N_4985,N_4609,N_4720);
xor U4986 (N_4986,N_4763,N_4737);
and U4987 (N_4987,N_4722,N_4792);
nor U4988 (N_4988,N_4752,N_4799);
and U4989 (N_4989,N_4665,N_4679);
or U4990 (N_4990,N_4700,N_4614);
or U4991 (N_4991,N_4649,N_4689);
nor U4992 (N_4992,N_4612,N_4640);
xor U4993 (N_4993,N_4745,N_4668);
nor U4994 (N_4994,N_4722,N_4603);
and U4995 (N_4995,N_4765,N_4697);
and U4996 (N_4996,N_4644,N_4759);
and U4997 (N_4997,N_4671,N_4774);
nand U4998 (N_4998,N_4637,N_4685);
xnor U4999 (N_4999,N_4750,N_4770);
nand UO_0 (O_0,N_4850,N_4958);
xor UO_1 (O_1,N_4874,N_4954);
or UO_2 (O_2,N_4839,N_4911);
and UO_3 (O_3,N_4878,N_4826);
nor UO_4 (O_4,N_4897,N_4886);
and UO_5 (O_5,N_4900,N_4905);
nor UO_6 (O_6,N_4936,N_4914);
xor UO_7 (O_7,N_4857,N_4965);
xnor UO_8 (O_8,N_4992,N_4985);
and UO_9 (O_9,N_4805,N_4903);
nor UO_10 (O_10,N_4823,N_4801);
nand UO_11 (O_11,N_4959,N_4972);
xor UO_12 (O_12,N_4849,N_4929);
nand UO_13 (O_13,N_4993,N_4918);
xor UO_14 (O_14,N_4916,N_4837);
and UO_15 (O_15,N_4810,N_4835);
and UO_16 (O_16,N_4994,N_4830);
nor UO_17 (O_17,N_4833,N_4844);
or UO_18 (O_18,N_4983,N_4875);
and UO_19 (O_19,N_4933,N_4901);
nand UO_20 (O_20,N_4802,N_4871);
nand UO_21 (O_21,N_4962,N_4975);
or UO_22 (O_22,N_4980,N_4991);
and UO_23 (O_23,N_4892,N_4872);
nand UO_24 (O_24,N_4814,N_4937);
and UO_25 (O_25,N_4820,N_4949);
nand UO_26 (O_26,N_4856,N_4968);
and UO_27 (O_27,N_4957,N_4928);
nand UO_28 (O_28,N_4907,N_4974);
nor UO_29 (O_29,N_4909,N_4910);
xnor UO_30 (O_30,N_4862,N_4990);
or UO_31 (O_31,N_4843,N_4899);
or UO_32 (O_32,N_4915,N_4881);
nor UO_33 (O_33,N_4888,N_4829);
or UO_34 (O_34,N_4824,N_4950);
or UO_35 (O_35,N_4867,N_4969);
nand UO_36 (O_36,N_4931,N_4825);
xor UO_37 (O_37,N_4893,N_4869);
nor UO_38 (O_38,N_4848,N_4828);
xor UO_39 (O_39,N_4940,N_4836);
nor UO_40 (O_40,N_4923,N_4986);
nor UO_41 (O_41,N_4966,N_4847);
nand UO_42 (O_42,N_4941,N_4832);
and UO_43 (O_43,N_4819,N_4976);
xor UO_44 (O_44,N_4834,N_4948);
nor UO_45 (O_45,N_4908,N_4803);
and UO_46 (O_46,N_4852,N_4863);
nand UO_47 (O_47,N_4859,N_4996);
and UO_48 (O_48,N_4998,N_4880);
or UO_49 (O_49,N_4815,N_4841);
xnor UO_50 (O_50,N_4804,N_4979);
or UO_51 (O_51,N_4939,N_4812);
and UO_52 (O_52,N_4807,N_4861);
nand UO_53 (O_53,N_4842,N_4906);
xnor UO_54 (O_54,N_4868,N_4919);
xnor UO_55 (O_55,N_4921,N_4953);
xnor UO_56 (O_56,N_4951,N_4989);
or UO_57 (O_57,N_4858,N_4838);
nand UO_58 (O_58,N_4973,N_4865);
nand UO_59 (O_59,N_4866,N_4938);
xor UO_60 (O_60,N_4811,N_4821);
or UO_61 (O_61,N_4891,N_4942);
xor UO_62 (O_62,N_4944,N_4932);
and UO_63 (O_63,N_4877,N_4890);
or UO_64 (O_64,N_4920,N_4925);
nor UO_65 (O_65,N_4884,N_4896);
or UO_66 (O_66,N_4873,N_4943);
nor UO_67 (O_67,N_4851,N_4902);
nand UO_68 (O_68,N_4883,N_4935);
nand UO_69 (O_69,N_4971,N_4882);
xor UO_70 (O_70,N_4984,N_4822);
and UO_71 (O_71,N_4978,N_4870);
nor UO_72 (O_72,N_4917,N_4970);
xor UO_73 (O_73,N_4955,N_4952);
xnor UO_74 (O_74,N_4816,N_4831);
nor UO_75 (O_75,N_4895,N_4961);
nor UO_76 (O_76,N_4960,N_4889);
nor UO_77 (O_77,N_4876,N_4904);
nor UO_78 (O_78,N_4840,N_4945);
nor UO_79 (O_79,N_4845,N_4887);
and UO_80 (O_80,N_4864,N_4995);
or UO_81 (O_81,N_4926,N_4846);
xnor UO_82 (O_82,N_4981,N_4809);
or UO_83 (O_83,N_4808,N_4860);
or UO_84 (O_84,N_4817,N_4997);
and UO_85 (O_85,N_4947,N_4854);
and UO_86 (O_86,N_4924,N_4894);
nor UO_87 (O_87,N_4913,N_4963);
xor UO_88 (O_88,N_4946,N_4956);
or UO_89 (O_89,N_4898,N_4927);
and UO_90 (O_90,N_4806,N_4922);
and UO_91 (O_91,N_4977,N_4930);
and UO_92 (O_92,N_4934,N_4885);
or UO_93 (O_93,N_4818,N_4813);
and UO_94 (O_94,N_4879,N_4853);
or UO_95 (O_95,N_4967,N_4999);
nand UO_96 (O_96,N_4988,N_4855);
or UO_97 (O_97,N_4800,N_4912);
or UO_98 (O_98,N_4982,N_4827);
and UO_99 (O_99,N_4964,N_4987);
and UO_100 (O_100,N_4804,N_4832);
xnor UO_101 (O_101,N_4842,N_4984);
and UO_102 (O_102,N_4996,N_4927);
or UO_103 (O_103,N_4891,N_4958);
and UO_104 (O_104,N_4854,N_4804);
nor UO_105 (O_105,N_4857,N_4801);
nor UO_106 (O_106,N_4818,N_4973);
and UO_107 (O_107,N_4898,N_4811);
and UO_108 (O_108,N_4827,N_4876);
xnor UO_109 (O_109,N_4928,N_4898);
and UO_110 (O_110,N_4877,N_4948);
and UO_111 (O_111,N_4918,N_4900);
and UO_112 (O_112,N_4816,N_4870);
xnor UO_113 (O_113,N_4845,N_4815);
xnor UO_114 (O_114,N_4958,N_4990);
nand UO_115 (O_115,N_4947,N_4920);
nor UO_116 (O_116,N_4933,N_4840);
xor UO_117 (O_117,N_4854,N_4894);
and UO_118 (O_118,N_4871,N_4839);
nor UO_119 (O_119,N_4995,N_4945);
nand UO_120 (O_120,N_4861,N_4854);
nor UO_121 (O_121,N_4874,N_4939);
nand UO_122 (O_122,N_4889,N_4817);
and UO_123 (O_123,N_4914,N_4868);
and UO_124 (O_124,N_4800,N_4933);
xor UO_125 (O_125,N_4995,N_4854);
or UO_126 (O_126,N_4849,N_4980);
nand UO_127 (O_127,N_4925,N_4873);
or UO_128 (O_128,N_4973,N_4925);
or UO_129 (O_129,N_4929,N_4857);
xnor UO_130 (O_130,N_4903,N_4978);
nand UO_131 (O_131,N_4948,N_4981);
xnor UO_132 (O_132,N_4935,N_4989);
nand UO_133 (O_133,N_4926,N_4806);
xnor UO_134 (O_134,N_4880,N_4913);
or UO_135 (O_135,N_4908,N_4852);
and UO_136 (O_136,N_4967,N_4889);
or UO_137 (O_137,N_4909,N_4857);
xnor UO_138 (O_138,N_4858,N_4941);
and UO_139 (O_139,N_4905,N_4988);
nand UO_140 (O_140,N_4863,N_4996);
or UO_141 (O_141,N_4899,N_4973);
nand UO_142 (O_142,N_4915,N_4874);
xor UO_143 (O_143,N_4947,N_4942);
xor UO_144 (O_144,N_4968,N_4886);
nand UO_145 (O_145,N_4826,N_4871);
xnor UO_146 (O_146,N_4910,N_4836);
xnor UO_147 (O_147,N_4887,N_4801);
nand UO_148 (O_148,N_4829,N_4929);
and UO_149 (O_149,N_4943,N_4956);
nand UO_150 (O_150,N_4899,N_4867);
or UO_151 (O_151,N_4838,N_4997);
and UO_152 (O_152,N_4859,N_4867);
or UO_153 (O_153,N_4910,N_4892);
nand UO_154 (O_154,N_4994,N_4800);
xor UO_155 (O_155,N_4992,N_4940);
or UO_156 (O_156,N_4973,N_4869);
nand UO_157 (O_157,N_4812,N_4966);
and UO_158 (O_158,N_4877,N_4807);
xor UO_159 (O_159,N_4846,N_4822);
or UO_160 (O_160,N_4857,N_4999);
or UO_161 (O_161,N_4852,N_4932);
or UO_162 (O_162,N_4942,N_4834);
or UO_163 (O_163,N_4813,N_4906);
xnor UO_164 (O_164,N_4942,N_4949);
nand UO_165 (O_165,N_4996,N_4860);
xor UO_166 (O_166,N_4938,N_4968);
nor UO_167 (O_167,N_4924,N_4847);
xnor UO_168 (O_168,N_4864,N_4857);
or UO_169 (O_169,N_4801,N_4816);
nor UO_170 (O_170,N_4907,N_4815);
nor UO_171 (O_171,N_4888,N_4841);
nand UO_172 (O_172,N_4808,N_4828);
or UO_173 (O_173,N_4910,N_4863);
nor UO_174 (O_174,N_4914,N_4944);
or UO_175 (O_175,N_4809,N_4982);
or UO_176 (O_176,N_4860,N_4855);
or UO_177 (O_177,N_4947,N_4926);
nor UO_178 (O_178,N_4832,N_4809);
nand UO_179 (O_179,N_4969,N_4805);
nor UO_180 (O_180,N_4962,N_4995);
or UO_181 (O_181,N_4936,N_4847);
xor UO_182 (O_182,N_4860,N_4850);
nor UO_183 (O_183,N_4992,N_4979);
and UO_184 (O_184,N_4995,N_4946);
nand UO_185 (O_185,N_4885,N_4930);
and UO_186 (O_186,N_4931,N_4982);
and UO_187 (O_187,N_4903,N_4923);
nand UO_188 (O_188,N_4879,N_4968);
and UO_189 (O_189,N_4968,N_4876);
and UO_190 (O_190,N_4902,N_4975);
or UO_191 (O_191,N_4911,N_4881);
or UO_192 (O_192,N_4897,N_4915);
nand UO_193 (O_193,N_4850,N_4858);
xor UO_194 (O_194,N_4962,N_4993);
nor UO_195 (O_195,N_4892,N_4819);
xnor UO_196 (O_196,N_4982,N_4880);
xor UO_197 (O_197,N_4816,N_4823);
xor UO_198 (O_198,N_4966,N_4886);
nor UO_199 (O_199,N_4801,N_4970);
nor UO_200 (O_200,N_4860,N_4889);
nor UO_201 (O_201,N_4853,N_4945);
xor UO_202 (O_202,N_4868,N_4985);
xor UO_203 (O_203,N_4982,N_4974);
nand UO_204 (O_204,N_4879,N_4904);
or UO_205 (O_205,N_4831,N_4931);
or UO_206 (O_206,N_4820,N_4914);
xnor UO_207 (O_207,N_4994,N_4919);
nand UO_208 (O_208,N_4869,N_4802);
nor UO_209 (O_209,N_4805,N_4954);
xnor UO_210 (O_210,N_4891,N_4990);
nand UO_211 (O_211,N_4908,N_4807);
xor UO_212 (O_212,N_4976,N_4824);
nand UO_213 (O_213,N_4948,N_4843);
and UO_214 (O_214,N_4952,N_4909);
and UO_215 (O_215,N_4800,N_4955);
or UO_216 (O_216,N_4959,N_4873);
nor UO_217 (O_217,N_4902,N_4912);
and UO_218 (O_218,N_4933,N_4997);
nand UO_219 (O_219,N_4890,N_4904);
xnor UO_220 (O_220,N_4945,N_4913);
or UO_221 (O_221,N_4903,N_4947);
nand UO_222 (O_222,N_4875,N_4890);
or UO_223 (O_223,N_4875,N_4855);
nor UO_224 (O_224,N_4868,N_4906);
xor UO_225 (O_225,N_4849,N_4875);
or UO_226 (O_226,N_4821,N_4846);
xor UO_227 (O_227,N_4878,N_4862);
xnor UO_228 (O_228,N_4840,N_4903);
nor UO_229 (O_229,N_4905,N_4898);
and UO_230 (O_230,N_4960,N_4968);
or UO_231 (O_231,N_4839,N_4836);
or UO_232 (O_232,N_4827,N_4878);
nor UO_233 (O_233,N_4877,N_4853);
nand UO_234 (O_234,N_4912,N_4857);
xor UO_235 (O_235,N_4912,N_4808);
nand UO_236 (O_236,N_4817,N_4806);
or UO_237 (O_237,N_4883,N_4903);
nand UO_238 (O_238,N_4852,N_4893);
nand UO_239 (O_239,N_4895,N_4927);
nand UO_240 (O_240,N_4939,N_4878);
and UO_241 (O_241,N_4950,N_4870);
and UO_242 (O_242,N_4904,N_4867);
and UO_243 (O_243,N_4897,N_4847);
nor UO_244 (O_244,N_4937,N_4944);
nor UO_245 (O_245,N_4860,N_4939);
nor UO_246 (O_246,N_4827,N_4856);
or UO_247 (O_247,N_4845,N_4842);
nor UO_248 (O_248,N_4910,N_4868);
and UO_249 (O_249,N_4801,N_4822);
xnor UO_250 (O_250,N_4900,N_4825);
and UO_251 (O_251,N_4856,N_4901);
and UO_252 (O_252,N_4844,N_4930);
xnor UO_253 (O_253,N_4852,N_4907);
nand UO_254 (O_254,N_4878,N_4814);
nor UO_255 (O_255,N_4828,N_4812);
and UO_256 (O_256,N_4905,N_4966);
or UO_257 (O_257,N_4999,N_4948);
and UO_258 (O_258,N_4975,N_4831);
nor UO_259 (O_259,N_4857,N_4861);
or UO_260 (O_260,N_4927,N_4900);
or UO_261 (O_261,N_4986,N_4936);
nor UO_262 (O_262,N_4982,N_4989);
nor UO_263 (O_263,N_4833,N_4896);
nor UO_264 (O_264,N_4841,N_4858);
xnor UO_265 (O_265,N_4895,N_4855);
nor UO_266 (O_266,N_4984,N_4921);
nor UO_267 (O_267,N_4849,N_4837);
and UO_268 (O_268,N_4863,N_4840);
nor UO_269 (O_269,N_4921,N_4958);
and UO_270 (O_270,N_4984,N_4840);
or UO_271 (O_271,N_4960,N_4974);
nand UO_272 (O_272,N_4997,N_4936);
nand UO_273 (O_273,N_4988,N_4951);
or UO_274 (O_274,N_4901,N_4920);
nand UO_275 (O_275,N_4979,N_4827);
and UO_276 (O_276,N_4863,N_4880);
and UO_277 (O_277,N_4891,N_4824);
and UO_278 (O_278,N_4869,N_4888);
and UO_279 (O_279,N_4892,N_4817);
nor UO_280 (O_280,N_4950,N_4905);
xnor UO_281 (O_281,N_4989,N_4862);
or UO_282 (O_282,N_4933,N_4888);
nand UO_283 (O_283,N_4865,N_4966);
or UO_284 (O_284,N_4818,N_4914);
and UO_285 (O_285,N_4878,N_4866);
or UO_286 (O_286,N_4928,N_4829);
nand UO_287 (O_287,N_4850,N_4864);
xor UO_288 (O_288,N_4938,N_4800);
xor UO_289 (O_289,N_4808,N_4965);
nand UO_290 (O_290,N_4853,N_4913);
and UO_291 (O_291,N_4898,N_4994);
and UO_292 (O_292,N_4869,N_4849);
and UO_293 (O_293,N_4809,N_4879);
and UO_294 (O_294,N_4953,N_4962);
nand UO_295 (O_295,N_4964,N_4831);
and UO_296 (O_296,N_4995,N_4862);
nor UO_297 (O_297,N_4973,N_4847);
nor UO_298 (O_298,N_4854,N_4965);
nand UO_299 (O_299,N_4945,N_4965);
nand UO_300 (O_300,N_4897,N_4868);
xor UO_301 (O_301,N_4948,N_4840);
xor UO_302 (O_302,N_4867,N_4937);
or UO_303 (O_303,N_4806,N_4936);
xnor UO_304 (O_304,N_4997,N_4834);
nor UO_305 (O_305,N_4926,N_4837);
and UO_306 (O_306,N_4907,N_4933);
or UO_307 (O_307,N_4828,N_4837);
nor UO_308 (O_308,N_4828,N_4880);
nor UO_309 (O_309,N_4926,N_4943);
xor UO_310 (O_310,N_4845,N_4942);
xnor UO_311 (O_311,N_4934,N_4985);
nor UO_312 (O_312,N_4943,N_4883);
nand UO_313 (O_313,N_4880,N_4916);
nor UO_314 (O_314,N_4981,N_4900);
nor UO_315 (O_315,N_4959,N_4804);
or UO_316 (O_316,N_4950,N_4841);
and UO_317 (O_317,N_4926,N_4928);
or UO_318 (O_318,N_4820,N_4995);
and UO_319 (O_319,N_4883,N_4868);
nand UO_320 (O_320,N_4952,N_4984);
xor UO_321 (O_321,N_4945,N_4878);
xnor UO_322 (O_322,N_4877,N_4830);
or UO_323 (O_323,N_4810,N_4885);
or UO_324 (O_324,N_4840,N_4977);
xor UO_325 (O_325,N_4955,N_4961);
and UO_326 (O_326,N_4946,N_4994);
nand UO_327 (O_327,N_4811,N_4868);
and UO_328 (O_328,N_4957,N_4906);
and UO_329 (O_329,N_4977,N_4835);
xor UO_330 (O_330,N_4895,N_4921);
nor UO_331 (O_331,N_4934,N_4972);
or UO_332 (O_332,N_4819,N_4953);
nand UO_333 (O_333,N_4927,N_4959);
nor UO_334 (O_334,N_4897,N_4935);
nand UO_335 (O_335,N_4945,N_4827);
nand UO_336 (O_336,N_4986,N_4932);
nor UO_337 (O_337,N_4897,N_4953);
or UO_338 (O_338,N_4952,N_4998);
nand UO_339 (O_339,N_4962,N_4969);
nor UO_340 (O_340,N_4867,N_4956);
nand UO_341 (O_341,N_4885,N_4980);
and UO_342 (O_342,N_4826,N_4930);
and UO_343 (O_343,N_4987,N_4967);
nand UO_344 (O_344,N_4859,N_4841);
and UO_345 (O_345,N_4830,N_4800);
nand UO_346 (O_346,N_4927,N_4963);
xnor UO_347 (O_347,N_4862,N_4972);
nand UO_348 (O_348,N_4806,N_4944);
nand UO_349 (O_349,N_4854,N_4971);
xnor UO_350 (O_350,N_4892,N_4834);
or UO_351 (O_351,N_4972,N_4944);
nand UO_352 (O_352,N_4846,N_4921);
nor UO_353 (O_353,N_4906,N_4870);
xnor UO_354 (O_354,N_4890,N_4821);
xor UO_355 (O_355,N_4889,N_4849);
xnor UO_356 (O_356,N_4820,N_4854);
nand UO_357 (O_357,N_4922,N_4955);
nand UO_358 (O_358,N_4933,N_4851);
xor UO_359 (O_359,N_4862,N_4956);
nor UO_360 (O_360,N_4995,N_4948);
xor UO_361 (O_361,N_4910,N_4883);
or UO_362 (O_362,N_4873,N_4855);
and UO_363 (O_363,N_4920,N_4894);
nor UO_364 (O_364,N_4911,N_4922);
or UO_365 (O_365,N_4983,N_4831);
and UO_366 (O_366,N_4950,N_4807);
xor UO_367 (O_367,N_4983,N_4807);
or UO_368 (O_368,N_4824,N_4848);
and UO_369 (O_369,N_4874,N_4811);
and UO_370 (O_370,N_4935,N_4962);
nand UO_371 (O_371,N_4863,N_4812);
xor UO_372 (O_372,N_4810,N_4921);
nand UO_373 (O_373,N_4975,N_4828);
nor UO_374 (O_374,N_4956,N_4925);
or UO_375 (O_375,N_4836,N_4840);
and UO_376 (O_376,N_4976,N_4805);
or UO_377 (O_377,N_4844,N_4805);
xor UO_378 (O_378,N_4904,N_4897);
nand UO_379 (O_379,N_4875,N_4924);
or UO_380 (O_380,N_4842,N_4980);
and UO_381 (O_381,N_4836,N_4977);
nand UO_382 (O_382,N_4823,N_4879);
nand UO_383 (O_383,N_4843,N_4831);
nor UO_384 (O_384,N_4910,N_4822);
nand UO_385 (O_385,N_4967,N_4865);
nor UO_386 (O_386,N_4907,N_4813);
or UO_387 (O_387,N_4960,N_4886);
and UO_388 (O_388,N_4875,N_4884);
nor UO_389 (O_389,N_4962,N_4868);
xnor UO_390 (O_390,N_4919,N_4905);
and UO_391 (O_391,N_4874,N_4966);
nor UO_392 (O_392,N_4925,N_4812);
or UO_393 (O_393,N_4890,N_4813);
or UO_394 (O_394,N_4829,N_4967);
nand UO_395 (O_395,N_4922,N_4944);
xor UO_396 (O_396,N_4983,N_4817);
nand UO_397 (O_397,N_4903,N_4813);
xor UO_398 (O_398,N_4953,N_4883);
and UO_399 (O_399,N_4818,N_4894);
nor UO_400 (O_400,N_4949,N_4884);
and UO_401 (O_401,N_4848,N_4910);
or UO_402 (O_402,N_4916,N_4902);
nor UO_403 (O_403,N_4984,N_4883);
nand UO_404 (O_404,N_4807,N_4947);
nor UO_405 (O_405,N_4930,N_4904);
or UO_406 (O_406,N_4957,N_4893);
nand UO_407 (O_407,N_4866,N_4863);
and UO_408 (O_408,N_4860,N_4911);
and UO_409 (O_409,N_4918,N_4899);
nand UO_410 (O_410,N_4954,N_4993);
nand UO_411 (O_411,N_4908,N_4845);
and UO_412 (O_412,N_4989,N_4851);
xnor UO_413 (O_413,N_4887,N_4925);
or UO_414 (O_414,N_4867,N_4959);
or UO_415 (O_415,N_4983,N_4851);
or UO_416 (O_416,N_4874,N_4873);
nor UO_417 (O_417,N_4991,N_4955);
and UO_418 (O_418,N_4975,N_4804);
nor UO_419 (O_419,N_4997,N_4857);
xnor UO_420 (O_420,N_4817,N_4931);
and UO_421 (O_421,N_4806,N_4973);
nand UO_422 (O_422,N_4806,N_4965);
and UO_423 (O_423,N_4940,N_4919);
nand UO_424 (O_424,N_4880,N_4867);
nor UO_425 (O_425,N_4940,N_4802);
or UO_426 (O_426,N_4815,N_4809);
xor UO_427 (O_427,N_4889,N_4885);
xor UO_428 (O_428,N_4882,N_4897);
nand UO_429 (O_429,N_4975,N_4848);
xnor UO_430 (O_430,N_4847,N_4990);
and UO_431 (O_431,N_4844,N_4967);
xor UO_432 (O_432,N_4828,N_4961);
and UO_433 (O_433,N_4831,N_4926);
nand UO_434 (O_434,N_4805,N_4807);
xnor UO_435 (O_435,N_4929,N_4968);
nand UO_436 (O_436,N_4967,N_4862);
xnor UO_437 (O_437,N_4877,N_4909);
nand UO_438 (O_438,N_4844,N_4952);
and UO_439 (O_439,N_4957,N_4815);
nor UO_440 (O_440,N_4997,N_4958);
and UO_441 (O_441,N_4826,N_4838);
nor UO_442 (O_442,N_4892,N_4810);
xor UO_443 (O_443,N_4850,N_4819);
xor UO_444 (O_444,N_4903,N_4842);
xnor UO_445 (O_445,N_4941,N_4885);
or UO_446 (O_446,N_4896,N_4811);
nor UO_447 (O_447,N_4830,N_4838);
nor UO_448 (O_448,N_4803,N_4914);
and UO_449 (O_449,N_4934,N_4924);
and UO_450 (O_450,N_4950,N_4806);
and UO_451 (O_451,N_4870,N_4912);
or UO_452 (O_452,N_4850,N_4879);
xnor UO_453 (O_453,N_4935,N_4889);
xnor UO_454 (O_454,N_4920,N_4923);
and UO_455 (O_455,N_4845,N_4993);
or UO_456 (O_456,N_4813,N_4909);
nand UO_457 (O_457,N_4817,N_4834);
or UO_458 (O_458,N_4855,N_4828);
nor UO_459 (O_459,N_4919,N_4800);
xnor UO_460 (O_460,N_4861,N_4968);
and UO_461 (O_461,N_4829,N_4832);
and UO_462 (O_462,N_4812,N_4827);
xor UO_463 (O_463,N_4966,N_4912);
nand UO_464 (O_464,N_4913,N_4847);
nand UO_465 (O_465,N_4979,N_4947);
xor UO_466 (O_466,N_4824,N_4905);
or UO_467 (O_467,N_4945,N_4836);
or UO_468 (O_468,N_4866,N_4888);
xnor UO_469 (O_469,N_4966,N_4878);
and UO_470 (O_470,N_4842,N_4994);
nor UO_471 (O_471,N_4853,N_4818);
nand UO_472 (O_472,N_4973,N_4963);
nor UO_473 (O_473,N_4819,N_4806);
or UO_474 (O_474,N_4972,N_4987);
nor UO_475 (O_475,N_4875,N_4912);
xnor UO_476 (O_476,N_4945,N_4944);
xor UO_477 (O_477,N_4942,N_4974);
or UO_478 (O_478,N_4968,N_4822);
nor UO_479 (O_479,N_4885,N_4890);
nand UO_480 (O_480,N_4976,N_4818);
nand UO_481 (O_481,N_4841,N_4992);
nand UO_482 (O_482,N_4803,N_4979);
or UO_483 (O_483,N_4845,N_4945);
xor UO_484 (O_484,N_4979,N_4860);
nand UO_485 (O_485,N_4973,N_4814);
nand UO_486 (O_486,N_4965,N_4819);
nand UO_487 (O_487,N_4851,N_4944);
nand UO_488 (O_488,N_4925,N_4846);
and UO_489 (O_489,N_4850,N_4805);
or UO_490 (O_490,N_4838,N_4874);
or UO_491 (O_491,N_4931,N_4966);
nor UO_492 (O_492,N_4992,N_4950);
or UO_493 (O_493,N_4998,N_4884);
nor UO_494 (O_494,N_4865,N_4921);
xnor UO_495 (O_495,N_4915,N_4956);
or UO_496 (O_496,N_4824,N_4959);
xnor UO_497 (O_497,N_4844,N_4881);
xnor UO_498 (O_498,N_4901,N_4982);
xor UO_499 (O_499,N_4923,N_4998);
nand UO_500 (O_500,N_4823,N_4825);
nand UO_501 (O_501,N_4874,N_4900);
or UO_502 (O_502,N_4829,N_4930);
xor UO_503 (O_503,N_4943,N_4971);
or UO_504 (O_504,N_4842,N_4993);
xnor UO_505 (O_505,N_4908,N_4935);
and UO_506 (O_506,N_4888,N_4959);
and UO_507 (O_507,N_4842,N_4861);
and UO_508 (O_508,N_4986,N_4962);
and UO_509 (O_509,N_4852,N_4805);
nor UO_510 (O_510,N_4900,N_4963);
xnor UO_511 (O_511,N_4875,N_4992);
nand UO_512 (O_512,N_4933,N_4893);
and UO_513 (O_513,N_4909,N_4942);
or UO_514 (O_514,N_4812,N_4829);
and UO_515 (O_515,N_4855,N_4885);
nor UO_516 (O_516,N_4874,N_4967);
xnor UO_517 (O_517,N_4941,N_4988);
nor UO_518 (O_518,N_4971,N_4998);
nor UO_519 (O_519,N_4958,N_4845);
or UO_520 (O_520,N_4895,N_4904);
xor UO_521 (O_521,N_4994,N_4819);
xor UO_522 (O_522,N_4886,N_4836);
xnor UO_523 (O_523,N_4819,N_4949);
and UO_524 (O_524,N_4872,N_4802);
and UO_525 (O_525,N_4865,N_4859);
nor UO_526 (O_526,N_4951,N_4878);
or UO_527 (O_527,N_4886,N_4972);
nor UO_528 (O_528,N_4952,N_4866);
nand UO_529 (O_529,N_4808,N_4966);
nand UO_530 (O_530,N_4944,N_4916);
xnor UO_531 (O_531,N_4892,N_4927);
nor UO_532 (O_532,N_4807,N_4848);
or UO_533 (O_533,N_4953,N_4899);
nor UO_534 (O_534,N_4966,N_4930);
xor UO_535 (O_535,N_4977,N_4903);
and UO_536 (O_536,N_4801,N_4998);
xor UO_537 (O_537,N_4971,N_4886);
or UO_538 (O_538,N_4876,N_4938);
or UO_539 (O_539,N_4977,N_4961);
or UO_540 (O_540,N_4810,N_4919);
or UO_541 (O_541,N_4825,N_4859);
nor UO_542 (O_542,N_4954,N_4879);
xor UO_543 (O_543,N_4946,N_4925);
and UO_544 (O_544,N_4931,N_4951);
xnor UO_545 (O_545,N_4970,N_4919);
nor UO_546 (O_546,N_4966,N_4827);
and UO_547 (O_547,N_4900,N_4929);
xnor UO_548 (O_548,N_4978,N_4914);
xor UO_549 (O_549,N_4869,N_4975);
nand UO_550 (O_550,N_4884,N_4984);
or UO_551 (O_551,N_4972,N_4993);
or UO_552 (O_552,N_4805,N_4829);
or UO_553 (O_553,N_4978,N_4951);
xnor UO_554 (O_554,N_4829,N_4858);
or UO_555 (O_555,N_4918,N_4910);
nor UO_556 (O_556,N_4942,N_4875);
xnor UO_557 (O_557,N_4879,N_4949);
xnor UO_558 (O_558,N_4951,N_4831);
or UO_559 (O_559,N_4861,N_4902);
or UO_560 (O_560,N_4941,N_4985);
nand UO_561 (O_561,N_4912,N_4953);
or UO_562 (O_562,N_4960,N_4946);
and UO_563 (O_563,N_4984,N_4801);
xor UO_564 (O_564,N_4956,N_4812);
xnor UO_565 (O_565,N_4812,N_4848);
nor UO_566 (O_566,N_4866,N_4873);
nor UO_567 (O_567,N_4944,N_4992);
and UO_568 (O_568,N_4847,N_4930);
nor UO_569 (O_569,N_4819,N_4832);
xor UO_570 (O_570,N_4818,N_4936);
or UO_571 (O_571,N_4958,N_4941);
and UO_572 (O_572,N_4942,N_4865);
nor UO_573 (O_573,N_4850,N_4892);
or UO_574 (O_574,N_4863,N_4813);
nor UO_575 (O_575,N_4840,N_4822);
nor UO_576 (O_576,N_4902,N_4810);
and UO_577 (O_577,N_4936,N_4932);
nand UO_578 (O_578,N_4813,N_4947);
and UO_579 (O_579,N_4860,N_4899);
nor UO_580 (O_580,N_4864,N_4941);
xor UO_581 (O_581,N_4884,N_4809);
nand UO_582 (O_582,N_4874,N_4879);
or UO_583 (O_583,N_4874,N_4819);
xor UO_584 (O_584,N_4807,N_4882);
nor UO_585 (O_585,N_4828,N_4983);
nand UO_586 (O_586,N_4896,N_4804);
and UO_587 (O_587,N_4850,N_4970);
and UO_588 (O_588,N_4950,N_4909);
nand UO_589 (O_589,N_4832,N_4818);
nor UO_590 (O_590,N_4943,N_4860);
nand UO_591 (O_591,N_4862,N_4854);
nor UO_592 (O_592,N_4971,N_4890);
or UO_593 (O_593,N_4838,N_4926);
xor UO_594 (O_594,N_4999,N_4832);
xnor UO_595 (O_595,N_4890,N_4882);
or UO_596 (O_596,N_4995,N_4917);
and UO_597 (O_597,N_4962,N_4978);
and UO_598 (O_598,N_4900,N_4950);
or UO_599 (O_599,N_4968,N_4974);
and UO_600 (O_600,N_4841,N_4866);
and UO_601 (O_601,N_4857,N_4844);
nand UO_602 (O_602,N_4848,N_4998);
nand UO_603 (O_603,N_4946,N_4836);
or UO_604 (O_604,N_4851,N_4959);
nor UO_605 (O_605,N_4902,N_4841);
or UO_606 (O_606,N_4814,N_4889);
nand UO_607 (O_607,N_4816,N_4931);
and UO_608 (O_608,N_4883,N_4860);
and UO_609 (O_609,N_4963,N_4866);
xnor UO_610 (O_610,N_4861,N_4868);
or UO_611 (O_611,N_4890,N_4841);
nor UO_612 (O_612,N_4855,N_4979);
and UO_613 (O_613,N_4972,N_4872);
nand UO_614 (O_614,N_4935,N_4818);
xnor UO_615 (O_615,N_4937,N_4884);
xor UO_616 (O_616,N_4957,N_4853);
xor UO_617 (O_617,N_4900,N_4980);
nor UO_618 (O_618,N_4961,N_4844);
nand UO_619 (O_619,N_4918,N_4892);
and UO_620 (O_620,N_4858,N_4999);
or UO_621 (O_621,N_4940,N_4999);
and UO_622 (O_622,N_4887,N_4986);
xor UO_623 (O_623,N_4848,N_4999);
xnor UO_624 (O_624,N_4928,N_4856);
and UO_625 (O_625,N_4991,N_4903);
nand UO_626 (O_626,N_4826,N_4955);
nor UO_627 (O_627,N_4816,N_4999);
xnor UO_628 (O_628,N_4861,N_4954);
and UO_629 (O_629,N_4967,N_4935);
and UO_630 (O_630,N_4972,N_4940);
nand UO_631 (O_631,N_4901,N_4824);
nand UO_632 (O_632,N_4823,N_4871);
and UO_633 (O_633,N_4910,N_4838);
nor UO_634 (O_634,N_4923,N_4984);
nor UO_635 (O_635,N_4984,N_4857);
or UO_636 (O_636,N_4821,N_4926);
or UO_637 (O_637,N_4994,N_4972);
or UO_638 (O_638,N_4922,N_4903);
nand UO_639 (O_639,N_4981,N_4936);
nor UO_640 (O_640,N_4966,N_4805);
xnor UO_641 (O_641,N_4933,N_4966);
nor UO_642 (O_642,N_4869,N_4989);
xor UO_643 (O_643,N_4941,N_4952);
and UO_644 (O_644,N_4970,N_4909);
nor UO_645 (O_645,N_4944,N_4907);
nor UO_646 (O_646,N_4954,N_4963);
nor UO_647 (O_647,N_4986,N_4806);
nand UO_648 (O_648,N_4926,N_4935);
xnor UO_649 (O_649,N_4820,N_4940);
nand UO_650 (O_650,N_4964,N_4839);
xor UO_651 (O_651,N_4881,N_4842);
and UO_652 (O_652,N_4878,N_4996);
nor UO_653 (O_653,N_4986,N_4839);
and UO_654 (O_654,N_4876,N_4958);
xnor UO_655 (O_655,N_4945,N_4962);
xnor UO_656 (O_656,N_4939,N_4926);
nand UO_657 (O_657,N_4849,N_4844);
or UO_658 (O_658,N_4992,N_4820);
xor UO_659 (O_659,N_4963,N_4875);
nor UO_660 (O_660,N_4803,N_4813);
and UO_661 (O_661,N_4958,N_4916);
nand UO_662 (O_662,N_4825,N_4916);
xor UO_663 (O_663,N_4852,N_4850);
xor UO_664 (O_664,N_4971,N_4825);
or UO_665 (O_665,N_4901,N_4993);
nand UO_666 (O_666,N_4924,N_4807);
xnor UO_667 (O_667,N_4841,N_4993);
or UO_668 (O_668,N_4983,N_4909);
and UO_669 (O_669,N_4918,N_4975);
nand UO_670 (O_670,N_4958,N_4934);
xor UO_671 (O_671,N_4897,N_4971);
xor UO_672 (O_672,N_4876,N_4854);
nand UO_673 (O_673,N_4825,N_4944);
xnor UO_674 (O_674,N_4851,N_4814);
xor UO_675 (O_675,N_4985,N_4959);
nand UO_676 (O_676,N_4810,N_4991);
nand UO_677 (O_677,N_4960,N_4954);
or UO_678 (O_678,N_4831,N_4969);
nand UO_679 (O_679,N_4946,N_4919);
and UO_680 (O_680,N_4978,N_4873);
nor UO_681 (O_681,N_4852,N_4815);
nand UO_682 (O_682,N_4858,N_4846);
nor UO_683 (O_683,N_4867,N_4825);
and UO_684 (O_684,N_4952,N_4883);
and UO_685 (O_685,N_4886,N_4976);
or UO_686 (O_686,N_4874,N_4961);
nand UO_687 (O_687,N_4888,N_4825);
xnor UO_688 (O_688,N_4949,N_4839);
and UO_689 (O_689,N_4841,N_4967);
and UO_690 (O_690,N_4855,N_4812);
and UO_691 (O_691,N_4898,N_4980);
or UO_692 (O_692,N_4823,N_4947);
nor UO_693 (O_693,N_4965,N_4823);
nor UO_694 (O_694,N_4951,N_4887);
nand UO_695 (O_695,N_4939,N_4995);
or UO_696 (O_696,N_4889,N_4856);
nor UO_697 (O_697,N_4941,N_4882);
xnor UO_698 (O_698,N_4851,N_4856);
and UO_699 (O_699,N_4957,N_4995);
nand UO_700 (O_700,N_4962,N_4835);
xnor UO_701 (O_701,N_4863,N_4991);
and UO_702 (O_702,N_4999,N_4991);
or UO_703 (O_703,N_4927,N_4809);
xor UO_704 (O_704,N_4814,N_4884);
xor UO_705 (O_705,N_4937,N_4900);
and UO_706 (O_706,N_4903,N_4907);
nor UO_707 (O_707,N_4828,N_4931);
and UO_708 (O_708,N_4866,N_4883);
and UO_709 (O_709,N_4965,N_4839);
and UO_710 (O_710,N_4915,N_4875);
nor UO_711 (O_711,N_4963,N_4956);
or UO_712 (O_712,N_4880,N_4829);
xnor UO_713 (O_713,N_4889,N_4922);
and UO_714 (O_714,N_4986,N_4935);
xor UO_715 (O_715,N_4985,N_4966);
nor UO_716 (O_716,N_4820,N_4839);
or UO_717 (O_717,N_4851,N_4889);
xnor UO_718 (O_718,N_4950,N_4813);
nor UO_719 (O_719,N_4854,N_4996);
xor UO_720 (O_720,N_4815,N_4807);
xor UO_721 (O_721,N_4810,N_4949);
and UO_722 (O_722,N_4845,N_4935);
or UO_723 (O_723,N_4905,N_4817);
nand UO_724 (O_724,N_4993,N_4959);
nor UO_725 (O_725,N_4965,N_4835);
xnor UO_726 (O_726,N_4918,N_4999);
and UO_727 (O_727,N_4951,N_4835);
xnor UO_728 (O_728,N_4895,N_4858);
nor UO_729 (O_729,N_4994,N_4993);
and UO_730 (O_730,N_4852,N_4934);
xnor UO_731 (O_731,N_4890,N_4999);
nand UO_732 (O_732,N_4937,N_4852);
and UO_733 (O_733,N_4917,N_4964);
or UO_734 (O_734,N_4806,N_4994);
and UO_735 (O_735,N_4917,N_4825);
or UO_736 (O_736,N_4859,N_4889);
nand UO_737 (O_737,N_4987,N_4934);
xor UO_738 (O_738,N_4917,N_4860);
xor UO_739 (O_739,N_4845,N_4994);
and UO_740 (O_740,N_4879,N_4963);
nor UO_741 (O_741,N_4924,N_4981);
nand UO_742 (O_742,N_4866,N_4874);
and UO_743 (O_743,N_4802,N_4873);
nor UO_744 (O_744,N_4865,N_4896);
nor UO_745 (O_745,N_4991,N_4933);
or UO_746 (O_746,N_4938,N_4851);
or UO_747 (O_747,N_4902,N_4936);
nor UO_748 (O_748,N_4847,N_4832);
and UO_749 (O_749,N_4887,N_4863);
xor UO_750 (O_750,N_4943,N_4831);
xor UO_751 (O_751,N_4876,N_4845);
or UO_752 (O_752,N_4865,N_4960);
xor UO_753 (O_753,N_4891,N_4884);
or UO_754 (O_754,N_4863,N_4921);
and UO_755 (O_755,N_4866,N_4815);
xnor UO_756 (O_756,N_4840,N_4922);
nand UO_757 (O_757,N_4825,N_4810);
xnor UO_758 (O_758,N_4818,N_4890);
and UO_759 (O_759,N_4974,N_4804);
nand UO_760 (O_760,N_4940,N_4969);
and UO_761 (O_761,N_4901,N_4927);
nor UO_762 (O_762,N_4922,N_4954);
or UO_763 (O_763,N_4861,N_4865);
or UO_764 (O_764,N_4800,N_4869);
or UO_765 (O_765,N_4940,N_4987);
and UO_766 (O_766,N_4867,N_4967);
nand UO_767 (O_767,N_4873,N_4875);
xnor UO_768 (O_768,N_4923,N_4993);
and UO_769 (O_769,N_4972,N_4966);
or UO_770 (O_770,N_4854,N_4938);
nand UO_771 (O_771,N_4806,N_4913);
nor UO_772 (O_772,N_4990,N_4878);
nand UO_773 (O_773,N_4980,N_4930);
xor UO_774 (O_774,N_4845,N_4964);
nand UO_775 (O_775,N_4804,N_4867);
nand UO_776 (O_776,N_4852,N_4857);
xnor UO_777 (O_777,N_4978,N_4801);
and UO_778 (O_778,N_4826,N_4921);
nor UO_779 (O_779,N_4996,N_4896);
or UO_780 (O_780,N_4966,N_4862);
nor UO_781 (O_781,N_4956,N_4822);
nand UO_782 (O_782,N_4875,N_4935);
or UO_783 (O_783,N_4914,N_4869);
or UO_784 (O_784,N_4919,N_4852);
or UO_785 (O_785,N_4918,N_4813);
xnor UO_786 (O_786,N_4816,N_4807);
nand UO_787 (O_787,N_4957,N_4962);
nand UO_788 (O_788,N_4946,N_4865);
nand UO_789 (O_789,N_4805,N_4864);
nand UO_790 (O_790,N_4851,N_4982);
nand UO_791 (O_791,N_4850,N_4853);
and UO_792 (O_792,N_4919,N_4969);
xnor UO_793 (O_793,N_4813,N_4821);
nor UO_794 (O_794,N_4885,N_4946);
xor UO_795 (O_795,N_4894,N_4947);
xnor UO_796 (O_796,N_4803,N_4962);
xnor UO_797 (O_797,N_4896,N_4840);
and UO_798 (O_798,N_4998,N_4897);
nor UO_799 (O_799,N_4899,N_4948);
and UO_800 (O_800,N_4916,N_4864);
nor UO_801 (O_801,N_4964,N_4899);
xnor UO_802 (O_802,N_4964,N_4924);
nor UO_803 (O_803,N_4906,N_4954);
and UO_804 (O_804,N_4906,N_4815);
or UO_805 (O_805,N_4922,N_4937);
nand UO_806 (O_806,N_4980,N_4838);
nand UO_807 (O_807,N_4945,N_4830);
nor UO_808 (O_808,N_4882,N_4852);
and UO_809 (O_809,N_4996,N_4966);
or UO_810 (O_810,N_4882,N_4999);
nand UO_811 (O_811,N_4945,N_4849);
xnor UO_812 (O_812,N_4997,N_4967);
xor UO_813 (O_813,N_4893,N_4953);
nand UO_814 (O_814,N_4995,N_4965);
or UO_815 (O_815,N_4895,N_4899);
nor UO_816 (O_816,N_4885,N_4839);
nand UO_817 (O_817,N_4865,N_4816);
nor UO_818 (O_818,N_4849,N_4973);
nand UO_819 (O_819,N_4901,N_4839);
xor UO_820 (O_820,N_4966,N_4887);
xnor UO_821 (O_821,N_4975,N_4865);
or UO_822 (O_822,N_4976,N_4897);
and UO_823 (O_823,N_4858,N_4940);
and UO_824 (O_824,N_4864,N_4869);
and UO_825 (O_825,N_4999,N_4814);
and UO_826 (O_826,N_4912,N_4929);
nand UO_827 (O_827,N_4912,N_4919);
and UO_828 (O_828,N_4945,N_4907);
nand UO_829 (O_829,N_4840,N_4912);
nor UO_830 (O_830,N_4923,N_4828);
nand UO_831 (O_831,N_4987,N_4894);
and UO_832 (O_832,N_4908,N_4974);
nand UO_833 (O_833,N_4886,N_4890);
xnor UO_834 (O_834,N_4808,N_4992);
and UO_835 (O_835,N_4925,N_4931);
and UO_836 (O_836,N_4947,N_4887);
or UO_837 (O_837,N_4933,N_4842);
or UO_838 (O_838,N_4822,N_4852);
nor UO_839 (O_839,N_4902,N_4914);
nand UO_840 (O_840,N_4911,N_4912);
nor UO_841 (O_841,N_4983,N_4907);
xnor UO_842 (O_842,N_4853,N_4992);
nand UO_843 (O_843,N_4953,N_4886);
nor UO_844 (O_844,N_4868,N_4976);
or UO_845 (O_845,N_4984,N_4998);
nand UO_846 (O_846,N_4954,N_4885);
and UO_847 (O_847,N_4973,N_4953);
xnor UO_848 (O_848,N_4803,N_4985);
nor UO_849 (O_849,N_4821,N_4928);
nand UO_850 (O_850,N_4960,N_4874);
xnor UO_851 (O_851,N_4806,N_4873);
nor UO_852 (O_852,N_4959,N_4839);
or UO_853 (O_853,N_4901,N_4847);
and UO_854 (O_854,N_4845,N_4978);
and UO_855 (O_855,N_4822,N_4951);
nor UO_856 (O_856,N_4920,N_4839);
nor UO_857 (O_857,N_4854,N_4856);
xor UO_858 (O_858,N_4921,N_4989);
nor UO_859 (O_859,N_4882,N_4952);
xor UO_860 (O_860,N_4876,N_4872);
or UO_861 (O_861,N_4865,N_4927);
xnor UO_862 (O_862,N_4873,N_4971);
nand UO_863 (O_863,N_4827,N_4865);
or UO_864 (O_864,N_4988,N_4998);
or UO_865 (O_865,N_4888,N_4938);
xor UO_866 (O_866,N_4994,N_4951);
xnor UO_867 (O_867,N_4928,N_4937);
or UO_868 (O_868,N_4830,N_4964);
nor UO_869 (O_869,N_4800,N_4953);
and UO_870 (O_870,N_4949,N_4844);
and UO_871 (O_871,N_4908,N_4814);
nand UO_872 (O_872,N_4850,N_4876);
xor UO_873 (O_873,N_4850,N_4901);
nor UO_874 (O_874,N_4942,N_4880);
nand UO_875 (O_875,N_4878,N_4976);
nand UO_876 (O_876,N_4901,N_4916);
or UO_877 (O_877,N_4964,N_4968);
nand UO_878 (O_878,N_4870,N_4822);
nand UO_879 (O_879,N_4994,N_4945);
and UO_880 (O_880,N_4872,N_4848);
xor UO_881 (O_881,N_4892,N_4881);
nand UO_882 (O_882,N_4958,N_4863);
xor UO_883 (O_883,N_4974,N_4957);
and UO_884 (O_884,N_4984,N_4802);
xor UO_885 (O_885,N_4877,N_4858);
or UO_886 (O_886,N_4973,N_4976);
nand UO_887 (O_887,N_4853,N_4912);
xor UO_888 (O_888,N_4807,N_4951);
xnor UO_889 (O_889,N_4964,N_4986);
or UO_890 (O_890,N_4832,N_4869);
and UO_891 (O_891,N_4969,N_4844);
nor UO_892 (O_892,N_4824,N_4803);
nand UO_893 (O_893,N_4922,N_4849);
nor UO_894 (O_894,N_4879,N_4984);
and UO_895 (O_895,N_4889,N_4983);
xor UO_896 (O_896,N_4989,N_4868);
nand UO_897 (O_897,N_4941,N_4948);
and UO_898 (O_898,N_4986,N_4912);
nor UO_899 (O_899,N_4899,N_4988);
or UO_900 (O_900,N_4845,N_4921);
xor UO_901 (O_901,N_4963,N_4849);
nor UO_902 (O_902,N_4847,N_4831);
or UO_903 (O_903,N_4945,N_4938);
and UO_904 (O_904,N_4855,N_4844);
and UO_905 (O_905,N_4838,N_4973);
nor UO_906 (O_906,N_4829,N_4915);
nand UO_907 (O_907,N_4817,N_4826);
xor UO_908 (O_908,N_4929,N_4896);
xor UO_909 (O_909,N_4988,N_4985);
or UO_910 (O_910,N_4977,N_4960);
xor UO_911 (O_911,N_4901,N_4946);
nor UO_912 (O_912,N_4812,N_4817);
nand UO_913 (O_913,N_4855,N_4997);
or UO_914 (O_914,N_4843,N_4860);
nor UO_915 (O_915,N_4997,N_4803);
and UO_916 (O_916,N_4890,N_4957);
nand UO_917 (O_917,N_4989,N_4836);
nand UO_918 (O_918,N_4829,N_4873);
nor UO_919 (O_919,N_4850,N_4932);
nor UO_920 (O_920,N_4984,N_4981);
or UO_921 (O_921,N_4835,N_4909);
nand UO_922 (O_922,N_4882,N_4820);
and UO_923 (O_923,N_4999,N_4973);
nor UO_924 (O_924,N_4844,N_4809);
and UO_925 (O_925,N_4875,N_4967);
and UO_926 (O_926,N_4853,N_4849);
and UO_927 (O_927,N_4806,N_4807);
nor UO_928 (O_928,N_4922,N_4852);
nor UO_929 (O_929,N_4990,N_4830);
nand UO_930 (O_930,N_4979,N_4811);
xor UO_931 (O_931,N_4976,N_4943);
nand UO_932 (O_932,N_4862,N_4818);
nor UO_933 (O_933,N_4892,N_4843);
and UO_934 (O_934,N_4834,N_4879);
nand UO_935 (O_935,N_4983,N_4932);
nor UO_936 (O_936,N_4817,N_4808);
and UO_937 (O_937,N_4990,N_4902);
xor UO_938 (O_938,N_4815,N_4991);
nor UO_939 (O_939,N_4836,N_4847);
or UO_940 (O_940,N_4844,N_4823);
nor UO_941 (O_941,N_4817,N_4908);
or UO_942 (O_942,N_4983,N_4802);
nor UO_943 (O_943,N_4941,N_4812);
or UO_944 (O_944,N_4809,N_4953);
nor UO_945 (O_945,N_4927,N_4857);
nor UO_946 (O_946,N_4936,N_4917);
and UO_947 (O_947,N_4939,N_4958);
xor UO_948 (O_948,N_4836,N_4972);
or UO_949 (O_949,N_4938,N_4998);
nor UO_950 (O_950,N_4912,N_4824);
nor UO_951 (O_951,N_4837,N_4923);
or UO_952 (O_952,N_4845,N_4847);
nand UO_953 (O_953,N_4857,N_4956);
and UO_954 (O_954,N_4919,N_4851);
and UO_955 (O_955,N_4962,N_4845);
or UO_956 (O_956,N_4906,N_4995);
nor UO_957 (O_957,N_4893,N_4994);
nor UO_958 (O_958,N_4817,N_4994);
nand UO_959 (O_959,N_4853,N_4831);
and UO_960 (O_960,N_4918,N_4871);
and UO_961 (O_961,N_4806,N_4939);
or UO_962 (O_962,N_4923,N_4881);
nand UO_963 (O_963,N_4921,N_4858);
or UO_964 (O_964,N_4945,N_4834);
or UO_965 (O_965,N_4985,N_4891);
and UO_966 (O_966,N_4869,N_4857);
and UO_967 (O_967,N_4948,N_4891);
nand UO_968 (O_968,N_4855,N_4849);
xnor UO_969 (O_969,N_4899,N_4929);
nor UO_970 (O_970,N_4868,N_4986);
xnor UO_971 (O_971,N_4997,N_4881);
and UO_972 (O_972,N_4888,N_4941);
or UO_973 (O_973,N_4925,N_4855);
or UO_974 (O_974,N_4816,N_4875);
or UO_975 (O_975,N_4841,N_4878);
and UO_976 (O_976,N_4944,N_4975);
nand UO_977 (O_977,N_4964,N_4842);
nand UO_978 (O_978,N_4840,N_4846);
nand UO_979 (O_979,N_4898,N_4949);
nor UO_980 (O_980,N_4971,N_4962);
and UO_981 (O_981,N_4864,N_4907);
and UO_982 (O_982,N_4922,N_4833);
and UO_983 (O_983,N_4811,N_4968);
nor UO_984 (O_984,N_4940,N_4966);
nor UO_985 (O_985,N_4983,N_4893);
nor UO_986 (O_986,N_4894,N_4831);
nand UO_987 (O_987,N_4928,N_4891);
xnor UO_988 (O_988,N_4817,N_4865);
xnor UO_989 (O_989,N_4886,N_4915);
and UO_990 (O_990,N_4807,N_4969);
and UO_991 (O_991,N_4922,N_4842);
or UO_992 (O_992,N_4818,N_4921);
xor UO_993 (O_993,N_4980,N_4953);
nand UO_994 (O_994,N_4825,N_4966);
xnor UO_995 (O_995,N_4922,N_4885);
or UO_996 (O_996,N_4803,N_4954);
nand UO_997 (O_997,N_4846,N_4968);
and UO_998 (O_998,N_4909,N_4802);
and UO_999 (O_999,N_4863,N_4867);
endmodule